magic
tech sky130A
magscale 1 2
timestamp 1762784779
<< viali >>
rect 2973 42789 3007 42823
rect 3617 42789 3651 42823
rect 7573 42789 7607 42823
rect 7665 42789 7699 42823
rect 8769 42789 8803 42823
rect 1133 42721 1167 42755
rect 1225 42721 1259 42755
rect 1492 42721 1526 42755
rect 4537 42721 4571 42755
rect 5457 42721 5491 42755
rect 5641 42721 5675 42755
rect 7476 42721 7510 42755
rect 7848 42721 7882 42755
rect 7941 42721 7975 42755
rect 8033 42721 8067 42755
rect 8217 42721 8251 42755
rect 8401 42721 8435 42755
rect 8494 42721 8528 42755
rect 8677 42721 8711 42755
rect 8866 42721 8900 42755
rect 9137 42721 9171 42755
rect 10057 42721 10091 42755
rect 10517 42721 10551 42755
rect 11069 42721 11103 42755
rect 11345 42721 11379 42755
rect 11437 42721 11471 42755
rect 11621 42721 11655 42755
rect 12265 42721 12299 42755
rect 4445 42653 4479 42687
rect 4813 42653 4847 42687
rect 6377 42653 6411 42687
rect 7205 42653 7239 42687
rect 9689 42653 9723 42687
rect 10241 42653 10275 42687
rect 10333 42653 10367 42687
rect 11989 42653 12023 42687
rect 3433 42585 3467 42619
rect 11253 42585 11287 42619
rect 949 42517 983 42551
rect 2605 42517 2639 42551
rect 2881 42517 2915 42551
rect 3801 42517 3835 42551
rect 5641 42517 5675 42551
rect 5825 42517 5859 42551
rect 6561 42517 6595 42551
rect 7297 42517 7331 42551
rect 8217 42517 8251 42551
rect 9045 42517 9079 42551
rect 9873 42517 9907 42551
rect 10701 42517 10735 42551
rect 11805 42517 11839 42551
rect 12081 42517 12115 42551
rect 12173 42517 12207 42551
rect 2973 42313 3007 42347
rect 5273 42313 5307 42347
rect 8677 42313 8711 42347
rect 4905 42245 4939 42279
rect 7845 42245 7879 42279
rect 10885 42245 10919 42279
rect 8493 42177 8527 42211
rect 857 42109 891 42143
rect 1005 42109 1039 42143
rect 1133 42109 1167 42143
rect 1363 42109 1397 42143
rect 1593 42109 1627 42143
rect 3433 42109 3467 42143
rect 4077 42109 4111 42143
rect 4170 42109 4204 42143
rect 4353 42109 4387 42143
rect 4445 42109 4479 42143
rect 4542 42109 4576 42143
rect 4813 42109 4847 42143
rect 5089 42109 5123 42143
rect 5365 42109 5399 42143
rect 5632 42109 5666 42143
rect 6929 42109 6963 42143
rect 7665 42109 7699 42143
rect 7757 42109 7791 42143
rect 7941 42109 7975 42143
rect 8585 42109 8619 42143
rect 9137 42109 9171 42143
rect 9321 42109 9355 42143
rect 9505 42109 9539 42143
rect 9689 42109 9723 42143
rect 10149 42109 10183 42143
rect 12265 42109 12299 42143
rect 1225 42041 1259 42075
rect 1860 42041 1894 42075
rect 8861 42041 8895 42075
rect 8953 42041 8987 42075
rect 9045 42041 9079 42075
rect 10425 42041 10459 42075
rect 12020 42041 12054 42075
rect 1501 41973 1535 42007
rect 3985 41973 4019 42007
rect 4721 41973 4755 42007
rect 6745 41973 6779 42007
rect 7481 41973 7515 42007
rect 8125 41973 8159 42007
rect 9873 41973 9907 42007
rect 10057 41973 10091 42007
rect 10517 41973 10551 42007
rect 1225 41769 1259 41803
rect 6101 41769 6135 41803
rect 9229 41769 9263 41803
rect 12081 41769 12115 41803
rect 12265 41769 12299 41803
rect 2145 41701 2179 41735
rect 4506 41701 4540 41735
rect 9045 41701 9079 41735
rect 10548 41701 10582 41735
rect 949 41633 983 41667
rect 1133 41633 1167 41667
rect 2237 41633 2271 41667
rect 2504 41633 2538 41667
rect 3893 41633 3927 41667
rect 4169 41633 4203 41667
rect 5825 41633 5859 41667
rect 6009 41633 6043 41667
rect 8033 41633 8067 41667
rect 8309 41633 8343 41667
rect 8861 41633 8895 41667
rect 11253 41633 11287 41667
rect 11345 41633 11379 41667
rect 11437 41633 11471 41667
rect 11621 41633 11655 41667
rect 1593 41565 1627 41599
rect 4077 41565 4111 41599
rect 4261 41565 4295 41599
rect 6653 41565 6687 41599
rect 10793 41565 10827 41599
rect 11713 41565 11747 41599
rect 1409 41497 1443 41531
rect 3709 41497 3743 41531
rect 3617 41429 3651 41463
rect 5641 41429 5675 41463
rect 5917 41429 5951 41463
rect 9413 41429 9447 41463
rect 10977 41429 11011 41463
rect 12081 41429 12115 41463
rect 11805 41225 11839 41259
rect 7573 41157 7607 41191
rect 8033 41157 8067 41191
rect 8401 41157 8435 41191
rect 857 41089 891 41123
rect 1409 41089 1443 41123
rect 7665 41089 7699 41123
rect 11989 41089 12023 41123
rect 1041 41021 1075 41055
rect 1225 41021 1259 41055
rect 1685 41021 1719 41055
rect 3709 41021 3743 41055
rect 5365 41021 5399 41055
rect 6837 41021 6871 41055
rect 7297 41021 7331 41055
rect 7481 41021 7515 41055
rect 7757 41021 7791 41055
rect 8033 41021 8067 41055
rect 8217 41021 8251 41055
rect 8677 41021 8711 41055
rect 9321 41021 9355 41055
rect 9413 41021 9447 41055
rect 10425 41021 10459 41055
rect 10692 41021 10726 41055
rect 12173 41021 12207 41055
rect 12265 41021 12299 41055
rect 3065 40953 3099 40987
rect 3525 40953 3559 40987
rect 3976 40953 4010 40987
rect 5632 40953 5666 40987
rect 7021 40953 7055 40987
rect 8401 40953 8435 40987
rect 8585 40953 8619 40987
rect 9965 40953 9999 40987
rect 10149 40953 10183 40987
rect 3433 40885 3467 40919
rect 5089 40885 5123 40919
rect 6745 40885 6779 40919
rect 7205 40885 7239 40919
rect 7941 40885 7975 40919
rect 8769 40885 8803 40919
rect 10333 40885 10367 40919
rect 11989 40885 12023 40919
rect 1225 40681 1259 40715
rect 1685 40681 1719 40715
rect 5457 40681 5491 40715
rect 5089 40613 5123 40647
rect 5181 40613 5215 40647
rect 1409 40545 1443 40579
rect 2329 40545 2363 40579
rect 2585 40545 2619 40579
rect 4031 40545 4065 40579
rect 4169 40545 4203 40579
rect 4261 40545 4295 40579
rect 4389 40545 4423 40579
rect 4537 40545 4571 40579
rect 4813 40545 4847 40579
rect 4906 40545 4940 40579
rect 5278 40545 5312 40579
rect 6653 40545 6687 40579
rect 7389 40545 7423 40579
rect 7573 40545 7607 40579
rect 8309 40545 8343 40579
rect 8677 40545 8711 40579
rect 9137 40545 9171 40579
rect 9597 40545 9631 40579
rect 10977 40545 11011 40579
rect 11253 40545 11287 40579
rect 11437 40545 11471 40579
rect 11529 40545 11563 40579
rect 11621 40545 11655 40579
rect 12081 40545 12115 40579
rect 2145 40477 2179 40511
rect 6561 40477 6595 40511
rect 7757 40477 7791 40511
rect 1777 40409 1811 40443
rect 3893 40409 3927 40443
rect 10149 40409 10183 40443
rect 3709 40341 3743 40375
rect 5917 40341 5951 40375
rect 7297 40341 7331 40375
rect 7481 40341 7515 40375
rect 11069 40341 11103 40375
rect 11897 40341 11931 40375
rect 12173 40341 12207 40375
rect 2145 40137 2179 40171
rect 2329 40137 2363 40171
rect 2513 40137 2547 40171
rect 6469 40137 6503 40171
rect 7757 40137 7791 40171
rect 8125 40137 8159 40171
rect 8493 40137 8527 40171
rect 9137 40137 9171 40171
rect 9689 40137 9723 40171
rect 10609 40137 10643 40171
rect 1409 40069 1443 40103
rect 8861 40069 8895 40103
rect 3801 40001 3835 40035
rect 5089 40001 5123 40035
rect 8217 40001 8251 40035
rect 12265 40001 12299 40035
rect 1133 39933 1167 39967
rect 1225 39933 1259 39967
rect 1409 39933 1443 39967
rect 1501 39933 1535 39967
rect 1685 39933 1719 39967
rect 1869 39933 1903 39967
rect 2663 39933 2697 39967
rect 2973 39933 3007 39967
rect 3065 39933 3099 39967
rect 4261 39933 4295 39967
rect 4353 39933 4387 39967
rect 4446 39933 4480 39967
rect 4629 39933 4663 39967
rect 4859 39933 4893 39967
rect 5356 39933 5390 39967
rect 7389 39933 7423 39967
rect 7573 39933 7607 39967
rect 7941 39933 7975 39967
rect 8401 39933 8435 39967
rect 8677 39933 8711 39967
rect 9045 39933 9079 39967
rect 9229 39933 9263 39967
rect 1961 39865 1995 39899
rect 3709 39865 3743 39899
rect 4721 39865 4755 39899
rect 9505 39865 9539 39899
rect 10149 39865 10183 39899
rect 10425 39865 10459 39899
rect 11998 39865 12032 39899
rect 949 39797 983 39831
rect 2171 39797 2205 39831
rect 3249 39797 3283 39831
rect 3617 39797 3651 39831
rect 4169 39797 4203 39831
rect 4997 39797 5031 39831
rect 6561 39797 6595 39831
rect 9705 39797 9739 39831
rect 9873 39797 9907 39831
rect 10057 39797 10091 39831
rect 10625 39797 10659 39831
rect 10793 39797 10827 39831
rect 10885 39797 10919 39831
rect 3709 39593 3743 39627
rect 2574 39525 2608 39559
rect 11437 39525 11471 39559
rect 1133 39457 1167 39491
rect 1593 39457 1627 39491
rect 1869 39457 1903 39491
rect 2053 39457 2087 39491
rect 2329 39457 2363 39491
rect 4077 39457 4111 39491
rect 5641 39457 5675 39491
rect 6561 39457 6595 39491
rect 8493 39457 8527 39491
rect 9075 39457 9109 39491
rect 9229 39457 9263 39491
rect 9321 39457 9355 39491
rect 9588 39457 9622 39491
rect 11713 39457 11747 39491
rect 11989 39457 12023 39491
rect 2145 39389 2179 39423
rect 4169 39389 4203 39423
rect 5917 39389 5951 39423
rect 7113 39389 7147 39423
rect 7849 39389 7883 39423
rect 8217 39389 8251 39423
rect 8677 39389 8711 39423
rect 11529 39389 11563 39423
rect 1409 39321 1443 39355
rect 4997 39321 5031 39355
rect 6469 39321 6503 39355
rect 8861 39321 8895 39355
rect 10701 39321 10735 39355
rect 11161 39321 11195 39355
rect 11897 39321 11931 39355
rect 949 39253 983 39287
rect 1685 39253 1719 39287
rect 3893 39253 3927 39287
rect 4813 39253 4847 39287
rect 6745 39253 6779 39287
rect 8309 39253 8343 39287
rect 10977 39253 11011 39287
rect 12173 39253 12207 39287
rect 3065 39049 3099 39083
rect 9965 39049 9999 39083
rect 10517 39049 10551 39083
rect 3893 38981 3927 39015
rect 7205 38981 7239 39015
rect 7481 38981 7515 39015
rect 8125 38981 8159 39015
rect 8769 38981 8803 39015
rect 9597 38981 9631 39015
rect 1593 38913 1627 38947
rect 3341 38913 3375 38947
rect 8401 38913 8435 38947
rect 8677 38913 8711 38947
rect 10793 38913 10827 38947
rect 1133 38845 1167 38879
rect 1225 38845 1259 38879
rect 1409 38845 1443 38879
rect 1685 38845 1719 38879
rect 3617 38845 3651 38879
rect 5825 38845 5859 38879
rect 7297 38845 7331 38879
rect 7941 38845 7975 38879
rect 8585 38845 8619 38879
rect 8861 38845 8895 38879
rect 9413 38845 9447 38879
rect 10090 38845 10124 38879
rect 10609 38845 10643 38879
rect 1952 38777 1986 38811
rect 4169 38777 4203 38811
rect 5733 38777 5767 38811
rect 6092 38777 6126 38811
rect 9045 38777 9079 38811
rect 11060 38777 11094 38811
rect 949 38709 983 38743
rect 3525 38709 3559 38743
rect 3709 38709 3743 38743
rect 7849 38709 7883 38743
rect 9229 38709 9263 38743
rect 9321 38709 9355 38743
rect 10149 38709 10183 38743
rect 12173 38709 12207 38743
rect 5181 38505 5215 38539
rect 7205 38505 7239 38539
rect 8401 38505 8435 38539
rect 11345 38505 11379 38539
rect 6070 38437 6104 38471
rect 10425 38437 10459 38471
rect 10625 38437 10659 38471
rect 10977 38437 11011 38471
rect 11989 38437 12023 38471
rect 1409 38369 1443 38403
rect 1593 38369 1627 38403
rect 2053 38369 2087 38403
rect 2309 38369 2343 38403
rect 3525 38369 3559 38403
rect 3709 38369 3743 38403
rect 3801 38369 3835 38403
rect 4068 38369 4102 38403
rect 5457 38369 5491 38403
rect 5549 38369 5583 38403
rect 5825 38369 5859 38403
rect 8217 38369 8251 38403
rect 9045 38369 9079 38403
rect 9321 38369 9355 38403
rect 9597 38369 9631 38403
rect 9781 38369 9815 38403
rect 10149 38369 10183 38403
rect 11161 38369 11195 38403
rect 11253 38369 11287 38403
rect 11805 38369 11839 38403
rect 12081 38369 12115 38403
rect 12265 38369 12299 38403
rect 949 38301 983 38335
rect 1685 38301 1719 38335
rect 5273 38301 5307 38335
rect 7297 38301 7331 38335
rect 8033 38301 8067 38335
rect 8769 38301 8803 38335
rect 9413 38301 9447 38335
rect 11621 38301 11655 38335
rect 3433 38233 3467 38267
rect 8493 38233 8527 38267
rect 9137 38233 9171 38267
rect 9505 38233 9539 38267
rect 11529 38233 11563 38267
rect 3617 38165 3651 38199
rect 7941 38165 7975 38199
rect 8677 38165 8711 38199
rect 9873 38165 9907 38199
rect 10333 38165 10367 38199
rect 10609 38165 10643 38199
rect 10793 38165 10827 38199
rect 12173 38165 12207 38199
rect 4813 37961 4847 37995
rect 5549 37961 5583 37995
rect 6377 37961 6411 37995
rect 9321 37961 9355 37995
rect 3249 37893 3283 37927
rect 5641 37893 5675 37927
rect 8677 37893 8711 37927
rect 2605 37825 2639 37859
rect 3065 37825 3099 37859
rect 3893 37825 3927 37859
rect 857 37757 891 37791
rect 2697 37757 2731 37791
rect 4169 37757 4203 37791
rect 4262 37757 4296 37791
rect 4675 37757 4709 37791
rect 4997 37757 5031 37791
rect 6285 37757 6319 37791
rect 7757 37757 7791 37791
rect 8033 37757 8067 37791
rect 8217 37757 8251 37791
rect 8401 37757 8435 37791
rect 8585 37757 8619 37791
rect 8769 37757 8803 37791
rect 8861 37757 8895 37791
rect 9137 37757 9171 37791
rect 9597 37757 9631 37791
rect 11805 37757 11839 37791
rect 11897 37757 11931 37791
rect 11989 37757 12023 37791
rect 1124 37689 1158 37723
rect 4445 37689 4479 37723
rect 4537 37689 4571 37723
rect 7490 37689 7524 37723
rect 2237 37621 2271 37655
rect 3617 37621 3651 37655
rect 3709 37621 3743 37655
rect 7849 37621 7883 37655
rect 9045 37621 9079 37655
rect 12173 37621 12207 37655
rect 949 37417 983 37451
rect 5825 37417 5859 37451
rect 7205 37417 7239 37451
rect 7573 37417 7607 37451
rect 8861 37417 8895 37451
rect 10333 37417 10367 37451
rect 12173 37417 12207 37451
rect 4261 37349 4295 37383
rect 7665 37349 7699 37383
rect 11437 37349 11471 37383
rect 11897 37349 11931 37383
rect 1041 37281 1075 37315
rect 1133 37281 1167 37315
rect 1225 37281 1259 37315
rect 1409 37281 1443 37315
rect 1685 37281 1719 37315
rect 1941 37281 1975 37315
rect 3525 37281 3559 37315
rect 3617 37281 3651 37315
rect 3801 37281 3835 37315
rect 4537 37281 4571 37315
rect 5089 37281 5123 37315
rect 5273 37281 5307 37315
rect 5549 37281 5583 37315
rect 6469 37281 6503 37315
rect 6929 37281 6963 37315
rect 8217 37281 8251 37315
rect 8309 37281 8343 37315
rect 8677 37281 8711 37315
rect 8769 37281 8803 37315
rect 8953 37281 8987 37315
rect 9045 37281 9079 37315
rect 11161 37281 11195 37315
rect 11529 37281 11563 37315
rect 11713 37281 11747 37315
rect 11989 37281 12023 37315
rect 4629 37213 4663 37247
rect 4905 37213 4939 37247
rect 5365 37213 5399 37247
rect 7021 37213 7055 37247
rect 7849 37213 7883 37247
rect 11253 37213 11287 37247
rect 1593 37145 1627 37179
rect 5457 37145 5491 37179
rect 6561 37145 6595 37179
rect 3065 37077 3099 37111
rect 8033 37077 8067 37111
rect 8217 37077 8251 37111
rect 10977 37077 11011 37111
rect 11161 37077 11195 37111
rect 3249 36873 3283 36907
rect 7297 36873 7331 36907
rect 8217 36873 8251 36907
rect 8769 36873 8803 36907
rect 6929 36805 6963 36839
rect 7757 36805 7791 36839
rect 9413 36805 9447 36839
rect 1409 36737 1443 36771
rect 6009 36737 6043 36771
rect 7205 36737 7239 36771
rect 8125 36737 8159 36771
rect 9045 36737 9079 36771
rect 9229 36737 9263 36771
rect 10333 36737 10367 36771
rect 10885 36737 10919 36771
rect 1317 36669 1351 36703
rect 1685 36669 1719 36703
rect 4629 36669 4663 36703
rect 4721 36669 4755 36703
rect 5365 36669 5399 36703
rect 5733 36669 5767 36703
rect 5917 36669 5951 36703
rect 7297 36669 7331 36703
rect 7481 36669 7515 36703
rect 7941 36669 7975 36703
rect 8217 36669 8251 36703
rect 8392 36647 8426 36681
rect 8493 36669 8527 36703
rect 8949 36669 8983 36703
rect 9137 36669 9171 36703
rect 9413 36669 9447 36703
rect 9689 36669 9723 36703
rect 10241 36669 10275 36703
rect 10793 36669 10827 36703
rect 3065 36601 3099 36635
rect 4384 36601 4418 36635
rect 5181 36601 5215 36635
rect 8677 36601 8711 36635
rect 11152 36601 11186 36635
rect 1133 36533 1167 36567
rect 5917 36533 5951 36567
rect 6653 36533 6687 36567
rect 6745 36533 6779 36567
rect 7665 36533 7699 36567
rect 8578 36533 8612 36567
rect 9597 36533 9631 36567
rect 9781 36533 9815 36567
rect 10149 36533 10183 36567
rect 10701 36533 10735 36567
rect 12265 36533 12299 36567
rect 5825 36329 5859 36363
rect 6285 36329 6319 36363
rect 7573 36329 7607 36363
rect 8585 36329 8619 36363
rect 10977 36329 11011 36363
rect 11713 36329 11747 36363
rect 4528 36261 4562 36295
rect 7481 36261 7515 36295
rect 8125 36261 8159 36295
rect 9137 36261 9171 36295
rect 1133 36193 1167 36227
rect 1317 36193 1351 36227
rect 1593 36193 1627 36227
rect 3801 36193 3835 36227
rect 4261 36193 4295 36227
rect 6193 36193 6227 36227
rect 6653 36193 6687 36227
rect 6837 36193 6871 36227
rect 6929 36193 6963 36227
rect 7113 36193 7147 36227
rect 7757 36193 7791 36227
rect 8401 36193 8435 36227
rect 8861 36193 8895 36227
rect 9781 36193 9815 36227
rect 9873 36193 9907 36227
rect 10425 36193 10459 36227
rect 11161 36193 11195 36227
rect 11253 36193 11287 36227
rect 11345 36193 11379 36227
rect 11463 36193 11497 36227
rect 11897 36193 11931 36227
rect 11989 36193 12023 36227
rect 6377 36125 6411 36159
rect 8033 36125 8067 36159
rect 8309 36125 8343 36159
rect 9045 36125 9079 36159
rect 9589 36125 9623 36159
rect 9689 36125 9723 36159
rect 10333 36125 10367 36159
rect 10793 36125 10827 36159
rect 11621 36125 11655 36159
rect 1501 36057 1535 36091
rect 7297 36057 7331 36091
rect 8677 36057 8711 36091
rect 949 35989 983 36023
rect 3985 35989 4019 36023
rect 5641 35989 5675 36023
rect 6745 35989 6779 36023
rect 7941 35989 7975 36023
rect 8401 35989 8435 36023
rect 8861 35989 8895 36023
rect 9413 35989 9447 36023
rect 949 35785 983 35819
rect 1593 35785 1627 35819
rect 5825 35785 5859 35819
rect 7757 35785 7791 35819
rect 9505 35785 9539 35819
rect 9689 35785 9723 35819
rect 10241 35785 10275 35819
rect 10425 35785 10459 35819
rect 5733 35717 5767 35751
rect 7481 35717 7515 35751
rect 9321 35717 9355 35751
rect 10149 35717 10183 35751
rect 10885 35717 10919 35751
rect 3709 35649 3743 35683
rect 3893 35649 3927 35683
rect 4353 35649 4387 35683
rect 6837 35649 6871 35683
rect 7113 35649 7147 35683
rect 8953 35649 8987 35683
rect 9781 35649 9815 35683
rect 10517 35649 10551 35683
rect 4077 35581 4111 35615
rect 4261 35581 4295 35615
rect 6009 35581 6043 35615
rect 6101 35581 6135 35615
rect 6193 35581 6227 35615
rect 6469 35581 6503 35615
rect 6745 35581 6779 35615
rect 7941 35581 7975 35615
rect 9137 35581 9171 35615
rect 9413 35581 9447 35615
rect 9689 35581 9723 35615
rect 9965 35581 9999 35615
rect 10425 35581 10459 35615
rect 12265 35581 12299 35615
rect 3065 35513 3099 35547
rect 4620 35513 4654 35547
rect 6331 35513 6365 35547
rect 7297 35513 7331 35547
rect 8125 35513 8159 35547
rect 8401 35513 8435 35547
rect 8585 35513 8619 35547
rect 10701 35513 10735 35547
rect 11998 35513 12032 35547
rect 3249 35445 3283 35479
rect 3617 35445 3651 35479
rect 4261 35445 4295 35479
rect 949 35241 983 35275
rect 2237 35241 2271 35275
rect 3709 35241 3743 35275
rect 4077 35241 4111 35275
rect 4537 35241 4571 35275
rect 6009 35241 6043 35275
rect 6653 35241 6687 35275
rect 3350 35173 3384 35207
rect 5273 35173 5307 35207
rect 7665 35173 7699 35207
rect 9137 35173 9171 35207
rect 12049 35173 12083 35207
rect 12265 35173 12299 35207
rect 1041 35105 1075 35139
rect 1133 35105 1167 35139
rect 1593 35105 1627 35139
rect 1777 35105 1811 35139
rect 3617 35105 3651 35139
rect 4721 35105 4755 35139
rect 4997 35105 5031 35139
rect 5181 35105 5215 35139
rect 5457 35105 5491 35139
rect 5549 35105 5583 35139
rect 5825 35105 5859 35139
rect 6009 35105 6043 35139
rect 6101 35105 6135 35139
rect 6837 35105 6871 35139
rect 7021 35105 7055 35139
rect 7113 35105 7147 35139
rect 7481 35105 7515 35139
rect 7849 35105 7883 35139
rect 8493 35105 8527 35139
rect 8769 35105 8803 35139
rect 8953 35105 8987 35139
rect 9505 35105 9539 35139
rect 9597 35105 9631 35139
rect 10241 35105 10275 35139
rect 11161 35105 11195 35139
rect 11253 35105 11287 35139
rect 11437 35105 11471 35139
rect 11621 35105 11655 35139
rect 1869 35037 1903 35071
rect 4169 35037 4203 35071
rect 4261 35037 4295 35071
rect 6377 35037 6411 35071
rect 7205 35037 7239 35071
rect 8309 35037 8343 35071
rect 9689 35037 9723 35071
rect 9781 35037 9815 35071
rect 10149 35037 10183 35071
rect 10609 34969 10643 35003
rect 11805 34969 11839 35003
rect 5273 34901 5307 34935
rect 7297 34901 7331 34935
rect 7941 34901 7975 34935
rect 8677 34901 8711 34935
rect 9965 34901 9999 34935
rect 10977 34901 11011 34935
rect 11897 34901 11931 34935
rect 12081 34901 12115 34935
rect 949 34697 983 34731
rect 4537 34697 4571 34731
rect 5825 34697 5859 34731
rect 6745 34697 6779 34731
rect 8861 34697 8895 34731
rect 2513 34629 2547 34663
rect 6929 34629 6963 34663
rect 10425 34629 10459 34663
rect 10517 34629 10551 34663
rect 2973 34561 3007 34595
rect 3801 34561 3835 34595
rect 4997 34561 5031 34595
rect 5181 34561 5215 34595
rect 5457 34561 5491 34595
rect 2329 34493 2363 34527
rect 2881 34493 2915 34527
rect 4169 34493 4203 34527
rect 5089 34493 5123 34527
rect 5273 34493 5307 34527
rect 6377 34493 6411 34527
rect 6469 34493 6503 34527
rect 6561 34493 6595 34527
rect 6837 34493 6871 34527
rect 7021 34493 7055 34527
rect 7389 34493 7423 34527
rect 7665 34493 7699 34527
rect 8217 34493 8251 34527
rect 8585 34493 8619 34527
rect 8677 34493 8711 34527
rect 8953 34493 8987 34527
rect 9045 34493 9079 34527
rect 10517 34493 10551 34527
rect 10701 34493 10735 34527
rect 11998 34493 12032 34527
rect 12265 34493 12299 34527
rect 2062 34425 2096 34459
rect 4537 34425 4571 34459
rect 5825 34425 5859 34459
rect 9312 34425 9346 34459
rect 3249 34357 3283 34391
rect 3617 34357 3651 34391
rect 3709 34357 3743 34391
rect 4721 34357 4755 34391
rect 4813 34357 4847 34391
rect 6009 34357 6043 34391
rect 8401 34357 8435 34391
rect 10885 34357 10919 34391
rect 949 34153 983 34187
rect 3617 34153 3651 34187
rect 11437 34153 11471 34187
rect 1133 34085 1167 34119
rect 2504 34085 2538 34119
rect 3801 34085 3835 34119
rect 11897 34085 11931 34119
rect 4031 34051 4065 34085
rect 1041 34017 1075 34051
rect 1593 34017 1627 34051
rect 1777 34017 1811 34051
rect 2237 34017 2271 34051
rect 4261 34017 4295 34051
rect 4528 34017 4562 34051
rect 6009 34017 6043 34051
rect 6265 34017 6299 34051
rect 7481 34017 7515 34051
rect 7665 34017 7699 34051
rect 8125 34017 8159 34051
rect 8401 34017 8435 34051
rect 9321 34017 9355 34051
rect 9597 34017 9631 34051
rect 9689 34017 9723 34051
rect 9781 34017 9815 34051
rect 9873 34017 9907 34051
rect 10069 34039 10103 34073
rect 11667 34051 11701 34085
rect 10333 34017 10367 34051
rect 10425 34017 10459 34051
rect 11253 34017 11287 34051
rect 12173 34017 12207 34051
rect 1869 33949 1903 33983
rect 7849 33949 7883 33983
rect 10517 33949 10551 33983
rect 10609 33949 10643 33983
rect 10977 33949 11011 33983
rect 9413 33881 9447 33915
rect 10149 33881 10183 33915
rect 11069 33881 11103 33915
rect 11529 33881 11563 33915
rect 3985 33813 4019 33847
rect 4169 33813 4203 33847
rect 5641 33813 5675 33847
rect 7389 33813 7423 33847
rect 7573 33813 7607 33847
rect 9137 33813 9171 33847
rect 11713 33813 11747 33847
rect 12081 33813 12115 33847
rect 857 33609 891 33643
rect 3617 33609 3651 33643
rect 6377 33609 6411 33643
rect 11897 33609 11931 33643
rect 5181 33541 5215 33575
rect 7481 33541 7515 33575
rect 8217 33541 8251 33575
rect 11989 33541 12023 33575
rect 2237 33473 2271 33507
rect 2513 33473 2547 33507
rect 3433 33473 3467 33507
rect 3801 33473 3835 33507
rect 5457 33473 5491 33507
rect 5733 33473 5767 33507
rect 2697 33405 2731 33439
rect 3709 33405 3743 33439
rect 4068 33405 4102 33439
rect 6561 33405 6595 33439
rect 6745 33405 6779 33439
rect 6837 33405 6871 33439
rect 7297 33405 7331 33439
rect 7481 33405 7515 33439
rect 7941 33405 7975 33439
rect 9514 33405 9548 33439
rect 9781 33405 9815 33439
rect 10517 33405 10551 33439
rect 10784 33405 10818 33439
rect 12265 33405 12299 33439
rect 1970 33337 2004 33371
rect 6929 33337 6963 33371
rect 7113 33337 7147 33371
rect 7757 33337 7791 33371
rect 8217 33337 8251 33371
rect 9965 33337 9999 33371
rect 10333 33337 10367 33371
rect 11989 33337 12023 33371
rect 2605 33269 2639 33303
rect 3065 33269 3099 33303
rect 3433 33269 3467 33303
rect 7665 33269 7699 33303
rect 8033 33269 8067 33303
rect 8401 33269 8435 33303
rect 12173 33269 12207 33303
rect 4169 33065 4203 33099
rect 4905 33065 4939 33099
rect 6745 33065 6779 33099
rect 7297 33065 7331 33099
rect 8033 33065 8067 33099
rect 8493 33065 8527 33099
rect 11069 33065 11103 33099
rect 1133 32997 1167 33031
rect 2964 32997 2998 33031
rect 5549 32997 5583 33031
rect 857 32929 891 32963
rect 2349 32929 2383 32963
rect 2605 32929 2639 32963
rect 4905 32929 4939 32963
rect 5089 32929 5123 32963
rect 5365 32929 5399 32963
rect 5825 32929 5859 32963
rect 5963 32929 5997 32963
rect 6285 32929 6319 32963
rect 6653 32929 6687 32963
rect 6837 32929 6871 32963
rect 7021 32929 7055 32963
rect 7205 32929 7239 32963
rect 7389 32929 7423 32963
rect 7481 32929 7515 32963
rect 7573 32929 7607 32963
rect 7941 32929 7975 32963
rect 8125 32929 8159 32963
rect 8217 32929 8251 32963
rect 8677 32929 8711 32963
rect 9137 32929 9171 32963
rect 9321 32929 9355 32963
rect 10537 32929 10571 32963
rect 10793 32929 10827 32963
rect 11253 32929 11287 32963
rect 11713 32929 11747 32963
rect 1133 32861 1167 32895
rect 2697 32861 2731 32895
rect 4813 32861 4847 32895
rect 5181 32861 5215 32895
rect 8493 32861 8527 32895
rect 11437 32861 11471 32895
rect 12265 32861 12299 32895
rect 949 32793 983 32827
rect 6193 32793 6227 32827
rect 6469 32793 6503 32827
rect 8309 32793 8343 32827
rect 1225 32725 1259 32759
rect 4077 32725 4111 32759
rect 6101 32725 6135 32759
rect 7757 32725 7791 32759
rect 8953 32725 8987 32759
rect 9229 32725 9263 32759
rect 9413 32725 9447 32759
rect 3249 32521 3283 32555
rect 5917 32521 5951 32555
rect 6653 32521 6687 32555
rect 6745 32521 6779 32555
rect 6929 32521 6963 32555
rect 9229 32521 9263 32555
rect 9505 32521 9539 32555
rect 10333 32521 10367 32555
rect 1501 32453 1535 32487
rect 4077 32453 4111 32487
rect 5181 32453 5215 32487
rect 5273 32453 5307 32487
rect 7205 32453 7239 32487
rect 8677 32453 8711 32487
rect 8861 32453 8895 32487
rect 9413 32453 9447 32487
rect 6009 32385 6043 32419
rect 6377 32385 6411 32419
rect 6469 32385 6503 32419
rect 7849 32385 7883 32419
rect 8033 32385 8067 32419
rect 8125 32385 8159 32419
rect 9781 32385 9815 32419
rect 9873 32385 9907 32419
rect 9965 32385 9999 32419
rect 949 32317 983 32351
rect 1225 32317 1259 32351
rect 2697 32317 2731 32351
rect 2973 32317 3007 32351
rect 3433 32317 3467 32351
rect 3525 32317 3559 32351
rect 3893 32317 3927 32351
rect 4353 32317 4387 32351
rect 4445 32317 4479 32351
rect 4629 32317 4663 32351
rect 4813 32317 4847 32351
rect 5089 32317 5123 32351
rect 5365 32317 5399 32351
rect 6101 32317 6135 32351
rect 7389 32317 7423 32351
rect 7573 32317 7607 32351
rect 7941 32317 7975 32351
rect 8493 32317 8527 32351
rect 9689 32317 9723 32351
rect 10149 32317 10183 32351
rect 10517 32317 10551 32351
rect 12265 32317 12299 32351
rect 1777 32249 1811 32283
rect 2237 32249 2271 32283
rect 2605 32249 2639 32283
rect 5549 32249 5583 32283
rect 5733 32249 5767 32283
rect 7113 32249 7147 32283
rect 9229 32249 9263 32283
rect 1041 32181 1075 32215
rect 1685 32181 1719 32215
rect 4169 32181 4203 32215
rect 4721 32181 4755 32215
rect 4905 32181 4939 32215
rect 6285 32181 6319 32215
rect 6913 32181 6947 32215
rect 7665 32181 7699 32215
rect 6009 31977 6043 32011
rect 8033 31977 8067 32011
rect 949 31909 983 31943
rect 2329 31909 2363 31943
rect 3525 31909 3559 31943
rect 4905 31909 4939 31943
rect 6561 31909 6595 31943
rect 8861 31909 8895 31943
rect 1409 31841 1443 31875
rect 1593 31841 1627 31875
rect 2053 31841 2087 31875
rect 2237 31841 2271 31875
rect 2605 31841 2639 31875
rect 2881 31841 2915 31875
rect 3709 31841 3743 31875
rect 4261 31841 4295 31875
rect 4537 31841 4571 31875
rect 5089 31841 5123 31875
rect 5181 31841 5215 31875
rect 5457 31841 5491 31875
rect 5549 31841 5583 31875
rect 5825 31841 5859 31875
rect 6285 31841 6319 31875
rect 6653 31841 6687 31875
rect 7021 31841 7055 31875
rect 7389 31841 7423 31875
rect 7481 31841 7515 31875
rect 7757 31841 7791 31875
rect 7849 31841 7883 31875
rect 8033 31841 8067 31875
rect 8309 31841 8343 31875
rect 8493 31841 8527 31875
rect 8585 31841 8619 31875
rect 8769 31831 8803 31865
rect 9045 31841 9079 31875
rect 9321 31841 9355 31875
rect 9577 31841 9611 31875
rect 10977 31841 11011 31875
rect 11161 31841 11195 31875
rect 11713 31841 11747 31875
rect 12081 31841 12115 31875
rect 1685 31773 1719 31807
rect 3249 31773 3283 31807
rect 3985 31773 4019 31807
rect 5365 31773 5399 31807
rect 6377 31773 6411 31807
rect 11897 31773 11931 31807
rect 12265 31773 12299 31807
rect 6101 31705 6135 31739
rect 8401 31705 8435 31739
rect 2237 31637 2271 31671
rect 3893 31637 3927 31671
rect 4077 31637 4111 31671
rect 4445 31637 4479 31671
rect 6561 31637 6595 31671
rect 7205 31637 7239 31671
rect 7665 31637 7699 31671
rect 8125 31637 8159 31671
rect 9229 31637 9263 31671
rect 10701 31637 10735 31671
rect 11161 31637 11195 31671
rect 857 31433 891 31467
rect 3433 31433 3467 31467
rect 5457 31433 5491 31467
rect 6101 31433 6135 31467
rect 10425 31433 10459 31467
rect 2421 31365 2455 31399
rect 5181 31365 5215 31399
rect 3249 31297 3283 31331
rect 10885 31297 10919 31331
rect 1970 31229 2004 31263
rect 2237 31229 2271 31263
rect 2697 31229 2731 31263
rect 2789 31229 2823 31263
rect 3709 31229 3743 31263
rect 3801 31229 3835 31263
rect 4068 31229 4102 31263
rect 5641 31229 5675 31263
rect 5733 31229 5767 31263
rect 5917 31229 5951 31263
rect 6009 31207 6043 31241
rect 6377 31229 6411 31263
rect 6469 31229 6503 31263
rect 6561 31229 6595 31263
rect 6653 31229 6687 31263
rect 6837 31229 6871 31263
rect 7113 31229 7147 31263
rect 7297 31229 7331 31263
rect 7389 31229 7423 31263
rect 7481 31229 7515 31263
rect 8033 31229 8067 31263
rect 8401 31229 8435 31263
rect 9045 31229 9079 31263
rect 10517 31229 10551 31263
rect 11152 31229 11186 31263
rect 2421 31161 2455 31195
rect 2605 31161 2639 31195
rect 2973 31161 3007 31195
rect 8217 31161 8251 31195
rect 8677 31161 8711 31195
rect 9312 31161 9346 31195
rect 3617 31093 3651 31127
rect 7757 31093 7791 31127
rect 7849 31093 7883 31127
rect 10701 31093 10735 31127
rect 12265 31093 12299 31127
rect 5089 30889 5123 30923
rect 5917 30889 5951 30923
rect 6745 30889 6779 30923
rect 6837 30889 6871 30923
rect 8953 30889 8987 30923
rect 9597 30889 9631 30923
rect 11069 30889 11103 30923
rect 11897 30889 11931 30923
rect 3976 30821 4010 30855
rect 7297 30821 7331 30855
rect 9229 30821 9263 30855
rect 9321 30821 9355 30855
rect 9749 30821 9783 30855
rect 9965 30821 9999 30855
rect 10425 30821 10459 30855
rect 1970 30753 2004 30787
rect 2329 30753 2363 30787
rect 2513 30753 2547 30787
rect 2789 30753 2823 30787
rect 3249 30753 3283 30787
rect 3525 30753 3559 30787
rect 5365 30753 5399 30787
rect 5641 30753 5675 30787
rect 6101 30753 6135 30787
rect 6469 30753 6503 30787
rect 6561 30753 6595 30787
rect 7021 30753 7055 30787
rect 7481 30753 7515 30787
rect 7665 30753 7699 30787
rect 7849 30753 7883 30787
rect 8125 30753 8159 30787
rect 8217 30753 8251 30787
rect 9137 30753 9171 30787
rect 9505 30753 9539 30787
rect 10057 30753 10091 30787
rect 10150 30753 10184 30787
rect 10793 30753 10827 30787
rect 11253 30753 11287 30787
rect 11805 30753 11839 30787
rect 12173 30753 12207 30787
rect 2237 30685 2271 30719
rect 3709 30685 3743 30719
rect 5549 30685 5583 30719
rect 7205 30685 7239 30719
rect 8585 30685 8619 30719
rect 10517 30685 10551 30719
rect 10701 30685 10735 30719
rect 11437 30685 11471 30719
rect 11897 30685 11931 30719
rect 12081 30617 12115 30651
rect 857 30549 891 30583
rect 2697 30549 2731 30583
rect 3065 30549 3099 30583
rect 3433 30549 3467 30583
rect 5181 30549 5215 30583
rect 5549 30549 5583 30583
rect 6193 30549 6227 30583
rect 7021 30549 7055 30583
rect 9781 30549 9815 30583
rect 10609 30549 10643 30583
rect 11621 30549 11655 30583
rect 2053 30345 2087 30379
rect 2881 30345 2915 30379
rect 5457 30345 5491 30379
rect 5917 30345 5951 30379
rect 6193 30345 6227 30379
rect 6745 30345 6779 30379
rect 7113 30345 7147 30379
rect 7481 30345 7515 30379
rect 10885 30345 10919 30379
rect 7665 30277 7699 30311
rect 8769 30277 8803 30311
rect 9689 30277 9723 30311
rect 10241 30277 10275 30311
rect 10701 30277 10735 30311
rect 2697 30209 2731 30243
rect 3617 30209 3651 30243
rect 9413 30209 9447 30243
rect 10517 30209 10551 30243
rect 12265 30209 12299 30243
rect 1225 30141 1259 30175
rect 1317 30141 1351 30175
rect 1501 30141 1535 30175
rect 2237 30141 2271 30175
rect 2421 30141 2455 30175
rect 2513 30141 2547 30175
rect 2973 30141 3007 30175
rect 3433 30141 3467 30175
rect 3525 30141 3559 30175
rect 3709 30141 3743 30175
rect 3893 30141 3927 30175
rect 4261 30141 4295 30175
rect 4629 30141 4663 30175
rect 5181 30141 5215 30175
rect 5641 30141 5675 30175
rect 5825 30141 5859 30175
rect 6009 30141 6043 30175
rect 6101 30141 6135 30175
rect 6285 30141 6319 30175
rect 6561 30141 6595 30175
rect 7113 30141 7147 30175
rect 7297 30141 7331 30175
rect 7573 30141 7607 30175
rect 7757 30141 7791 30175
rect 8125 30141 8159 30175
rect 8401 30141 8435 30175
rect 8861 30141 8895 30175
rect 8953 30141 8987 30175
rect 9045 30141 9079 30175
rect 9321 30141 9355 30175
rect 9781 30141 9815 30175
rect 10333 30141 10367 30175
rect 10793 30141 10827 30175
rect 1961 30073 1995 30107
rect 2697 30073 2731 30107
rect 6377 30073 6411 30107
rect 8585 30073 8619 30107
rect 11998 30073 12032 30107
rect 3249 30005 3283 30039
rect 4077 30005 4111 30039
rect 4445 30005 4479 30039
rect 4813 30005 4847 30039
rect 5089 30005 5123 30039
rect 7941 30005 7975 30039
rect 9965 30005 9999 30039
rect 10517 30005 10551 30039
rect 1041 29801 1075 29835
rect 1501 29801 1535 29835
rect 1777 29801 1811 29835
rect 2966 29801 3000 29835
rect 3433 29801 3467 29835
rect 3617 29801 3651 29835
rect 4997 29801 5031 29835
rect 6837 29801 6871 29835
rect 8033 29801 8067 29835
rect 10057 29801 10091 29835
rect 10241 29801 10275 29835
rect 10977 29801 11011 29835
rect 11881 29801 11915 29835
rect 1685 29733 1719 29767
rect 3068 29733 3102 29767
rect 6653 29733 6687 29767
rect 10701 29733 10735 29767
rect 12081 29733 12115 29767
rect 1225 29665 1259 29699
rect 1409 29665 1443 29699
rect 1961 29665 1995 29699
rect 2421 29665 2455 29699
rect 2605 29665 2639 29699
rect 2789 29665 2823 29699
rect 2881 29665 2915 29699
rect 3157 29665 3191 29699
rect 3709 29665 3743 29699
rect 3801 29665 3835 29699
rect 3893 29665 3927 29699
rect 4261 29665 4295 29699
rect 4721 29665 4755 29699
rect 4905 29665 4939 29699
rect 5273 29665 5307 29699
rect 5457 29665 5491 29699
rect 5825 29665 5859 29699
rect 5963 29665 5997 29699
rect 7021 29665 7055 29699
rect 7665 29665 7699 29699
rect 7849 29665 7883 29699
rect 9045 29665 9079 29699
rect 9229 29665 9263 29699
rect 10149 29665 10183 29699
rect 10333 29665 10367 29699
rect 10609 29665 10643 29699
rect 10793 29665 10827 29699
rect 11621 29665 11655 29699
rect 2145 29597 2179 29631
rect 2237 29597 2271 29631
rect 2697 29597 2731 29631
rect 3433 29597 3467 29631
rect 4077 29597 4111 29631
rect 7205 29597 7239 29631
rect 1685 29529 1719 29563
rect 3801 29529 3835 29563
rect 6193 29529 6227 29563
rect 3249 29461 3283 29495
rect 4353 29461 4387 29495
rect 4721 29461 4755 29495
rect 5365 29461 5399 29495
rect 6561 29461 6595 29495
rect 7665 29461 7699 29495
rect 11713 29461 11747 29495
rect 11897 29461 11931 29495
rect 2329 29257 2363 29291
rect 2973 29257 3007 29291
rect 4537 29257 4571 29291
rect 10425 29257 10459 29291
rect 11069 29257 11103 29291
rect 11437 29257 11471 29291
rect 11529 29257 11563 29291
rect 11897 29257 11931 29291
rect 7757 29189 7791 29223
rect 9965 29189 9999 29223
rect 1777 29121 1811 29155
rect 4813 29121 4847 29155
rect 5825 29121 5859 29155
rect 8585 29121 8619 29155
rect 9505 29121 9539 29155
rect 9873 29121 9907 29155
rect 10793 29121 10827 29155
rect 11805 29121 11839 29155
rect 11989 29121 12023 29155
rect 1501 29053 1535 29087
rect 1685 29053 1719 29087
rect 2513 29053 2547 29087
rect 2789 29053 2823 29087
rect 2881 29053 2915 29087
rect 3065 29053 3099 29087
rect 3525 29053 3559 29087
rect 3709 29053 3743 29087
rect 4445 29053 4479 29087
rect 5273 29053 5307 29087
rect 5365 29053 5399 29087
rect 6101 29053 6135 29087
rect 6745 29053 6779 29087
rect 8217 29053 8251 29087
rect 8769 29053 8803 29087
rect 9413 29053 9447 29087
rect 10333 29053 10367 29087
rect 10425 29053 10459 29087
rect 10609 29053 10643 29087
rect 10701 29053 10735 29087
rect 10977 29053 11011 29087
rect 11161 29053 11195 29087
rect 11253 29053 11287 29087
rect 11437 29053 11471 29087
rect 11529 29053 11563 29087
rect 11713 29053 11747 29087
rect 12081 29053 12115 29087
rect 1041 28985 1075 29019
rect 2697 28985 2731 29019
rect 4905 28985 4939 29019
rect 6009 28985 6043 29019
rect 6469 28985 6503 29019
rect 6837 28985 6871 29019
rect 7205 28985 7239 29019
rect 3341 28917 3375 28951
rect 7573 28917 7607 28951
rect 8125 28917 8159 28951
rect 8677 28917 8711 28951
rect 9137 28917 9171 28951
rect 9781 28917 9815 28951
rect 3433 28713 3467 28747
rect 4261 28713 4295 28747
rect 5365 28713 5399 28747
rect 8677 28713 8711 28747
rect 9781 28713 9815 28747
rect 12173 28713 12207 28747
rect 2329 28645 2363 28679
rect 4537 28645 4571 28679
rect 6193 28645 6227 28679
rect 8861 28645 8895 28679
rect 10057 28645 10091 28679
rect 10609 28645 10643 28679
rect 11897 28645 11931 28679
rect 1113 28577 1147 28611
rect 2789 28577 2823 28611
rect 2973 28577 3007 28611
rect 3617 28577 3651 28611
rect 3801 28577 3835 28611
rect 3893 28577 3927 28611
rect 4629 28577 4663 28611
rect 4997 28577 5031 28611
rect 5917 28577 5951 28611
rect 6837 28577 6871 28611
rect 7205 28577 7239 28611
rect 7665 28577 7699 28611
rect 7941 28577 7975 28611
rect 8125 28577 8159 28611
rect 8217 28577 8251 28611
rect 8493 28577 8527 28611
rect 9137 28577 9171 28611
rect 9321 28577 9355 28611
rect 9597 28577 9631 28611
rect 9873 28577 9907 28611
rect 10425 28577 10459 28611
rect 10793 28577 10827 28611
rect 10977 28577 11011 28611
rect 11161 28577 11195 28611
rect 11253 28577 11287 28611
rect 11437 28577 11471 28611
rect 11529 28577 11563 28611
rect 11713 28577 11747 28611
rect 11805 28577 11839 28611
rect 12081 28577 12115 28611
rect 12265 28577 12299 28611
rect 857 28509 891 28543
rect 3065 28509 3099 28543
rect 7757 28509 7791 28543
rect 2237 28441 2271 28475
rect 7481 28441 7515 28475
rect 7849 28441 7883 28475
rect 8309 28441 8343 28475
rect 10241 28441 10275 28475
rect 5549 28373 5583 28407
rect 6009 28373 6043 28407
rect 8953 28373 8987 28407
rect 9137 28373 9171 28407
rect 9413 28373 9447 28407
rect 11069 28373 11103 28407
rect 11345 28373 11379 28407
rect 11621 28373 11655 28407
rect 857 28169 891 28203
rect 2605 28169 2639 28203
rect 4445 28169 4479 28203
rect 6193 28169 6227 28203
rect 7205 28169 7239 28203
rect 7941 28169 7975 28203
rect 9229 28169 9263 28203
rect 2237 28033 2271 28067
rect 3525 28033 3559 28067
rect 6653 28033 6687 28067
rect 6745 28033 6779 28067
rect 10057 28033 10091 28067
rect 10333 28033 10367 28067
rect 10977 28033 11011 28067
rect 11437 28033 11471 28067
rect 2789 27965 2823 27999
rect 2973 27965 3007 27999
rect 3065 27965 3099 27999
rect 3985 27965 4019 27999
rect 4261 27965 4295 27999
rect 4445 27965 4479 27999
rect 5457 27965 5491 27999
rect 6561 27965 6595 27999
rect 7021 27965 7055 27999
rect 7205 27965 7239 27999
rect 7481 27965 7515 27999
rect 7665 27965 7699 27999
rect 7757 27965 7791 27999
rect 8953 27965 8987 27999
rect 9045 27965 9079 27999
rect 9321 27965 9355 27999
rect 9597 27965 9631 27999
rect 9873 27965 9907 27999
rect 9965 27965 9999 27999
rect 10149 27965 10183 27999
rect 10425 27965 10459 27999
rect 10885 27965 10919 27999
rect 11069 27965 11103 27999
rect 11345 27965 11379 27999
rect 11805 27965 11839 27999
rect 11897 27965 11931 27999
rect 12081 27965 12115 27999
rect 1970 27897 2004 27931
rect 3893 27897 3927 27931
rect 4997 27897 5031 27931
rect 5089 27897 5123 27931
rect 8033 27897 8067 27931
rect 8401 27897 8435 27931
rect 8585 27897 8619 27931
rect 9413 27897 9447 27931
rect 3801 27829 3835 27863
rect 4721 27829 4755 27863
rect 5825 27829 5859 27863
rect 6009 27829 6043 27863
rect 7297 27829 7331 27863
rect 8769 27829 8803 27863
rect 9781 27829 9815 27863
rect 10793 27829 10827 27863
rect 11713 27829 11747 27863
rect 12265 27829 12299 27863
rect 3617 27625 3651 27659
rect 8125 27625 8159 27659
rect 8585 27625 8619 27659
rect 11069 27625 11103 27659
rect 2145 27557 2179 27591
rect 3249 27557 3283 27591
rect 8493 27557 8527 27591
rect 9873 27557 9907 27591
rect 11989 27557 12023 27591
rect 1317 27489 1351 27523
rect 1501 27489 1535 27523
rect 1777 27489 1811 27523
rect 2053 27489 2087 27523
rect 2329 27489 2363 27523
rect 2513 27489 2547 27523
rect 2605 27489 2639 27523
rect 2881 27489 2915 27523
rect 3065 27489 3099 27523
rect 3157 27489 3191 27523
rect 3433 27489 3467 27523
rect 3709 27489 3743 27523
rect 4353 27489 4387 27523
rect 4537 27489 4571 27523
rect 5089 27489 5123 27523
rect 5181 27489 5215 27523
rect 5365 27489 5399 27523
rect 6101 27489 6135 27523
rect 6837 27489 6871 27523
rect 7021 27489 7055 27523
rect 7389 27489 7423 27523
rect 8033 27489 8067 27523
rect 9321 27489 9355 27523
rect 9413 27489 9447 27523
rect 9597 27489 9631 27523
rect 9689 27489 9723 27523
rect 10517 27489 10551 27523
rect 10701 27489 10735 27523
rect 10793 27489 10827 27523
rect 10977 27489 11011 27523
rect 11161 27489 11195 27523
rect 11437 27489 11471 27523
rect 11897 27489 11931 27523
rect 12081 27489 12115 27523
rect 7205 27421 7239 27455
rect 7481 27421 7515 27455
rect 7573 27421 7607 27455
rect 7665 27421 7699 27455
rect 8677 27421 8711 27455
rect 10333 27421 10367 27455
rect 11529 27421 11563 27455
rect 1961 27353 1995 27387
rect 2697 27353 2731 27387
rect 4721 27353 4755 27387
rect 4905 27353 4939 27387
rect 5273 27353 5307 27387
rect 9137 27353 9171 27387
rect 1133 27285 1167 27319
rect 1593 27285 1627 27319
rect 6193 27285 6227 27319
rect 6929 27285 6963 27319
rect 7941 27285 7975 27319
rect 9965 27285 9999 27319
rect 11713 27285 11747 27319
rect 4629 27081 4663 27115
rect 7757 27081 7791 27115
rect 9229 27081 9263 27115
rect 10793 27081 10827 27115
rect 11161 27081 11195 27115
rect 4537 27013 4571 27047
rect 8585 27013 8619 27047
rect 8861 27013 8895 27047
rect 11437 27013 11471 27047
rect 4169 26945 4203 26979
rect 6101 26945 6135 26979
rect 6285 26945 6319 26979
rect 9781 26945 9815 26979
rect 11713 26945 11747 26979
rect 1317 26877 1351 26911
rect 1501 26877 1535 26911
rect 1593 26877 1627 26911
rect 4935 26877 4969 26911
rect 5089 26877 5123 26911
rect 6009 26877 6043 26911
rect 6193 26877 6227 26911
rect 6745 26877 6779 26911
rect 7113 26877 7147 26911
rect 7297 26877 7331 26911
rect 7389 26877 7423 26911
rect 7481 26877 7515 26911
rect 7665 26877 7699 26911
rect 7941 26877 7975 26911
rect 8217 26877 8251 26911
rect 8401 26877 8435 26911
rect 8585 26877 8619 26911
rect 8769 26877 8803 26911
rect 8953 26877 8987 26911
rect 9045 26877 9079 26911
rect 9689 26877 9723 26911
rect 9965 26877 9999 26911
rect 10609 26877 10643 26911
rect 11069 26877 11103 26911
rect 11253 26877 11287 26911
rect 11805 26877 11839 26911
rect 857 26809 891 26843
rect 10425 26809 10459 26843
rect 4721 26741 4755 26775
rect 5825 26741 5859 26775
rect 6561 26741 6595 26775
rect 6929 26741 6963 26775
rect 8125 26741 8159 26775
rect 9321 26741 9355 26775
rect 10149 26741 10183 26775
rect 2519 26537 2553 26571
rect 6009 26537 6043 26571
rect 7205 26537 7239 26571
rect 8953 26537 8987 26571
rect 2789 26469 2823 26503
rect 2973 26469 3007 26503
rect 4353 26469 4387 26503
rect 857 26401 891 26435
rect 1124 26401 1158 26435
rect 2421 26401 2455 26435
rect 2605 26401 2639 26435
rect 2697 26401 2731 26435
rect 3065 26401 3099 26435
rect 3985 26401 4019 26435
rect 4813 26401 4847 26435
rect 4997 26401 5031 26435
rect 5365 26401 5399 26435
rect 6285 26401 6319 26435
rect 6561 26401 6595 26435
rect 6837 26401 6871 26435
rect 7481 26401 7515 26435
rect 7573 26401 7607 26435
rect 7665 26401 7699 26435
rect 7849 26401 7883 26435
rect 7941 26401 7975 26435
rect 8217 26401 8251 26435
rect 8401 26401 8435 26435
rect 8493 26391 8527 26425
rect 8585 26401 8619 26435
rect 8769 26401 8803 26435
rect 9229 26401 9263 26435
rect 9321 26401 9355 26435
rect 9413 26401 9447 26435
rect 9597 26401 9631 26435
rect 4905 26333 4939 26367
rect 5273 26333 5307 26367
rect 5457 26333 5491 26367
rect 5549 26333 5583 26367
rect 6745 26333 6779 26367
rect 9045 26333 9079 26367
rect 9505 26333 9539 26367
rect 2237 26265 2271 26299
rect 2789 26265 2823 26299
rect 8217 26265 8251 26299
rect 9137 26265 9171 26299
rect 4353 26197 4387 26231
rect 4537 26197 4571 26231
rect 5089 26197 5123 26231
rect 6469 26197 6503 26231
rect 7297 26197 7331 26231
rect 2421 25993 2455 26027
rect 2605 25993 2639 26027
rect 4813 25993 4847 26027
rect 6653 25993 6687 26027
rect 2329 25925 2363 25959
rect 10701 25925 10735 25959
rect 1041 25857 1075 25891
rect 2513 25857 2547 25891
rect 3525 25857 3559 25891
rect 5917 25857 5951 25891
rect 6101 25857 6135 25891
rect 6193 25857 6227 25891
rect 7021 25857 7055 25891
rect 10241 25857 10275 25891
rect 1501 25789 1535 25823
rect 1685 25789 1719 25823
rect 1777 25789 1811 25823
rect 2237 25789 2271 25823
rect 2789 25789 2823 25823
rect 2973 25789 3007 25823
rect 3065 25789 3099 25823
rect 3709 25789 3743 25823
rect 3985 25789 4019 25823
rect 4169 25789 4203 25823
rect 4537 25789 4571 25823
rect 4629 25789 4663 25823
rect 5457 25789 5491 25823
rect 6009 25789 6043 25823
rect 6683 25789 6717 25823
rect 6837 25789 6871 25823
rect 6929 25789 6963 25823
rect 7113 25789 7147 25823
rect 8585 25789 8619 25823
rect 9321 25789 9355 25823
rect 9505 25789 9539 25823
rect 10425 25789 10459 25823
rect 10517 25789 10551 25823
rect 10885 25789 10919 25823
rect 11161 25789 11195 25823
rect 11345 25789 11379 25823
rect 11897 25789 11931 25823
rect 11989 25789 12023 25823
rect 8769 25721 8803 25755
rect 3893 25653 3927 25687
rect 5641 25653 5675 25687
rect 6377 25653 6411 25687
rect 9413 25653 9447 25687
rect 10241 25653 10275 25687
rect 11253 25653 11287 25687
rect 12173 25653 12207 25687
rect 857 25449 891 25483
rect 2881 25449 2915 25483
rect 3157 25449 3191 25483
rect 6653 25449 6687 25483
rect 7389 25449 7423 25483
rect 9229 25449 9263 25483
rect 10333 25449 10367 25483
rect 10609 25449 10643 25483
rect 10977 25449 11011 25483
rect 2697 25381 2731 25415
rect 5181 25381 5215 25415
rect 9689 25381 9723 25415
rect 10425 25381 10459 25415
rect 1970 25313 2004 25347
rect 2237 25313 2271 25347
rect 2605 25313 2639 25347
rect 2973 25313 3007 25347
rect 3341 25313 3375 25347
rect 3525 25313 3559 25347
rect 4813 25313 4847 25347
rect 4997 25313 5031 25347
rect 6929 25313 6963 25347
rect 7021 25313 7055 25347
rect 7113 25313 7147 25347
rect 7297 25313 7331 25347
rect 7665 25313 7699 25347
rect 7941 25313 7975 25347
rect 8585 25313 8619 25347
rect 9413 25313 9447 25347
rect 9965 25313 9999 25347
rect 10701 25313 10735 25347
rect 11345 25313 11379 25347
rect 11989 25313 12023 25347
rect 2329 25245 2363 25279
rect 7389 25245 7423 25279
rect 7849 25245 7883 25279
rect 8493 25245 8527 25279
rect 8953 25245 8987 25279
rect 9505 25245 9539 25279
rect 10057 25245 10091 25279
rect 11253 25245 11287 25279
rect 11897 25245 11931 25279
rect 2513 25177 2547 25211
rect 8309 25177 8343 25211
rect 10425 25177 10459 25211
rect 11621 25177 11655 25211
rect 2421 25109 2455 25143
rect 2697 25109 2731 25143
rect 7573 25109 7607 25143
rect 9689 25109 9723 25143
rect 3341 24905 3375 24939
rect 6561 24905 6595 24939
rect 7021 24905 7055 24939
rect 7849 24905 7883 24939
rect 7941 24905 7975 24939
rect 9413 24905 9447 24939
rect 10241 24905 10275 24939
rect 5365 24837 5399 24871
rect 7389 24769 7423 24803
rect 7481 24769 7515 24803
rect 8493 24769 8527 24803
rect 9505 24769 9539 24803
rect 10701 24769 10735 24803
rect 11161 24769 11195 24803
rect 11437 24769 11471 24803
rect 12173 24769 12207 24803
rect 1501 24701 1535 24735
rect 1685 24701 1719 24735
rect 1777 24701 1811 24735
rect 2145 24701 2179 24735
rect 2329 24701 2363 24735
rect 2421 24701 2455 24735
rect 2605 24701 2639 24735
rect 3525 24701 3559 24735
rect 3892 24701 3926 24735
rect 3985 24701 4019 24735
rect 4445 24701 4479 24735
rect 4813 24701 4847 24735
rect 5549 24701 5583 24735
rect 5733 24701 5767 24735
rect 5917 24701 5951 24735
rect 6193 24701 6227 24735
rect 6469 24701 6503 24735
rect 6745 24701 6779 24735
rect 6837 24701 6871 24735
rect 7113 24701 7147 24735
rect 7297 24701 7331 24735
rect 7665 24701 7699 24735
rect 8217 24701 8251 24735
rect 8401 24701 8435 24735
rect 8769 24701 8803 24735
rect 8953 24701 8987 24735
rect 9045 24701 9079 24735
rect 9137 24701 9171 24735
rect 9781 24701 9815 24735
rect 9873 24701 9907 24735
rect 9965 24701 9999 24735
rect 10149 24701 10183 24735
rect 10609 24701 10643 24735
rect 11069 24701 11103 24735
rect 11897 24701 11931 24735
rect 11989 24701 12023 24735
rect 12081 24701 12115 24735
rect 1041 24633 1075 24667
rect 2513 24633 2547 24667
rect 6009 24633 6043 24667
rect 6377 24633 6411 24667
rect 7941 24633 7975 24667
rect 2237 24565 2271 24599
rect 3617 24565 3651 24599
rect 5825 24565 5859 24599
rect 8125 24565 8159 24599
rect 11713 24565 11747 24599
rect 2421 24361 2455 24395
rect 3617 24361 3651 24395
rect 4813 24361 4847 24395
rect 7573 24361 7607 24395
rect 8401 24361 8435 24395
rect 9229 24361 9263 24395
rect 4997 24293 5031 24327
rect 6745 24293 6779 24327
rect 6929 24293 6963 24327
rect 857 24225 891 24259
rect 1124 24225 1158 24259
rect 2605 24225 2639 24259
rect 2789 24225 2823 24259
rect 3341 24225 3375 24259
rect 3709 24225 3743 24259
rect 3801 24225 3835 24259
rect 3985 24225 4019 24259
rect 4169 24225 4203 24259
rect 4353 24225 4387 24259
rect 5181 24225 5215 24259
rect 5457 24225 5491 24259
rect 5549 24225 5583 24259
rect 5825 24225 5859 24259
rect 6009 24225 6043 24259
rect 6285 24225 6319 24259
rect 6469 24225 6503 24259
rect 6561 24225 6595 24259
rect 7021 24225 7055 24259
rect 7205 24225 7239 24259
rect 7297 24225 7331 24259
rect 7389 24225 7423 24259
rect 7665 24225 7699 24259
rect 7849 24225 7883 24259
rect 8217 24225 8251 24259
rect 8493 24225 8527 24259
rect 9137 24225 9171 24259
rect 9321 24225 9355 24259
rect 9689 24225 9723 24259
rect 10241 24225 10275 24259
rect 10333 24225 10367 24259
rect 10425 24225 10459 24259
rect 11161 24225 11195 24259
rect 11621 24225 11655 24259
rect 11805 24225 11839 24259
rect 3525 24157 3559 24191
rect 6193 24157 6227 24191
rect 7941 24157 7975 24191
rect 8033 24157 8067 24191
rect 10517 24157 10551 24191
rect 10977 24157 11011 24191
rect 11345 24157 11379 24191
rect 11713 24157 11747 24191
rect 11897 24157 11931 24191
rect 3433 24089 3467 24123
rect 4629 24089 4663 24123
rect 8585 24089 8619 24123
rect 10057 24089 10091 24123
rect 2237 24021 2271 24055
rect 4077 24021 4111 24055
rect 5365 24021 5399 24055
rect 6377 24021 6411 24055
rect 9873 24021 9907 24055
rect 11437 24021 11471 24055
rect 5549 23817 5583 23851
rect 5825 23817 5859 23851
rect 10149 23817 10183 23851
rect 11989 23817 12023 23851
rect 3065 23749 3099 23783
rect 4445 23749 4479 23783
rect 1685 23681 1719 23715
rect 3709 23681 3743 23715
rect 3893 23681 3927 23715
rect 5273 23681 5307 23715
rect 6469 23681 6503 23715
rect 6628 23681 6662 23715
rect 6745 23681 6779 23715
rect 7021 23681 7055 23715
rect 1133 23613 1167 23647
rect 1409 23613 1443 23647
rect 3617 23613 3651 23647
rect 4077 23613 4111 23647
rect 4261 23613 4295 23647
rect 4537 23613 4571 23647
rect 4629 23613 4663 23647
rect 4905 23613 4939 23647
rect 5089 23613 5123 23647
rect 5181 23613 5215 23647
rect 5365 23613 5399 23647
rect 5733 23613 5767 23647
rect 7481 23613 7515 23647
rect 7665 23613 7699 23647
rect 10057 23613 10091 23647
rect 10241 23613 10275 23647
rect 11713 23613 11747 23647
rect 11805 23613 11839 23647
rect 12081 23613 12115 23647
rect 12265 23613 12299 23647
rect 1952 23545 1986 23579
rect 4353 23545 4387 23579
rect 3249 23477 3283 23511
rect 4169 23477 4203 23511
rect 5089 23477 5123 23511
rect 12173 23477 12207 23511
rect 2237 23273 2271 23307
rect 11345 23273 11379 23307
rect 12173 23273 12207 23307
rect 2789 23205 2823 23239
rect 4445 23205 4479 23239
rect 5457 23205 5491 23239
rect 7205 23205 7239 23239
rect 8677 23205 8711 23239
rect 11897 23205 11931 23239
rect 857 23137 891 23171
rect 1124 23137 1158 23171
rect 2329 23137 2363 23171
rect 4537 23137 4571 23171
rect 4721 23137 4755 23171
rect 4813 23137 4847 23171
rect 5089 23137 5123 23171
rect 5825 23137 5859 23171
rect 6009 23137 6043 23171
rect 6377 23137 6411 23171
rect 6745 23137 6779 23171
rect 6929 23137 6963 23171
rect 7021 23137 7055 23171
rect 7389 23137 7423 23171
rect 7481 23137 7515 23171
rect 7665 23137 7699 23171
rect 7849 23137 7883 23171
rect 8033 23137 8067 23171
rect 8309 23137 8343 23171
rect 8585 23137 8619 23171
rect 8861 23137 8895 23171
rect 9321 23137 9355 23171
rect 10057 23137 10091 23171
rect 10241 23137 10275 23171
rect 10609 23137 10643 23171
rect 10793 23137 10827 23171
rect 11161 23137 11195 23171
rect 11437 23137 11471 23171
rect 11529 23137 11563 23171
rect 11713 23137 11747 23171
rect 11989 23137 12023 23171
rect 4905 23069 4939 23103
rect 6101 23069 6135 23103
rect 6193 23069 6227 23103
rect 7757 23069 7791 23103
rect 9597 23069 9631 23103
rect 5641 23001 5675 23035
rect 9045 23001 9079 23035
rect 9505 23001 9539 23035
rect 10977 23001 11011 23035
rect 2513 22933 2547 22967
rect 5273 22933 5307 22967
rect 6561 22933 6595 22967
rect 6929 22933 6963 22967
rect 8217 22933 8251 22967
rect 8401 22933 8435 22967
rect 9137 22933 9171 22967
rect 10149 22933 10183 22967
rect 10609 22933 10643 22967
rect 3801 22729 3835 22763
rect 4353 22729 4387 22763
rect 5365 22729 5399 22763
rect 6929 22729 6963 22763
rect 8861 22729 8895 22763
rect 10057 22729 10091 22763
rect 10977 22729 11011 22763
rect 11437 22729 11471 22763
rect 1041 22661 1075 22695
rect 2513 22661 2547 22695
rect 4905 22661 4939 22695
rect 12173 22661 12207 22695
rect 1317 22593 1351 22627
rect 2053 22593 2087 22627
rect 3525 22593 3559 22627
rect 5733 22593 5767 22627
rect 9873 22593 9907 22627
rect 10701 22593 10735 22627
rect 1225 22525 1259 22559
rect 1777 22525 1811 22559
rect 1961 22525 1995 22559
rect 2697 22525 2731 22559
rect 2789 22525 2823 22559
rect 2973 22525 3007 22559
rect 3065 22525 3099 22559
rect 3433 22525 3467 22559
rect 4077 22525 4111 22559
rect 4169 22525 4203 22559
rect 4445 22525 4479 22559
rect 5641 22525 5675 22559
rect 6377 22525 6411 22559
rect 8217 22525 8251 22559
rect 8401 22525 8435 22559
rect 8769 22525 8803 22559
rect 9045 22525 9079 22559
rect 9137 22525 9171 22559
rect 9781 22525 9815 22559
rect 10057 22525 10091 22559
rect 10241 22525 10275 22559
rect 10609 22525 10643 22559
rect 11069 22525 11103 22559
rect 11345 22525 11379 22559
rect 3893 22457 3927 22491
rect 4537 22457 4571 22491
rect 6193 22457 6227 22491
rect 11253 22457 11287 22491
rect 11713 22457 11747 22491
rect 12173 22457 12207 22491
rect 4997 22389 5031 22423
rect 6009 22389 6043 22423
rect 8585 22389 8619 22423
rect 9321 22389 9355 22423
rect 9413 22389 9447 22423
rect 11345 22389 11379 22423
rect 11621 22389 11655 22423
rect 5273 22185 5307 22219
rect 10793 22185 10827 22219
rect 11345 22185 11379 22219
rect 11529 22185 11563 22219
rect 11713 22185 11747 22219
rect 3249 22117 3283 22151
rect 10057 22117 10091 22151
rect 10241 22117 10275 22151
rect 3617 22049 3651 22083
rect 3709 22049 3743 22083
rect 4077 22049 4111 22083
rect 4261 22049 4295 22083
rect 4537 22049 4571 22083
rect 4905 22049 4939 22083
rect 5181 22049 5215 22083
rect 5457 22049 5491 22083
rect 6791 22049 6825 22083
rect 8125 22049 8159 22083
rect 8217 22049 8251 22083
rect 8493 22049 8527 22083
rect 8953 22049 8987 22083
rect 9045 22049 9079 22083
rect 9142 22049 9176 22083
rect 9321 22049 9355 22083
rect 9872 22049 9906 22083
rect 9965 22049 9999 22083
rect 10333 22049 10367 22083
rect 10517 22049 10551 22083
rect 10609 22049 10643 22083
rect 11161 22049 11195 22083
rect 11437 22049 11471 22083
rect 11710 22049 11744 22083
rect 12081 22049 12115 22083
rect 6653 21981 6687 22015
rect 6929 21981 6963 22015
rect 7205 21981 7239 22015
rect 7665 21981 7699 22015
rect 7849 21981 7883 22015
rect 8401 21981 8435 22015
rect 12173 21981 12207 22015
rect 3893 21913 3927 21947
rect 6009 21913 6043 21947
rect 1041 21845 1075 21879
rect 1961 21845 1995 21879
rect 3433 21845 3467 21879
rect 4077 21845 4111 21879
rect 4353 21845 4387 21879
rect 4721 21845 4755 21879
rect 5641 21845 5675 21879
rect 7941 21845 7975 21879
rect 8677 21845 8711 21879
rect 9781 21845 9815 21879
rect 10333 21845 10367 21879
rect 10977 21845 11011 21879
rect 3893 21641 3927 21675
rect 4445 21641 4479 21675
rect 5549 21641 5583 21675
rect 5825 21641 5859 21675
rect 7205 21641 7239 21675
rect 8401 21641 8435 21675
rect 2789 21573 2823 21607
rect 5733 21573 5767 21607
rect 6561 21573 6595 21607
rect 6653 21573 6687 21607
rect 7297 21573 7331 21607
rect 9965 21573 9999 21607
rect 10057 21573 10091 21607
rect 2881 21505 2915 21539
rect 3341 21505 3375 21539
rect 4721 21505 4755 21539
rect 7389 21505 7423 21539
rect 7941 21505 7975 21539
rect 8217 21505 8251 21539
rect 1409 21437 1443 21471
rect 2145 21437 2179 21471
rect 2605 21437 2639 21471
rect 3617 21437 3651 21471
rect 3801 21437 3835 21471
rect 3985 21437 4019 21471
rect 4261 21437 4295 21471
rect 4537 21437 4571 21471
rect 4635 21437 4669 21471
rect 4813 21437 4847 21471
rect 5825 21437 5859 21471
rect 6101 21437 6135 21471
rect 6469 21437 6503 21471
rect 6745 21437 6779 21471
rect 7113 21437 7147 21471
rect 7849 21437 7883 21471
rect 8585 21437 8619 21471
rect 8677 21437 8711 21471
rect 8861 21437 8895 21471
rect 8953 21437 8987 21471
rect 9689 21437 9723 21471
rect 9781 21437 9815 21471
rect 10057 21437 10091 21471
rect 10241 21437 10275 21471
rect 10333 21437 10367 21471
rect 11897 21437 11931 21471
rect 12081 21437 12115 21471
rect 1133 21369 1167 21403
rect 4077 21369 4111 21403
rect 5365 21369 5399 21403
rect 5565 21369 5599 21403
rect 9965 21369 9999 21403
rect 2421 21301 2455 21335
rect 6009 21301 6043 21335
rect 6285 21301 6319 21335
rect 11713 21301 11747 21335
rect 2421 21097 2455 21131
rect 2973 21097 3007 21131
rect 5457 21097 5491 21131
rect 7757 21097 7791 21131
rect 11529 21097 11563 21131
rect 1970 20961 2004 20995
rect 2605 20961 2639 20995
rect 2789 20961 2823 20995
rect 3157 20961 3191 20995
rect 3341 20961 3375 20995
rect 3709 20961 3743 20995
rect 3893 20961 3927 20995
rect 4261 20961 4295 20995
rect 4445 20961 4479 20995
rect 4629 20961 4663 20995
rect 4813 20961 4847 20995
rect 5273 20961 5307 20995
rect 5549 20961 5583 20995
rect 5825 20961 5859 20995
rect 6745 20961 6779 20995
rect 6929 20961 6963 20995
rect 7389 20961 7423 20995
rect 7481 20961 7515 20995
rect 11069 20961 11103 20995
rect 11253 20961 11287 20995
rect 11345 20961 11379 20995
rect 11437 20961 11471 20995
rect 11621 20961 11655 20995
rect 2237 20893 2271 20927
rect 2893 20893 2927 20927
rect 3433 20893 3467 20927
rect 4537 20893 4571 20927
rect 4721 20893 4755 20927
rect 7113 20893 7147 20927
rect 7297 20893 7331 20927
rect 7757 20893 7791 20927
rect 4077 20825 4111 20859
rect 6009 20825 6043 20859
rect 7205 20825 7239 20859
rect 857 20757 891 20791
rect 3525 20757 3559 20791
rect 5089 20757 5123 20791
rect 6929 20757 6963 20791
rect 7573 20757 7607 20791
rect 11161 20757 11195 20791
rect 5641 20553 5675 20587
rect 7665 20553 7699 20587
rect 7941 20553 7975 20587
rect 8769 20553 8803 20587
rect 9873 20553 9907 20587
rect 11253 20553 11287 20587
rect 2697 20485 2731 20519
rect 4813 20485 4847 20519
rect 5917 20485 5951 20519
rect 6009 20485 6043 20519
rect 11713 20485 11747 20519
rect 857 20417 891 20451
rect 1593 20417 1627 20451
rect 2789 20417 2823 20451
rect 3617 20417 3651 20451
rect 3709 20417 3743 20451
rect 4445 20417 4479 20451
rect 6561 20417 6595 20451
rect 7205 20417 7239 20451
rect 8953 20417 8987 20451
rect 10057 20417 10091 20451
rect 10885 20417 10919 20451
rect 1317 20349 1351 20383
rect 1501 20349 1535 20383
rect 2513 20349 2547 20383
rect 3433 20349 3467 20383
rect 4261 20349 4295 20383
rect 4537 20349 4571 20383
rect 4629 20349 4663 20383
rect 5825 20349 5859 20383
rect 6101 20349 6135 20383
rect 6469 20349 6503 20383
rect 6653 20349 6687 20383
rect 6745 20349 6779 20383
rect 7113 20349 7147 20383
rect 7389 20349 7423 20383
rect 7481 20349 7515 20383
rect 7757 20349 7791 20383
rect 8401 20349 8435 20383
rect 8585 20349 8619 20383
rect 8677 20349 8711 20383
rect 9045 20349 9079 20383
rect 9138 20349 9172 20383
rect 9510 20349 9544 20383
rect 10149 20349 10183 20383
rect 10977 20349 11011 20383
rect 4077 20281 4111 20315
rect 8953 20281 8987 20315
rect 9321 20281 9355 20315
rect 9413 20281 9447 20315
rect 11529 20281 11563 20315
rect 2329 20213 2363 20247
rect 3249 20213 3283 20247
rect 6285 20213 6319 20247
rect 8493 20213 8527 20247
rect 9689 20213 9723 20247
rect 949 20009 983 20043
rect 2697 20009 2731 20043
rect 3433 20009 3467 20043
rect 3801 20009 3835 20043
rect 4077 20009 4111 20043
rect 6929 20009 6963 20043
rect 11345 20009 11379 20043
rect 2513 19941 2547 19975
rect 6193 19941 6227 19975
rect 10701 19941 10735 19975
rect 11897 19941 11931 19975
rect 1133 19873 1167 19907
rect 2145 19873 2179 19907
rect 2789 19873 2823 19907
rect 3138 19863 3172 19897
rect 3249 19873 3283 19907
rect 3525 19873 3559 19907
rect 3617 19873 3651 19907
rect 3893 19873 3927 19907
rect 3985 19873 4019 19907
rect 4169 19873 4203 19907
rect 4445 19873 4479 19907
rect 4721 19873 4755 19907
rect 4813 19873 4847 19907
rect 4997 19873 5031 19907
rect 5365 19873 5399 19907
rect 5825 19873 5859 19907
rect 6561 19873 6595 19907
rect 7113 19873 7147 19907
rect 7205 19873 7239 19907
rect 7481 19873 7515 19907
rect 7849 19873 7883 19907
rect 7941 19873 7975 19907
rect 8033 19873 8067 19907
rect 8217 19873 8251 19907
rect 8677 19873 8711 19907
rect 9321 19873 9355 19907
rect 10057 19873 10091 19907
rect 10333 19873 10367 19907
rect 10517 19873 10551 19907
rect 10609 19873 10643 19907
rect 10793 19873 10827 19907
rect 11161 19873 11195 19907
rect 11437 19873 11471 19907
rect 11713 19873 11747 19907
rect 11989 19873 12023 19907
rect 1317 19805 1351 19839
rect 1409 19805 1443 19839
rect 2421 19805 2455 19839
rect 2881 19805 2915 19839
rect 4629 19805 4663 19839
rect 7389 19805 7423 19839
rect 8769 19805 8803 19839
rect 8953 19805 8987 19839
rect 9229 19805 9263 19839
rect 9781 19805 9815 19839
rect 2329 19737 2363 19771
rect 3065 19737 3099 19771
rect 3249 19737 3283 19771
rect 8309 19737 8343 19771
rect 11529 19737 11563 19771
rect 1961 19669 1995 19703
rect 2513 19669 2547 19703
rect 2973 19669 3007 19703
rect 3617 19669 3651 19703
rect 4261 19669 4295 19703
rect 5181 19669 5215 19703
rect 6745 19669 6779 19703
rect 7573 19669 7607 19703
rect 9689 19669 9723 19703
rect 9873 19669 9907 19703
rect 10241 19669 10275 19703
rect 10517 19669 10551 19703
rect 10977 19669 11011 19703
rect 1409 19465 1443 19499
rect 2513 19465 2547 19499
rect 7481 19465 7515 19499
rect 7757 19465 7791 19499
rect 9413 19465 9447 19499
rect 10793 19465 10827 19499
rect 11805 19465 11839 19499
rect 9689 19397 9723 19431
rect 6193 19329 6227 19363
rect 8769 19329 8803 19363
rect 9137 19329 9171 19363
rect 1593 19261 1627 19295
rect 1777 19261 1811 19295
rect 1869 19261 1903 19295
rect 2237 19261 2271 19295
rect 5549 19261 5583 19295
rect 5733 19261 5767 19295
rect 6469 19261 6503 19295
rect 6586 19261 6620 19295
rect 6745 19261 6779 19295
rect 7481 19261 7515 19295
rect 7665 19261 7699 19295
rect 7941 19261 7975 19295
rect 8125 19261 8159 19295
rect 8217 19261 8251 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 8677 19261 8711 19295
rect 8953 19261 8987 19295
rect 9321 19261 9355 19295
rect 9498 19261 9532 19295
rect 9873 19261 9907 19295
rect 10241 19261 10275 19295
rect 10517 19261 10551 19295
rect 10609 19261 10643 19295
rect 10885 19261 10919 19295
rect 11713 19261 11747 19295
rect 11989 19261 12023 19295
rect 2513 19193 2547 19227
rect 9965 19193 9999 19227
rect 10057 19193 10091 19227
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 11529 19193 11563 19227
rect 2329 19125 2363 19159
rect 7389 19125 7423 19159
rect 12173 19125 12207 19159
rect 2053 18921 2087 18955
rect 7941 18921 7975 18955
rect 9597 18921 9631 18955
rect 9781 18921 9815 18955
rect 12173 18921 12207 18955
rect 3249 18853 3283 18887
rect 4445 18853 4479 18887
rect 5457 18853 5491 18887
rect 10333 18853 10367 18887
rect 1409 18785 1443 18819
rect 1593 18785 1627 18819
rect 2237 18785 2271 18819
rect 2605 18785 2639 18819
rect 2789 18785 2823 18819
rect 2973 18785 3007 18819
rect 3065 18785 3099 18819
rect 3157 18785 3191 18819
rect 3433 18785 3467 18819
rect 3617 18785 3651 18819
rect 3801 18785 3835 18819
rect 4629 18785 4663 18819
rect 4997 18785 5031 18819
rect 5181 18785 5215 18819
rect 5273 18785 5307 18819
rect 5641 18785 5675 18819
rect 5825 18785 5859 18819
rect 6862 18785 6896 18819
rect 7021 18785 7055 18819
rect 8125 18785 8159 18819
rect 8309 18785 8343 18819
rect 8401 18785 8435 18819
rect 8585 18785 8619 18819
rect 9505 18785 9539 18819
rect 9689 18785 9723 18819
rect 9965 18785 9999 18819
rect 10241 18785 10275 18819
rect 10517 18785 10551 18819
rect 10609 18785 10643 18819
rect 11621 18785 11655 18819
rect 12081 18785 12115 18819
rect 12265 18785 12299 18819
rect 949 18717 983 18751
rect 1685 18717 1719 18751
rect 2513 18717 2547 18751
rect 4813 18717 4847 18751
rect 4905 18717 4939 18751
rect 6009 18717 6043 18751
rect 6469 18717 6503 18751
rect 6745 18717 6779 18751
rect 7757 18717 7791 18751
rect 10149 18717 10183 18751
rect 11529 18717 11563 18751
rect 11989 18717 12023 18751
rect 8217 18649 8251 18683
rect 10333 18649 10367 18683
rect 2421 18581 2455 18615
rect 3433 18581 3467 18615
rect 3709 18581 3743 18615
rect 7665 18581 7699 18615
rect 8769 18581 8803 18615
rect 857 18377 891 18411
rect 2329 18377 2363 18411
rect 3893 18377 3927 18411
rect 7573 18377 7607 18411
rect 8401 18377 8435 18411
rect 10425 18377 10459 18411
rect 11989 18377 12023 18411
rect 2697 18309 2731 18343
rect 9137 18309 9171 18343
rect 11253 18309 11287 18343
rect 11897 18309 11931 18343
rect 3525 18241 3559 18275
rect 3617 18241 3651 18275
rect 3801 18241 3835 18275
rect 8769 18241 8803 18275
rect 1981 18173 2015 18207
rect 2237 18173 2271 18207
rect 2513 18173 2547 18207
rect 2789 18173 2823 18207
rect 3341 18173 3375 18207
rect 3433 18173 3467 18207
rect 4169 18173 4203 18207
rect 4261 18173 4295 18207
rect 4445 18173 4479 18207
rect 6745 18173 6779 18207
rect 7665 18173 7699 18207
rect 7849 18173 7883 18207
rect 8585 18173 8619 18207
rect 8677 18173 8711 18207
rect 8861 18173 8895 18207
rect 9321 18173 9355 18207
rect 9413 18173 9447 18207
rect 10333 18173 10367 18207
rect 10517 18173 10551 18207
rect 10977 18173 11011 18207
rect 11253 18173 11287 18207
rect 11713 18173 11747 18207
rect 11989 18173 12023 18207
rect 3893 18105 3927 18139
rect 6561 18105 6595 18139
rect 7205 18105 7239 18139
rect 7389 18105 7423 18139
rect 9137 18105 9171 18139
rect 4077 18037 4111 18071
rect 4353 18037 4387 18071
rect 6929 18037 6963 18071
rect 8033 18037 8067 18071
rect 11069 18037 11103 18071
rect 2973 17833 3007 17867
rect 9597 17833 9631 17867
rect 10793 17833 10827 17867
rect 11805 17833 11839 17867
rect 4997 17765 5031 17799
rect 6837 17765 6871 17799
rect 7021 17765 7055 17799
rect 7481 17765 7515 17799
rect 8677 17765 8711 17799
rect 9321 17765 9355 17799
rect 1981 17697 2015 17731
rect 2513 17697 2547 17731
rect 2789 17697 2823 17731
rect 3065 17697 3099 17731
rect 3525 17697 3559 17731
rect 3617 17697 3651 17731
rect 3985 17697 4019 17731
rect 4261 17697 4295 17731
rect 4721 17697 4755 17731
rect 5181 17697 5215 17731
rect 5365 17697 5399 17731
rect 5825 17697 5859 17731
rect 6009 17697 6043 17731
rect 6193 17697 6227 17731
rect 6377 17697 6411 17731
rect 7665 17697 7699 17731
rect 7849 17697 7883 17731
rect 7941 17697 7975 17731
rect 8217 17697 8251 17731
rect 8493 17697 8527 17731
rect 8953 17697 8987 17731
rect 9101 17697 9135 17731
rect 9229 17697 9263 17731
rect 9418 17697 9452 17731
rect 9873 17697 9907 17731
rect 10149 17697 10183 17731
rect 10609 17697 10643 17731
rect 11345 17697 11379 17731
rect 11713 17697 11747 17731
rect 2237 17629 2271 17663
rect 3341 17629 3375 17663
rect 3433 17629 3467 17663
rect 4077 17629 4111 17663
rect 4169 17629 4203 17663
rect 6101 17629 6135 17663
rect 6653 17629 6687 17663
rect 8033 17629 8067 17663
rect 9689 17629 9723 17663
rect 9965 17629 9999 17663
rect 10057 17629 10091 17663
rect 10333 17629 10367 17663
rect 11437 17629 11471 17663
rect 8861 17561 8895 17595
rect 10977 17561 11011 17595
rect 857 17493 891 17527
rect 2329 17493 2363 17527
rect 2697 17493 2731 17527
rect 3157 17493 3191 17527
rect 3801 17493 3835 17527
rect 4537 17493 4571 17527
rect 6561 17493 6595 17527
rect 7205 17493 7239 17527
rect 8401 17493 8435 17527
rect 10425 17493 10459 17527
rect 2513 17289 2547 17323
rect 4261 17289 4295 17323
rect 5273 17289 5307 17323
rect 6377 17289 6411 17323
rect 6561 17289 6595 17323
rect 2605 17221 2639 17255
rect 5457 17221 5491 17255
rect 10425 17221 10459 17255
rect 1225 17153 1259 17187
rect 7021 17153 7055 17187
rect 8769 17153 8803 17187
rect 9965 17153 9999 17187
rect 11529 17153 11563 17187
rect 1317 17085 1351 17119
rect 1501 17085 1535 17119
rect 2237 17085 2271 17119
rect 2513 17085 2547 17119
rect 2605 17085 2639 17119
rect 2881 17085 2915 17119
rect 4169 17085 4203 17119
rect 4353 17085 4387 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 5365 17085 5399 17119
rect 5641 17085 5675 17119
rect 5825 17085 5859 17119
rect 6101 17085 6135 17119
rect 6193 17085 6227 17119
rect 6469 17085 6503 17119
rect 6745 17085 6779 17119
rect 6837 17085 6871 17119
rect 7113 17085 7147 17119
rect 7665 17085 7699 17119
rect 7849 17085 7883 17119
rect 7941 17085 7975 17119
rect 8033 17085 8067 17119
rect 8217 17085 8251 17119
rect 8401 17085 8435 17119
rect 8585 17085 8619 17119
rect 8677 17085 8711 17119
rect 8953 17085 8987 17119
rect 9505 17085 9539 17119
rect 9781 17085 9815 17119
rect 10057 17085 10091 17119
rect 10609 17085 10643 17119
rect 10793 17085 10827 17119
rect 11437 17085 11471 17119
rect 11713 17085 11747 17119
rect 12081 17085 12115 17119
rect 1961 17017 1995 17051
rect 2329 17017 2363 17051
rect 2789 17017 2823 17051
rect 10701 17017 10735 17051
rect 10885 17017 10919 17051
rect 11897 17017 11931 17051
rect 4813 16949 4847 16983
rect 5917 16949 5951 16983
rect 7481 16949 7515 16983
rect 9137 16949 9171 16983
rect 9321 16949 9355 16983
rect 9689 16949 9723 16983
rect 11161 16949 11195 16983
rect 3801 16745 3835 16779
rect 4261 16745 4295 16779
rect 8217 16745 8251 16779
rect 8769 16745 8803 16779
rect 9689 16745 9723 16779
rect 10241 16745 10275 16779
rect 11345 16745 11379 16779
rect 949 16677 983 16711
rect 3985 16677 4019 16711
rect 4169 16677 4203 16711
rect 4997 16677 5031 16711
rect 5641 16677 5675 16711
rect 9781 16677 9815 16711
rect 10701 16677 10735 16711
rect 1409 16609 1443 16643
rect 1593 16609 1627 16643
rect 4537 16609 4571 16643
rect 5273 16609 5307 16643
rect 5365 16609 5399 16643
rect 6285 16609 6319 16643
rect 6653 16609 6687 16643
rect 6837 16609 6871 16643
rect 7297 16609 7331 16643
rect 7481 16609 7515 16643
rect 7665 16609 7699 16643
rect 7849 16609 7883 16643
rect 8309 16609 8343 16643
rect 8585 16609 8619 16643
rect 8769 16609 8803 16643
rect 8861 16609 8895 16643
rect 8953 16609 8987 16643
rect 9045 16609 9079 16643
rect 9505 16609 9539 16643
rect 10517 16609 10551 16643
rect 11253 16609 11287 16643
rect 11437 16609 11471 16643
rect 11805 16609 11839 16643
rect 11989 16609 12023 16643
rect 12081 16609 12115 16643
rect 1685 16541 1719 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 4997 16541 5031 16575
rect 5641 16541 5675 16575
rect 6469 16541 6503 16575
rect 6561 16541 6595 16575
rect 7573 16541 7607 16575
rect 9321 16541 9355 16575
rect 5181 16473 5215 16507
rect 10057 16473 10091 16507
rect 10333 16473 10367 16507
rect 5457 16405 5491 16439
rect 6101 16405 6135 16439
rect 7113 16405 7147 16439
rect 11805 16405 11839 16439
rect 2237 16201 2271 16235
rect 2789 16201 2823 16235
rect 6193 16201 6227 16235
rect 8033 16201 8067 16235
rect 8953 16201 8987 16235
rect 9781 16201 9815 16235
rect 11621 16201 11655 16235
rect 11989 16201 12023 16235
rect 10057 16133 10091 16167
rect 2881 16065 2915 16099
rect 857 15997 891 16031
rect 2605 15997 2639 16031
rect 5825 15997 5859 16031
rect 6009 15997 6043 16031
rect 6561 15997 6595 16031
rect 6837 15997 6871 16031
rect 7021 15997 7055 16031
rect 7113 15997 7147 16031
rect 7205 15997 7239 16031
rect 7389 15997 7423 16031
rect 7849 15997 7883 16031
rect 8401 15997 8435 16031
rect 8493 15997 8527 16031
rect 8677 15997 8711 16031
rect 8769 15997 8803 16031
rect 9413 15997 9447 16031
rect 10333 15997 10367 16031
rect 11345 15997 11379 16031
rect 11529 15997 11563 16031
rect 11805 15997 11839 16031
rect 12081 15997 12115 16031
rect 1124 15929 1158 15963
rect 7665 15929 7699 15963
rect 9965 15929 9999 15963
rect 10057 15929 10091 15963
rect 2421 15861 2455 15895
rect 6653 15861 6687 15895
rect 7573 15861 7607 15895
rect 9321 15861 9355 15895
rect 9597 15861 9631 15895
rect 9760 15861 9794 15895
rect 10241 15861 10275 15895
rect 11529 15861 11563 15895
rect 1685 15657 1719 15691
rect 1777 15657 1811 15691
rect 3525 15657 3559 15691
rect 3893 15657 3927 15691
rect 7297 15657 7331 15691
rect 8493 15657 8527 15691
rect 8677 15657 8711 15691
rect 10793 15657 10827 15691
rect 11345 15657 11379 15691
rect 12081 15657 12115 15691
rect 3157 15589 3191 15623
rect 10977 15589 11011 15623
rect 1501 15521 1535 15555
rect 1961 15521 1995 15555
rect 2513 15521 2547 15555
rect 2697 15521 2731 15555
rect 2789 15521 2823 15555
rect 3341 15521 3375 15555
rect 4997 15521 5031 15555
rect 5181 15521 5215 15555
rect 5917 15521 5951 15555
rect 6101 15521 6135 15555
rect 6193 15521 6227 15555
rect 6377 15521 6411 15555
rect 6469 15521 6503 15555
rect 7205 15521 7239 15555
rect 7389 15521 7423 15555
rect 7665 15521 7699 15555
rect 7757 15521 7791 15555
rect 7941 15521 7975 15555
rect 8033 15521 8067 15555
rect 8125 15521 8159 15555
rect 8618 15521 8652 15555
rect 9045 15521 9079 15555
rect 9137 15521 9171 15555
rect 9229 15521 9263 15555
rect 9413 15521 9447 15555
rect 10149 15521 10183 15555
rect 11161 15521 11195 15555
rect 11621 15521 11655 15555
rect 12081 15521 12115 15555
rect 12265 15521 12299 15555
rect 1225 15453 1259 15487
rect 2237 15453 2271 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 9597 15453 9631 15487
rect 9873 15453 9907 15487
rect 11713 15453 11747 15487
rect 2145 15385 2179 15419
rect 7481 15385 7515 15419
rect 8309 15385 8343 15419
rect 11989 15385 12023 15419
rect 1317 15317 1351 15351
rect 2329 15317 2363 15351
rect 2973 15317 3007 15351
rect 5089 15317 5123 15351
rect 4261 15113 4295 15147
rect 9413 15113 9447 15147
rect 3249 15045 3283 15079
rect 3893 15045 3927 15079
rect 4813 15045 4847 15079
rect 5641 15045 5675 15079
rect 10517 15045 10551 15079
rect 2237 14977 2271 15011
rect 6101 14977 6135 15011
rect 7481 14977 7515 15011
rect 7573 14977 7607 15011
rect 8401 14977 8435 15011
rect 8677 14977 8711 15011
rect 9781 14977 9815 15011
rect 10149 14977 10183 15011
rect 10609 14977 10643 15011
rect 11713 14977 11747 15011
rect 3525 14909 3559 14943
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 4537 14909 4571 14943
rect 5089 14909 5123 14943
rect 5273 14909 5307 14943
rect 5457 14909 5491 14943
rect 5733 14909 5767 14943
rect 6193 14909 6227 14943
rect 7297 14909 7331 14943
rect 7389 14909 7423 14943
rect 8769 14909 8803 14943
rect 9321 14909 9355 14943
rect 9597 14909 9631 14943
rect 9689 14909 9723 14943
rect 9873 14909 9907 14943
rect 10057 14909 10091 14943
rect 10885 14909 10919 14943
rect 11161 14909 11195 14943
rect 11253 14909 11287 14943
rect 11345 14909 11379 14943
rect 12081 14909 12115 14943
rect 1970 14841 2004 14875
rect 3249 14841 3283 14875
rect 3893 14841 3927 14875
rect 4813 14841 4847 14875
rect 7941 14841 7975 14875
rect 857 14773 891 14807
rect 3433 14773 3467 14807
rect 4077 14773 4111 14807
rect 4445 14773 4479 14807
rect 4997 14773 5031 14807
rect 5365 14773 5399 14807
rect 6561 14773 6595 14807
rect 7113 14773 7147 14807
rect 7849 14773 7883 14807
rect 9137 14773 9171 14807
rect 10701 14773 10735 14807
rect 11069 14773 11103 14807
rect 11437 14773 11471 14807
rect 11897 14773 11931 14807
rect 4445 14569 4479 14603
rect 5825 14569 5859 14603
rect 6469 14569 6503 14603
rect 11621 14569 11655 14603
rect 4261 14501 4295 14535
rect 857 14433 891 14467
rect 1317 14433 1351 14467
rect 1501 14433 1535 14467
rect 1593 14433 1627 14467
rect 2145 14433 2179 14467
rect 2329 14433 2363 14467
rect 2697 14433 2731 14467
rect 3065 14433 3099 14467
rect 3157 14433 3191 14467
rect 3341 14433 3375 14467
rect 3433 14433 3467 14467
rect 3617 14433 3651 14467
rect 4537 14433 4571 14467
rect 5273 14433 5307 14467
rect 6009 14433 6043 14467
rect 6102 14433 6136 14467
rect 6653 14433 6687 14467
rect 6929 14433 6963 14467
rect 7389 14433 7423 14467
rect 7481 14433 7515 14467
rect 7665 14433 7699 14467
rect 8125 14433 8159 14467
rect 8493 14433 8527 14467
rect 8677 14433 8711 14467
rect 9229 14433 9263 14467
rect 9873 14433 9907 14467
rect 10149 14433 10183 14467
rect 10333 14433 10367 14467
rect 11161 14433 11195 14467
rect 11805 14433 11839 14467
rect 11989 14433 12023 14467
rect 12081 14433 12115 14467
rect 2421 14365 2455 14399
rect 2973 14365 3007 14399
rect 4905 14365 4939 14399
rect 5089 14365 5123 14399
rect 5181 14365 5215 14399
rect 5365 14365 5399 14399
rect 6193 14365 6227 14399
rect 6285 14365 6319 14399
rect 7849 14365 7883 14399
rect 8309 14365 8343 14399
rect 8401 14365 8435 14399
rect 8769 14365 8803 14399
rect 8953 14365 8987 14399
rect 9045 14365 9079 14399
rect 9137 14365 9171 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 11253 14365 11287 14399
rect 11529 14365 11563 14399
rect 2513 14297 2547 14331
rect 2881 14297 2915 14331
rect 3433 14297 3467 14331
rect 4261 14297 4295 14331
rect 6745 14297 6779 14331
rect 6837 14297 6871 14331
rect 7941 14297 7975 14331
rect 1961 14229 1995 14263
rect 3341 14229 3375 14263
rect 10333 14229 10367 14263
rect 10609 14229 10643 14263
rect 1593 14025 1627 14059
rect 5549 14025 5583 14059
rect 6101 14025 6135 14059
rect 6837 14025 6871 14059
rect 10149 14025 10183 14059
rect 12081 14025 12115 14059
rect 1961 13957 1995 13991
rect 2697 13957 2731 13991
rect 9965 13957 9999 13991
rect 11805 13957 11839 13991
rect 2605 13889 2639 13923
rect 11069 13889 11103 13923
rect 1777 13821 1811 13855
rect 2053 13821 2087 13855
rect 2145 13821 2179 13855
rect 2329 13821 2363 13855
rect 2513 13821 2547 13855
rect 2973 13821 3007 13855
rect 5181 13821 5215 13855
rect 5733 13821 5767 13855
rect 6561 13821 6595 13855
rect 6837 13821 6871 13855
rect 10517 13821 10551 13855
rect 10701 13821 10735 13855
rect 10793 13821 10827 13855
rect 10885 13821 10919 13855
rect 11161 13821 11195 13855
rect 11897 13821 11931 13855
rect 12081 13821 12115 13855
rect 2697 13753 2731 13787
rect 2881 13753 2915 13787
rect 5365 13753 5399 13787
rect 5917 13753 5951 13787
rect 9689 13753 9723 13787
rect 11437 13753 11471 13787
rect 11621 13753 11655 13787
rect 6653 13685 6687 13719
rect 10701 13685 10735 13719
rect 2421 13481 2455 13515
rect 2789 13481 2823 13515
rect 6561 13481 6595 13515
rect 8953 13481 8987 13515
rect 10977 13481 11011 13515
rect 2605 13413 2639 13447
rect 1970 13345 2004 13379
rect 2329 13345 2363 13379
rect 2697 13345 2731 13379
rect 2881 13345 2915 13379
rect 3801 13345 3835 13379
rect 4813 13345 4847 13379
rect 6469 13345 6503 13379
rect 6745 13345 6779 13379
rect 8861 13345 8895 13379
rect 9137 13345 9171 13379
rect 10977 13345 11011 13379
rect 11161 13345 11195 13379
rect 2237 13277 2271 13311
rect 3893 13277 3927 13311
rect 2605 13209 2639 13243
rect 857 13141 891 13175
rect 4169 13141 4203 13175
rect 4629 13141 4663 13175
rect 6929 13141 6963 13175
rect 9137 13141 9171 13175
rect 2605 12937 2639 12971
rect 6285 12937 6319 12971
rect 9413 12937 9447 12971
rect 9965 12937 9999 12971
rect 5549 12869 5583 12903
rect 6193 12869 6227 12903
rect 7573 12869 7607 12903
rect 8493 12869 8527 12903
rect 11989 12869 12023 12903
rect 1593 12801 1627 12835
rect 2513 12801 2547 12835
rect 5273 12801 5307 12835
rect 5917 12801 5951 12835
rect 7297 12801 7331 12835
rect 7665 12801 7699 12835
rect 8677 12801 8711 12835
rect 9597 12801 9631 12835
rect 11713 12801 11747 12835
rect 1317 12733 1351 12767
rect 1501 12733 1535 12767
rect 2697 12733 2731 12767
rect 2789 12733 2823 12767
rect 4169 12733 4203 12767
rect 4353 12733 4387 12767
rect 4445 12733 4479 12767
rect 4537 12733 4571 12767
rect 5181 12733 5215 12767
rect 5825 12733 5859 12767
rect 6469 12733 6503 12767
rect 6561 12733 6595 12767
rect 6745 12733 6779 12767
rect 6837 12733 6871 12767
rect 7205 12733 7239 12767
rect 7849 12733 7883 12767
rect 7941 12733 7975 12767
rect 8125 12733 8159 12767
rect 8217 12733 8251 12767
rect 8401 12733 8435 12767
rect 8769 12733 8803 12767
rect 8917 12733 8951 12767
rect 9137 12733 9171 12767
rect 9275 12733 9309 12767
rect 9689 12733 9723 12767
rect 11621 12733 11655 12767
rect 857 12665 891 12699
rect 8677 12665 8711 12699
rect 9045 12665 9079 12699
rect 4813 12597 4847 12631
rect 3065 12393 3099 12427
rect 4629 12393 4663 12427
rect 6009 12393 6043 12427
rect 11805 12393 11839 12427
rect 1409 12325 1443 12359
rect 1225 12257 1259 12291
rect 1869 12257 1903 12291
rect 2053 12257 2087 12291
rect 2789 12257 2823 12291
rect 3341 12257 3375 12291
rect 4077 12257 4111 12291
rect 4169 12257 4203 12291
rect 4261 12257 4295 12291
rect 4445 12257 4479 12291
rect 4537 12257 4571 12291
rect 4721 12257 4755 12291
rect 4997 12257 5031 12291
rect 5457 12257 5491 12291
rect 5641 12257 5675 12291
rect 6193 12257 6227 12291
rect 6377 12257 6411 12291
rect 6469 12257 6503 12291
rect 6561 12257 6595 12291
rect 6745 12257 6779 12291
rect 6837 12257 6871 12291
rect 7297 12257 7331 12291
rect 7573 12257 7607 12291
rect 7665 12257 7699 12291
rect 7849 12257 7883 12291
rect 8033 12257 8067 12291
rect 8217 12257 8251 12291
rect 8861 12257 8895 12291
rect 9505 12257 9539 12291
rect 9965 12257 9999 12291
rect 10057 12257 10091 12291
rect 10241 12257 10275 12291
rect 10977 12257 11011 12291
rect 11161 12257 11195 12291
rect 11437 12257 11471 12291
rect 12081 12257 12115 12291
rect 12173 12257 12207 12291
rect 2145 12189 2179 12223
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 3709 12189 3743 12223
rect 5089 12189 5123 12223
rect 7941 12189 7975 12223
rect 8953 12189 8987 12223
rect 9137 12189 9171 12223
rect 9413 12189 9447 12223
rect 11345 12189 11379 12223
rect 11897 12189 11931 12223
rect 3801 12121 3835 12155
rect 5549 12121 5583 12155
rect 9873 12121 9907 12155
rect 1041 12053 1075 12087
rect 2881 12053 2915 12087
rect 5365 12053 5399 12087
rect 7021 12053 7055 12087
rect 7113 12053 7147 12087
rect 7481 12053 7515 12087
rect 8401 12053 8435 12087
rect 8493 12053 8527 12087
rect 10425 12053 10459 12087
rect 11069 12053 11103 12087
rect 11989 12053 12023 12087
rect 2697 11849 2731 11883
rect 6285 11849 6319 11883
rect 7665 11849 7699 11883
rect 8493 11849 8527 11883
rect 8861 11849 8895 11883
rect 9781 11849 9815 11883
rect 11437 11849 11471 11883
rect 11713 11849 11747 11883
rect 5825 11781 5859 11815
rect 4353 11713 4387 11747
rect 4721 11713 4755 11747
rect 5549 11713 5583 11747
rect 6653 11713 6687 11747
rect 8401 11713 8435 11747
rect 10793 11713 10827 11747
rect 1225 11645 1259 11679
rect 1317 11645 1351 11679
rect 3985 11645 4019 11679
rect 4629 11645 4663 11679
rect 4813 11645 4847 11679
rect 4905 11645 4939 11679
rect 5457 11645 5491 11679
rect 6469 11645 6503 11679
rect 6745 11645 6779 11679
rect 6929 11645 6963 11679
rect 7021 11645 7055 11679
rect 7113 11645 7147 11679
rect 7297 11645 7331 11679
rect 7849 11645 7883 11679
rect 8125 11645 8159 11679
rect 8585 11645 8619 11679
rect 8677 11645 8711 11679
rect 8769 11645 8803 11679
rect 8953 11645 8987 11679
rect 9413 11645 9447 11679
rect 9597 11645 9631 11679
rect 9873 11645 9907 11679
rect 10057 11645 10091 11679
rect 10241 11645 10275 11679
rect 10885 11645 10919 11679
rect 11345 11645 11379 11679
rect 11529 11645 11563 11679
rect 11621 11645 11655 11679
rect 11805 11645 11839 11679
rect 1584 11577 1618 11611
rect 4169 11577 4203 11611
rect 10609 11577 10643 11611
rect 1041 11509 1075 11543
rect 4445 11509 4479 11543
rect 7481 11509 7515 11543
rect 8033 11509 8067 11543
rect 9965 11509 9999 11543
rect 10425 11509 10459 11543
rect 11253 11509 11287 11543
rect 5273 11305 5307 11339
rect 6929 11305 6963 11339
rect 7941 11305 7975 11339
rect 9413 11305 9447 11339
rect 1970 11169 2004 11203
rect 2329 11169 2363 11203
rect 5089 11169 5123 11203
rect 5365 11169 5399 11203
rect 6009 11169 6043 11203
rect 6101 11169 6135 11203
rect 6285 11169 6319 11203
rect 6377 11169 6411 11203
rect 6837 11169 6871 11203
rect 7021 11169 7055 11203
rect 7849 11169 7883 11203
rect 8033 11169 8067 11203
rect 9781 11169 9815 11203
rect 10057 11169 10091 11203
rect 10241 11169 10275 11203
rect 10333 11169 10367 11203
rect 10425 11169 10459 11203
rect 11345 11169 11379 11203
rect 2237 11101 2271 11135
rect 9597 11101 9631 11135
rect 9689 11101 9723 11135
rect 9873 11101 9907 11135
rect 10701 11101 10735 11135
rect 11253 11101 11287 11135
rect 857 11033 891 11067
rect 2513 11033 2547 11067
rect 4905 11033 4939 11067
rect 5825 10965 5859 10999
rect 10977 10965 11011 10999
rect 2329 10761 2363 10795
rect 3065 10761 3099 10795
rect 3525 10761 3559 10795
rect 6377 10761 6411 10795
rect 9505 10761 9539 10795
rect 10057 10761 10091 10795
rect 11805 10761 11839 10795
rect 3893 10693 3927 10727
rect 9137 10693 9171 10727
rect 1041 10625 1075 10659
rect 1777 10625 1811 10659
rect 3617 10625 3651 10659
rect 6101 10625 6135 10659
rect 6285 10625 6319 10659
rect 7573 10625 7607 10659
rect 10977 10625 11011 10659
rect 1501 10557 1535 10591
rect 1685 10557 1719 10591
rect 2789 10557 2823 10591
rect 3525 10557 3559 10591
rect 4169 10557 4203 10591
rect 4261 10557 4295 10591
rect 4445 10557 4479 10591
rect 4537 10557 4571 10591
rect 6009 10557 6043 10591
rect 6561 10557 6595 10591
rect 6653 10557 6687 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 7389 10557 7423 10591
rect 7481 10557 7515 10591
rect 7665 10557 7699 10591
rect 9965 10557 9999 10591
rect 10149 10557 10183 10591
rect 10885 10557 10919 10591
rect 11345 10557 11379 10591
rect 11621 10557 11655 10591
rect 2881 10489 2915 10523
rect 3065 10489 3099 10523
rect 7205 10489 7239 10523
rect 8769 10489 8803 10523
rect 9689 10489 9723 10523
rect 9873 10489 9907 10523
rect 3985 10421 4019 10455
rect 6285 10421 6319 10455
rect 7021 10421 7055 10455
rect 9229 10421 9263 10455
rect 11253 10421 11287 10455
rect 11437 10421 11471 10455
rect 8217 10217 8251 10251
rect 9137 10217 9171 10251
rect 9597 10217 9631 10251
rect 1970 10149 2004 10183
rect 5089 10149 5123 10183
rect 9229 10149 9263 10183
rect 11529 10149 11563 10183
rect 3341 10081 3375 10115
rect 3709 10081 3743 10115
rect 4537 10081 4571 10115
rect 4629 10081 4663 10115
rect 4813 10081 4847 10115
rect 4997 10081 5031 10115
rect 5273 10081 5307 10115
rect 7573 10081 7607 10115
rect 7849 10081 7883 10115
rect 8309 10081 8343 10115
rect 8493 10081 8527 10115
rect 8769 10081 8803 10115
rect 9413 10081 9447 10115
rect 9689 10081 9723 10115
rect 9781 10081 9815 10115
rect 9965 10081 9999 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 11713 10081 11747 10115
rect 11897 10081 11931 10115
rect 11989 10081 12023 10115
rect 2237 10013 2271 10047
rect 3985 10013 4019 10047
rect 4721 10013 4755 10047
rect 7757 10013 7791 10047
rect 8401 10013 8435 10047
rect 8677 10013 8711 10047
rect 12173 10013 12207 10047
rect 10977 9945 11011 9979
rect 857 9877 891 9911
rect 4353 9877 4387 9911
rect 5457 9877 5491 9911
rect 6285 9877 6319 9911
rect 9781 9877 9815 9911
rect 12081 9877 12115 9911
rect 7757 9673 7791 9707
rect 8861 9673 8895 9707
rect 10517 9673 10551 9707
rect 12265 9673 12299 9707
rect 3249 9605 3283 9639
rect 3893 9605 3927 9639
rect 6653 9605 6687 9639
rect 7665 9605 7699 9639
rect 1225 9537 1259 9571
rect 1961 9537 1995 9571
rect 2421 9537 2455 9571
rect 3709 9537 3743 9571
rect 4813 9537 4847 9571
rect 5457 9537 5491 9571
rect 5733 9537 5767 9571
rect 6929 9537 6963 9571
rect 8493 9537 8527 9571
rect 9321 9537 9355 9571
rect 10149 9537 10183 9571
rect 1685 9469 1719 9503
rect 1869 9469 1903 9503
rect 2513 9469 2547 9503
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 4353 9469 4387 9503
rect 4721 9469 4755 9503
rect 5365 9469 5399 9503
rect 6285 9469 6319 9503
rect 7021 9469 7055 9503
rect 7297 9469 7331 9503
rect 7451 9469 7485 9503
rect 8033 9469 8067 9503
rect 8585 9469 8619 9503
rect 10057 9469 10091 9503
rect 10609 9469 10643 9503
rect 10885 9469 10919 9503
rect 7757 9401 7791 9435
rect 11152 9401 11186 9435
rect 2881 9333 2915 9367
rect 4261 9333 4295 9367
rect 5089 9333 5123 9367
rect 7941 9333 7975 9367
rect 3893 9129 3927 9163
rect 4353 9129 4387 9163
rect 6653 9129 6687 9163
rect 6929 9129 6963 9163
rect 9137 9129 9171 9163
rect 9505 9129 9539 9163
rect 12173 9129 12207 9163
rect 3801 9061 3835 9095
rect 8769 9061 8803 9095
rect 9781 9061 9815 9095
rect 1869 8993 1903 9027
rect 4261 8993 4295 9027
rect 4629 8993 4663 9027
rect 4721 8993 4755 9027
rect 4905 8993 4939 9027
rect 5641 8993 5675 9027
rect 6285 8993 6319 9027
rect 6561 8993 6595 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 7021 8993 7055 9027
rect 7941 8993 7975 9027
rect 9321 8993 9355 9027
rect 9597 8993 9631 9027
rect 9965 8993 9999 9027
rect 10425 8993 10459 9027
rect 10609 8993 10643 9027
rect 11161 8993 11195 9027
rect 11621 8993 11655 9027
rect 11805 8993 11839 9027
rect 12081 8993 12115 9027
rect 12265 8993 12299 9027
rect 4169 8925 4203 8959
rect 4353 8925 4387 8959
rect 5825 8925 5859 8959
rect 7205 8925 7239 8959
rect 8033 8925 8067 8959
rect 10701 8925 10735 8959
rect 11253 8925 11287 8959
rect 5917 8857 5951 8891
rect 8493 8857 8527 8891
rect 10149 8857 10183 8891
rect 11529 8857 11563 8891
rect 2329 8789 2363 8823
rect 4169 8789 4203 8823
rect 4537 8789 4571 8823
rect 4813 8789 4847 8823
rect 5549 8789 5583 8823
rect 8309 8789 8343 8823
rect 10241 8789 10275 8823
rect 11989 8789 12023 8823
rect 2421 8585 2455 8619
rect 3249 8585 3283 8619
rect 5549 8585 5583 8619
rect 6653 8585 6687 8619
rect 7757 8585 7791 8619
rect 10609 8585 10643 8619
rect 11253 8585 11287 8619
rect 11621 8585 11655 8619
rect 3065 8517 3099 8551
rect 4353 8517 4387 8551
rect 6561 8517 6595 8551
rect 11437 8517 11471 8551
rect 2605 8449 2639 8483
rect 3433 8449 3467 8483
rect 3893 8449 3927 8483
rect 6469 8449 6503 8483
rect 1593 8381 1627 8415
rect 1777 8381 1811 8415
rect 1869 8381 1903 8415
rect 2237 8381 2271 8415
rect 2421 8381 2455 8415
rect 2697 8381 2731 8415
rect 3525 8381 3559 8415
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 4169 8381 4203 8415
rect 4445 8381 4479 8415
rect 4905 8381 4939 8415
rect 4997 8381 5031 8415
rect 5181 8381 5215 8415
rect 5273 8381 5307 8415
rect 5365 8381 5399 8415
rect 5825 8381 5859 8415
rect 6009 8381 6043 8415
rect 6101 8381 6135 8415
rect 6193 8381 6227 8415
rect 6377 8381 6411 8415
rect 6745 8381 6779 8415
rect 7481 8381 7515 8415
rect 7757 8381 7791 8415
rect 9045 8381 9079 8415
rect 9229 8381 9263 8415
rect 9321 8381 9355 8415
rect 9505 8381 9539 8415
rect 10517 8381 10551 8415
rect 10701 8381 10735 8415
rect 10793 8381 10827 8415
rect 10977 8381 11011 8415
rect 1133 8313 1167 8347
rect 5641 8313 5675 8347
rect 7573 8313 7607 8347
rect 9413 8313 9447 8347
rect 11069 8313 11103 8347
rect 11897 8313 11931 8347
rect 9229 8245 9263 8279
rect 10793 8245 10827 8279
rect 11279 8245 11313 8279
rect 857 8041 891 8075
rect 2329 8041 2363 8075
rect 3985 8041 4019 8075
rect 5273 8041 5307 8075
rect 6193 8041 6227 8075
rect 8769 8041 8803 8075
rect 9505 8041 9539 8075
rect 1970 7973 2004 8007
rect 4813 7973 4847 8007
rect 8585 7973 8619 8007
rect 10149 7973 10183 8007
rect 10333 7973 10367 8007
rect 11897 7973 11931 8007
rect 2605 7905 2639 7939
rect 3157 7905 3191 7939
rect 4261 7905 4295 7939
rect 4721 7905 4755 7939
rect 5007 7905 5041 7939
rect 5457 7905 5491 7939
rect 5641 7905 5675 7939
rect 6009 7905 6043 7939
rect 7113 7905 7147 7939
rect 7297 7905 7331 7939
rect 7389 7905 7423 7939
rect 8401 7905 8435 7939
rect 9045 7905 9079 7939
rect 9873 7905 9907 7939
rect 11161 7905 11195 7939
rect 11621 7905 11655 7939
rect 11713 7905 11747 7939
rect 11989 7905 12023 7939
rect 12173 7905 12207 7939
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 3249 7837 3283 7871
rect 4169 7837 4203 7871
rect 5825 7837 5859 7871
rect 9137 7837 9171 7871
rect 9413 7837 9447 7871
rect 9781 7837 9815 7871
rect 11069 7837 11103 7871
rect 11529 7837 11563 7871
rect 11897 7837 11931 7871
rect 2513 7701 2547 7735
rect 4629 7701 4663 7735
rect 4997 7701 5031 7735
rect 6929 7701 6963 7735
rect 11989 7701 12023 7735
rect 2421 7497 2455 7531
rect 2789 7497 2823 7531
rect 7297 7497 7331 7531
rect 8953 7497 8987 7531
rect 12265 7497 12299 7531
rect 4905 7429 4939 7463
rect 5089 7429 5123 7463
rect 5549 7429 5583 7463
rect 9137 7429 9171 7463
rect 4629 7361 4663 7395
rect 7941 7361 7975 7395
rect 8217 7361 8251 7395
rect 8677 7361 8711 7395
rect 9321 7361 9355 7395
rect 10885 7361 10919 7395
rect 2237 7293 2271 7327
rect 2329 7293 2363 7327
rect 2513 7293 2547 7327
rect 2605 7293 2639 7327
rect 2789 7293 2823 7327
rect 5365 7293 5399 7327
rect 5549 7293 5583 7327
rect 5641 7293 5675 7327
rect 5825 7293 5859 7327
rect 6377 7293 6411 7327
rect 6561 7293 6595 7327
rect 6653 7293 6687 7327
rect 6837 7293 6871 7327
rect 6929 7293 6963 7327
rect 7021 7293 7055 7327
rect 7849 7293 7883 7327
rect 8585 7293 8619 7327
rect 9045 7293 9079 7327
rect 11152 7293 11186 7327
rect 1992 7225 2026 7259
rect 5733 7225 5767 7259
rect 857 7157 891 7191
rect 6561 7157 6595 7191
rect 9321 7157 9355 7191
rect 7573 6953 7607 6987
rect 8033 6953 8067 6987
rect 8953 6953 8987 6987
rect 10701 6953 10735 6987
rect 1409 6817 1443 6851
rect 1593 6817 1627 6851
rect 1685 6817 1719 6851
rect 2329 6817 2363 6851
rect 3065 6817 3099 6851
rect 3985 6817 4019 6851
rect 4077 6817 4111 6851
rect 4169 6817 4203 6851
rect 4353 6817 4387 6851
rect 4445 6817 4479 6851
rect 4629 6817 4663 6851
rect 4721 6817 4755 6851
rect 4813 6817 4847 6851
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 5641 6817 5675 6851
rect 6101 6817 6135 6851
rect 6561 6817 6595 6851
rect 7205 6817 7239 6851
rect 7665 6817 7699 6851
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 8309 6817 8343 6851
rect 8493 6817 8527 6851
rect 8677 6817 8711 6851
rect 8769 6817 8803 6851
rect 9045 6817 9079 6851
rect 9597 6817 9631 6851
rect 9781 6817 9815 6851
rect 10057 6817 10091 6851
rect 10241 6817 10275 6851
rect 10517 6817 10551 6851
rect 10793 6817 10827 6851
rect 11345 6817 11379 6851
rect 949 6749 983 6783
rect 2053 6749 2087 6783
rect 3709 6749 3743 6783
rect 5089 6749 5123 6783
rect 5825 6749 5859 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 6929 6749 6963 6783
rect 7113 6749 7147 6783
rect 9873 6749 9907 6783
rect 10977 6749 11011 6783
rect 11253 6749 11287 6783
rect 2237 6681 2271 6715
rect 5181 6681 5215 6715
rect 6009 6681 6043 6715
rect 2145 6613 2179 6647
rect 2973 6613 3007 6647
rect 5917 6613 5951 6647
rect 8769 6613 8803 6647
rect 9689 6613 9723 6647
rect 10333 6613 10367 6647
rect 2513 6409 2547 6443
rect 3065 6409 3099 6443
rect 4629 6409 4663 6443
rect 4905 6409 4939 6443
rect 5641 6409 5675 6443
rect 6837 6409 6871 6443
rect 7021 6409 7055 6443
rect 7205 6409 7239 6443
rect 9505 6409 9539 6443
rect 10701 6409 10735 6443
rect 3525 6273 3559 6307
rect 3801 6273 3835 6307
rect 10333 6273 10367 6307
rect 857 6205 891 6239
rect 1041 6205 1075 6239
rect 1133 6205 1167 6239
rect 2789 6205 2823 6239
rect 3065 6205 3099 6239
rect 3433 6205 3467 6239
rect 4169 6205 4203 6239
rect 4261 6205 4295 6239
rect 4445 6205 4479 6239
rect 4721 6205 4755 6239
rect 4905 6205 4939 6239
rect 5641 6205 5675 6239
rect 5825 6205 5859 6239
rect 6469 6205 6503 6239
rect 6653 6205 6687 6239
rect 6929 6205 6963 6239
rect 7113 6205 7147 6239
rect 7205 6205 7239 6239
rect 7389 6205 7423 6239
rect 9689 6205 9723 6239
rect 9781 6205 9815 6239
rect 10241 6205 10275 6239
rect 949 6137 983 6171
rect 1378 6137 1412 6171
rect 9505 6137 9539 6171
rect 10669 6137 10703 6171
rect 10885 6137 10919 6171
rect 2881 6069 2915 6103
rect 9873 6069 9907 6103
rect 10517 6069 10551 6103
rect 1685 5865 1719 5899
rect 2145 5865 2179 5899
rect 2973 5865 3007 5899
rect 3525 5865 3559 5899
rect 9689 5865 9723 5899
rect 9965 5865 9999 5899
rect 2605 5797 2639 5831
rect 2697 5797 2731 5831
rect 3065 5797 3099 5831
rect 10149 5797 10183 5831
rect 10333 5797 10367 5831
rect 1869 5729 1903 5763
rect 2053 5729 2087 5763
rect 2145 5729 2179 5763
rect 2329 5729 2363 5763
rect 2513 5729 2547 5763
rect 2881 5729 2915 5763
rect 2973 5729 3007 5763
rect 3249 5729 3283 5763
rect 3433 5729 3467 5763
rect 3525 5729 3559 5763
rect 3709 5729 3743 5763
rect 9321 5729 9355 5763
rect 9229 5661 9263 5695
rect 2789 5321 2823 5355
rect 4169 5321 4203 5355
rect 4721 5321 4755 5355
rect 5181 5321 5215 5355
rect 8033 5321 8067 5355
rect 11345 5321 11379 5355
rect 3985 5253 4019 5287
rect 6929 5253 6963 5287
rect 7757 5253 7791 5287
rect 7941 5253 7975 5287
rect 9045 5253 9079 5287
rect 3709 5185 3743 5219
rect 8125 5185 8159 5219
rect 8677 5185 8711 5219
rect 11161 5185 11195 5219
rect 2329 5117 2363 5151
rect 2513 5117 2547 5151
rect 2605 5117 2639 5151
rect 3065 5117 3099 5151
rect 3617 5117 3651 5151
rect 4353 5117 4387 5151
rect 4629 5117 4663 5151
rect 4721 5117 4755 5151
rect 4905 5117 4939 5151
rect 5365 5117 5399 5151
rect 5549 5117 5583 5151
rect 5641 5117 5675 5151
rect 6101 5117 6135 5151
rect 7113 5117 7147 5151
rect 7297 5117 7331 5151
rect 7389 5117 7423 5151
rect 7481 5117 7515 5151
rect 7849 5117 7883 5151
rect 8585 5117 8619 5151
rect 9321 5117 9355 5151
rect 11437 5117 11471 5151
rect 2421 5049 2455 5083
rect 5917 5049 5951 5083
rect 7573 5049 7607 5083
rect 7757 5049 7791 5083
rect 9045 5049 9079 5083
rect 11529 5049 11563 5083
rect 11713 5049 11747 5083
rect 2973 4981 3007 5015
rect 4537 4981 4571 5015
rect 5733 4981 5767 5015
rect 8953 4981 8987 5015
rect 9229 4981 9263 5015
rect 11161 4981 11195 5015
rect 3157 4777 3191 4811
rect 3433 4777 3467 4811
rect 4261 4777 4295 4811
rect 6561 4777 6595 4811
rect 7665 4777 7699 4811
rect 9045 4777 9079 4811
rect 11145 4777 11179 4811
rect 2973 4709 3007 4743
rect 9597 4709 9631 4743
rect 11345 4709 11379 4743
rect 2789 4641 2823 4675
rect 3249 4641 3283 4675
rect 3433 4641 3467 4675
rect 4537 4641 4571 4675
rect 4904 4641 4938 4675
rect 4997 4641 5031 4675
rect 5273 4641 5307 4675
rect 6193 4641 6227 4675
rect 6745 4641 6779 4675
rect 6837 4641 6871 4675
rect 7297 4641 7331 4675
rect 8033 4641 8067 4675
rect 8677 4641 8711 4675
rect 9413 4641 9447 4675
rect 10609 4641 10643 4675
rect 10793 4641 10827 4675
rect 11621 4641 11655 4675
rect 12173 4641 12207 4675
rect 4261 4573 4295 4607
rect 4629 4573 4663 4607
rect 5181 4573 5215 4607
rect 6101 4573 6135 4607
rect 7389 4573 7423 4607
rect 8125 4573 8159 4607
rect 8585 4573 8619 4607
rect 10701 4573 10735 4607
rect 11805 4573 11839 4607
rect 5641 4505 5675 4539
rect 8401 4505 8435 4539
rect 11989 4505 12023 4539
rect 4445 4437 4479 4471
rect 7021 4437 7055 4471
rect 9781 4437 9815 4471
rect 10977 4437 11011 4471
rect 11170 4437 11204 4471
rect 11437 4437 11471 4471
rect 2789 4233 2823 4267
rect 4353 4233 4387 4267
rect 5273 4233 5307 4267
rect 5825 4233 5859 4267
rect 7297 4233 7331 4267
rect 8125 4233 8159 4267
rect 8769 4233 8803 4267
rect 12265 4233 12299 4267
rect 6101 4165 6135 4199
rect 10241 4165 10275 4199
rect 4169 4097 4203 4131
rect 4905 4097 4939 4131
rect 5641 4097 5675 4131
rect 6009 4097 6043 4131
rect 7021 4097 7055 4131
rect 8401 4097 8435 4131
rect 9873 4097 9907 4131
rect 10149 4097 10183 4131
rect 10517 4097 10551 4131
rect 10885 4097 10919 4131
rect 1409 4029 1443 4063
rect 4077 4029 4111 4063
rect 4629 4029 4663 4063
rect 4813 4029 4847 4063
rect 5089 4029 5123 4063
rect 5549 4029 5583 4063
rect 6929 4029 6963 4063
rect 7573 4029 7607 4063
rect 7849 4029 7883 4063
rect 8033 4029 8067 4063
rect 8217 4029 8251 4063
rect 8585 4029 8619 4063
rect 9229 4029 9263 4063
rect 9505 4029 9539 4063
rect 9781 4029 9815 4063
rect 10609 4029 10643 4063
rect 11152 4029 11186 4063
rect 1676 3961 1710 3995
rect 4721 3961 4755 3995
rect 6469 3961 6503 3995
rect 7757 3961 7791 3995
rect 9045 3961 9079 3995
rect 9413 3961 9447 3995
rect 7389 3893 7423 3927
rect 1685 3689 1719 3723
rect 2697 3689 2731 3723
rect 5181 3689 5215 3723
rect 5273 3689 5307 3723
rect 7297 3689 7331 3723
rect 8585 3689 8619 3723
rect 9597 3689 9631 3723
rect 10057 3689 10091 3723
rect 1225 3621 1259 3655
rect 1441 3621 1475 3655
rect 1869 3621 1903 3655
rect 2329 3621 2363 3655
rect 3525 3621 3559 3655
rect 7205 3621 7239 3655
rect 11345 3621 11379 3655
rect 11621 3621 11655 3655
rect 11989 3621 12023 3655
rect 2513 3553 2547 3587
rect 2789 3553 2823 3587
rect 3341 3553 3375 3587
rect 3801 3553 3835 3587
rect 4261 3553 4295 3587
rect 4445 3553 4479 3587
rect 4629 3553 4663 3587
rect 4721 3553 4755 3587
rect 4813 3553 4847 3587
rect 4906 3553 4940 3587
rect 5273 3553 5307 3587
rect 5457 3553 5491 3587
rect 6837 3553 6871 3587
rect 7021 3553 7055 3587
rect 7572 3553 7606 3587
rect 7665 3553 7699 3587
rect 8493 3553 8527 3587
rect 8677 3553 8711 3587
rect 8769 3553 8803 3587
rect 8953 3553 8987 3587
rect 9321 3553 9355 3587
rect 9413 3553 9447 3587
rect 9689 3553 9723 3587
rect 9782 3553 9816 3587
rect 11805 3553 11839 3587
rect 2237 3485 2271 3519
rect 3157 3485 3191 3519
rect 3709 3485 3743 3519
rect 8861 3485 8895 3519
rect 1593 3417 1627 3451
rect 10977 3417 11011 3451
rect 1409 3349 1443 3383
rect 1869 3349 1903 3383
rect 4077 3349 4111 3383
rect 11345 3349 11379 3383
rect 11529 3349 11563 3383
rect 4537 3145 4571 3179
rect 12265 3145 12299 3179
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 2421 3009 2455 3043
rect 2881 3009 2915 3043
rect 10885 3009 10919 3043
rect 1869 2941 1903 2975
rect 2513 2941 2547 2975
rect 4169 2941 4203 2975
rect 6561 2941 6595 2975
rect 6745 2941 6779 2975
rect 11152 2941 11186 2975
rect 4353 2873 4387 2907
rect 6653 2805 6687 2839
rect 3525 2601 3559 2635
rect 6837 2601 6871 2635
rect 7465 2601 7499 2635
rect 10333 2601 10367 2635
rect 6009 2533 6043 2567
rect 7665 2533 7699 2567
rect 9229 2533 9263 2567
rect 2513 2465 2547 2499
rect 3157 2465 3191 2499
rect 5825 2465 5859 2499
rect 6469 2465 6503 2499
rect 7021 2465 7055 2499
rect 7205 2465 7239 2499
rect 8033 2465 8067 2499
rect 8677 2465 8711 2499
rect 8861 2465 8895 2499
rect 9137 2465 9171 2499
rect 9321 2465 9355 2499
rect 9505 2465 9539 2499
rect 9965 2465 9999 2499
rect 10609 2465 10643 2499
rect 2421 2397 2455 2431
rect 3065 2397 3099 2431
rect 6561 2397 6595 2431
rect 7757 2397 7791 2431
rect 10057 2397 10091 2431
rect 2881 2329 2915 2363
rect 7297 2329 7331 2363
rect 10425 2329 10459 2363
rect 6193 2261 6227 2295
rect 7205 2261 7239 2295
rect 7481 2261 7515 2295
rect 8677 2261 8711 2295
rect 9597 2261 9631 2295
rect 3249 2057 3283 2091
rect 3985 2057 4019 2091
rect 8217 2057 8251 2091
rect 9781 2057 9815 2091
rect 2605 1989 2639 2023
rect 4905 1989 4939 2023
rect 5549 1989 5583 2023
rect 2513 1921 2547 1955
rect 3709 1921 3743 1955
rect 4445 1921 4479 1955
rect 5089 1921 5123 1955
rect 5641 1921 5675 1955
rect 2237 1853 2271 1887
rect 2329 1853 2363 1887
rect 2881 1853 2915 1887
rect 3433 1853 3467 1887
rect 3617 1853 3651 1887
rect 3801 1853 3835 1887
rect 4537 1853 4571 1887
rect 5181 1853 5215 1887
rect 5825 1853 5859 1887
rect 6009 1853 6043 1887
rect 6285 1853 6319 1887
rect 6561 1853 6595 1887
rect 6745 1853 6779 1887
rect 6837 1853 6871 1887
rect 8401 1853 8435 1887
rect 10057 1853 10091 1887
rect 10333 1853 10367 1887
rect 10517 1853 10551 1887
rect 10793 1853 10827 1887
rect 10977 1853 11011 1887
rect 11069 1853 11103 1887
rect 11253 1853 11287 1887
rect 2513 1785 2547 1819
rect 2605 1785 2639 1819
rect 7104 1785 7138 1819
rect 8668 1785 8702 1819
rect 11161 1785 11195 1819
rect 2789 1717 2823 1751
rect 6101 1717 6135 1751
rect 9873 1717 9907 1751
rect 10609 1717 10643 1751
rect 3157 1513 3191 1547
rect 5273 1513 5307 1547
rect 7389 1513 7423 1547
rect 8125 1513 8159 1547
rect 8401 1513 8435 1547
rect 8585 1513 8619 1547
rect 9321 1513 9355 1547
rect 10425 1513 10459 1547
rect 10609 1513 10643 1547
rect 2044 1445 2078 1479
rect 3617 1377 3651 1411
rect 4261 1377 4295 1411
rect 4905 1377 4939 1411
rect 5457 1367 5491 1401
rect 5641 1377 5675 1411
rect 6009 1377 6043 1411
rect 6285 1377 6319 1411
rect 6745 1377 6779 1411
rect 7573 1377 7607 1411
rect 7665 1377 7699 1411
rect 7941 1377 7975 1411
rect 8217 1377 8251 1411
rect 8861 1377 8895 1411
rect 9137 1377 9171 1411
rect 9597 1377 9631 1411
rect 10057 1377 10091 1411
rect 10241 1377 10275 1411
rect 10517 1377 10551 1411
rect 10609 1377 10643 1411
rect 10793 1377 10827 1411
rect 1777 1309 1811 1343
rect 3709 1309 3743 1343
rect 4169 1309 4203 1343
rect 4629 1309 4663 1343
rect 4813 1309 4847 1343
rect 6193 1309 6227 1343
rect 6837 1309 6871 1343
rect 7389 1309 7423 1343
rect 7757 1309 7791 1343
rect 8585 1309 8619 1343
rect 8953 1309 8987 1343
rect 9689 1309 9723 1343
rect 5825 1241 5859 1275
rect 8769 1241 8803 1275
rect 3985 1173 4019 1207
rect 5549 1173 5583 1207
rect 7021 1173 7055 1207
rect 9873 1173 9907 1207
rect 3801 969 3835 1003
rect 6193 969 6227 1003
rect 6653 969 6687 1003
rect 9597 969 9631 1003
rect 4077 833 4111 867
rect 3249 765 3283 799
rect 3617 765 3651 799
rect 3709 765 3743 799
rect 3893 765 3927 799
rect 3985 765 4019 799
rect 4169 765 4203 799
rect 6101 765 6135 799
rect 6285 765 6319 799
rect 6653 765 6687 799
rect 6837 765 6871 799
rect 9413 765 9447 799
rect 9597 765 9631 799
rect 3433 697 3467 731
<< metal1 >>
rect 7190 43324 7196 43376
rect 7248 43364 7254 43376
rect 10042 43364 10048 43376
rect 7248 43336 10048 43364
rect 7248 43324 7254 43336
rect 10042 43324 10048 43336
rect 10100 43324 10106 43376
rect 2958 43120 2964 43172
rect 3016 43160 3022 43172
rect 8662 43160 8668 43172
rect 3016 43132 8668 43160
rect 3016 43120 3022 43132
rect 8662 43120 8668 43132
rect 8720 43120 8726 43172
rect 7466 43052 7472 43104
rect 7524 43092 7530 43104
rect 9950 43092 9956 43104
rect 7524 43064 9956 43092
rect 7524 43052 7530 43064
rect 9950 43052 9956 43064
rect 10008 43052 10014 43104
rect 552 43002 12604 43024
rect 552 42950 4322 43002
rect 4374 42950 4386 43002
rect 4438 42950 4450 43002
rect 4502 42950 4514 43002
rect 4566 42950 4578 43002
rect 4630 42950 10722 43002
rect 10774 42950 10786 43002
rect 10838 42950 10850 43002
rect 10902 42950 10914 43002
rect 10966 42950 10978 43002
rect 11030 42950 12604 43002
rect 552 42928 12604 42950
rect 8294 42888 8300 42900
rect 2976 42860 8300 42888
rect 2976 42829 3004 42860
rect 8294 42848 8300 42860
rect 8352 42848 8358 42900
rect 8772 42860 12020 42888
rect 2961 42823 3019 42829
rect 2961 42789 2973 42823
rect 3007 42789 3019 42823
rect 2961 42783 3019 42789
rect 3605 42823 3663 42829
rect 3605 42789 3617 42823
rect 3651 42820 3663 42823
rect 6638 42820 6644 42832
rect 3651 42792 6644 42820
rect 3651 42789 3663 42792
rect 3605 42783 3663 42789
rect 6638 42780 6644 42792
rect 6696 42780 6702 42832
rect 7561 42823 7619 42829
rect 7561 42820 7573 42823
rect 6748 42792 7573 42820
rect 14 42712 20 42764
rect 72 42752 78 42764
rect 1121 42755 1179 42761
rect 1121 42752 1133 42755
rect 72 42724 1133 42752
rect 72 42712 78 42724
rect 1121 42721 1133 42724
rect 1167 42721 1179 42755
rect 1121 42715 1179 42721
rect 1213 42755 1271 42761
rect 1213 42721 1225 42755
rect 1259 42752 1271 42755
rect 1302 42752 1308 42764
rect 1259 42724 1308 42752
rect 1259 42721 1271 42724
rect 1213 42715 1271 42721
rect 1302 42712 1308 42724
rect 1360 42712 1366 42764
rect 1486 42761 1492 42764
rect 1480 42715 1492 42761
rect 1486 42712 1492 42715
rect 1544 42712 1550 42764
rect 4246 42712 4252 42764
rect 4304 42752 4310 42764
rect 4525 42755 4583 42761
rect 4525 42752 4537 42755
rect 4304 42724 4537 42752
rect 4304 42712 4310 42724
rect 4525 42721 4537 42724
rect 4571 42721 4583 42755
rect 4525 42715 4583 42721
rect 5350 42712 5356 42764
rect 5408 42752 5414 42764
rect 5445 42755 5503 42761
rect 5445 42752 5457 42755
rect 5408 42724 5457 42752
rect 5408 42712 5414 42724
rect 5445 42721 5457 42724
rect 5491 42721 5503 42755
rect 5445 42715 5503 42721
rect 5629 42755 5687 42761
rect 5629 42721 5641 42755
rect 5675 42752 5687 42755
rect 6178 42752 6184 42764
rect 5675 42724 6184 42752
rect 5675 42721 5687 42724
rect 5629 42715 5687 42721
rect 6178 42712 6184 42724
rect 6236 42712 6242 42764
rect 6270 42712 6276 42764
rect 6328 42752 6334 42764
rect 6748 42752 6776 42792
rect 7561 42789 7573 42792
rect 7607 42789 7619 42823
rect 7561 42783 7619 42789
rect 7653 42823 7711 42829
rect 7653 42789 7665 42823
rect 7699 42820 7711 42823
rect 7742 42820 7748 42832
rect 7699 42792 7748 42820
rect 7699 42789 7711 42792
rect 7653 42783 7711 42789
rect 7742 42780 7748 42792
rect 7800 42780 7806 42832
rect 8772 42829 8800 42860
rect 8757 42823 8815 42829
rect 7852 42792 8616 42820
rect 7466 42761 7472 42764
rect 7464 42752 7472 42761
rect 6328 42724 6776 42752
rect 7427 42724 7472 42752
rect 6328 42712 6334 42724
rect 7464 42715 7472 42724
rect 7466 42712 7472 42715
rect 7524 42712 7530 42764
rect 7852 42761 7880 42792
rect 7836 42755 7894 42761
rect 7836 42721 7848 42755
rect 7882 42721 7894 42755
rect 7836 42715 7894 42721
rect 7926 42712 7932 42764
rect 7984 42712 7990 42764
rect 8018 42712 8024 42764
rect 8076 42712 8082 42764
rect 8205 42755 8263 42761
rect 8205 42721 8217 42755
rect 8251 42721 8263 42755
rect 8205 42715 8263 42721
rect 8389 42755 8447 42761
rect 8389 42721 8401 42755
rect 8435 42721 8447 42755
rect 8389 42715 8447 42721
rect 4433 42687 4491 42693
rect 4433 42653 4445 42687
rect 4479 42653 4491 42687
rect 4433 42647 4491 42653
rect 4801 42687 4859 42693
rect 4801 42653 4813 42687
rect 4847 42684 4859 42687
rect 4890 42684 4896 42696
rect 4847 42656 4896 42684
rect 4847 42653 4859 42656
rect 4801 42647 4859 42653
rect 3142 42576 3148 42628
rect 3200 42616 3206 42628
rect 3421 42619 3479 42625
rect 3421 42616 3433 42619
rect 3200 42588 3433 42616
rect 3200 42576 3206 42588
rect 3421 42585 3433 42588
rect 3467 42585 3479 42619
rect 4448 42616 4476 42647
rect 4890 42644 4896 42656
rect 4948 42644 4954 42696
rect 5258 42644 5264 42696
rect 5316 42684 5322 42696
rect 6365 42687 6423 42693
rect 6365 42684 6377 42687
rect 5316 42656 6377 42684
rect 5316 42644 5322 42656
rect 6365 42653 6377 42656
rect 6411 42653 6423 42687
rect 6365 42647 6423 42653
rect 7193 42687 7251 42693
rect 7193 42653 7205 42687
rect 7239 42684 7251 42687
rect 7282 42684 7288 42696
rect 7239 42656 7288 42684
rect 7239 42653 7251 42656
rect 7193 42647 7251 42653
rect 7282 42644 7288 42656
rect 7340 42644 7346 42696
rect 8110 42644 8116 42696
rect 8168 42684 8174 42696
rect 8220 42684 8248 42715
rect 8168 42656 8248 42684
rect 8168 42644 8174 42656
rect 8294 42644 8300 42696
rect 8352 42684 8358 42696
rect 8404 42684 8432 42715
rect 8478 42712 8484 42764
rect 8536 42712 8542 42764
rect 8352 42656 8432 42684
rect 8588 42684 8616 42792
rect 8757 42789 8769 42823
rect 8803 42789 8815 42823
rect 9030 42820 9036 42832
rect 8757 42783 8815 42789
rect 8869 42792 9036 42820
rect 8662 42712 8668 42764
rect 8720 42712 8726 42764
rect 8869 42761 8897 42792
rect 9030 42780 9036 42792
rect 9088 42780 9094 42832
rect 11698 42820 11704 42832
rect 11348 42792 11704 42820
rect 8854 42755 8912 42761
rect 8854 42721 8866 42755
rect 8900 42721 8912 42755
rect 9125 42755 9183 42761
rect 9125 42752 9137 42755
rect 8854 42715 8912 42721
rect 8956 42724 9137 42752
rect 8956 42684 8984 42724
rect 9125 42721 9137 42724
rect 9171 42721 9183 42755
rect 9125 42715 9183 42721
rect 10042 42712 10048 42764
rect 10100 42712 10106 42764
rect 10505 42755 10563 42761
rect 10505 42721 10517 42755
rect 10551 42752 10563 42755
rect 10778 42752 10784 42764
rect 10551 42724 10784 42752
rect 10551 42721 10563 42724
rect 10505 42715 10563 42721
rect 10778 42712 10784 42724
rect 10836 42712 10842 42764
rect 11057 42755 11115 42761
rect 11057 42721 11069 42755
rect 11103 42752 11115 42755
rect 11146 42752 11152 42764
rect 11103 42724 11152 42752
rect 11103 42721 11115 42724
rect 11057 42715 11115 42721
rect 11146 42712 11152 42724
rect 11204 42712 11210 42764
rect 11348 42761 11376 42792
rect 11698 42780 11704 42792
rect 11756 42780 11762 42832
rect 11333 42755 11391 42761
rect 11333 42721 11345 42755
rect 11379 42721 11391 42755
rect 11333 42715 11391 42721
rect 11425 42755 11483 42761
rect 11425 42721 11437 42755
rect 11471 42721 11483 42755
rect 11425 42715 11483 42721
rect 11609 42755 11667 42761
rect 11609 42721 11621 42755
rect 11655 42721 11667 42755
rect 11609 42715 11667 42721
rect 8588 42656 8984 42684
rect 8352 42644 8358 42656
rect 9674 42644 9680 42696
rect 9732 42644 9738 42696
rect 9766 42644 9772 42696
rect 9824 42684 9830 42696
rect 10229 42687 10287 42693
rect 10229 42684 10241 42687
rect 9824 42656 10241 42684
rect 9824 42644 9830 42656
rect 10229 42653 10241 42656
rect 10275 42653 10287 42687
rect 10229 42647 10287 42653
rect 10321 42687 10379 42693
rect 10321 42653 10333 42687
rect 10367 42653 10379 42687
rect 11440 42684 11468 42715
rect 10321 42647 10379 42653
rect 11256 42656 11468 42684
rect 4448 42588 7328 42616
rect 3421 42579 3479 42585
rect 934 42508 940 42560
rect 992 42508 998 42560
rect 2590 42508 2596 42560
rect 2648 42508 2654 42560
rect 2866 42508 2872 42560
rect 2924 42508 2930 42560
rect 3789 42551 3847 42557
rect 3789 42517 3801 42551
rect 3835 42548 3847 42551
rect 4062 42548 4068 42560
rect 3835 42520 4068 42548
rect 3835 42517 3847 42520
rect 3789 42511 3847 42517
rect 4062 42508 4068 42520
rect 4120 42508 4126 42560
rect 5626 42508 5632 42560
rect 5684 42508 5690 42560
rect 5810 42508 5816 42560
rect 5868 42508 5874 42560
rect 6546 42508 6552 42560
rect 6604 42508 6610 42560
rect 7300 42557 7328 42588
rect 9398 42576 9404 42628
rect 9456 42616 9462 42628
rect 10336 42616 10364 42647
rect 11256 42628 11284 42656
rect 9456 42588 10364 42616
rect 9456 42576 9462 42588
rect 10870 42576 10876 42628
rect 10928 42616 10934 42628
rect 10928 42588 11192 42616
rect 10928 42576 10934 42588
rect 7285 42551 7343 42557
rect 7285 42517 7297 42551
rect 7331 42517 7343 42551
rect 7285 42511 7343 42517
rect 8202 42508 8208 42560
rect 8260 42508 8266 42560
rect 8386 42508 8392 42560
rect 8444 42548 8450 42560
rect 9033 42551 9091 42557
rect 9033 42548 9045 42551
rect 8444 42520 9045 42548
rect 8444 42508 8450 42520
rect 9033 42517 9045 42520
rect 9079 42517 9091 42551
rect 9033 42511 9091 42517
rect 9122 42508 9128 42560
rect 9180 42548 9186 42560
rect 9861 42551 9919 42557
rect 9861 42548 9873 42551
rect 9180 42520 9873 42548
rect 9180 42508 9186 42520
rect 9861 42517 9873 42520
rect 9907 42517 9919 42551
rect 9861 42511 9919 42517
rect 10689 42551 10747 42557
rect 10689 42517 10701 42551
rect 10735 42548 10747 42551
rect 10962 42548 10968 42560
rect 10735 42520 10968 42548
rect 10735 42517 10747 42520
rect 10689 42511 10747 42517
rect 10962 42508 10968 42520
rect 11020 42508 11026 42560
rect 11164 42548 11192 42588
rect 11238 42576 11244 42628
rect 11296 42576 11302 42628
rect 11624 42548 11652 42715
rect 11992 42693 12020 42860
rect 12066 42712 12072 42764
rect 12124 42752 12130 42764
rect 12253 42755 12311 42761
rect 12253 42752 12265 42755
rect 12124 42724 12265 42752
rect 12124 42712 12130 42724
rect 12253 42721 12265 42724
rect 12299 42721 12311 42755
rect 12253 42715 12311 42721
rect 11977 42687 12035 42693
rect 11977 42653 11989 42687
rect 12023 42684 12035 42687
rect 12158 42684 12164 42696
rect 12023 42656 12164 42684
rect 12023 42653 12035 42656
rect 11977 42647 12035 42653
rect 12158 42644 12164 42656
rect 12216 42644 12222 42696
rect 11164 42520 11652 42548
rect 11790 42508 11796 42560
rect 11848 42508 11854 42560
rect 11882 42508 11888 42560
rect 11940 42548 11946 42560
rect 12069 42551 12127 42557
rect 12069 42548 12081 42551
rect 11940 42520 12081 42548
rect 11940 42508 11946 42520
rect 12069 42517 12081 42520
rect 12115 42517 12127 42551
rect 12069 42511 12127 42517
rect 12161 42551 12219 42557
rect 12161 42517 12173 42551
rect 12207 42548 12219 42551
rect 12434 42548 12440 42560
rect 12207 42520 12440 42548
rect 12207 42517 12219 42520
rect 12161 42511 12219 42517
rect 12434 42508 12440 42520
rect 12492 42508 12498 42560
rect 552 42458 12604 42480
rect 552 42406 3662 42458
rect 3714 42406 3726 42458
rect 3778 42406 3790 42458
rect 3842 42406 3854 42458
rect 3906 42406 3918 42458
rect 3970 42406 10062 42458
rect 10114 42406 10126 42458
rect 10178 42406 10190 42458
rect 10242 42406 10254 42458
rect 10306 42406 10318 42458
rect 10370 42406 12604 42458
rect 552 42384 12604 42406
rect 1228 42316 2535 42344
rect 842 42100 848 42152
rect 900 42100 906 42152
rect 1026 42149 1032 42152
rect 993 42143 1032 42149
rect 993 42109 1005 42143
rect 993 42103 1032 42109
rect 1026 42100 1032 42103
rect 1084 42100 1090 42152
rect 1121 42143 1179 42149
rect 1121 42109 1133 42143
rect 1167 42140 1179 42143
rect 1228 42140 1256 42316
rect 2507 42276 2535 42316
rect 2958 42304 2964 42356
rect 3016 42304 3022 42356
rect 4154 42344 4160 42356
rect 3068 42316 4160 42344
rect 3068 42276 3096 42316
rect 4154 42304 4160 42316
rect 4212 42304 4218 42356
rect 5258 42304 5264 42356
rect 5316 42304 5322 42356
rect 5350 42304 5356 42356
rect 5408 42344 5414 42356
rect 5718 42344 5724 42356
rect 5408 42316 5724 42344
rect 5408 42304 5414 42316
rect 5718 42304 5724 42316
rect 5776 42304 5782 42356
rect 6914 42304 6920 42356
rect 6972 42344 6978 42356
rect 8386 42344 8392 42356
rect 6972 42316 8392 42344
rect 6972 42304 6978 42316
rect 8386 42304 8392 42316
rect 8444 42304 8450 42356
rect 8665 42347 8723 42353
rect 8665 42313 8677 42347
rect 8711 42344 8723 42347
rect 9122 42344 9128 42356
rect 8711 42316 9128 42344
rect 8711 42313 8723 42316
rect 8665 42307 8723 42313
rect 9122 42304 9128 42316
rect 9180 42304 9186 42356
rect 2507 42248 3096 42276
rect 3786 42236 3792 42288
rect 3844 42276 3850 42288
rect 7834 42285 7840 42288
rect 4893 42279 4951 42285
rect 4893 42276 4905 42279
rect 3844 42248 4905 42276
rect 3844 42236 3850 42248
rect 4893 42245 4905 42248
rect 4939 42245 4951 42279
rect 4893 42239 4951 42245
rect 7833 42239 7840 42285
rect 7892 42276 7898 42288
rect 7892 42248 9720 42276
rect 4246 42208 4252 42220
rect 4080 42180 4252 42208
rect 1167 42112 1256 42140
rect 1351 42143 1409 42149
rect 1167 42109 1179 42112
rect 1121 42103 1179 42109
rect 1351 42109 1363 42143
rect 1397 42140 1409 42143
rect 1397 42112 1532 42140
rect 1397 42109 1409 42112
rect 1351 42103 1409 42109
rect 1210 42032 1216 42084
rect 1268 42032 1274 42084
rect 1504 42072 1532 42112
rect 1578 42100 1584 42152
rect 1636 42100 1642 42152
rect 2130 42140 2136 42152
rect 1780 42112 2136 42140
rect 1780 42072 1808 42112
rect 2130 42100 2136 42112
rect 2188 42100 2194 42152
rect 3421 42143 3479 42149
rect 3421 42109 3433 42143
rect 3467 42140 3479 42143
rect 3970 42140 3976 42152
rect 3467 42112 3976 42140
rect 3467 42109 3479 42112
rect 3421 42103 3479 42109
rect 3970 42100 3976 42112
rect 4028 42100 4034 42152
rect 4080 42149 4108 42180
rect 4246 42168 4252 42180
rect 4304 42168 4310 42220
rect 4908 42208 4936 42239
rect 7834 42236 7840 42239
rect 7892 42236 7898 42248
rect 8481 42211 8539 42217
rect 8481 42208 8493 42211
rect 4448 42180 4752 42208
rect 4908 42180 5488 42208
rect 4065 42143 4123 42149
rect 4065 42109 4077 42143
rect 4111 42109 4123 42143
rect 4065 42103 4123 42109
rect 4154 42100 4160 42152
rect 4212 42140 4218 42152
rect 4212 42112 4257 42140
rect 4212 42100 4218 42112
rect 4338 42100 4344 42152
rect 4396 42100 4402 42152
rect 4448 42149 4476 42180
rect 4433 42143 4491 42149
rect 4433 42109 4445 42143
rect 4479 42109 4491 42143
rect 4433 42103 4491 42109
rect 4530 42143 4588 42149
rect 4530 42109 4542 42143
rect 4576 42140 4588 42143
rect 4576 42112 4660 42140
rect 4576 42109 4588 42112
rect 4530 42103 4588 42109
rect 1854 42081 1860 42084
rect 1504 42044 1808 42072
rect 1848 42035 1860 42081
rect 1854 42032 1860 42035
rect 1912 42032 1918 42084
rect 3142 42032 3148 42084
rect 3200 42072 3206 42084
rect 3200 42044 4476 42072
rect 3200 42032 3206 42044
rect 1489 42007 1547 42013
rect 1489 41973 1501 42007
rect 1535 42004 1547 42007
rect 2866 42004 2872 42016
rect 1535 41976 2872 42004
rect 1535 41973 1547 41976
rect 1489 41967 1547 41973
rect 2866 41964 2872 41976
rect 2924 41964 2930 42016
rect 3973 42007 4031 42013
rect 3973 41973 3985 42007
rect 4019 42004 4031 42007
rect 4154 42004 4160 42016
rect 4019 41976 4160 42004
rect 4019 41973 4031 41976
rect 3973 41967 4031 41973
rect 4154 41964 4160 41976
rect 4212 41964 4218 42016
rect 4448 42004 4476 42044
rect 4632 42004 4660 42112
rect 4724 42072 4752 42180
rect 4798 42100 4804 42152
rect 4856 42100 4862 42152
rect 5074 42100 5080 42152
rect 5132 42100 5138 42152
rect 5166 42100 5172 42152
rect 5224 42140 5230 42152
rect 5353 42143 5411 42149
rect 5353 42140 5365 42143
rect 5224 42112 5365 42140
rect 5224 42100 5230 42112
rect 5353 42109 5365 42112
rect 5399 42109 5411 42143
rect 5353 42103 5411 42109
rect 5258 42072 5264 42084
rect 4724 42044 5264 42072
rect 5258 42032 5264 42044
rect 5316 42032 5322 42084
rect 5460 42072 5488 42180
rect 7760 42180 8493 42208
rect 7760 42152 7788 42180
rect 8481 42177 8493 42180
rect 8527 42208 8539 42211
rect 8527 42180 9536 42208
rect 8527 42177 8539 42180
rect 8481 42171 8539 42177
rect 5620 42143 5678 42149
rect 5620 42109 5632 42143
rect 5666 42140 5678 42143
rect 6546 42140 6552 42152
rect 5666 42112 6552 42140
rect 5666 42109 5678 42112
rect 5620 42103 5678 42109
rect 6546 42100 6552 42112
rect 6604 42100 6610 42152
rect 6917 42143 6975 42149
rect 6917 42109 6929 42143
rect 6963 42140 6975 42143
rect 7190 42140 7196 42152
rect 6963 42112 7196 42140
rect 6963 42109 6975 42112
rect 6917 42103 6975 42109
rect 6822 42072 6828 42084
rect 5460 42044 6828 42072
rect 6822 42032 6828 42044
rect 6880 42032 6886 42084
rect 4448 41976 4660 42004
rect 4709 42007 4767 42013
rect 4709 41973 4721 42007
rect 4755 42004 4767 42007
rect 5442 42004 5448 42016
rect 4755 41976 5448 42004
rect 4755 41973 4767 41976
rect 4709 41967 4767 41973
rect 5442 41964 5448 41976
rect 5500 41964 5506 42016
rect 6454 41964 6460 42016
rect 6512 42004 6518 42016
rect 6733 42007 6791 42013
rect 6733 42004 6745 42007
rect 6512 41976 6745 42004
rect 6512 41964 6518 41976
rect 6733 41973 6745 41976
rect 6779 42004 6791 42007
rect 6932 42004 6960 42103
rect 7190 42100 7196 42112
rect 7248 42100 7254 42152
rect 7466 42100 7472 42152
rect 7524 42140 7530 42152
rect 7653 42143 7711 42149
rect 7653 42140 7665 42143
rect 7524 42112 7665 42140
rect 7524 42100 7530 42112
rect 7653 42109 7665 42112
rect 7699 42109 7711 42143
rect 7653 42103 7711 42109
rect 7742 42100 7748 42152
rect 7800 42100 7806 42152
rect 7926 42100 7932 42152
rect 7984 42140 7990 42152
rect 8110 42140 8116 42152
rect 7984 42112 8116 42140
rect 7984 42100 7990 42112
rect 8110 42100 8116 42112
rect 8168 42100 8174 42152
rect 8386 42100 8392 42152
rect 8444 42140 8450 42152
rect 8573 42143 8631 42149
rect 8573 42140 8585 42143
rect 8444 42112 8585 42140
rect 8444 42100 8450 42112
rect 8573 42109 8585 42112
rect 8619 42109 8631 42143
rect 8573 42103 8631 42109
rect 8754 42100 8760 42152
rect 8812 42140 8818 42152
rect 9125 42143 9183 42149
rect 9125 42140 9137 42143
rect 8812 42112 9137 42140
rect 8812 42100 8818 42112
rect 9125 42109 9137 42112
rect 9171 42109 9183 42143
rect 9125 42103 9183 42109
rect 9214 42100 9220 42152
rect 9272 42140 9278 42152
rect 9508 42149 9536 42180
rect 9692 42149 9720 42248
rect 9766 42236 9772 42288
rect 9824 42276 9830 42288
rect 10870 42276 10876 42288
rect 9824 42248 10876 42276
rect 9824 42236 9830 42248
rect 10870 42236 10876 42248
rect 10928 42236 10934 42288
rect 9309 42143 9367 42149
rect 9309 42140 9321 42143
rect 9272 42112 9321 42140
rect 9272 42100 9278 42112
rect 9309 42109 9321 42112
rect 9355 42109 9367 42143
rect 9309 42103 9367 42109
rect 9493 42143 9551 42149
rect 9493 42109 9505 42143
rect 9539 42109 9551 42143
rect 9493 42103 9551 42109
rect 9677 42143 9735 42149
rect 9677 42109 9689 42143
rect 9723 42109 9735 42143
rect 9677 42103 9735 42109
rect 9950 42100 9956 42152
rect 10008 42140 10014 42152
rect 10137 42143 10195 42149
rect 10137 42140 10149 42143
rect 10008 42112 10149 42140
rect 10008 42100 10014 42112
rect 10137 42109 10149 42112
rect 10183 42109 10195 42143
rect 10137 42103 10195 42109
rect 10594 42100 10600 42152
rect 10652 42140 10658 42152
rect 12250 42140 12256 42152
rect 10652 42112 12256 42140
rect 10652 42100 10658 42112
rect 12250 42100 12256 42112
rect 12308 42100 12314 42152
rect 7006 42032 7012 42084
rect 7064 42072 7070 42084
rect 8018 42072 8024 42084
rect 7064 42044 8024 42072
rect 7064 42032 7070 42044
rect 8018 42032 8024 42044
rect 8076 42032 8082 42084
rect 8846 42032 8852 42084
rect 8904 42032 8910 42084
rect 8938 42032 8944 42084
rect 8996 42032 9002 42084
rect 9033 42075 9091 42081
rect 9033 42041 9045 42075
rect 9079 42041 9091 42075
rect 9033 42035 9091 42041
rect 6779 41976 6960 42004
rect 7469 42007 7527 42013
rect 6779 41973 6791 41976
rect 6733 41967 6791 41973
rect 7469 41973 7481 42007
rect 7515 42004 7527 42007
rect 7558 42004 7564 42016
rect 7515 41976 7564 42004
rect 7515 41973 7527 41976
rect 7469 41967 7527 41973
rect 7558 41964 7564 41976
rect 7616 41964 7622 42016
rect 8110 41964 8116 42016
rect 8168 41964 8174 42016
rect 8478 41964 8484 42016
rect 8536 42004 8542 42016
rect 9048 42004 9076 42035
rect 10410 42032 10416 42084
rect 10468 42032 10474 42084
rect 10778 42032 10784 42084
rect 10836 42072 10842 42084
rect 11514 42072 11520 42084
rect 10836 42044 11520 42072
rect 10836 42032 10842 42044
rect 11514 42032 11520 42044
rect 11572 42032 11578 42084
rect 12008 42075 12066 42081
rect 12008 42041 12020 42075
rect 12054 42072 12066 42075
rect 12054 42044 12664 42072
rect 12054 42041 12066 42044
rect 12008 42035 12066 42041
rect 8536 41976 9076 42004
rect 8536 41964 8542 41976
rect 9858 41964 9864 42016
rect 9916 41964 9922 42016
rect 10042 41964 10048 42016
rect 10100 41964 10106 42016
rect 10502 41964 10508 42016
rect 10560 41964 10566 42016
rect 552 41914 12604 41936
rect 552 41862 4322 41914
rect 4374 41862 4386 41914
rect 4438 41862 4450 41914
rect 4502 41862 4514 41914
rect 4566 41862 4578 41914
rect 4630 41862 10722 41914
rect 10774 41862 10786 41914
rect 10838 41862 10850 41914
rect 10902 41862 10914 41914
rect 10966 41862 10978 41914
rect 11030 41862 12604 41914
rect 552 41840 12604 41862
rect 1026 41760 1032 41812
rect 1084 41760 1090 41812
rect 1213 41803 1271 41809
rect 1213 41769 1225 41803
rect 1259 41800 1271 41803
rect 1854 41800 1860 41812
rect 1259 41772 1860 41800
rect 1259 41769 1271 41772
rect 1213 41763 1271 41769
rect 1854 41760 1860 41772
rect 1912 41760 1918 41812
rect 2590 41800 2596 41812
rect 1964 41772 2596 41800
rect 1044 41732 1072 41760
rect 1964 41732 1992 41772
rect 2590 41760 2596 41772
rect 2648 41760 2654 41812
rect 4798 41760 4804 41812
rect 4856 41800 4862 41812
rect 6089 41803 6147 41809
rect 6089 41800 6101 41803
rect 4856 41772 6101 41800
rect 4856 41760 4862 41772
rect 6089 41769 6101 41772
rect 6135 41769 6147 41803
rect 6089 41763 6147 41769
rect 7024 41772 8616 41800
rect 1044 41704 1992 41732
rect 2133 41735 2191 41741
rect 2133 41701 2145 41735
rect 2179 41732 2191 41735
rect 4494 41735 4552 41741
rect 4494 41732 4506 41735
rect 2179 41704 4506 41732
rect 2179 41701 2191 41704
rect 2133 41695 2191 41701
rect 4494 41701 4506 41704
rect 4540 41701 4552 41735
rect 4494 41695 4552 41701
rect 5626 41692 5632 41744
rect 5684 41732 5690 41744
rect 6730 41732 6736 41744
rect 5684 41704 6736 41732
rect 5684 41692 5690 41704
rect 6730 41692 6736 41704
rect 6788 41692 6794 41744
rect 937 41667 995 41673
rect 937 41633 949 41667
rect 983 41664 995 41667
rect 1026 41664 1032 41676
rect 983 41636 1032 41664
rect 983 41633 995 41636
rect 937 41627 995 41633
rect 1026 41624 1032 41636
rect 1084 41624 1090 41676
rect 1121 41667 1179 41673
rect 1121 41633 1133 41667
rect 1167 41633 1179 41667
rect 1121 41627 1179 41633
rect 1136 41460 1164 41627
rect 1302 41624 1308 41676
rect 1360 41664 1366 41676
rect 2225 41667 2283 41673
rect 2225 41664 2237 41667
rect 1360 41636 2237 41664
rect 1360 41624 1366 41636
rect 2225 41633 2237 41636
rect 2271 41664 2283 41667
rect 2314 41664 2320 41676
rect 2271 41636 2320 41664
rect 2271 41633 2283 41636
rect 2225 41627 2283 41633
rect 2314 41624 2320 41636
rect 2372 41624 2378 41676
rect 2498 41673 2504 41676
rect 2492 41627 2504 41673
rect 2498 41624 2504 41627
rect 2556 41624 2562 41676
rect 2866 41624 2872 41676
rect 2924 41664 2930 41676
rect 3881 41667 3939 41673
rect 3881 41664 3893 41667
rect 2924 41636 3893 41664
rect 2924 41624 2930 41636
rect 3881 41633 3893 41636
rect 3927 41633 3939 41667
rect 3881 41627 3939 41633
rect 4154 41624 4160 41676
rect 4212 41624 4218 41676
rect 5813 41667 5871 41673
rect 5813 41633 5825 41667
rect 5859 41664 5871 41667
rect 5902 41664 5908 41676
rect 5859 41636 5908 41664
rect 5859 41633 5871 41636
rect 5813 41627 5871 41633
rect 5902 41624 5908 41636
rect 5960 41624 5966 41676
rect 5994 41624 6000 41676
rect 6052 41624 6058 41676
rect 7024 41664 7052 41772
rect 7374 41692 7380 41744
rect 7432 41692 7438 41744
rect 8478 41732 8484 41744
rect 8036 41704 8484 41732
rect 8036 41673 8064 41704
rect 8478 41692 8484 41704
rect 8536 41692 8542 41744
rect 8588 41732 8616 41772
rect 9214 41760 9220 41812
rect 9272 41760 9278 41812
rect 10778 41760 10784 41812
rect 10836 41760 10842 41812
rect 11790 41760 11796 41812
rect 11848 41800 11854 41812
rect 12069 41803 12127 41809
rect 12069 41800 12081 41803
rect 11848 41772 12081 41800
rect 11848 41760 11854 41772
rect 12069 41769 12081 41772
rect 12115 41769 12127 41803
rect 12069 41763 12127 41769
rect 12253 41803 12311 41809
rect 12253 41769 12265 41803
rect 12299 41800 12311 41803
rect 12636 41800 12664 42044
rect 12299 41772 12664 41800
rect 12299 41769 12311 41772
rect 12253 41763 12311 41769
rect 9033 41735 9091 41741
rect 9033 41732 9045 41735
rect 8588 41704 9045 41732
rect 9033 41701 9045 41704
rect 9079 41732 9091 41735
rect 10536 41735 10594 41741
rect 9079 41704 9674 41732
rect 9079 41701 9091 41704
rect 9033 41695 9091 41701
rect 6104 41636 7052 41664
rect 8021 41667 8079 41673
rect 1581 41599 1639 41605
rect 1581 41565 1593 41599
rect 1627 41565 1639 41599
rect 1581 41559 1639 41565
rect 1397 41531 1455 41537
rect 1397 41497 1409 41531
rect 1443 41528 1455 41531
rect 1486 41528 1492 41540
rect 1443 41500 1492 41528
rect 1443 41497 1455 41500
rect 1397 41491 1455 41497
rect 1486 41488 1492 41500
rect 1544 41488 1550 41540
rect 1596 41528 1624 41559
rect 3326 41556 3332 41608
rect 3384 41596 3390 41608
rect 3786 41596 3792 41608
rect 3384 41568 3792 41596
rect 3384 41556 3390 41568
rect 3786 41556 3792 41568
rect 3844 41596 3850 41608
rect 4065 41599 4123 41605
rect 4065 41596 4077 41599
rect 3844 41568 4077 41596
rect 3844 41556 3850 41568
rect 4065 41565 4077 41568
rect 4111 41565 4123 41599
rect 4065 41559 4123 41565
rect 4246 41556 4252 41608
rect 4304 41556 4310 41608
rect 5718 41556 5724 41608
rect 5776 41596 5782 41608
rect 6104 41596 6132 41636
rect 8021 41633 8033 41667
rect 8067 41633 8079 41667
rect 8021 41627 8079 41633
rect 8110 41624 8116 41676
rect 8168 41664 8174 41676
rect 8297 41667 8355 41673
rect 8297 41664 8309 41667
rect 8168 41636 8309 41664
rect 8168 41624 8174 41636
rect 8297 41633 8309 41636
rect 8343 41633 8355 41667
rect 8297 41627 8355 41633
rect 8662 41624 8668 41676
rect 8720 41664 8726 41676
rect 8849 41667 8907 41673
rect 8849 41664 8861 41667
rect 8720 41636 8861 41664
rect 8720 41624 8726 41636
rect 8849 41633 8861 41636
rect 8895 41633 8907 41667
rect 9646 41664 9674 41704
rect 10536 41701 10548 41735
rect 10582 41732 10594 41735
rect 10796 41732 10824 41760
rect 10582 41704 10824 41732
rect 10582 41701 10594 41704
rect 10536 41695 10594 41701
rect 10870 41692 10876 41744
rect 10928 41732 10934 41744
rect 11054 41732 11060 41744
rect 10928 41704 11060 41732
rect 10928 41692 10934 41704
rect 11054 41692 11060 41704
rect 11112 41732 11118 41744
rect 11112 41704 11376 41732
rect 11112 41692 11118 41704
rect 11348 41673 11376 41704
rect 11241 41667 11299 41673
rect 10704 41664 10824 41667
rect 11241 41664 11253 41667
rect 9646 41639 11253 41664
rect 9646 41636 10732 41639
rect 10796 41636 11253 41639
rect 8849 41627 8907 41633
rect 5776 41568 6132 41596
rect 5776 41556 5782 41568
rect 6178 41556 6184 41608
rect 6236 41596 6242 41608
rect 6641 41599 6699 41605
rect 6641 41596 6653 41599
rect 6236 41568 6653 41596
rect 6236 41556 6242 41568
rect 6641 41565 6653 41568
rect 6687 41596 6699 41599
rect 7190 41596 7196 41608
rect 6687 41568 7196 41596
rect 6687 41565 6699 41568
rect 6641 41559 6699 41565
rect 7190 41556 7196 41568
rect 7248 41556 7254 41608
rect 10781 41599 10839 41605
rect 10781 41565 10793 41599
rect 10827 41565 10839 41599
rect 10781 41559 10839 41565
rect 3697 41531 3755 41537
rect 3697 41528 3709 41531
rect 1596 41500 2268 41528
rect 1854 41460 1860 41472
rect 1136 41432 1860 41460
rect 1854 41420 1860 41432
rect 1912 41420 1918 41472
rect 2240 41460 2268 41500
rect 3252 41500 3709 41528
rect 3252 41460 3280 41500
rect 3697 41497 3709 41500
rect 3743 41497 3755 41531
rect 3697 41491 3755 41497
rect 3970 41488 3976 41540
rect 4028 41528 4034 41540
rect 4028 41500 4292 41528
rect 4028 41488 4034 41500
rect 2240 41432 3280 41460
rect 3510 41420 3516 41472
rect 3568 41460 3574 41472
rect 3605 41463 3663 41469
rect 3605 41460 3617 41463
rect 3568 41432 3617 41460
rect 3568 41420 3574 41432
rect 3605 41429 3617 41432
rect 3651 41429 3663 41463
rect 4264 41460 4292 41500
rect 6362 41488 6368 41540
rect 6420 41528 6426 41540
rect 9030 41528 9036 41540
rect 6420 41500 9036 41528
rect 6420 41488 6426 41500
rect 9030 41488 9036 41500
rect 9088 41528 9094 41540
rect 9088 41500 9904 41528
rect 9088 41488 9094 41500
rect 5626 41460 5632 41472
rect 4264 41432 5632 41460
rect 3605 41423 3663 41429
rect 5626 41420 5632 41432
rect 5684 41420 5690 41472
rect 5905 41463 5963 41469
rect 5905 41429 5917 41463
rect 5951 41460 5963 41463
rect 7098 41460 7104 41472
rect 5951 41432 7104 41460
rect 5951 41429 5963 41432
rect 5905 41423 5963 41429
rect 7098 41420 7104 41432
rect 7156 41420 7162 41472
rect 7190 41420 7196 41472
rect 7248 41460 7254 41472
rect 8662 41460 8668 41472
rect 7248 41432 8668 41460
rect 7248 41420 7254 41432
rect 8662 41420 8668 41432
rect 8720 41420 8726 41472
rect 9398 41420 9404 41472
rect 9456 41420 9462 41472
rect 9876 41460 9904 41500
rect 10042 41460 10048 41472
rect 9876 41432 10048 41460
rect 10042 41420 10048 41432
rect 10100 41420 10106 41472
rect 10594 41420 10600 41472
rect 10652 41460 10658 41472
rect 10787 41460 10815 41559
rect 10980 41528 11008 41636
rect 11241 41633 11253 41636
rect 11287 41633 11299 41667
rect 11241 41627 11299 41633
rect 11333 41667 11391 41673
rect 11333 41633 11345 41667
rect 11379 41633 11391 41667
rect 11333 41627 11391 41633
rect 11425 41667 11483 41673
rect 11425 41633 11437 41667
rect 11471 41633 11483 41667
rect 11425 41627 11483 41633
rect 11609 41667 11667 41673
rect 11609 41633 11621 41667
rect 11655 41664 11667 41667
rect 11655 41636 12112 41664
rect 11655 41633 11667 41636
rect 11609 41627 11667 41633
rect 11054 41556 11060 41608
rect 11112 41596 11118 41608
rect 11440 41596 11468 41627
rect 11112 41568 11468 41596
rect 11112 41556 11118 41568
rect 11514 41556 11520 41608
rect 11572 41596 11578 41608
rect 11701 41599 11759 41605
rect 11701 41596 11713 41599
rect 11572 41568 11713 41596
rect 11572 41556 11578 41568
rect 11701 41565 11713 41568
rect 11747 41565 11759 41599
rect 11701 41559 11759 41565
rect 10980 41500 11560 41528
rect 11532 41472 11560 41500
rect 10652 41432 10815 41460
rect 10652 41420 10658 41432
rect 10962 41420 10968 41472
rect 11020 41420 11026 41472
rect 11514 41420 11520 41472
rect 11572 41420 11578 41472
rect 12084 41469 12112 41636
rect 12069 41463 12127 41469
rect 12069 41429 12081 41463
rect 12115 41460 12127 41463
rect 12526 41460 12532 41472
rect 12115 41432 12532 41460
rect 12115 41429 12127 41432
rect 12069 41423 12127 41429
rect 12526 41420 12532 41432
rect 12584 41420 12590 41472
rect 552 41370 12604 41392
rect 552 41318 3662 41370
rect 3714 41318 3726 41370
rect 3778 41318 3790 41370
rect 3842 41318 3854 41370
rect 3906 41318 3918 41370
rect 3970 41318 10062 41370
rect 10114 41318 10126 41370
rect 10178 41318 10190 41370
rect 10242 41318 10254 41370
rect 10306 41318 10318 41370
rect 10370 41318 12604 41370
rect 552 41296 12604 41318
rect 1210 41216 1216 41268
rect 1268 41256 1274 41268
rect 2682 41256 2688 41268
rect 1268 41228 2688 41256
rect 1268 41216 1274 41228
rect 2682 41216 2688 41228
rect 2740 41216 2746 41268
rect 5074 41216 5080 41268
rect 5132 41256 5138 41268
rect 6914 41256 6920 41268
rect 5132 41228 6920 41256
rect 5132 41216 5138 41228
rect 6914 41216 6920 41228
rect 6972 41216 6978 41268
rect 7024 41228 8156 41256
rect 6638 41148 6644 41200
rect 6696 41148 6702 41200
rect 6730 41148 6736 41200
rect 6788 41188 6794 41200
rect 7024 41188 7052 41228
rect 6788 41160 7052 41188
rect 7561 41191 7619 41197
rect 6788 41148 6794 41160
rect 7561 41157 7573 41191
rect 7607 41188 7619 41191
rect 7742 41188 7748 41200
rect 7607 41160 7748 41188
rect 7607 41157 7619 41160
rect 7561 41151 7619 41157
rect 7742 41148 7748 41160
rect 7800 41148 7806 41200
rect 8018 41148 8024 41200
rect 8076 41148 8082 41200
rect 845 41123 903 41129
rect 845 41089 857 41123
rect 891 41120 903 41123
rect 1118 41120 1124 41132
rect 891 41092 1124 41120
rect 891 41089 903 41092
rect 845 41083 903 41089
rect 1118 41080 1124 41092
rect 1176 41080 1182 41132
rect 1302 41080 1308 41132
rect 1360 41120 1366 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 1360 41092 1409 41120
rect 1360 41080 1366 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 6656 41120 6684 41148
rect 8128 41132 8156 41228
rect 11514 41216 11520 41268
rect 11572 41256 11578 41268
rect 11793 41259 11851 41265
rect 11793 41256 11805 41259
rect 11572 41228 11805 41256
rect 11572 41216 11578 41228
rect 11793 41225 11805 41228
rect 11839 41225 11851 41259
rect 11793 41219 11851 41225
rect 8389 41191 8447 41197
rect 8389 41157 8401 41191
rect 8435 41188 8447 41191
rect 8435 41160 9444 41188
rect 8435 41157 8447 41160
rect 8389 41151 8447 41157
rect 7653 41123 7711 41129
rect 6656 41092 7604 41120
rect 1397 41083 1455 41089
rect 1029 41055 1087 41061
rect 1029 41021 1041 41055
rect 1075 41021 1087 41055
rect 1029 41015 1087 41021
rect 1213 41055 1271 41061
rect 1213 41021 1225 41055
rect 1259 41052 1271 41055
rect 1486 41052 1492 41064
rect 1259 41024 1492 41052
rect 1259 41021 1271 41024
rect 1213 41015 1271 41021
rect 1044 40984 1072 41015
rect 1486 41012 1492 41024
rect 1544 41012 1550 41064
rect 1673 41055 1731 41061
rect 1673 41021 1685 41055
rect 1719 41052 1731 41055
rect 1762 41052 1768 41064
rect 1719 41024 1768 41052
rect 1719 41021 1731 41024
rect 1673 41015 1731 41021
rect 1762 41012 1768 41024
rect 1820 41012 1826 41064
rect 2314 41012 2320 41064
rect 2372 41052 2378 41064
rect 3697 41055 3755 41061
rect 3697 41052 3709 41055
rect 2372 41024 3709 41052
rect 2372 41012 2378 41024
rect 3697 41021 3709 41024
rect 3743 41052 3755 41055
rect 4246 41052 4252 41064
rect 3743 41024 4252 41052
rect 3743 41021 3755 41024
rect 3697 41015 3755 41021
rect 4246 41012 4252 41024
rect 4304 41052 4310 41064
rect 5074 41052 5080 41064
rect 4304 41024 5080 41052
rect 4304 41012 4310 41024
rect 5074 41012 5080 41024
rect 5132 41052 5138 41064
rect 5353 41055 5411 41061
rect 5353 41052 5365 41055
rect 5132 41024 5365 41052
rect 5132 41012 5138 41024
rect 5353 41021 5365 41024
rect 5399 41021 5411 41055
rect 5353 41015 5411 41021
rect 5902 41012 5908 41064
rect 5960 41052 5966 41064
rect 6638 41052 6644 41064
rect 5960 41024 6644 41052
rect 5960 41012 5966 41024
rect 6638 41012 6644 41024
rect 6696 41052 6702 41064
rect 6825 41055 6883 41061
rect 6825 41052 6837 41055
rect 6696 41024 6837 41052
rect 6696 41012 6702 41024
rect 6825 41021 6837 41024
rect 6871 41021 6883 41055
rect 7190 41052 7196 41064
rect 6825 41015 6883 41021
rect 7024 41024 7196 41052
rect 1394 40984 1400 40996
rect 1044 40956 1400 40984
rect 1394 40944 1400 40956
rect 1452 40944 1458 40996
rect 3050 40944 3056 40996
rect 3108 40944 3114 40996
rect 3513 40987 3571 40993
rect 3513 40953 3525 40987
rect 3559 40953 3571 40987
rect 3513 40947 3571 40953
rect 3964 40987 4022 40993
rect 3964 40953 3976 40987
rect 4010 40984 4022 40987
rect 4062 40984 4068 40996
rect 4010 40956 4068 40984
rect 4010 40953 4022 40956
rect 3964 40947 4022 40953
rect 2130 40876 2136 40928
rect 2188 40916 2194 40928
rect 2590 40916 2596 40928
rect 2188 40888 2596 40916
rect 2188 40876 2194 40888
rect 2590 40876 2596 40888
rect 2648 40876 2654 40928
rect 3418 40876 3424 40928
rect 3476 40876 3482 40928
rect 3528 40916 3556 40947
rect 4062 40944 4068 40956
rect 4120 40944 4126 40996
rect 5620 40987 5678 40993
rect 5000 40956 5580 40984
rect 5000 40916 5028 40956
rect 5552 40928 5580 40956
rect 5620 40953 5632 40987
rect 5666 40984 5678 40987
rect 5810 40984 5816 40996
rect 5666 40956 5816 40984
rect 5666 40953 5678 40956
rect 5620 40947 5678 40953
rect 5810 40944 5816 40956
rect 5868 40944 5874 40996
rect 6086 40944 6092 40996
rect 6144 40984 6150 40996
rect 7024 40993 7052 41024
rect 7190 41012 7196 41024
rect 7248 41012 7254 41064
rect 7285 41055 7343 41061
rect 7285 41021 7297 41055
rect 7331 41052 7343 41055
rect 7374 41052 7380 41064
rect 7331 41024 7380 41052
rect 7331 41021 7343 41024
rect 7285 41015 7343 41021
rect 7374 41012 7380 41024
rect 7432 41012 7438 41064
rect 7466 41012 7472 41064
rect 7524 41012 7530 41064
rect 7576 41052 7604 41092
rect 7653 41089 7665 41123
rect 7699 41120 7711 41123
rect 7834 41120 7840 41132
rect 7699 41092 7840 41120
rect 7699 41089 7711 41092
rect 7653 41083 7711 41089
rect 7834 41080 7840 41092
rect 7892 41080 7898 41132
rect 8110 41080 8116 41132
rect 8168 41080 8174 41132
rect 7745 41055 7803 41061
rect 7745 41052 7757 41055
rect 7576 41024 7757 41052
rect 7745 41021 7757 41024
rect 7791 41052 7803 41055
rect 7926 41052 7932 41064
rect 7791 41024 7932 41052
rect 7791 41021 7803 41024
rect 7745 41015 7803 41021
rect 7926 41012 7932 41024
rect 7984 41012 7990 41064
rect 8021 41055 8079 41061
rect 8021 41021 8033 41055
rect 8067 41021 8079 41055
rect 8128 41052 8156 41080
rect 8205 41055 8263 41061
rect 8205 41052 8217 41055
rect 8128 41024 8217 41052
rect 8021 41015 8079 41021
rect 8205 41021 8217 41024
rect 8251 41021 8263 41055
rect 8205 41015 8263 41021
rect 8665 41055 8723 41061
rect 8665 41021 8677 41055
rect 8711 41052 8723 41055
rect 8938 41052 8944 41064
rect 8711 41024 8944 41052
rect 8711 41021 8723 41024
rect 8665 41015 8723 41021
rect 7009 40987 7067 40993
rect 7009 40984 7021 40987
rect 6144 40956 7021 40984
rect 6144 40944 6150 40956
rect 7009 40953 7021 40956
rect 7055 40953 7067 40987
rect 7484 40984 7512 41012
rect 7009 40947 7067 40953
rect 7116 40956 7512 40984
rect 3528 40888 5028 40916
rect 5077 40919 5135 40925
rect 5077 40885 5089 40919
rect 5123 40916 5135 40919
rect 5166 40916 5172 40928
rect 5123 40888 5172 40916
rect 5123 40885 5135 40888
rect 5077 40879 5135 40885
rect 5166 40876 5172 40888
rect 5224 40876 5230 40928
rect 5534 40876 5540 40928
rect 5592 40876 5598 40928
rect 5994 40876 6000 40928
rect 6052 40916 6058 40928
rect 6178 40916 6184 40928
rect 6052 40888 6184 40916
rect 6052 40876 6058 40888
rect 6178 40876 6184 40888
rect 6236 40916 6242 40928
rect 6733 40919 6791 40925
rect 6733 40916 6745 40919
rect 6236 40888 6745 40916
rect 6236 40876 6242 40888
rect 6733 40885 6745 40888
rect 6779 40885 6791 40919
rect 6733 40879 6791 40885
rect 6822 40876 6828 40928
rect 6880 40916 6886 40928
rect 7116 40916 7144 40956
rect 6880 40888 7144 40916
rect 7193 40919 7251 40925
rect 6880 40876 6886 40888
rect 7193 40885 7205 40919
rect 7239 40916 7251 40919
rect 7374 40916 7380 40928
rect 7239 40888 7380 40916
rect 7239 40885 7251 40888
rect 7193 40879 7251 40885
rect 7374 40876 7380 40888
rect 7432 40876 7438 40928
rect 7929 40919 7987 40925
rect 7929 40885 7941 40919
rect 7975 40916 7987 40919
rect 8036 40916 8064 41015
rect 8938 41012 8944 41024
rect 8996 41052 9002 41064
rect 8996 41024 9260 41052
rect 8996 41012 9002 41024
rect 8386 40944 8392 40996
rect 8444 40944 8450 40996
rect 8573 40987 8631 40993
rect 8573 40953 8585 40987
rect 8619 40984 8631 40987
rect 8846 40984 8852 40996
rect 8619 40956 8852 40984
rect 8619 40953 8631 40956
rect 8573 40947 8631 40953
rect 8846 40944 8852 40956
rect 8904 40984 8910 40996
rect 8904 40956 9168 40984
rect 8904 40944 8910 40956
rect 9140 40928 9168 40956
rect 8294 40916 8300 40928
rect 7975 40888 8300 40916
rect 7975 40885 7987 40888
rect 7929 40879 7987 40885
rect 8294 40876 8300 40888
rect 8352 40876 8358 40928
rect 8478 40876 8484 40928
rect 8536 40916 8542 40928
rect 8757 40919 8815 40925
rect 8757 40916 8769 40919
rect 8536 40888 8769 40916
rect 8536 40876 8542 40888
rect 8757 40885 8769 40888
rect 8803 40885 8815 40919
rect 8757 40879 8815 40885
rect 9122 40876 9128 40928
rect 9180 40876 9186 40928
rect 9232 40916 9260 41024
rect 9306 41012 9312 41064
rect 9364 41012 9370 41064
rect 9416 41061 9444 41160
rect 11977 41123 12035 41129
rect 11977 41089 11989 41123
rect 12023 41120 12035 41123
rect 12618 41120 12624 41132
rect 12023 41092 12624 41120
rect 12023 41089 12035 41092
rect 11977 41083 12035 41089
rect 12618 41080 12624 41092
rect 12676 41080 12682 41132
rect 9401 41055 9459 41061
rect 9401 41021 9413 41055
rect 9447 41021 9459 41055
rect 9401 41015 9459 41021
rect 10413 41055 10471 41061
rect 10413 41021 10425 41055
rect 10459 41052 10471 41055
rect 10502 41052 10508 41064
rect 10459 41024 10508 41052
rect 10459 41021 10471 41024
rect 10413 41015 10471 41021
rect 10502 41012 10508 41024
rect 10560 41012 10566 41064
rect 10680 41055 10738 41061
rect 10680 41021 10692 41055
rect 10726 41052 10738 41055
rect 10962 41052 10968 41064
rect 10726 41024 10968 41052
rect 10726 41021 10738 41024
rect 10680 41015 10738 41021
rect 10962 41012 10968 41024
rect 11020 41012 11026 41064
rect 11146 41012 11152 41064
rect 11204 41012 11210 41064
rect 12158 41012 12164 41064
rect 12216 41012 12222 41064
rect 12253 41055 12311 41061
rect 12253 41021 12265 41055
rect 12299 41021 12311 41055
rect 12253 41015 12311 41021
rect 9950 40944 9956 40996
rect 10008 40944 10014 40996
rect 10042 40944 10048 40996
rect 10100 40984 10106 40996
rect 10137 40987 10195 40993
rect 10137 40984 10149 40987
rect 10100 40956 10149 40984
rect 10100 40944 10106 40956
rect 10137 40953 10149 40956
rect 10183 40984 10195 40987
rect 11164 40984 11192 41012
rect 10183 40956 11192 40984
rect 10183 40953 10195 40956
rect 10137 40947 10195 40953
rect 11790 40944 11796 40996
rect 11848 40984 11854 40996
rect 12268 40984 12296 41015
rect 11848 40956 12296 40984
rect 11848 40944 11854 40956
rect 10321 40919 10379 40925
rect 10321 40916 10333 40919
rect 9232 40888 10333 40916
rect 10321 40885 10333 40888
rect 10367 40885 10379 40919
rect 10321 40879 10379 40885
rect 11146 40876 11152 40928
rect 11204 40916 11210 40928
rect 11977 40919 12035 40925
rect 11977 40916 11989 40919
rect 11204 40888 11989 40916
rect 11204 40876 11210 40888
rect 11977 40885 11989 40888
rect 12023 40885 12035 40919
rect 11977 40879 12035 40885
rect 552 40826 12604 40848
rect 552 40774 4322 40826
rect 4374 40774 4386 40826
rect 4438 40774 4450 40826
rect 4502 40774 4514 40826
rect 4566 40774 4578 40826
rect 4630 40774 10722 40826
rect 10774 40774 10786 40826
rect 10838 40774 10850 40826
rect 10902 40774 10914 40826
rect 10966 40774 10978 40826
rect 11030 40774 12604 40826
rect 552 40752 12604 40774
rect 1210 40672 1216 40724
rect 1268 40672 1274 40724
rect 1394 40672 1400 40724
rect 1452 40712 1458 40724
rect 1673 40715 1731 40721
rect 1673 40712 1685 40715
rect 1452 40684 1685 40712
rect 1452 40672 1458 40684
rect 1673 40681 1685 40684
rect 1719 40712 1731 40715
rect 2498 40712 2504 40724
rect 1719 40684 2504 40712
rect 1719 40681 1731 40684
rect 1673 40675 1731 40681
rect 2498 40672 2504 40684
rect 2556 40672 2562 40724
rect 4154 40672 4160 40724
rect 4212 40712 4218 40724
rect 5445 40715 5503 40721
rect 4212 40684 5212 40712
rect 4212 40672 4218 40684
rect 3234 40604 3240 40656
rect 3292 40604 3298 40656
rect 3510 40604 3516 40656
rect 3568 40644 3574 40656
rect 3568 40616 4936 40644
rect 3568 40604 3574 40616
rect 1302 40536 1308 40588
rect 1360 40576 1366 40588
rect 1397 40579 1455 40585
rect 1397 40576 1409 40579
rect 1360 40548 1409 40576
rect 1360 40536 1366 40548
rect 1397 40545 1409 40548
rect 1443 40545 1455 40579
rect 1397 40539 1455 40545
rect 2314 40536 2320 40588
rect 2372 40536 2378 40588
rect 2406 40536 2412 40588
rect 2464 40576 2470 40588
rect 2573 40579 2631 40585
rect 2573 40576 2585 40579
rect 2464 40548 2585 40576
rect 2464 40536 2470 40548
rect 2573 40545 2585 40548
rect 2619 40545 2631 40579
rect 3252 40576 3280 40604
rect 4019 40579 4077 40585
rect 4019 40576 4031 40579
rect 3252 40548 4031 40576
rect 2573 40539 2631 40545
rect 4019 40545 4031 40548
rect 4065 40545 4077 40579
rect 4019 40539 4077 40545
rect 4154 40536 4160 40588
rect 4212 40536 4218 40588
rect 4246 40536 4252 40588
rect 4304 40536 4310 40588
rect 4377 40579 4435 40585
rect 4377 40576 4389 40579
rect 4356 40545 4389 40576
rect 4423 40545 4435 40579
rect 4356 40539 4435 40545
rect 2130 40468 2136 40520
rect 2188 40468 2194 40520
rect 3326 40468 3332 40520
rect 3384 40508 3390 40520
rect 4356 40508 4384 40539
rect 4522 40536 4528 40588
rect 4580 40576 4586 40588
rect 4908 40585 4936 40616
rect 4982 40604 4988 40656
rect 5040 40644 5046 40656
rect 5184 40653 5212 40684
rect 5445 40681 5457 40715
rect 5491 40712 5503 40715
rect 8662 40712 8668 40724
rect 5491 40684 8668 40712
rect 5491 40681 5503 40684
rect 5445 40675 5503 40681
rect 8662 40672 8668 40684
rect 8720 40672 8726 40724
rect 11514 40672 11520 40724
rect 11572 40672 11578 40724
rect 5077 40647 5135 40653
rect 5077 40644 5089 40647
rect 5040 40616 5089 40644
rect 5040 40604 5046 40616
rect 5077 40613 5089 40616
rect 5123 40613 5135 40647
rect 5077 40607 5135 40613
rect 5169 40647 5227 40653
rect 5169 40613 5181 40647
rect 5215 40644 5227 40647
rect 5534 40644 5540 40656
rect 5215 40616 5540 40644
rect 5215 40613 5227 40616
rect 5169 40607 5227 40613
rect 5534 40604 5540 40616
rect 5592 40604 5598 40656
rect 6822 40644 6828 40656
rect 6472 40616 6828 40644
rect 4801 40579 4859 40585
rect 4801 40576 4813 40579
rect 4580 40548 4813 40576
rect 4580 40536 4586 40548
rect 4801 40545 4813 40548
rect 4847 40545 4859 40579
rect 4801 40539 4859 40545
rect 4894 40579 4952 40585
rect 4894 40545 4906 40579
rect 4940 40545 4952 40579
rect 4894 40539 4952 40545
rect 4614 40508 4620 40520
rect 3384 40480 4384 40508
rect 4449 40480 4620 40508
rect 3384 40468 3390 40480
rect 1486 40400 1492 40452
rect 1544 40440 1550 40452
rect 1762 40440 1768 40452
rect 1544 40412 1768 40440
rect 1544 40400 1550 40412
rect 1762 40400 1768 40412
rect 1820 40400 1826 40452
rect 3881 40443 3939 40449
rect 3881 40440 3893 40443
rect 3344 40412 3893 40440
rect 2222 40332 2228 40384
rect 2280 40372 2286 40384
rect 3344 40372 3372 40412
rect 3881 40409 3893 40412
rect 3927 40409 3939 40443
rect 3881 40403 3939 40409
rect 4246 40400 4252 40452
rect 4304 40440 4310 40452
rect 4449 40440 4477 40480
rect 4614 40468 4620 40480
rect 4672 40508 4678 40520
rect 5000 40508 5028 40604
rect 5258 40536 5264 40588
rect 5316 40585 5322 40588
rect 5316 40576 5324 40585
rect 5316 40548 5361 40576
rect 5316 40539 5324 40548
rect 5316 40536 5322 40539
rect 5442 40536 5448 40588
rect 5500 40576 5506 40588
rect 6178 40576 6184 40588
rect 5500 40548 6184 40576
rect 5500 40536 5506 40548
rect 6178 40536 6184 40548
rect 6236 40536 6242 40588
rect 4672 40480 5028 40508
rect 4672 40468 4678 40480
rect 6472 40440 6500 40616
rect 6822 40604 6828 40616
rect 6880 40604 6886 40656
rect 7098 40604 7104 40656
rect 7156 40644 7162 40656
rect 7156 40616 7604 40644
rect 7156 40604 7162 40616
rect 6638 40536 6644 40588
rect 6696 40536 6702 40588
rect 7374 40536 7380 40588
rect 7432 40536 7438 40588
rect 7576 40585 7604 40616
rect 7650 40604 7656 40656
rect 7708 40644 7714 40656
rect 8018 40644 8024 40656
rect 7708 40616 8024 40644
rect 7708 40604 7714 40616
rect 8018 40604 8024 40616
rect 8076 40604 8082 40656
rect 8202 40604 8208 40656
rect 8260 40604 8266 40656
rect 9858 40644 9864 40656
rect 8680 40616 9864 40644
rect 7561 40579 7619 40585
rect 7561 40545 7573 40579
rect 7607 40576 7619 40579
rect 8220 40576 8248 40604
rect 8680 40585 8708 40616
rect 9858 40604 9864 40616
rect 9916 40604 9922 40656
rect 11532 40644 11560 40672
rect 12526 40644 12532 40656
rect 11256 40616 12532 40644
rect 8297 40579 8355 40585
rect 8297 40576 8309 40579
rect 7607 40548 7880 40576
rect 8220 40548 8309 40576
rect 7607 40545 7619 40548
rect 7561 40539 7619 40545
rect 6549 40511 6607 40517
rect 6549 40477 6561 40511
rect 6595 40477 6607 40511
rect 6549 40471 6607 40477
rect 4304 40412 4477 40440
rect 5000 40412 6500 40440
rect 6564 40440 6592 40471
rect 7466 40468 7472 40520
rect 7524 40508 7530 40520
rect 7745 40511 7803 40517
rect 7745 40508 7757 40511
rect 7524 40480 7757 40508
rect 7524 40468 7530 40480
rect 7745 40477 7757 40480
rect 7791 40477 7803 40511
rect 7852 40508 7880 40548
rect 8297 40545 8309 40548
rect 8343 40545 8355 40579
rect 8297 40539 8355 40545
rect 8665 40579 8723 40585
rect 8665 40545 8677 40579
rect 8711 40545 8723 40579
rect 8665 40539 8723 40545
rect 9122 40536 9128 40588
rect 9180 40536 9186 40588
rect 9214 40536 9220 40588
rect 9272 40576 9278 40588
rect 9582 40576 9588 40588
rect 9272 40548 9588 40576
rect 9272 40536 9278 40548
rect 9582 40536 9588 40548
rect 9640 40536 9646 40588
rect 9766 40536 9772 40588
rect 9824 40576 9830 40588
rect 11256 40585 11284 40616
rect 12526 40604 12532 40616
rect 12584 40604 12590 40656
rect 10965 40579 11023 40585
rect 10965 40576 10977 40579
rect 9824 40548 10977 40576
rect 9824 40536 9830 40548
rect 10965 40545 10977 40548
rect 11011 40545 11023 40579
rect 10965 40539 11023 40545
rect 11241 40579 11299 40585
rect 11241 40545 11253 40579
rect 11287 40545 11299 40579
rect 11241 40539 11299 40545
rect 11422 40536 11428 40588
rect 11480 40536 11486 40588
rect 11517 40579 11575 40585
rect 11517 40545 11529 40579
rect 11563 40545 11575 40579
rect 11517 40539 11575 40545
rect 11609 40579 11667 40585
rect 11609 40545 11621 40579
rect 11655 40576 11667 40579
rect 12069 40579 12127 40585
rect 11655 40548 11836 40576
rect 11655 40545 11667 40548
rect 11609 40539 11667 40545
rect 8754 40508 8760 40520
rect 7852 40480 8760 40508
rect 7745 40471 7803 40477
rect 8754 40468 8760 40480
rect 8812 40468 8818 40520
rect 11330 40468 11336 40520
rect 11388 40508 11394 40520
rect 11532 40508 11560 40539
rect 11698 40508 11704 40520
rect 11388 40480 11704 40508
rect 11388 40468 11394 40480
rect 11698 40468 11704 40480
rect 11756 40468 11762 40520
rect 7650 40440 7656 40452
rect 6564 40412 7656 40440
rect 4304 40400 4310 40412
rect 5000 40384 5028 40412
rect 7650 40400 7656 40412
rect 7708 40400 7714 40452
rect 8386 40400 8392 40452
rect 8444 40440 8450 40452
rect 10137 40443 10195 40449
rect 10137 40440 10149 40443
rect 8444 40412 10149 40440
rect 8444 40400 8450 40412
rect 10137 40409 10149 40412
rect 10183 40409 10195 40443
rect 10137 40403 10195 40409
rect 10686 40400 10692 40452
rect 10744 40440 10750 40452
rect 11238 40440 11244 40452
rect 10744 40412 11244 40440
rect 10744 40400 10750 40412
rect 11238 40400 11244 40412
rect 11296 40440 11302 40452
rect 11808 40440 11836 40548
rect 12069 40545 12081 40579
rect 12115 40576 12127 40579
rect 12342 40576 12348 40588
rect 12115 40548 12348 40576
rect 12115 40545 12127 40548
rect 12069 40539 12127 40545
rect 12342 40536 12348 40548
rect 12400 40536 12406 40588
rect 11296 40412 11836 40440
rect 11296 40400 11302 40412
rect 2280 40344 3372 40372
rect 3697 40375 3755 40381
rect 2280 40332 2286 40344
rect 3697 40341 3709 40375
rect 3743 40372 3755 40375
rect 4430 40372 4436 40384
rect 3743 40344 4436 40372
rect 3743 40341 3755 40344
rect 3697 40335 3755 40341
rect 4430 40332 4436 40344
rect 4488 40332 4494 40384
rect 4982 40332 4988 40384
rect 5040 40332 5046 40384
rect 5902 40332 5908 40384
rect 5960 40332 5966 40384
rect 7282 40332 7288 40384
rect 7340 40332 7346 40384
rect 7466 40332 7472 40384
rect 7524 40372 7530 40384
rect 7926 40372 7932 40384
rect 7524 40344 7932 40372
rect 7524 40332 7530 40344
rect 7926 40332 7932 40344
rect 7984 40332 7990 40384
rect 9214 40332 9220 40384
rect 9272 40372 9278 40384
rect 11057 40375 11115 40381
rect 11057 40372 11069 40375
rect 9272 40344 11069 40372
rect 9272 40332 9278 40344
rect 11057 40341 11069 40344
rect 11103 40341 11115 40375
rect 11057 40335 11115 40341
rect 11882 40332 11888 40384
rect 11940 40332 11946 40384
rect 12066 40332 12072 40384
rect 12124 40372 12130 40384
rect 12161 40375 12219 40381
rect 12161 40372 12173 40375
rect 12124 40344 12173 40372
rect 12124 40332 12130 40344
rect 12161 40341 12173 40344
rect 12207 40341 12219 40375
rect 12161 40335 12219 40341
rect 552 40282 12604 40304
rect 552 40230 3662 40282
rect 3714 40230 3726 40282
rect 3778 40230 3790 40282
rect 3842 40230 3854 40282
rect 3906 40230 3918 40282
rect 3970 40230 10062 40282
rect 10114 40230 10126 40282
rect 10178 40230 10190 40282
rect 10242 40230 10254 40282
rect 10306 40230 10318 40282
rect 10370 40230 12604 40282
rect 552 40208 12604 40230
rect 1762 40128 1768 40180
rect 1820 40168 1826 40180
rect 2130 40168 2136 40180
rect 1820 40140 2136 40168
rect 1820 40128 1826 40140
rect 2130 40128 2136 40140
rect 2188 40128 2194 40180
rect 2317 40171 2375 40177
rect 2317 40137 2329 40171
rect 2363 40168 2375 40171
rect 2406 40168 2412 40180
rect 2363 40140 2412 40168
rect 2363 40137 2375 40140
rect 2317 40131 2375 40137
rect 2406 40128 2412 40140
rect 2464 40128 2470 40180
rect 2498 40128 2504 40180
rect 2556 40128 2562 40180
rect 3050 40128 3056 40180
rect 3108 40168 3114 40180
rect 3694 40168 3700 40180
rect 3108 40140 3700 40168
rect 3108 40128 3114 40140
rect 3694 40128 3700 40140
rect 3752 40128 3758 40180
rect 6457 40171 6515 40177
rect 6457 40137 6469 40171
rect 6503 40168 6515 40171
rect 6638 40168 6644 40180
rect 6503 40140 6644 40168
rect 6503 40137 6515 40140
rect 6457 40131 6515 40137
rect 6638 40128 6644 40140
rect 6696 40128 6702 40180
rect 7650 40128 7656 40180
rect 7708 40168 7714 40180
rect 7745 40171 7803 40177
rect 7745 40168 7757 40171
rect 7708 40140 7757 40168
rect 7708 40128 7714 40140
rect 7745 40137 7757 40140
rect 7791 40137 7803 40171
rect 7745 40131 7803 40137
rect 8113 40171 8171 40177
rect 8113 40137 8125 40171
rect 8159 40168 8171 40171
rect 8202 40168 8208 40180
rect 8159 40140 8208 40168
rect 8159 40137 8171 40140
rect 8113 40131 8171 40137
rect 8202 40128 8208 40140
rect 8260 40168 8266 40180
rect 8481 40171 8539 40177
rect 8481 40168 8493 40171
rect 8260 40140 8493 40168
rect 8260 40128 8266 40140
rect 8481 40137 8493 40140
rect 8527 40137 8539 40171
rect 8481 40131 8539 40137
rect 9122 40128 9128 40180
rect 9180 40128 9186 40180
rect 9677 40171 9735 40177
rect 9677 40137 9689 40171
rect 9723 40168 9735 40171
rect 10502 40168 10508 40180
rect 9723 40140 10508 40168
rect 9723 40137 9735 40140
rect 9677 40131 9735 40137
rect 10502 40128 10508 40140
rect 10560 40128 10566 40180
rect 10597 40171 10655 40177
rect 10597 40137 10609 40171
rect 10643 40168 10655 40171
rect 10686 40168 10692 40180
rect 10643 40140 10692 40168
rect 10643 40137 10655 40140
rect 10597 40131 10655 40137
rect 10686 40128 10692 40140
rect 10744 40128 10750 40180
rect 1397 40103 1455 40109
rect 1397 40069 1409 40103
rect 1443 40100 1455 40103
rect 2038 40100 2044 40112
rect 1443 40072 2044 40100
rect 1443 40069 1455 40072
rect 1397 40063 1455 40069
rect 2038 40060 2044 40072
rect 2096 40060 2102 40112
rect 4154 40100 4160 40112
rect 3804 40072 4160 40100
rect 1946 40032 1952 40044
rect 1412 40004 1952 40032
rect 1026 39924 1032 39976
rect 1084 39964 1090 39976
rect 1121 39967 1179 39973
rect 1121 39964 1133 39967
rect 1084 39936 1133 39964
rect 1084 39924 1090 39936
rect 1121 39933 1133 39936
rect 1167 39933 1179 39967
rect 1121 39927 1179 39933
rect 1210 39924 1216 39976
rect 1268 39924 1274 39976
rect 1412 39973 1440 40004
rect 1946 39992 1952 40004
rect 2004 39992 2010 40044
rect 2406 40032 2412 40044
rect 2148 40004 2412 40032
rect 1397 39967 1455 39973
rect 1397 39933 1409 39967
rect 1443 39933 1455 39967
rect 1397 39927 1455 39933
rect 1489 39967 1547 39973
rect 1489 39933 1501 39967
rect 1535 39933 1547 39967
rect 1673 39967 1731 39973
rect 1673 39966 1685 39967
rect 1489 39927 1547 39933
rect 1596 39938 1685 39966
rect 1504 39896 1532 39927
rect 1136 39868 1532 39896
rect 1136 39840 1164 39868
rect 934 39788 940 39840
rect 992 39788 998 39840
rect 1118 39788 1124 39840
rect 1176 39788 1182 39840
rect 1486 39788 1492 39840
rect 1544 39828 1550 39840
rect 1596 39828 1624 39938
rect 1673 39933 1685 39938
rect 1719 39933 1731 39967
rect 1673 39927 1731 39933
rect 1857 39967 1915 39973
rect 1857 39933 1869 39967
rect 1903 39964 1915 39967
rect 2148 39964 2176 40004
rect 2406 39992 2412 40004
rect 2464 39992 2470 40044
rect 3804 40041 3832 40072
rect 4154 40060 4160 40072
rect 4212 40060 4218 40112
rect 4982 40100 4988 40112
rect 4356 40072 4988 40100
rect 3789 40035 3847 40041
rect 3789 40032 3801 40035
rect 2700 40004 3801 40032
rect 2700 39976 2728 40004
rect 3789 40001 3801 40004
rect 3835 40001 3847 40035
rect 4356 40032 4384 40072
rect 4982 40060 4988 40072
rect 5040 40060 5046 40112
rect 7374 40060 7380 40112
rect 7432 40100 7438 40112
rect 8849 40103 8907 40109
rect 8849 40100 8861 40103
rect 7432 40072 8861 40100
rect 7432 40060 7438 40072
rect 8849 40069 8861 40072
rect 8895 40069 8907 40103
rect 11054 40100 11060 40112
rect 8849 40063 8907 40069
rect 10428 40072 11060 40100
rect 10428 40044 10456 40072
rect 11054 40060 11060 40072
rect 11112 40060 11118 40112
rect 3789 39995 3847 40001
rect 4264 40004 4384 40032
rect 2682 39973 2688 39976
rect 1903 39936 2176 39964
rect 2651 39967 2688 39973
rect 1903 39933 1915 39936
rect 1857 39927 1915 39933
rect 2651 39933 2663 39967
rect 2651 39927 2688 39933
rect 2682 39924 2688 39927
rect 2740 39924 2746 39976
rect 2958 39924 2964 39976
rect 3016 39924 3022 39976
rect 3053 39967 3111 39973
rect 3053 39933 3065 39967
rect 3099 39964 3111 39967
rect 3528 39964 3740 39966
rect 4154 39964 4160 39976
rect 3099 39938 4160 39964
rect 3099 39936 3556 39938
rect 3712 39936 4160 39938
rect 3099 39933 3111 39936
rect 3053 39927 3111 39933
rect 4154 39924 4160 39936
rect 4212 39924 4218 39976
rect 4264 39973 4292 40004
rect 4522 39992 4528 40044
rect 4580 40032 4586 40044
rect 4580 40004 5028 40032
rect 4580 39992 4586 40004
rect 4249 39967 4307 39973
rect 4249 39933 4261 39967
rect 4295 39933 4307 39967
rect 4249 39927 4307 39933
rect 4338 39924 4344 39976
rect 4396 39924 4402 39976
rect 4430 39924 4436 39976
rect 4488 39964 4494 39976
rect 4488 39936 4533 39964
rect 4488 39924 4494 39936
rect 4614 39924 4620 39976
rect 4672 39924 4678 39976
rect 4890 39973 4896 39976
rect 4847 39967 4896 39973
rect 4847 39933 4859 39967
rect 4893 39933 4896 39967
rect 4847 39927 4896 39933
rect 4890 39924 4896 39927
rect 4948 39924 4954 39976
rect 5000 39964 5028 40004
rect 5074 39992 5080 40044
rect 5132 39992 5138 40044
rect 7282 39992 7288 40044
rect 7340 40032 7346 40044
rect 8205 40035 8263 40041
rect 8205 40032 8217 40035
rect 7340 40004 8217 40032
rect 7340 39992 7346 40004
rect 8205 40001 8217 40004
rect 8251 40001 8263 40035
rect 8205 39995 8263 40001
rect 10410 39992 10416 40044
rect 10468 39992 10474 40044
rect 11238 40032 11244 40044
rect 10529 40004 11244 40032
rect 5344 39967 5402 39973
rect 5000 39936 5309 39964
rect 1949 39899 2007 39905
rect 1949 39865 1961 39899
rect 1995 39896 2007 39899
rect 2038 39896 2044 39908
rect 1995 39868 2044 39896
rect 1995 39865 2007 39868
rect 1949 39859 2007 39865
rect 2038 39856 2044 39868
rect 2096 39856 2102 39908
rect 3142 39856 3148 39908
rect 3200 39896 3206 39908
rect 3200 39868 3372 39896
rect 3200 39856 3206 39868
rect 2159 39831 2217 39837
rect 2159 39828 2171 39831
rect 1544 39800 2171 39828
rect 1544 39788 1550 39800
rect 2159 39797 2171 39800
rect 2205 39828 2217 39831
rect 2958 39828 2964 39840
rect 2205 39800 2964 39828
rect 2205 39797 2217 39800
rect 2159 39791 2217 39797
rect 2958 39788 2964 39800
rect 3016 39828 3022 39840
rect 3237 39831 3295 39837
rect 3237 39828 3249 39831
rect 3016 39800 3249 39828
rect 3016 39788 3022 39800
rect 3237 39797 3249 39800
rect 3283 39797 3295 39831
rect 3344 39828 3372 39868
rect 3694 39856 3700 39908
rect 3752 39856 3758 39908
rect 3605 39831 3663 39837
rect 3605 39828 3617 39831
rect 3344 39800 3617 39828
rect 3237 39791 3295 39797
rect 3605 39797 3617 39800
rect 3651 39797 3663 39831
rect 3605 39791 3663 39797
rect 4157 39831 4215 39837
rect 4157 39797 4169 39831
rect 4203 39828 4215 39831
rect 4522 39828 4528 39840
rect 4203 39800 4528 39828
rect 4203 39797 4215 39800
rect 4157 39791 4215 39797
rect 4522 39788 4528 39800
rect 4580 39788 4586 39840
rect 4632 39828 4660 39924
rect 4709 39899 4767 39905
rect 4709 39865 4721 39899
rect 4755 39896 4767 39899
rect 5281 39896 5309 39936
rect 5344 39933 5356 39967
rect 5390 39964 5402 39967
rect 5902 39964 5908 39976
rect 5390 39936 5908 39964
rect 5390 39933 5402 39936
rect 5344 39927 5402 39933
rect 5902 39924 5908 39936
rect 5960 39924 5966 39976
rect 7006 39964 7012 39976
rect 6012 39936 7012 39964
rect 6012 39896 6040 39936
rect 7006 39924 7012 39936
rect 7064 39924 7070 39976
rect 7377 39967 7435 39973
rect 7377 39933 7389 39967
rect 7423 39964 7435 39967
rect 7466 39964 7472 39976
rect 7423 39936 7472 39964
rect 7423 39933 7435 39936
rect 7377 39927 7435 39933
rect 7466 39924 7472 39936
rect 7524 39924 7530 39976
rect 7558 39924 7564 39976
rect 7616 39924 7622 39976
rect 7929 39967 7987 39973
rect 7929 39933 7941 39967
rect 7975 39933 7987 39967
rect 7929 39927 7987 39933
rect 8389 39967 8447 39973
rect 8389 39933 8401 39967
rect 8435 39933 8447 39967
rect 8389 39927 8447 39933
rect 4755 39868 5120 39896
rect 5281 39868 6040 39896
rect 4755 39865 4767 39868
rect 4709 39859 4767 39865
rect 4798 39828 4804 39840
rect 4632 39800 4804 39828
rect 4798 39788 4804 39800
rect 4856 39788 4862 39840
rect 4982 39788 4988 39840
rect 5040 39788 5046 39840
rect 5092 39828 5120 39868
rect 6178 39856 6184 39908
rect 6236 39896 6242 39908
rect 7944 39896 7972 39927
rect 6236 39868 7972 39896
rect 6236 39856 6242 39868
rect 5350 39828 5356 39840
rect 5092 39800 5356 39828
rect 5350 39788 5356 39800
rect 5408 39788 5414 39840
rect 6362 39788 6368 39840
rect 6420 39828 6426 39840
rect 6549 39831 6607 39837
rect 6549 39828 6561 39831
rect 6420 39800 6561 39828
rect 6420 39788 6426 39800
rect 6549 39797 6561 39800
rect 6595 39797 6607 39831
rect 6549 39791 6607 39797
rect 7190 39788 7196 39840
rect 7248 39828 7254 39840
rect 7650 39828 7656 39840
rect 7248 39800 7656 39828
rect 7248 39788 7254 39800
rect 7650 39788 7656 39800
rect 7708 39788 7714 39840
rect 7742 39788 7748 39840
rect 7800 39828 7806 39840
rect 8404 39828 8432 39927
rect 8662 39924 8668 39976
rect 8720 39924 8726 39976
rect 8938 39924 8944 39976
rect 8996 39964 9002 39976
rect 9033 39967 9091 39973
rect 9033 39964 9045 39967
rect 8996 39936 9045 39964
rect 8996 39924 9002 39936
rect 9033 39933 9045 39936
rect 9079 39933 9091 39967
rect 9033 39927 9091 39933
rect 9214 39924 9220 39976
rect 9272 39924 9278 39976
rect 9674 39924 9680 39976
rect 9732 39964 9738 39976
rect 9732 39936 10272 39964
rect 9732 39924 9738 39936
rect 10244 39908 10272 39936
rect 9306 39856 9312 39908
rect 9364 39896 9370 39908
rect 9493 39899 9551 39905
rect 9493 39896 9505 39899
rect 9364 39868 9505 39896
rect 9364 39856 9370 39868
rect 9493 39865 9505 39868
rect 9539 39865 9551 39899
rect 9493 39859 9551 39865
rect 10134 39856 10140 39908
rect 10192 39856 10198 39908
rect 10226 39856 10232 39908
rect 10284 39896 10290 39908
rect 10413 39899 10471 39905
rect 10413 39896 10425 39899
rect 10284 39868 10425 39896
rect 10284 39856 10290 39868
rect 10413 39865 10425 39868
rect 10459 39865 10471 39899
rect 10413 39859 10471 39865
rect 7800 39800 8432 39828
rect 7800 39788 7806 39800
rect 9674 39788 9680 39840
rect 9732 39837 9738 39840
rect 9732 39831 9751 39837
rect 9739 39797 9751 39831
rect 9732 39791 9751 39797
rect 9732 39788 9738 39791
rect 9858 39788 9864 39840
rect 9916 39788 9922 39840
rect 10042 39788 10048 39840
rect 10100 39788 10106 39840
rect 10529 39828 10557 40004
rect 11238 39992 11244 40004
rect 11296 39992 11302 40044
rect 12250 39992 12256 40044
rect 12308 39992 12314 40044
rect 11054 39896 11060 39908
rect 10796 39868 11060 39896
rect 10796 39837 10824 39868
rect 11054 39856 11060 39868
rect 11112 39896 11118 39908
rect 11606 39896 11612 39908
rect 11112 39868 11612 39896
rect 11112 39856 11118 39868
rect 11606 39856 11612 39868
rect 11664 39856 11670 39908
rect 11882 39856 11888 39908
rect 11940 39896 11946 39908
rect 11986 39899 12044 39905
rect 11986 39896 11998 39899
rect 11940 39868 11998 39896
rect 11940 39856 11946 39868
rect 11986 39865 11998 39868
rect 12032 39865 12044 39899
rect 11986 39859 12044 39865
rect 10613 39831 10671 39837
rect 10613 39828 10625 39831
rect 10529 39800 10625 39828
rect 10613 39797 10625 39800
rect 10659 39797 10671 39831
rect 10613 39791 10671 39797
rect 10781 39831 10839 39837
rect 10781 39797 10793 39831
rect 10827 39797 10839 39831
rect 10781 39791 10839 39797
rect 10870 39788 10876 39840
rect 10928 39788 10934 39840
rect 11238 39788 11244 39840
rect 11296 39828 11302 39840
rect 12066 39828 12072 39840
rect 11296 39800 12072 39828
rect 11296 39788 11302 39800
rect 12066 39788 12072 39800
rect 12124 39788 12130 39840
rect 552 39738 12604 39760
rect 552 39686 4322 39738
rect 4374 39686 4386 39738
rect 4438 39686 4450 39738
rect 4502 39686 4514 39738
rect 4566 39686 4578 39738
rect 4630 39686 10722 39738
rect 10774 39686 10786 39738
rect 10838 39686 10850 39738
rect 10902 39686 10914 39738
rect 10966 39686 10978 39738
rect 11030 39686 12604 39738
rect 552 39664 12604 39686
rect 2774 39624 2780 39636
rect 1136 39596 2780 39624
rect 1136 39497 1164 39596
rect 2774 39584 2780 39596
rect 2832 39584 2838 39636
rect 3697 39627 3755 39633
rect 3697 39593 3709 39627
rect 3743 39624 3755 39627
rect 4706 39624 4712 39636
rect 3743 39596 4712 39624
rect 3743 39593 3755 39596
rect 3697 39587 3755 39593
rect 4706 39584 4712 39596
rect 4764 39584 4770 39636
rect 4982 39584 4988 39636
rect 5040 39624 5046 39636
rect 10226 39624 10232 39636
rect 5040 39596 8524 39624
rect 5040 39584 5046 39596
rect 2406 39556 2412 39568
rect 2056 39528 2412 39556
rect 1121 39491 1179 39497
rect 1121 39457 1133 39491
rect 1167 39457 1179 39491
rect 1121 39451 1179 39457
rect 1486 39448 1492 39500
rect 1544 39488 1550 39500
rect 1581 39491 1639 39497
rect 1581 39488 1593 39491
rect 1544 39460 1593 39488
rect 1544 39448 1550 39460
rect 1581 39457 1593 39460
rect 1627 39457 1639 39491
rect 1581 39451 1639 39457
rect 1854 39448 1860 39500
rect 1912 39448 1918 39500
rect 2056 39497 2084 39528
rect 2406 39516 2412 39528
rect 2464 39556 2470 39568
rect 2562 39559 2620 39565
rect 2562 39556 2574 39559
rect 2464 39528 2574 39556
rect 2464 39516 2470 39528
rect 2562 39525 2574 39528
rect 2608 39525 2620 39559
rect 5074 39556 5080 39568
rect 2562 39519 2620 39525
rect 2746 39528 5080 39556
rect 2041 39491 2099 39497
rect 2041 39457 2053 39491
rect 2087 39457 2099 39491
rect 2041 39451 2099 39457
rect 2314 39448 2320 39500
rect 2372 39448 2378 39500
rect 2746 39488 2774 39528
rect 5074 39516 5080 39528
rect 5132 39516 5138 39568
rect 5644 39528 8340 39556
rect 2424 39460 2774 39488
rect 658 39380 664 39432
rect 716 39420 722 39432
rect 716 39392 1532 39420
rect 716 39380 722 39392
rect 1394 39312 1400 39364
rect 1452 39312 1458 39364
rect 1504 39352 1532 39392
rect 1762 39380 1768 39432
rect 1820 39420 1826 39432
rect 2133 39423 2191 39429
rect 2133 39420 2145 39423
rect 1820 39392 2145 39420
rect 1820 39380 1826 39392
rect 2133 39389 2145 39392
rect 2179 39389 2191 39423
rect 2424 39420 2452 39460
rect 3050 39448 3056 39500
rect 3108 39488 3114 39500
rect 4065 39491 4123 39497
rect 4065 39488 4077 39491
rect 3108 39460 4077 39488
rect 3108 39448 3114 39460
rect 4065 39457 4077 39460
rect 4111 39457 4123 39491
rect 4065 39451 4123 39457
rect 4246 39448 4252 39500
rect 4304 39488 4310 39500
rect 4706 39488 4712 39500
rect 4304 39460 4712 39488
rect 4304 39448 4310 39460
rect 4706 39448 4712 39460
rect 4764 39448 4770 39500
rect 5644 39497 5672 39528
rect 5629 39491 5687 39497
rect 5629 39457 5641 39491
rect 5675 39457 5687 39491
rect 5629 39451 5687 39457
rect 6178 39448 6184 39500
rect 6236 39488 6242 39500
rect 6549 39491 6607 39497
rect 6549 39488 6561 39491
rect 6236 39460 6561 39488
rect 6236 39448 6242 39460
rect 6549 39457 6561 39460
rect 6595 39457 6607 39491
rect 6549 39451 6607 39457
rect 7742 39448 7748 39500
rect 7800 39448 7806 39500
rect 2133 39383 2191 39389
rect 2240 39392 2452 39420
rect 2240 39352 2268 39392
rect 3418 39380 3424 39432
rect 3476 39420 3482 39432
rect 4157 39423 4215 39429
rect 4157 39420 4169 39423
rect 3476 39392 4169 39420
rect 3476 39380 3482 39392
rect 4157 39389 4169 39392
rect 4203 39389 4215 39423
rect 4157 39383 4215 39389
rect 5902 39380 5908 39432
rect 5960 39380 5966 39432
rect 7101 39423 7159 39429
rect 7101 39389 7113 39423
rect 7147 39420 7159 39423
rect 7558 39420 7564 39432
rect 7147 39392 7564 39420
rect 7147 39389 7159 39392
rect 7101 39383 7159 39389
rect 7558 39380 7564 39392
rect 7616 39380 7622 39432
rect 7834 39380 7840 39432
rect 7892 39380 7898 39432
rect 8205 39423 8263 39429
rect 8205 39389 8217 39423
rect 8251 39389 8263 39423
rect 8312 39420 8340 39528
rect 8496 39497 8524 39596
rect 9078 39596 10232 39624
rect 8481 39491 8539 39497
rect 8481 39457 8493 39491
rect 8527 39457 8539 39491
rect 8481 39451 8539 39457
rect 8846 39448 8852 39500
rect 8904 39488 8910 39500
rect 9078 39497 9106 39596
rect 10226 39584 10232 39596
rect 10284 39624 10290 39636
rect 11146 39624 11152 39636
rect 10284 39596 11152 39624
rect 10284 39584 10290 39596
rect 11146 39584 11152 39596
rect 11204 39584 11210 39636
rect 9858 39516 9864 39568
rect 9916 39556 9922 39568
rect 11425 39559 11483 39565
rect 11425 39556 11437 39559
rect 9916 39528 11437 39556
rect 9916 39516 9922 39528
rect 11425 39525 11437 39528
rect 11471 39525 11483 39559
rect 12066 39556 12072 39568
rect 11425 39519 11483 39525
rect 11716 39528 12072 39556
rect 9063 39491 9121 39497
rect 9063 39488 9075 39491
rect 8904 39460 9075 39488
rect 8904 39448 8910 39460
rect 9063 39457 9075 39460
rect 9109 39457 9121 39491
rect 9063 39451 9121 39457
rect 9217 39491 9275 39497
rect 9217 39457 9229 39491
rect 9263 39457 9275 39491
rect 9217 39451 9275 39457
rect 9309 39491 9367 39497
rect 9309 39457 9321 39491
rect 9355 39488 9367 39491
rect 9398 39488 9404 39500
rect 9355 39460 9404 39488
rect 9355 39457 9367 39460
rect 9309 39451 9367 39457
rect 8665 39423 8723 39429
rect 8665 39420 8677 39423
rect 8312 39392 8677 39420
rect 8205 39383 8263 39389
rect 8665 39389 8677 39392
rect 8711 39389 8723 39423
rect 8665 39383 8723 39389
rect 1504 39324 2268 39352
rect 4062 39312 4068 39364
rect 4120 39352 4126 39364
rect 4985 39355 5043 39361
rect 4985 39352 4997 39355
rect 4120 39324 4997 39352
rect 4120 39312 4126 39324
rect 4985 39321 4997 39324
rect 5031 39321 5043 39355
rect 4985 39315 5043 39321
rect 6457 39355 6515 39361
rect 6457 39321 6469 39355
rect 6503 39352 6515 39355
rect 8220 39352 8248 39383
rect 6503 39324 8248 39352
rect 6503 39321 6515 39324
rect 6457 39315 6515 39321
rect 8570 39312 8576 39364
rect 8628 39352 8634 39364
rect 8849 39355 8907 39361
rect 8849 39352 8861 39355
rect 8628 39324 8861 39352
rect 8628 39312 8634 39324
rect 8849 39321 8861 39324
rect 8895 39321 8907 39355
rect 8849 39315 8907 39321
rect 934 39244 940 39296
rect 992 39244 998 39296
rect 1673 39287 1731 39293
rect 1673 39253 1685 39287
rect 1719 39284 1731 39287
rect 1946 39284 1952 39296
rect 1719 39256 1952 39284
rect 1719 39253 1731 39256
rect 1673 39247 1731 39253
rect 1946 39244 1952 39256
rect 2004 39244 2010 39296
rect 3050 39244 3056 39296
rect 3108 39284 3114 39296
rect 3881 39287 3939 39293
rect 3881 39284 3893 39287
rect 3108 39256 3893 39284
rect 3108 39244 3114 39256
rect 3881 39253 3893 39256
rect 3927 39253 3939 39287
rect 3881 39247 3939 39253
rect 4246 39244 4252 39296
rect 4304 39284 4310 39296
rect 4801 39287 4859 39293
rect 4801 39284 4813 39287
rect 4304 39256 4813 39284
rect 4304 39244 4310 39256
rect 4801 39253 4813 39256
rect 4847 39253 4859 39287
rect 4801 39247 4859 39253
rect 6638 39244 6644 39296
rect 6696 39284 6702 39296
rect 6733 39287 6791 39293
rect 6733 39284 6745 39287
rect 6696 39256 6745 39284
rect 6696 39244 6702 39256
rect 6733 39253 6745 39256
rect 6779 39253 6791 39287
rect 6733 39247 6791 39253
rect 7190 39244 7196 39296
rect 7248 39284 7254 39296
rect 7742 39284 7748 39296
rect 7248 39256 7748 39284
rect 7248 39244 7254 39256
rect 7742 39244 7748 39256
rect 7800 39244 7806 39296
rect 8202 39244 8208 39296
rect 8260 39284 8266 39296
rect 8297 39287 8355 39293
rect 8297 39284 8309 39287
rect 8260 39256 8309 39284
rect 8260 39244 8266 39256
rect 8297 39253 8309 39256
rect 8343 39253 8355 39287
rect 8297 39247 8355 39253
rect 8938 39244 8944 39296
rect 8996 39284 9002 39296
rect 9232 39284 9260 39451
rect 9398 39448 9404 39460
rect 9456 39448 9462 39500
rect 9576 39491 9634 39497
rect 9576 39457 9588 39491
rect 9622 39488 9634 39491
rect 9950 39488 9956 39500
rect 9622 39460 9956 39488
rect 9622 39457 9634 39460
rect 9576 39451 9634 39457
rect 9950 39448 9956 39460
rect 10008 39448 10014 39500
rect 10318 39448 10324 39500
rect 10376 39488 10382 39500
rect 11716 39497 11744 39528
rect 12066 39516 12072 39528
rect 12124 39516 12130 39568
rect 11701 39491 11759 39497
rect 10376 39460 11652 39488
rect 10376 39448 10382 39460
rect 11624 39432 11652 39460
rect 11701 39457 11713 39491
rect 11747 39457 11759 39491
rect 11701 39451 11759 39457
rect 11977 39491 12035 39497
rect 11977 39457 11989 39491
rect 12023 39457 12035 39491
rect 11977 39451 12035 39457
rect 11517 39423 11575 39429
rect 11517 39420 11529 39423
rect 10888 39392 11529 39420
rect 10686 39312 10692 39364
rect 10744 39312 10750 39364
rect 10888 39284 10916 39392
rect 11517 39389 11529 39392
rect 11563 39389 11575 39423
rect 11517 39383 11575 39389
rect 11149 39355 11207 39361
rect 11149 39321 11161 39355
rect 11195 39352 11207 39355
rect 11238 39352 11244 39364
rect 11195 39324 11244 39352
rect 11195 39321 11207 39324
rect 11149 39315 11207 39321
rect 11238 39312 11244 39324
rect 11296 39312 11302 39364
rect 11422 39312 11428 39364
rect 11480 39352 11486 39364
rect 11532 39352 11560 39383
rect 11606 39380 11612 39432
rect 11664 39420 11670 39432
rect 11992 39420 12020 39451
rect 11664 39392 12020 39420
rect 11664 39380 11670 39392
rect 11790 39352 11796 39364
rect 11480 39324 11796 39352
rect 11480 39312 11486 39324
rect 11790 39312 11796 39324
rect 11848 39312 11854 39364
rect 11885 39355 11943 39361
rect 11885 39321 11897 39355
rect 11931 39352 11943 39355
rect 12434 39352 12440 39364
rect 11931 39324 12440 39352
rect 11931 39321 11943 39324
rect 11885 39315 11943 39321
rect 12434 39312 12440 39324
rect 12492 39312 12498 39364
rect 8996 39256 10916 39284
rect 8996 39244 9002 39256
rect 10962 39244 10968 39296
rect 11020 39244 11026 39296
rect 12161 39287 12219 39293
rect 12161 39253 12173 39287
rect 12207 39284 12219 39287
rect 12342 39284 12348 39296
rect 12207 39256 12348 39284
rect 12207 39253 12219 39256
rect 12161 39247 12219 39253
rect 12342 39244 12348 39256
rect 12400 39244 12406 39296
rect 552 39194 12604 39216
rect 552 39142 3662 39194
rect 3714 39142 3726 39194
rect 3778 39142 3790 39194
rect 3842 39142 3854 39194
rect 3906 39142 3918 39194
rect 3970 39142 10062 39194
rect 10114 39142 10126 39194
rect 10178 39142 10190 39194
rect 10242 39142 10254 39194
rect 10306 39142 10318 39194
rect 10370 39142 12604 39194
rect 552 39120 12604 39142
rect 3053 39083 3111 39089
rect 3053 39049 3065 39083
rect 3099 39080 3111 39083
rect 3326 39080 3332 39092
rect 3099 39052 3332 39080
rect 3099 39049 3111 39052
rect 3053 39043 3111 39049
rect 3326 39040 3332 39052
rect 3384 39040 3390 39092
rect 3510 39040 3516 39092
rect 3568 39080 3574 39092
rect 3568 39052 8064 39080
rect 3568 39040 3574 39052
rect 934 38972 940 39024
rect 992 39012 998 39024
rect 992 38984 1348 39012
rect 992 38972 998 38984
rect 474 38836 480 38888
rect 532 38876 538 38888
rect 1121 38879 1179 38885
rect 1121 38876 1133 38879
rect 532 38848 1133 38876
rect 532 38836 538 38848
rect 1121 38845 1133 38848
rect 1167 38845 1179 38879
rect 1121 38839 1179 38845
rect 1213 38879 1271 38885
rect 1213 38845 1225 38879
rect 1259 38845 1271 38879
rect 1213 38839 1271 38845
rect 1228 38808 1256 38839
rect 1136 38780 1256 38808
rect 1320 38808 1348 38984
rect 3878 38972 3884 39024
rect 3936 38972 3942 39024
rect 7190 38972 7196 39024
rect 7248 38972 7254 39024
rect 7374 38972 7380 39024
rect 7432 39012 7438 39024
rect 7469 39015 7527 39021
rect 7469 39012 7481 39015
rect 7432 38984 7481 39012
rect 7432 38972 7438 38984
rect 7469 38981 7481 38984
rect 7515 38981 7527 39015
rect 8036 39012 8064 39052
rect 9858 39040 9864 39092
rect 9916 39040 9922 39092
rect 9950 39040 9956 39092
rect 10008 39040 10014 39092
rect 10505 39083 10563 39089
rect 10505 39049 10517 39083
rect 10551 39080 10563 39083
rect 10962 39080 10968 39092
rect 10551 39052 10968 39080
rect 10551 39049 10563 39052
rect 10505 39043 10563 39049
rect 10962 39040 10968 39052
rect 11020 39040 11026 39092
rect 8113 39015 8171 39021
rect 8113 39012 8125 39015
rect 8036 38984 8125 39012
rect 7469 38975 7527 38981
rect 8113 38981 8125 38984
rect 8159 38981 8171 39015
rect 8113 38975 8171 38981
rect 8294 38972 8300 39024
rect 8352 39012 8358 39024
rect 8757 39015 8815 39021
rect 8757 39012 8769 39015
rect 8352 38984 8769 39012
rect 8352 38972 8358 38984
rect 8757 38981 8769 38984
rect 8803 38981 8815 39015
rect 8757 38975 8815 38981
rect 9582 38972 9588 39024
rect 9640 38972 9646 39024
rect 9876 39012 9904 39040
rect 10042 39012 10048 39024
rect 9876 38984 10048 39012
rect 10042 38972 10048 38984
rect 10100 38972 10106 39024
rect 10594 38972 10600 39024
rect 10652 39012 10658 39024
rect 10652 38984 10824 39012
rect 10652 38972 10658 38984
rect 1581 38947 1639 38953
rect 1581 38913 1593 38947
rect 1627 38944 1639 38947
rect 1627 38916 1808 38944
rect 1627 38913 1639 38916
rect 1581 38907 1639 38913
rect 1394 38836 1400 38888
rect 1452 38836 1458 38888
rect 1673 38879 1731 38885
rect 1673 38876 1685 38879
rect 1504 38848 1685 38876
rect 1504 38808 1532 38848
rect 1673 38845 1685 38848
rect 1719 38845 1731 38879
rect 1780 38878 1808 38916
rect 2682 38904 2688 38956
rect 2740 38944 2746 38956
rect 3329 38947 3387 38953
rect 3329 38944 3341 38947
rect 2740 38916 3341 38944
rect 2740 38904 2746 38916
rect 3329 38913 3341 38916
rect 3375 38913 3387 38947
rect 4154 38944 4160 38956
rect 3329 38907 3387 38913
rect 4080 38916 4160 38944
rect 1780 38850 2084 38878
rect 1673 38839 1731 38845
rect 1946 38817 1952 38820
rect 1940 38808 1952 38817
rect 1320 38780 1532 38808
rect 1907 38780 1952 38808
rect 1136 38752 1164 38780
rect 1940 38771 1952 38780
rect 1946 38768 1952 38771
rect 2004 38768 2010 38820
rect 2056 38808 2084 38850
rect 2774 38836 2780 38888
rect 2832 38876 2838 38888
rect 3605 38879 3663 38885
rect 3605 38876 3617 38879
rect 2832 38848 3617 38876
rect 2832 38836 2838 38848
rect 3605 38845 3617 38848
rect 3651 38845 3663 38879
rect 3605 38839 3663 38845
rect 2130 38808 2136 38820
rect 2056 38780 2136 38808
rect 2130 38768 2136 38780
rect 2188 38768 2194 38820
rect 474 38700 480 38752
rect 532 38740 538 38752
rect 937 38743 995 38749
rect 937 38740 949 38743
rect 532 38712 949 38740
rect 532 38700 538 38712
rect 937 38709 949 38712
rect 983 38709 995 38743
rect 937 38703 995 38709
rect 1118 38700 1124 38752
rect 1176 38700 1182 38752
rect 3510 38700 3516 38752
rect 3568 38700 3574 38752
rect 3697 38743 3755 38749
rect 3697 38709 3709 38743
rect 3743 38740 3755 38743
rect 4080 38740 4108 38916
rect 4154 38904 4160 38916
rect 4212 38904 4218 38956
rect 5074 38904 5080 38956
rect 5132 38944 5138 38956
rect 5132 38916 5948 38944
rect 5132 38904 5138 38916
rect 5810 38876 5816 38888
rect 4172 38848 5816 38876
rect 4172 38820 4200 38848
rect 5810 38836 5816 38848
rect 5868 38836 5874 38888
rect 5920 38876 5948 38916
rect 7650 38904 7656 38956
rect 7708 38944 7714 38956
rect 8389 38947 8447 38953
rect 8389 38944 8401 38947
rect 7708 38916 8401 38944
rect 7708 38904 7714 38916
rect 8389 38913 8401 38916
rect 8435 38913 8447 38947
rect 8389 38907 8447 38913
rect 8662 38904 8668 38956
rect 8720 38904 8726 38956
rect 9490 38904 9496 38956
rect 9548 38944 9554 38956
rect 10796 38953 10824 38984
rect 10781 38947 10839 38953
rect 10781 38944 10793 38947
rect 9548 38916 10793 38944
rect 9548 38904 9554 38916
rect 10781 38913 10793 38916
rect 10827 38913 10839 38947
rect 10781 38907 10839 38913
rect 7285 38879 7343 38885
rect 7285 38876 7297 38879
rect 5920 38848 7297 38876
rect 7285 38845 7297 38848
rect 7331 38845 7343 38879
rect 7285 38839 7343 38845
rect 7742 38836 7748 38888
rect 7800 38876 7806 38888
rect 7929 38879 7987 38885
rect 7929 38876 7941 38879
rect 7800 38848 7941 38876
rect 7800 38836 7806 38848
rect 7929 38845 7941 38848
rect 7975 38845 7987 38879
rect 7929 38839 7987 38845
rect 8018 38836 8024 38888
rect 8076 38876 8082 38888
rect 8573 38879 8631 38885
rect 8573 38876 8585 38879
rect 8076 38848 8585 38876
rect 8076 38836 8082 38848
rect 8573 38845 8585 38848
rect 8619 38845 8631 38879
rect 8573 38839 8631 38845
rect 8754 38836 8760 38888
rect 8812 38876 8818 38888
rect 8849 38879 8907 38885
rect 8849 38876 8861 38879
rect 8812 38848 8861 38876
rect 8812 38836 8818 38848
rect 8849 38845 8861 38848
rect 8895 38845 8907 38879
rect 9401 38879 9459 38885
rect 9401 38876 9413 38879
rect 8849 38839 8907 38845
rect 8956 38848 9413 38876
rect 4154 38768 4160 38820
rect 4212 38768 4218 38820
rect 6086 38817 6092 38820
rect 5721 38811 5779 38817
rect 5721 38777 5733 38811
rect 5767 38777 5779 38811
rect 5721 38771 5779 38777
rect 6080 38771 6092 38817
rect 5074 38740 5080 38752
rect 3743 38712 5080 38740
rect 3743 38709 3755 38712
rect 3697 38703 3755 38709
rect 5074 38700 5080 38712
rect 5132 38700 5138 38752
rect 5736 38740 5764 38771
rect 6086 38768 6092 38771
rect 6144 38768 6150 38820
rect 7558 38768 7564 38820
rect 7616 38808 7622 38820
rect 8956 38808 8984 38848
rect 9401 38845 9413 38848
rect 9447 38845 9459 38879
rect 9401 38839 9459 38845
rect 9766 38836 9772 38888
rect 9824 38876 9830 38888
rect 10078 38879 10136 38885
rect 10078 38876 10090 38879
rect 9824 38848 10090 38876
rect 9824 38836 9830 38848
rect 10078 38845 10090 38848
rect 10124 38845 10136 38879
rect 10078 38839 10136 38845
rect 10318 38836 10324 38888
rect 10376 38876 10382 38888
rect 10597 38879 10655 38885
rect 10597 38876 10609 38879
rect 10376 38848 10609 38876
rect 10376 38836 10382 38848
rect 10597 38845 10609 38848
rect 10643 38845 10655 38879
rect 10597 38839 10655 38845
rect 7616 38780 8984 38808
rect 7616 38768 7622 38780
rect 9030 38768 9036 38820
rect 9088 38768 9094 38820
rect 11048 38811 11106 38817
rect 9416 38780 10456 38808
rect 9416 38752 9444 38780
rect 10428 38752 10456 38780
rect 11048 38777 11060 38811
rect 11094 38808 11106 38811
rect 11882 38808 11888 38820
rect 11094 38780 11888 38808
rect 11094 38777 11106 38780
rect 11048 38771 11106 38777
rect 11882 38768 11888 38780
rect 11940 38768 11946 38820
rect 7190 38740 7196 38752
rect 5736 38712 7196 38740
rect 7190 38700 7196 38712
rect 7248 38700 7254 38752
rect 7374 38700 7380 38752
rect 7432 38740 7438 38752
rect 7650 38740 7656 38752
rect 7432 38712 7656 38740
rect 7432 38700 7438 38712
rect 7650 38700 7656 38712
rect 7708 38700 7714 38752
rect 7742 38700 7748 38752
rect 7800 38740 7806 38752
rect 7837 38743 7895 38749
rect 7837 38740 7849 38743
rect 7800 38712 7849 38740
rect 7800 38700 7806 38712
rect 7837 38709 7849 38712
rect 7883 38740 7895 38743
rect 8018 38740 8024 38752
rect 7883 38712 8024 38740
rect 7883 38709 7895 38712
rect 7837 38703 7895 38709
rect 8018 38700 8024 38712
rect 8076 38700 8082 38752
rect 8938 38700 8944 38752
rect 8996 38740 9002 38752
rect 9217 38743 9275 38749
rect 9217 38740 9229 38743
rect 8996 38712 9229 38740
rect 8996 38700 9002 38712
rect 9217 38709 9229 38712
rect 9263 38709 9275 38743
rect 9217 38703 9275 38709
rect 9306 38700 9312 38752
rect 9364 38700 9370 38752
rect 9398 38700 9404 38752
rect 9456 38700 9462 38752
rect 10134 38700 10140 38752
rect 10192 38700 10198 38752
rect 10410 38700 10416 38752
rect 10468 38740 10474 38752
rect 11974 38740 11980 38752
rect 10468 38712 11980 38740
rect 10468 38700 10474 38712
rect 11974 38700 11980 38712
rect 12032 38740 12038 38752
rect 12161 38743 12219 38749
rect 12161 38740 12173 38743
rect 12032 38712 12173 38740
rect 12032 38700 12038 38712
rect 12161 38709 12173 38712
rect 12207 38740 12219 38743
rect 12250 38740 12256 38752
rect 12207 38712 12256 38740
rect 12207 38709 12219 38712
rect 12161 38703 12219 38709
rect 12250 38700 12256 38712
rect 12308 38700 12314 38752
rect 552 38650 12604 38672
rect 552 38598 4322 38650
rect 4374 38598 4386 38650
rect 4438 38598 4450 38650
rect 4502 38598 4514 38650
rect 4566 38598 4578 38650
rect 4630 38598 10722 38650
rect 10774 38598 10786 38650
rect 10838 38598 10850 38650
rect 10902 38598 10914 38650
rect 10966 38598 10978 38650
rect 11030 38598 12604 38650
rect 552 38576 12604 38598
rect 1394 38496 1400 38548
rect 1452 38536 1458 38548
rect 2222 38536 2228 38548
rect 1452 38508 2228 38536
rect 1452 38496 1458 38508
rect 2222 38496 2228 38508
rect 2280 38496 2286 38548
rect 2314 38496 2320 38548
rect 2372 38536 2378 38548
rect 4154 38536 4160 38548
rect 2372 38508 4160 38536
rect 2372 38496 2378 38508
rect 290 38428 296 38480
rect 348 38468 354 38480
rect 1670 38468 1676 38480
rect 348 38440 1676 38468
rect 348 38428 354 38440
rect 1670 38428 1676 38440
rect 1728 38428 1734 38480
rect 2332 38468 2360 38496
rect 2056 38440 2360 38468
rect 1397 38403 1455 38409
rect 1397 38369 1409 38403
rect 1443 38400 1455 38403
rect 1486 38400 1492 38412
rect 1443 38372 1492 38400
rect 1443 38369 1455 38372
rect 1397 38363 1455 38369
rect 1486 38360 1492 38372
rect 1544 38360 1550 38412
rect 1581 38403 1639 38409
rect 1581 38369 1593 38403
rect 1627 38400 1639 38403
rect 1946 38400 1952 38412
rect 1627 38372 1952 38400
rect 1627 38369 1639 38372
rect 1581 38363 1639 38369
rect 1946 38360 1952 38372
rect 2004 38360 2010 38412
rect 2056 38409 2084 38440
rect 3804 38412 3832 38508
rect 4154 38496 4160 38508
rect 4212 38496 4218 38548
rect 4338 38496 4344 38548
rect 4396 38536 4402 38548
rect 4890 38536 4896 38548
rect 4396 38508 4896 38536
rect 4396 38496 4402 38508
rect 4890 38496 4896 38508
rect 4948 38496 4954 38548
rect 5169 38539 5227 38545
rect 5169 38505 5181 38539
rect 5215 38536 5227 38539
rect 5258 38536 5264 38548
rect 5215 38508 5264 38536
rect 5215 38505 5227 38508
rect 5169 38499 5227 38505
rect 5258 38496 5264 38508
rect 5316 38496 5322 38548
rect 7193 38539 7251 38545
rect 7193 38505 7205 38539
rect 7239 38505 7251 38539
rect 7193 38499 7251 38505
rect 8389 38539 8447 38545
rect 8389 38505 8401 38539
rect 8435 38536 8447 38539
rect 9030 38536 9036 38548
rect 8435 38508 9036 38536
rect 8435 38505 8447 38508
rect 8389 38499 8447 38505
rect 3896 38440 5304 38468
rect 2041 38403 2099 38409
rect 2041 38369 2053 38403
rect 2087 38369 2099 38403
rect 2041 38363 2099 38369
rect 2130 38360 2136 38412
rect 2188 38400 2194 38412
rect 2297 38403 2355 38409
rect 2297 38400 2309 38403
rect 2188 38372 2309 38400
rect 2188 38360 2194 38372
rect 2297 38369 2309 38372
rect 2343 38369 2355 38403
rect 2297 38363 2355 38369
rect 3513 38403 3571 38409
rect 3513 38369 3525 38403
rect 3559 38369 3571 38403
rect 3513 38363 3571 38369
rect 934 38292 940 38344
rect 992 38292 998 38344
rect 1673 38335 1731 38341
rect 1673 38301 1685 38335
rect 1719 38301 1731 38335
rect 3528 38332 3556 38363
rect 3694 38360 3700 38412
rect 3752 38360 3758 38412
rect 3786 38360 3792 38412
rect 3844 38360 3850 38412
rect 3896 38332 3924 38440
rect 4062 38409 4068 38412
rect 4056 38363 4068 38409
rect 4062 38360 4068 38363
rect 4120 38360 4126 38412
rect 4430 38360 4436 38412
rect 4488 38400 4494 38412
rect 5276 38400 5304 38440
rect 5350 38428 5356 38480
rect 5408 38468 5414 38480
rect 6058 38471 6116 38477
rect 6058 38468 6070 38471
rect 5408 38440 6070 38468
rect 5408 38428 5414 38440
rect 6058 38437 6070 38440
rect 6104 38437 6116 38471
rect 6058 38431 6116 38437
rect 6454 38428 6460 38480
rect 6512 38468 6518 38480
rect 7208 38468 7236 38499
rect 9030 38496 9036 38508
rect 9088 38496 9094 38548
rect 9306 38536 9312 38548
rect 9133 38508 9312 38536
rect 9133 38468 9161 38508
rect 9306 38496 9312 38508
rect 9364 38496 9370 38548
rect 10226 38536 10232 38548
rect 9600 38508 10232 38536
rect 6512 38440 9161 38468
rect 6512 38428 6518 38440
rect 9600 38412 9628 38508
rect 10226 38496 10232 38508
rect 10284 38496 10290 38548
rect 10502 38496 10508 38548
rect 10560 38536 10566 38548
rect 10560 38508 11100 38536
rect 10560 38496 10566 38508
rect 10410 38468 10416 38480
rect 10152 38440 10416 38468
rect 5445 38403 5503 38409
rect 4488 38372 4844 38400
rect 5276 38372 5396 38400
rect 4488 38360 4494 38372
rect 4816 38344 4844 38372
rect 3528 38304 3924 38332
rect 1673 38295 1731 38301
rect 1688 38196 1716 38295
rect 4798 38292 4804 38344
rect 4856 38332 4862 38344
rect 5261 38335 5319 38341
rect 5261 38332 5273 38335
rect 4856 38304 5273 38332
rect 4856 38292 4862 38304
rect 5261 38301 5273 38304
rect 5307 38301 5319 38335
rect 5261 38295 5319 38301
rect 3418 38224 3424 38276
rect 3476 38224 3482 38276
rect 5368 38264 5396 38372
rect 5445 38369 5457 38403
rect 5491 38369 5503 38403
rect 5445 38363 5503 38369
rect 5460 38332 5488 38363
rect 5534 38360 5540 38412
rect 5592 38360 5598 38412
rect 5810 38360 5816 38412
rect 5868 38360 5874 38412
rect 7926 38360 7932 38412
rect 7984 38400 7990 38412
rect 8205 38403 8263 38409
rect 8205 38400 8217 38403
rect 7984 38372 8217 38400
rect 7984 38360 7990 38372
rect 8205 38369 8217 38372
rect 8251 38369 8263 38403
rect 9030 38400 9036 38412
rect 8205 38363 8263 38369
rect 8496 38372 9036 38400
rect 5626 38332 5632 38344
rect 5460 38304 5632 38332
rect 5626 38292 5632 38304
rect 5684 38292 5690 38344
rect 7098 38292 7104 38344
rect 7156 38332 7162 38344
rect 7285 38335 7343 38341
rect 7285 38332 7297 38335
rect 7156 38304 7297 38332
rect 7156 38292 7162 38304
rect 7285 38301 7297 38304
rect 7331 38301 7343 38335
rect 7285 38295 7343 38301
rect 7834 38292 7840 38344
rect 7892 38332 7898 38344
rect 8021 38335 8079 38341
rect 8021 38332 8033 38335
rect 7892 38304 8033 38332
rect 7892 38292 7898 38304
rect 8021 38301 8033 38304
rect 8067 38332 8079 38335
rect 8294 38332 8300 38344
rect 8067 38304 8300 38332
rect 8067 38301 8079 38304
rect 8021 38295 8079 38301
rect 8294 38292 8300 38304
rect 8352 38332 8358 38344
rect 8496 38332 8524 38372
rect 9030 38360 9036 38372
rect 9088 38360 9094 38412
rect 9309 38403 9367 38409
rect 9309 38369 9321 38403
rect 9355 38398 9367 38403
rect 9416 38398 9536 38400
rect 9355 38372 9536 38398
rect 9355 38370 9444 38372
rect 9355 38369 9367 38370
rect 9309 38363 9367 38369
rect 8352 38304 8524 38332
rect 8352 38292 8358 38304
rect 8662 38292 8668 38344
rect 8720 38332 8726 38344
rect 8757 38335 8815 38341
rect 8757 38332 8769 38335
rect 8720 38304 8769 38332
rect 8720 38292 8726 38304
rect 8757 38301 8769 38304
rect 8803 38332 8815 38335
rect 9401 38335 9459 38341
rect 9401 38332 9413 38335
rect 8803 38304 9413 38332
rect 8803 38301 8815 38304
rect 8757 38295 8815 38301
rect 9401 38301 9413 38304
rect 9447 38301 9459 38335
rect 9508 38332 9536 38372
rect 9582 38360 9588 38412
rect 9640 38360 9646 38412
rect 9766 38360 9772 38412
rect 9824 38360 9830 38412
rect 9858 38360 9864 38412
rect 9916 38400 9922 38412
rect 10042 38400 10048 38412
rect 9916 38372 10048 38400
rect 9916 38360 9922 38372
rect 10042 38360 10048 38372
rect 10100 38360 10106 38412
rect 10152 38409 10180 38440
rect 10410 38428 10416 38440
rect 10468 38428 10474 38480
rect 10594 38428 10600 38480
rect 10652 38477 10658 38480
rect 10652 38471 10671 38477
rect 10659 38437 10671 38471
rect 10652 38431 10671 38437
rect 10652 38428 10658 38431
rect 10962 38428 10968 38480
rect 11020 38428 11026 38480
rect 11072 38468 11100 38508
rect 11146 38496 11152 38548
rect 11204 38536 11210 38548
rect 11333 38539 11391 38545
rect 11333 38536 11345 38539
rect 11204 38508 11345 38536
rect 11204 38496 11210 38508
rect 11333 38505 11345 38508
rect 11379 38536 11391 38539
rect 11698 38536 11704 38548
rect 11379 38508 11704 38536
rect 11379 38505 11391 38508
rect 11333 38499 11391 38505
rect 11698 38496 11704 38508
rect 11756 38496 11762 38548
rect 11977 38471 12035 38477
rect 11977 38468 11989 38471
rect 11072 38440 11989 38468
rect 11977 38437 11989 38440
rect 12023 38468 12035 38471
rect 12023 38440 12296 38468
rect 12023 38437 12035 38440
rect 11977 38431 12035 38437
rect 10137 38403 10195 38409
rect 10137 38369 10149 38403
rect 10183 38369 10195 38403
rect 10137 38363 10195 38369
rect 11149 38403 11207 38409
rect 11149 38369 11161 38403
rect 11195 38369 11207 38403
rect 11149 38363 11207 38369
rect 9784 38332 9812 38360
rect 11164 38332 11192 38363
rect 11238 38360 11244 38412
rect 11296 38360 11302 38412
rect 11793 38403 11851 38409
rect 11793 38369 11805 38403
rect 11839 38400 11851 38403
rect 11839 38372 11912 38400
rect 11839 38369 11851 38372
rect 11793 38363 11851 38369
rect 11422 38332 11428 38344
rect 9508 38304 9812 38332
rect 10612 38304 11428 38332
rect 9401 38295 9459 38301
rect 5810 38264 5816 38276
rect 5368 38236 5816 38264
rect 5810 38224 5816 38236
rect 5868 38224 5874 38276
rect 7742 38224 7748 38276
rect 7800 38264 7806 38276
rect 8481 38267 8539 38273
rect 8481 38264 8493 38267
rect 7800 38236 8493 38264
rect 7800 38224 7806 38236
rect 8481 38233 8493 38236
rect 8527 38233 8539 38267
rect 8481 38227 8539 38233
rect 8570 38224 8576 38276
rect 8628 38264 8634 38276
rect 9125 38267 9183 38273
rect 9125 38264 9137 38267
rect 8628 38236 9137 38264
rect 8628 38224 8634 38236
rect 9125 38233 9137 38236
rect 9171 38233 9183 38267
rect 9493 38267 9551 38273
rect 9493 38264 9505 38267
rect 9125 38227 9183 38233
rect 9232 38236 9505 38264
rect 3234 38196 3240 38208
rect 1688 38168 3240 38196
rect 3234 38156 3240 38168
rect 3292 38156 3298 38208
rect 3605 38199 3663 38205
rect 3605 38165 3617 38199
rect 3651 38196 3663 38199
rect 7098 38196 7104 38208
rect 3651 38168 7104 38196
rect 3651 38165 3663 38168
rect 3605 38159 3663 38165
rect 7098 38156 7104 38168
rect 7156 38156 7162 38208
rect 7650 38156 7656 38208
rect 7708 38196 7714 38208
rect 7929 38199 7987 38205
rect 7929 38196 7941 38199
rect 7708 38168 7941 38196
rect 7708 38156 7714 38168
rect 7929 38165 7941 38168
rect 7975 38165 7987 38199
rect 7929 38159 7987 38165
rect 8662 38156 8668 38208
rect 8720 38156 8726 38208
rect 8754 38156 8760 38208
rect 8812 38196 8818 38208
rect 9232 38196 9260 38236
rect 9493 38233 9505 38236
rect 9539 38233 9551 38267
rect 9493 38227 9551 38233
rect 8812 38168 9260 38196
rect 8812 38156 8818 38168
rect 9398 38156 9404 38208
rect 9456 38196 9462 38208
rect 9861 38199 9919 38205
rect 9861 38196 9873 38199
rect 9456 38168 9873 38196
rect 9456 38156 9462 38168
rect 9861 38165 9873 38168
rect 9907 38165 9919 38199
rect 9861 38159 9919 38165
rect 10321 38199 10379 38205
rect 10321 38165 10333 38199
rect 10367 38196 10379 38199
rect 10502 38196 10508 38208
rect 10367 38168 10508 38196
rect 10367 38165 10379 38168
rect 10321 38159 10379 38165
rect 10502 38156 10508 38168
rect 10560 38156 10566 38208
rect 10612 38205 10640 38304
rect 11422 38292 11428 38304
rect 11480 38292 11486 38344
rect 11609 38335 11667 38341
rect 11609 38301 11621 38335
rect 11655 38332 11667 38335
rect 11884 38332 11912 38372
rect 12066 38360 12072 38412
rect 12124 38360 12130 38412
rect 12268 38409 12296 38440
rect 12253 38403 12311 38409
rect 12253 38369 12265 38403
rect 12299 38369 12311 38403
rect 12253 38363 12311 38369
rect 12710 38332 12716 38344
rect 11655 38304 11836 38332
rect 11884 38304 12716 38332
rect 11655 38301 11667 38304
rect 11609 38295 11667 38301
rect 11808 38276 11836 38304
rect 12710 38292 12716 38304
rect 12768 38292 12774 38344
rect 10686 38224 10692 38276
rect 10744 38264 10750 38276
rect 10744 38236 10916 38264
rect 10744 38224 10750 38236
rect 10597 38199 10655 38205
rect 10597 38165 10609 38199
rect 10643 38165 10655 38199
rect 10597 38159 10655 38165
rect 10778 38156 10784 38208
rect 10836 38156 10842 38208
rect 10888 38196 10916 38236
rect 11146 38224 11152 38276
rect 11204 38264 11210 38276
rect 11517 38267 11575 38273
rect 11517 38264 11529 38267
rect 11204 38236 11529 38264
rect 11204 38224 11210 38236
rect 11517 38233 11529 38236
rect 11563 38233 11575 38267
rect 11517 38227 11575 38233
rect 11790 38224 11796 38276
rect 11848 38224 11854 38276
rect 12161 38199 12219 38205
rect 12161 38196 12173 38199
rect 10888 38168 12173 38196
rect 12161 38165 12173 38168
rect 12207 38165 12219 38199
rect 12161 38159 12219 38165
rect 552 38106 12604 38128
rect 552 38054 3662 38106
rect 3714 38054 3726 38106
rect 3778 38054 3790 38106
rect 3842 38054 3854 38106
rect 3906 38054 3918 38106
rect 3970 38054 10062 38106
rect 10114 38054 10126 38106
rect 10178 38054 10190 38106
rect 10242 38054 10254 38106
rect 10306 38054 10318 38106
rect 10370 38054 12604 38106
rect 552 38032 12604 38054
rect 1026 37952 1032 38004
rect 1084 37992 1090 38004
rect 2038 37992 2044 38004
rect 1084 37964 2044 37992
rect 1084 37952 1090 37964
rect 2038 37952 2044 37964
rect 2096 37952 2102 38004
rect 3970 37952 3976 38004
rect 4028 37992 4034 38004
rect 4706 37992 4712 38004
rect 4028 37964 4712 37992
rect 4028 37952 4034 37964
rect 4706 37952 4712 37964
rect 4764 37952 4770 38004
rect 4801 37995 4859 38001
rect 4801 37961 4813 37995
rect 4847 37992 4859 37995
rect 5258 37992 5264 38004
rect 4847 37964 5264 37992
rect 4847 37961 4859 37964
rect 4801 37955 4859 37961
rect 5258 37952 5264 37964
rect 5316 37952 5322 38004
rect 5350 37952 5356 38004
rect 5408 37992 5414 38004
rect 5537 37995 5595 38001
rect 5537 37992 5549 37995
rect 5408 37964 5549 37992
rect 5408 37952 5414 37964
rect 5537 37961 5549 37964
rect 5583 37961 5595 37995
rect 5537 37955 5595 37961
rect 6365 37995 6423 38001
rect 6365 37961 6377 37995
rect 6411 37992 6423 37995
rect 6822 37992 6828 38004
rect 6411 37964 6828 37992
rect 6411 37961 6423 37964
rect 6365 37955 6423 37961
rect 6822 37952 6828 37964
rect 6880 37952 6886 38004
rect 7098 37952 7104 38004
rect 7156 37992 7162 38004
rect 9309 37995 9367 38001
rect 7156 37964 8708 37992
rect 7156 37952 7162 37964
rect 2866 37884 2872 37936
rect 2924 37924 2930 37936
rect 3237 37927 3295 37933
rect 3237 37924 3249 37927
rect 2924 37896 3249 37924
rect 2924 37884 2930 37896
rect 3237 37893 3249 37896
rect 3283 37893 3295 37927
rect 4522 37924 4528 37936
rect 3237 37887 3295 37893
rect 3896 37896 4528 37924
rect 2590 37816 2596 37868
rect 2648 37816 2654 37868
rect 3053 37859 3111 37865
rect 3053 37825 3065 37859
rect 3099 37856 3111 37859
rect 3326 37856 3332 37868
rect 3099 37828 3332 37856
rect 3099 37825 3111 37828
rect 3053 37819 3111 37825
rect 3326 37816 3332 37828
rect 3384 37816 3390 37868
rect 3896 37865 3924 37896
rect 4522 37884 4528 37896
rect 4580 37924 4586 37936
rect 5442 37924 5448 37936
rect 4580 37896 5448 37924
rect 4580 37884 4586 37896
rect 5442 37884 5448 37896
rect 5500 37884 5506 37936
rect 5629 37927 5687 37933
rect 5629 37893 5641 37927
rect 5675 37924 5687 37927
rect 6086 37924 6092 37936
rect 5675 37896 6092 37924
rect 5675 37893 5687 37896
rect 5629 37887 5687 37893
rect 6086 37884 6092 37896
rect 6144 37884 6150 37936
rect 8680 37933 8708 37964
rect 9309 37961 9321 37995
rect 9355 37992 9367 37995
rect 9355 37964 11183 37992
rect 9355 37961 9367 37964
rect 9309 37955 9367 37961
rect 8665 37927 8723 37933
rect 8665 37893 8677 37927
rect 8711 37893 8723 37927
rect 11155 37924 11183 37964
rect 11238 37952 11244 38004
rect 11296 37992 11302 38004
rect 11790 37992 11796 38004
rect 11296 37964 11796 37992
rect 11296 37952 11302 37964
rect 11790 37952 11796 37964
rect 11848 37952 11854 38004
rect 12618 37924 12624 37936
rect 11155 37896 12624 37924
rect 8665 37887 8723 37893
rect 12618 37884 12624 37896
rect 12676 37884 12682 37936
rect 3881 37859 3939 37865
rect 3881 37825 3893 37859
rect 3927 37825 3939 37859
rect 3881 37819 3939 37825
rect 7668 37828 8432 37856
rect 845 37791 903 37797
rect 845 37757 857 37791
rect 891 37788 903 37791
rect 1578 37788 1584 37800
rect 891 37760 1584 37788
rect 891 37757 903 37760
rect 845 37751 903 37757
rect 1578 37748 1584 37760
rect 1636 37748 1642 37800
rect 2498 37748 2504 37800
rect 2556 37788 2562 37800
rect 2685 37791 2743 37797
rect 2685 37788 2697 37791
rect 2556 37760 2697 37788
rect 2556 37748 2562 37760
rect 2685 37757 2697 37760
rect 2731 37757 2743 37791
rect 3786 37788 3792 37800
rect 2685 37751 2743 37757
rect 2792 37760 3792 37788
rect 1118 37729 1124 37732
rect 1112 37720 1124 37729
rect 1079 37692 1124 37720
rect 1112 37683 1124 37692
rect 1118 37680 1124 37683
rect 1176 37680 1182 37732
rect 1670 37680 1676 37732
rect 1728 37720 1734 37732
rect 2792 37720 2820 37760
rect 3786 37748 3792 37760
rect 3844 37748 3850 37800
rect 3970 37748 3976 37800
rect 4028 37788 4034 37800
rect 4157 37791 4215 37797
rect 4157 37788 4169 37791
rect 4028 37760 4169 37788
rect 4028 37748 4034 37760
rect 4157 37757 4169 37760
rect 4203 37757 4215 37791
rect 4157 37751 4215 37757
rect 4246 37748 4252 37800
rect 4304 37788 4310 37800
rect 4663 37791 4721 37797
rect 4304 37760 4349 37788
rect 4304 37748 4310 37760
rect 4663 37757 4675 37791
rect 4709 37790 4721 37791
rect 4798 37790 4804 37800
rect 4709 37762 4804 37790
rect 4709 37757 4721 37762
rect 4663 37751 4721 37757
rect 4798 37748 4804 37762
rect 4856 37748 4862 37800
rect 4985 37791 5043 37797
rect 4985 37757 4997 37791
rect 5031 37788 5043 37791
rect 5350 37788 5356 37800
rect 5031 37760 5356 37788
rect 5031 37757 5043 37760
rect 4985 37751 5043 37757
rect 5350 37748 5356 37760
rect 5408 37748 5414 37800
rect 6273 37791 6331 37797
rect 6273 37757 6285 37791
rect 6319 37788 6331 37791
rect 6638 37788 6644 37800
rect 6319 37760 6644 37788
rect 6319 37757 6331 37760
rect 6273 37751 6331 37757
rect 6638 37748 6644 37760
rect 6696 37748 6702 37800
rect 6914 37748 6920 37800
rect 6972 37788 6978 37800
rect 7668 37788 7696 37828
rect 6972 37760 7696 37788
rect 7745 37791 7803 37797
rect 6972 37748 6978 37760
rect 7745 37757 7757 37791
rect 7791 37788 7803 37791
rect 8021 37791 8079 37797
rect 7791 37760 7972 37788
rect 7791 37757 7803 37760
rect 7745 37751 7803 37757
rect 3050 37720 3056 37732
rect 1728 37692 2820 37720
rect 2884 37692 3056 37720
rect 1728 37680 1734 37692
rect 2884 37664 2912 37692
rect 3050 37680 3056 37692
rect 3108 37720 3114 37732
rect 3108 37692 4293 37720
rect 3108 37680 3114 37692
rect 1210 37612 1216 37664
rect 1268 37652 1274 37664
rect 1854 37652 1860 37664
rect 1268 37624 1860 37652
rect 1268 37612 1274 37624
rect 1854 37612 1860 37624
rect 1912 37612 1918 37664
rect 2222 37612 2228 37664
rect 2280 37612 2286 37664
rect 2866 37612 2872 37664
rect 2924 37612 2930 37664
rect 3510 37612 3516 37664
rect 3568 37652 3574 37664
rect 3605 37655 3663 37661
rect 3605 37652 3617 37655
rect 3568 37624 3617 37652
rect 3568 37612 3574 37624
rect 3605 37621 3617 37624
rect 3651 37621 3663 37655
rect 3605 37615 3663 37621
rect 3694 37612 3700 37664
rect 3752 37612 3758 37664
rect 4265 37652 4293 37692
rect 4430 37680 4436 37732
rect 4488 37680 4494 37732
rect 4522 37680 4528 37732
rect 4580 37680 4586 37732
rect 5534 37680 5540 37732
rect 5592 37720 5598 37732
rect 7098 37720 7104 37732
rect 5592 37692 7104 37720
rect 5592 37680 5598 37692
rect 7098 37680 7104 37692
rect 7156 37680 7162 37732
rect 7190 37680 7196 37732
rect 7248 37720 7254 37732
rect 7478 37723 7536 37729
rect 7478 37720 7490 37723
rect 7248 37692 7490 37720
rect 7248 37680 7254 37692
rect 7478 37689 7490 37692
rect 7524 37689 7536 37723
rect 7478 37683 7536 37689
rect 4614 37652 4620 37664
rect 4265 37624 4620 37652
rect 4614 37612 4620 37624
rect 4672 37612 4678 37664
rect 5718 37612 5724 37664
rect 5776 37652 5782 37664
rect 5902 37652 5908 37664
rect 5776 37624 5908 37652
rect 5776 37612 5782 37624
rect 5902 37612 5908 37624
rect 5960 37612 5966 37664
rect 7834 37612 7840 37664
rect 7892 37612 7898 37664
rect 7944 37652 7972 37760
rect 8021 37757 8033 37791
rect 8067 37757 8079 37791
rect 8021 37751 8079 37757
rect 8036 37720 8064 37751
rect 8202 37748 8208 37800
rect 8260 37748 8266 37800
rect 8404 37797 8432 37828
rect 9048 37828 9628 37856
rect 8389 37791 8447 37797
rect 8389 37757 8401 37791
rect 8435 37788 8447 37791
rect 8478 37788 8484 37800
rect 8435 37760 8484 37788
rect 8435 37757 8447 37760
rect 8389 37751 8447 37757
rect 8478 37748 8484 37760
rect 8536 37748 8542 37800
rect 8570 37748 8576 37800
rect 8628 37748 8634 37800
rect 8662 37748 8668 37800
rect 8720 37788 8726 37800
rect 8757 37791 8815 37797
rect 8757 37788 8769 37791
rect 8720 37760 8769 37788
rect 8720 37748 8726 37760
rect 8757 37757 8769 37760
rect 8803 37757 8815 37791
rect 8757 37751 8815 37757
rect 8849 37791 8907 37797
rect 8849 37757 8861 37791
rect 8895 37788 8907 37791
rect 8938 37788 8944 37800
rect 8895 37760 8944 37788
rect 8895 37757 8907 37760
rect 8849 37751 8907 37757
rect 8938 37748 8944 37760
rect 8996 37748 9002 37800
rect 8588 37720 8616 37748
rect 9048 37720 9076 37828
rect 9600 37800 9628 37828
rect 10778 37816 10784 37868
rect 10836 37856 10842 37868
rect 10836 37828 11928 37856
rect 10836 37816 10842 37828
rect 9125 37791 9183 37797
rect 9125 37757 9137 37791
rect 9171 37788 9183 37791
rect 9214 37788 9220 37800
rect 9171 37760 9220 37788
rect 9171 37757 9183 37760
rect 9125 37751 9183 37757
rect 9214 37748 9220 37760
rect 9272 37748 9278 37800
rect 9582 37748 9588 37800
rect 9640 37748 9646 37800
rect 11790 37748 11796 37800
rect 11848 37748 11854 37800
rect 11900 37797 11928 37828
rect 11885 37791 11943 37797
rect 11885 37757 11897 37791
rect 11931 37757 11943 37791
rect 11885 37751 11943 37757
rect 11977 37791 12035 37797
rect 11977 37757 11989 37791
rect 12023 37788 12035 37791
rect 12066 37788 12072 37800
rect 12023 37760 12072 37788
rect 12023 37757 12035 37760
rect 11977 37751 12035 37757
rect 8036 37692 8616 37720
rect 8676 37692 9076 37720
rect 8676 37652 8704 37692
rect 9306 37680 9312 37732
rect 9364 37720 9370 37732
rect 11992 37720 12020 37751
rect 12066 37748 12072 37760
rect 12124 37748 12130 37800
rect 9364 37692 12020 37720
rect 9364 37680 9370 37692
rect 7944 37624 8704 37652
rect 9033 37655 9091 37661
rect 9033 37621 9045 37655
rect 9079 37652 9091 37655
rect 9214 37652 9220 37664
rect 9079 37624 9220 37652
rect 9079 37621 9091 37624
rect 9033 37615 9091 37621
rect 9214 37612 9220 37624
rect 9272 37612 9278 37664
rect 10410 37612 10416 37664
rect 10468 37652 10474 37664
rect 12161 37655 12219 37661
rect 12161 37652 12173 37655
rect 10468 37624 12173 37652
rect 10468 37612 10474 37624
rect 12161 37621 12173 37624
rect 12207 37621 12219 37655
rect 12161 37615 12219 37621
rect 552 37562 12604 37584
rect 552 37510 4322 37562
rect 4374 37510 4386 37562
rect 4438 37510 4450 37562
rect 4502 37510 4514 37562
rect 4566 37510 4578 37562
rect 4630 37510 10722 37562
rect 10774 37510 10786 37562
rect 10838 37510 10850 37562
rect 10902 37510 10914 37562
rect 10966 37510 10978 37562
rect 11030 37510 12604 37562
rect 552 37488 12604 37510
rect 842 37408 848 37460
rect 900 37448 906 37460
rect 937 37451 995 37457
rect 937 37448 949 37451
rect 900 37420 949 37448
rect 900 37408 906 37420
rect 937 37417 949 37420
rect 983 37417 995 37451
rect 5813 37451 5871 37457
rect 5813 37448 5825 37451
rect 937 37411 995 37417
rect 1136 37420 5825 37448
rect 1026 37272 1032 37324
rect 1084 37272 1090 37324
rect 1136 37321 1164 37420
rect 5813 37417 5825 37420
rect 5859 37417 5871 37451
rect 5813 37411 5871 37417
rect 5902 37408 5908 37460
rect 5960 37448 5966 37460
rect 5960 37420 7144 37448
rect 5960 37408 5966 37420
rect 1486 37340 1492 37392
rect 1544 37380 1550 37392
rect 4249 37383 4307 37389
rect 4249 37380 4261 37383
rect 1544 37352 4261 37380
rect 1544 37340 1550 37352
rect 4249 37349 4261 37352
rect 4295 37349 4307 37383
rect 4249 37343 4307 37349
rect 4356 37352 5304 37380
rect 1121 37315 1179 37321
rect 1121 37281 1133 37315
rect 1167 37281 1179 37315
rect 1121 37275 1179 37281
rect 1210 37272 1216 37324
rect 1268 37272 1274 37324
rect 1394 37272 1400 37324
rect 1452 37272 1458 37324
rect 1578 37272 1584 37324
rect 1636 37312 1642 37324
rect 1673 37315 1731 37321
rect 1673 37312 1685 37315
rect 1636 37284 1685 37312
rect 1636 37272 1642 37284
rect 1673 37281 1685 37284
rect 1719 37281 1731 37315
rect 1673 37275 1731 37281
rect 1762 37272 1768 37324
rect 1820 37312 1826 37324
rect 1929 37315 1987 37321
rect 1929 37312 1941 37315
rect 1820 37284 1941 37312
rect 1820 37272 1826 37284
rect 1929 37281 1941 37284
rect 1975 37281 1987 37315
rect 1929 37275 1987 37281
rect 2222 37272 2228 37324
rect 2280 37312 2286 37324
rect 3513 37315 3571 37321
rect 3513 37312 3525 37315
rect 2280 37284 3525 37312
rect 2280 37272 2286 37284
rect 3513 37281 3525 37284
rect 3559 37281 3571 37315
rect 3513 37275 3571 37281
rect 3602 37272 3608 37324
rect 3660 37272 3666 37324
rect 3786 37272 3792 37324
rect 3844 37272 3850 37324
rect 4356 37312 4384 37352
rect 3896 37284 4384 37312
rect 4525 37315 4583 37321
rect 1581 37179 1639 37185
rect 1581 37145 1593 37179
rect 1627 37176 1639 37179
rect 1670 37176 1676 37188
rect 1627 37148 1676 37176
rect 1627 37145 1639 37148
rect 1581 37139 1639 37145
rect 1670 37136 1676 37148
rect 1728 37136 1734 37188
rect 2682 37136 2688 37188
rect 2740 37176 2746 37188
rect 3896 37176 3924 37284
rect 4525 37281 4537 37315
rect 4571 37281 4583 37315
rect 4525 37275 4583 37281
rect 4154 37204 4160 37256
rect 4212 37244 4218 37256
rect 4540 37244 4568 37275
rect 5074 37272 5080 37324
rect 5132 37272 5138 37324
rect 5276 37321 5304 37352
rect 6822 37340 6828 37392
rect 6880 37380 6886 37392
rect 6880 37352 7052 37380
rect 6880 37340 6886 37352
rect 5261 37315 5319 37321
rect 5261 37281 5273 37315
rect 5307 37281 5319 37315
rect 5261 37275 5319 37281
rect 5534 37272 5540 37324
rect 5592 37272 5598 37324
rect 6454 37272 6460 37324
rect 6512 37272 6518 37324
rect 6546 37272 6552 37324
rect 6604 37312 6610 37324
rect 6914 37312 6920 37324
rect 6604 37284 6920 37312
rect 6604 37272 6610 37284
rect 6914 37272 6920 37284
rect 6972 37272 6978 37324
rect 4212 37216 4568 37244
rect 4617 37247 4675 37253
rect 4212 37204 4218 37216
rect 4617 37213 4629 37247
rect 4663 37213 4675 37247
rect 4617 37207 4675 37213
rect 2740 37148 3924 37176
rect 2740 37136 2746 37148
rect 4430 37136 4436 37188
rect 4488 37176 4494 37188
rect 4632 37176 4660 37207
rect 4798 37204 4804 37256
rect 4856 37244 4862 37256
rect 7024 37253 7052 37352
rect 7116 37312 7144 37420
rect 7190 37408 7196 37460
rect 7248 37408 7254 37460
rect 7561 37451 7619 37457
rect 7561 37417 7573 37451
rect 7607 37448 7619 37451
rect 7834 37448 7840 37460
rect 7607 37420 7840 37448
rect 7607 37417 7619 37420
rect 7561 37411 7619 37417
rect 7834 37408 7840 37420
rect 7892 37408 7898 37460
rect 8846 37408 8852 37460
rect 8904 37408 8910 37460
rect 9582 37408 9588 37460
rect 9640 37448 9646 37460
rect 10321 37451 10379 37457
rect 10321 37448 10333 37451
rect 9640 37420 10333 37448
rect 9640 37408 9646 37420
rect 10321 37417 10333 37420
rect 10367 37448 10379 37451
rect 10870 37448 10876 37460
rect 10367 37420 10876 37448
rect 10367 37417 10379 37420
rect 10321 37411 10379 37417
rect 10870 37408 10876 37420
rect 10928 37408 10934 37460
rect 11146 37408 11152 37460
rect 11204 37448 11210 37460
rect 12161 37451 12219 37457
rect 12161 37448 12173 37451
rect 11204 37420 12173 37448
rect 11204 37408 11210 37420
rect 12161 37417 12173 37420
rect 12207 37417 12219 37451
rect 12161 37411 12219 37417
rect 7650 37340 7656 37392
rect 7708 37340 7714 37392
rect 9674 37380 9680 37392
rect 8588 37352 9680 37380
rect 8205 37315 8263 37321
rect 8205 37312 8217 37315
rect 7116 37284 8217 37312
rect 8205 37281 8217 37284
rect 8251 37281 8263 37315
rect 8205 37275 8263 37281
rect 4893 37247 4951 37253
rect 4893 37244 4905 37247
rect 4856 37216 4905 37244
rect 4856 37204 4862 37216
rect 4893 37213 4905 37216
rect 4939 37244 4951 37247
rect 5353 37247 5411 37253
rect 5353 37244 5365 37247
rect 4939 37216 5365 37244
rect 4939 37213 4951 37216
rect 4893 37207 4951 37213
rect 5353 37213 5365 37216
rect 5399 37213 5411 37247
rect 5353 37207 5411 37213
rect 7009 37247 7067 37253
rect 7009 37213 7021 37247
rect 7055 37213 7067 37247
rect 7009 37207 7067 37213
rect 7837 37247 7895 37253
rect 7837 37213 7849 37247
rect 7883 37244 7895 37247
rect 8110 37244 8116 37256
rect 7883 37216 8116 37244
rect 7883 37213 7895 37216
rect 7837 37207 7895 37213
rect 8110 37204 8116 37216
rect 8168 37204 8174 37256
rect 8220 37244 8248 37275
rect 8294 37272 8300 37324
rect 8352 37272 8358 37324
rect 8588 37312 8616 37352
rect 9674 37340 9680 37352
rect 9732 37340 9738 37392
rect 11238 37340 11244 37392
rect 11296 37340 11302 37392
rect 11425 37383 11483 37389
rect 11425 37349 11437 37383
rect 11471 37380 11483 37383
rect 11790 37380 11796 37392
rect 11471 37352 11796 37380
rect 11471 37349 11483 37352
rect 11425 37343 11483 37349
rect 11790 37340 11796 37352
rect 11848 37380 11854 37392
rect 11885 37383 11943 37389
rect 11885 37380 11897 37383
rect 11848 37352 11897 37380
rect 11848 37340 11854 37352
rect 11885 37349 11897 37352
rect 11931 37349 11943 37383
rect 11885 37343 11943 37349
rect 8496 37284 8616 37312
rect 8665 37315 8723 37321
rect 8496 37244 8524 37284
rect 8665 37281 8677 37315
rect 8711 37281 8723 37315
rect 8665 37275 8723 37281
rect 8220 37216 8524 37244
rect 8680 37244 8708 37275
rect 8754 37272 8760 37324
rect 8812 37272 8818 37324
rect 8846 37272 8852 37324
rect 8904 37312 8910 37324
rect 8941 37315 8999 37321
rect 8941 37312 8953 37315
rect 8904 37284 8953 37312
rect 8904 37272 8910 37284
rect 8941 37281 8953 37284
rect 8987 37281 8999 37315
rect 8941 37275 8999 37281
rect 9033 37315 9091 37321
rect 9033 37281 9045 37315
rect 9079 37312 9091 37315
rect 9582 37312 9588 37324
rect 9079 37284 9588 37312
rect 9079 37281 9091 37284
rect 9033 37275 9091 37281
rect 9582 37272 9588 37284
rect 9640 37272 9646 37324
rect 10318 37272 10324 37324
rect 10376 37272 10382 37324
rect 11149 37315 11207 37321
rect 11149 37281 11161 37315
rect 11195 37312 11207 37315
rect 11256 37312 11284 37340
rect 11195 37284 11284 37312
rect 11517 37315 11575 37321
rect 11195 37281 11207 37284
rect 11149 37275 11207 37281
rect 11517 37281 11529 37315
rect 11563 37281 11575 37315
rect 11517 37275 11575 37281
rect 8864 37244 8892 37272
rect 8680 37216 8892 37244
rect 10336 37244 10364 37272
rect 10336 37216 11008 37244
rect 4488 37148 4660 37176
rect 5445 37179 5503 37185
rect 4488 37136 4494 37148
rect 5445 37145 5457 37179
rect 5491 37145 5503 37179
rect 5445 37139 5503 37145
rect 3050 37068 3056 37120
rect 3108 37068 3114 37120
rect 3326 37068 3332 37120
rect 3384 37108 3390 37120
rect 5460 37108 5488 37139
rect 5534 37136 5540 37188
rect 5592 37176 5598 37188
rect 6549 37179 6607 37185
rect 6549 37176 6561 37179
rect 5592 37148 6561 37176
rect 5592 37136 5598 37148
rect 6549 37145 6561 37148
rect 6595 37145 6607 37179
rect 6549 37139 6607 37145
rect 7282 37136 7288 37188
rect 7340 37176 7346 37188
rect 7650 37176 7656 37188
rect 7340 37148 7656 37176
rect 7340 37136 7346 37148
rect 7650 37136 7656 37148
rect 7708 37176 7714 37188
rect 7708 37148 8248 37176
rect 7708 37136 7714 37148
rect 3384 37080 5488 37108
rect 3384 37068 3390 37080
rect 8018 37068 8024 37120
rect 8076 37068 8082 37120
rect 8220 37117 8248 37148
rect 8386 37136 8392 37188
rect 8444 37176 8450 37188
rect 9030 37176 9036 37188
rect 8444 37148 9036 37176
rect 8444 37136 8450 37148
rect 9030 37136 9036 37148
rect 9088 37136 9094 37188
rect 10980 37176 11008 37216
rect 11238 37204 11244 37256
rect 11296 37204 11302 37256
rect 11422 37204 11428 37256
rect 11480 37244 11486 37256
rect 11532 37244 11560 37275
rect 11698 37272 11704 37324
rect 11756 37272 11762 37324
rect 11974 37272 11980 37324
rect 12032 37272 12038 37324
rect 12526 37244 12532 37256
rect 11480 37216 12532 37244
rect 11480 37204 11486 37216
rect 12526 37204 12532 37216
rect 12584 37204 12590 37256
rect 11698 37176 11704 37188
rect 10980 37148 11704 37176
rect 11698 37136 11704 37148
rect 11756 37136 11762 37188
rect 8205 37111 8263 37117
rect 8205 37077 8217 37111
rect 8251 37077 8263 37111
rect 8205 37071 8263 37077
rect 8570 37068 8576 37120
rect 8628 37108 8634 37120
rect 9122 37108 9128 37120
rect 8628 37080 9128 37108
rect 8628 37068 8634 37080
rect 9122 37068 9128 37080
rect 9180 37108 9186 37120
rect 9398 37108 9404 37120
rect 9180 37080 9404 37108
rect 9180 37068 9186 37080
rect 9398 37068 9404 37080
rect 9456 37068 9462 37120
rect 9766 37068 9772 37120
rect 9824 37108 9830 37120
rect 10965 37111 11023 37117
rect 10965 37108 10977 37111
rect 9824 37080 10977 37108
rect 9824 37068 9830 37080
rect 10965 37077 10977 37080
rect 11011 37077 11023 37111
rect 10965 37071 11023 37077
rect 11146 37068 11152 37120
rect 11204 37108 11210 37120
rect 12710 37108 12716 37120
rect 11204 37080 12716 37108
rect 11204 37068 11210 37080
rect 12710 37068 12716 37080
rect 12768 37068 12774 37120
rect 552 37018 12604 37040
rect 552 36966 3662 37018
rect 3714 36966 3726 37018
rect 3778 36966 3790 37018
rect 3842 36966 3854 37018
rect 3906 36966 3918 37018
rect 3970 36966 10062 37018
rect 10114 36966 10126 37018
rect 10178 36966 10190 37018
rect 10242 36966 10254 37018
rect 10306 36966 10318 37018
rect 10370 36966 12604 37018
rect 552 36944 12604 36966
rect 1394 36864 1400 36916
rect 1452 36904 1458 36916
rect 3142 36904 3148 36916
rect 1452 36876 3148 36904
rect 1452 36864 1458 36876
rect 3142 36864 3148 36876
rect 3200 36864 3206 36916
rect 3234 36864 3240 36916
rect 3292 36864 3298 36916
rect 3878 36864 3884 36916
rect 3936 36904 3942 36916
rect 7285 36907 7343 36913
rect 7285 36904 7297 36907
rect 3936 36876 7297 36904
rect 3936 36864 3942 36876
rect 3050 36796 3056 36848
rect 3108 36836 3114 36848
rect 3510 36836 3516 36848
rect 3108 36808 3516 36836
rect 3108 36796 3114 36808
rect 3510 36796 3516 36808
rect 3568 36796 3574 36848
rect 1397 36771 1455 36777
rect 1397 36737 1409 36771
rect 1443 36768 1455 36771
rect 1578 36768 1584 36780
rect 1443 36740 1584 36768
rect 1443 36737 1455 36740
rect 1397 36731 1455 36737
rect 1578 36728 1584 36740
rect 1636 36728 1642 36780
rect 2774 36728 2780 36780
rect 2832 36768 2838 36780
rect 3142 36768 3148 36780
rect 2832 36740 3148 36768
rect 2832 36728 2838 36740
rect 3142 36728 3148 36740
rect 3200 36728 3206 36780
rect 198 36660 204 36712
rect 256 36700 262 36712
rect 1118 36700 1124 36712
rect 256 36672 1124 36700
rect 256 36660 262 36672
rect 1118 36660 1124 36672
rect 1176 36700 1182 36712
rect 1305 36703 1363 36709
rect 1305 36700 1317 36703
rect 1176 36672 1317 36700
rect 1176 36660 1182 36672
rect 1305 36669 1317 36672
rect 1351 36669 1363 36703
rect 1305 36663 1363 36669
rect 1673 36703 1731 36709
rect 1673 36669 1685 36703
rect 1719 36700 1731 36703
rect 1762 36700 1768 36712
rect 1719 36672 1768 36700
rect 1719 36669 1731 36672
rect 1673 36663 1731 36669
rect 1762 36660 1768 36672
rect 1820 36660 1826 36712
rect 4724 36709 4752 36876
rect 7285 36873 7297 36876
rect 7331 36873 7343 36907
rect 7285 36867 7343 36873
rect 7650 36864 7656 36916
rect 7708 36904 7714 36916
rect 8205 36907 8263 36913
rect 8205 36904 8217 36907
rect 7708 36876 8217 36904
rect 7708 36864 7714 36876
rect 8205 36873 8217 36876
rect 8251 36904 8263 36907
rect 8294 36904 8300 36916
rect 8251 36876 8300 36904
rect 8251 36873 8263 36876
rect 8205 36867 8263 36873
rect 8294 36864 8300 36876
rect 8352 36864 8358 36916
rect 8570 36864 8576 36916
rect 8628 36864 8634 36916
rect 8662 36864 8668 36916
rect 8720 36864 8726 36916
rect 8754 36864 8760 36916
rect 8812 36864 8818 36916
rect 9214 36864 9220 36916
rect 9272 36904 9278 36916
rect 9272 36876 9536 36904
rect 9272 36864 9278 36876
rect 4890 36796 4896 36848
rect 4948 36836 4954 36848
rect 6730 36836 6736 36848
rect 4948 36808 6736 36836
rect 4948 36796 4954 36808
rect 6730 36796 6736 36808
rect 6788 36796 6794 36848
rect 6917 36839 6975 36845
rect 6917 36805 6929 36839
rect 6963 36836 6975 36839
rect 7098 36836 7104 36848
rect 6963 36808 7104 36836
rect 6963 36805 6975 36808
rect 6917 36799 6975 36805
rect 7098 36796 7104 36808
rect 7156 36796 7162 36848
rect 7745 36839 7803 36845
rect 7745 36805 7757 36839
rect 7791 36836 7803 36839
rect 8386 36836 8392 36848
rect 7791 36808 8392 36836
rect 7791 36805 7803 36808
rect 7745 36799 7803 36805
rect 8386 36796 8392 36808
rect 8444 36796 8450 36848
rect 8588 36836 8616 36864
rect 8496 36808 8616 36836
rect 5442 36728 5448 36780
rect 5500 36768 5506 36780
rect 5997 36771 6055 36777
rect 5997 36768 6009 36771
rect 5500 36740 6009 36768
rect 5500 36728 5506 36740
rect 5997 36737 6009 36740
rect 6043 36737 6055 36771
rect 5997 36731 6055 36737
rect 6086 36728 6092 36780
rect 6144 36768 6150 36780
rect 6546 36768 6552 36780
rect 6144 36740 6552 36768
rect 6144 36728 6150 36740
rect 6546 36728 6552 36740
rect 6604 36768 6610 36780
rect 7193 36771 7251 36777
rect 7193 36768 7205 36771
rect 6604 36740 7205 36768
rect 6604 36728 6610 36740
rect 7193 36737 7205 36740
rect 7239 36737 7251 36771
rect 8113 36771 8171 36777
rect 7193 36731 7251 36737
rect 7760 36740 8064 36768
rect 7760 36712 7788 36740
rect 4617 36703 4675 36709
rect 4617 36700 4629 36703
rect 4264 36672 4629 36700
rect 4264 36644 4292 36672
rect 4617 36669 4629 36672
rect 4663 36669 4675 36703
rect 4617 36663 4675 36669
rect 4709 36703 4767 36709
rect 4709 36669 4721 36703
rect 4755 36669 4767 36703
rect 4709 36663 4767 36669
rect 4982 36660 4988 36712
rect 5040 36700 5046 36712
rect 5353 36703 5411 36709
rect 5353 36700 5365 36703
rect 5040 36672 5365 36700
rect 5040 36660 5046 36672
rect 5353 36669 5365 36672
rect 5399 36669 5411 36703
rect 5353 36663 5411 36669
rect 5721 36703 5779 36709
rect 5721 36669 5733 36703
rect 5767 36669 5779 36703
rect 5721 36663 5779 36669
rect 5905 36703 5963 36709
rect 5905 36669 5917 36703
rect 5951 36700 5963 36703
rect 7006 36700 7012 36712
rect 5951 36672 7012 36700
rect 5951 36669 5963 36672
rect 5905 36663 5963 36669
rect 3050 36592 3056 36644
rect 3108 36592 3114 36644
rect 4246 36592 4252 36644
rect 4304 36592 4310 36644
rect 4338 36592 4344 36644
rect 4396 36641 4402 36644
rect 4396 36635 4430 36641
rect 4418 36632 4430 36635
rect 4418 36604 4752 36632
rect 4418 36601 4430 36604
rect 4396 36595 4430 36601
rect 4396 36592 4402 36595
rect 4724 36576 4752 36604
rect 5074 36592 5080 36644
rect 5132 36632 5138 36644
rect 5169 36635 5227 36641
rect 5169 36632 5181 36635
rect 5132 36604 5181 36632
rect 5132 36592 5138 36604
rect 5169 36601 5181 36604
rect 5215 36632 5227 36635
rect 5626 36632 5632 36644
rect 5215 36604 5632 36632
rect 5215 36601 5227 36604
rect 5169 36595 5227 36601
rect 5626 36592 5632 36604
rect 5684 36592 5690 36644
rect 5736 36632 5764 36663
rect 7006 36660 7012 36672
rect 7064 36660 7070 36712
rect 7282 36660 7288 36712
rect 7340 36660 7346 36712
rect 7466 36660 7472 36712
rect 7524 36660 7530 36712
rect 7742 36660 7748 36712
rect 7800 36660 7806 36712
rect 7834 36660 7840 36712
rect 7892 36702 7898 36712
rect 7929 36703 7987 36709
rect 7929 36702 7941 36703
rect 7892 36674 7941 36702
rect 7892 36660 7898 36674
rect 7929 36669 7941 36674
rect 7975 36669 7987 36703
rect 8036 36700 8064 36740
rect 8113 36737 8125 36771
rect 8159 36768 8171 36771
rect 8159 36740 8432 36768
rect 8159 36737 8171 36740
rect 8113 36731 8171 36737
rect 8205 36703 8263 36709
rect 8205 36700 8217 36703
rect 8036 36672 8217 36700
rect 7929 36663 7987 36669
rect 8205 36669 8217 36672
rect 8251 36669 8263 36703
rect 8404 36687 8432 36740
rect 8496 36709 8524 36808
rect 8676 36768 8704 36864
rect 8938 36836 8944 36848
rect 8869 36808 8944 36836
rect 8754 36768 8760 36780
rect 8676 36740 8760 36768
rect 8754 36728 8760 36740
rect 8812 36728 8818 36780
rect 8481 36703 8539 36709
rect 8205 36663 8263 36669
rect 8380 36681 8438 36687
rect 8380 36647 8392 36681
rect 8426 36647 8438 36681
rect 8481 36669 8493 36703
rect 8527 36669 8539 36703
rect 8481 36663 8539 36669
rect 8380 36644 8438 36647
rect 7098 36632 7104 36644
rect 5736 36604 7104 36632
rect 7098 36592 7104 36604
rect 7156 36592 7162 36644
rect 8380 36641 8392 36644
rect 8386 36592 8392 36641
rect 8444 36592 8450 36644
rect 382 36524 388 36576
rect 440 36564 446 36576
rect 1121 36567 1179 36573
rect 1121 36564 1133 36567
rect 440 36536 1133 36564
rect 440 36524 446 36536
rect 1121 36533 1133 36536
rect 1167 36533 1179 36567
rect 1121 36527 1179 36533
rect 3786 36524 3792 36576
rect 3844 36564 3850 36576
rect 4522 36564 4528 36576
rect 3844 36536 4528 36564
rect 3844 36524 3850 36536
rect 4522 36524 4528 36536
rect 4580 36524 4586 36576
rect 4706 36524 4712 36576
rect 4764 36524 4770 36576
rect 5902 36524 5908 36576
rect 5960 36524 5966 36576
rect 6270 36524 6276 36576
rect 6328 36564 6334 36576
rect 6641 36567 6699 36573
rect 6641 36564 6653 36567
rect 6328 36536 6653 36564
rect 6328 36524 6334 36536
rect 6641 36533 6653 36536
rect 6687 36533 6699 36567
rect 6641 36527 6699 36533
rect 6730 36524 6736 36576
rect 6788 36564 6794 36576
rect 7282 36564 7288 36576
rect 6788 36536 7288 36564
rect 6788 36524 6794 36536
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 7650 36524 7656 36576
rect 7708 36524 7714 36576
rect 7742 36524 7748 36576
rect 7800 36564 7806 36576
rect 8496 36564 8524 36663
rect 8658 36626 8664 36678
rect 8716 36641 8722 36678
rect 8716 36626 8723 36641
rect 8665 36601 8677 36626
rect 8711 36601 8723 36626
rect 8665 36595 8723 36601
rect 7800 36536 8524 36564
rect 8566 36567 8624 36573
rect 7800 36524 7806 36536
rect 8566 36533 8578 36567
rect 8612 36564 8624 36567
rect 8869 36564 8897 36808
rect 8938 36796 8944 36808
rect 8996 36796 9002 36848
rect 9122 36796 9128 36848
rect 9180 36836 9186 36848
rect 9401 36839 9459 36845
rect 9401 36836 9413 36839
rect 9180 36808 9413 36836
rect 9180 36796 9186 36808
rect 9401 36805 9413 36808
rect 9447 36805 9459 36839
rect 9401 36799 9459 36805
rect 9030 36728 9036 36780
rect 9088 36728 9094 36780
rect 9217 36771 9275 36777
rect 9217 36737 9229 36771
rect 9263 36768 9275 36771
rect 9508 36768 9536 36876
rect 11238 36864 11244 36916
rect 11296 36904 11302 36916
rect 11790 36904 11796 36916
rect 11296 36876 11796 36904
rect 11296 36864 11302 36876
rect 11790 36864 11796 36876
rect 11848 36864 11854 36916
rect 9674 36796 9680 36848
rect 9732 36796 9738 36848
rect 9263 36740 9536 36768
rect 9692 36768 9720 36796
rect 10318 36768 10324 36780
rect 9692 36740 10324 36768
rect 9263 36737 9275 36740
rect 9217 36731 9275 36737
rect 10318 36728 10324 36740
rect 10376 36728 10382 36780
rect 10594 36728 10600 36780
rect 10652 36768 10658 36780
rect 10870 36768 10876 36780
rect 10652 36740 10876 36768
rect 10652 36728 10658 36740
rect 10870 36728 10876 36740
rect 10928 36728 10934 36780
rect 8937 36703 8995 36709
rect 8937 36669 8949 36703
rect 8983 36700 8995 36703
rect 9125 36703 9183 36709
rect 8983 36672 9076 36700
rect 8983 36669 8995 36672
rect 8937 36663 8995 36669
rect 9048 36644 9076 36672
rect 9125 36669 9137 36703
rect 9171 36669 9183 36703
rect 9125 36663 9183 36669
rect 9030 36592 9036 36644
rect 9088 36592 9094 36644
rect 8612 36536 8897 36564
rect 9140 36564 9168 36663
rect 9398 36660 9404 36712
rect 9456 36660 9462 36712
rect 9677 36703 9735 36709
rect 9677 36669 9689 36703
rect 9723 36700 9735 36703
rect 10229 36703 10287 36709
rect 9723 36672 9996 36700
rect 9723 36669 9735 36672
rect 9677 36663 9735 36669
rect 9416 36632 9444 36660
rect 9968 36632 9996 36672
rect 10229 36669 10241 36703
rect 10275 36700 10287 36703
rect 10410 36700 10416 36712
rect 10275 36672 10416 36700
rect 10275 36669 10287 36672
rect 10229 36663 10287 36669
rect 10410 36660 10416 36672
rect 10468 36660 10474 36712
rect 10781 36703 10839 36709
rect 10781 36669 10793 36703
rect 10827 36700 10839 36703
rect 11974 36700 11980 36712
rect 10827 36672 11980 36700
rect 10827 36669 10839 36672
rect 10781 36663 10839 36669
rect 11974 36660 11980 36672
rect 12032 36660 12038 36712
rect 11146 36641 11152 36644
rect 9416 36604 9904 36632
rect 9968 36604 10815 36632
rect 9876 36576 9904 36604
rect 9398 36564 9404 36576
rect 9140 36536 9404 36564
rect 8612 36533 8624 36536
rect 8566 36527 8624 36533
rect 9398 36524 9404 36536
rect 9456 36524 9462 36576
rect 9490 36524 9496 36576
rect 9548 36564 9554 36576
rect 9585 36567 9643 36573
rect 9585 36564 9597 36567
rect 9548 36536 9597 36564
rect 9548 36524 9554 36536
rect 9585 36533 9597 36536
rect 9631 36533 9643 36567
rect 9585 36527 9643 36533
rect 9766 36524 9772 36576
rect 9824 36524 9830 36576
rect 9858 36524 9864 36576
rect 9916 36524 9922 36576
rect 9950 36524 9956 36576
rect 10008 36564 10014 36576
rect 10137 36567 10195 36573
rect 10137 36564 10149 36567
rect 10008 36536 10149 36564
rect 10008 36524 10014 36536
rect 10137 36533 10149 36536
rect 10183 36533 10195 36567
rect 10137 36527 10195 36533
rect 10410 36524 10416 36576
rect 10468 36564 10474 36576
rect 10689 36567 10747 36573
rect 10689 36564 10701 36567
rect 10468 36536 10701 36564
rect 10468 36524 10474 36536
rect 10689 36533 10701 36536
rect 10735 36533 10747 36567
rect 10787 36564 10815 36604
rect 11140 36595 11152 36641
rect 11146 36592 11152 36595
rect 11204 36592 11210 36644
rect 11238 36564 11244 36576
rect 10787 36536 11244 36564
rect 10689 36527 10747 36533
rect 11238 36524 11244 36536
rect 11296 36524 11302 36576
rect 12066 36524 12072 36576
rect 12124 36564 12130 36576
rect 12253 36567 12311 36573
rect 12253 36564 12265 36567
rect 12124 36536 12265 36564
rect 12124 36524 12130 36536
rect 12253 36533 12265 36536
rect 12299 36533 12311 36567
rect 12253 36527 12311 36533
rect 552 36474 12604 36496
rect 552 36422 4322 36474
rect 4374 36422 4386 36474
rect 4438 36422 4450 36474
rect 4502 36422 4514 36474
rect 4566 36422 4578 36474
rect 4630 36422 10722 36474
rect 10774 36422 10786 36474
rect 10838 36422 10850 36474
rect 10902 36422 10914 36474
rect 10966 36422 10978 36474
rect 11030 36422 12604 36474
rect 552 36400 12604 36422
rect 3510 36320 3516 36372
rect 3568 36360 3574 36372
rect 4798 36360 4804 36372
rect 3568 36332 4804 36360
rect 3568 36320 3574 36332
rect 4798 36320 4804 36332
rect 4856 36320 4862 36372
rect 5813 36363 5871 36369
rect 5813 36329 5825 36363
rect 5859 36329 5871 36363
rect 5813 36323 5871 36329
rect 4516 36295 4574 36301
rect 4516 36261 4528 36295
rect 4562 36292 4574 36295
rect 5828 36292 5856 36323
rect 6270 36320 6276 36372
rect 6328 36320 6334 36372
rect 6638 36320 6644 36372
rect 6696 36360 6702 36372
rect 7561 36363 7619 36369
rect 7561 36360 7573 36363
rect 6696 36332 7573 36360
rect 6696 36320 6702 36332
rect 7561 36329 7573 36332
rect 7607 36329 7619 36363
rect 7561 36323 7619 36329
rect 8573 36363 8631 36369
rect 8573 36329 8585 36363
rect 8619 36360 8631 36363
rect 10318 36360 10324 36372
rect 8619 36329 8635 36360
rect 8573 36323 8635 36329
rect 4562 36264 5856 36292
rect 4562 36261 4574 36264
rect 4516 36255 4574 36261
rect 5902 36252 5908 36304
rect 5960 36292 5966 36304
rect 6730 36292 6736 36304
rect 5960 36264 6736 36292
rect 5960 36252 5966 36264
rect 6730 36252 6736 36264
rect 6788 36292 6794 36304
rect 6788 36264 6960 36292
rect 6788 36252 6794 36264
rect 106 36184 112 36236
rect 164 36224 170 36236
rect 290 36224 296 36236
rect 164 36196 296 36224
rect 164 36184 170 36196
rect 290 36184 296 36196
rect 348 36224 354 36236
rect 1026 36224 1032 36236
rect 348 36196 1032 36224
rect 348 36184 354 36196
rect 1026 36184 1032 36196
rect 1084 36224 1090 36236
rect 1121 36227 1179 36233
rect 1121 36224 1133 36227
rect 1084 36196 1133 36224
rect 1084 36184 1090 36196
rect 1121 36193 1133 36196
rect 1167 36193 1179 36227
rect 1121 36187 1179 36193
rect 1305 36227 1363 36233
rect 1305 36193 1317 36227
rect 1351 36224 1363 36227
rect 1486 36224 1492 36236
rect 1351 36196 1492 36224
rect 1351 36193 1363 36196
rect 1305 36187 1363 36193
rect 1486 36184 1492 36196
rect 1544 36184 1550 36236
rect 1578 36184 1584 36236
rect 1636 36184 1642 36236
rect 3510 36184 3516 36236
rect 3568 36224 3574 36236
rect 3789 36227 3847 36233
rect 3789 36224 3801 36227
rect 3568 36196 3801 36224
rect 3568 36184 3574 36196
rect 3789 36193 3801 36196
rect 3835 36224 3847 36227
rect 4154 36224 4160 36236
rect 3835 36196 4160 36224
rect 3835 36193 3847 36196
rect 3789 36187 3847 36193
rect 4154 36184 4160 36196
rect 4212 36184 4218 36236
rect 4246 36184 4252 36236
rect 4304 36184 4310 36236
rect 4338 36184 4344 36236
rect 4396 36224 4402 36236
rect 5626 36224 5632 36236
rect 4396 36196 5632 36224
rect 4396 36184 4402 36196
rect 5626 36184 5632 36196
rect 5684 36184 5690 36236
rect 6181 36227 6239 36233
rect 6181 36193 6193 36227
rect 6227 36224 6239 36227
rect 6546 36224 6552 36236
rect 6227 36196 6552 36224
rect 6227 36193 6239 36196
rect 6181 36187 6239 36193
rect 6546 36184 6552 36196
rect 6604 36184 6610 36236
rect 6638 36184 6644 36236
rect 6696 36184 6702 36236
rect 6932 36233 6960 36264
rect 7006 36252 7012 36304
rect 7064 36292 7070 36304
rect 7469 36295 7527 36301
rect 7469 36292 7481 36295
rect 7064 36264 7481 36292
rect 7064 36252 7070 36264
rect 7469 36261 7481 36264
rect 7515 36261 7527 36295
rect 7469 36255 7527 36261
rect 8018 36252 8024 36304
rect 8076 36292 8082 36304
rect 8113 36295 8171 36301
rect 8113 36292 8125 36295
rect 8076 36264 8125 36292
rect 8076 36252 8082 36264
rect 8113 36261 8125 36264
rect 8159 36261 8171 36295
rect 8113 36255 8171 36261
rect 8202 36252 8208 36304
rect 8260 36292 8266 36304
rect 8607 36292 8635 36323
rect 9140 36332 10324 36360
rect 8754 36292 8760 36304
rect 8260 36264 8524 36292
rect 8607 36264 8760 36292
rect 8260 36252 8266 36264
rect 6825 36227 6883 36233
rect 6825 36193 6837 36227
rect 6871 36193 6883 36227
rect 6825 36187 6883 36193
rect 6917 36227 6975 36233
rect 6917 36193 6929 36227
rect 6963 36193 6975 36227
rect 6917 36187 6975 36193
rect 7101 36227 7159 36233
rect 7101 36193 7113 36227
rect 7147 36224 7159 36227
rect 7374 36224 7380 36236
rect 7147 36196 7380 36224
rect 7147 36193 7159 36196
rect 7101 36187 7159 36193
rect 750 36116 756 36168
rect 808 36156 814 36168
rect 3970 36156 3976 36168
rect 808 36128 3976 36156
rect 808 36116 814 36128
rect 3970 36116 3976 36128
rect 4028 36116 4034 36168
rect 6362 36116 6368 36168
rect 6420 36116 6426 36168
rect 6454 36116 6460 36168
rect 6512 36156 6518 36168
rect 6656 36156 6684 36184
rect 6512 36128 6684 36156
rect 6512 36116 6518 36128
rect 1489 36091 1547 36097
rect 1489 36057 1501 36091
rect 1535 36088 1547 36091
rect 1946 36088 1952 36100
rect 1535 36060 1952 36088
rect 1535 36057 1547 36060
rect 1489 36051 1547 36057
rect 1946 36048 1952 36060
rect 2004 36048 2010 36100
rect 3786 36048 3792 36100
rect 3844 36088 3850 36100
rect 4154 36088 4160 36100
rect 3844 36060 4160 36088
rect 3844 36048 3850 36060
rect 4154 36048 4160 36060
rect 4212 36048 4218 36100
rect 5810 36048 5816 36100
rect 5868 36088 5874 36100
rect 6840 36088 6868 36187
rect 7374 36184 7380 36196
rect 7432 36184 7438 36236
rect 7745 36227 7803 36233
rect 7745 36193 7757 36227
rect 7791 36193 7803 36227
rect 7745 36187 7803 36193
rect 7006 36116 7012 36168
rect 7064 36156 7070 36168
rect 7760 36156 7788 36187
rect 7834 36184 7840 36236
rect 7892 36224 7898 36236
rect 8389 36227 8447 36233
rect 8389 36224 8401 36227
rect 7892 36196 8401 36224
rect 7892 36184 7898 36196
rect 8389 36193 8401 36196
rect 8435 36193 8447 36227
rect 8389 36187 8447 36193
rect 7064 36128 7788 36156
rect 7064 36116 7070 36128
rect 7926 36116 7932 36168
rect 7984 36156 7990 36168
rect 8021 36159 8079 36165
rect 8021 36156 8033 36159
rect 7984 36128 8033 36156
rect 7984 36116 7990 36128
rect 8021 36125 8033 36128
rect 8067 36125 8079 36159
rect 8297 36159 8355 36165
rect 8297 36156 8309 36159
rect 8021 36119 8079 36125
rect 8220 36128 8309 36156
rect 8220 36100 8248 36128
rect 8297 36125 8309 36128
rect 8343 36125 8355 36159
rect 8297 36119 8355 36125
rect 5868 36060 6868 36088
rect 7285 36091 7343 36097
rect 5868 36048 5874 36060
rect 6472 36032 6500 36060
rect 7285 36057 7297 36091
rect 7331 36088 7343 36091
rect 7834 36088 7840 36100
rect 7331 36060 7840 36088
rect 7331 36057 7343 36060
rect 7285 36051 7343 36057
rect 7834 36048 7840 36060
rect 7892 36048 7898 36100
rect 8202 36048 8208 36100
rect 8260 36048 8266 36100
rect 8496 36088 8524 36264
rect 8754 36252 8760 36264
rect 8812 36252 8818 36304
rect 8938 36252 8944 36304
rect 8996 36252 9002 36304
rect 9140 36301 9168 36332
rect 10318 36320 10324 36332
rect 10376 36320 10382 36372
rect 10410 36320 10416 36372
rect 10468 36360 10474 36372
rect 10686 36360 10692 36372
rect 10468 36332 10692 36360
rect 10468 36320 10474 36332
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 10965 36363 11023 36369
rect 10965 36329 10977 36363
rect 11011 36360 11023 36363
rect 11146 36360 11152 36372
rect 11011 36332 11152 36360
rect 11011 36329 11023 36332
rect 10965 36323 11023 36329
rect 11146 36320 11152 36332
rect 11204 36320 11210 36372
rect 11701 36363 11759 36369
rect 11701 36329 11713 36363
rect 11747 36360 11759 36363
rect 12158 36360 12164 36372
rect 11747 36332 12164 36360
rect 11747 36329 11759 36332
rect 11701 36323 11759 36329
rect 12158 36320 12164 36332
rect 12216 36320 12222 36372
rect 9125 36295 9183 36301
rect 9125 36261 9137 36295
rect 9171 36261 9183 36295
rect 10226 36292 10232 36304
rect 9125 36255 9183 36261
rect 9784 36264 10232 36292
rect 8849 36227 8907 36233
rect 8849 36193 8861 36227
rect 8895 36224 8907 36227
rect 8956 36224 8984 36252
rect 9398 36224 9404 36236
rect 8895 36196 9404 36224
rect 8895 36193 8907 36196
rect 8849 36187 8907 36193
rect 9398 36184 9404 36196
rect 9456 36224 9462 36236
rect 9784 36233 9812 36264
rect 10226 36252 10232 36264
rect 10284 36252 10290 36304
rect 10428 36264 11652 36292
rect 10428 36236 10456 36264
rect 9769 36227 9827 36233
rect 9769 36224 9781 36227
rect 9456 36196 9781 36224
rect 9456 36184 9462 36196
rect 9769 36193 9781 36196
rect 9815 36193 9827 36227
rect 9769 36187 9827 36193
rect 9861 36227 9919 36233
rect 9861 36193 9873 36227
rect 9907 36224 9919 36227
rect 10134 36224 10140 36236
rect 9907 36196 10140 36224
rect 9907 36193 9919 36196
rect 9861 36187 9919 36193
rect 10134 36184 10140 36196
rect 10192 36184 10198 36236
rect 10410 36184 10416 36236
rect 10468 36184 10474 36236
rect 11149 36227 11207 36233
rect 11149 36224 11161 36227
rect 10796 36196 11161 36224
rect 8570 36116 8576 36168
rect 8628 36156 8634 36168
rect 9033 36159 9091 36165
rect 9033 36156 9045 36159
rect 8628 36128 9045 36156
rect 8628 36116 8634 36128
rect 9033 36125 9045 36128
rect 9079 36125 9091 36159
rect 9033 36119 9091 36125
rect 8665 36091 8723 36097
rect 8665 36088 8677 36091
rect 8496 36060 8677 36088
rect 8665 36057 8677 36060
rect 8711 36057 8723 36091
rect 9048 36088 9076 36119
rect 9306 36116 9312 36168
rect 9364 36156 9370 36168
rect 9577 36159 9635 36165
rect 9577 36156 9589 36159
rect 9364 36128 9589 36156
rect 9364 36116 9370 36128
rect 9577 36125 9589 36128
rect 9623 36125 9635 36159
rect 9577 36119 9635 36125
rect 9674 36116 9680 36168
rect 9732 36116 9738 36168
rect 10042 36116 10048 36168
rect 10100 36156 10106 36168
rect 10796 36165 10824 36196
rect 11149 36193 11161 36196
rect 11195 36193 11207 36227
rect 11149 36187 11207 36193
rect 11241 36227 11299 36233
rect 11241 36193 11253 36227
rect 11287 36193 11299 36227
rect 11241 36187 11299 36193
rect 11333 36227 11391 36233
rect 11333 36193 11345 36227
rect 11379 36193 11391 36227
rect 11451 36227 11509 36233
rect 11451 36224 11463 36227
rect 11333 36187 11391 36193
rect 11440 36193 11463 36224
rect 11497 36193 11509 36227
rect 11440 36187 11509 36193
rect 10321 36159 10379 36165
rect 10321 36156 10333 36159
rect 10100 36128 10333 36156
rect 10100 36116 10106 36128
rect 10321 36125 10333 36128
rect 10367 36125 10379 36159
rect 10321 36119 10379 36125
rect 10781 36159 10839 36165
rect 10781 36125 10793 36159
rect 10827 36125 10839 36159
rect 10781 36119 10839 36125
rect 10134 36088 10140 36100
rect 9048 36060 10140 36088
rect 8665 36051 8723 36057
rect 10134 36048 10140 36060
rect 10192 36048 10198 36100
rect 10336 36088 10364 36119
rect 10962 36116 10968 36168
rect 11020 36156 11026 36168
rect 11256 36156 11284 36187
rect 11020 36128 11284 36156
rect 11020 36116 11026 36128
rect 11146 36088 11152 36100
rect 10336 36060 11152 36088
rect 11146 36048 11152 36060
rect 11204 36048 11210 36100
rect 934 35980 940 36032
rect 992 35980 998 36032
rect 3418 35980 3424 36032
rect 3476 36020 3482 36032
rect 3878 36020 3884 36032
rect 3476 35992 3884 36020
rect 3476 35980 3482 35992
rect 3878 35980 3884 35992
rect 3936 36020 3942 36032
rect 3973 36023 4031 36029
rect 3973 36020 3985 36023
rect 3936 35992 3985 36020
rect 3936 35980 3942 35992
rect 3973 35989 3985 35992
rect 4019 35989 4031 36023
rect 3973 35983 4031 35989
rect 5442 35980 5448 36032
rect 5500 36020 5506 36032
rect 5629 36023 5687 36029
rect 5629 36020 5641 36023
rect 5500 35992 5641 36020
rect 5500 35980 5506 35992
rect 5629 35989 5641 35992
rect 5675 35989 5687 36023
rect 5629 35983 5687 35989
rect 6454 35980 6460 36032
rect 6512 35980 6518 36032
rect 6733 36023 6791 36029
rect 6733 35989 6745 36023
rect 6779 36020 6791 36023
rect 7374 36020 7380 36032
rect 6779 35992 7380 36020
rect 6779 35989 6791 35992
rect 6733 35983 6791 35989
rect 7374 35980 7380 35992
rect 7432 35980 7438 36032
rect 7929 36023 7987 36029
rect 7929 35989 7941 36023
rect 7975 36020 7987 36023
rect 8110 36020 8116 36032
rect 7975 35992 8116 36020
rect 7975 35989 7987 35992
rect 7929 35983 7987 35989
rect 8110 35980 8116 35992
rect 8168 35980 8174 36032
rect 8386 35980 8392 36032
rect 8444 35980 8450 36032
rect 8478 35980 8484 36032
rect 8536 36020 8542 36032
rect 8846 36020 8852 36032
rect 8536 35992 8852 36020
rect 8536 35980 8542 35992
rect 8846 35980 8852 35992
rect 8904 35980 8910 36032
rect 9122 35980 9128 36032
rect 9180 36020 9186 36032
rect 9401 36023 9459 36029
rect 9401 36020 9413 36023
rect 9180 35992 9413 36020
rect 9180 35980 9186 35992
rect 9401 35989 9413 35992
rect 9447 35989 9459 36023
rect 9401 35983 9459 35989
rect 10318 35980 10324 36032
rect 10376 36020 10382 36032
rect 10502 36020 10508 36032
rect 10376 35992 10508 36020
rect 10376 35980 10382 35992
rect 10502 35980 10508 35992
rect 10560 35980 10566 36032
rect 11349 36020 11377 36187
rect 11440 36088 11468 36187
rect 11624 36165 11652 36264
rect 11882 36184 11888 36236
rect 11940 36184 11946 36236
rect 11974 36184 11980 36236
rect 12032 36184 12038 36236
rect 11609 36159 11667 36165
rect 11609 36125 11621 36159
rect 11655 36156 11667 36159
rect 12066 36156 12072 36168
rect 11655 36128 12072 36156
rect 11655 36125 11667 36128
rect 11609 36119 11667 36125
rect 12066 36116 12072 36128
rect 12124 36116 12130 36168
rect 11698 36088 11704 36100
rect 11440 36060 11704 36088
rect 11698 36048 11704 36060
rect 11756 36088 11762 36100
rect 12710 36088 12716 36100
rect 11756 36060 12716 36088
rect 11756 36048 11762 36060
rect 12710 36048 12716 36060
rect 12768 36048 12774 36100
rect 12158 36020 12164 36032
rect 11349 35992 12164 36020
rect 12158 35980 12164 35992
rect 12216 36020 12222 36032
rect 12618 36020 12624 36032
rect 12216 35992 12624 36020
rect 12216 35980 12222 35992
rect 12618 35980 12624 35992
rect 12676 35980 12682 36032
rect 552 35930 12604 35952
rect 552 35878 3662 35930
rect 3714 35878 3726 35930
rect 3778 35878 3790 35930
rect 3842 35878 3854 35930
rect 3906 35878 3918 35930
rect 3970 35878 10062 35930
rect 10114 35878 10126 35930
rect 10178 35878 10190 35930
rect 10242 35878 10254 35930
rect 10306 35878 10318 35930
rect 10370 35878 12604 35930
rect 552 35856 12604 35878
rect 937 35819 995 35825
rect 937 35785 949 35819
rect 983 35816 995 35819
rect 1026 35816 1032 35828
rect 983 35788 1032 35816
rect 983 35785 995 35788
rect 937 35779 995 35785
rect 1026 35776 1032 35788
rect 1084 35776 1090 35828
rect 1578 35776 1584 35828
rect 1636 35776 1642 35828
rect 2406 35776 2412 35828
rect 2464 35816 2470 35828
rect 2682 35816 2688 35828
rect 2464 35788 2688 35816
rect 2464 35776 2470 35788
rect 2682 35776 2688 35788
rect 2740 35776 2746 35828
rect 5813 35819 5871 35825
rect 5813 35785 5825 35819
rect 5859 35816 5871 35819
rect 6362 35816 6368 35828
rect 5859 35788 6368 35816
rect 5859 35785 5871 35788
rect 5813 35779 5871 35785
rect 6362 35776 6368 35788
rect 6420 35776 6426 35828
rect 6730 35776 6736 35828
rect 6788 35776 6794 35828
rect 7098 35776 7104 35828
rect 7156 35816 7162 35828
rect 7745 35819 7803 35825
rect 7745 35816 7757 35819
rect 7156 35788 7757 35816
rect 7156 35776 7162 35788
rect 7745 35785 7757 35788
rect 7791 35785 7803 35819
rect 7745 35779 7803 35785
rect 8386 35776 8392 35828
rect 8444 35816 8450 35828
rect 9493 35819 9551 35825
rect 9493 35816 9505 35819
rect 8444 35788 9505 35816
rect 8444 35776 8450 35788
rect 9493 35785 9505 35788
rect 9539 35785 9551 35819
rect 9493 35779 9551 35785
rect 9674 35776 9680 35828
rect 9732 35776 9738 35828
rect 9950 35776 9956 35828
rect 10008 35816 10014 35828
rect 10229 35819 10287 35825
rect 10229 35816 10241 35819
rect 10008 35788 10241 35816
rect 10008 35776 10014 35788
rect 10229 35785 10241 35788
rect 10275 35785 10287 35819
rect 10229 35779 10287 35785
rect 10410 35776 10416 35828
rect 10468 35776 10474 35828
rect 11514 35816 11520 35828
rect 10704 35788 11520 35816
rect 3050 35708 3056 35760
rect 3108 35748 3114 35760
rect 3786 35748 3792 35760
rect 3108 35720 3792 35748
rect 3108 35708 3114 35720
rect 3786 35708 3792 35720
rect 3844 35708 3850 35760
rect 4062 35708 4068 35760
rect 4120 35748 4126 35760
rect 5721 35751 5779 35757
rect 4120 35720 4384 35748
rect 4120 35708 4126 35720
rect 1946 35640 1952 35692
rect 2004 35680 2010 35692
rect 2498 35680 2504 35692
rect 2004 35652 2504 35680
rect 2004 35640 2010 35652
rect 2498 35640 2504 35652
rect 2556 35680 2562 35692
rect 2682 35680 2688 35692
rect 2556 35652 2688 35680
rect 2556 35640 2562 35652
rect 2682 35640 2688 35652
rect 2740 35680 2746 35692
rect 3697 35683 3755 35689
rect 3697 35680 3709 35683
rect 2740 35652 3709 35680
rect 2740 35640 2746 35652
rect 3697 35649 3709 35652
rect 3743 35649 3755 35683
rect 3697 35643 3755 35649
rect 3878 35640 3884 35692
rect 3936 35640 3942 35692
rect 3970 35640 3976 35692
rect 4028 35680 4034 35692
rect 4356 35689 4384 35720
rect 5721 35717 5733 35751
rect 5767 35748 5779 35751
rect 6178 35748 6184 35760
rect 5767 35720 6184 35748
rect 5767 35717 5779 35720
rect 5721 35711 5779 35717
rect 6178 35708 6184 35720
rect 6236 35708 6242 35760
rect 4341 35683 4399 35689
rect 4028 35652 4292 35680
rect 4028 35640 4034 35652
rect 1762 35572 1768 35624
rect 1820 35612 1826 35624
rect 2774 35612 2780 35624
rect 1820 35584 2780 35612
rect 1820 35572 1826 35584
rect 2774 35572 2780 35584
rect 2832 35572 2838 35624
rect 4264 35621 4292 35652
rect 4341 35649 4353 35683
rect 4387 35649 4399 35683
rect 4341 35643 4399 35649
rect 6105 35652 6684 35680
rect 4065 35615 4123 35621
rect 4065 35581 4077 35615
rect 4111 35581 4123 35615
rect 4065 35575 4123 35581
rect 4249 35615 4307 35621
rect 4249 35581 4261 35615
rect 4295 35581 4307 35615
rect 4249 35575 4307 35581
rect 3050 35504 3056 35556
rect 3108 35504 3114 35556
rect 4080 35544 4108 35575
rect 5718 35572 5724 35624
rect 5776 35612 5782 35624
rect 6105 35621 6133 35652
rect 6656 35624 6684 35652
rect 5997 35615 6055 35621
rect 5997 35612 6009 35615
rect 5776 35584 6009 35612
rect 5776 35572 5782 35584
rect 5997 35581 6009 35584
rect 6043 35581 6055 35615
rect 5997 35575 6055 35581
rect 6089 35615 6147 35621
rect 6089 35581 6101 35615
rect 6135 35581 6147 35615
rect 6089 35575 6147 35581
rect 6178 35572 6184 35624
rect 6236 35572 6242 35624
rect 6454 35572 6460 35624
rect 6512 35572 6518 35624
rect 6638 35572 6644 35624
rect 6696 35572 6702 35624
rect 6748 35621 6776 35776
rect 7282 35748 7288 35760
rect 7024 35720 7288 35748
rect 6825 35683 6883 35689
rect 6825 35649 6837 35683
rect 6871 35680 6883 35683
rect 7024 35680 7052 35720
rect 7282 35708 7288 35720
rect 7340 35708 7346 35760
rect 7466 35708 7472 35760
rect 7524 35708 7530 35760
rect 9306 35708 9312 35760
rect 9364 35708 9370 35760
rect 9692 35748 9720 35776
rect 10137 35751 10195 35757
rect 9692 35720 10088 35748
rect 6871 35652 7052 35680
rect 7101 35683 7159 35689
rect 6871 35649 6883 35652
rect 6825 35643 6883 35649
rect 7101 35649 7113 35683
rect 7147 35649 7159 35683
rect 7101 35643 7159 35649
rect 8941 35683 8999 35689
rect 8941 35649 8953 35683
rect 8987 35680 8999 35683
rect 9769 35683 9827 35689
rect 8987 35652 9444 35680
rect 8987 35649 8999 35652
rect 8941 35643 8999 35649
rect 6733 35615 6791 35621
rect 6733 35581 6745 35615
rect 6779 35581 6791 35615
rect 7116 35612 7144 35643
rect 7190 35612 7196 35624
rect 7116 35584 7196 35612
rect 6733 35575 6791 35581
rect 7190 35572 7196 35584
rect 7248 35572 7254 35624
rect 7929 35615 7987 35621
rect 7929 35581 7941 35615
rect 7975 35612 7987 35615
rect 8754 35612 8760 35624
rect 7975 35584 8760 35612
rect 7975 35581 7987 35584
rect 7929 35575 7987 35581
rect 8754 35572 8760 35584
rect 8812 35612 8818 35624
rect 9122 35612 9128 35624
rect 8812 35584 9128 35612
rect 8812 35572 8818 35584
rect 9122 35572 9128 35584
rect 9180 35572 9186 35624
rect 9416 35621 9444 35652
rect 9769 35649 9781 35683
rect 9815 35649 9827 35683
rect 10060 35680 10088 35720
rect 10137 35717 10149 35751
rect 10183 35748 10195 35751
rect 10704 35748 10732 35788
rect 11514 35776 11520 35788
rect 11572 35816 11578 35828
rect 11882 35816 11888 35828
rect 11572 35788 11888 35816
rect 11572 35776 11578 35788
rect 11882 35776 11888 35788
rect 11940 35776 11946 35828
rect 10183 35720 10732 35748
rect 10183 35717 10195 35720
rect 10137 35711 10195 35717
rect 10870 35708 10876 35760
rect 10928 35708 10934 35760
rect 10226 35680 10232 35692
rect 10060 35652 10232 35680
rect 9769 35643 9827 35649
rect 9401 35615 9459 35621
rect 9401 35581 9413 35615
rect 9447 35612 9459 35615
rect 9490 35612 9496 35624
rect 9447 35584 9496 35612
rect 9447 35581 9459 35584
rect 9401 35575 9459 35581
rect 9490 35572 9496 35584
rect 9548 35572 9554 35624
rect 9674 35572 9680 35624
rect 9732 35572 9738 35624
rect 4608 35547 4666 35553
rect 4080 35516 4568 35544
rect 3234 35436 3240 35488
rect 3292 35436 3298 35488
rect 3602 35436 3608 35488
rect 3660 35436 3666 35488
rect 4249 35479 4307 35485
rect 4249 35445 4261 35479
rect 4295 35476 4307 35479
rect 4338 35476 4344 35488
rect 4295 35448 4344 35476
rect 4295 35445 4307 35448
rect 4249 35439 4307 35445
rect 4338 35436 4344 35448
rect 4396 35436 4402 35488
rect 4540 35476 4568 35516
rect 4608 35513 4620 35547
rect 4654 35544 4666 35547
rect 4706 35544 4712 35556
rect 4654 35516 4712 35544
rect 4654 35513 4666 35516
rect 4608 35507 4666 35513
rect 4706 35504 4712 35516
rect 4764 35504 4770 35556
rect 4982 35504 4988 35556
rect 5040 35544 5046 35556
rect 5626 35544 5632 35556
rect 5040 35516 5632 35544
rect 5040 35504 5046 35516
rect 5626 35504 5632 35516
rect 5684 35504 5690 35556
rect 6319 35547 6377 35553
rect 6319 35513 6331 35547
rect 6365 35513 6377 35547
rect 6319 35507 6377 35513
rect 5994 35476 6000 35488
rect 4540 35448 6000 35476
rect 5994 35436 6000 35448
rect 6052 35436 6058 35488
rect 6178 35436 6184 35488
rect 6236 35476 6242 35488
rect 6334 35476 6362 35507
rect 7282 35504 7288 35556
rect 7340 35504 7346 35556
rect 8110 35504 8116 35556
rect 8168 35504 8174 35556
rect 8202 35504 8208 35556
rect 8260 35544 8266 35556
rect 8389 35547 8447 35553
rect 8389 35544 8401 35547
rect 8260 35516 8401 35544
rect 8260 35504 8266 35516
rect 8389 35513 8401 35516
rect 8435 35513 8447 35547
rect 8389 35507 8447 35513
rect 8570 35504 8576 35556
rect 8628 35504 8634 35556
rect 8846 35504 8852 35556
rect 8904 35544 8910 35556
rect 9784 35544 9812 35643
rect 10226 35640 10232 35652
rect 10284 35640 10290 35692
rect 10318 35640 10324 35692
rect 10376 35680 10382 35692
rect 10505 35683 10563 35689
rect 10505 35680 10517 35683
rect 10376 35652 10517 35680
rect 10376 35640 10382 35652
rect 10505 35649 10517 35652
rect 10551 35649 10563 35683
rect 10505 35643 10563 35649
rect 9858 35572 9864 35624
rect 9916 35612 9922 35624
rect 9953 35615 10011 35621
rect 9953 35612 9965 35615
rect 9916 35584 9965 35612
rect 9916 35572 9922 35584
rect 9953 35581 9965 35584
rect 9999 35581 10011 35615
rect 9953 35575 10011 35581
rect 10134 35572 10140 35624
rect 10192 35612 10198 35624
rect 10413 35615 10471 35621
rect 10413 35612 10425 35615
rect 10192 35584 10425 35612
rect 10192 35572 10198 35584
rect 10413 35581 10425 35584
rect 10459 35581 10471 35615
rect 10413 35575 10471 35581
rect 10594 35572 10600 35624
rect 10652 35612 10658 35624
rect 12253 35615 12311 35621
rect 12253 35612 12265 35615
rect 10652 35584 12265 35612
rect 10652 35572 10658 35584
rect 12253 35581 12265 35584
rect 12299 35581 12311 35615
rect 12253 35575 12311 35581
rect 10042 35544 10048 35556
rect 8904 35516 10048 35544
rect 8904 35504 8910 35516
rect 10042 35504 10048 35516
rect 10100 35504 10106 35556
rect 10502 35504 10508 35556
rect 10560 35544 10566 35556
rect 10689 35547 10747 35553
rect 10689 35544 10701 35547
rect 10560 35516 10701 35544
rect 10560 35504 10566 35516
rect 10689 35513 10701 35516
rect 10735 35513 10747 35547
rect 10689 35507 10747 35513
rect 11986 35547 12044 35553
rect 11986 35513 11998 35547
rect 12032 35513 12044 35547
rect 11986 35507 12044 35513
rect 6236 35448 6362 35476
rect 6236 35436 6242 35448
rect 8662 35436 8668 35488
rect 8720 35476 8726 35488
rect 9306 35476 9312 35488
rect 8720 35448 9312 35476
rect 8720 35436 8726 35448
rect 9306 35436 9312 35448
rect 9364 35476 9370 35488
rect 10870 35476 10876 35488
rect 9364 35448 10876 35476
rect 9364 35436 9370 35448
rect 10870 35436 10876 35448
rect 10928 35476 10934 35488
rect 11882 35476 11888 35488
rect 10928 35448 11888 35476
rect 10928 35436 10934 35448
rect 11882 35436 11888 35448
rect 11940 35436 11946 35488
rect 11992 35476 12020 35507
rect 12066 35476 12072 35488
rect 11992 35448 12072 35476
rect 12066 35436 12072 35448
rect 12124 35436 12130 35488
rect 552 35386 12604 35408
rect 552 35334 4322 35386
rect 4374 35334 4386 35386
rect 4438 35334 4450 35386
rect 4502 35334 4514 35386
rect 4566 35334 4578 35386
rect 4630 35334 10722 35386
rect 10774 35334 10786 35386
rect 10838 35334 10850 35386
rect 10902 35334 10914 35386
rect 10966 35334 10978 35386
rect 11030 35334 12604 35386
rect 552 35312 12604 35334
rect 658 35232 664 35284
rect 716 35272 722 35284
rect 937 35275 995 35281
rect 937 35272 949 35275
rect 716 35244 949 35272
rect 716 35232 722 35244
rect 937 35241 949 35244
rect 983 35241 995 35275
rect 937 35235 995 35241
rect 1118 35232 1124 35284
rect 1176 35232 1182 35284
rect 1486 35232 1492 35284
rect 1544 35272 1550 35284
rect 2225 35275 2283 35281
rect 2225 35272 2237 35275
rect 1544 35244 2237 35272
rect 1544 35232 1550 35244
rect 2225 35241 2237 35244
rect 2271 35241 2283 35275
rect 2225 35235 2283 35241
rect 2774 35232 2780 35284
rect 2832 35272 2838 35284
rect 3697 35275 3755 35281
rect 3697 35272 3709 35275
rect 2832 35244 3709 35272
rect 2832 35232 2838 35244
rect 3697 35241 3709 35244
rect 3743 35241 3755 35275
rect 3697 35235 3755 35241
rect 4062 35232 4068 35284
rect 4120 35232 4126 35284
rect 4154 35232 4160 35284
rect 4212 35272 4218 35284
rect 4338 35272 4344 35284
rect 4212 35244 4344 35272
rect 4212 35232 4218 35244
rect 4338 35232 4344 35244
rect 4396 35232 4402 35284
rect 4525 35275 4583 35281
rect 4525 35241 4537 35275
rect 4571 35272 4583 35275
rect 4706 35272 4712 35284
rect 4571 35244 4712 35272
rect 4571 35241 4583 35244
rect 4525 35235 4583 35241
rect 4706 35232 4712 35244
rect 4764 35232 4770 35284
rect 4816 35244 5396 35272
rect 1026 35096 1032 35148
rect 1084 35096 1090 35148
rect 1136 35145 1164 35232
rect 2130 35204 2136 35216
rect 1596 35176 2136 35204
rect 1121 35139 1179 35145
rect 1121 35105 1133 35139
rect 1167 35105 1179 35139
rect 1121 35099 1179 35105
rect 1486 35096 1492 35148
rect 1544 35136 1550 35148
rect 1596 35145 1624 35176
rect 2130 35164 2136 35176
rect 2188 35164 2194 35216
rect 3234 35164 3240 35216
rect 3292 35204 3298 35216
rect 3338 35207 3396 35213
rect 3338 35204 3350 35207
rect 3292 35176 3350 35204
rect 3292 35164 3298 35176
rect 3338 35173 3350 35176
rect 3384 35173 3396 35207
rect 4246 35204 4252 35216
rect 3338 35167 3396 35173
rect 3620 35176 4252 35204
rect 1581 35139 1639 35145
rect 1581 35136 1593 35139
rect 1544 35108 1593 35136
rect 1544 35096 1550 35108
rect 1581 35105 1593 35108
rect 1627 35105 1639 35139
rect 1581 35099 1639 35105
rect 1762 35096 1768 35148
rect 1820 35096 1826 35148
rect 1946 35096 1952 35148
rect 2004 35136 2010 35148
rect 3620 35145 3648 35176
rect 4246 35164 4252 35176
rect 4304 35164 4310 35216
rect 4816 35204 4844 35244
rect 5261 35207 5319 35213
rect 5261 35204 5273 35207
rect 4387 35176 4844 35204
rect 5092 35176 5273 35204
rect 3605 35139 3663 35145
rect 2004 35108 3556 35136
rect 2004 35096 2010 35108
rect 1210 35028 1216 35080
rect 1268 35068 1274 35080
rect 1857 35071 1915 35077
rect 1857 35068 1869 35071
rect 1268 35040 1869 35068
rect 1268 35028 1274 35040
rect 1857 35037 1869 35040
rect 1903 35037 1915 35071
rect 3528 35068 3556 35108
rect 3605 35105 3617 35139
rect 3651 35105 3663 35139
rect 3605 35099 3663 35105
rect 3878 35096 3884 35148
rect 3936 35136 3942 35148
rect 4387 35136 4415 35176
rect 3936 35108 4415 35136
rect 4709 35139 4767 35145
rect 3936 35096 3942 35108
rect 3786 35068 3792 35080
rect 3528 35040 3792 35068
rect 1857 35031 1915 35037
rect 3786 35028 3792 35040
rect 3844 35068 3850 35080
rect 4264 35077 4292 35108
rect 4709 35105 4721 35139
rect 4755 35136 4767 35139
rect 4890 35136 4896 35148
rect 4755 35108 4896 35136
rect 4755 35105 4767 35108
rect 4709 35099 4767 35105
rect 4890 35096 4896 35108
rect 4948 35096 4954 35148
rect 4985 35139 5043 35145
rect 4985 35105 4997 35139
rect 5031 35105 5043 35139
rect 4985 35099 5043 35105
rect 4157 35071 4215 35077
rect 4157 35068 4169 35071
rect 3844 35040 4169 35068
rect 3844 35028 3850 35040
rect 4157 35037 4169 35040
rect 4203 35037 4215 35071
rect 4157 35031 4215 35037
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35037 4307 35071
rect 4249 35031 4307 35037
rect 4338 35028 4344 35080
rect 4396 35068 4402 35080
rect 5000 35068 5028 35099
rect 4396 35040 5028 35068
rect 4396 35028 4402 35040
rect 5092 35000 5120 35176
rect 5261 35173 5273 35176
rect 5307 35173 5319 35207
rect 5261 35167 5319 35173
rect 5169 35139 5227 35145
rect 5169 35105 5181 35139
rect 5215 35136 5227 35139
rect 5368 35136 5396 35244
rect 5994 35232 6000 35284
rect 6052 35232 6058 35284
rect 6454 35232 6460 35284
rect 6512 35272 6518 35284
rect 6641 35275 6699 35281
rect 6641 35272 6653 35275
rect 6512 35244 6653 35272
rect 6512 35232 6518 35244
rect 6641 35241 6653 35244
rect 6687 35241 6699 35275
rect 6641 35235 6699 35241
rect 6730 35232 6736 35284
rect 6788 35272 6794 35284
rect 6788 35244 9168 35272
rect 6788 35232 6794 35244
rect 6270 35204 6276 35216
rect 6012 35176 6276 35204
rect 5215 35108 5396 35136
rect 5445 35139 5503 35145
rect 5215 35105 5227 35108
rect 5169 35099 5227 35105
rect 3988 34972 5120 35000
rect 5276 35000 5304 35108
rect 5445 35105 5457 35139
rect 5491 35105 5503 35139
rect 5445 35099 5503 35105
rect 5460 35068 5488 35099
rect 5534 35096 5540 35148
rect 5592 35096 5598 35148
rect 5810 35096 5816 35148
rect 5868 35096 5874 35148
rect 6012 35145 6040 35176
rect 6270 35164 6276 35176
rect 6328 35164 6334 35216
rect 6546 35164 6552 35216
rect 6604 35204 6610 35216
rect 9140 35213 9168 35244
rect 9490 35232 9496 35284
rect 9548 35232 9554 35284
rect 9674 35232 9680 35284
rect 9732 35272 9738 35284
rect 9732 35244 11376 35272
rect 9732 35232 9738 35244
rect 7653 35207 7711 35213
rect 7653 35204 7665 35207
rect 6604 35176 7665 35204
rect 6604 35164 6610 35176
rect 7653 35173 7665 35176
rect 7699 35173 7711 35207
rect 7653 35167 7711 35173
rect 9125 35207 9183 35213
rect 9125 35173 9137 35207
rect 9171 35173 9183 35207
rect 9508 35204 9536 35232
rect 9950 35204 9956 35216
rect 9508 35176 9956 35204
rect 9125 35167 9183 35173
rect 5997 35139 6055 35145
rect 5997 35105 6009 35139
rect 6043 35105 6055 35139
rect 5997 35099 6055 35105
rect 6089 35139 6147 35145
rect 6089 35105 6101 35139
rect 6135 35105 6147 35139
rect 6089 35099 6147 35105
rect 6825 35139 6883 35145
rect 6825 35105 6837 35139
rect 6871 35105 6883 35139
rect 6825 35099 6883 35105
rect 5460 35040 5580 35068
rect 5442 35000 5448 35012
rect 5276 34972 5448 35000
rect 1118 34892 1124 34944
rect 1176 34932 1182 34944
rect 3988 34932 4016 34972
rect 5442 34960 5448 34972
rect 5500 34960 5506 35012
rect 1176 34904 4016 34932
rect 1176 34892 1182 34904
rect 4706 34892 4712 34944
rect 4764 34932 4770 34944
rect 4982 34932 4988 34944
rect 4764 34904 4988 34932
rect 4764 34892 4770 34904
rect 4982 34892 4988 34904
rect 5040 34892 5046 34944
rect 5258 34892 5264 34944
rect 5316 34892 5322 34944
rect 5552 34932 5580 35040
rect 5626 35028 5632 35080
rect 5684 35068 5690 35080
rect 6104 35068 6132 35099
rect 5684 35040 6132 35068
rect 6365 35071 6423 35077
rect 5684 35028 5690 35040
rect 6365 35037 6377 35071
rect 6411 35037 6423 35071
rect 6365 35031 6423 35037
rect 6380 35000 6408 35031
rect 6546 35028 6552 35080
rect 6604 35068 6610 35080
rect 6840 35068 6868 35099
rect 6914 35096 6920 35148
rect 6972 35136 6978 35148
rect 7009 35139 7067 35145
rect 7009 35136 7021 35139
rect 6972 35108 7021 35136
rect 6972 35096 6978 35108
rect 7009 35105 7021 35108
rect 7055 35105 7067 35139
rect 7009 35099 7067 35105
rect 7098 35096 7104 35148
rect 7156 35096 7162 35148
rect 7466 35096 7472 35148
rect 7524 35096 7530 35148
rect 7558 35096 7564 35148
rect 7616 35136 7622 35148
rect 7837 35139 7895 35145
rect 7837 35136 7849 35139
rect 7616 35108 7849 35136
rect 7616 35096 7622 35108
rect 7837 35105 7849 35108
rect 7883 35105 7895 35139
rect 7837 35099 7895 35105
rect 8478 35096 8484 35148
rect 8536 35136 8542 35148
rect 8757 35139 8815 35145
rect 8757 35136 8769 35139
rect 8536 35108 8769 35136
rect 8536 35096 8542 35108
rect 8757 35105 8769 35108
rect 8803 35105 8815 35139
rect 8757 35099 8815 35105
rect 8941 35139 8999 35145
rect 8941 35105 8953 35139
rect 8987 35136 8999 35139
rect 9306 35136 9312 35148
rect 8987 35108 9312 35136
rect 8987 35105 8999 35108
rect 8941 35099 8999 35105
rect 9306 35096 9312 35108
rect 9364 35096 9370 35148
rect 9398 35096 9404 35148
rect 9456 35136 9462 35148
rect 9600 35145 9628 35176
rect 9950 35164 9956 35176
rect 10008 35204 10014 35216
rect 10134 35204 10140 35216
rect 10008 35176 10140 35204
rect 10008 35164 10014 35176
rect 10134 35164 10140 35176
rect 10192 35164 10198 35216
rect 10410 35164 10416 35216
rect 10468 35204 10474 35216
rect 11348 35204 11376 35244
rect 11790 35232 11796 35284
rect 11848 35272 11854 35284
rect 12158 35272 12164 35284
rect 11848 35244 12164 35272
rect 11848 35232 11854 35244
rect 12158 35232 12164 35244
rect 12216 35232 12222 35284
rect 11974 35204 11980 35216
rect 10468 35176 11284 35204
rect 11348 35176 11980 35204
rect 10468 35164 10474 35176
rect 9493 35139 9551 35145
rect 9493 35136 9505 35139
rect 9456 35108 9505 35136
rect 9456 35096 9462 35108
rect 9493 35105 9505 35108
rect 9539 35105 9551 35139
rect 9493 35099 9551 35105
rect 9585 35139 9643 35145
rect 9585 35105 9597 35139
rect 9631 35105 9643 35139
rect 10153 35134 10181 35164
rect 10229 35139 10287 35145
rect 10229 35134 10241 35139
rect 10153 35106 10241 35134
rect 9585 35099 9643 35105
rect 10229 35105 10241 35106
rect 10275 35105 10287 35139
rect 10229 35099 10287 35105
rect 11146 35096 11152 35148
rect 11204 35096 11210 35148
rect 11256 35145 11284 35176
rect 11974 35164 11980 35176
rect 12032 35213 12038 35216
rect 12032 35207 12095 35213
rect 12032 35173 12049 35207
rect 12083 35173 12095 35207
rect 12032 35167 12095 35173
rect 12032 35164 12038 35167
rect 12250 35164 12256 35216
rect 12308 35164 12314 35216
rect 11241 35139 11299 35145
rect 11241 35105 11253 35139
rect 11287 35105 11299 35139
rect 11241 35099 11299 35105
rect 11422 35096 11428 35148
rect 11480 35096 11486 35148
rect 11609 35139 11667 35145
rect 11609 35105 11621 35139
rect 11655 35105 11667 35139
rect 11609 35099 11667 35105
rect 7193 35071 7251 35077
rect 7193 35068 7205 35071
rect 6604 35040 7205 35068
rect 6604 35028 6610 35040
rect 7193 35037 7205 35040
rect 7239 35037 7251 35071
rect 7193 35031 7251 35037
rect 7374 35028 7380 35080
rect 7432 35068 7438 35080
rect 8297 35071 8355 35077
rect 8297 35068 8309 35071
rect 7432 35040 8309 35068
rect 7432 35028 7438 35040
rect 8297 35037 8309 35040
rect 8343 35037 8355 35071
rect 9674 35068 9680 35080
rect 8297 35031 8355 35037
rect 8772 35040 9680 35068
rect 6638 35000 6644 35012
rect 6380 34972 6644 35000
rect 6638 34960 6644 34972
rect 6696 34960 6702 35012
rect 6730 34960 6736 35012
rect 6788 35000 6794 35012
rect 7466 35000 7472 35012
rect 6788 34972 7472 35000
rect 6788 34960 6794 34972
rect 7466 34960 7472 34972
rect 7524 34960 7530 35012
rect 7742 34960 7748 35012
rect 7800 35000 7806 35012
rect 8772 35000 8800 35040
rect 9674 35028 9680 35040
rect 9732 35028 9738 35080
rect 9769 35071 9827 35077
rect 9769 35037 9781 35071
rect 9815 35037 9827 35071
rect 9769 35031 9827 35037
rect 7800 34972 8800 35000
rect 7800 34960 7806 34972
rect 8846 34960 8852 35012
rect 8904 35000 8910 35012
rect 9784 35000 9812 35031
rect 9858 35028 9864 35080
rect 9916 35068 9922 35080
rect 10137 35071 10195 35077
rect 10137 35068 10149 35071
rect 9916 35040 10149 35068
rect 9916 35028 9922 35040
rect 10137 35037 10149 35040
rect 10183 35037 10195 35071
rect 10137 35031 10195 35037
rect 10597 35003 10655 35009
rect 8904 34972 10088 35000
rect 8904 34960 8910 34972
rect 6362 34932 6368 34944
rect 5552 34904 6368 34932
rect 6362 34892 6368 34904
rect 6420 34892 6426 34944
rect 6914 34892 6920 34944
rect 6972 34932 6978 34944
rect 7282 34932 7288 34944
rect 6972 34904 7288 34932
rect 6972 34892 6978 34904
rect 7282 34892 7288 34904
rect 7340 34892 7346 34944
rect 7926 34892 7932 34944
rect 7984 34892 7990 34944
rect 8665 34935 8723 34941
rect 8665 34901 8677 34935
rect 8711 34932 8723 34935
rect 9306 34932 9312 34944
rect 8711 34904 9312 34932
rect 8711 34901 8723 34904
rect 8665 34895 8723 34901
rect 9306 34892 9312 34904
rect 9364 34892 9370 34944
rect 9858 34892 9864 34944
rect 9916 34932 9922 34944
rect 9953 34935 10011 34941
rect 9953 34932 9965 34935
rect 9916 34904 9965 34932
rect 9916 34892 9922 34904
rect 9953 34901 9965 34904
rect 9999 34901 10011 34935
rect 10060 34932 10088 34972
rect 10597 34969 10609 35003
rect 10643 35000 10655 35003
rect 11624 35000 11652 35099
rect 11882 35028 11888 35080
rect 11940 35068 11946 35080
rect 11940 35040 12112 35068
rect 11940 35028 11946 35040
rect 10643 34972 11652 35000
rect 11793 35003 11851 35009
rect 10643 34969 10655 34972
rect 10597 34963 10655 34969
rect 11793 34969 11805 35003
rect 11839 35000 11851 35003
rect 11974 35000 11980 35012
rect 11839 34972 11980 35000
rect 11839 34969 11851 34972
rect 11793 34963 11851 34969
rect 11974 34960 11980 34972
rect 12032 34960 12038 35012
rect 10965 34935 11023 34941
rect 10965 34932 10977 34935
rect 10060 34904 10977 34932
rect 9953 34895 10011 34901
rect 10965 34901 10977 34904
rect 11011 34901 11023 34935
rect 10965 34895 11023 34901
rect 11330 34892 11336 34944
rect 11388 34932 11394 34944
rect 12084 34941 12112 35040
rect 11885 34935 11943 34941
rect 11885 34932 11897 34935
rect 11388 34904 11897 34932
rect 11388 34892 11394 34904
rect 11885 34901 11897 34904
rect 11931 34901 11943 34935
rect 11885 34895 11943 34901
rect 12069 34935 12127 34941
rect 12069 34901 12081 34935
rect 12115 34901 12127 34935
rect 12069 34895 12127 34901
rect 552 34842 12604 34864
rect 552 34790 3662 34842
rect 3714 34790 3726 34842
rect 3778 34790 3790 34842
rect 3842 34790 3854 34842
rect 3906 34790 3918 34842
rect 3970 34790 10062 34842
rect 10114 34790 10126 34842
rect 10178 34790 10190 34842
rect 10242 34790 10254 34842
rect 10306 34790 10318 34842
rect 10370 34790 12604 34842
rect 552 34768 12604 34790
rect 937 34731 995 34737
rect 937 34697 949 34731
rect 983 34728 995 34731
rect 1210 34728 1216 34740
rect 983 34700 1216 34728
rect 983 34697 995 34700
rect 937 34691 995 34697
rect 1210 34688 1216 34700
rect 1268 34688 1274 34740
rect 1394 34688 1400 34740
rect 1452 34688 1458 34740
rect 2038 34688 2044 34740
rect 2096 34728 2102 34740
rect 2590 34728 2596 34740
rect 2096 34700 2596 34728
rect 2096 34688 2102 34700
rect 2590 34688 2596 34700
rect 2648 34688 2654 34740
rect 3418 34688 3424 34740
rect 3476 34728 3482 34740
rect 3694 34728 3700 34740
rect 3476 34700 3700 34728
rect 3476 34688 3482 34700
rect 3694 34688 3700 34700
rect 3752 34688 3758 34740
rect 4525 34731 4583 34737
rect 4525 34697 4537 34731
rect 4571 34728 4583 34731
rect 5350 34728 5356 34740
rect 4571 34700 4936 34728
rect 4571 34697 4583 34700
rect 4525 34691 4583 34697
rect 1412 34660 1440 34688
rect 400 34632 1440 34660
rect 400 34536 428 34632
rect 2406 34620 2412 34672
rect 2464 34660 2470 34672
rect 2501 34663 2559 34669
rect 2501 34660 2513 34663
rect 2464 34632 2513 34660
rect 2464 34620 2470 34632
rect 2501 34629 2513 34632
rect 2547 34629 2559 34663
rect 4706 34660 4712 34672
rect 2501 34623 2559 34629
rect 2884 34632 4712 34660
rect 382 34484 388 34536
rect 440 34484 446 34536
rect 1578 34484 1584 34536
rect 1636 34524 1642 34536
rect 2222 34524 2228 34536
rect 1636 34496 2228 34524
rect 1636 34484 1642 34496
rect 2222 34484 2228 34496
rect 2280 34524 2286 34536
rect 2884 34533 2912 34632
rect 4706 34620 4712 34632
rect 4764 34620 4770 34672
rect 2961 34595 3019 34601
rect 2961 34561 2973 34595
rect 3007 34592 3019 34595
rect 3050 34592 3056 34604
rect 3007 34564 3056 34592
rect 3007 34561 3019 34564
rect 2961 34555 3019 34561
rect 3050 34552 3056 34564
rect 3108 34552 3114 34604
rect 3786 34552 3792 34604
rect 3844 34552 3850 34604
rect 4246 34592 4252 34604
rect 3896 34564 4252 34592
rect 2317 34527 2375 34533
rect 2317 34524 2329 34527
rect 2280 34496 2329 34524
rect 2280 34484 2286 34496
rect 2317 34493 2329 34496
rect 2363 34493 2375 34527
rect 2317 34487 2375 34493
rect 2869 34527 2927 34533
rect 2869 34493 2881 34527
rect 2915 34493 2927 34527
rect 2869 34487 2927 34493
rect 1762 34416 1768 34468
rect 1820 34456 1826 34468
rect 2050 34459 2108 34465
rect 2050 34456 2062 34459
rect 1820 34428 2062 34456
rect 1820 34416 1826 34428
rect 2050 34425 2062 34428
rect 2096 34425 2108 34459
rect 2332 34456 2360 34487
rect 3510 34456 3516 34468
rect 2332 34428 3516 34456
rect 2050 34419 2108 34425
rect 3510 34416 3516 34428
rect 3568 34456 3574 34468
rect 3896 34456 3924 34564
rect 4246 34552 4252 34564
rect 4304 34552 4310 34604
rect 4157 34527 4215 34533
rect 4157 34493 4169 34527
rect 4203 34493 4215 34527
rect 4908 34524 4936 34700
rect 5000 34700 5356 34728
rect 5000 34601 5028 34700
rect 5350 34688 5356 34700
rect 5408 34688 5414 34740
rect 5810 34688 5816 34740
rect 5868 34688 5874 34740
rect 6733 34731 6791 34737
rect 6733 34697 6745 34731
rect 6779 34728 6791 34731
rect 7098 34728 7104 34740
rect 6779 34700 7104 34728
rect 6779 34697 6791 34700
rect 6733 34691 6791 34697
rect 7098 34688 7104 34700
rect 7156 34688 7162 34740
rect 8849 34731 8907 34737
rect 8849 34697 8861 34731
rect 8895 34728 8907 34731
rect 10134 34728 10140 34740
rect 8895 34700 10140 34728
rect 8895 34697 8907 34700
rect 8849 34691 8907 34697
rect 10134 34688 10140 34700
rect 10192 34688 10198 34740
rect 5994 34660 6000 34672
rect 5184 34632 6000 34660
rect 5184 34601 5212 34632
rect 5994 34620 6000 34632
rect 6052 34620 6058 34672
rect 6917 34663 6975 34669
rect 6917 34629 6929 34663
rect 6963 34660 6975 34663
rect 10413 34663 10471 34669
rect 10413 34660 10425 34663
rect 6963 34632 9076 34660
rect 6963 34629 6975 34632
rect 6917 34623 6975 34629
rect 4985 34595 5043 34601
rect 4985 34561 4997 34595
rect 5031 34561 5043 34595
rect 4985 34555 5043 34561
rect 5169 34595 5227 34601
rect 5169 34561 5181 34595
rect 5215 34561 5227 34595
rect 5169 34555 5227 34561
rect 5445 34595 5503 34601
rect 5445 34561 5457 34595
rect 5491 34592 5503 34595
rect 5534 34592 5540 34604
rect 5491 34564 5540 34592
rect 5491 34561 5503 34564
rect 5445 34555 5503 34561
rect 5534 34552 5540 34564
rect 5592 34552 5598 34604
rect 5902 34552 5908 34604
rect 5960 34592 5966 34604
rect 8846 34592 8852 34604
rect 5960 34564 6592 34592
rect 5960 34552 5966 34564
rect 4157 34487 4215 34493
rect 4264 34496 4936 34524
rect 3568 34428 3924 34456
rect 3568 34416 3574 34428
rect 4062 34416 4068 34468
rect 4120 34456 4126 34468
rect 4172 34456 4200 34487
rect 4120 34428 4200 34456
rect 4120 34416 4126 34428
rect 566 34348 572 34400
rect 624 34388 630 34400
rect 1854 34388 1860 34400
rect 624 34360 1860 34388
rect 624 34348 630 34360
rect 1854 34348 1860 34360
rect 1912 34348 1918 34400
rect 3234 34348 3240 34400
rect 3292 34348 3298 34400
rect 3418 34348 3424 34400
rect 3476 34388 3482 34400
rect 3605 34391 3663 34397
rect 3605 34388 3617 34391
rect 3476 34360 3617 34388
rect 3476 34348 3482 34360
rect 3605 34357 3617 34360
rect 3651 34357 3663 34391
rect 3605 34351 3663 34357
rect 3694 34348 3700 34400
rect 3752 34348 3758 34400
rect 4154 34348 4160 34400
rect 4212 34388 4218 34400
rect 4264 34388 4292 34496
rect 4525 34459 4583 34465
rect 4525 34425 4537 34459
rect 4571 34456 4583 34459
rect 4571 34428 4844 34456
rect 4571 34425 4583 34428
rect 4525 34419 4583 34425
rect 4212 34360 4292 34388
rect 4212 34348 4218 34360
rect 4706 34348 4712 34400
rect 4764 34348 4770 34400
rect 4816 34397 4844 34428
rect 4801 34391 4859 34397
rect 4801 34357 4813 34391
rect 4847 34357 4859 34391
rect 4908 34388 4936 34496
rect 5077 34527 5135 34533
rect 5077 34493 5089 34527
rect 5123 34493 5135 34527
rect 5077 34487 5135 34493
rect 5261 34527 5319 34533
rect 5261 34493 5273 34527
rect 5307 34524 5319 34527
rect 5920 34524 5948 34552
rect 5307 34496 5948 34524
rect 5307 34493 5319 34496
rect 5261 34487 5319 34493
rect 5092 34456 5120 34487
rect 6362 34484 6368 34536
rect 6420 34484 6426 34536
rect 6454 34484 6460 34536
rect 6512 34484 6518 34536
rect 6564 34533 6592 34564
rect 6840 34564 8852 34592
rect 6840 34533 6868 34564
rect 8846 34552 8852 34564
rect 8904 34552 8910 34604
rect 9048 34592 9076 34632
rect 10060 34632 10425 34660
rect 9048 34564 9161 34592
rect 6549 34527 6607 34533
rect 6549 34493 6561 34527
rect 6595 34493 6607 34527
rect 6549 34487 6607 34493
rect 6825 34527 6883 34533
rect 6825 34493 6837 34527
rect 6871 34493 6883 34527
rect 6825 34487 6883 34493
rect 7009 34527 7067 34533
rect 7009 34493 7021 34527
rect 7055 34493 7067 34527
rect 7009 34487 7067 34493
rect 5534 34456 5540 34468
rect 5092 34428 5540 34456
rect 5534 34416 5540 34428
rect 5592 34416 5598 34468
rect 5813 34459 5871 34465
rect 5813 34425 5825 34459
rect 5859 34456 5871 34459
rect 6730 34456 6736 34468
rect 5859 34428 6736 34456
rect 5859 34425 5871 34428
rect 5813 34419 5871 34425
rect 5828 34388 5856 34419
rect 6730 34416 6736 34428
rect 6788 34416 6794 34468
rect 6914 34416 6920 34468
rect 6972 34456 6978 34468
rect 7024 34456 7052 34487
rect 7374 34484 7380 34536
rect 7432 34484 7438 34536
rect 7650 34484 7656 34536
rect 7708 34484 7714 34536
rect 8202 34484 8208 34536
rect 8260 34484 8266 34536
rect 8573 34527 8631 34533
rect 8573 34524 8585 34527
rect 8312 34496 8585 34524
rect 7742 34456 7748 34468
rect 6972 34428 7748 34456
rect 6972 34416 6978 34428
rect 7742 34416 7748 34428
rect 7800 34416 7806 34468
rect 8018 34416 8024 34468
rect 8076 34456 8082 34468
rect 8312 34456 8340 34496
rect 8573 34493 8585 34496
rect 8619 34493 8631 34527
rect 8573 34487 8631 34493
rect 8665 34527 8723 34533
rect 8665 34493 8677 34527
rect 8711 34524 8723 34527
rect 8754 34524 8760 34536
rect 8711 34496 8760 34524
rect 8711 34493 8723 34496
rect 8665 34487 8723 34493
rect 8754 34484 8760 34496
rect 8812 34484 8818 34536
rect 8938 34484 8944 34536
rect 8996 34484 9002 34536
rect 9030 34484 9036 34536
rect 9088 34484 9094 34536
rect 9133 34524 9161 34564
rect 9766 34524 9772 34536
rect 9133 34496 9772 34524
rect 9766 34484 9772 34496
rect 9824 34484 9830 34536
rect 10060 34524 10088 34632
rect 10413 34629 10425 34632
rect 10459 34629 10471 34663
rect 10413 34623 10471 34629
rect 10428 34592 10456 34623
rect 10502 34620 10508 34672
rect 10560 34620 10566 34672
rect 10428 34564 10732 34592
rect 10704 34533 10732 34564
rect 9876 34496 10088 34524
rect 10505 34527 10563 34533
rect 8076 34428 8340 34456
rect 9300 34459 9358 34465
rect 8076 34416 8082 34428
rect 9300 34425 9312 34459
rect 9346 34456 9358 34459
rect 9398 34456 9404 34468
rect 9346 34428 9404 34456
rect 9346 34425 9358 34428
rect 9300 34419 9358 34425
rect 9398 34416 9404 34428
rect 9456 34416 9462 34468
rect 9490 34416 9496 34468
rect 9548 34456 9554 34468
rect 9876 34456 9904 34496
rect 10505 34493 10517 34527
rect 10551 34493 10563 34527
rect 10505 34487 10563 34493
rect 10689 34527 10747 34533
rect 10689 34493 10701 34527
rect 10735 34493 10747 34527
rect 10689 34487 10747 34493
rect 9548 34428 9904 34456
rect 9548 34416 9554 34428
rect 9950 34416 9956 34468
rect 10008 34456 10014 34468
rect 10410 34456 10416 34468
rect 10008 34428 10416 34456
rect 10008 34416 10014 34428
rect 10410 34416 10416 34428
rect 10468 34456 10474 34468
rect 10520 34456 10548 34487
rect 11974 34484 11980 34536
rect 12032 34533 12038 34536
rect 12032 34524 12044 34533
rect 12032 34496 12077 34524
rect 12032 34487 12044 34496
rect 12032 34484 12038 34487
rect 12250 34484 12256 34536
rect 12308 34484 12314 34536
rect 10468 34428 10916 34456
rect 10468 34416 10474 34428
rect 4908 34360 5856 34388
rect 5997 34391 6055 34397
rect 4801 34351 4859 34357
rect 5997 34357 6009 34391
rect 6043 34388 6055 34391
rect 6086 34388 6092 34400
rect 6043 34360 6092 34388
rect 6043 34357 6055 34360
rect 5997 34351 6055 34357
rect 6086 34348 6092 34360
rect 6144 34348 6150 34400
rect 6362 34348 6368 34400
rect 6420 34388 6426 34400
rect 7006 34388 7012 34400
rect 6420 34360 7012 34388
rect 6420 34348 6426 34360
rect 7006 34348 7012 34360
rect 7064 34348 7070 34400
rect 7834 34348 7840 34400
rect 7892 34388 7898 34400
rect 8389 34391 8447 34397
rect 8389 34388 8401 34391
rect 7892 34360 8401 34388
rect 7892 34348 7898 34360
rect 8389 34357 8401 34360
rect 8435 34357 8447 34391
rect 8389 34351 8447 34357
rect 9674 34348 9680 34400
rect 9732 34388 9738 34400
rect 10594 34388 10600 34400
rect 9732 34360 10600 34388
rect 9732 34348 9738 34360
rect 10594 34348 10600 34360
rect 10652 34348 10658 34400
rect 10888 34397 10916 34428
rect 11606 34416 11612 34468
rect 11664 34456 11670 34468
rect 11664 34428 12020 34456
rect 11664 34416 11670 34428
rect 11992 34400 12020 34428
rect 10873 34391 10931 34397
rect 10873 34357 10885 34391
rect 10919 34357 10931 34391
rect 10873 34351 10931 34357
rect 11146 34348 11152 34400
rect 11204 34388 11210 34400
rect 11790 34388 11796 34400
rect 11204 34360 11796 34388
rect 11204 34348 11210 34360
rect 11790 34348 11796 34360
rect 11848 34348 11854 34400
rect 11974 34348 11980 34400
rect 12032 34348 12038 34400
rect 552 34298 12604 34320
rect 552 34246 4322 34298
rect 4374 34246 4386 34298
rect 4438 34246 4450 34298
rect 4502 34246 4514 34298
rect 4566 34246 4578 34298
rect 4630 34246 10722 34298
rect 10774 34246 10786 34298
rect 10838 34246 10850 34298
rect 10902 34246 10914 34298
rect 10966 34246 10978 34298
rect 11030 34246 12604 34298
rect 552 34224 12604 34246
rect 937 34187 995 34193
rect 937 34153 949 34187
rect 983 34184 995 34187
rect 3326 34184 3332 34196
rect 983 34156 3332 34184
rect 983 34153 995 34156
rect 937 34147 995 34153
rect 3326 34144 3332 34156
rect 3384 34144 3390 34196
rect 3602 34144 3608 34196
rect 3660 34144 3666 34196
rect 6270 34184 6276 34196
rect 3804 34156 6276 34184
rect 842 34076 848 34128
rect 900 34116 906 34128
rect 1121 34119 1179 34125
rect 1121 34116 1133 34119
rect 900 34088 1133 34116
rect 900 34076 906 34088
rect 1121 34085 1133 34088
rect 1167 34085 1179 34119
rect 1121 34079 1179 34085
rect 1210 34076 1216 34128
rect 1268 34116 1274 34128
rect 2492 34119 2550 34125
rect 1268 34088 2360 34116
rect 1268 34076 1274 34088
rect 1026 34008 1032 34060
rect 1084 34008 1090 34060
rect 1486 34008 1492 34060
rect 1544 34048 1550 34060
rect 1581 34051 1639 34057
rect 1581 34048 1593 34051
rect 1544 34020 1593 34048
rect 1544 34008 1550 34020
rect 1581 34017 1593 34020
rect 1627 34017 1639 34051
rect 1581 34011 1639 34017
rect 1765 34051 1823 34057
rect 1765 34017 1777 34051
rect 1811 34048 1823 34051
rect 1946 34048 1952 34060
rect 1811 34020 1952 34048
rect 1811 34017 1823 34020
rect 1765 34011 1823 34017
rect 1946 34008 1952 34020
rect 2004 34008 2010 34060
rect 2222 34008 2228 34060
rect 2280 34008 2286 34060
rect 2332 34048 2360 34088
rect 2492 34085 2504 34119
rect 2538 34116 2550 34119
rect 3234 34116 3240 34128
rect 2538 34088 3240 34116
rect 2538 34085 2550 34088
rect 2492 34079 2550 34085
rect 3234 34076 3240 34088
rect 3292 34076 3298 34128
rect 3804 34125 3832 34156
rect 6270 34144 6276 34156
rect 6328 34144 6334 34196
rect 6638 34144 6644 34196
rect 6696 34184 6702 34196
rect 7558 34184 7564 34196
rect 6696 34156 7564 34184
rect 6696 34144 6702 34156
rect 7558 34144 7564 34156
rect 7616 34144 7622 34196
rect 7650 34144 7656 34196
rect 7708 34184 7714 34196
rect 9674 34184 9680 34196
rect 7708 34156 9680 34184
rect 7708 34144 7714 34156
rect 9674 34144 9680 34156
rect 9732 34144 9738 34196
rect 11238 34184 11244 34196
rect 9968 34156 11244 34184
rect 3789 34119 3847 34125
rect 3789 34116 3801 34119
rect 3344 34088 3801 34116
rect 3344 34048 3372 34088
rect 3789 34085 3801 34088
rect 3835 34085 3847 34119
rect 9030 34116 9036 34128
rect 3789 34079 3847 34085
rect 4019 34085 4077 34091
rect 4019 34082 4031 34085
rect 4004 34060 4031 34082
rect 2332 34020 3372 34048
rect 3418 34008 3424 34060
rect 3476 34048 3482 34060
rect 3970 34048 3976 34060
rect 3476 34020 3976 34048
rect 3476 34008 3482 34020
rect 3970 34008 3976 34020
rect 4028 34051 4031 34060
rect 4065 34051 4077 34085
rect 4264 34088 9036 34116
rect 4264 34057 4292 34088
rect 4522 34057 4528 34060
rect 4028 34045 4077 34051
rect 4249 34051 4307 34057
rect 4028 34008 4034 34045
rect 4249 34017 4261 34051
rect 4295 34017 4307 34051
rect 4516 34048 4528 34057
rect 4483 34020 4528 34048
rect 4249 34011 4307 34017
rect 4516 34011 4528 34020
rect 4522 34008 4528 34011
rect 4580 34008 4586 34060
rect 6012 34057 6040 34088
rect 9030 34076 9036 34088
rect 9088 34076 9094 34128
rect 9968 34116 9996 34156
rect 9232 34088 9996 34116
rect 5997 34051 6055 34057
rect 5997 34017 6009 34051
rect 6043 34017 6055 34051
rect 5997 34011 6055 34017
rect 6086 34008 6092 34060
rect 6144 34048 6150 34060
rect 6253 34051 6311 34057
rect 6253 34048 6265 34051
rect 6144 34020 6265 34048
rect 6144 34008 6150 34020
rect 6253 34017 6265 34020
rect 6299 34017 6311 34051
rect 6253 34011 6311 34017
rect 7374 34008 7380 34060
rect 7432 34048 7438 34060
rect 7469 34051 7527 34057
rect 7469 34048 7481 34051
rect 7432 34020 7481 34048
rect 7432 34008 7438 34020
rect 7469 34017 7481 34020
rect 7515 34017 7527 34051
rect 7469 34011 7527 34017
rect 7653 34051 7711 34057
rect 7653 34017 7665 34051
rect 7699 34017 7711 34051
rect 7653 34011 7711 34017
rect 14 33940 20 33992
rect 72 33980 78 33992
rect 842 33980 848 33992
rect 72 33952 848 33980
rect 72 33940 78 33952
rect 842 33940 848 33952
rect 900 33940 906 33992
rect 1857 33983 1915 33989
rect 1857 33949 1869 33983
rect 1903 33949 1915 33983
rect 1857 33943 1915 33949
rect 1872 33912 1900 33943
rect 5626 33940 5632 33992
rect 5684 33940 5690 33992
rect 4246 33912 4252 33924
rect 492 33884 1900 33912
rect 3896 33884 4252 33912
rect 492 33640 520 33884
rect 2406 33804 2412 33856
rect 2464 33844 2470 33856
rect 3896 33844 3924 33884
rect 4246 33872 4252 33884
rect 4304 33872 4310 33924
rect 2464 33816 3924 33844
rect 2464 33804 2470 33816
rect 3970 33804 3976 33856
rect 4028 33804 4034 33856
rect 4062 33804 4068 33856
rect 4120 33844 4126 33856
rect 5644 33853 5672 33940
rect 7668 33912 7696 34011
rect 8110 34008 8116 34060
rect 8168 34048 8174 34060
rect 8168 34020 8294 34048
rect 8168 34008 8174 34020
rect 7837 33983 7895 33989
rect 7837 33949 7849 33983
rect 7883 33980 7895 33983
rect 8018 33980 8024 33992
rect 7883 33952 8024 33980
rect 7883 33949 7895 33952
rect 7837 33943 7895 33949
rect 8018 33940 8024 33952
rect 8076 33940 8082 33992
rect 8266 33980 8294 34020
rect 8386 34008 8392 34060
rect 8444 34008 8450 34060
rect 9232 34048 9260 34088
rect 10042 34076 10048 34128
rect 10100 34082 10106 34128
rect 10100 34076 10121 34082
rect 10057 34073 10121 34076
rect 8680 34038 9260 34048
rect 8496 34020 9260 34038
rect 9309 34051 9367 34057
rect 8496 34010 8708 34020
rect 9309 34017 9321 34051
rect 9355 34048 9367 34051
rect 9490 34048 9496 34060
rect 9355 34020 9496 34048
rect 9355 34017 9367 34020
rect 9309 34011 9367 34017
rect 8496 33980 8524 34010
rect 9490 34008 9496 34020
rect 9548 34008 9554 34060
rect 9582 34008 9588 34060
rect 9640 34008 9646 34060
rect 9674 34008 9680 34060
rect 9732 34008 9738 34060
rect 9766 34008 9772 34060
rect 9824 34008 9830 34060
rect 9858 34008 9864 34060
rect 9916 34008 9922 34060
rect 10057 34039 10069 34073
rect 10103 34042 10121 34073
rect 10336 34057 10364 34156
rect 11238 34144 11244 34156
rect 11296 34144 11302 34196
rect 11422 34144 11428 34196
rect 11480 34144 11486 34196
rect 11655 34085 11713 34091
rect 10321 34051 10379 34057
rect 10103 34039 10115 34042
rect 10057 34033 10115 34039
rect 10321 34017 10333 34051
rect 10367 34017 10379 34051
rect 10321 34011 10379 34017
rect 10410 34008 10416 34060
rect 10468 34008 10474 34060
rect 11146 34008 11152 34060
rect 11204 34048 11210 34060
rect 11241 34051 11299 34057
rect 11241 34048 11253 34051
rect 11204 34020 11253 34048
rect 11204 34008 11210 34020
rect 11241 34017 11253 34020
rect 11287 34017 11299 34051
rect 11655 34051 11667 34085
rect 11701 34051 11713 34085
rect 11882 34076 11888 34128
rect 11940 34076 11946 34128
rect 11655 34045 11713 34051
rect 12161 34051 12219 34057
rect 11241 34011 11299 34017
rect 8266 33952 8524 33980
rect 9600 33980 9628 34008
rect 10505 33983 10563 33989
rect 10505 33980 10517 33983
rect 9600 33952 10517 33980
rect 10505 33949 10517 33952
rect 10551 33949 10563 33983
rect 10505 33943 10563 33949
rect 10594 33940 10600 33992
rect 10652 33940 10658 33992
rect 10778 33940 10784 33992
rect 10836 33980 10842 33992
rect 10965 33983 11023 33989
rect 10965 33980 10977 33983
rect 10836 33952 10977 33980
rect 10836 33940 10842 33952
rect 10965 33949 10977 33952
rect 11011 33980 11023 33983
rect 11330 33980 11336 33992
rect 11011 33952 11336 33980
rect 11011 33949 11023 33952
rect 10965 33943 11023 33949
rect 11330 33940 11336 33952
rect 11388 33980 11394 33992
rect 11684 33980 11712 34045
rect 12161 34017 12173 34051
rect 12207 34017 12219 34051
rect 12161 34011 12219 34017
rect 11388 33952 11712 33980
rect 11388 33940 11394 33952
rect 8478 33912 8484 33924
rect 7668 33884 8484 33912
rect 8478 33872 8484 33884
rect 8536 33872 8542 33924
rect 9398 33872 9404 33924
rect 9456 33872 9462 33924
rect 10134 33872 10140 33924
rect 10192 33872 10198 33924
rect 11054 33872 11060 33924
rect 11112 33872 11118 33924
rect 11146 33872 11152 33924
rect 11204 33912 11210 33924
rect 11517 33915 11575 33921
rect 11517 33912 11529 33915
rect 11204 33884 11529 33912
rect 11204 33872 11210 33884
rect 11517 33881 11529 33884
rect 11563 33881 11575 33915
rect 12176 33912 12204 34011
rect 11517 33875 11575 33881
rect 11624 33884 12204 33912
rect 4157 33847 4215 33853
rect 4157 33844 4169 33847
rect 4120 33816 4169 33844
rect 4120 33804 4126 33816
rect 4157 33813 4169 33816
rect 4203 33813 4215 33847
rect 4157 33807 4215 33813
rect 5629 33847 5687 33853
rect 5629 33813 5641 33847
rect 5675 33813 5687 33847
rect 5629 33807 5687 33813
rect 7374 33804 7380 33856
rect 7432 33804 7438 33856
rect 7561 33847 7619 33853
rect 7561 33813 7573 33847
rect 7607 33844 7619 33847
rect 7742 33844 7748 33856
rect 7607 33816 7748 33844
rect 7607 33813 7619 33816
rect 7561 33807 7619 33813
rect 7742 33804 7748 33816
rect 7800 33804 7806 33856
rect 9125 33847 9183 33853
rect 9125 33813 9137 33847
rect 9171 33844 9183 33847
rect 9858 33844 9864 33856
rect 9171 33816 9864 33844
rect 9171 33813 9183 33816
rect 9125 33807 9183 33813
rect 9858 33804 9864 33816
rect 9916 33804 9922 33856
rect 11422 33804 11428 33856
rect 11480 33844 11486 33856
rect 11624 33844 11652 33884
rect 11480 33816 11652 33844
rect 11480 33804 11486 33816
rect 11698 33804 11704 33856
rect 11756 33804 11762 33856
rect 11790 33804 11796 33856
rect 11848 33844 11854 33856
rect 12069 33847 12127 33853
rect 12069 33844 12081 33847
rect 11848 33816 12081 33844
rect 11848 33804 11854 33816
rect 12069 33813 12081 33816
rect 12115 33813 12127 33847
rect 12069 33807 12127 33813
rect 552 33754 12604 33776
rect 552 33702 3662 33754
rect 3714 33702 3726 33754
rect 3778 33702 3790 33754
rect 3842 33702 3854 33754
rect 3906 33702 3918 33754
rect 3970 33702 10062 33754
rect 10114 33702 10126 33754
rect 10178 33702 10190 33754
rect 10242 33702 10254 33754
rect 10306 33702 10318 33754
rect 10370 33702 12604 33754
rect 552 33680 12604 33702
rect 845 33643 903 33649
rect 845 33640 857 33643
rect 492 33612 857 33640
rect 845 33609 857 33612
rect 891 33609 903 33643
rect 845 33603 903 33609
rect 2038 33600 2044 33652
rect 2096 33640 2102 33652
rect 2866 33640 2872 33652
rect 2096 33612 2872 33640
rect 2096 33600 2102 33612
rect 2866 33600 2872 33612
rect 2924 33600 2930 33652
rect 3605 33643 3663 33649
rect 3605 33609 3617 33643
rect 3651 33640 3663 33643
rect 4062 33640 4068 33652
rect 3651 33612 4068 33640
rect 3651 33609 3663 33612
rect 3605 33603 3663 33609
rect 4062 33600 4068 33612
rect 4120 33600 4126 33652
rect 5810 33600 5816 33652
rect 5868 33640 5874 33652
rect 6365 33643 6423 33649
rect 6365 33640 6377 33643
rect 5868 33612 6377 33640
rect 5868 33600 5874 33612
rect 6365 33609 6377 33612
rect 6411 33609 6423 33643
rect 7926 33640 7932 33652
rect 6365 33603 6423 33609
rect 7208 33612 7932 33640
rect 5169 33575 5227 33581
rect 5169 33541 5181 33575
rect 5215 33572 5227 33575
rect 6638 33572 6644 33584
rect 5215 33544 6644 33572
rect 5215 33541 5227 33544
rect 5169 33535 5227 33541
rect 6638 33532 6644 33544
rect 6696 33532 6702 33584
rect 2222 33464 2228 33516
rect 2280 33464 2286 33516
rect 2498 33464 2504 33516
rect 2556 33464 2562 33516
rect 3421 33507 3479 33513
rect 3421 33473 3433 33507
rect 3467 33473 3479 33507
rect 3421 33467 3479 33473
rect 2314 33396 2320 33448
rect 2372 33436 2378 33448
rect 2685 33439 2743 33445
rect 2685 33436 2697 33439
rect 2372 33408 2697 33436
rect 2372 33396 2378 33408
rect 2685 33405 2697 33408
rect 2731 33436 2743 33439
rect 3050 33436 3056 33448
rect 2731 33408 3056 33436
rect 2731 33405 2743 33408
rect 2685 33399 2743 33405
rect 3050 33396 3056 33408
rect 3108 33396 3114 33448
rect 1946 33328 1952 33380
rect 2004 33377 2010 33380
rect 2004 33368 2016 33377
rect 3142 33368 3148 33380
rect 2004 33340 2049 33368
rect 2148 33340 3148 33368
rect 2004 33331 2016 33340
rect 2004 33328 2010 33331
rect 1486 33260 1492 33312
rect 1544 33300 1550 33312
rect 2148 33300 2176 33340
rect 3142 33328 3148 33340
rect 3200 33368 3206 33380
rect 3436 33368 3464 33467
rect 3510 33464 3516 33516
rect 3568 33504 3574 33516
rect 3789 33507 3847 33513
rect 3789 33504 3801 33507
rect 3568 33476 3801 33504
rect 3568 33464 3574 33476
rect 3789 33473 3801 33476
rect 3835 33473 3847 33507
rect 3789 33467 3847 33473
rect 5442 33464 5448 33516
rect 5500 33464 5506 33516
rect 5721 33507 5779 33513
rect 5721 33473 5733 33507
rect 5767 33504 5779 33507
rect 5994 33504 6000 33516
rect 5767 33476 6000 33504
rect 5767 33473 5779 33476
rect 5721 33467 5779 33473
rect 3694 33396 3700 33448
rect 3752 33396 3758 33448
rect 4056 33439 4114 33445
rect 4056 33405 4068 33439
rect 4102 33436 4114 33439
rect 5258 33436 5264 33448
rect 4102 33408 5264 33436
rect 4102 33405 4114 33408
rect 4056 33399 4114 33405
rect 5258 33396 5264 33408
rect 5316 33396 5322 33448
rect 4154 33368 4160 33380
rect 3200 33340 4160 33368
rect 3200 33328 3206 33340
rect 4154 33328 4160 33340
rect 4212 33328 4218 33380
rect 5736 33368 5764 33467
rect 5994 33464 6000 33476
rect 6052 33464 6058 33516
rect 6270 33464 6276 33516
rect 6328 33504 6334 33516
rect 7098 33504 7104 33516
rect 6328 33476 7104 33504
rect 6328 33464 6334 33476
rect 7098 33464 7104 33476
rect 7156 33464 7162 33516
rect 6362 33396 6368 33448
rect 6420 33436 6426 33448
rect 6549 33439 6607 33445
rect 6549 33436 6561 33439
rect 6420 33408 6561 33436
rect 6420 33396 6426 33408
rect 6549 33405 6561 33408
rect 6595 33405 6607 33439
rect 6549 33399 6607 33405
rect 5276 33340 5764 33368
rect 6564 33368 6592 33399
rect 6638 33396 6644 33448
rect 6696 33436 6702 33448
rect 6733 33439 6791 33445
rect 6733 33436 6745 33439
rect 6696 33408 6745 33436
rect 6696 33396 6702 33408
rect 6733 33405 6745 33408
rect 6779 33405 6791 33439
rect 6733 33399 6791 33405
rect 6825 33439 6883 33445
rect 6825 33405 6837 33439
rect 6871 33436 6883 33439
rect 7208 33436 7236 33612
rect 7926 33600 7932 33612
rect 7984 33600 7990 33652
rect 10134 33640 10140 33652
rect 8128 33612 10140 33640
rect 7469 33575 7527 33581
rect 7469 33541 7481 33575
rect 7515 33572 7527 33575
rect 8128 33572 8156 33612
rect 10134 33600 10140 33612
rect 10192 33600 10198 33652
rect 11882 33600 11888 33652
rect 11940 33600 11946 33652
rect 7515 33544 8156 33572
rect 8205 33575 8263 33581
rect 7515 33541 7527 33544
rect 7469 33535 7527 33541
rect 8205 33541 8217 33575
rect 8251 33572 8263 33575
rect 11977 33575 12035 33581
rect 8251 33544 8800 33572
rect 8251 33541 8263 33544
rect 8205 33535 8263 33541
rect 7484 33476 8609 33504
rect 7484 33445 7512 33476
rect 6871 33408 7236 33436
rect 7285 33439 7343 33445
rect 6871 33405 6883 33408
rect 6825 33399 6883 33405
rect 6917 33371 6975 33377
rect 6917 33368 6929 33371
rect 6564 33340 6929 33368
rect 5276 33312 5304 33340
rect 6917 33337 6929 33340
rect 6963 33337 6975 33371
rect 6917 33331 6975 33337
rect 1544 33272 2176 33300
rect 1544 33260 1550 33272
rect 2590 33260 2596 33312
rect 2648 33260 2654 33312
rect 3050 33260 3056 33312
rect 3108 33260 3114 33312
rect 3421 33303 3479 33309
rect 3421 33269 3433 33303
rect 3467 33300 3479 33303
rect 4246 33300 4252 33312
rect 3467 33272 4252 33300
rect 3467 33269 3479 33272
rect 3421 33263 3479 33269
rect 4246 33260 4252 33272
rect 4304 33260 4310 33312
rect 5258 33260 5264 33312
rect 5316 33260 5322 33312
rect 5350 33260 5356 33312
rect 5408 33300 5414 33312
rect 7024 33300 7052 33408
rect 7285 33405 7297 33439
rect 7331 33436 7343 33439
rect 7469 33439 7527 33445
rect 7331 33408 7420 33436
rect 7331 33405 7343 33408
rect 7285 33399 7343 33405
rect 7101 33371 7159 33377
rect 7101 33337 7113 33371
rect 7147 33337 7159 33371
rect 7392 33368 7420 33408
rect 7469 33405 7481 33439
rect 7515 33405 7527 33439
rect 7469 33399 7527 33405
rect 7650 33396 7656 33448
rect 7708 33396 7714 33448
rect 7926 33396 7932 33448
rect 7984 33396 7990 33448
rect 8386 33436 8392 33448
rect 8128 33408 8392 33436
rect 7668 33368 7696 33396
rect 7392 33340 7696 33368
rect 7745 33371 7803 33377
rect 7101 33331 7159 33337
rect 7745 33337 7757 33371
rect 7791 33368 7803 33371
rect 8128 33368 8156 33408
rect 8386 33396 8392 33408
rect 8444 33396 8450 33448
rect 7791 33340 8156 33368
rect 8205 33371 8263 33377
rect 7791 33337 7803 33340
rect 7745 33331 7803 33337
rect 8205 33337 8217 33371
rect 8251 33368 8263 33371
rect 8478 33368 8484 33380
rect 8251 33340 8484 33368
rect 8251 33337 8263 33340
rect 8205 33331 8263 33337
rect 5408 33272 7052 33300
rect 7116 33300 7144 33331
rect 8478 33328 8484 33340
rect 8536 33328 8542 33380
rect 8581 33368 8609 33476
rect 8772 33436 8800 33544
rect 11977 33541 11989 33575
rect 12023 33541 12035 33575
rect 11977 33535 12035 33541
rect 9502 33439 9560 33445
rect 9502 33436 9514 33439
rect 8772 33408 9514 33436
rect 9502 33405 9514 33408
rect 9548 33405 9560 33439
rect 9502 33399 9560 33405
rect 9769 33439 9827 33445
rect 9769 33405 9781 33439
rect 9815 33436 9827 33439
rect 10502 33436 10508 33448
rect 9815 33408 10508 33436
rect 9815 33405 9827 33408
rect 9769 33399 9827 33405
rect 10502 33396 10508 33408
rect 10560 33396 10566 33448
rect 10772 33439 10830 33445
rect 10772 33405 10784 33439
rect 10818 33436 10830 33439
rect 11992 33436 12020 33535
rect 10818 33408 12020 33436
rect 12253 33439 12311 33445
rect 10818 33405 10830 33408
rect 10772 33399 10830 33405
rect 12253 33405 12265 33439
rect 12299 33436 12311 33439
rect 12526 33436 12532 33448
rect 12299 33408 12532 33436
rect 12299 33405 12311 33408
rect 12253 33399 12311 33405
rect 12526 33396 12532 33408
rect 12584 33396 12590 33448
rect 9674 33368 9680 33380
rect 8581 33340 9680 33368
rect 9674 33328 9680 33340
rect 9732 33328 9738 33380
rect 9950 33328 9956 33380
rect 10008 33328 10014 33380
rect 10226 33328 10232 33380
rect 10284 33368 10290 33380
rect 10321 33371 10379 33377
rect 10321 33368 10333 33371
rect 10284 33340 10333 33368
rect 10284 33328 10290 33340
rect 10321 33337 10333 33340
rect 10367 33337 10379 33371
rect 10321 33331 10379 33337
rect 11974 33328 11980 33380
rect 12032 33328 12038 33380
rect 7374 33300 7380 33312
rect 7116 33272 7380 33300
rect 5408 33260 5414 33272
rect 7374 33260 7380 33272
rect 7432 33260 7438 33312
rect 7558 33260 7564 33312
rect 7616 33300 7622 33312
rect 7653 33303 7711 33309
rect 7653 33300 7665 33303
rect 7616 33272 7665 33300
rect 7616 33260 7622 33272
rect 7653 33269 7665 33272
rect 7699 33300 7711 33303
rect 8021 33303 8079 33309
rect 8021 33300 8033 33303
rect 7699 33272 8033 33300
rect 7699 33269 7711 33272
rect 7653 33263 7711 33269
rect 8021 33269 8033 33272
rect 8067 33269 8079 33303
rect 8021 33263 8079 33269
rect 8389 33303 8447 33309
rect 8389 33269 8401 33303
rect 8435 33300 8447 33303
rect 8662 33300 8668 33312
rect 8435 33272 8668 33300
rect 8435 33269 8447 33272
rect 8389 33263 8447 33269
rect 8662 33260 8668 33272
rect 8720 33260 8726 33312
rect 12158 33260 12164 33312
rect 12216 33260 12222 33312
rect 552 33210 12604 33232
rect 552 33158 4322 33210
rect 4374 33158 4386 33210
rect 4438 33158 4450 33210
rect 4502 33158 4514 33210
rect 4566 33158 4578 33210
rect 4630 33158 10722 33210
rect 10774 33158 10786 33210
rect 10838 33158 10850 33210
rect 10902 33158 10914 33210
rect 10966 33158 10978 33210
rect 11030 33158 12604 33210
rect 552 33136 12604 33158
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 4157 33099 4215 33105
rect 4157 33096 4169 33099
rect 2924 33068 4169 33096
rect 2924 33056 2930 33068
rect 4157 33065 4169 33068
rect 4203 33065 4215 33099
rect 4157 33059 4215 33065
rect 4890 33056 4896 33108
rect 4948 33056 4954 33108
rect 6454 33056 6460 33108
rect 6512 33096 6518 33108
rect 6733 33099 6791 33105
rect 6733 33096 6745 33099
rect 6512 33068 6745 33096
rect 6512 33056 6518 33068
rect 6733 33065 6745 33068
rect 6779 33096 6791 33099
rect 7006 33096 7012 33108
rect 6779 33068 7012 33096
rect 6779 33065 6791 33068
rect 6733 33059 6791 33065
rect 7006 33056 7012 33068
rect 7064 33056 7070 33108
rect 7098 33056 7104 33108
rect 7156 33096 7162 33108
rect 7156 33068 7236 33096
rect 7156 33056 7162 33068
rect 1118 32988 1124 33040
rect 1176 32988 1182 33040
rect 2222 32988 2228 33040
rect 2280 33028 2286 33040
rect 2952 33031 3010 33037
rect 2280 33000 2636 33028
rect 2280 32988 2286 33000
rect 845 32963 903 32969
rect 845 32929 857 32963
rect 891 32960 903 32963
rect 1210 32960 1216 32972
rect 891 32932 1216 32960
rect 891 32929 903 32932
rect 845 32923 903 32929
rect 1210 32920 1216 32932
rect 1268 32920 1274 32972
rect 2337 32963 2395 32969
rect 2337 32929 2349 32963
rect 2383 32960 2395 32963
rect 2498 32960 2504 32972
rect 2383 32932 2504 32960
rect 2383 32929 2395 32932
rect 2337 32923 2395 32929
rect 2498 32920 2504 32932
rect 2556 32920 2562 32972
rect 2608 32969 2636 33000
rect 2952 32997 2964 33031
rect 2998 33028 3010 33031
rect 3050 33028 3056 33040
rect 2998 33000 3056 33028
rect 2998 32997 3010 33000
rect 2952 32991 3010 32997
rect 3050 32988 3056 33000
rect 3108 32988 3114 33040
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 5537 33031 5595 33037
rect 5537 33028 5549 33031
rect 3476 33000 5549 33028
rect 3476 32988 3482 33000
rect 5537 32997 5549 33000
rect 5583 32997 5595 33031
rect 7208 33028 7236 33068
rect 7282 33056 7288 33108
rect 7340 33056 7346 33108
rect 7926 33056 7932 33108
rect 7984 33096 7990 33108
rect 8021 33099 8079 33105
rect 8021 33096 8033 33099
rect 7984 33068 8033 33096
rect 7984 33056 7990 33068
rect 8021 33065 8033 33068
rect 8067 33065 8079 33099
rect 8021 33059 8079 33065
rect 8478 33056 8484 33108
rect 8536 33056 8542 33108
rect 9306 33056 9312 33108
rect 9364 33096 9370 33108
rect 9766 33096 9772 33108
rect 9364 33068 9772 33096
rect 9364 33056 9370 33068
rect 9766 33056 9772 33068
rect 9824 33056 9830 33108
rect 10502 33056 10508 33108
rect 10560 33096 10566 33108
rect 10560 33068 10824 33096
rect 10560 33056 10566 33068
rect 5537 32991 5595 32997
rect 5736 33000 7144 33028
rect 7208 33000 7512 33028
rect 2593 32963 2651 32969
rect 2593 32929 2605 32963
rect 2639 32929 2651 32963
rect 2593 32923 2651 32929
rect 4890 32920 4896 32972
rect 4948 32920 4954 32972
rect 5077 32963 5135 32969
rect 5077 32929 5089 32963
rect 5123 32929 5135 32963
rect 5077 32923 5135 32929
rect 1121 32895 1179 32901
rect 1121 32861 1133 32895
rect 1167 32892 1179 32895
rect 1486 32892 1492 32904
rect 1167 32864 1492 32892
rect 1167 32861 1179 32864
rect 1121 32855 1179 32861
rect 1486 32852 1492 32864
rect 1544 32852 1550 32904
rect 2682 32852 2688 32904
rect 2740 32852 2746 32904
rect 4801 32895 4859 32901
rect 4801 32861 4813 32895
rect 4847 32892 4859 32895
rect 4982 32892 4988 32904
rect 4847 32864 4988 32892
rect 4847 32861 4859 32864
rect 4801 32855 4859 32861
rect 937 32827 995 32833
rect 937 32793 949 32827
rect 983 32824 995 32827
rect 983 32796 1716 32824
rect 983 32793 995 32796
rect 937 32787 995 32793
rect 1213 32759 1271 32765
rect 1213 32725 1225 32759
rect 1259 32756 1271 32759
rect 1486 32756 1492 32768
rect 1259 32728 1492 32756
rect 1259 32725 1271 32728
rect 1213 32719 1271 32725
rect 1486 32716 1492 32728
rect 1544 32716 1550 32768
rect 1688 32756 1716 32796
rect 3694 32784 3700 32836
rect 3752 32824 3758 32836
rect 4430 32824 4436 32836
rect 3752 32796 4436 32824
rect 3752 32784 3758 32796
rect 4430 32784 4436 32796
rect 4488 32784 4494 32836
rect 3418 32756 3424 32768
rect 1688 32728 3424 32756
rect 3418 32716 3424 32728
rect 3476 32716 3482 32768
rect 4065 32759 4123 32765
rect 4065 32725 4077 32759
rect 4111 32756 4123 32759
rect 4816 32756 4844 32855
rect 4982 32852 4988 32864
rect 5040 32852 5046 32904
rect 5092 32824 5120 32923
rect 5350 32920 5356 32972
rect 5408 32920 5414 32972
rect 5736 32960 5764 33000
rect 5460 32932 5764 32960
rect 5460 32904 5488 32932
rect 5810 32920 5816 32972
rect 5868 32920 5874 32972
rect 5951 32963 6009 32969
rect 5951 32929 5963 32963
rect 5997 32960 6009 32963
rect 6178 32960 6184 32972
rect 5997 32932 6184 32960
rect 5997 32929 6009 32932
rect 5951 32923 6009 32929
rect 6178 32920 6184 32932
rect 6236 32920 6242 32972
rect 6273 32963 6331 32969
rect 6273 32929 6285 32963
rect 6319 32960 6331 32963
rect 6454 32960 6460 32972
rect 6319 32932 6460 32960
rect 6319 32929 6331 32932
rect 6273 32923 6331 32929
rect 6454 32920 6460 32932
rect 6512 32920 6518 32972
rect 6638 32920 6644 32972
rect 6696 32920 6702 32972
rect 6822 32920 6828 32972
rect 6880 32920 6886 32972
rect 6914 32920 6920 32972
rect 6972 32960 6978 32972
rect 7009 32963 7067 32969
rect 7009 32960 7021 32963
rect 6972 32932 7021 32960
rect 6972 32920 6978 32932
rect 7009 32929 7021 32932
rect 7055 32929 7067 32963
rect 7116 32960 7144 33000
rect 7193 32963 7251 32969
rect 7193 32960 7205 32963
rect 7116 32932 7205 32960
rect 7009 32923 7067 32929
rect 7193 32929 7205 32932
rect 7239 32929 7251 32963
rect 7193 32923 7251 32929
rect 7282 32920 7288 32972
rect 7340 32960 7346 32972
rect 7484 32969 7512 33000
rect 7944 33000 9260 33028
rect 7944 32969 7972 33000
rect 7377 32963 7435 32969
rect 7377 32960 7389 32963
rect 7340 32932 7389 32960
rect 7340 32920 7346 32932
rect 7377 32929 7389 32932
rect 7423 32929 7435 32963
rect 7377 32923 7435 32929
rect 7469 32963 7527 32969
rect 7469 32929 7481 32963
rect 7515 32929 7527 32963
rect 7469 32923 7527 32929
rect 7561 32963 7619 32969
rect 7561 32929 7573 32963
rect 7607 32929 7619 32963
rect 7561 32923 7619 32929
rect 7929 32963 7987 32969
rect 7929 32929 7941 32963
rect 7975 32929 7987 32963
rect 7929 32923 7987 32929
rect 5169 32895 5227 32901
rect 5169 32861 5181 32895
rect 5215 32892 5227 32895
rect 5442 32892 5448 32904
rect 5215 32864 5448 32892
rect 5215 32861 5227 32864
rect 5169 32855 5227 32861
rect 5442 32852 5448 32864
rect 5500 32852 5506 32904
rect 5534 32852 5540 32904
rect 5592 32892 5598 32904
rect 7576 32892 7604 32923
rect 8110 32920 8116 32972
rect 8168 32920 8174 32972
rect 8205 32963 8263 32969
rect 8205 32929 8217 32963
rect 8251 32929 8263 32963
rect 8205 32923 8263 32929
rect 5592 32864 7604 32892
rect 5592 32852 5598 32864
rect 7650 32852 7656 32904
rect 7708 32892 7714 32904
rect 8220 32892 8248 32923
rect 8662 32920 8668 32972
rect 8720 32920 8726 32972
rect 8754 32920 8760 32972
rect 8812 32960 8818 32972
rect 9125 32963 9183 32969
rect 9125 32960 9137 32963
rect 8812 32932 9137 32960
rect 8812 32920 8818 32932
rect 9125 32929 9137 32932
rect 9171 32929 9183 32963
rect 9125 32923 9183 32929
rect 7708 32864 8248 32892
rect 8481 32895 8539 32901
rect 7708 32852 7714 32864
rect 8481 32861 8493 32895
rect 8527 32892 8539 32895
rect 8527 32864 9168 32892
rect 8527 32861 8539 32864
rect 8481 32855 8539 32861
rect 9140 32836 9168 32864
rect 5350 32824 5356 32836
rect 5092 32796 5356 32824
rect 5350 32784 5356 32796
rect 5408 32784 5414 32836
rect 6181 32827 6239 32833
rect 6181 32793 6193 32827
rect 6227 32824 6239 32827
rect 6457 32827 6515 32833
rect 6457 32824 6469 32827
rect 6227 32796 6469 32824
rect 6227 32793 6239 32796
rect 6181 32787 6239 32793
rect 6457 32793 6469 32796
rect 6503 32793 6515 32827
rect 6457 32787 6515 32793
rect 6914 32784 6920 32836
rect 6972 32824 6978 32836
rect 7466 32824 7472 32836
rect 6972 32796 7472 32824
rect 6972 32784 6978 32796
rect 7466 32784 7472 32796
rect 7524 32784 7530 32836
rect 7926 32784 7932 32836
rect 7984 32824 7990 32836
rect 8297 32827 8355 32833
rect 8297 32824 8309 32827
rect 7984 32796 8309 32824
rect 7984 32784 7990 32796
rect 8297 32793 8309 32796
rect 8343 32793 8355 32827
rect 8297 32787 8355 32793
rect 9122 32784 9128 32836
rect 9180 32784 9186 32836
rect 4111 32728 4844 32756
rect 4111 32725 4123 32728
rect 4065 32719 4123 32725
rect 6086 32716 6092 32768
rect 6144 32716 6150 32768
rect 6730 32716 6736 32768
rect 6788 32756 6794 32768
rect 7098 32756 7104 32768
rect 6788 32728 7104 32756
rect 6788 32716 6794 32728
rect 7098 32716 7104 32728
rect 7156 32756 7162 32768
rect 7745 32759 7803 32765
rect 7745 32756 7757 32759
rect 7156 32728 7757 32756
rect 7156 32716 7162 32728
rect 7745 32725 7757 32728
rect 7791 32725 7803 32759
rect 7745 32719 7803 32725
rect 8386 32716 8392 32768
rect 8444 32756 8450 32768
rect 8938 32756 8944 32768
rect 8444 32728 8944 32756
rect 8444 32716 8450 32728
rect 8938 32716 8944 32728
rect 8996 32716 9002 32768
rect 9232 32765 9260 33000
rect 9858 32988 9864 33040
rect 9916 33028 9922 33040
rect 10686 33028 10692 33040
rect 9916 33000 10692 33028
rect 9916 32988 9922 33000
rect 10686 32988 10692 33000
rect 10744 32988 10750 33040
rect 10796 33028 10824 33068
rect 10870 33056 10876 33108
rect 10928 33096 10934 33108
rect 11057 33099 11115 33105
rect 11057 33096 11069 33099
rect 10928 33068 11069 33096
rect 10928 33056 10934 33068
rect 11057 33065 11069 33068
rect 11103 33096 11115 33099
rect 12710 33096 12716 33108
rect 11103 33068 12716 33096
rect 11103 33065 11115 33068
rect 11057 33059 11115 33065
rect 12710 33056 12716 33068
rect 12768 33056 12774 33108
rect 12250 33028 12256 33040
rect 10796 33000 12256 33028
rect 9309 32963 9367 32969
rect 9309 32929 9321 32963
rect 9355 32960 9367 32963
rect 9582 32960 9588 32972
rect 9355 32932 9588 32960
rect 9355 32929 9367 32932
rect 9309 32923 9367 32929
rect 9582 32920 9588 32932
rect 9640 32920 9646 32972
rect 10796 32969 10824 33000
rect 12250 32988 12256 33000
rect 12308 32988 12314 33040
rect 10525 32963 10583 32969
rect 10525 32929 10537 32963
rect 10571 32960 10583 32963
rect 10781 32963 10839 32969
rect 10571 32932 10732 32960
rect 10571 32929 10583 32932
rect 10525 32923 10583 32929
rect 10704 32892 10732 32932
rect 10781 32929 10793 32963
rect 10827 32929 10839 32963
rect 10781 32923 10839 32929
rect 11241 32963 11299 32969
rect 11241 32929 11253 32963
rect 11287 32960 11299 32963
rect 11330 32960 11336 32972
rect 11287 32932 11336 32960
rect 11287 32929 11299 32932
rect 11241 32923 11299 32929
rect 11330 32920 11336 32932
rect 11388 32920 11394 32972
rect 11701 32963 11759 32969
rect 11701 32929 11713 32963
rect 11747 32960 11759 32963
rect 11882 32960 11888 32972
rect 11747 32932 11888 32960
rect 11747 32929 11759 32932
rect 11701 32923 11759 32929
rect 11882 32920 11888 32932
rect 11940 32920 11946 32972
rect 11146 32892 11152 32904
rect 10704 32864 11152 32892
rect 11146 32852 11152 32864
rect 11204 32852 11210 32904
rect 11425 32895 11483 32901
rect 11425 32861 11437 32895
rect 11471 32861 11483 32895
rect 11425 32855 11483 32861
rect 11440 32824 11468 32855
rect 12158 32852 12164 32904
rect 12216 32892 12222 32904
rect 12253 32895 12311 32901
rect 12253 32892 12265 32895
rect 12216 32864 12265 32892
rect 12216 32852 12222 32864
rect 12253 32861 12265 32864
rect 12299 32861 12311 32895
rect 12253 32855 12311 32861
rect 11698 32824 11704 32836
rect 11440 32796 11704 32824
rect 11698 32784 11704 32796
rect 11756 32784 11762 32836
rect 9217 32759 9275 32765
rect 9217 32725 9229 32759
rect 9263 32756 9275 32759
rect 9306 32756 9312 32768
rect 9263 32728 9312 32756
rect 9263 32725 9275 32728
rect 9217 32719 9275 32725
rect 9306 32716 9312 32728
rect 9364 32716 9370 32768
rect 9401 32759 9459 32765
rect 9401 32725 9413 32759
rect 9447 32756 9459 32759
rect 9490 32756 9496 32768
rect 9447 32728 9496 32756
rect 9447 32725 9459 32728
rect 9401 32719 9459 32725
rect 9490 32716 9496 32728
rect 9548 32716 9554 32768
rect 10134 32716 10140 32768
rect 10192 32756 10198 32768
rect 11330 32756 11336 32768
rect 10192 32728 11336 32756
rect 10192 32716 10198 32728
rect 11330 32716 11336 32728
rect 11388 32716 11394 32768
rect 552 32666 12604 32688
rect 552 32614 3662 32666
rect 3714 32614 3726 32666
rect 3778 32614 3790 32666
rect 3842 32614 3854 32666
rect 3906 32614 3918 32666
rect 3970 32614 10062 32666
rect 10114 32614 10126 32666
rect 10178 32614 10190 32666
rect 10242 32614 10254 32666
rect 10306 32614 10318 32666
rect 10370 32614 12604 32666
rect 552 32592 12604 32614
rect 1118 32512 1124 32564
rect 1176 32552 1182 32564
rect 2130 32552 2136 32564
rect 1176 32524 2136 32552
rect 1176 32512 1182 32524
rect 2130 32512 2136 32524
rect 2188 32512 2194 32564
rect 2498 32512 2504 32564
rect 2556 32552 2562 32564
rect 3237 32555 3295 32561
rect 3237 32552 3249 32555
rect 2556 32524 3249 32552
rect 2556 32512 2562 32524
rect 3237 32521 3249 32524
rect 3283 32521 3295 32555
rect 4890 32552 4896 32564
rect 3237 32515 3295 32521
rect 3896 32524 4896 32552
rect 1486 32444 1492 32496
rect 1544 32444 1550 32496
rect 3896 32416 3924 32524
rect 4890 32512 4896 32524
rect 4948 32512 4954 32564
rect 5534 32552 5540 32564
rect 5184 32524 5540 32552
rect 5184 32493 5212 32524
rect 5534 32512 5540 32524
rect 5592 32512 5598 32564
rect 5905 32555 5963 32561
rect 5905 32521 5917 32555
rect 5951 32552 5963 32555
rect 6086 32552 6092 32564
rect 5951 32524 6092 32552
rect 5951 32521 5963 32524
rect 5905 32515 5963 32521
rect 6086 32512 6092 32524
rect 6144 32512 6150 32564
rect 6638 32512 6644 32564
rect 6696 32512 6702 32564
rect 6733 32555 6791 32561
rect 6733 32521 6745 32555
rect 6779 32552 6791 32555
rect 6822 32552 6828 32564
rect 6779 32524 6828 32552
rect 6779 32521 6791 32524
rect 6733 32515 6791 32521
rect 6822 32512 6828 32524
rect 6880 32512 6886 32564
rect 6917 32555 6975 32561
rect 6917 32521 6929 32555
rect 6963 32552 6975 32555
rect 7098 32552 7104 32564
rect 6963 32524 7104 32552
rect 6963 32521 6975 32524
rect 6917 32515 6975 32521
rect 7098 32512 7104 32524
rect 7156 32512 7162 32564
rect 7926 32512 7932 32564
rect 7984 32552 7990 32564
rect 9217 32555 9275 32561
rect 7984 32524 8892 32552
rect 7984 32512 7990 32524
rect 4065 32487 4123 32493
rect 4065 32453 4077 32487
rect 4111 32484 4123 32487
rect 5169 32487 5227 32493
rect 4111 32456 4936 32484
rect 4111 32453 4123 32456
rect 4065 32447 4123 32453
rect 952 32388 3924 32416
rect 952 32357 980 32388
rect 4246 32376 4252 32428
rect 4304 32416 4310 32428
rect 4304 32388 4660 32416
rect 4304 32376 4310 32388
rect 937 32351 995 32357
rect 937 32317 949 32351
rect 983 32317 995 32351
rect 937 32311 995 32317
rect 1210 32308 1216 32360
rect 1268 32348 1274 32360
rect 2685 32351 2743 32357
rect 2685 32348 2697 32351
rect 1268 32320 2697 32348
rect 1268 32308 1274 32320
rect 2685 32317 2697 32320
rect 2731 32317 2743 32351
rect 2685 32311 2743 32317
rect 2961 32351 3019 32357
rect 2961 32317 2973 32351
rect 3007 32348 3019 32351
rect 3326 32348 3332 32360
rect 3007 32320 3332 32348
rect 3007 32317 3019 32320
rect 2961 32311 3019 32317
rect 3326 32308 3332 32320
rect 3384 32348 3390 32360
rect 3421 32351 3479 32357
rect 3421 32348 3433 32351
rect 3384 32320 3433 32348
rect 3384 32308 3390 32320
rect 3421 32317 3433 32320
rect 3467 32317 3479 32351
rect 3421 32311 3479 32317
rect 3513 32351 3571 32357
rect 3513 32317 3525 32351
rect 3559 32317 3571 32351
rect 3513 32311 3571 32317
rect 1765 32283 1823 32289
rect 1765 32280 1777 32283
rect 1412 32252 1777 32280
rect 1412 32224 1440 32252
rect 1765 32249 1777 32252
rect 1811 32249 1823 32283
rect 1765 32243 1823 32249
rect 2225 32283 2283 32289
rect 2225 32249 2237 32283
rect 2271 32249 2283 32283
rect 2225 32243 2283 32249
rect 1026 32172 1032 32224
rect 1084 32172 1090 32224
rect 1394 32172 1400 32224
rect 1452 32172 1458 32224
rect 1673 32215 1731 32221
rect 1673 32181 1685 32215
rect 1719 32212 1731 32215
rect 2240 32212 2268 32243
rect 2406 32240 2412 32292
rect 2464 32280 2470 32292
rect 2593 32283 2651 32289
rect 2593 32280 2605 32283
rect 2464 32252 2605 32280
rect 2464 32240 2470 32252
rect 2593 32249 2605 32252
rect 2639 32280 2651 32283
rect 3528 32280 3556 32311
rect 3602 32308 3608 32360
rect 3660 32348 3666 32360
rect 3881 32351 3939 32357
rect 3881 32348 3893 32351
rect 3660 32320 3893 32348
rect 3660 32308 3666 32320
rect 3881 32317 3893 32320
rect 3927 32317 3939 32351
rect 3881 32311 3939 32317
rect 4062 32308 4068 32360
rect 4120 32348 4126 32360
rect 4341 32351 4399 32357
rect 4341 32348 4353 32351
rect 4120 32320 4353 32348
rect 4120 32308 4126 32320
rect 4341 32317 4353 32320
rect 4387 32317 4399 32351
rect 4341 32311 4399 32317
rect 4430 32308 4436 32360
rect 4488 32308 4494 32360
rect 4632 32357 4660 32388
rect 4617 32351 4675 32357
rect 4617 32317 4629 32351
rect 4663 32317 4675 32351
rect 4617 32311 4675 32317
rect 4801 32351 4859 32357
rect 4801 32317 4813 32351
rect 4847 32317 4859 32351
rect 4908 32348 4936 32456
rect 5169 32453 5181 32487
rect 5215 32453 5227 32487
rect 5169 32447 5227 32453
rect 5261 32487 5319 32493
rect 5261 32453 5273 32487
rect 5307 32484 5319 32487
rect 5350 32484 5356 32496
rect 5307 32456 5356 32484
rect 5307 32453 5319 32456
rect 5261 32447 5319 32453
rect 5350 32444 5356 32456
rect 5408 32484 5414 32496
rect 5408 32456 6040 32484
rect 5408 32444 5414 32456
rect 4982 32376 4988 32428
rect 5040 32416 5046 32428
rect 6012 32425 6040 32456
rect 6270 32444 6276 32496
rect 6328 32444 6334 32496
rect 7006 32444 7012 32496
rect 7064 32484 7070 32496
rect 7193 32487 7251 32493
rect 7193 32484 7205 32487
rect 7064 32456 7205 32484
rect 7064 32444 7070 32456
rect 7193 32453 7205 32456
rect 7239 32453 7251 32487
rect 8294 32484 8300 32496
rect 7193 32447 7251 32453
rect 8036 32456 8300 32484
rect 5997 32419 6055 32425
rect 5040 32388 5396 32416
rect 5040 32376 5046 32388
rect 5368 32357 5396 32388
rect 5997 32385 6009 32419
rect 6043 32416 6055 32419
rect 6178 32416 6184 32428
rect 6043 32388 6184 32416
rect 6043 32385 6055 32388
rect 5997 32379 6055 32385
rect 6178 32376 6184 32388
rect 6236 32376 6242 32428
rect 6288 32416 6316 32444
rect 6365 32419 6423 32425
rect 6365 32416 6377 32419
rect 6288 32388 6377 32416
rect 6365 32385 6377 32388
rect 6411 32385 6423 32419
rect 6365 32379 6423 32385
rect 5077 32351 5135 32357
rect 5077 32348 5089 32351
rect 4908 32320 5089 32348
rect 4801 32311 4859 32317
rect 5077 32317 5089 32320
rect 5123 32317 5135 32351
rect 5077 32311 5135 32317
rect 5353 32351 5411 32357
rect 5353 32317 5365 32351
rect 5399 32317 5411 32351
rect 5353 32311 5411 32317
rect 6089 32351 6147 32357
rect 6089 32317 6101 32351
rect 6135 32348 6147 32351
rect 6270 32348 6276 32360
rect 6135 32320 6276 32348
rect 6135 32317 6147 32320
rect 6089 32311 6147 32317
rect 4816 32280 4844 32311
rect 2639 32252 3556 32280
rect 4172 32252 4844 32280
rect 5092 32280 5120 32311
rect 6270 32308 6276 32320
rect 6328 32308 6334 32360
rect 5537 32283 5595 32289
rect 5537 32280 5549 32283
rect 5092 32252 5549 32280
rect 2639 32249 2651 32252
rect 2593 32243 2651 32249
rect 4172 32224 4200 32252
rect 5537 32249 5549 32252
rect 5583 32249 5595 32283
rect 5537 32243 5595 32249
rect 5721 32283 5779 32289
rect 5721 32249 5733 32283
rect 5767 32280 5779 32283
rect 6178 32280 6184 32292
rect 5767 32252 6184 32280
rect 5767 32249 5779 32252
rect 5721 32243 5779 32249
rect 1719 32184 2268 32212
rect 1719 32181 1731 32184
rect 1673 32175 1731 32181
rect 3234 32172 3240 32224
rect 3292 32212 3298 32224
rect 3786 32212 3792 32224
rect 3292 32184 3792 32212
rect 3292 32172 3298 32184
rect 3786 32172 3792 32184
rect 3844 32172 3850 32224
rect 4154 32172 4160 32224
rect 4212 32172 4218 32224
rect 4246 32172 4252 32224
rect 4304 32212 4310 32224
rect 4709 32215 4767 32221
rect 4709 32212 4721 32215
rect 4304 32184 4721 32212
rect 4304 32172 4310 32184
rect 4709 32181 4721 32184
rect 4755 32181 4767 32215
rect 4709 32175 4767 32181
rect 4893 32215 4951 32221
rect 4893 32181 4905 32215
rect 4939 32212 4951 32215
rect 5074 32212 5080 32224
rect 4939 32184 5080 32212
rect 4939 32181 4951 32184
rect 4893 32175 4951 32181
rect 5074 32172 5080 32184
rect 5132 32172 5138 32224
rect 5552 32212 5580 32243
rect 6178 32240 6184 32252
rect 6236 32280 6242 32292
rect 6380 32280 6408 32379
rect 6454 32376 6460 32428
rect 6512 32416 6518 32428
rect 6512 32388 7696 32416
rect 6512 32376 6518 32388
rect 6236 32252 6408 32280
rect 6748 32280 6776 32388
rect 6822 32308 6828 32360
rect 6880 32348 6886 32360
rect 7377 32351 7435 32357
rect 7377 32348 7389 32351
rect 6880 32320 7389 32348
rect 6880 32308 6886 32320
rect 7377 32317 7389 32320
rect 7423 32317 7435 32351
rect 7377 32311 7435 32317
rect 7558 32308 7564 32360
rect 7616 32308 7622 32360
rect 7668 32348 7696 32388
rect 7834 32376 7840 32428
rect 7892 32376 7898 32428
rect 8036 32425 8064 32456
rect 8294 32444 8300 32456
rect 8352 32484 8358 32496
rect 8570 32484 8576 32496
rect 8352 32456 8576 32484
rect 8352 32444 8358 32456
rect 8570 32444 8576 32456
rect 8628 32484 8634 32496
rect 8665 32487 8723 32493
rect 8665 32484 8677 32487
rect 8628 32456 8677 32484
rect 8628 32444 8634 32456
rect 8665 32453 8677 32456
rect 8711 32484 8723 32487
rect 8754 32484 8760 32496
rect 8711 32456 8760 32484
rect 8711 32453 8723 32456
rect 8665 32447 8723 32453
rect 8754 32444 8760 32456
rect 8812 32444 8818 32496
rect 8864 32493 8892 32524
rect 9217 32521 9229 32555
rect 9263 32552 9275 32555
rect 9493 32555 9551 32561
rect 9493 32552 9505 32555
rect 9263 32524 9505 32552
rect 9263 32521 9275 32524
rect 9217 32515 9275 32521
rect 9493 32521 9505 32524
rect 9539 32521 9551 32555
rect 9493 32515 9551 32521
rect 9582 32512 9588 32564
rect 9640 32552 9646 32564
rect 10321 32555 10379 32561
rect 10321 32552 10333 32555
rect 9640 32524 10333 32552
rect 9640 32512 9646 32524
rect 10321 32521 10333 32524
rect 10367 32552 10379 32555
rect 10594 32552 10600 32564
rect 10367 32524 10600 32552
rect 10367 32521 10379 32524
rect 10321 32515 10379 32521
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 8849 32487 8907 32493
rect 8849 32453 8861 32487
rect 8895 32453 8907 32487
rect 8849 32447 8907 32453
rect 9398 32444 9404 32496
rect 9456 32444 9462 32496
rect 8021 32419 8079 32425
rect 8021 32385 8033 32419
rect 8067 32385 8079 32419
rect 8021 32379 8079 32385
rect 8113 32419 8171 32425
rect 8113 32385 8125 32419
rect 8159 32416 8171 32419
rect 8159 32388 8609 32416
rect 8159 32385 8171 32388
rect 8113 32379 8171 32385
rect 7929 32351 7987 32357
rect 7929 32348 7941 32351
rect 7668 32320 7941 32348
rect 7852 32292 7880 32320
rect 7929 32317 7941 32320
rect 7975 32317 7987 32351
rect 7929 32311 7987 32317
rect 7006 32280 7012 32292
rect 6748 32252 7012 32280
rect 6236 32240 6242 32252
rect 7006 32240 7012 32252
rect 7064 32240 7070 32292
rect 7101 32283 7159 32289
rect 7101 32249 7113 32283
rect 7147 32280 7159 32283
rect 7147 32252 7770 32280
rect 7147 32249 7159 32252
rect 7101 32243 7159 32249
rect 5902 32212 5908 32224
rect 5552 32184 5908 32212
rect 5902 32172 5908 32184
rect 5960 32212 5966 32224
rect 6273 32215 6331 32221
rect 6273 32212 6285 32215
rect 5960 32184 6285 32212
rect 5960 32172 5966 32184
rect 6273 32181 6285 32184
rect 6319 32212 6331 32215
rect 6546 32212 6552 32224
rect 6319 32184 6552 32212
rect 6319 32181 6331 32184
rect 6273 32175 6331 32181
rect 6546 32172 6552 32184
rect 6604 32172 6610 32224
rect 6901 32215 6959 32221
rect 6901 32181 6913 32215
rect 6947 32212 6959 32215
rect 7282 32212 7288 32224
rect 6947 32184 7288 32212
rect 6947 32181 6959 32184
rect 6901 32175 6959 32181
rect 7282 32172 7288 32184
rect 7340 32172 7346 32224
rect 7466 32172 7472 32224
rect 7524 32212 7530 32224
rect 7653 32215 7711 32221
rect 7653 32212 7665 32215
rect 7524 32184 7665 32212
rect 7524 32172 7530 32184
rect 7653 32181 7665 32184
rect 7699 32181 7711 32215
rect 7742 32212 7770 32252
rect 7834 32240 7840 32292
rect 7892 32240 7898 32292
rect 7926 32212 7932 32224
rect 7742 32184 7932 32212
rect 7653 32175 7711 32181
rect 7926 32172 7932 32184
rect 7984 32212 7990 32224
rect 8128 32212 8156 32379
rect 8481 32351 8539 32357
rect 8481 32317 8493 32351
rect 8527 32317 8539 32351
rect 8581 32348 8609 32388
rect 8938 32376 8944 32428
rect 8996 32416 9002 32428
rect 9600 32416 9628 32512
rect 9674 32444 9680 32496
rect 9732 32484 9738 32496
rect 10226 32484 10232 32496
rect 9732 32456 10232 32484
rect 9732 32444 9738 32456
rect 10226 32444 10232 32456
rect 10284 32444 10290 32496
rect 9769 32419 9827 32425
rect 9769 32416 9781 32419
rect 8996 32388 9781 32416
rect 8996 32376 9002 32388
rect 9769 32385 9781 32388
rect 9815 32385 9827 32419
rect 9769 32379 9827 32385
rect 9858 32376 9864 32428
rect 9916 32376 9922 32428
rect 9953 32419 10011 32425
rect 9953 32385 9965 32419
rect 9999 32416 10011 32419
rect 11790 32416 11796 32428
rect 9999 32388 11796 32416
rect 9999 32385 10011 32388
rect 9953 32379 10011 32385
rect 8581 32320 9343 32348
rect 8481 32311 8539 32317
rect 7984 32184 8156 32212
rect 8496 32212 8524 32311
rect 9122 32240 9128 32292
rect 9180 32280 9186 32292
rect 9217 32283 9275 32289
rect 9217 32280 9229 32283
rect 9180 32252 9229 32280
rect 9180 32240 9186 32252
rect 9217 32249 9229 32252
rect 9263 32249 9275 32283
rect 9315 32280 9343 32320
rect 9674 32308 9680 32360
rect 9732 32308 9738 32360
rect 9968 32348 9996 32379
rect 11790 32376 11796 32388
rect 11848 32376 11854 32428
rect 9784 32320 9996 32348
rect 10137 32351 10195 32357
rect 9784 32280 9812 32320
rect 10137 32317 10149 32351
rect 10183 32317 10195 32351
rect 10137 32311 10195 32317
rect 9315 32252 9812 32280
rect 10152 32280 10180 32311
rect 10226 32308 10232 32360
rect 10284 32348 10290 32360
rect 10505 32351 10563 32357
rect 10505 32348 10517 32351
rect 10284 32320 10517 32348
rect 10284 32308 10290 32320
rect 10505 32317 10517 32320
rect 10551 32317 10563 32351
rect 10505 32311 10563 32317
rect 12250 32308 12256 32360
rect 12308 32308 12314 32360
rect 10594 32280 10600 32292
rect 10152 32252 10600 32280
rect 9217 32243 9275 32249
rect 10594 32240 10600 32252
rect 10652 32240 10658 32292
rect 10134 32212 10140 32224
rect 8496 32184 10140 32212
rect 7984 32172 7990 32184
rect 10134 32172 10140 32184
rect 10192 32212 10198 32224
rect 11514 32212 11520 32224
rect 10192 32184 11520 32212
rect 10192 32172 10198 32184
rect 11514 32172 11520 32184
rect 11572 32172 11578 32224
rect 11882 32172 11888 32224
rect 11940 32212 11946 32224
rect 12158 32212 12164 32224
rect 11940 32184 12164 32212
rect 11940 32172 11946 32184
rect 12158 32172 12164 32184
rect 12216 32172 12222 32224
rect 552 32122 12604 32144
rect 552 32070 4322 32122
rect 4374 32070 4386 32122
rect 4438 32070 4450 32122
rect 4502 32070 4514 32122
rect 4566 32070 4578 32122
rect 4630 32070 10722 32122
rect 10774 32070 10786 32122
rect 10838 32070 10850 32122
rect 10902 32070 10914 32122
rect 10966 32070 10978 32122
rect 11030 32070 12604 32122
rect 552 32048 12604 32070
rect 566 31968 572 32020
rect 624 32008 630 32020
rect 1670 32008 1676 32020
rect 624 31980 796 32008
rect 624 31968 630 31980
rect 382 31832 388 31884
rect 440 31872 446 31884
rect 566 31872 572 31884
rect 440 31844 572 31872
rect 440 31832 446 31844
rect 566 31832 572 31844
rect 624 31832 630 31884
rect 768 31816 796 31980
rect 1504 31980 1676 32008
rect 842 31900 848 31952
rect 900 31940 906 31952
rect 937 31943 995 31949
rect 937 31940 949 31943
rect 900 31912 949 31940
rect 900 31900 906 31912
rect 937 31909 949 31912
rect 983 31909 995 31943
rect 937 31903 995 31909
rect 1026 31900 1032 31952
rect 1084 31940 1090 31952
rect 1504 31940 1532 31980
rect 1670 31968 1676 31980
rect 1728 31968 1734 32020
rect 2038 31968 2044 32020
rect 2096 31968 2102 32020
rect 2332 31980 3740 32008
rect 1084 31912 1532 31940
rect 2056 31940 2084 31968
rect 2332 31952 2360 31980
rect 2056 31912 2268 31940
rect 1084 31900 1090 31912
rect 2240 31884 2268 31912
rect 2314 31900 2320 31952
rect 2372 31900 2378 31952
rect 2406 31900 2412 31952
rect 2464 31940 2470 31952
rect 3513 31943 3571 31949
rect 3513 31940 3525 31943
rect 2464 31912 3525 31940
rect 2464 31900 2470 31912
rect 3513 31909 3525 31912
rect 3559 31909 3571 31943
rect 3513 31903 3571 31909
rect 1210 31832 1216 31884
rect 1268 31872 1274 31884
rect 1397 31875 1455 31881
rect 1397 31872 1409 31875
rect 1268 31844 1409 31872
rect 1268 31832 1274 31844
rect 1397 31841 1409 31844
rect 1443 31841 1455 31875
rect 1397 31835 1455 31841
rect 1581 31875 1639 31881
rect 1581 31841 1593 31875
rect 1627 31872 1639 31875
rect 1946 31872 1952 31884
rect 1627 31844 1952 31872
rect 1627 31841 1639 31844
rect 1581 31835 1639 31841
rect 1946 31832 1952 31844
rect 2004 31832 2010 31884
rect 2041 31875 2099 31881
rect 2041 31841 2053 31875
rect 2087 31872 2099 31875
rect 2130 31872 2136 31884
rect 2087 31844 2136 31872
rect 2087 31841 2099 31844
rect 2041 31835 2099 31841
rect 2130 31832 2136 31844
rect 2188 31832 2194 31884
rect 2222 31832 2228 31884
rect 2280 31832 2286 31884
rect 2590 31832 2596 31884
rect 2648 31832 2654 31884
rect 2866 31832 2872 31884
rect 2924 31832 2930 31884
rect 3712 31881 3740 31980
rect 5442 31968 5448 32020
rect 5500 32008 5506 32020
rect 5902 32008 5908 32020
rect 5500 31980 5908 32008
rect 5500 31968 5506 31980
rect 5902 31968 5908 31980
rect 5960 31968 5966 32020
rect 5997 32011 6055 32017
rect 5997 31977 6009 32011
rect 6043 32008 6055 32011
rect 6638 32008 6644 32020
rect 6043 31980 6644 32008
rect 6043 31977 6055 31980
rect 5997 31971 6055 31977
rect 6638 31968 6644 31980
rect 6696 31968 6702 32020
rect 7006 31968 7012 32020
rect 7064 32008 7070 32020
rect 7064 31980 7880 32008
rect 7064 31968 7070 31980
rect 3786 31900 3792 31952
rect 3844 31940 3850 31952
rect 4893 31943 4951 31949
rect 4893 31940 4905 31943
rect 3844 31912 4905 31940
rect 3844 31900 3850 31912
rect 4893 31909 4905 31912
rect 4939 31909 4951 31943
rect 6086 31940 6092 31952
rect 4893 31903 4951 31909
rect 5184 31912 6092 31940
rect 3697 31875 3755 31881
rect 3068 31844 3372 31872
rect 750 31764 756 31816
rect 808 31764 814 31816
rect 1486 31764 1492 31816
rect 1544 31804 1550 31816
rect 1673 31807 1731 31813
rect 1673 31804 1685 31807
rect 1544 31776 1685 31804
rect 1544 31764 1550 31776
rect 1673 31773 1685 31776
rect 1719 31773 1731 31807
rect 1673 31767 1731 31773
rect 2498 31764 2504 31816
rect 2556 31804 2562 31816
rect 3068 31804 3096 31844
rect 2556 31776 3096 31804
rect 2556 31764 2562 31776
rect 3234 31764 3240 31816
rect 3292 31764 3298 31816
rect 3344 31736 3372 31844
rect 3697 31841 3709 31875
rect 3743 31841 3755 31875
rect 4249 31875 4307 31881
rect 4249 31872 4261 31875
rect 3697 31835 3755 31841
rect 3804 31844 4261 31872
rect 3418 31764 3424 31816
rect 3476 31804 3482 31816
rect 3804 31804 3832 31844
rect 4249 31841 4261 31844
rect 4295 31841 4307 31875
rect 4249 31835 4307 31841
rect 4525 31875 4583 31881
rect 4525 31841 4537 31875
rect 4571 31872 4583 31875
rect 4614 31872 4620 31884
rect 4571 31844 4620 31872
rect 4571 31841 4583 31844
rect 4525 31835 4583 31841
rect 4614 31832 4620 31844
rect 4672 31872 4678 31884
rect 4982 31872 4988 31884
rect 4672 31844 4988 31872
rect 4672 31832 4678 31844
rect 4982 31832 4988 31844
rect 5040 31832 5046 31884
rect 5074 31832 5080 31884
rect 5132 31832 5138 31884
rect 5184 31881 5212 31912
rect 6086 31900 6092 31912
rect 6144 31900 6150 31952
rect 6362 31900 6368 31952
rect 6420 31900 6426 31952
rect 6549 31943 6607 31949
rect 6549 31909 6561 31943
rect 6595 31940 6607 31943
rect 6730 31940 6736 31952
rect 6595 31912 6736 31940
rect 6595 31909 6607 31912
rect 6549 31903 6607 31909
rect 6730 31900 6736 31912
rect 6788 31900 6794 31952
rect 7558 31940 7564 31952
rect 7392 31912 7564 31940
rect 5169 31875 5227 31881
rect 5169 31841 5181 31875
rect 5215 31841 5227 31875
rect 5169 31835 5227 31841
rect 5442 31832 5448 31884
rect 5500 31832 5506 31884
rect 5534 31832 5540 31884
rect 5592 31832 5598 31884
rect 5813 31875 5871 31881
rect 5813 31841 5825 31875
rect 5859 31872 5871 31875
rect 5994 31872 6000 31884
rect 5859 31844 6000 31872
rect 5859 31841 5871 31844
rect 5813 31835 5871 31841
rect 5994 31832 6000 31844
rect 6052 31832 6058 31884
rect 6270 31832 6276 31884
rect 6328 31832 6334 31884
rect 6380 31872 6408 31900
rect 6380 31844 6592 31872
rect 3973 31807 4031 31813
rect 3973 31804 3985 31807
rect 3476 31776 3832 31804
rect 3896 31776 3985 31804
rect 3476 31764 3482 31776
rect 3896 31736 3924 31776
rect 3973 31773 3985 31776
rect 4019 31773 4031 31807
rect 3973 31767 4031 31773
rect 5350 31764 5356 31816
rect 5408 31764 5414 31816
rect 6362 31764 6368 31816
rect 6420 31764 6426 31816
rect 6454 31764 6460 31816
rect 6512 31764 6518 31816
rect 6564 31804 6592 31844
rect 6638 31832 6644 31884
rect 6696 31832 6702 31884
rect 7392 31881 7420 31912
rect 7558 31900 7564 31912
rect 7616 31900 7622 31952
rect 7852 31881 7880 31980
rect 7926 31968 7932 32020
rect 7984 31968 7990 32020
rect 8021 32011 8079 32017
rect 8021 31977 8033 32011
rect 8067 32008 8079 32011
rect 8110 32008 8116 32020
rect 8067 31980 8116 32008
rect 8067 31977 8079 31980
rect 8021 31971 8079 31977
rect 8110 31968 8116 31980
rect 8168 31968 8174 32020
rect 8202 31968 8208 32020
rect 8260 32008 8266 32020
rect 8478 32008 8484 32020
rect 8260 31980 8484 32008
rect 8260 31968 8266 31980
rect 8478 31968 8484 31980
rect 8536 31968 8542 32020
rect 8570 31968 8576 32020
rect 8628 32008 8634 32020
rect 8628 31980 9076 32008
rect 8628 31968 8634 31980
rect 7009 31875 7067 31881
rect 7009 31872 7021 31875
rect 6748 31844 7021 31872
rect 6748 31804 6776 31844
rect 7009 31841 7021 31844
rect 7055 31841 7067 31875
rect 7009 31835 7067 31841
rect 7377 31875 7435 31881
rect 7377 31841 7389 31875
rect 7423 31841 7435 31875
rect 7377 31835 7435 31841
rect 7469 31875 7527 31881
rect 7469 31841 7481 31875
rect 7515 31841 7527 31875
rect 7469 31835 7527 31841
rect 7745 31875 7803 31881
rect 7745 31841 7757 31875
rect 7791 31841 7803 31875
rect 7745 31835 7803 31841
rect 7837 31875 7895 31881
rect 7837 31841 7849 31875
rect 7883 31841 7895 31875
rect 7944 31872 7972 31968
rect 8386 31900 8392 31952
rect 8444 31940 8450 31952
rect 8754 31940 8760 31952
rect 8444 31912 8524 31940
rect 8444 31900 8450 31912
rect 8021 31875 8079 31881
rect 8021 31872 8033 31875
rect 7944 31844 8033 31872
rect 7837 31835 7895 31841
rect 8021 31841 8033 31844
rect 8067 31841 8079 31875
rect 8294 31872 8300 31884
rect 8021 31835 8079 31841
rect 8220 31844 8300 31872
rect 6564 31776 6776 31804
rect 1228 31708 2912 31736
rect 3344 31708 3924 31736
rect 1228 31680 1256 31708
rect 1210 31628 1216 31680
rect 1268 31628 1274 31680
rect 2225 31671 2283 31677
rect 2225 31637 2237 31671
rect 2271 31668 2283 31671
rect 2774 31668 2780 31680
rect 2271 31640 2780 31668
rect 2271 31637 2283 31640
rect 2225 31631 2283 31637
rect 2774 31628 2780 31640
rect 2832 31628 2838 31680
rect 2884 31668 2912 31708
rect 4154 31696 4160 31748
rect 4212 31736 4218 31748
rect 4212 31708 4476 31736
rect 4212 31696 4218 31708
rect 4448 31680 4476 31708
rect 4706 31696 4712 31748
rect 4764 31736 4770 31748
rect 5442 31736 5448 31748
rect 4764 31708 5448 31736
rect 4764 31696 4770 31708
rect 5442 31696 5448 31708
rect 5500 31696 5506 31748
rect 6089 31739 6147 31745
rect 6089 31705 6101 31739
rect 6135 31736 6147 31739
rect 6472 31736 6500 31764
rect 6135 31708 6500 31736
rect 6135 31705 6147 31708
rect 6089 31699 6147 31705
rect 7006 31696 7012 31748
rect 7064 31736 7070 31748
rect 7484 31736 7512 31835
rect 7760 31804 7788 31835
rect 7926 31804 7932 31816
rect 7760 31776 7932 31804
rect 7926 31764 7932 31776
rect 7984 31764 7990 31816
rect 8220 31736 8248 31844
rect 8294 31832 8300 31844
rect 8352 31872 8358 31884
rect 8496 31881 8524 31912
rect 8680 31912 8760 31940
rect 8481 31875 8539 31881
rect 8352 31844 8397 31872
rect 8352 31832 8358 31844
rect 8481 31841 8493 31875
rect 8527 31841 8539 31875
rect 8481 31835 8539 31841
rect 8570 31832 8576 31884
rect 8628 31832 8634 31884
rect 7064 31708 7512 31736
rect 7944 31708 8248 31736
rect 8389 31739 8447 31745
rect 7064 31696 7070 31708
rect 7944 31680 7972 31708
rect 8389 31705 8401 31739
rect 8435 31736 8447 31739
rect 8680 31736 8708 31912
rect 8754 31900 8760 31912
rect 8812 31900 8818 31952
rect 8849 31943 8907 31949
rect 8849 31909 8861 31943
rect 8895 31940 8907 31943
rect 8938 31940 8944 31952
rect 8895 31912 8944 31940
rect 8895 31909 8907 31912
rect 8849 31903 8907 31909
rect 8938 31900 8944 31912
rect 8996 31900 9002 31952
rect 9048 31881 9076 31980
rect 9490 31968 9496 32020
rect 9548 32008 9554 32020
rect 9548 31980 12080 32008
rect 9548 31968 9554 31980
rect 10870 31940 10876 31952
rect 9324 31912 10876 31940
rect 9033 31875 9091 31881
rect 8757 31865 8815 31871
rect 8757 31831 8769 31865
rect 8803 31831 8815 31865
rect 9033 31841 9045 31875
rect 9079 31841 9091 31875
rect 9033 31835 9091 31841
rect 8757 31825 8815 31831
rect 8772 31748 8800 31825
rect 8938 31764 8944 31816
rect 8996 31804 9002 31816
rect 9048 31804 9076 31835
rect 9122 31832 9128 31884
rect 9180 31872 9186 31884
rect 9324 31881 9352 31912
rect 10870 31900 10876 31912
rect 10928 31900 10934 31952
rect 12052 31940 12080 31980
rect 12052 31912 12112 31940
rect 9309 31875 9367 31881
rect 9309 31872 9321 31875
rect 9180 31844 9321 31872
rect 9180 31832 9186 31844
rect 9309 31841 9321 31844
rect 9355 31841 9367 31875
rect 9309 31835 9367 31841
rect 9398 31832 9404 31884
rect 9456 31872 9462 31884
rect 9565 31875 9623 31881
rect 9565 31872 9577 31875
rect 9456 31844 9577 31872
rect 9456 31832 9462 31844
rect 9565 31841 9577 31844
rect 9611 31841 9623 31875
rect 9565 31835 9623 31841
rect 10962 31832 10968 31884
rect 11020 31832 11026 31884
rect 11149 31875 11207 31881
rect 11149 31841 11161 31875
rect 11195 31872 11207 31875
rect 11606 31872 11612 31884
rect 11195 31844 11612 31872
rect 11195 31841 11207 31844
rect 11149 31835 11207 31841
rect 11606 31832 11612 31844
rect 11664 31832 11670 31884
rect 11701 31875 11759 31881
rect 11701 31841 11713 31875
rect 11747 31841 11759 31875
rect 11701 31835 11759 31841
rect 11716 31804 11744 31835
rect 11790 31832 11796 31884
rect 11848 31872 11854 31884
rect 12084 31881 12112 31912
rect 12069 31875 12127 31881
rect 11848 31844 12020 31872
rect 11848 31832 11854 31844
rect 8996 31776 9076 31804
rect 11440 31776 11744 31804
rect 11885 31807 11943 31813
rect 8996 31764 9002 31776
rect 8435 31708 8708 31736
rect 8435 31705 8447 31708
rect 8389 31699 8447 31705
rect 8754 31696 8760 31748
rect 8812 31696 8818 31748
rect 10870 31696 10876 31748
rect 10928 31736 10934 31748
rect 11440 31736 11468 31776
rect 11885 31773 11897 31807
rect 11931 31773 11943 31807
rect 11992 31804 12020 31844
rect 12069 31841 12081 31875
rect 12115 31841 12127 31875
rect 12069 31835 12127 31841
rect 12253 31807 12311 31813
rect 12253 31804 12265 31807
rect 11992 31776 12265 31804
rect 11885 31767 11943 31773
rect 12253 31773 12265 31776
rect 12299 31804 12311 31807
rect 12526 31804 12532 31816
rect 12299 31776 12532 31804
rect 12299 31773 12311 31776
rect 12253 31767 12311 31773
rect 10928 31708 11468 31736
rect 10928 31696 10934 31708
rect 3881 31671 3939 31677
rect 3881 31668 3893 31671
rect 2884 31640 3893 31668
rect 3881 31637 3893 31640
rect 3927 31637 3939 31671
rect 3881 31631 3939 31637
rect 4062 31628 4068 31680
rect 4120 31628 4126 31680
rect 4430 31628 4436 31680
rect 4488 31628 4494 31680
rect 5902 31628 5908 31680
rect 5960 31668 5966 31680
rect 6549 31671 6607 31677
rect 6549 31668 6561 31671
rect 5960 31640 6561 31668
rect 5960 31628 5966 31640
rect 6549 31637 6561 31640
rect 6595 31668 6607 31671
rect 7098 31668 7104 31680
rect 6595 31640 7104 31668
rect 6595 31637 6607 31640
rect 6549 31631 6607 31637
rect 7098 31628 7104 31640
rect 7156 31628 7162 31680
rect 7193 31671 7251 31677
rect 7193 31637 7205 31671
rect 7239 31668 7251 31671
rect 7282 31668 7288 31680
rect 7239 31640 7288 31668
rect 7239 31637 7251 31640
rect 7193 31631 7251 31637
rect 7282 31628 7288 31640
rect 7340 31628 7346 31680
rect 7558 31628 7564 31680
rect 7616 31668 7622 31680
rect 7653 31671 7711 31677
rect 7653 31668 7665 31671
rect 7616 31640 7665 31668
rect 7616 31628 7622 31640
rect 7653 31637 7665 31640
rect 7699 31637 7711 31671
rect 7653 31631 7711 31637
rect 7926 31628 7932 31680
rect 7984 31628 7990 31680
rect 8113 31671 8171 31677
rect 8113 31637 8125 31671
rect 8159 31668 8171 31671
rect 8202 31668 8208 31680
rect 8159 31640 8208 31668
rect 8159 31637 8171 31640
rect 8113 31631 8171 31637
rect 8202 31628 8208 31640
rect 8260 31628 8266 31680
rect 8294 31628 8300 31680
rect 8352 31668 8358 31680
rect 9217 31671 9275 31677
rect 9217 31668 9229 31671
rect 8352 31640 9229 31668
rect 8352 31628 8358 31640
rect 9217 31637 9229 31640
rect 9263 31637 9275 31671
rect 9217 31631 9275 31637
rect 10686 31628 10692 31680
rect 10744 31628 10750 31680
rect 11146 31628 11152 31680
rect 11204 31628 11210 31680
rect 11440 31668 11468 31708
rect 11514 31696 11520 31748
rect 11572 31736 11578 31748
rect 11900 31736 11928 31767
rect 12526 31764 12532 31776
rect 12584 31764 12590 31816
rect 12342 31736 12348 31748
rect 11572 31708 12348 31736
rect 11572 31696 11578 31708
rect 12342 31696 12348 31708
rect 12400 31696 12406 31748
rect 12250 31668 12256 31680
rect 11440 31640 12256 31668
rect 12250 31628 12256 31640
rect 12308 31628 12314 31680
rect 552 31578 12604 31600
rect 552 31526 3662 31578
rect 3714 31526 3726 31578
rect 3778 31526 3790 31578
rect 3842 31526 3854 31578
rect 3906 31526 3918 31578
rect 3970 31526 10062 31578
rect 10114 31526 10126 31578
rect 10178 31526 10190 31578
rect 10242 31526 10254 31578
rect 10306 31526 10318 31578
rect 10370 31526 12604 31578
rect 552 31504 12604 31526
rect 845 31467 903 31473
rect 845 31433 857 31467
rect 891 31464 903 31467
rect 1486 31464 1492 31476
rect 891 31436 1492 31464
rect 891 31433 903 31436
rect 845 31427 903 31433
rect 1486 31424 1492 31436
rect 1544 31424 1550 31476
rect 2222 31424 2228 31476
rect 2280 31464 2286 31476
rect 3234 31464 3240 31476
rect 2280 31436 3240 31464
rect 2280 31424 2286 31436
rect 3234 31424 3240 31436
rect 3292 31424 3298 31476
rect 3418 31424 3424 31476
rect 3476 31424 3482 31476
rect 5350 31424 5356 31476
rect 5408 31464 5414 31476
rect 5445 31467 5503 31473
rect 5445 31464 5457 31467
rect 5408 31436 5457 31464
rect 5408 31424 5414 31436
rect 5445 31433 5457 31436
rect 5491 31433 5503 31467
rect 5445 31427 5503 31433
rect 5810 31424 5816 31476
rect 5868 31424 5874 31476
rect 6089 31467 6147 31473
rect 6089 31433 6101 31467
rect 6135 31464 6147 31467
rect 6914 31464 6920 31476
rect 6135 31436 6920 31464
rect 6135 31433 6147 31436
rect 6089 31427 6147 31433
rect 6914 31424 6920 31436
rect 6972 31424 6978 31476
rect 8938 31424 8944 31476
rect 8996 31464 9002 31476
rect 10134 31464 10140 31476
rect 8996 31436 10140 31464
rect 8996 31424 9002 31436
rect 10134 31424 10140 31436
rect 10192 31424 10198 31476
rect 10410 31424 10416 31476
rect 10468 31424 10474 31476
rect 2409 31399 2467 31405
rect 2409 31365 2421 31399
rect 2455 31365 2467 31399
rect 2682 31396 2688 31408
rect 2409 31359 2467 31365
rect 2608 31368 2688 31396
rect 2424 31328 2452 31359
rect 2148 31300 2452 31328
rect 1946 31220 1952 31272
rect 2004 31269 2010 31272
rect 2004 31260 2016 31269
rect 2004 31232 2049 31260
rect 2004 31223 2016 31232
rect 2004 31220 2010 31223
rect 1670 31152 1676 31204
rect 1728 31192 1734 31204
rect 2148 31192 2176 31300
rect 2222 31220 2228 31272
rect 2280 31260 2286 31272
rect 2608 31260 2636 31368
rect 2682 31356 2688 31368
rect 2740 31356 2746 31408
rect 5169 31399 5227 31405
rect 5169 31365 5181 31399
rect 5215 31396 5227 31399
rect 5534 31396 5540 31408
rect 5215 31368 5540 31396
rect 5215 31365 5227 31368
rect 5169 31359 5227 31365
rect 5534 31356 5540 31368
rect 5592 31356 5598 31408
rect 5828 31396 5856 31424
rect 5828 31368 6316 31396
rect 3142 31288 3148 31340
rect 3200 31328 3206 31340
rect 3237 31331 3295 31337
rect 3237 31328 3249 31331
rect 3200 31300 3249 31328
rect 3200 31288 3206 31300
rect 3237 31297 3249 31300
rect 3283 31297 3295 31331
rect 5810 31328 5816 31340
rect 3237 31291 3295 31297
rect 5644 31300 5816 31328
rect 2280 31232 2636 31260
rect 2280 31220 2286 31232
rect 2682 31220 2688 31272
rect 2740 31220 2746 31272
rect 2777 31263 2835 31269
rect 2777 31229 2789 31263
rect 2823 31260 2835 31263
rect 3326 31260 3332 31272
rect 2823 31232 3332 31260
rect 2823 31229 2835 31232
rect 2777 31223 2835 31229
rect 3326 31220 3332 31232
rect 3384 31220 3390 31272
rect 3697 31263 3755 31269
rect 3697 31229 3709 31263
rect 3743 31229 3755 31263
rect 3697 31223 3755 31229
rect 1728 31164 2176 31192
rect 2409 31195 2467 31201
rect 1728 31152 1734 31164
rect 2409 31161 2421 31195
rect 2455 31161 2467 31195
rect 2409 31155 2467 31161
rect 1486 31084 1492 31136
rect 1544 31124 1550 31136
rect 2424 31124 2452 31155
rect 2498 31152 2504 31204
rect 2556 31192 2562 31204
rect 2593 31195 2651 31201
rect 2593 31192 2605 31195
rect 2556 31164 2605 31192
rect 2556 31152 2562 31164
rect 2593 31161 2605 31164
rect 2639 31161 2651 31195
rect 2593 31155 2651 31161
rect 2961 31195 3019 31201
rect 2961 31161 2973 31195
rect 3007 31192 3019 31195
rect 3142 31192 3148 31204
rect 3007 31164 3148 31192
rect 3007 31161 3019 31164
rect 2961 31155 3019 31161
rect 3142 31152 3148 31164
rect 3200 31152 3206 31204
rect 3712 31192 3740 31223
rect 3786 31220 3792 31272
rect 3844 31220 3850 31272
rect 4056 31263 4114 31269
rect 4056 31229 4068 31263
rect 4102 31260 4114 31263
rect 4522 31260 4528 31272
rect 4102 31232 4528 31260
rect 4102 31229 4114 31232
rect 4056 31223 4114 31229
rect 4522 31220 4528 31232
rect 4580 31220 4586 31272
rect 5644 31269 5672 31300
rect 5810 31288 5816 31300
rect 5868 31288 5874 31340
rect 5994 31288 6000 31340
rect 6052 31288 6058 31340
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31229 5687 31263
rect 5629 31223 5687 31229
rect 5721 31263 5779 31269
rect 5721 31229 5733 31263
rect 5767 31260 5779 31263
rect 5905 31263 5963 31269
rect 5767 31232 5856 31260
rect 5767 31229 5779 31232
rect 5721 31223 5779 31229
rect 5828 31204 5856 31232
rect 5905 31229 5917 31263
rect 5951 31229 5963 31263
rect 6012 31247 6040 31288
rect 6288 31260 6316 31368
rect 7190 31356 7196 31408
rect 7248 31356 7254 31408
rect 7208 31328 7236 31356
rect 7208 31300 8432 31328
rect 6365 31263 6423 31269
rect 6365 31260 6377 31263
rect 5905 31223 5963 31229
rect 5997 31241 6055 31247
rect 4430 31192 4436 31204
rect 3712 31164 4436 31192
rect 4430 31152 4436 31164
rect 4488 31152 4494 31204
rect 5810 31152 5816 31204
rect 5868 31152 5874 31204
rect 3050 31124 3056 31136
rect 1544 31096 3056 31124
rect 1544 31084 1550 31096
rect 3050 31084 3056 31096
rect 3108 31084 3114 31136
rect 3605 31127 3663 31133
rect 3605 31093 3617 31127
rect 3651 31124 3663 31127
rect 4614 31124 4620 31136
rect 3651 31096 4620 31124
rect 3651 31093 3663 31096
rect 3605 31087 3663 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 5258 31084 5264 31136
rect 5316 31124 5322 31136
rect 5920 31124 5948 31223
rect 5997 31207 6009 31241
rect 6043 31207 6055 31241
rect 6288 31232 6377 31260
rect 6365 31229 6377 31232
rect 6411 31229 6423 31263
rect 6365 31223 6423 31229
rect 6454 31220 6460 31272
rect 6512 31220 6518 31272
rect 6546 31220 6552 31272
rect 6604 31220 6610 31272
rect 6641 31263 6699 31269
rect 6641 31229 6653 31263
rect 6687 31260 6699 31263
rect 6730 31260 6736 31272
rect 6687 31232 6736 31260
rect 6687 31229 6699 31232
rect 6641 31223 6699 31229
rect 6730 31220 6736 31232
rect 6788 31220 6794 31272
rect 6825 31263 6883 31269
rect 6825 31229 6837 31263
rect 6871 31260 6883 31263
rect 6914 31260 6920 31272
rect 6871 31232 6920 31260
rect 6871 31229 6883 31232
rect 6825 31223 6883 31229
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 7101 31263 7159 31269
rect 7101 31229 7113 31263
rect 7147 31260 7159 31263
rect 7190 31260 7196 31272
rect 7147 31232 7196 31260
rect 7147 31229 7159 31232
rect 7101 31223 7159 31229
rect 7190 31220 7196 31232
rect 7248 31220 7254 31272
rect 7282 31220 7288 31272
rect 7340 31220 7346 31272
rect 7392 31269 7420 31300
rect 7377 31263 7435 31269
rect 7377 31229 7389 31263
rect 7423 31229 7435 31263
rect 7377 31223 7435 31229
rect 7469 31263 7527 31269
rect 7469 31229 7481 31263
rect 7515 31260 7527 31263
rect 7650 31260 7656 31272
rect 7515 31232 7656 31260
rect 7515 31229 7527 31232
rect 7469 31223 7527 31229
rect 7650 31220 7656 31232
rect 7708 31220 7714 31272
rect 8021 31263 8079 31269
rect 8021 31229 8033 31263
rect 8067 31260 8079 31263
rect 8110 31260 8116 31272
rect 8067 31232 8116 31260
rect 8067 31229 8079 31232
rect 8021 31223 8079 31229
rect 8110 31220 8116 31232
rect 8168 31220 8174 31272
rect 8404 31269 8432 31300
rect 10870 31288 10876 31340
rect 10928 31288 10934 31340
rect 8389 31263 8447 31269
rect 8389 31229 8401 31263
rect 8435 31229 8447 31263
rect 8389 31223 8447 31229
rect 9033 31263 9091 31269
rect 9033 31229 9045 31263
rect 9079 31260 9091 31263
rect 9122 31260 9128 31272
rect 9079 31232 9128 31260
rect 9079 31229 9091 31232
rect 9033 31223 9091 31229
rect 9122 31220 9128 31232
rect 9180 31220 9186 31272
rect 9766 31220 9772 31272
rect 9824 31260 9830 31272
rect 11146 31269 11152 31272
rect 10505 31263 10563 31269
rect 10505 31260 10517 31263
rect 9824 31232 10517 31260
rect 9824 31220 9830 31232
rect 10505 31229 10517 31232
rect 10551 31229 10563 31263
rect 11140 31260 11152 31269
rect 11107 31232 11152 31260
rect 10505 31223 10563 31229
rect 11140 31223 11152 31232
rect 11146 31220 11152 31223
rect 11204 31220 11210 31272
rect 5997 31201 6055 31207
rect 6932 31192 6960 31220
rect 7558 31192 7564 31204
rect 6932 31164 7564 31192
rect 7558 31152 7564 31164
rect 7616 31152 7622 31204
rect 7668 31192 7696 31220
rect 8205 31195 8263 31201
rect 8205 31192 8217 31195
rect 7668 31164 8217 31192
rect 8205 31161 8217 31164
rect 8251 31192 8263 31195
rect 8294 31192 8300 31204
rect 8251 31164 8300 31192
rect 8251 31161 8263 31164
rect 8205 31155 8263 31161
rect 8294 31152 8300 31164
rect 8352 31152 8358 31204
rect 8665 31195 8723 31201
rect 8665 31161 8677 31195
rect 8711 31192 8723 31195
rect 8938 31192 8944 31204
rect 8711 31164 8944 31192
rect 8711 31161 8723 31164
rect 8665 31155 8723 31161
rect 8938 31152 8944 31164
rect 8996 31152 9002 31204
rect 9300 31195 9358 31201
rect 9300 31161 9312 31195
rect 9346 31192 9358 31195
rect 9582 31192 9588 31204
rect 9346 31164 9588 31192
rect 9346 31161 9358 31164
rect 9300 31155 9358 31161
rect 9582 31152 9588 31164
rect 9640 31152 9646 31204
rect 7006 31124 7012 31136
rect 5316 31096 7012 31124
rect 5316 31084 5322 31096
rect 7006 31084 7012 31096
rect 7064 31084 7070 31136
rect 7650 31084 7656 31136
rect 7708 31124 7714 31136
rect 7745 31127 7803 31133
rect 7745 31124 7757 31127
rect 7708 31096 7757 31124
rect 7708 31084 7714 31096
rect 7745 31093 7757 31096
rect 7791 31093 7803 31127
rect 7745 31087 7803 31093
rect 7834 31084 7840 31136
rect 7892 31084 7898 31136
rect 9122 31084 9128 31136
rect 9180 31124 9186 31136
rect 10689 31127 10747 31133
rect 10689 31124 10701 31127
rect 9180 31096 10701 31124
rect 9180 31084 9186 31096
rect 10689 31093 10701 31096
rect 10735 31124 10747 31127
rect 11146 31124 11152 31136
rect 10735 31096 11152 31124
rect 10735 31093 10747 31096
rect 10689 31087 10747 31093
rect 11146 31084 11152 31096
rect 11204 31084 11210 31136
rect 11422 31084 11428 31136
rect 11480 31124 11486 31136
rect 12253 31127 12311 31133
rect 12253 31124 12265 31127
rect 11480 31096 12265 31124
rect 11480 31084 11486 31096
rect 12253 31093 12265 31096
rect 12299 31124 12311 31127
rect 12299 31096 12756 31124
rect 12299 31093 12311 31096
rect 12253 31087 12311 31093
rect 552 31034 12604 31056
rect 552 30982 4322 31034
rect 4374 30982 4386 31034
rect 4438 30982 4450 31034
rect 4502 30982 4514 31034
rect 4566 30982 4578 31034
rect 4630 30982 10722 31034
rect 10774 30982 10786 31034
rect 10838 30982 10850 31034
rect 10902 30982 10914 31034
rect 10966 30982 10978 31034
rect 11030 30982 12604 31034
rect 552 30960 12604 30982
rect 2774 30880 2780 30932
rect 2832 30920 2838 30932
rect 2832 30892 3372 30920
rect 2832 30880 2838 30892
rect 934 30812 940 30864
rect 992 30852 998 30864
rect 2590 30852 2596 30864
rect 992 30824 2596 30852
rect 992 30812 998 30824
rect 2590 30812 2596 30824
rect 2648 30852 2654 30864
rect 2648 30824 2820 30852
rect 2648 30812 2654 30824
rect 1394 30744 1400 30796
rect 1452 30784 1458 30796
rect 1958 30787 2016 30793
rect 1958 30784 1970 30787
rect 1452 30756 1970 30784
rect 1452 30744 1458 30756
rect 1958 30753 1970 30756
rect 2004 30784 2016 30787
rect 2317 30787 2375 30793
rect 2317 30784 2329 30787
rect 2004 30756 2329 30784
rect 2004 30753 2016 30756
rect 1958 30747 2016 30753
rect 2317 30753 2329 30756
rect 2363 30753 2375 30787
rect 2317 30747 2375 30753
rect 2406 30744 2412 30796
rect 2464 30784 2470 30796
rect 2792 30793 2820 30824
rect 2501 30787 2559 30793
rect 2501 30784 2513 30787
rect 2464 30756 2513 30784
rect 2464 30744 2470 30756
rect 2501 30753 2513 30756
rect 2547 30753 2559 30787
rect 2501 30747 2559 30753
rect 2777 30787 2835 30793
rect 2777 30753 2789 30787
rect 2823 30753 2835 30787
rect 2777 30747 2835 30753
rect 3142 30744 3148 30796
rect 3200 30784 3206 30796
rect 3237 30787 3295 30793
rect 3237 30784 3249 30787
rect 3200 30756 3249 30784
rect 3200 30744 3206 30756
rect 3237 30753 3249 30756
rect 3283 30753 3295 30787
rect 3344 30784 3372 30892
rect 3510 30880 3516 30932
rect 3568 30920 3574 30932
rect 4430 30920 4436 30932
rect 3568 30892 4436 30920
rect 3568 30880 3574 30892
rect 4430 30880 4436 30892
rect 4488 30880 4494 30932
rect 4706 30880 4712 30932
rect 4764 30920 4770 30932
rect 5077 30923 5135 30929
rect 5077 30920 5089 30923
rect 4764 30892 5089 30920
rect 4764 30880 4770 30892
rect 5077 30889 5089 30892
rect 5123 30920 5135 30923
rect 5166 30920 5172 30932
rect 5123 30892 5172 30920
rect 5123 30889 5135 30892
rect 5077 30883 5135 30889
rect 5166 30880 5172 30892
rect 5224 30880 5230 30932
rect 5350 30880 5356 30932
rect 5408 30920 5414 30932
rect 5905 30923 5963 30929
rect 5905 30920 5917 30923
rect 5408 30892 5917 30920
rect 5408 30880 5414 30892
rect 5905 30889 5917 30892
rect 5951 30889 5963 30923
rect 5905 30883 5963 30889
rect 3964 30855 4022 30861
rect 3964 30821 3976 30855
rect 4010 30852 4022 30855
rect 4062 30852 4068 30864
rect 4010 30824 4068 30852
rect 4010 30821 4022 30824
rect 3964 30815 4022 30821
rect 4062 30812 4068 30824
rect 4120 30812 4126 30864
rect 5920 30852 5948 30883
rect 6454 30880 6460 30932
rect 6512 30920 6518 30932
rect 6733 30923 6791 30929
rect 6733 30920 6745 30923
rect 6512 30892 6745 30920
rect 6512 30880 6518 30892
rect 6733 30889 6745 30892
rect 6779 30889 6791 30923
rect 6733 30883 6791 30889
rect 6825 30923 6883 30929
rect 6825 30889 6837 30923
rect 6871 30920 6883 30923
rect 7098 30920 7104 30932
rect 6871 30892 7104 30920
rect 6871 30889 6883 30892
rect 6825 30883 6883 30889
rect 7098 30880 7104 30892
rect 7156 30880 7162 30932
rect 7834 30920 7840 30932
rect 7300 30892 7840 30920
rect 7300 30861 7328 30892
rect 7834 30880 7840 30892
rect 7892 30880 7898 30932
rect 8570 30880 8576 30932
rect 8628 30920 8634 30932
rect 8941 30923 8999 30929
rect 8941 30920 8953 30923
rect 8628 30892 8953 30920
rect 8628 30880 8634 30892
rect 8941 30889 8953 30892
rect 8987 30889 8999 30923
rect 8941 30883 8999 30889
rect 9582 30880 9588 30932
rect 9640 30880 9646 30932
rect 9876 30892 10456 30920
rect 7285 30855 7343 30861
rect 5920 30824 6500 30852
rect 6472 30796 6500 30824
rect 6561 30824 7236 30852
rect 3510 30784 3516 30796
rect 3344 30756 3516 30784
rect 3237 30747 3295 30753
rect 3510 30744 3516 30756
rect 3568 30744 3574 30796
rect 3786 30784 3792 30796
rect 3712 30756 3792 30784
rect 2222 30676 2228 30728
rect 2280 30716 2286 30728
rect 3712 30725 3740 30756
rect 3786 30744 3792 30756
rect 3844 30744 3850 30796
rect 5350 30744 5356 30796
rect 5408 30744 5414 30796
rect 5629 30787 5687 30793
rect 5629 30753 5641 30787
rect 5675 30784 5687 30787
rect 6089 30787 6147 30793
rect 5675 30756 6040 30784
rect 5675 30753 5687 30756
rect 5629 30747 5687 30753
rect 3697 30719 3755 30725
rect 3697 30716 3709 30719
rect 2280 30688 3709 30716
rect 2280 30676 2286 30688
rect 3697 30685 3709 30688
rect 3743 30685 3755 30719
rect 3697 30679 3755 30685
rect 5258 30676 5264 30728
rect 5316 30716 5322 30728
rect 5537 30719 5595 30725
rect 5537 30716 5549 30719
rect 5316 30688 5549 30716
rect 5316 30676 5322 30688
rect 5537 30685 5549 30688
rect 5583 30685 5595 30719
rect 5537 30679 5595 30685
rect 6012 30660 6040 30756
rect 6089 30753 6101 30787
rect 6135 30784 6147 30787
rect 6362 30784 6368 30796
rect 6135 30756 6368 30784
rect 6135 30753 6147 30756
rect 6089 30747 6147 30753
rect 6362 30744 6368 30756
rect 6420 30744 6426 30796
rect 6454 30744 6460 30796
rect 6512 30744 6518 30796
rect 6561 30793 6589 30824
rect 6549 30787 6607 30793
rect 6549 30753 6561 30787
rect 6595 30753 6607 30787
rect 6549 30747 6607 30753
rect 7006 30744 7012 30796
rect 7064 30744 7070 30796
rect 7208 30784 7236 30824
rect 7285 30821 7297 30855
rect 7331 30821 7343 30855
rect 8662 30852 8668 30864
rect 7285 30815 7343 30821
rect 7392 30824 8668 30852
rect 7392 30784 7420 30824
rect 8662 30812 8668 30824
rect 8720 30812 8726 30864
rect 8846 30852 8852 30864
rect 8772 30824 8852 30852
rect 7208 30756 7420 30784
rect 7466 30744 7472 30796
rect 7524 30744 7530 30796
rect 7650 30744 7656 30796
rect 7708 30744 7714 30796
rect 7834 30744 7840 30796
rect 7892 30744 7898 30796
rect 8110 30744 8116 30796
rect 8168 30744 8174 30796
rect 8202 30744 8208 30796
rect 8260 30744 8266 30796
rect 7193 30719 7251 30725
rect 7193 30685 7205 30719
rect 7239 30685 7251 30719
rect 7193 30679 7251 30685
rect 5994 30608 6000 30660
rect 6052 30648 6058 30660
rect 7208 30648 7236 30679
rect 7282 30676 7288 30728
rect 7340 30716 7346 30728
rect 7558 30716 7564 30728
rect 7340 30688 7564 30716
rect 7340 30676 7346 30688
rect 7558 30676 7564 30688
rect 7616 30716 7622 30728
rect 8573 30719 8631 30725
rect 8573 30716 8585 30719
rect 7616 30688 8585 30716
rect 7616 30676 7622 30688
rect 8573 30685 8585 30688
rect 8619 30685 8631 30719
rect 8573 30679 8631 30685
rect 8662 30676 8668 30728
rect 8720 30716 8726 30728
rect 8772 30716 8800 30824
rect 8846 30812 8852 30824
rect 8904 30852 8910 30864
rect 9217 30855 9275 30861
rect 9217 30852 9229 30855
rect 8904 30824 9229 30852
rect 8904 30812 8910 30824
rect 9217 30821 9229 30824
rect 9263 30821 9275 30855
rect 9217 30815 9275 30821
rect 9306 30812 9312 30864
rect 9364 30852 9370 30864
rect 9737 30855 9795 30861
rect 9737 30852 9749 30855
rect 9364 30824 9749 30852
rect 9364 30812 9370 30824
rect 9737 30821 9749 30824
rect 9783 30821 9795 30855
rect 9737 30815 9795 30821
rect 9122 30744 9128 30796
rect 9180 30744 9186 30796
rect 9493 30787 9551 30793
rect 9493 30753 9505 30787
rect 9539 30784 9551 30787
rect 9876 30784 9904 30892
rect 9953 30855 10011 30861
rect 9953 30821 9965 30855
rect 9999 30852 10011 30855
rect 10226 30852 10232 30864
rect 9999 30824 10232 30852
rect 9999 30821 10011 30824
rect 9953 30815 10011 30821
rect 10226 30812 10232 30824
rect 10284 30812 10290 30864
rect 10428 30861 10456 30892
rect 10594 30880 10600 30932
rect 10652 30920 10658 30932
rect 11057 30923 11115 30929
rect 11057 30920 11069 30923
rect 10652 30892 11069 30920
rect 10652 30880 10658 30892
rect 11057 30889 11069 30892
rect 11103 30889 11115 30923
rect 11057 30883 11115 30889
rect 11606 30880 11612 30932
rect 11664 30920 11670 30932
rect 11885 30923 11943 30929
rect 11885 30920 11897 30923
rect 11664 30892 11897 30920
rect 11664 30880 11670 30892
rect 11885 30889 11897 30892
rect 11931 30889 11943 30923
rect 11885 30883 11943 30889
rect 10413 30855 10471 30861
rect 10413 30821 10425 30855
rect 10459 30852 10471 30855
rect 10686 30852 10692 30864
rect 10459 30824 10692 30852
rect 10459 30821 10471 30824
rect 10413 30815 10471 30821
rect 10686 30812 10692 30824
rect 10744 30812 10750 30864
rect 11698 30852 11704 30864
rect 10796 30824 11704 30852
rect 9539 30756 9904 30784
rect 9539 30753 9551 30756
rect 9493 30747 9551 30753
rect 10042 30744 10048 30796
rect 10100 30744 10106 30796
rect 10134 30744 10140 30796
rect 10192 30744 10198 30796
rect 10796 30793 10824 30824
rect 11698 30812 11704 30824
rect 11756 30812 11762 30864
rect 10781 30787 10839 30793
rect 10781 30753 10793 30787
rect 10827 30753 10839 30787
rect 10781 30747 10839 30753
rect 11241 30787 11299 30793
rect 11241 30753 11253 30787
rect 11287 30784 11299 30787
rect 11330 30784 11336 30796
rect 11287 30756 11336 30784
rect 11287 30753 11299 30756
rect 11241 30747 11299 30753
rect 11330 30744 11336 30756
rect 11388 30744 11394 30796
rect 11606 30744 11612 30796
rect 11664 30784 11670 30796
rect 11793 30787 11851 30793
rect 11793 30784 11805 30787
rect 11664 30756 11805 30784
rect 11664 30744 11670 30756
rect 11793 30753 11805 30756
rect 11839 30753 11851 30787
rect 11793 30747 11851 30753
rect 12161 30787 12219 30793
rect 12161 30753 12173 30787
rect 12207 30784 12219 30787
rect 12728 30784 12756 31096
rect 12207 30756 12756 30784
rect 12207 30753 12219 30756
rect 12161 30747 12219 30753
rect 9398 30716 9404 30728
rect 8720 30688 8800 30716
rect 8864 30688 9404 30716
rect 8720 30676 8726 30688
rect 7466 30648 7472 30660
rect 6052 30620 7052 30648
rect 7208 30620 7472 30648
rect 6052 30608 6058 30620
rect 14 30540 20 30592
rect 72 30580 78 30592
rect 566 30580 572 30592
rect 72 30552 572 30580
rect 72 30540 78 30552
rect 566 30540 572 30552
rect 624 30540 630 30592
rect 842 30540 848 30592
rect 900 30540 906 30592
rect 1854 30540 1860 30592
rect 1912 30580 1918 30592
rect 2685 30583 2743 30589
rect 2685 30580 2697 30583
rect 1912 30552 2697 30580
rect 1912 30540 1918 30552
rect 2685 30549 2697 30552
rect 2731 30549 2743 30583
rect 2685 30543 2743 30549
rect 2866 30540 2872 30592
rect 2924 30580 2930 30592
rect 3053 30583 3111 30589
rect 3053 30580 3065 30583
rect 2924 30552 3065 30580
rect 2924 30540 2930 30552
rect 3053 30549 3065 30552
rect 3099 30549 3111 30583
rect 3053 30543 3111 30549
rect 3421 30583 3479 30589
rect 3421 30549 3433 30583
rect 3467 30580 3479 30583
rect 4614 30580 4620 30592
rect 3467 30552 4620 30580
rect 3467 30549 3479 30552
rect 3421 30543 3479 30549
rect 4614 30540 4620 30552
rect 4672 30540 4678 30592
rect 4706 30540 4712 30592
rect 4764 30580 4770 30592
rect 5169 30583 5227 30589
rect 5169 30580 5181 30583
rect 4764 30552 5181 30580
rect 4764 30540 4770 30552
rect 5169 30549 5181 30552
rect 5215 30549 5227 30583
rect 5169 30543 5227 30549
rect 5534 30540 5540 30592
rect 5592 30540 5598 30592
rect 5718 30540 5724 30592
rect 5776 30580 5782 30592
rect 7024 30589 7052 30620
rect 7466 30608 7472 30620
rect 7524 30608 7530 30660
rect 7650 30608 7656 30660
rect 7708 30648 7714 30660
rect 7834 30648 7840 30660
rect 7708 30620 7840 30648
rect 7708 30608 7714 30620
rect 7834 30608 7840 30620
rect 7892 30648 7898 30660
rect 8864 30648 8892 30688
rect 9398 30676 9404 30688
rect 9456 30676 9462 30728
rect 9858 30676 9864 30728
rect 9916 30716 9922 30728
rect 10505 30719 10563 30725
rect 10505 30716 10517 30719
rect 9916 30688 10517 30716
rect 9916 30676 9922 30688
rect 10505 30685 10517 30688
rect 10551 30685 10563 30719
rect 10505 30679 10563 30685
rect 10689 30719 10747 30725
rect 10689 30685 10701 30719
rect 10735 30716 10747 30719
rect 10962 30716 10968 30728
rect 10735 30688 10968 30716
rect 10735 30685 10747 30688
rect 10689 30679 10747 30685
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 7892 30620 8892 30648
rect 7892 30608 7898 30620
rect 8938 30608 8944 30660
rect 8996 30648 9002 30660
rect 9582 30648 9588 30660
rect 8996 30620 9588 30648
rect 8996 30608 9002 30620
rect 9582 30608 9588 30620
rect 9640 30608 9646 30660
rect 11348 30648 11376 30744
rect 11422 30676 11428 30728
rect 11480 30676 11486 30728
rect 11882 30676 11888 30728
rect 11940 30676 11946 30728
rect 12342 30676 12348 30728
rect 12400 30716 12406 30728
rect 12618 30716 12624 30728
rect 12400 30688 12624 30716
rect 12400 30676 12406 30688
rect 12618 30676 12624 30688
rect 12676 30676 12682 30728
rect 12069 30651 12127 30657
rect 12069 30648 12081 30651
rect 11348 30620 12081 30648
rect 11900 30592 11928 30620
rect 12069 30617 12081 30620
rect 12115 30617 12127 30651
rect 12069 30611 12127 30617
rect 6181 30583 6239 30589
rect 6181 30580 6193 30583
rect 5776 30552 6193 30580
rect 5776 30540 5782 30552
rect 6181 30549 6193 30552
rect 6227 30549 6239 30583
rect 6181 30543 6239 30549
rect 7009 30583 7067 30589
rect 7009 30549 7021 30583
rect 7055 30549 7067 30583
rect 7009 30543 7067 30549
rect 8294 30540 8300 30592
rect 8352 30580 8358 30592
rect 9769 30583 9827 30589
rect 9769 30580 9781 30583
rect 8352 30552 9781 30580
rect 8352 30540 8358 30552
rect 9769 30549 9781 30552
rect 9815 30549 9827 30583
rect 9769 30543 9827 30549
rect 10410 30540 10416 30592
rect 10468 30580 10474 30592
rect 10597 30583 10655 30589
rect 10597 30580 10609 30583
rect 10468 30552 10609 30580
rect 10468 30540 10474 30552
rect 10597 30549 10609 30552
rect 10643 30549 10655 30583
rect 10597 30543 10655 30549
rect 11609 30583 11667 30589
rect 11609 30549 11621 30583
rect 11655 30580 11667 30583
rect 11698 30580 11704 30592
rect 11655 30552 11704 30580
rect 11655 30549 11667 30552
rect 11609 30543 11667 30549
rect 11698 30540 11704 30552
rect 11756 30540 11762 30592
rect 11882 30540 11888 30592
rect 11940 30540 11946 30592
rect 552 30490 12604 30512
rect 552 30438 3662 30490
rect 3714 30438 3726 30490
rect 3778 30438 3790 30490
rect 3842 30438 3854 30490
rect 3906 30438 3918 30490
rect 3970 30438 10062 30490
rect 10114 30438 10126 30490
rect 10178 30438 10190 30490
rect 10242 30438 10254 30490
rect 10306 30438 10318 30490
rect 10370 30438 12604 30490
rect 552 30416 12604 30438
rect 584 30348 1256 30376
rect 584 30320 612 30348
rect 566 30268 572 30320
rect 624 30268 630 30320
rect 658 30268 664 30320
rect 716 30308 722 30320
rect 1118 30308 1124 30320
rect 716 30280 1124 30308
rect 716 30268 722 30280
rect 1118 30268 1124 30280
rect 1176 30268 1182 30320
rect 1228 30308 1256 30348
rect 1946 30336 1952 30388
rect 2004 30376 2010 30388
rect 2041 30379 2099 30385
rect 2041 30376 2053 30379
rect 2004 30348 2053 30376
rect 2004 30336 2010 30348
rect 2041 30345 2053 30348
rect 2087 30345 2099 30379
rect 2869 30379 2927 30385
rect 2041 30339 2099 30345
rect 2332 30348 2820 30376
rect 2332 30308 2360 30348
rect 1228 30280 1348 30308
rect 1320 30240 1348 30280
rect 1964 30280 2360 30308
rect 1320 30212 1532 30240
rect 842 30132 848 30184
rect 900 30172 906 30184
rect 1213 30175 1271 30181
rect 1213 30172 1225 30175
rect 900 30144 1225 30172
rect 900 30132 906 30144
rect 1213 30141 1225 30144
rect 1259 30141 1271 30175
rect 1213 30135 1271 30141
rect 1305 30175 1363 30181
rect 1305 30141 1317 30175
rect 1351 30172 1363 30175
rect 1394 30172 1400 30184
rect 1351 30144 1400 30172
rect 1351 30141 1363 30144
rect 1305 30135 1363 30141
rect 1394 30132 1400 30144
rect 1452 30132 1458 30184
rect 1504 30181 1532 30212
rect 1489 30175 1547 30181
rect 1489 30141 1501 30175
rect 1535 30141 1547 30175
rect 1489 30135 1547 30141
rect 1118 30064 1124 30116
rect 1176 30104 1182 30116
rect 1964 30113 1992 30280
rect 2406 30268 2412 30320
rect 2464 30268 2470 30320
rect 2792 30308 2820 30348
rect 2869 30345 2881 30379
rect 2915 30376 2927 30379
rect 3786 30376 3792 30388
rect 2915 30348 3792 30376
rect 2915 30345 2927 30348
rect 2869 30339 2927 30345
rect 3786 30336 3792 30348
rect 3844 30336 3850 30388
rect 5445 30379 5503 30385
rect 3896 30348 4108 30376
rect 3896 30308 3924 30348
rect 2792 30280 3924 30308
rect 2424 30240 2452 30268
rect 2682 30240 2688 30252
rect 2424 30212 2688 30240
rect 2682 30200 2688 30212
rect 2740 30200 2746 30252
rect 3234 30200 3240 30252
rect 3292 30240 3298 30252
rect 3605 30248 3663 30249
rect 3353 30243 3663 30248
rect 3353 30240 3617 30243
rect 3292 30220 3617 30240
rect 3292 30212 3381 30220
rect 3292 30200 3298 30212
rect 3605 30209 3617 30220
rect 3651 30209 3663 30243
rect 4080 30240 4108 30348
rect 5445 30345 5457 30379
rect 5491 30376 5503 30379
rect 5626 30376 5632 30388
rect 5491 30348 5632 30376
rect 5491 30345 5503 30348
rect 5445 30339 5503 30345
rect 5626 30336 5632 30348
rect 5684 30336 5690 30388
rect 5905 30379 5963 30385
rect 5905 30345 5917 30379
rect 5951 30376 5963 30379
rect 5994 30376 6000 30388
rect 5951 30348 6000 30376
rect 5951 30345 5963 30348
rect 5905 30339 5963 30345
rect 5994 30336 6000 30348
rect 6052 30336 6058 30388
rect 6181 30379 6239 30385
rect 6181 30345 6193 30379
rect 6227 30376 6239 30379
rect 6546 30376 6552 30388
rect 6227 30348 6552 30376
rect 6227 30345 6239 30348
rect 6181 30339 6239 30345
rect 6546 30336 6552 30348
rect 6604 30336 6610 30388
rect 6730 30336 6736 30388
rect 6788 30336 6794 30388
rect 7006 30336 7012 30388
rect 7064 30376 7070 30388
rect 7101 30379 7159 30385
rect 7101 30376 7113 30379
rect 7064 30348 7113 30376
rect 7064 30336 7070 30348
rect 7101 30345 7113 30348
rect 7147 30345 7159 30379
rect 7101 30339 7159 30345
rect 7190 30336 7196 30388
rect 7248 30376 7254 30388
rect 7469 30379 7527 30385
rect 7469 30376 7481 30379
rect 7248 30348 7481 30376
rect 7248 30336 7254 30348
rect 7469 30345 7481 30348
rect 7515 30345 7527 30379
rect 7469 30339 7527 30345
rect 7834 30336 7840 30388
rect 7892 30376 7898 30388
rect 9490 30376 9496 30388
rect 7892 30348 9496 30376
rect 7892 30336 7898 30348
rect 9490 30336 9496 30348
rect 9548 30336 9554 30388
rect 10778 30376 10784 30388
rect 10520 30348 10784 30376
rect 4154 30268 4160 30320
rect 4212 30308 4218 30320
rect 4706 30308 4712 30320
rect 4212 30280 4712 30308
rect 4212 30268 4218 30280
rect 4706 30268 4712 30280
rect 4764 30268 4770 30320
rect 5810 30308 5816 30320
rect 5644 30280 5816 30308
rect 4080 30212 4660 30240
rect 3605 30203 3663 30209
rect 2225 30175 2283 30181
rect 2225 30141 2237 30175
rect 2271 30172 2283 30175
rect 2314 30172 2320 30184
rect 2271 30144 2320 30172
rect 2271 30141 2283 30144
rect 2225 30135 2283 30141
rect 2314 30132 2320 30144
rect 2372 30132 2378 30184
rect 2406 30132 2412 30184
rect 2464 30132 2470 30184
rect 2501 30175 2559 30181
rect 2501 30141 2513 30175
rect 2547 30172 2559 30175
rect 2590 30172 2596 30184
rect 2547 30144 2596 30172
rect 2547 30141 2559 30144
rect 2501 30135 2559 30141
rect 2590 30132 2596 30144
rect 2648 30132 2654 30184
rect 2961 30175 3019 30181
rect 2961 30172 2973 30175
rect 2792 30144 2973 30172
rect 2792 30116 2820 30144
rect 2961 30141 2973 30144
rect 3007 30141 3019 30175
rect 2961 30135 3019 30141
rect 3326 30132 3332 30184
rect 3384 30174 3390 30184
rect 3421 30175 3479 30181
rect 3421 30174 3433 30175
rect 3384 30146 3433 30174
rect 3384 30132 3390 30146
rect 3421 30141 3433 30146
rect 3467 30141 3479 30175
rect 3421 30135 3479 30141
rect 3513 30175 3571 30181
rect 3513 30141 3525 30175
rect 3559 30141 3571 30175
rect 3513 30135 3571 30141
rect 1949 30107 2007 30113
rect 1949 30104 1961 30107
rect 1176 30076 1961 30104
rect 1176 30064 1182 30076
rect 1949 30073 1961 30076
rect 1995 30073 2007 30107
rect 1949 30067 2007 30073
rect 2682 30064 2688 30116
rect 2740 30064 2746 30116
rect 2774 30064 2780 30116
rect 2832 30064 2838 30116
rect 1394 29996 1400 30048
rect 1452 30036 1458 30048
rect 3237 30039 3295 30045
rect 3237 30036 3249 30039
rect 1452 30008 3249 30036
rect 1452 29996 1458 30008
rect 3237 30005 3249 30008
rect 3283 30005 3295 30039
rect 3237 29999 3295 30005
rect 3418 29996 3424 30048
rect 3476 30036 3482 30048
rect 3528 30036 3556 30135
rect 3476 30008 3556 30036
rect 3620 30036 3648 30203
rect 3694 30132 3700 30184
rect 3752 30132 3758 30184
rect 3881 30175 3939 30181
rect 3881 30141 3893 30175
rect 3927 30174 3939 30175
rect 3927 30172 4007 30174
rect 4154 30172 4160 30184
rect 3927 30146 4160 30172
rect 3927 30141 3939 30146
rect 3979 30144 4160 30146
rect 3881 30135 3939 30141
rect 4154 30132 4160 30144
rect 4212 30132 4218 30184
rect 4249 30175 4307 30181
rect 4249 30141 4261 30175
rect 4295 30172 4307 30175
rect 4430 30172 4436 30184
rect 4295 30144 4436 30172
rect 4295 30141 4307 30144
rect 4249 30135 4307 30141
rect 4430 30132 4436 30144
rect 4488 30132 4494 30184
rect 4632 30181 4660 30212
rect 4617 30175 4675 30181
rect 4617 30141 4629 30175
rect 4663 30141 4675 30175
rect 4617 30135 4675 30141
rect 4982 30132 4988 30184
rect 5040 30172 5046 30184
rect 5169 30175 5227 30181
rect 5169 30172 5181 30175
rect 5040 30144 5181 30172
rect 5040 30132 5046 30144
rect 5169 30141 5181 30144
rect 5215 30141 5227 30175
rect 5169 30135 5227 30141
rect 5534 30132 5540 30184
rect 5592 30132 5598 30184
rect 5644 30181 5672 30280
rect 5810 30268 5816 30280
rect 5868 30268 5874 30320
rect 6914 30268 6920 30320
rect 6972 30308 6978 30320
rect 7653 30311 7711 30317
rect 7653 30308 7665 30311
rect 6972 30280 7665 30308
rect 6972 30268 6978 30280
rect 7653 30277 7665 30280
rect 7699 30277 7711 30311
rect 7653 30271 7711 30277
rect 8754 30268 8760 30320
rect 8812 30268 8818 30320
rect 9677 30311 9735 30317
rect 9677 30308 9689 30311
rect 9600 30280 9689 30308
rect 6730 30240 6736 30252
rect 6012 30212 6736 30240
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30141 5687 30175
rect 5629 30135 5687 30141
rect 5718 30132 5724 30184
rect 5776 30172 5782 30184
rect 6012 30181 6040 30212
rect 6730 30200 6736 30212
rect 6788 30200 6794 30252
rect 7926 30240 7932 30252
rect 7576 30212 7932 30240
rect 5813 30175 5871 30181
rect 5813 30172 5825 30175
rect 5776 30144 5825 30172
rect 5776 30132 5782 30144
rect 5813 30141 5825 30144
rect 5859 30141 5871 30175
rect 5813 30135 5871 30141
rect 5997 30175 6055 30181
rect 5997 30141 6009 30175
rect 6043 30141 6055 30175
rect 5997 30135 6055 30141
rect 6089 30175 6147 30181
rect 6089 30141 6101 30175
rect 6135 30141 6147 30175
rect 6089 30135 6147 30141
rect 3970 30064 3976 30116
rect 4028 30064 4034 30116
rect 5552 30104 5580 30132
rect 6104 30104 6132 30135
rect 6270 30132 6276 30184
rect 6328 30132 6334 30184
rect 6549 30175 6607 30181
rect 6549 30141 6561 30175
rect 6595 30172 6607 30175
rect 6638 30172 6644 30184
rect 6595 30144 6644 30172
rect 6595 30141 6607 30144
rect 6549 30135 6607 30141
rect 6638 30132 6644 30144
rect 6696 30132 6702 30184
rect 7098 30132 7104 30184
rect 7156 30132 7162 30184
rect 7282 30132 7288 30184
rect 7340 30172 7346 30184
rect 7576 30181 7604 30212
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 9398 30200 9404 30252
rect 9456 30200 9462 30252
rect 9490 30200 9496 30252
rect 9548 30240 9554 30252
rect 9600 30240 9628 30280
rect 9677 30277 9689 30280
rect 9723 30277 9735 30311
rect 9677 30271 9735 30277
rect 10226 30268 10232 30320
rect 10284 30268 10290 30320
rect 10520 30249 10548 30348
rect 10778 30336 10784 30348
rect 10836 30336 10842 30388
rect 10873 30379 10931 30385
rect 10873 30345 10885 30379
rect 10919 30376 10931 30379
rect 11606 30376 11612 30388
rect 10919 30348 11612 30376
rect 10919 30345 10931 30348
rect 10873 30339 10931 30345
rect 11606 30336 11612 30348
rect 11664 30336 11670 30388
rect 10594 30268 10600 30320
rect 10652 30308 10658 30320
rect 10689 30311 10747 30317
rect 10689 30308 10701 30311
rect 10652 30280 10701 30308
rect 10652 30268 10658 30280
rect 10689 30277 10701 30280
rect 10735 30277 10747 30311
rect 10689 30271 10747 30277
rect 10505 30243 10563 30249
rect 9548 30212 9628 30240
rect 9692 30212 10456 30240
rect 9548 30200 9554 30212
rect 7561 30175 7619 30181
rect 7561 30172 7573 30175
rect 7340 30144 7573 30172
rect 7340 30132 7346 30144
rect 7561 30141 7573 30144
rect 7607 30141 7619 30175
rect 7561 30135 7619 30141
rect 7745 30175 7803 30181
rect 7745 30141 7757 30175
rect 7791 30172 7803 30175
rect 7834 30172 7840 30184
rect 7791 30144 7840 30172
rect 7791 30141 7803 30144
rect 7745 30135 7803 30141
rect 4632 30076 5120 30104
rect 5552 30076 6132 30104
rect 6365 30107 6423 30113
rect 3878 30036 3884 30048
rect 3620 30008 3884 30036
rect 3476 29996 3482 30008
rect 3878 29996 3884 30008
rect 3936 29996 3942 30048
rect 3988 30036 4016 30064
rect 4632 30048 4660 30076
rect 4065 30039 4123 30045
rect 4065 30036 4077 30039
rect 3988 30008 4077 30036
rect 4065 30005 4077 30008
rect 4111 30005 4123 30039
rect 4065 29999 4123 30005
rect 4433 30039 4491 30045
rect 4433 30005 4445 30039
rect 4479 30036 4491 30039
rect 4522 30036 4528 30048
rect 4479 30008 4528 30036
rect 4479 30005 4491 30008
rect 4433 29999 4491 30005
rect 4522 29996 4528 30008
rect 4580 29996 4586 30048
rect 4614 29996 4620 30048
rect 4672 29996 4678 30048
rect 4798 29996 4804 30048
rect 4856 29996 4862 30048
rect 5092 30045 5120 30076
rect 6365 30073 6377 30107
rect 6411 30104 6423 30107
rect 6914 30104 6920 30116
rect 6411 30076 6920 30104
rect 6411 30073 6423 30076
rect 6365 30067 6423 30073
rect 6914 30064 6920 30076
rect 6972 30064 6978 30116
rect 7006 30064 7012 30116
rect 7064 30104 7070 30116
rect 7760 30104 7788 30135
rect 7834 30132 7840 30144
rect 7892 30132 7898 30184
rect 8110 30132 8116 30184
rect 8168 30132 8174 30184
rect 8389 30175 8447 30181
rect 8389 30172 8401 30175
rect 8220 30144 8401 30172
rect 7064 30076 7788 30104
rect 7064 30064 7070 30076
rect 5077 30039 5135 30045
rect 5077 30005 5089 30039
rect 5123 30005 5135 30039
rect 5077 29999 5135 30005
rect 5534 29996 5540 30048
rect 5592 30036 5598 30048
rect 7929 30039 7987 30045
rect 7929 30036 7941 30039
rect 5592 30008 7941 30036
rect 5592 29996 5598 30008
rect 7929 30005 7941 30008
rect 7975 30005 7987 30039
rect 8220 30036 8248 30144
rect 8389 30141 8401 30144
rect 8435 30141 8447 30175
rect 8389 30135 8447 30141
rect 8478 30132 8484 30184
rect 8536 30172 8542 30184
rect 8536 30144 8800 30172
rect 8536 30132 8542 30144
rect 8294 30064 8300 30116
rect 8352 30104 8358 30116
rect 8573 30107 8631 30113
rect 8573 30104 8585 30107
rect 8352 30076 8585 30104
rect 8352 30064 8358 30076
rect 8573 30073 8585 30076
rect 8619 30073 8631 30107
rect 8772 30104 8800 30144
rect 8846 30132 8852 30184
rect 8904 30132 8910 30184
rect 8938 30132 8944 30184
rect 8996 30132 9002 30184
rect 9033 30175 9091 30181
rect 9033 30141 9045 30175
rect 9079 30172 9091 30175
rect 9214 30172 9220 30184
rect 9079 30144 9220 30172
rect 9079 30141 9091 30144
rect 9033 30135 9091 30141
rect 9214 30132 9220 30144
rect 9272 30132 9278 30184
rect 9309 30175 9367 30181
rect 9309 30141 9321 30175
rect 9355 30172 9367 30175
rect 9692 30172 9720 30212
rect 9355 30144 9720 30172
rect 9769 30175 9827 30181
rect 9355 30141 9367 30144
rect 9309 30135 9367 30141
rect 9769 30141 9781 30175
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 9784 30104 9812 30135
rect 9950 30132 9956 30184
rect 10008 30172 10014 30184
rect 10321 30175 10379 30181
rect 10321 30172 10333 30175
rect 10008 30144 10333 30172
rect 10008 30132 10014 30144
rect 10321 30141 10333 30144
rect 10367 30141 10379 30175
rect 10428 30172 10456 30212
rect 10505 30209 10517 30243
rect 10551 30209 10563 30243
rect 10505 30203 10563 30209
rect 10612 30212 10916 30240
rect 10612 30172 10640 30212
rect 10428 30144 10640 30172
rect 10781 30175 10839 30181
rect 10321 30135 10379 30141
rect 10781 30141 10793 30175
rect 10827 30141 10839 30175
rect 10888 30172 10916 30212
rect 12250 30200 12256 30252
rect 12308 30200 12314 30252
rect 11698 30172 11704 30184
rect 10888 30144 11704 30172
rect 10781 30135 10839 30141
rect 10226 30104 10232 30116
rect 8772 30076 9812 30104
rect 9876 30076 10232 30104
rect 8573 30067 8631 30073
rect 8846 30036 8852 30048
rect 8220 30008 8852 30036
rect 7929 29999 7987 30005
rect 8846 29996 8852 30008
rect 8904 29996 8910 30048
rect 9214 29996 9220 30048
rect 9272 30036 9278 30048
rect 9876 30036 9904 30076
rect 10226 30064 10232 30076
rect 10284 30064 10290 30116
rect 9272 30008 9904 30036
rect 9272 29996 9278 30008
rect 9950 29996 9956 30048
rect 10008 29996 10014 30048
rect 10318 29996 10324 30048
rect 10376 30036 10382 30048
rect 10505 30039 10563 30045
rect 10505 30036 10517 30039
rect 10376 30008 10517 30036
rect 10376 29996 10382 30008
rect 10505 30005 10517 30008
rect 10551 30005 10563 30039
rect 10796 30036 10824 30135
rect 11698 30132 11704 30144
rect 11756 30132 11762 30184
rect 11514 30064 11520 30116
rect 11572 30104 11578 30116
rect 11986 30107 12044 30113
rect 11986 30104 11998 30107
rect 11572 30076 11998 30104
rect 11572 30064 11578 30076
rect 11986 30073 11998 30076
rect 12032 30073 12044 30107
rect 11986 30067 12044 30073
rect 12250 30036 12256 30048
rect 10796 30008 12256 30036
rect 10505 29999 10563 30005
rect 12250 29996 12256 30008
rect 12308 29996 12314 30048
rect 552 29946 12604 29968
rect 552 29894 4322 29946
rect 4374 29894 4386 29946
rect 4438 29894 4450 29946
rect 4502 29894 4514 29946
rect 4566 29894 4578 29946
rect 4630 29894 10722 29946
rect 10774 29894 10786 29946
rect 10838 29894 10850 29946
rect 10902 29894 10914 29946
rect 10966 29894 10978 29946
rect 11030 29894 12604 29946
rect 552 29872 12604 29894
rect 474 29792 480 29844
rect 532 29832 538 29844
rect 1029 29835 1087 29841
rect 1029 29832 1041 29835
rect 532 29804 1041 29832
rect 532 29792 538 29804
rect 1029 29801 1041 29804
rect 1075 29801 1087 29835
rect 1029 29795 1087 29801
rect 1486 29792 1492 29844
rect 1544 29792 1550 29844
rect 1762 29792 1768 29844
rect 1820 29792 1826 29844
rect 2130 29792 2136 29844
rect 2188 29832 2194 29844
rect 2314 29832 2320 29844
rect 2188 29804 2320 29832
rect 2188 29792 2194 29804
rect 2314 29792 2320 29804
rect 2372 29792 2378 29844
rect 2406 29792 2412 29844
rect 2464 29832 2470 29844
rect 2954 29835 3012 29841
rect 2954 29832 2966 29835
rect 2464 29804 2966 29832
rect 2464 29792 2470 29804
rect 2954 29801 2966 29804
rect 3000 29801 3012 29835
rect 2954 29795 3012 29801
rect 3421 29835 3479 29841
rect 3421 29801 3433 29835
rect 3467 29832 3479 29835
rect 3510 29832 3516 29844
rect 3467 29804 3516 29832
rect 3467 29801 3479 29804
rect 3421 29795 3479 29801
rect 3510 29792 3516 29804
rect 3568 29792 3574 29844
rect 3605 29835 3663 29841
rect 3605 29801 3617 29835
rect 3651 29832 3663 29835
rect 3786 29832 3792 29844
rect 3651 29804 3792 29832
rect 3651 29801 3663 29804
rect 3605 29795 3663 29801
rect 3786 29792 3792 29804
rect 3844 29792 3850 29844
rect 4154 29832 4160 29844
rect 3988 29804 4160 29832
rect 1670 29724 1676 29776
rect 1728 29724 1734 29776
rect 2682 29724 2688 29776
rect 2740 29724 2746 29776
rect 3056 29767 3114 29773
rect 3056 29733 3068 29767
rect 3102 29733 3114 29767
rect 3988 29764 4016 29804
rect 4154 29792 4160 29804
rect 4212 29792 4218 29844
rect 4982 29792 4988 29844
rect 5040 29792 5046 29844
rect 5442 29792 5448 29844
rect 5500 29792 5506 29844
rect 5718 29792 5724 29844
rect 5776 29832 5782 29844
rect 6086 29832 6092 29844
rect 5776 29804 6092 29832
rect 5776 29792 5782 29804
rect 6086 29792 6092 29804
rect 6144 29832 6150 29844
rect 6825 29835 6883 29841
rect 6825 29832 6837 29835
rect 6144 29804 6837 29832
rect 6144 29792 6150 29804
rect 6825 29801 6837 29804
rect 6871 29801 6883 29835
rect 6825 29795 6883 29801
rect 7098 29792 7104 29844
rect 7156 29832 7162 29844
rect 7650 29832 7656 29844
rect 7156 29804 7656 29832
rect 7156 29792 7162 29804
rect 7650 29792 7656 29804
rect 7708 29792 7714 29844
rect 8021 29835 8079 29841
rect 8021 29801 8033 29835
rect 8067 29832 8079 29835
rect 8110 29832 8116 29844
rect 8067 29804 8116 29832
rect 8067 29801 8079 29804
rect 8021 29795 8079 29801
rect 8110 29792 8116 29804
rect 8168 29792 8174 29844
rect 9398 29792 9404 29844
rect 9456 29832 9462 29844
rect 10045 29835 10103 29841
rect 10045 29832 10057 29835
rect 9456 29804 10057 29832
rect 9456 29792 9462 29804
rect 10045 29801 10057 29804
rect 10091 29801 10103 29835
rect 10045 29795 10103 29801
rect 10134 29792 10140 29844
rect 10192 29832 10198 29844
rect 10229 29835 10287 29841
rect 10229 29832 10241 29835
rect 10192 29804 10241 29832
rect 10192 29792 10198 29804
rect 10229 29801 10241 29804
rect 10275 29801 10287 29835
rect 10229 29795 10287 29801
rect 10318 29792 10324 29844
rect 10376 29832 10382 29844
rect 10502 29832 10508 29844
rect 10376 29804 10508 29832
rect 10376 29792 10382 29804
rect 10502 29792 10508 29804
rect 10560 29792 10566 29844
rect 11882 29841 11888 29844
rect 10965 29835 11023 29841
rect 10965 29801 10977 29835
rect 11011 29832 11023 29835
rect 11869 29835 11888 29841
rect 11011 29804 11192 29832
rect 11011 29801 11023 29804
rect 10965 29795 11023 29801
rect 3056 29727 3114 29733
rect 3528 29736 4016 29764
rect 1026 29656 1032 29708
rect 1084 29696 1090 29708
rect 1213 29699 1271 29705
rect 1213 29696 1225 29699
rect 1084 29668 1225 29696
rect 1084 29656 1090 29668
rect 1213 29665 1225 29668
rect 1259 29665 1271 29699
rect 1213 29659 1271 29665
rect 1394 29656 1400 29708
rect 1452 29656 1458 29708
rect 1949 29699 2007 29705
rect 1949 29665 1961 29699
rect 1995 29696 2007 29699
rect 1995 29668 2360 29696
rect 1995 29665 2007 29668
rect 1949 29659 2007 29665
rect 1762 29588 1768 29640
rect 1820 29628 1826 29640
rect 2133 29631 2191 29637
rect 2133 29628 2145 29631
rect 1820 29600 2145 29628
rect 1820 29588 1826 29600
rect 2133 29597 2145 29600
rect 2179 29628 2191 29631
rect 2225 29631 2283 29637
rect 2225 29628 2237 29631
rect 2179 29600 2237 29628
rect 2179 29597 2191 29600
rect 2133 29591 2191 29597
rect 2225 29597 2237 29600
rect 2271 29597 2283 29631
rect 2225 29591 2283 29597
rect 2332 29572 2360 29668
rect 2406 29656 2412 29708
rect 2464 29656 2470 29708
rect 2498 29656 2504 29708
rect 2556 29696 2562 29708
rect 2593 29699 2651 29705
rect 2593 29696 2605 29699
rect 2556 29668 2605 29696
rect 2556 29656 2562 29668
rect 2593 29665 2605 29668
rect 2639 29665 2651 29699
rect 2693 29696 2721 29724
rect 2777 29699 2835 29705
rect 2777 29696 2789 29699
rect 2693 29668 2789 29696
rect 2593 29659 2651 29665
rect 2777 29665 2789 29668
rect 2823 29665 2835 29699
rect 2777 29659 2835 29665
rect 2869 29699 2927 29705
rect 2869 29665 2881 29699
rect 2915 29665 2927 29699
rect 3068 29696 3096 29727
rect 3142 29696 3148 29708
rect 3068 29668 3148 29696
rect 2869 29659 2927 29665
rect 2682 29588 2688 29640
rect 2740 29588 2746 29640
rect 2884 29628 2912 29659
rect 3142 29656 3148 29668
rect 3200 29656 3206 29708
rect 3528 29696 3556 29736
rect 4062 29724 4068 29776
rect 4120 29764 4126 29776
rect 5460 29764 5488 29792
rect 6641 29767 6699 29773
rect 4120 29736 4752 29764
rect 4120 29724 4126 29736
rect 3252 29668 3556 29696
rect 3252 29628 3280 29668
rect 3602 29656 3608 29708
rect 3660 29696 3666 29708
rect 3697 29699 3755 29705
rect 3697 29696 3709 29699
rect 3660 29668 3709 29696
rect 3660 29656 3666 29668
rect 3697 29665 3709 29668
rect 3743 29665 3755 29699
rect 3697 29659 3755 29665
rect 3789 29699 3847 29705
rect 3789 29665 3801 29699
rect 3835 29665 3847 29699
rect 3789 29659 3847 29665
rect 3881 29699 3939 29705
rect 3881 29665 3893 29699
rect 3927 29696 3939 29699
rect 3927 29668 4016 29696
rect 3927 29665 3939 29668
rect 3881 29659 3939 29665
rect 2884 29600 3280 29628
rect 3418 29588 3424 29640
rect 3476 29588 3482 29640
rect 3804 29628 3832 29659
rect 3988 29640 4016 29668
rect 4246 29656 4252 29708
rect 4304 29656 4310 29708
rect 4724 29705 4752 29736
rect 4908 29736 6307 29764
rect 4908 29705 4936 29736
rect 4709 29699 4767 29705
rect 4709 29665 4721 29699
rect 4755 29665 4767 29699
rect 4709 29659 4767 29665
rect 4893 29699 4951 29705
rect 4893 29665 4905 29699
rect 4939 29665 4951 29699
rect 4893 29659 4951 29665
rect 5261 29699 5319 29705
rect 5261 29665 5273 29699
rect 5307 29696 5319 29699
rect 5350 29696 5356 29708
rect 5307 29668 5356 29696
rect 5307 29665 5319 29668
rect 5261 29659 5319 29665
rect 5350 29656 5356 29668
rect 5408 29656 5414 29708
rect 5445 29699 5503 29705
rect 5445 29665 5457 29699
rect 5491 29665 5503 29699
rect 5445 29659 5503 29665
rect 3804 29600 3912 29628
rect 1673 29563 1731 29569
rect 1673 29529 1685 29563
rect 1719 29560 1731 29563
rect 1854 29560 1860 29572
rect 1719 29532 1860 29560
rect 1719 29529 1731 29532
rect 1673 29523 1731 29529
rect 1854 29520 1860 29532
rect 1912 29520 1918 29572
rect 2314 29520 2320 29572
rect 2372 29520 2378 29572
rect 3789 29563 3847 29569
rect 3789 29560 3801 29563
rect 2792 29532 3801 29560
rect 382 29452 388 29504
rect 440 29492 446 29504
rect 2792 29492 2820 29532
rect 3789 29529 3801 29532
rect 3835 29529 3847 29563
rect 3884 29560 3912 29600
rect 3970 29588 3976 29640
rect 4028 29588 4034 29640
rect 4065 29631 4123 29637
rect 4065 29597 4077 29631
rect 4111 29628 4123 29631
rect 5074 29628 5080 29640
rect 4111 29600 5080 29628
rect 4111 29597 4123 29600
rect 4065 29591 4123 29597
rect 5074 29588 5080 29600
rect 5132 29588 5138 29640
rect 5460 29628 5488 29659
rect 5810 29656 5816 29708
rect 5868 29656 5874 29708
rect 5902 29656 5908 29708
rect 5960 29705 5966 29708
rect 5960 29699 6009 29705
rect 5960 29665 5963 29699
rect 5997 29696 6009 29699
rect 6086 29696 6092 29708
rect 5997 29668 6092 29696
rect 5997 29666 6010 29668
rect 5997 29665 6009 29666
rect 5960 29659 6009 29665
rect 5960 29656 5966 29659
rect 6086 29656 6092 29668
rect 6144 29656 6150 29708
rect 6178 29628 6184 29651
rect 5460 29600 6184 29628
rect 6178 29599 6184 29600
rect 6236 29599 6242 29651
rect 6279 29628 6307 29736
rect 6641 29733 6653 29767
rect 6687 29764 6699 29767
rect 7374 29764 7380 29776
rect 6687 29736 7380 29764
rect 6687 29733 6699 29736
rect 6641 29727 6699 29733
rect 7374 29724 7380 29736
rect 7432 29724 7438 29776
rect 8938 29724 8944 29776
rect 8996 29764 9002 29776
rect 10689 29767 10747 29773
rect 8996 29736 10272 29764
rect 8996 29724 9002 29736
rect 6546 29656 6552 29708
rect 6604 29696 6610 29708
rect 7009 29699 7067 29705
rect 7009 29696 7021 29699
rect 6604 29668 7021 29696
rect 6604 29656 6610 29668
rect 7009 29665 7021 29668
rect 7055 29665 7067 29699
rect 7653 29699 7711 29705
rect 7653 29696 7665 29699
rect 7009 29659 7067 29665
rect 7392 29668 7665 29696
rect 7392 29640 7420 29668
rect 7653 29665 7665 29668
rect 7699 29696 7711 29699
rect 7742 29696 7748 29708
rect 7699 29668 7748 29696
rect 7699 29665 7711 29668
rect 7653 29659 7711 29665
rect 7742 29656 7748 29668
rect 7800 29656 7806 29708
rect 7837 29699 7895 29705
rect 7837 29665 7849 29699
rect 7883 29696 7895 29699
rect 7926 29696 7932 29708
rect 7883 29668 7932 29696
rect 7883 29665 7895 29668
rect 7837 29659 7895 29665
rect 7926 29656 7932 29668
rect 7984 29656 7990 29708
rect 8110 29656 8116 29708
rect 8168 29696 8174 29708
rect 8478 29696 8484 29708
rect 8168 29668 8484 29696
rect 8168 29656 8174 29668
rect 8478 29656 8484 29668
rect 8536 29696 8542 29708
rect 9033 29699 9091 29705
rect 9033 29696 9045 29699
rect 8536 29668 9045 29696
rect 8536 29656 8542 29668
rect 9033 29665 9045 29668
rect 9079 29665 9091 29699
rect 9033 29659 9091 29665
rect 9214 29656 9220 29708
rect 9272 29656 9278 29708
rect 9674 29656 9680 29708
rect 9732 29696 9738 29708
rect 10137 29699 10195 29705
rect 10137 29696 10149 29699
rect 9732 29668 10149 29696
rect 9732 29656 9738 29668
rect 10137 29665 10149 29668
rect 10183 29665 10195 29699
rect 10244 29696 10272 29736
rect 10689 29733 10701 29767
rect 10735 29764 10747 29767
rect 10735 29736 11100 29764
rect 10735 29733 10747 29736
rect 10689 29727 10747 29733
rect 11072 29708 11100 29736
rect 10321 29699 10379 29705
rect 10321 29696 10333 29699
rect 10244 29668 10333 29696
rect 10137 29659 10195 29665
rect 10321 29665 10333 29668
rect 10367 29665 10379 29699
rect 10321 29659 10379 29665
rect 10594 29656 10600 29708
rect 10652 29656 10658 29708
rect 10781 29699 10839 29705
rect 10781 29665 10793 29699
rect 10827 29665 10839 29699
rect 10781 29659 10839 29665
rect 6914 29628 6920 29640
rect 6279 29600 6920 29628
rect 6914 29588 6920 29600
rect 6972 29588 6978 29640
rect 7193 29631 7251 29637
rect 7193 29597 7205 29631
rect 7239 29597 7251 29631
rect 7193 29591 7251 29597
rect 3884 29532 4200 29560
rect 3789 29523 3847 29529
rect 4172 29504 4200 29532
rect 4798 29520 4804 29572
rect 4856 29560 4862 29572
rect 5258 29560 5264 29572
rect 4856 29532 5264 29560
rect 4856 29520 4862 29532
rect 5258 29520 5264 29532
rect 5316 29560 5322 29572
rect 6181 29563 6239 29569
rect 6181 29560 6193 29563
rect 5316 29532 6193 29560
rect 5316 29520 5322 29532
rect 6181 29529 6193 29532
rect 6227 29529 6239 29563
rect 7208 29560 7236 29591
rect 7374 29588 7380 29640
rect 7432 29588 7438 29640
rect 7944 29628 7972 29656
rect 7944 29600 10180 29628
rect 7558 29560 7564 29572
rect 6181 29523 6239 29529
rect 6472 29532 7564 29560
rect 440 29464 2820 29492
rect 440 29452 446 29464
rect 2866 29452 2872 29504
rect 2924 29492 2930 29504
rect 3237 29495 3295 29501
rect 3237 29492 3249 29495
rect 2924 29464 3249 29492
rect 2924 29452 2930 29464
rect 3237 29461 3249 29464
rect 3283 29461 3295 29495
rect 3237 29455 3295 29461
rect 4154 29452 4160 29504
rect 4212 29492 4218 29504
rect 4341 29495 4399 29501
rect 4341 29492 4353 29495
rect 4212 29464 4353 29492
rect 4212 29452 4218 29464
rect 4341 29461 4353 29464
rect 4387 29461 4399 29495
rect 4341 29455 4399 29461
rect 4614 29452 4620 29504
rect 4672 29492 4678 29504
rect 4709 29495 4767 29501
rect 4709 29492 4721 29495
rect 4672 29464 4721 29492
rect 4672 29452 4678 29464
rect 4709 29461 4721 29464
rect 4755 29461 4767 29495
rect 4709 29455 4767 29461
rect 5350 29452 5356 29504
rect 5408 29452 5414 29504
rect 5626 29452 5632 29504
rect 5684 29492 5690 29504
rect 6086 29492 6092 29504
rect 5684 29464 6092 29492
rect 5684 29452 5690 29464
rect 6086 29452 6092 29464
rect 6144 29492 6150 29504
rect 6472 29492 6500 29532
rect 7558 29520 7564 29532
rect 7616 29520 7622 29572
rect 7834 29520 7840 29572
rect 7892 29560 7898 29572
rect 10152 29560 10180 29600
rect 10226 29588 10232 29640
rect 10284 29628 10290 29640
rect 10787 29628 10815 29659
rect 11054 29656 11060 29708
rect 11112 29656 11118 29708
rect 10284 29600 10815 29628
rect 11164 29628 11192 29804
rect 11869 29801 11881 29835
rect 11869 29795 11888 29801
rect 11882 29792 11888 29795
rect 11940 29792 11946 29844
rect 11698 29724 11704 29776
rect 11756 29764 11762 29776
rect 12069 29767 12127 29773
rect 12069 29764 12081 29767
rect 11756 29736 12081 29764
rect 11756 29724 11762 29736
rect 12069 29733 12081 29736
rect 12115 29733 12127 29767
rect 12069 29727 12127 29733
rect 11606 29656 11612 29708
rect 11664 29656 11670 29708
rect 12250 29628 12256 29640
rect 11164 29600 12256 29628
rect 10284 29588 10290 29600
rect 12250 29588 12256 29600
rect 12308 29588 12314 29640
rect 11330 29560 11336 29572
rect 7892 29532 9720 29560
rect 10152 29532 11336 29560
rect 7892 29520 7898 29532
rect 6144 29464 6500 29492
rect 6144 29452 6150 29464
rect 6546 29452 6552 29504
rect 6604 29452 6610 29504
rect 7653 29495 7711 29501
rect 7653 29461 7665 29495
rect 7699 29492 7711 29495
rect 8202 29492 8208 29504
rect 7699 29464 8208 29492
rect 7699 29461 7711 29464
rect 7653 29455 7711 29461
rect 8202 29452 8208 29464
rect 8260 29452 8266 29504
rect 9692 29492 9720 29532
rect 11330 29520 11336 29532
rect 11388 29560 11394 29572
rect 11388 29532 11928 29560
rect 11388 29520 11394 29532
rect 10778 29492 10784 29504
rect 9692 29464 10784 29492
rect 10778 29452 10784 29464
rect 10836 29452 10842 29504
rect 11606 29452 11612 29504
rect 11664 29492 11670 29504
rect 11900 29501 11928 29532
rect 11701 29495 11759 29501
rect 11701 29492 11713 29495
rect 11664 29464 11713 29492
rect 11664 29452 11670 29464
rect 11701 29461 11713 29464
rect 11747 29461 11759 29495
rect 11701 29455 11759 29461
rect 11885 29495 11943 29501
rect 11885 29461 11897 29495
rect 11931 29461 11943 29495
rect 11885 29455 11943 29461
rect 552 29402 12604 29424
rect 552 29350 3662 29402
rect 3714 29350 3726 29402
rect 3778 29350 3790 29402
rect 3842 29350 3854 29402
rect 3906 29350 3918 29402
rect 3970 29350 10062 29402
rect 10114 29350 10126 29402
rect 10178 29350 10190 29402
rect 10242 29350 10254 29402
rect 10306 29350 10318 29402
rect 10370 29350 12604 29402
rect 552 29328 12604 29350
rect 2314 29248 2320 29300
rect 2372 29248 2378 29300
rect 2866 29248 2872 29300
rect 2924 29288 2930 29300
rect 2961 29291 3019 29297
rect 2961 29288 2973 29291
rect 2924 29260 2973 29288
rect 2924 29248 2930 29260
rect 2961 29257 2973 29260
rect 3007 29257 3019 29291
rect 2961 29251 3019 29257
rect 4525 29291 4583 29297
rect 4525 29257 4537 29291
rect 4571 29288 4583 29291
rect 5074 29288 5080 29300
rect 4571 29260 5080 29288
rect 4571 29257 4583 29260
rect 4525 29251 4583 29257
rect 5074 29248 5080 29260
rect 5132 29248 5138 29300
rect 8754 29248 8760 29300
rect 8812 29288 8818 29300
rect 10413 29291 10471 29297
rect 8812 29260 10181 29288
rect 8812 29248 8818 29260
rect 1578 29180 1584 29232
rect 1636 29220 1642 29232
rect 1854 29220 1860 29232
rect 1636 29192 1860 29220
rect 1636 29180 1642 29192
rect 1854 29180 1860 29192
rect 1912 29180 1918 29232
rect 1946 29180 1952 29232
rect 2004 29220 2010 29232
rect 5534 29220 5540 29232
rect 2004 29192 2912 29220
rect 2004 29180 2010 29192
rect 934 29112 940 29164
rect 992 29152 998 29164
rect 1765 29155 1823 29161
rect 1765 29152 1777 29155
rect 992 29124 1777 29152
rect 992 29112 998 29124
rect 1765 29121 1777 29124
rect 1811 29121 1823 29155
rect 1765 29115 1823 29121
rect 1489 29087 1547 29093
rect 1489 29053 1501 29087
rect 1535 29084 1547 29087
rect 1578 29084 1584 29096
rect 1535 29056 1584 29084
rect 1535 29053 1547 29056
rect 1489 29047 1547 29053
rect 1578 29044 1584 29056
rect 1636 29044 1642 29096
rect 1673 29087 1731 29093
rect 1673 29053 1685 29087
rect 1719 29084 1731 29087
rect 1946 29084 1952 29096
rect 1719 29056 1952 29084
rect 1719 29053 1731 29056
rect 1673 29047 1731 29053
rect 1946 29044 1952 29056
rect 2004 29044 2010 29096
rect 2498 29044 2504 29096
rect 2556 29044 2562 29096
rect 2590 29044 2596 29096
rect 2648 29084 2654 29096
rect 2884 29093 2912 29192
rect 3528 29192 5540 29220
rect 2777 29087 2835 29093
rect 2777 29084 2789 29087
rect 2648 29056 2789 29084
rect 2648 29044 2654 29056
rect 2777 29053 2789 29056
rect 2823 29053 2835 29087
rect 2777 29047 2835 29053
rect 2869 29087 2927 29093
rect 2869 29053 2881 29087
rect 2915 29053 2927 29087
rect 2869 29047 2927 29053
rect 2958 29044 2964 29096
rect 3016 29084 3022 29096
rect 3053 29087 3111 29093
rect 3053 29084 3065 29087
rect 3016 29056 3065 29084
rect 3016 29044 3022 29056
rect 3053 29053 3065 29056
rect 3099 29053 3111 29087
rect 3053 29047 3111 29053
rect 3418 29044 3424 29096
rect 3476 29084 3482 29096
rect 3528 29093 3556 29192
rect 5534 29180 5540 29192
rect 5592 29180 5598 29232
rect 7745 29223 7803 29229
rect 7745 29189 7757 29223
rect 7791 29220 7803 29223
rect 8478 29220 8484 29232
rect 7791 29192 8484 29220
rect 7791 29189 7803 29192
rect 7745 29183 7803 29189
rect 4798 29112 4804 29164
rect 4856 29112 4862 29164
rect 5626 29112 5632 29164
rect 5684 29152 5690 29164
rect 5813 29155 5871 29161
rect 5813 29152 5825 29155
rect 5684 29124 5825 29152
rect 5684 29112 5690 29124
rect 5813 29121 5825 29124
rect 5859 29152 5871 29155
rect 5994 29152 6000 29164
rect 5859 29124 6000 29152
rect 5859 29121 5871 29124
rect 5813 29115 5871 29121
rect 5994 29112 6000 29124
rect 6052 29112 6058 29164
rect 6104 29124 6302 29152
rect 3513 29087 3571 29093
rect 3513 29084 3525 29087
rect 3476 29056 3525 29084
rect 3476 29044 3482 29056
rect 3513 29053 3525 29056
rect 3559 29053 3571 29087
rect 3513 29047 3571 29053
rect 3694 29044 3700 29096
rect 3752 29084 3758 29096
rect 3970 29084 3976 29096
rect 3752 29056 3976 29084
rect 3752 29044 3758 29056
rect 3970 29044 3976 29056
rect 4028 29044 4034 29096
rect 4433 29087 4491 29093
rect 4433 29053 4445 29087
rect 4479 29084 4491 29087
rect 4706 29084 4712 29096
rect 4479 29056 4712 29084
rect 4479 29053 4491 29056
rect 4433 29047 4491 29053
rect 4706 29044 4712 29056
rect 4764 29084 4770 29096
rect 5166 29084 5172 29096
rect 4764 29056 5172 29084
rect 4764 29044 4770 29056
rect 5166 29044 5172 29056
rect 5224 29084 5230 29096
rect 5261 29087 5319 29093
rect 5261 29084 5273 29087
rect 5224 29056 5273 29084
rect 5224 29044 5230 29056
rect 5261 29053 5273 29056
rect 5307 29053 5319 29087
rect 5261 29047 5319 29053
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29084 5411 29087
rect 5718 29084 5724 29096
rect 5399 29056 5724 29084
rect 5399 29053 5411 29056
rect 5353 29047 5411 29053
rect 5718 29044 5724 29056
rect 5776 29044 5782 29096
rect 6104 29093 6132 29124
rect 6089 29087 6147 29093
rect 6089 29053 6101 29087
rect 6135 29053 6147 29087
rect 6089 29047 6147 29053
rect 1026 28976 1032 29028
rect 1084 28976 1090 29028
rect 2682 28976 2688 29028
rect 2740 28976 2746 29028
rect 4893 29019 4951 29025
rect 4893 29016 4905 29019
rect 4172 28988 4905 29016
rect 3329 28951 3387 28957
rect 3329 28917 3341 28951
rect 3375 28948 3387 28951
rect 3418 28948 3424 28960
rect 3375 28920 3424 28948
rect 3375 28917 3387 28920
rect 3329 28911 3387 28917
rect 3418 28908 3424 28920
rect 3476 28948 3482 28960
rect 3878 28948 3884 28960
rect 3476 28920 3884 28948
rect 3476 28908 3482 28920
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 3970 28908 3976 28960
rect 4028 28948 4034 28960
rect 4172 28948 4200 28988
rect 4893 28985 4905 28988
rect 4939 28985 4951 29019
rect 4893 28979 4951 28985
rect 5442 28976 5448 29028
rect 5500 29016 5506 29028
rect 5997 29019 6055 29025
rect 5997 29016 6009 29019
rect 5500 28988 6009 29016
rect 5500 28976 5506 28988
rect 5997 28985 6009 28988
rect 6043 28985 6055 29019
rect 5997 28979 6055 28985
rect 4028 28920 4200 28948
rect 4028 28908 4034 28920
rect 4246 28908 4252 28960
rect 4304 28948 4310 28960
rect 5626 28948 5632 28960
rect 4304 28920 5632 28948
rect 4304 28908 4310 28920
rect 5626 28908 5632 28920
rect 5684 28908 5690 28960
rect 5718 28908 5724 28960
rect 5776 28948 5782 28960
rect 6104 28948 6132 29047
rect 6362 29044 6368 29096
rect 6420 29084 6426 29096
rect 6638 29084 6644 29096
rect 6420 29056 6644 29084
rect 6420 29044 6426 29056
rect 6638 29044 6644 29056
rect 6696 29084 6702 29096
rect 6733 29087 6791 29093
rect 6733 29084 6745 29087
rect 6696 29056 6745 29084
rect 6696 29044 6702 29056
rect 6733 29053 6745 29056
rect 6779 29053 6791 29087
rect 6733 29047 6791 29053
rect 6914 29044 6920 29096
rect 6972 29084 6978 29096
rect 7760 29084 7788 29183
rect 8478 29180 8484 29192
rect 8536 29180 8542 29232
rect 9953 29223 10011 29229
rect 9953 29220 9965 29223
rect 9508 29192 9965 29220
rect 9508 29164 9536 29192
rect 9953 29189 9965 29192
rect 9999 29189 10011 29223
rect 9953 29183 10011 29189
rect 8573 29155 8631 29161
rect 8573 29121 8585 29155
rect 8619 29152 8631 29155
rect 9030 29152 9036 29164
rect 8619 29124 9036 29152
rect 8619 29121 8631 29124
rect 8573 29115 8631 29121
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 9490 29112 9496 29164
rect 9548 29112 9554 29164
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 9861 29155 9919 29161
rect 9861 29152 9873 29155
rect 9732 29124 9873 29152
rect 9732 29112 9738 29124
rect 9861 29121 9873 29124
rect 9907 29121 9919 29155
rect 10153 29152 10181 29260
rect 10413 29257 10425 29291
rect 10459 29288 10471 29291
rect 10962 29288 10968 29300
rect 10459 29260 10968 29288
rect 10459 29257 10471 29260
rect 10413 29251 10471 29257
rect 10962 29248 10968 29260
rect 11020 29248 11026 29300
rect 11054 29248 11060 29300
rect 11112 29248 11118 29300
rect 11330 29248 11336 29300
rect 11388 29288 11394 29300
rect 11425 29291 11483 29297
rect 11425 29288 11437 29291
rect 11388 29260 11437 29288
rect 11388 29248 11394 29260
rect 11425 29257 11437 29260
rect 11471 29257 11483 29291
rect 11425 29251 11483 29257
rect 11514 29248 11520 29300
rect 11572 29248 11578 29300
rect 11885 29291 11943 29297
rect 11885 29257 11897 29291
rect 11931 29288 11943 29291
rect 11974 29288 11980 29300
rect 11931 29260 11980 29288
rect 11931 29257 11943 29260
rect 11885 29251 11943 29257
rect 11974 29248 11980 29260
rect 12032 29248 12038 29300
rect 10502 29180 10508 29232
rect 10560 29220 10566 29232
rect 12710 29220 12716 29232
rect 10560 29192 11560 29220
rect 10560 29180 10566 29192
rect 10153 29124 10732 29152
rect 9861 29115 9919 29121
rect 6972 29056 7788 29084
rect 8205 29087 8263 29093
rect 6972 29044 6978 29056
rect 8205 29053 8217 29087
rect 8251 29084 8263 29087
rect 8662 29084 8668 29096
rect 8251 29056 8668 29084
rect 8251 29053 8263 29056
rect 8205 29047 8263 29053
rect 8662 29044 8668 29056
rect 8720 29044 8726 29096
rect 8754 29044 8760 29096
rect 8812 29044 8818 29096
rect 9401 29087 9459 29093
rect 9401 29053 9413 29087
rect 9447 29084 9459 29087
rect 10321 29087 10379 29093
rect 10321 29084 10333 29087
rect 9447 29056 10333 29084
rect 9447 29053 9459 29056
rect 9401 29047 9459 29053
rect 10321 29053 10333 29056
rect 10367 29053 10379 29087
rect 10321 29047 10379 29053
rect 6457 29019 6515 29025
rect 6457 28985 6469 29019
rect 6503 29016 6515 29019
rect 6503 28988 6684 29016
rect 6503 28985 6515 28988
rect 6457 28979 6515 28985
rect 5776 28920 6132 28948
rect 6656 28948 6684 28988
rect 6822 28976 6828 29028
rect 6880 28976 6886 29028
rect 7098 28976 7104 29028
rect 7156 29016 7162 29028
rect 7193 29019 7251 29025
rect 7193 29016 7205 29019
rect 7156 28988 7205 29016
rect 7156 28976 7162 28988
rect 7193 28985 7205 28988
rect 7239 28985 7251 29019
rect 8018 29016 8024 29028
rect 7193 28979 7251 28985
rect 7484 28988 8024 29016
rect 7484 28960 7512 28988
rect 8018 28976 8024 28988
rect 8076 28976 8082 29028
rect 9416 29016 9444 29047
rect 10410 29044 10416 29096
rect 10468 29044 10474 29096
rect 10594 29044 10600 29096
rect 10652 29044 10658 29096
rect 10704 29093 10732 29124
rect 10778 29112 10784 29164
rect 10836 29112 10842 29164
rect 10980 29124 11284 29152
rect 10980 29093 11008 29124
rect 11256 29096 11284 29124
rect 10689 29087 10747 29093
rect 10689 29053 10701 29087
rect 10735 29053 10747 29087
rect 10689 29047 10747 29053
rect 10965 29087 11023 29093
rect 10965 29053 10977 29087
rect 11011 29053 11023 29087
rect 10965 29047 11023 29053
rect 11149 29087 11207 29093
rect 11149 29053 11161 29087
rect 11195 29053 11207 29087
rect 11149 29047 11207 29053
rect 8220 28988 9444 29016
rect 9508 28988 9996 29016
rect 8220 28960 8248 28988
rect 7282 28948 7288 28960
rect 6656 28920 7288 28948
rect 5776 28908 5782 28920
rect 7282 28908 7288 28920
rect 7340 28908 7346 28960
rect 7466 28908 7472 28960
rect 7524 28908 7530 28960
rect 7558 28908 7564 28960
rect 7616 28908 7622 28960
rect 7834 28908 7840 28960
rect 7892 28948 7898 28960
rect 8113 28951 8171 28957
rect 8113 28948 8125 28951
rect 7892 28920 8125 28948
rect 7892 28908 7898 28920
rect 8113 28917 8125 28920
rect 8159 28917 8171 28951
rect 8113 28911 8171 28917
rect 8202 28908 8208 28960
rect 8260 28908 8266 28960
rect 8478 28908 8484 28960
rect 8536 28948 8542 28960
rect 8665 28951 8723 28957
rect 8665 28948 8677 28951
rect 8536 28920 8677 28948
rect 8536 28908 8542 28920
rect 8665 28917 8677 28920
rect 8711 28917 8723 28951
rect 8665 28911 8723 28917
rect 8846 28908 8852 28960
rect 8904 28948 8910 28960
rect 9125 28951 9183 28957
rect 9125 28948 9137 28951
rect 8904 28920 9137 28948
rect 8904 28908 8910 28920
rect 9125 28917 9137 28920
rect 9171 28917 9183 28951
rect 9125 28911 9183 28917
rect 9306 28908 9312 28960
rect 9364 28948 9370 28960
rect 9508 28948 9536 28988
rect 9364 28920 9536 28948
rect 9769 28951 9827 28957
rect 9364 28908 9370 28920
rect 9769 28917 9781 28951
rect 9815 28948 9827 28951
rect 9858 28948 9864 28960
rect 9815 28920 9864 28948
rect 9815 28917 9827 28920
rect 9769 28911 9827 28917
rect 9858 28908 9864 28920
rect 9916 28908 9922 28960
rect 9968 28948 9996 28988
rect 10042 28976 10048 29028
rect 10100 29016 10106 29028
rect 10502 29016 10508 29028
rect 10100 28988 10508 29016
rect 10100 28976 10106 28988
rect 10502 28976 10508 28988
rect 10560 28976 10566 29028
rect 11164 29016 11192 29047
rect 11238 29044 11244 29096
rect 11296 29044 11302 29096
rect 11422 29044 11428 29096
rect 11480 29044 11486 29096
rect 11532 29093 11560 29192
rect 11808 29192 12716 29220
rect 11808 29161 11836 29192
rect 12710 29180 12716 29192
rect 12768 29180 12774 29232
rect 11793 29155 11851 29161
rect 11793 29121 11805 29155
rect 11839 29121 11851 29155
rect 11793 29115 11851 29121
rect 11977 29155 12035 29161
rect 11977 29121 11989 29155
rect 12023 29152 12035 29155
rect 12526 29152 12532 29164
rect 12023 29124 12532 29152
rect 12023 29121 12035 29124
rect 11977 29115 12035 29121
rect 12526 29112 12532 29124
rect 12584 29112 12590 29164
rect 11517 29087 11575 29093
rect 11517 29053 11529 29087
rect 11563 29053 11575 29087
rect 11517 29047 11575 29053
rect 11606 29044 11612 29096
rect 11664 29084 11670 29096
rect 11701 29087 11759 29093
rect 11701 29084 11713 29087
rect 11664 29056 11713 29084
rect 11664 29044 11670 29056
rect 11701 29053 11713 29056
rect 11747 29053 11759 29087
rect 12069 29087 12127 29093
rect 12069 29084 12081 29087
rect 11701 29047 11759 29053
rect 11900 29056 12081 29084
rect 11790 29016 11796 29028
rect 11164 28988 11796 29016
rect 11790 28976 11796 28988
rect 11848 28976 11854 29028
rect 11900 28948 11928 29056
rect 12069 29053 12081 29056
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 9968 28920 11928 28948
rect 552 28858 12604 28880
rect 552 28806 4322 28858
rect 4374 28806 4386 28858
rect 4438 28806 4450 28858
rect 4502 28806 4514 28858
rect 4566 28806 4578 28858
rect 4630 28806 10722 28858
rect 10774 28806 10786 28858
rect 10838 28806 10850 28858
rect 10902 28806 10914 28858
rect 10966 28806 10978 28858
rect 11030 28806 12604 28858
rect 552 28784 12604 28806
rect 2682 28704 2688 28756
rect 2740 28744 2746 28756
rect 3421 28747 3479 28753
rect 3421 28744 3433 28747
rect 2740 28716 3433 28744
rect 2740 28704 2746 28716
rect 3421 28713 3433 28716
rect 3467 28713 3479 28747
rect 3421 28707 3479 28713
rect 4246 28704 4252 28756
rect 4304 28704 4310 28756
rect 5353 28747 5411 28753
rect 5353 28713 5365 28747
rect 5399 28744 5411 28747
rect 5534 28744 5540 28756
rect 5399 28716 5540 28744
rect 5399 28713 5411 28716
rect 5353 28707 5411 28713
rect 5534 28704 5540 28716
rect 5592 28744 5598 28756
rect 5902 28744 5908 28756
rect 5592 28716 5908 28744
rect 5592 28704 5598 28716
rect 5902 28704 5908 28716
rect 5960 28704 5966 28756
rect 7558 28704 7564 28756
rect 7616 28744 7622 28756
rect 7616 28716 8524 28744
rect 7616 28704 7622 28716
rect 2314 28636 2320 28688
rect 2372 28636 2378 28688
rect 2424 28648 3004 28676
rect 290 28568 296 28620
rect 348 28608 354 28620
rect 1101 28611 1159 28617
rect 1101 28608 1113 28611
rect 348 28580 1113 28608
rect 348 28568 354 28580
rect 1101 28577 1113 28580
rect 1147 28608 1159 28611
rect 2424 28608 2452 28648
rect 2976 28617 3004 28648
rect 3142 28636 3148 28688
rect 3200 28676 3206 28688
rect 3970 28676 3976 28688
rect 3200 28648 3976 28676
rect 3200 28636 3206 28648
rect 3970 28636 3976 28648
rect 4028 28636 4034 28688
rect 4525 28679 4583 28685
rect 4525 28645 4537 28679
rect 4571 28676 4583 28679
rect 4706 28676 4712 28688
rect 4571 28648 4712 28676
rect 4571 28645 4583 28648
rect 4525 28639 4583 28645
rect 4706 28636 4712 28648
rect 4764 28636 4770 28688
rect 5166 28676 5172 28688
rect 4908 28648 5172 28676
rect 1147 28580 2452 28608
rect 2777 28611 2835 28617
rect 1147 28577 1159 28580
rect 1101 28571 1159 28577
rect 2777 28577 2789 28611
rect 2823 28577 2835 28611
rect 2777 28571 2835 28577
rect 2961 28611 3019 28617
rect 2961 28577 2973 28611
rect 3007 28577 3019 28611
rect 3234 28608 3240 28620
rect 2961 28571 3019 28577
rect 3160 28580 3240 28608
rect 842 28500 848 28552
rect 900 28500 906 28552
rect 1854 28500 1860 28552
rect 1912 28540 1918 28552
rect 2792 28540 2820 28571
rect 1912 28512 2820 28540
rect 3053 28543 3111 28549
rect 1912 28500 1918 28512
rect 3053 28509 3065 28543
rect 3099 28509 3111 28543
rect 3053 28503 3111 28509
rect 2225 28475 2283 28481
rect 2225 28441 2237 28475
rect 2271 28472 2283 28475
rect 3068 28472 3096 28503
rect 2271 28444 3096 28472
rect 2271 28441 2283 28444
rect 2225 28435 2283 28441
rect 2866 28364 2872 28416
rect 2924 28404 2930 28416
rect 3160 28404 3188 28580
rect 3234 28568 3240 28580
rect 3292 28608 3298 28620
rect 3605 28611 3663 28617
rect 3605 28608 3617 28611
rect 3292 28580 3617 28608
rect 3292 28568 3298 28580
rect 3605 28577 3617 28580
rect 3651 28577 3663 28611
rect 3605 28571 3663 28577
rect 3786 28568 3792 28620
rect 3844 28568 3850 28620
rect 3878 28568 3884 28620
rect 3936 28568 3942 28620
rect 4617 28611 4675 28617
rect 4080 28580 4568 28608
rect 3234 28432 3240 28484
rect 3292 28472 3298 28484
rect 3804 28472 3832 28568
rect 3970 28500 3976 28552
rect 4028 28540 4034 28552
rect 4080 28540 4108 28580
rect 4540 28552 4568 28580
rect 4617 28577 4629 28611
rect 4663 28608 4675 28611
rect 4908 28608 4936 28648
rect 5166 28636 5172 28648
rect 5224 28676 5230 28688
rect 5718 28676 5724 28688
rect 5224 28648 5724 28676
rect 5224 28636 5230 28648
rect 5718 28636 5724 28648
rect 5776 28636 5782 28688
rect 6181 28679 6239 28685
rect 6181 28645 6193 28679
rect 6227 28676 6239 28679
rect 6270 28676 6276 28688
rect 6227 28648 6276 28676
rect 6227 28645 6239 28648
rect 6181 28639 6239 28645
rect 6270 28636 6276 28648
rect 6328 28636 6334 28688
rect 4663 28580 4936 28608
rect 4985 28611 5043 28617
rect 4663 28577 4675 28580
rect 4617 28571 4675 28577
rect 4985 28577 4997 28611
rect 5031 28608 5043 28611
rect 5810 28608 5816 28620
rect 5031 28580 5816 28608
rect 5031 28577 5043 28580
rect 4985 28571 5043 28577
rect 5810 28568 5816 28580
rect 5868 28568 5874 28620
rect 5905 28611 5963 28617
rect 5905 28577 5917 28611
rect 5951 28577 5963 28611
rect 5905 28571 5963 28577
rect 4028 28526 4108 28540
rect 4028 28512 4094 28526
rect 4028 28500 4034 28512
rect 4522 28500 4528 28552
rect 4580 28500 4586 28552
rect 3292 28444 3832 28472
rect 5920 28472 5948 28571
rect 5994 28568 6000 28620
rect 6052 28608 6058 28620
rect 6638 28608 6644 28620
rect 6052 28580 6644 28608
rect 6052 28568 6058 28580
rect 6638 28568 6644 28580
rect 6696 28608 6702 28620
rect 6825 28611 6883 28617
rect 6825 28608 6837 28611
rect 6696 28580 6837 28608
rect 6696 28568 6702 28580
rect 6825 28577 6837 28580
rect 6871 28577 6883 28611
rect 6825 28571 6883 28577
rect 7193 28611 7251 28617
rect 7193 28577 7205 28611
rect 7239 28608 7251 28611
rect 7466 28608 7472 28620
rect 7239 28580 7472 28608
rect 7239 28577 7251 28580
rect 7193 28571 7251 28577
rect 7466 28568 7472 28580
rect 7524 28568 7530 28620
rect 7668 28617 7696 28716
rect 7742 28636 7748 28688
rect 7800 28676 7806 28688
rect 7800 28648 8432 28676
rect 7800 28636 7806 28648
rect 7653 28611 7711 28617
rect 7653 28577 7665 28611
rect 7699 28577 7711 28611
rect 7653 28571 7711 28577
rect 7834 28568 7840 28620
rect 7892 28608 7898 28620
rect 8128 28617 8156 28648
rect 7929 28611 7987 28617
rect 7929 28608 7941 28611
rect 7892 28580 7941 28608
rect 7892 28568 7898 28580
rect 7929 28577 7941 28580
rect 7975 28577 7987 28611
rect 7929 28571 7987 28577
rect 8113 28611 8171 28617
rect 8113 28577 8125 28611
rect 8159 28577 8171 28611
rect 8113 28571 8171 28577
rect 8202 28568 8208 28620
rect 8260 28568 8266 28620
rect 6546 28540 6552 28552
rect 6288 28512 6552 28540
rect 6288 28472 6316 28512
rect 6546 28500 6552 28512
rect 6604 28500 6610 28552
rect 7745 28543 7803 28549
rect 7745 28509 7757 28543
rect 7791 28540 7803 28543
rect 8220 28540 8248 28568
rect 7791 28512 8248 28540
rect 7791 28509 7803 28512
rect 7745 28503 7803 28509
rect 5920 28444 6316 28472
rect 3292 28432 3298 28444
rect 6362 28432 6368 28484
rect 6420 28472 6426 28484
rect 7469 28475 7527 28481
rect 7469 28472 7481 28475
rect 6420 28444 7481 28472
rect 6420 28432 6426 28444
rect 7469 28441 7481 28444
rect 7515 28441 7527 28475
rect 7469 28435 7527 28441
rect 7834 28432 7840 28484
rect 7892 28472 7898 28484
rect 8297 28475 8355 28481
rect 8297 28472 8309 28475
rect 7892 28444 8309 28472
rect 7892 28432 7898 28444
rect 8297 28441 8309 28444
rect 8343 28441 8355 28475
rect 8404 28472 8432 28648
rect 8496 28617 8524 28716
rect 8662 28704 8668 28756
rect 8720 28744 8726 28756
rect 9582 28744 9588 28756
rect 8720 28716 9588 28744
rect 8720 28704 8726 28716
rect 9582 28704 9588 28716
rect 9640 28744 9646 28756
rect 9769 28747 9827 28753
rect 9769 28744 9781 28747
rect 9640 28716 9781 28744
rect 9640 28704 9646 28716
rect 9769 28713 9781 28716
rect 9815 28713 9827 28747
rect 11698 28744 11704 28756
rect 9769 28707 9827 28713
rect 11440 28716 11704 28744
rect 8846 28636 8852 28688
rect 8904 28636 8910 28688
rect 8938 28636 8944 28688
rect 8996 28676 9002 28688
rect 10045 28679 10103 28685
rect 10045 28676 10057 28679
rect 8996 28648 10057 28676
rect 8996 28636 9002 28648
rect 10045 28645 10057 28648
rect 10091 28645 10103 28679
rect 10045 28639 10103 28645
rect 10597 28679 10655 28685
rect 10597 28645 10609 28679
rect 10643 28676 10655 28679
rect 11440 28676 11468 28716
rect 11698 28704 11704 28716
rect 11756 28744 11762 28756
rect 11974 28744 11980 28756
rect 11756 28716 11980 28744
rect 11756 28704 11762 28716
rect 11974 28704 11980 28716
rect 12032 28704 12038 28756
rect 12066 28704 12072 28756
rect 12124 28744 12130 28756
rect 12161 28747 12219 28753
rect 12161 28744 12173 28747
rect 12124 28716 12173 28744
rect 12124 28704 12130 28716
rect 12161 28713 12173 28716
rect 12207 28713 12219 28747
rect 12161 28707 12219 28713
rect 11885 28679 11943 28685
rect 11885 28676 11897 28679
rect 10643 28648 11468 28676
rect 10643 28645 10655 28648
rect 10597 28639 10655 28645
rect 8481 28611 8539 28617
rect 8481 28577 8493 28611
rect 8527 28608 8539 28611
rect 8754 28608 8760 28620
rect 8527 28580 8760 28608
rect 8527 28577 8539 28580
rect 8481 28571 8539 28577
rect 8754 28568 8760 28580
rect 8812 28568 8818 28620
rect 9122 28568 9128 28620
rect 9180 28568 9186 28620
rect 9306 28568 9312 28620
rect 9364 28568 9370 28620
rect 9585 28611 9643 28617
rect 9585 28577 9597 28611
rect 9631 28608 9643 28611
rect 9674 28608 9680 28620
rect 9631 28580 9680 28608
rect 9631 28577 9643 28580
rect 9585 28571 9643 28577
rect 9674 28568 9680 28580
rect 9732 28568 9738 28620
rect 9858 28568 9864 28620
rect 9916 28568 9922 28620
rect 10413 28611 10471 28617
rect 10413 28577 10425 28611
rect 10459 28577 10471 28611
rect 10413 28571 10471 28577
rect 10781 28611 10839 28617
rect 10781 28577 10793 28611
rect 10827 28608 10839 28611
rect 10965 28611 11023 28617
rect 10965 28608 10977 28611
rect 10827 28580 10977 28608
rect 10827 28577 10839 28580
rect 10781 28571 10839 28577
rect 10965 28577 10977 28580
rect 11011 28577 11023 28611
rect 10965 28571 11023 28577
rect 11149 28611 11207 28617
rect 11149 28577 11161 28611
rect 11195 28577 11207 28611
rect 11149 28571 11207 28577
rect 9766 28500 9772 28552
rect 9824 28540 9830 28552
rect 10428 28540 10456 28571
rect 9824 28512 10456 28540
rect 9824 28500 9830 28512
rect 9674 28472 9680 28484
rect 8404 28444 9680 28472
rect 8297 28435 8355 28441
rect 9674 28432 9680 28444
rect 9732 28472 9738 28484
rect 10229 28475 10287 28481
rect 10229 28472 10241 28475
rect 9732 28444 10241 28472
rect 9732 28432 9738 28444
rect 10229 28441 10241 28444
rect 10275 28441 10287 28475
rect 11164 28472 11192 28571
rect 11238 28568 11244 28620
rect 11296 28568 11302 28620
rect 11440 28617 11468 28648
rect 11716 28648 11897 28676
rect 11716 28617 11744 28648
rect 11885 28645 11897 28648
rect 11931 28645 11943 28679
rect 11885 28639 11943 28645
rect 11425 28611 11483 28617
rect 11425 28577 11437 28611
rect 11471 28577 11483 28611
rect 11425 28571 11483 28577
rect 11517 28611 11575 28617
rect 11517 28577 11529 28611
rect 11563 28577 11575 28611
rect 11517 28571 11575 28577
rect 11701 28611 11759 28617
rect 11701 28577 11713 28611
rect 11747 28577 11759 28611
rect 11701 28571 11759 28577
rect 11793 28611 11851 28617
rect 11793 28577 11805 28611
rect 11839 28577 11851 28611
rect 11793 28571 11851 28577
rect 11532 28472 11560 28571
rect 11808 28540 11836 28571
rect 12066 28568 12072 28620
rect 12124 28568 12130 28620
rect 12253 28611 12311 28617
rect 12253 28577 12265 28611
rect 12299 28608 12311 28611
rect 12434 28608 12440 28620
rect 12299 28580 12440 28608
rect 12299 28577 12311 28580
rect 12253 28571 12311 28577
rect 12434 28568 12440 28580
rect 12492 28568 12498 28620
rect 11882 28540 11888 28552
rect 11808 28512 11888 28540
rect 11882 28500 11888 28512
rect 11940 28500 11946 28552
rect 12066 28472 12072 28484
rect 11164 28444 11376 28472
rect 11532 28444 12072 28472
rect 10229 28435 10287 28441
rect 11348 28416 11376 28444
rect 12066 28432 12072 28444
rect 12124 28432 12130 28484
rect 2924 28376 3188 28404
rect 5537 28407 5595 28413
rect 2924 28364 2930 28376
rect 5537 28373 5549 28407
rect 5583 28404 5595 28407
rect 5902 28404 5908 28416
rect 5583 28376 5908 28404
rect 5583 28373 5595 28376
rect 5537 28367 5595 28373
rect 5902 28364 5908 28376
rect 5960 28364 5966 28416
rect 5997 28407 6055 28413
rect 5997 28373 6009 28407
rect 6043 28404 6055 28407
rect 6270 28404 6276 28416
rect 6043 28376 6276 28404
rect 6043 28373 6055 28376
rect 5997 28367 6055 28373
rect 6270 28364 6276 28376
rect 6328 28364 6334 28416
rect 8570 28364 8576 28416
rect 8628 28404 8634 28416
rect 8941 28407 8999 28413
rect 8941 28404 8953 28407
rect 8628 28376 8953 28404
rect 8628 28364 8634 28376
rect 8941 28373 8953 28376
rect 8987 28373 8999 28407
rect 8941 28367 8999 28373
rect 9125 28407 9183 28413
rect 9125 28373 9137 28407
rect 9171 28404 9183 28407
rect 9214 28404 9220 28416
rect 9171 28376 9220 28404
rect 9171 28373 9183 28376
rect 9125 28367 9183 28373
rect 9214 28364 9220 28376
rect 9272 28364 9278 28416
rect 9401 28407 9459 28413
rect 9401 28373 9413 28407
rect 9447 28404 9459 28407
rect 9950 28404 9956 28416
rect 9447 28376 9956 28404
rect 9447 28373 9459 28376
rect 9401 28367 9459 28373
rect 9950 28364 9956 28376
rect 10008 28364 10014 28416
rect 10410 28364 10416 28416
rect 10468 28404 10474 28416
rect 11057 28407 11115 28413
rect 11057 28404 11069 28407
rect 10468 28376 11069 28404
rect 10468 28364 10474 28376
rect 11057 28373 11069 28376
rect 11103 28373 11115 28407
rect 11057 28367 11115 28373
rect 11330 28364 11336 28416
rect 11388 28364 11394 28416
rect 11422 28364 11428 28416
rect 11480 28404 11486 28416
rect 11609 28407 11667 28413
rect 11609 28404 11621 28407
rect 11480 28376 11621 28404
rect 11480 28364 11486 28376
rect 11609 28373 11621 28376
rect 11655 28373 11667 28407
rect 11609 28367 11667 28373
rect 552 28314 12604 28336
rect 552 28262 3662 28314
rect 3714 28262 3726 28314
rect 3778 28262 3790 28314
rect 3842 28262 3854 28314
rect 3906 28262 3918 28314
rect 3970 28262 10062 28314
rect 10114 28262 10126 28314
rect 10178 28262 10190 28314
rect 10242 28262 10254 28314
rect 10306 28262 10318 28314
rect 10370 28262 12604 28314
rect 552 28240 12604 28262
rect 845 28203 903 28209
rect 845 28169 857 28203
rect 891 28200 903 28203
rect 934 28200 940 28212
rect 891 28172 940 28200
rect 891 28169 903 28172
rect 845 28163 903 28169
rect 934 28160 940 28172
rect 992 28160 998 28212
rect 2590 28160 2596 28212
rect 2648 28160 2654 28212
rect 4430 28160 4436 28212
rect 4488 28160 4494 28212
rect 6178 28160 6184 28212
rect 6236 28160 6242 28212
rect 7193 28203 7251 28209
rect 7193 28169 7205 28203
rect 7239 28200 7251 28203
rect 7834 28200 7840 28212
rect 7239 28172 7840 28200
rect 7239 28169 7251 28172
rect 7193 28163 7251 28169
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 7926 28160 7932 28212
rect 7984 28200 7990 28212
rect 9030 28200 9036 28212
rect 7984 28172 9036 28200
rect 7984 28160 7990 28172
rect 9030 28160 9036 28172
rect 9088 28160 9094 28212
rect 9214 28160 9220 28212
rect 9272 28160 9278 28212
rect 10594 28160 10600 28212
rect 10652 28200 10658 28212
rect 11698 28200 11704 28212
rect 10652 28172 11704 28200
rect 10652 28160 10658 28172
rect 11698 28160 11704 28172
rect 11756 28160 11762 28212
rect 4154 28092 4160 28144
rect 4212 28132 4218 28144
rect 6822 28132 6828 28144
rect 4212 28104 4292 28132
rect 4212 28092 4218 28104
rect 2222 28064 2228 28076
rect 2148 28036 2228 28064
rect 1394 27956 1400 28008
rect 1452 27996 1458 28008
rect 2148 27996 2176 28036
rect 2222 28024 2228 28036
rect 2280 28024 2286 28076
rect 3418 28064 3424 28076
rect 2976 28036 3424 28064
rect 2976 28005 3004 28036
rect 3418 28024 3424 28036
rect 3476 28064 3482 28076
rect 3513 28067 3571 28073
rect 3513 28064 3525 28067
rect 3476 28036 3525 28064
rect 3476 28024 3482 28036
rect 3513 28033 3525 28036
rect 3559 28033 3571 28067
rect 3513 28027 3571 28033
rect 1452 27968 2176 27996
rect 2777 27999 2835 28005
rect 1452 27956 1458 27968
rect 2777 27965 2789 27999
rect 2823 27965 2835 27999
rect 2777 27959 2835 27965
rect 2961 27999 3019 28005
rect 2961 27965 2973 27999
rect 3007 27965 3019 27999
rect 2961 27959 3019 27965
rect 1946 27888 1952 27940
rect 2004 27937 2010 27940
rect 2004 27928 2016 27937
rect 2792 27928 2820 27959
rect 3050 27956 3056 28008
rect 3108 27956 3114 28008
rect 3973 27999 4031 28005
rect 3973 27965 3985 27999
rect 4019 27996 4031 27999
rect 4154 27996 4160 28008
rect 4019 27968 4160 27996
rect 4019 27965 4031 27968
rect 3973 27959 4031 27965
rect 4154 27956 4160 27968
rect 4212 27956 4218 28008
rect 4264 28005 4292 28104
rect 6572 28104 6828 28132
rect 4614 28024 4620 28076
rect 4672 28024 4678 28076
rect 6572 28064 6600 28104
rect 5750 28036 6600 28064
rect 6638 28024 6644 28076
rect 6696 28024 6702 28076
rect 6748 28073 6776 28104
rect 6822 28092 6828 28104
rect 6880 28092 6886 28144
rect 11146 28132 11152 28144
rect 7208 28104 11152 28132
rect 6733 28067 6791 28073
rect 6733 28033 6745 28067
rect 6779 28033 6791 28067
rect 6733 28027 6791 28033
rect 4249 27999 4307 28005
rect 4249 27965 4261 27999
rect 4295 27965 4307 27999
rect 4249 27959 4307 27965
rect 3142 27928 3148 27940
rect 2004 27900 2049 27928
rect 2792 27900 3148 27928
rect 2004 27891 2016 27900
rect 2004 27888 2010 27891
rect 3142 27888 3148 27900
rect 3200 27888 3206 27940
rect 3881 27931 3939 27937
rect 3881 27897 3893 27931
rect 3927 27928 3939 27931
rect 4062 27928 4068 27940
rect 3927 27900 4068 27928
rect 3927 27897 3939 27900
rect 3881 27891 3939 27897
rect 4062 27888 4068 27900
rect 4120 27888 4126 27940
rect 3050 27820 3056 27872
rect 3108 27860 3114 27872
rect 3789 27863 3847 27869
rect 3789 27860 3801 27863
rect 3108 27832 3801 27860
rect 3108 27820 3114 27832
rect 3789 27829 3801 27832
rect 3835 27829 3847 27863
rect 4264 27860 4292 27959
rect 4430 27956 4436 28008
rect 4488 27956 4494 28008
rect 4632 27996 4660 28024
rect 5166 27996 5172 28008
rect 4632 27968 5172 27996
rect 5166 27956 5172 27968
rect 5224 27956 5230 28008
rect 5445 27999 5503 28005
rect 5445 27965 5457 27999
rect 5491 27996 5503 27999
rect 5534 27996 5540 28008
rect 5491 27968 5540 27996
rect 5491 27965 5503 27968
rect 5445 27959 5503 27965
rect 5534 27956 5540 27968
rect 5592 27956 5598 28008
rect 5810 27956 5816 28008
rect 5868 27996 5874 28008
rect 6549 27999 6607 28005
rect 6549 27996 6561 27999
rect 5868 27968 6561 27996
rect 5868 27956 5874 27968
rect 6549 27965 6561 27968
rect 6595 27965 6607 27999
rect 6549 27959 6607 27965
rect 4338 27888 4344 27940
rect 4396 27928 4402 27940
rect 4985 27931 5043 27937
rect 4985 27928 4997 27931
rect 4396 27900 4997 27928
rect 4396 27888 4402 27900
rect 4985 27897 4997 27900
rect 5031 27897 5043 27931
rect 4985 27891 5043 27897
rect 5077 27931 5135 27937
rect 5077 27897 5089 27931
rect 5123 27928 5135 27931
rect 5258 27928 5264 27940
rect 5123 27900 5264 27928
rect 5123 27897 5135 27900
rect 5077 27891 5135 27897
rect 5258 27888 5264 27900
rect 5316 27888 5322 27940
rect 5828 27928 5856 27956
rect 5736 27900 5856 27928
rect 4614 27860 4620 27872
rect 4264 27832 4620 27860
rect 3789 27823 3847 27829
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 4709 27863 4767 27869
rect 4709 27829 4721 27863
rect 4755 27860 4767 27863
rect 5736 27860 5764 27900
rect 4755 27832 5764 27860
rect 4755 27829 4767 27832
rect 4709 27823 4767 27829
rect 5810 27820 5816 27872
rect 5868 27820 5874 27872
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 5997 27863 6055 27869
rect 5997 27860 6009 27863
rect 5960 27832 6009 27860
rect 5960 27820 5966 27832
rect 5997 27829 6009 27832
rect 6043 27829 6055 27863
rect 6748 27860 6776 28027
rect 7009 27999 7067 28005
rect 7009 27965 7021 27999
rect 7055 27996 7067 27999
rect 7098 27996 7104 28008
rect 7055 27968 7104 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 7208 28005 7236 28104
rect 7852 28076 7880 28104
rect 11146 28092 11152 28104
rect 11204 28092 11210 28144
rect 7282 28024 7288 28076
rect 7340 28064 7346 28076
rect 7340 28036 7696 28064
rect 7340 28024 7346 28036
rect 7668 28005 7696 28036
rect 7834 28024 7840 28076
rect 7892 28024 7898 28076
rect 10045 28067 10103 28073
rect 10045 28064 10057 28067
rect 8956 28036 10057 28064
rect 7193 27999 7251 28005
rect 7193 27965 7205 27999
rect 7239 27965 7251 27999
rect 7193 27959 7251 27965
rect 7469 27999 7527 28005
rect 7469 27965 7481 27999
rect 7515 27965 7527 27999
rect 7469 27959 7527 27965
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27965 7711 27999
rect 7653 27959 7711 27965
rect 7745 27999 7803 28005
rect 7745 27965 7757 27999
rect 7791 27996 7803 27999
rect 8294 27996 8300 28008
rect 7791 27968 8300 27996
rect 7791 27965 7803 27968
rect 7745 27959 7803 27965
rect 7484 27928 7512 27959
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 8956 28005 8984 28036
rect 10045 28033 10057 28036
rect 10091 28033 10103 28067
rect 10045 28027 10103 28033
rect 10321 28067 10379 28073
rect 10321 28033 10333 28067
rect 10367 28064 10379 28067
rect 10965 28067 11023 28073
rect 10965 28064 10977 28067
rect 10367 28036 10977 28064
rect 10367 28033 10379 28036
rect 10321 28027 10379 28033
rect 10965 28033 10977 28036
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 11422 28024 11428 28076
rect 11480 28024 11486 28076
rect 8941 27999 8999 28005
rect 8941 27965 8953 27999
rect 8987 27965 8999 27999
rect 8941 27959 8999 27965
rect 9033 27999 9091 28005
rect 9033 27965 9045 27999
rect 9079 27965 9091 27999
rect 9033 27959 9091 27965
rect 7926 27928 7932 27940
rect 7484 27900 7932 27928
rect 7926 27888 7932 27900
rect 7984 27888 7990 27940
rect 8018 27888 8024 27940
rect 8076 27888 8082 27940
rect 8386 27888 8392 27940
rect 8444 27888 8450 27940
rect 8570 27888 8576 27940
rect 8628 27888 8634 27940
rect 9048 27928 9076 27959
rect 9214 27956 9220 28008
rect 9272 27996 9278 28008
rect 9309 27999 9367 28005
rect 9309 27996 9321 27999
rect 9272 27968 9321 27996
rect 9272 27956 9278 27968
rect 9309 27965 9321 27968
rect 9355 27965 9367 27999
rect 9585 27999 9643 28005
rect 9585 27996 9597 27999
rect 9309 27959 9367 27965
rect 9508 27968 9597 27996
rect 9401 27931 9459 27937
rect 9401 27928 9413 27931
rect 9048 27900 9413 27928
rect 9401 27897 9413 27900
rect 9447 27897 9459 27931
rect 9401 27891 9459 27897
rect 7190 27860 7196 27872
rect 6748 27832 7196 27860
rect 5997 27823 6055 27829
rect 7190 27820 7196 27832
rect 7248 27820 7254 27872
rect 7282 27820 7288 27872
rect 7340 27820 7346 27872
rect 8754 27820 8760 27872
rect 8812 27820 8818 27872
rect 9030 27820 9036 27872
rect 9088 27860 9094 27872
rect 9508 27860 9536 27968
rect 9585 27965 9597 27968
rect 9631 27965 9643 27999
rect 9585 27959 9643 27965
rect 9858 27956 9864 28008
rect 9916 27996 9922 28008
rect 9953 27999 10011 28005
rect 9953 27996 9965 27999
rect 9916 27968 9965 27996
rect 9916 27956 9922 27968
rect 9953 27965 9965 27968
rect 9999 27965 10011 27999
rect 9953 27959 10011 27965
rect 10137 27999 10195 28005
rect 10137 27965 10149 27999
rect 10183 27965 10195 27999
rect 10137 27959 10195 27965
rect 10152 27928 10180 27959
rect 10410 27956 10416 28008
rect 10468 27956 10474 28008
rect 10502 27956 10508 28008
rect 10560 27996 10566 28008
rect 10873 27999 10931 28005
rect 10873 27996 10885 27999
rect 10560 27968 10885 27996
rect 10560 27956 10566 27968
rect 10873 27965 10885 27968
rect 10919 27965 10931 27999
rect 10873 27959 10931 27965
rect 11057 27999 11115 28005
rect 11057 27965 11069 27999
rect 11103 27996 11115 27999
rect 11238 27996 11244 28008
rect 11103 27968 11244 27996
rect 11103 27965 11115 27968
rect 11057 27959 11115 27965
rect 11238 27956 11244 27968
rect 11296 27956 11302 28008
rect 11330 27956 11336 28008
rect 11388 27996 11394 28008
rect 11793 27999 11851 28005
rect 11793 27996 11805 27999
rect 11388 27968 11805 27996
rect 11388 27956 11394 27968
rect 11793 27965 11805 27968
rect 11839 27965 11851 27999
rect 11793 27959 11851 27965
rect 11882 27956 11888 28008
rect 11940 27956 11946 28008
rect 12066 27956 12072 28008
rect 12124 27956 12130 28008
rect 9784 27900 10180 27928
rect 9088 27832 9536 27860
rect 9088 27820 9094 27832
rect 9582 27820 9588 27872
rect 9640 27860 9646 27872
rect 9784 27869 9812 27900
rect 9769 27863 9827 27869
rect 9769 27860 9781 27863
rect 9640 27832 9781 27860
rect 9640 27820 9646 27832
rect 9769 27829 9781 27832
rect 9815 27829 9827 27863
rect 9769 27823 9827 27829
rect 10594 27820 10600 27872
rect 10652 27860 10658 27872
rect 10781 27863 10839 27869
rect 10781 27860 10793 27863
rect 10652 27832 10793 27860
rect 10652 27820 10658 27832
rect 10781 27829 10793 27832
rect 10827 27829 10839 27863
rect 10781 27823 10839 27829
rect 11701 27863 11759 27869
rect 11701 27829 11713 27863
rect 11747 27860 11759 27863
rect 11790 27860 11796 27872
rect 11747 27832 11796 27860
rect 11747 27829 11759 27832
rect 11701 27823 11759 27829
rect 11790 27820 11796 27832
rect 11848 27820 11854 27872
rect 12250 27820 12256 27872
rect 12308 27820 12314 27872
rect 552 27770 12604 27792
rect 552 27718 4322 27770
rect 4374 27718 4386 27770
rect 4438 27718 4450 27770
rect 4502 27718 4514 27770
rect 4566 27718 4578 27770
rect 4630 27718 10722 27770
rect 10774 27718 10786 27770
rect 10838 27718 10850 27770
rect 10902 27718 10914 27770
rect 10966 27718 10978 27770
rect 11030 27718 12604 27770
rect 552 27696 12604 27718
rect 2498 27616 2504 27668
rect 2556 27616 2562 27668
rect 3418 27616 3424 27668
rect 3476 27656 3482 27668
rect 3605 27659 3663 27665
rect 3605 27656 3617 27659
rect 3476 27628 3617 27656
rect 3476 27616 3482 27628
rect 3605 27625 3617 27628
rect 3651 27625 3663 27659
rect 3605 27619 3663 27625
rect 4338 27616 4344 27668
rect 4396 27656 4402 27668
rect 4798 27656 4804 27668
rect 4396 27628 4804 27656
rect 4396 27616 4402 27628
rect 4798 27616 4804 27628
rect 4856 27616 4862 27668
rect 5258 27616 5264 27668
rect 5316 27656 5322 27668
rect 5718 27656 5724 27668
rect 5316 27628 5724 27656
rect 5316 27616 5322 27628
rect 5718 27616 5724 27628
rect 5776 27616 5782 27668
rect 6454 27616 6460 27668
rect 6512 27656 6518 27668
rect 7006 27656 7012 27668
rect 6512 27628 7012 27656
rect 6512 27616 6518 27628
rect 7006 27616 7012 27628
rect 7064 27616 7070 27668
rect 8113 27659 8171 27665
rect 8113 27625 8125 27659
rect 8159 27625 8171 27659
rect 8113 27619 8171 27625
rect 8573 27659 8631 27665
rect 8573 27625 8585 27659
rect 8619 27656 8631 27659
rect 8754 27656 8760 27668
rect 8619 27628 8760 27656
rect 8619 27625 8631 27628
rect 8573 27619 8631 27625
rect 2133 27591 2191 27597
rect 2133 27588 2145 27591
rect 1320 27560 2145 27588
rect 1320 27529 1348 27560
rect 2133 27557 2145 27560
rect 2179 27557 2191 27591
rect 2516 27588 2544 27616
rect 3237 27591 3295 27597
rect 3237 27588 3249 27591
rect 2133 27551 2191 27557
rect 2332 27560 2544 27588
rect 2608 27560 3249 27588
rect 1305 27523 1363 27529
rect 1305 27489 1317 27523
rect 1351 27489 1363 27523
rect 1305 27483 1363 27489
rect 1489 27523 1547 27529
rect 1489 27489 1501 27523
rect 1535 27520 1547 27523
rect 1762 27520 1768 27532
rect 1535 27492 1768 27520
rect 1535 27489 1547 27492
rect 1489 27483 1547 27489
rect 1762 27480 1768 27492
rect 1820 27480 1826 27532
rect 2332 27529 2360 27560
rect 2608 27529 2636 27560
rect 3237 27557 3249 27560
rect 3283 27557 3295 27591
rect 3237 27551 3295 27557
rect 4154 27548 4160 27600
rect 4212 27588 4218 27600
rect 8128 27588 8156 27619
rect 8754 27616 8760 27628
rect 8812 27616 8818 27668
rect 9306 27616 9312 27668
rect 9364 27656 9370 27668
rect 9364 27628 9444 27656
rect 9364 27616 9370 27628
rect 4212 27560 8156 27588
rect 8481 27591 8539 27597
rect 4212 27548 4218 27560
rect 8481 27557 8493 27591
rect 8527 27588 8539 27591
rect 8662 27588 8668 27600
rect 8527 27560 8668 27588
rect 8527 27557 8539 27560
rect 8481 27551 8539 27557
rect 8662 27548 8668 27560
rect 8720 27548 8726 27600
rect 8938 27548 8944 27600
rect 8996 27588 9002 27600
rect 8996 27560 9352 27588
rect 8996 27548 9002 27560
rect 2041 27523 2099 27529
rect 2041 27489 2053 27523
rect 2087 27520 2099 27523
rect 2317 27523 2375 27529
rect 2317 27520 2329 27523
rect 2087 27492 2329 27520
rect 2087 27489 2099 27492
rect 2041 27483 2099 27489
rect 2317 27489 2329 27492
rect 2363 27489 2375 27523
rect 2317 27483 2375 27489
rect 2501 27523 2559 27529
rect 2501 27489 2513 27523
rect 2547 27489 2559 27523
rect 2501 27483 2559 27489
rect 2593 27523 2651 27529
rect 2593 27489 2605 27523
rect 2639 27489 2651 27523
rect 2593 27483 2651 27489
rect 2516 27452 2544 27483
rect 2682 27480 2688 27532
rect 2740 27520 2746 27532
rect 2869 27523 2927 27529
rect 2869 27520 2881 27523
rect 2740 27492 2881 27520
rect 2740 27480 2746 27492
rect 2869 27489 2881 27492
rect 2915 27489 2927 27523
rect 2869 27483 2927 27489
rect 3050 27480 3056 27532
rect 3108 27480 3114 27532
rect 3142 27480 3148 27532
rect 3200 27520 3206 27532
rect 3418 27520 3424 27532
rect 3200 27492 3424 27520
rect 3200 27480 3206 27492
rect 3418 27480 3424 27492
rect 3476 27480 3482 27532
rect 3697 27523 3755 27529
rect 3697 27489 3709 27523
rect 3743 27489 3755 27523
rect 3697 27483 3755 27489
rect 2700 27452 2728 27480
rect 2516 27424 2728 27452
rect 3712 27452 3740 27483
rect 4338 27480 4344 27532
rect 4396 27480 4402 27532
rect 4525 27523 4583 27529
rect 4525 27489 4537 27523
rect 4571 27520 4583 27523
rect 4890 27520 4896 27532
rect 4571 27492 4896 27520
rect 4571 27489 4583 27492
rect 4525 27483 4583 27489
rect 4890 27480 4896 27492
rect 4948 27480 4954 27532
rect 5074 27480 5080 27532
rect 5132 27480 5138 27532
rect 5166 27480 5172 27532
rect 5224 27480 5230 27532
rect 5350 27480 5356 27532
rect 5408 27480 5414 27532
rect 6086 27480 6092 27532
rect 6144 27480 6150 27532
rect 6822 27480 6828 27532
rect 6880 27480 6886 27532
rect 7006 27480 7012 27532
rect 7064 27480 7070 27532
rect 7282 27480 7288 27532
rect 7340 27520 7346 27532
rect 7377 27523 7435 27529
rect 7377 27520 7389 27523
rect 7340 27492 7389 27520
rect 7340 27480 7346 27492
rect 7377 27489 7389 27492
rect 7423 27489 7435 27523
rect 8021 27523 8079 27529
rect 7377 27483 7435 27489
rect 7576 27492 7880 27520
rect 7576 27464 7604 27492
rect 7193 27455 7251 27461
rect 7193 27452 7205 27455
rect 3712 27424 7205 27452
rect 7193 27421 7205 27424
rect 7239 27421 7251 27455
rect 7193 27415 7251 27421
rect 7469 27455 7527 27461
rect 7469 27421 7481 27455
rect 7515 27421 7527 27455
rect 7469 27415 7527 27421
rect 1949 27387 2007 27393
rect 1949 27353 1961 27387
rect 1995 27384 2007 27387
rect 2685 27387 2743 27393
rect 2685 27384 2697 27387
rect 1995 27356 2697 27384
rect 1995 27353 2007 27356
rect 1949 27347 2007 27353
rect 2685 27353 2697 27356
rect 2731 27353 2743 27387
rect 2685 27347 2743 27353
rect 4614 27344 4620 27396
rect 4672 27384 4678 27396
rect 4709 27387 4767 27393
rect 4709 27384 4721 27387
rect 4672 27356 4721 27384
rect 4672 27344 4678 27356
rect 4709 27353 4721 27356
rect 4755 27353 4767 27387
rect 4709 27347 4767 27353
rect 4890 27344 4896 27396
rect 4948 27344 4954 27396
rect 5261 27387 5319 27393
rect 5261 27353 5273 27387
rect 5307 27384 5319 27387
rect 5442 27384 5448 27396
rect 5307 27356 5448 27384
rect 5307 27353 5319 27356
rect 5261 27347 5319 27353
rect 5442 27344 5448 27356
rect 5500 27344 5506 27396
rect 7484 27384 7512 27415
rect 7558 27412 7564 27464
rect 7616 27412 7622 27464
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 7742 27452 7748 27464
rect 7699 27424 7748 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 7742 27412 7748 27424
rect 7800 27412 7806 27464
rect 7852 27452 7880 27492
rect 8021 27489 8033 27523
rect 8067 27520 8079 27523
rect 8110 27520 8116 27532
rect 8067 27492 8116 27520
rect 8067 27489 8079 27492
rect 8021 27483 8079 27489
rect 8110 27480 8116 27492
rect 8168 27480 8174 27532
rect 8202 27480 8208 27532
rect 8260 27520 8266 27532
rect 9324 27529 9352 27560
rect 9416 27529 9444 27628
rect 9490 27616 9496 27668
rect 9548 27616 9554 27668
rect 9582 27616 9588 27668
rect 9640 27656 9646 27668
rect 9640 27616 9674 27656
rect 10226 27616 10232 27668
rect 10284 27656 10290 27668
rect 11057 27659 11115 27665
rect 10284 27628 11008 27656
rect 10284 27616 10290 27628
rect 9508 27588 9536 27616
rect 9646 27588 9674 27616
rect 9861 27591 9919 27597
rect 9861 27588 9873 27591
rect 9508 27560 9608 27588
rect 9646 27560 9873 27588
rect 9580 27529 9608 27560
rect 9861 27557 9873 27560
rect 9907 27557 9919 27591
rect 9861 27551 9919 27557
rect 10594 27548 10600 27600
rect 10652 27588 10658 27600
rect 10652 27560 10824 27588
rect 10652 27548 10658 27560
rect 9309 27523 9367 27529
rect 8260 27492 9260 27520
rect 8260 27480 8266 27492
rect 9232 27464 9260 27492
rect 9309 27489 9321 27523
rect 9355 27489 9367 27523
rect 9309 27483 9367 27489
rect 9401 27523 9459 27529
rect 9401 27489 9413 27523
rect 9447 27489 9459 27523
rect 9580 27523 9643 27529
rect 9580 27492 9597 27523
rect 9401 27483 9459 27489
rect 9585 27489 9597 27492
rect 9631 27489 9643 27523
rect 9585 27483 9643 27489
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 10796 27529 10824 27560
rect 10980 27529 11008 27628
rect 11057 27625 11069 27659
rect 11103 27656 11115 27659
rect 11882 27656 11888 27668
rect 11103 27628 11888 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 11882 27616 11888 27628
rect 11940 27616 11946 27668
rect 11977 27591 12035 27597
rect 11977 27588 11989 27591
rect 11440 27560 11989 27588
rect 10505 27523 10563 27529
rect 10505 27520 10517 27523
rect 9732 27492 10517 27520
rect 9732 27480 9738 27492
rect 10505 27489 10517 27492
rect 10551 27489 10563 27523
rect 10505 27483 10563 27489
rect 10689 27523 10747 27529
rect 10689 27489 10701 27523
rect 10735 27489 10747 27523
rect 10689 27483 10747 27489
rect 10781 27523 10839 27529
rect 10781 27489 10793 27523
rect 10827 27489 10839 27523
rect 10781 27483 10839 27489
rect 10965 27523 11023 27529
rect 10965 27489 10977 27523
rect 11011 27520 11023 27523
rect 11011 27492 11100 27520
rect 11011 27489 11023 27492
rect 10965 27483 11023 27489
rect 8665 27455 8723 27461
rect 8665 27452 8677 27455
rect 7852 27424 8677 27452
rect 8665 27421 8677 27424
rect 8711 27421 8723 27455
rect 8665 27415 8723 27421
rect 9214 27412 9220 27464
rect 9272 27452 9278 27464
rect 10321 27455 10379 27461
rect 10321 27452 10333 27455
rect 9272 27424 10333 27452
rect 9272 27412 9278 27424
rect 10321 27421 10333 27424
rect 10367 27421 10379 27455
rect 10321 27415 10379 27421
rect 9125 27387 9183 27393
rect 9125 27384 9137 27387
rect 7484 27356 9137 27384
rect 9125 27353 9137 27356
rect 9171 27353 9183 27387
rect 9125 27347 9183 27353
rect 9306 27344 9312 27396
rect 9364 27384 9370 27396
rect 10410 27384 10416 27396
rect 9364 27356 10416 27384
rect 9364 27344 9370 27356
rect 10410 27344 10416 27356
rect 10468 27384 10474 27396
rect 10704 27384 10732 27483
rect 11072 27464 11100 27492
rect 11146 27480 11152 27532
rect 11204 27480 11210 27532
rect 11238 27480 11244 27532
rect 11296 27520 11302 27532
rect 11440 27529 11468 27560
rect 11977 27557 11989 27560
rect 12023 27557 12035 27591
rect 11977 27551 12035 27557
rect 11425 27523 11483 27529
rect 11425 27520 11437 27523
rect 11296 27492 11437 27520
rect 11296 27480 11302 27492
rect 11425 27489 11437 27492
rect 11471 27489 11483 27523
rect 11425 27483 11483 27489
rect 11698 27480 11704 27532
rect 11756 27520 11762 27532
rect 11882 27520 11888 27532
rect 11756 27492 11888 27520
rect 11756 27480 11762 27492
rect 11882 27480 11888 27492
rect 11940 27480 11946 27532
rect 12069 27523 12127 27529
rect 12069 27489 12081 27523
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 11054 27412 11060 27464
rect 11112 27412 11118 27464
rect 11514 27412 11520 27464
rect 11572 27412 11578 27464
rect 11606 27412 11612 27464
rect 11664 27452 11670 27464
rect 12084 27452 12112 27483
rect 11664 27424 12112 27452
rect 11664 27412 11670 27424
rect 10468 27356 10732 27384
rect 10468 27344 10474 27356
rect 1121 27319 1179 27325
rect 1121 27285 1133 27319
rect 1167 27316 1179 27319
rect 1486 27316 1492 27328
rect 1167 27288 1492 27316
rect 1167 27285 1179 27288
rect 1121 27279 1179 27285
rect 1486 27276 1492 27288
rect 1544 27276 1550 27328
rect 1581 27319 1639 27325
rect 1581 27285 1593 27319
rect 1627 27316 1639 27319
rect 2038 27316 2044 27328
rect 1627 27288 2044 27316
rect 1627 27285 1639 27288
rect 1581 27279 1639 27285
rect 2038 27276 2044 27288
rect 2096 27276 2102 27328
rect 4338 27276 4344 27328
rect 4396 27316 4402 27328
rect 5166 27316 5172 27328
rect 4396 27288 5172 27316
rect 4396 27276 4402 27288
rect 5166 27276 5172 27288
rect 5224 27276 5230 27328
rect 6178 27276 6184 27328
rect 6236 27276 6242 27328
rect 6917 27319 6975 27325
rect 6917 27285 6929 27319
rect 6963 27316 6975 27319
rect 7006 27316 7012 27328
rect 6963 27288 7012 27316
rect 6963 27285 6975 27288
rect 6917 27279 6975 27285
rect 7006 27276 7012 27288
rect 7064 27276 7070 27328
rect 7098 27276 7104 27328
rect 7156 27316 7162 27328
rect 7929 27319 7987 27325
rect 7929 27316 7941 27319
rect 7156 27288 7941 27316
rect 7156 27276 7162 27288
rect 7929 27285 7941 27288
rect 7975 27285 7987 27319
rect 7929 27279 7987 27285
rect 8570 27276 8576 27328
rect 8628 27316 8634 27328
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 8628 27288 9965 27316
rect 8628 27276 8634 27288
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 11698 27276 11704 27328
rect 11756 27276 11762 27328
rect 552 27226 12604 27248
rect 552 27174 3662 27226
rect 3714 27174 3726 27226
rect 3778 27174 3790 27226
rect 3842 27174 3854 27226
rect 3906 27174 3918 27226
rect 3970 27174 10062 27226
rect 10114 27174 10126 27226
rect 10178 27174 10190 27226
rect 10242 27174 10254 27226
rect 10306 27174 10318 27226
rect 10370 27174 12604 27226
rect 552 27152 12604 27174
rect 1762 27072 1768 27124
rect 1820 27112 1826 27124
rect 2130 27112 2136 27124
rect 1820 27084 2136 27112
rect 1820 27072 1826 27084
rect 2130 27072 2136 27084
rect 2188 27072 2194 27124
rect 4617 27115 4675 27121
rect 4617 27081 4629 27115
rect 4663 27112 4675 27115
rect 6086 27112 6092 27124
rect 4663 27084 6092 27112
rect 4663 27081 4675 27084
rect 4617 27075 4675 27081
rect 6086 27072 6092 27084
rect 6144 27072 6150 27124
rect 7282 27072 7288 27124
rect 7340 27112 7346 27124
rect 7558 27112 7564 27124
rect 7340 27084 7564 27112
rect 7340 27072 7346 27084
rect 7558 27072 7564 27084
rect 7616 27072 7622 27124
rect 7742 27072 7748 27124
rect 7800 27072 7806 27124
rect 9122 27072 9128 27124
rect 9180 27112 9186 27124
rect 9217 27115 9275 27121
rect 9217 27112 9229 27115
rect 9180 27084 9229 27112
rect 9180 27072 9186 27084
rect 9217 27081 9229 27084
rect 9263 27081 9275 27115
rect 9217 27075 9275 27081
rect 10502 27072 10508 27124
rect 10560 27112 10566 27124
rect 10781 27115 10839 27121
rect 10781 27112 10793 27115
rect 10560 27084 10793 27112
rect 10560 27072 10566 27084
rect 10781 27081 10793 27084
rect 10827 27081 10839 27115
rect 10781 27075 10839 27081
rect 11149 27115 11207 27121
rect 11149 27081 11161 27115
rect 11195 27112 11207 27115
rect 12066 27112 12072 27124
rect 11195 27084 12072 27112
rect 11195 27081 11207 27084
rect 11149 27075 11207 27081
rect 12066 27072 12072 27084
rect 12124 27072 12130 27124
rect 658 27004 664 27056
rect 716 27044 722 27056
rect 1670 27044 1676 27056
rect 716 27016 1676 27044
rect 716 27004 722 27016
rect 1670 27004 1676 27016
rect 1728 27004 1734 27056
rect 4525 27047 4583 27053
rect 4525 27013 4537 27047
rect 4571 27044 4583 27047
rect 4706 27044 4712 27056
rect 4571 27016 4712 27044
rect 4571 27013 4583 27016
rect 4525 27007 4583 27013
rect 4706 27004 4712 27016
rect 4764 27004 4770 27056
rect 4982 27004 4988 27056
rect 5040 27004 5046 27056
rect 6178 27004 6184 27056
rect 6236 27044 6242 27056
rect 6236 27016 6776 27044
rect 6236 27004 6242 27016
rect 1854 26976 1860 26988
rect 1412 26948 1860 26976
rect 1305 26911 1363 26917
rect 1305 26877 1317 26911
rect 1351 26908 1363 26911
rect 1412 26908 1440 26948
rect 1854 26936 1860 26948
rect 1912 26936 1918 26988
rect 4154 26936 4160 26988
rect 4212 26976 4218 26988
rect 5000 26976 5028 27004
rect 4212 26948 5120 26976
rect 4212 26936 4218 26948
rect 1351 26880 1440 26908
rect 1351 26877 1363 26880
rect 1305 26871 1363 26877
rect 1486 26868 1492 26920
rect 1544 26868 1550 26920
rect 1581 26911 1639 26917
rect 1581 26877 1593 26911
rect 1627 26877 1639 26911
rect 1581 26871 1639 26877
rect 474 26800 480 26852
rect 532 26840 538 26852
rect 845 26843 903 26849
rect 845 26840 857 26843
rect 532 26812 857 26840
rect 532 26800 538 26812
rect 845 26809 857 26812
rect 891 26809 903 26843
rect 845 26803 903 26809
rect 1302 26732 1308 26784
rect 1360 26772 1366 26784
rect 1596 26772 1624 26871
rect 4798 26868 4804 26920
rect 4856 26908 4862 26920
rect 5092 26917 5120 26948
rect 5626 26936 5632 26988
rect 5684 26976 5690 26988
rect 6089 26979 6147 26985
rect 6089 26976 6101 26979
rect 5684 26948 6101 26976
rect 5684 26936 5690 26948
rect 6089 26945 6101 26948
rect 6135 26945 6147 26979
rect 6089 26939 6147 26945
rect 6273 26979 6331 26985
rect 6273 26945 6285 26979
rect 6319 26976 6331 26979
rect 6362 26976 6368 26988
rect 6319 26948 6368 26976
rect 6319 26945 6331 26948
rect 6273 26939 6331 26945
rect 6362 26936 6368 26948
rect 6420 26936 6426 26988
rect 4923 26911 4981 26917
rect 4923 26908 4935 26911
rect 4856 26880 4935 26908
rect 4856 26868 4862 26880
rect 4923 26877 4935 26880
rect 4969 26877 4981 26911
rect 4923 26871 4981 26877
rect 5077 26911 5135 26917
rect 5077 26877 5089 26911
rect 5123 26877 5135 26911
rect 5077 26871 5135 26877
rect 5994 26868 6000 26920
rect 6052 26868 6058 26920
rect 6178 26868 6184 26920
rect 6236 26868 6242 26920
rect 6748 26917 6776 27016
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 7190 27044 7196 27056
rect 6880 27016 7196 27044
rect 6880 27004 6886 27016
rect 7190 27004 7196 27016
rect 7248 27004 7254 27056
rect 8573 27047 8631 27053
rect 8573 27013 8585 27047
rect 8619 27044 8631 27047
rect 8849 27047 8907 27053
rect 8849 27044 8861 27047
rect 8619 27016 8861 27044
rect 8619 27013 8631 27016
rect 8573 27007 8631 27013
rect 8849 27013 8861 27016
rect 8895 27013 8907 27047
rect 8849 27007 8907 27013
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 11425 27047 11483 27053
rect 11425 27044 11437 27047
rect 8996 27016 11437 27044
rect 8996 27004 9002 27016
rect 11425 27013 11437 27016
rect 11471 27013 11483 27047
rect 11425 27007 11483 27013
rect 7006 26936 7012 26988
rect 7064 26976 7070 26988
rect 7064 26948 7696 26976
rect 7064 26936 7070 26948
rect 6733 26911 6791 26917
rect 6733 26877 6745 26911
rect 6779 26908 6791 26911
rect 6822 26908 6828 26920
rect 6779 26880 6828 26908
rect 6779 26877 6791 26880
rect 6733 26871 6791 26877
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 7098 26868 7104 26920
rect 7156 26868 7162 26920
rect 7285 26911 7343 26917
rect 7285 26877 7297 26911
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 7300 26840 7328 26871
rect 7374 26868 7380 26920
rect 7432 26868 7438 26920
rect 7466 26868 7472 26920
rect 7524 26868 7530 26920
rect 7668 26917 7696 26948
rect 7742 26936 7748 26988
rect 7800 26976 7806 26988
rect 7800 26948 9720 26976
rect 7800 26936 7806 26948
rect 7653 26911 7711 26917
rect 7653 26877 7665 26911
rect 7699 26877 7711 26911
rect 7653 26871 7711 26877
rect 7929 26911 7987 26917
rect 7929 26877 7941 26911
rect 7975 26908 7987 26911
rect 8018 26908 8024 26920
rect 7975 26880 8024 26908
rect 7975 26877 7987 26880
rect 7929 26871 7987 26877
rect 8018 26868 8024 26880
rect 8076 26868 8082 26920
rect 8205 26911 8263 26917
rect 8205 26877 8217 26911
rect 8251 26877 8263 26911
rect 8205 26871 8263 26877
rect 7558 26840 7564 26852
rect 6564 26812 7052 26840
rect 7300 26812 7564 26840
rect 1360 26744 1624 26772
rect 4709 26775 4767 26781
rect 1360 26732 1366 26744
rect 4709 26741 4721 26775
rect 4755 26772 4767 26775
rect 4798 26772 4804 26784
rect 4755 26744 4804 26772
rect 4755 26741 4767 26744
rect 4709 26735 4767 26741
rect 4798 26732 4804 26744
rect 4856 26732 4862 26784
rect 5350 26732 5356 26784
rect 5408 26772 5414 26784
rect 5813 26775 5871 26781
rect 5813 26772 5825 26775
rect 5408 26744 5825 26772
rect 5408 26732 5414 26744
rect 5813 26741 5825 26744
rect 5859 26741 5871 26775
rect 5813 26735 5871 26741
rect 6362 26732 6368 26784
rect 6420 26772 6426 26784
rect 6564 26781 6592 26812
rect 6549 26775 6607 26781
rect 6549 26772 6561 26775
rect 6420 26744 6561 26772
rect 6420 26732 6426 26744
rect 6549 26741 6561 26744
rect 6595 26741 6607 26775
rect 6549 26735 6607 26741
rect 6638 26732 6644 26784
rect 6696 26772 6702 26784
rect 6917 26775 6975 26781
rect 6917 26772 6929 26775
rect 6696 26744 6929 26772
rect 6696 26732 6702 26744
rect 6917 26741 6929 26744
rect 6963 26741 6975 26775
rect 7024 26772 7052 26812
rect 7558 26800 7564 26812
rect 7616 26800 7622 26852
rect 8220 26840 8248 26871
rect 8386 26868 8392 26920
rect 8444 26868 8450 26920
rect 8573 26911 8631 26917
rect 8573 26877 8585 26911
rect 8619 26908 8631 26911
rect 8662 26908 8668 26920
rect 8619 26880 8668 26908
rect 8619 26877 8631 26880
rect 8573 26871 8631 26877
rect 8662 26868 8668 26880
rect 8720 26868 8726 26920
rect 8757 26911 8815 26917
rect 8757 26877 8769 26911
rect 8803 26908 8815 26911
rect 8846 26908 8852 26920
rect 8803 26880 8852 26908
rect 8803 26877 8815 26880
rect 8757 26871 8815 26877
rect 8846 26868 8852 26880
rect 8904 26868 8910 26920
rect 8938 26868 8944 26920
rect 8996 26868 9002 26920
rect 9033 26911 9091 26917
rect 9033 26877 9045 26911
rect 9079 26908 9091 26911
rect 9214 26908 9220 26920
rect 9079 26880 9220 26908
rect 9079 26877 9091 26880
rect 9033 26871 9091 26877
rect 9214 26868 9220 26880
rect 9272 26868 9278 26920
rect 9692 26917 9720 26948
rect 9766 26936 9772 26988
rect 9824 26936 9830 26988
rect 11606 26976 11612 26988
rect 9876 26948 10456 26976
rect 9677 26911 9735 26917
rect 9677 26877 9689 26911
rect 9723 26908 9735 26911
rect 9876 26908 9904 26948
rect 9723 26880 9904 26908
rect 9953 26911 10011 26917
rect 9723 26877 9735 26880
rect 9677 26871 9735 26877
rect 9953 26877 9965 26911
rect 9999 26877 10011 26911
rect 9953 26871 10011 26877
rect 8478 26840 8484 26852
rect 8220 26812 8484 26840
rect 8478 26800 8484 26812
rect 8536 26800 8542 26852
rect 9232 26840 9260 26868
rect 9232 26812 9536 26840
rect 7926 26772 7932 26784
rect 7024 26744 7932 26772
rect 6917 26735 6975 26741
rect 7926 26732 7932 26744
rect 7984 26772 7990 26784
rect 8113 26775 8171 26781
rect 8113 26772 8125 26775
rect 7984 26744 8125 26772
rect 7984 26732 7990 26744
rect 8113 26741 8125 26744
rect 8159 26741 8171 26775
rect 8113 26735 8171 26741
rect 9309 26775 9367 26781
rect 9309 26741 9321 26775
rect 9355 26772 9367 26775
rect 9398 26772 9404 26784
rect 9355 26744 9404 26772
rect 9355 26741 9367 26744
rect 9309 26735 9367 26741
rect 9398 26732 9404 26744
rect 9456 26732 9462 26784
rect 9508 26772 9536 26812
rect 9766 26800 9772 26852
rect 9824 26840 9830 26852
rect 9968 26840 9996 26871
rect 10428 26849 10456 26948
rect 10612 26948 11612 26976
rect 10612 26917 10640 26948
rect 11606 26936 11612 26948
rect 11664 26936 11670 26988
rect 11698 26936 11704 26988
rect 11756 26936 11762 26988
rect 10597 26911 10655 26917
rect 10597 26877 10609 26911
rect 10643 26877 10655 26911
rect 10597 26871 10655 26877
rect 11054 26868 11060 26920
rect 11112 26868 11118 26920
rect 11146 26868 11152 26920
rect 11204 26908 11210 26920
rect 11241 26911 11299 26917
rect 11241 26908 11253 26911
rect 11204 26880 11253 26908
rect 11204 26868 11210 26880
rect 11241 26877 11253 26880
rect 11287 26877 11299 26911
rect 11241 26871 11299 26877
rect 9824 26812 9996 26840
rect 10413 26843 10471 26849
rect 9824 26800 9830 26812
rect 10413 26809 10425 26843
rect 10459 26840 10471 26843
rect 10502 26840 10508 26852
rect 10459 26812 10508 26840
rect 10459 26809 10471 26812
rect 10413 26803 10471 26809
rect 10502 26800 10508 26812
rect 10560 26800 10566 26852
rect 10137 26775 10195 26781
rect 10137 26772 10149 26775
rect 9508 26744 10149 26772
rect 10137 26741 10149 26744
rect 10183 26741 10195 26775
rect 11072 26772 11100 26868
rect 11256 26840 11284 26871
rect 11790 26868 11796 26920
rect 11848 26868 11854 26920
rect 12342 26840 12348 26852
rect 11256 26812 12348 26840
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 11330 26772 11336 26784
rect 11072 26744 11336 26772
rect 10137 26735 10195 26741
rect 11330 26732 11336 26744
rect 11388 26732 11394 26784
rect 552 26682 12604 26704
rect 552 26630 4322 26682
rect 4374 26630 4386 26682
rect 4438 26630 4450 26682
rect 4502 26630 4514 26682
rect 4566 26630 4578 26682
rect 4630 26630 10722 26682
rect 10774 26630 10786 26682
rect 10838 26630 10850 26682
rect 10902 26630 10914 26682
rect 10966 26630 10978 26682
rect 11030 26630 12604 26682
rect 552 26608 12604 26630
rect 1302 26528 1308 26580
rect 1360 26568 1366 26580
rect 2507 26571 2565 26577
rect 2507 26568 2519 26571
rect 1360 26540 1992 26568
rect 1360 26528 1366 26540
rect 1394 26500 1400 26512
rect 860 26472 1400 26500
rect 860 26441 888 26472
rect 1394 26460 1400 26472
rect 1452 26460 1458 26512
rect 845 26435 903 26441
rect 845 26401 857 26435
rect 891 26401 903 26435
rect 845 26395 903 26401
rect 1112 26435 1170 26441
rect 1112 26401 1124 26435
rect 1158 26432 1170 26435
rect 1486 26432 1492 26444
rect 1158 26404 1492 26432
rect 1158 26401 1170 26404
rect 1112 26395 1170 26401
rect 1486 26392 1492 26404
rect 1544 26392 1550 26444
rect 1964 26296 1992 26540
rect 2240 26540 2519 26568
rect 2130 26324 2136 26376
rect 2188 26364 2194 26376
rect 2240 26364 2268 26540
rect 2507 26537 2519 26540
rect 2553 26537 2565 26571
rect 5810 26568 5816 26580
rect 2507 26531 2565 26537
rect 2884 26540 5816 26568
rect 2314 26460 2320 26512
rect 2372 26500 2378 26512
rect 2777 26503 2835 26509
rect 2777 26500 2789 26503
rect 2372 26472 2789 26500
rect 2372 26460 2378 26472
rect 2777 26469 2789 26472
rect 2823 26469 2835 26503
rect 2777 26463 2835 26469
rect 2409 26435 2467 26441
rect 2409 26401 2421 26435
rect 2455 26432 2467 26435
rect 2498 26432 2504 26444
rect 2455 26404 2504 26432
rect 2455 26401 2467 26404
rect 2409 26395 2467 26401
rect 2498 26392 2504 26404
rect 2556 26392 2562 26444
rect 2590 26392 2596 26444
rect 2648 26392 2654 26444
rect 2685 26435 2743 26441
rect 2685 26401 2697 26435
rect 2731 26432 2743 26435
rect 2884 26432 2912 26540
rect 5810 26528 5816 26540
rect 5868 26528 5874 26580
rect 5997 26571 6055 26577
rect 5997 26537 6009 26571
rect 6043 26568 6055 26571
rect 6178 26568 6184 26580
rect 6043 26540 6184 26568
rect 6043 26537 6055 26540
rect 5997 26531 6055 26537
rect 6178 26528 6184 26540
rect 6236 26528 6242 26580
rect 7193 26571 7251 26577
rect 7193 26537 7205 26571
rect 7239 26568 7251 26571
rect 7374 26568 7380 26580
rect 7239 26540 7380 26568
rect 7239 26537 7251 26540
rect 7193 26531 7251 26537
rect 7374 26528 7380 26540
rect 7432 26528 7438 26580
rect 8938 26528 8944 26580
rect 8996 26528 9002 26580
rect 9214 26528 9220 26580
rect 9272 26568 9278 26580
rect 9272 26540 9352 26568
rect 9272 26528 9278 26540
rect 2958 26460 2964 26512
rect 3016 26460 3022 26512
rect 4154 26460 4160 26512
rect 4212 26500 4218 26512
rect 4341 26503 4399 26509
rect 4341 26500 4353 26503
rect 4212 26472 4353 26500
rect 4212 26460 4218 26472
rect 4341 26469 4353 26472
rect 4387 26469 4399 26503
rect 6638 26500 6644 26512
rect 4341 26463 4399 26469
rect 5000 26472 6644 26500
rect 2731 26404 2912 26432
rect 3053 26435 3111 26441
rect 2731 26401 2743 26404
rect 2685 26395 2743 26401
rect 3053 26401 3065 26435
rect 3099 26401 3111 26435
rect 3053 26395 3111 26401
rect 3973 26435 4031 26441
rect 3973 26401 3985 26435
rect 4019 26432 4031 26435
rect 4706 26432 4712 26444
rect 4019 26404 4712 26432
rect 4019 26401 4031 26404
rect 3973 26395 4031 26401
rect 3068 26364 3096 26395
rect 4706 26392 4712 26404
rect 4764 26392 4770 26444
rect 5000 26441 5028 26472
rect 6638 26460 6644 26472
rect 6696 26460 6702 26512
rect 9324 26500 9352 26540
rect 10502 26528 10508 26580
rect 10560 26568 10566 26580
rect 11882 26568 11888 26580
rect 10560 26540 11888 26568
rect 10560 26528 10566 26540
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 9324 26472 9628 26500
rect 4801 26435 4859 26441
rect 4801 26401 4813 26435
rect 4847 26401 4859 26435
rect 4801 26395 4859 26401
rect 4985 26435 5043 26441
rect 4985 26401 4997 26435
rect 5031 26401 5043 26435
rect 4985 26395 5043 26401
rect 2188 26336 2268 26364
rect 2424 26336 3096 26364
rect 2188 26324 2194 26336
rect 2225 26299 2283 26305
rect 2225 26296 2237 26299
rect 1964 26268 2237 26296
rect 2225 26265 2237 26268
rect 2271 26265 2283 26299
rect 2225 26259 2283 26265
rect 2424 26240 2452 26336
rect 2774 26256 2780 26308
rect 2832 26256 2838 26308
rect 3234 26256 3240 26308
rect 3292 26296 3298 26308
rect 3510 26296 3516 26308
rect 3292 26268 3516 26296
rect 3292 26256 3298 26268
rect 3510 26256 3516 26268
rect 3568 26256 3574 26308
rect 4816 26296 4844 26395
rect 5350 26392 5356 26444
rect 5408 26392 5414 26444
rect 6273 26435 6331 26441
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 6362 26432 6368 26444
rect 6319 26404 6368 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 4893 26367 4951 26373
rect 4893 26333 4905 26367
rect 4939 26364 4951 26367
rect 5261 26367 5319 26373
rect 5261 26364 5273 26367
rect 4939 26336 5273 26364
rect 4939 26333 4951 26336
rect 4893 26327 4951 26333
rect 5261 26333 5273 26336
rect 5307 26333 5319 26367
rect 5261 26327 5319 26333
rect 5442 26324 5448 26376
rect 5500 26324 5506 26376
rect 5534 26324 5540 26376
rect 5592 26324 5598 26376
rect 6288 26296 6316 26395
rect 6362 26392 6368 26404
rect 6420 26392 6426 26444
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 6825 26435 6883 26441
rect 6825 26432 6837 26435
rect 6595 26404 6837 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 6825 26401 6837 26404
rect 6871 26432 6883 26435
rect 7469 26435 7527 26441
rect 6871 26404 7431 26432
rect 6871 26401 6883 26404
rect 6825 26395 6883 26401
rect 6733 26367 6791 26373
rect 6733 26333 6745 26367
rect 6779 26364 6791 26367
rect 7098 26364 7104 26376
rect 6779 26336 7104 26364
rect 6779 26333 6791 26336
rect 6733 26327 6791 26333
rect 7098 26324 7104 26336
rect 7156 26324 7162 26376
rect 7282 26324 7288 26376
rect 7340 26324 7346 26376
rect 4816 26268 6316 26296
rect 6362 26256 6368 26308
rect 6420 26296 6426 26308
rect 7300 26296 7328 26324
rect 6420 26268 7328 26296
rect 6420 26256 6426 26268
rect 1486 26188 1492 26240
rect 1544 26228 1550 26240
rect 1854 26228 1860 26240
rect 1544 26200 1860 26228
rect 1544 26188 1550 26200
rect 1854 26188 1860 26200
rect 1912 26188 1918 26240
rect 2406 26188 2412 26240
rect 2464 26188 2470 26240
rect 4246 26188 4252 26240
rect 4304 26228 4310 26240
rect 4341 26231 4399 26237
rect 4341 26228 4353 26231
rect 4304 26200 4353 26228
rect 4304 26188 4310 26200
rect 4341 26197 4353 26200
rect 4387 26197 4399 26231
rect 4341 26191 4399 26197
rect 4522 26188 4528 26240
rect 4580 26188 4586 26240
rect 5074 26188 5080 26240
rect 5132 26188 5138 26240
rect 6457 26231 6515 26237
rect 6457 26197 6469 26231
rect 6503 26228 6515 26231
rect 6638 26228 6644 26240
rect 6503 26200 6644 26228
rect 6503 26197 6515 26200
rect 6457 26191 6515 26197
rect 6638 26188 6644 26200
rect 6696 26188 6702 26240
rect 6822 26188 6828 26240
rect 6880 26228 6886 26240
rect 7006 26228 7012 26240
rect 6880 26200 7012 26228
rect 6880 26188 6886 26200
rect 7006 26188 7012 26200
rect 7064 26188 7070 26240
rect 7282 26188 7288 26240
rect 7340 26188 7346 26240
rect 7403 26228 7431 26404
rect 7469 26401 7481 26435
rect 7515 26401 7527 26435
rect 7469 26395 7527 26401
rect 7561 26435 7619 26441
rect 7561 26401 7573 26435
rect 7607 26401 7619 26435
rect 7561 26395 7619 26401
rect 7653 26435 7711 26441
rect 7653 26401 7665 26435
rect 7699 26432 7711 26435
rect 7742 26432 7748 26444
rect 7699 26404 7748 26432
rect 7699 26401 7711 26404
rect 7653 26395 7711 26401
rect 7484 26296 7512 26395
rect 7576 26364 7604 26395
rect 7742 26392 7748 26404
rect 7800 26392 7806 26444
rect 7837 26435 7895 26441
rect 7837 26401 7849 26435
rect 7883 26401 7895 26435
rect 7837 26395 7895 26401
rect 7852 26364 7880 26395
rect 7926 26392 7932 26444
rect 7984 26392 7990 26444
rect 8202 26392 8208 26444
rect 8260 26392 8266 26444
rect 8389 26435 8447 26441
rect 8389 26401 8401 26435
rect 8435 26401 8447 26435
rect 8389 26395 8447 26401
rect 8481 26425 8539 26431
rect 7576 26336 7788 26364
rect 7852 26336 8248 26364
rect 7760 26308 7788 26336
rect 7650 26296 7656 26308
rect 7484 26268 7656 26296
rect 7650 26256 7656 26268
rect 7708 26256 7714 26308
rect 7742 26256 7748 26308
rect 7800 26256 7806 26308
rect 8220 26305 8248 26336
rect 8205 26299 8263 26305
rect 8205 26265 8217 26299
rect 8251 26265 8263 26299
rect 8205 26259 8263 26265
rect 8294 26228 8300 26240
rect 7403 26200 8300 26228
rect 8294 26188 8300 26200
rect 8352 26188 8358 26240
rect 8404 26228 8432 26395
rect 8481 26391 8493 26425
rect 8527 26391 8539 26425
rect 8570 26392 8576 26444
rect 8628 26392 8634 26444
rect 8754 26392 8760 26444
rect 8812 26392 8818 26444
rect 9122 26392 9128 26444
rect 9180 26432 9186 26444
rect 9324 26441 9352 26472
rect 9217 26435 9275 26441
rect 9217 26432 9229 26435
rect 9180 26404 9229 26432
rect 9180 26392 9186 26404
rect 9217 26401 9229 26404
rect 9263 26401 9275 26435
rect 9217 26395 9275 26401
rect 9309 26435 9367 26441
rect 9309 26401 9321 26435
rect 9355 26401 9367 26435
rect 9309 26395 9367 26401
rect 9398 26392 9404 26444
rect 9456 26392 9462 26444
rect 9600 26441 9628 26472
rect 9585 26435 9643 26441
rect 9585 26401 9597 26435
rect 9631 26401 9643 26435
rect 9585 26395 9643 26401
rect 8481 26385 8539 26391
rect 8496 26296 8524 26385
rect 8846 26324 8852 26376
rect 8904 26364 8910 26376
rect 9033 26367 9091 26373
rect 9033 26364 9045 26367
rect 8904 26336 9045 26364
rect 8904 26324 8910 26336
rect 9033 26333 9045 26336
rect 9079 26364 9091 26367
rect 9493 26367 9551 26373
rect 9493 26364 9505 26367
rect 9079 26336 9505 26364
rect 9079 26333 9091 26336
rect 9033 26327 9091 26333
rect 9493 26333 9505 26336
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9125 26299 9183 26305
rect 9125 26296 9137 26299
rect 8496 26268 9137 26296
rect 9125 26265 9137 26268
rect 9171 26265 9183 26299
rect 9125 26259 9183 26265
rect 8938 26228 8944 26240
rect 8404 26200 8944 26228
rect 8938 26188 8944 26200
rect 8996 26188 9002 26240
rect 552 26138 12604 26160
rect 552 26086 3662 26138
rect 3714 26086 3726 26138
rect 3778 26086 3790 26138
rect 3842 26086 3854 26138
rect 3906 26086 3918 26138
rect 3970 26086 10062 26138
rect 10114 26086 10126 26138
rect 10178 26086 10190 26138
rect 10242 26086 10254 26138
rect 10306 26086 10318 26138
rect 10370 26086 12604 26138
rect 552 26064 12604 26086
rect 2406 25984 2412 26036
rect 2464 25984 2470 26036
rect 2590 25984 2596 26036
rect 2648 25984 2654 26036
rect 4062 26024 4068 26036
rect 3068 25996 4068 26024
rect 2317 25959 2375 25965
rect 2317 25925 2329 25959
rect 2363 25956 2375 25959
rect 3068 25956 3096 25996
rect 4062 25984 4068 25996
rect 4120 25984 4126 26036
rect 4801 26027 4859 26033
rect 4801 25993 4813 26027
rect 4847 26024 4859 26027
rect 4982 26024 4988 26036
rect 4847 25996 4988 26024
rect 4847 25993 4859 25996
rect 4801 25987 4859 25993
rect 4982 25984 4988 25996
rect 5040 26024 5046 26036
rect 5626 26024 5632 26036
rect 5040 25996 5632 26024
rect 5040 25984 5046 25996
rect 5626 25984 5632 25996
rect 5684 25984 5690 26036
rect 5994 25984 6000 26036
rect 6052 26024 6058 26036
rect 6641 26027 6699 26033
rect 6641 26024 6653 26027
rect 6052 25996 6653 26024
rect 6052 25984 6058 25996
rect 6641 25993 6653 25996
rect 6687 25993 6699 26027
rect 6641 25987 6699 25993
rect 6822 25984 6828 26036
rect 6880 26024 6886 26036
rect 6880 25996 9674 26024
rect 6880 25984 6886 25996
rect 2363 25928 3096 25956
rect 2363 25925 2375 25928
rect 2317 25919 2375 25925
rect 3142 25916 3148 25968
rect 3200 25916 3206 25968
rect 7282 25956 7288 25968
rect 6104 25928 7288 25956
rect 1026 25848 1032 25900
rect 1084 25848 1090 25900
rect 1946 25888 1952 25900
rect 1688 25860 1952 25888
rect 1486 25780 1492 25832
rect 1544 25780 1550 25832
rect 1688 25829 1716 25860
rect 1946 25848 1952 25860
rect 2004 25848 2010 25900
rect 2501 25891 2559 25897
rect 2501 25857 2513 25891
rect 2547 25888 2559 25891
rect 2590 25888 2596 25900
rect 2547 25860 2596 25888
rect 2547 25857 2559 25860
rect 2501 25851 2559 25857
rect 2590 25848 2596 25860
rect 2648 25848 2654 25900
rect 3160 25888 3188 25916
rect 3513 25891 3571 25897
rect 3513 25888 3525 25891
rect 2976 25860 3188 25888
rect 3344 25860 3525 25888
rect 2976 25832 3004 25860
rect 1673 25823 1731 25829
rect 1673 25789 1685 25823
rect 1719 25789 1731 25823
rect 1673 25783 1731 25789
rect 1765 25823 1823 25829
rect 1765 25789 1777 25823
rect 1811 25789 1823 25823
rect 1765 25783 1823 25789
rect 2225 25823 2283 25829
rect 2225 25789 2237 25823
rect 2271 25789 2283 25823
rect 2225 25783 2283 25789
rect 2777 25823 2835 25829
rect 2777 25789 2789 25823
rect 2823 25820 2835 25823
rect 2866 25820 2872 25832
rect 2823 25792 2872 25820
rect 2823 25789 2835 25792
rect 2777 25783 2835 25789
rect 1780 25684 1808 25783
rect 492 25656 1808 25684
rect 2240 25684 2268 25783
rect 2866 25780 2872 25792
rect 2924 25780 2930 25832
rect 2958 25780 2964 25832
rect 3016 25780 3022 25832
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25820 3111 25823
rect 3142 25820 3148 25832
rect 3099 25792 3148 25820
rect 3099 25789 3111 25792
rect 3053 25783 3111 25789
rect 3142 25780 3148 25792
rect 3200 25780 3206 25832
rect 3344 25684 3372 25860
rect 3513 25857 3525 25860
rect 3559 25888 3571 25891
rect 5534 25888 5540 25900
rect 3559 25860 5540 25888
rect 3559 25857 3571 25860
rect 3513 25851 3571 25857
rect 5534 25848 5540 25860
rect 5592 25888 5598 25900
rect 6104 25897 6132 25928
rect 7282 25916 7288 25928
rect 7340 25916 7346 25968
rect 9646 25956 9674 25996
rect 10410 25984 10416 26036
rect 10468 26024 10474 26036
rect 10468 25996 10916 26024
rect 10468 25984 10474 25996
rect 10428 25956 10456 25984
rect 9646 25928 10456 25956
rect 10689 25959 10747 25965
rect 10689 25925 10701 25959
rect 10735 25925 10747 25959
rect 10689 25919 10747 25925
rect 5905 25891 5963 25897
rect 5905 25888 5917 25891
rect 5592 25860 5917 25888
rect 5592 25848 5598 25860
rect 5905 25857 5917 25860
rect 5951 25857 5963 25891
rect 5905 25851 5963 25857
rect 6089 25891 6147 25897
rect 6089 25857 6101 25891
rect 6135 25857 6147 25891
rect 6089 25851 6147 25857
rect 6181 25891 6239 25897
rect 6181 25857 6193 25891
rect 6227 25888 6239 25891
rect 7009 25891 7067 25897
rect 7009 25888 7021 25891
rect 6227 25860 7021 25888
rect 6227 25857 6239 25860
rect 6181 25851 6239 25857
rect 7009 25857 7021 25860
rect 7055 25857 7067 25891
rect 7009 25851 7067 25857
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 10229 25891 10287 25897
rect 10229 25888 10241 25891
rect 9916 25860 10241 25888
rect 9916 25848 9922 25860
rect 10229 25857 10241 25860
rect 10275 25888 10287 25891
rect 10704 25888 10732 25919
rect 10275 25860 10732 25888
rect 10275 25857 10287 25860
rect 10229 25851 10287 25857
rect 3418 25780 3424 25832
rect 3476 25820 3482 25832
rect 3694 25820 3700 25832
rect 3476 25792 3700 25820
rect 3476 25780 3482 25792
rect 3694 25780 3700 25792
rect 3752 25780 3758 25832
rect 3970 25780 3976 25832
rect 4028 25780 4034 25832
rect 4154 25780 4160 25832
rect 4212 25780 4218 25832
rect 4246 25780 4252 25832
rect 4304 25820 4310 25832
rect 4525 25823 4583 25829
rect 4525 25820 4537 25823
rect 4304 25792 4537 25820
rect 4304 25780 4310 25792
rect 4525 25789 4537 25792
rect 4571 25789 4583 25823
rect 4525 25783 4583 25789
rect 4617 25823 4675 25829
rect 4617 25789 4629 25823
rect 4663 25820 4675 25823
rect 4706 25820 4712 25832
rect 4663 25792 4712 25820
rect 4663 25789 4675 25792
rect 4617 25783 4675 25789
rect 4706 25780 4712 25792
rect 4764 25780 4770 25832
rect 5445 25823 5503 25829
rect 5445 25789 5457 25823
rect 5491 25789 5503 25823
rect 5997 25823 6055 25829
rect 5997 25820 6009 25823
rect 5445 25783 5503 25789
rect 5644 25792 6009 25820
rect 3510 25712 3516 25764
rect 3568 25752 3574 25764
rect 5460 25752 5488 25783
rect 5534 25752 5540 25764
rect 3568 25724 5540 25752
rect 3568 25712 3574 25724
rect 5534 25712 5540 25724
rect 5592 25712 5598 25764
rect 2240 25656 3372 25684
rect 492 25480 520 25656
rect 3418 25644 3424 25696
rect 3476 25684 3482 25696
rect 3881 25687 3939 25693
rect 3881 25684 3893 25687
rect 3476 25656 3893 25684
rect 3476 25644 3482 25656
rect 3881 25653 3893 25656
rect 3927 25653 3939 25687
rect 3881 25647 3939 25653
rect 5166 25644 5172 25696
rect 5224 25684 5230 25696
rect 5442 25684 5448 25696
rect 5224 25656 5448 25684
rect 5224 25644 5230 25656
rect 5442 25644 5448 25656
rect 5500 25684 5506 25696
rect 5644 25693 5672 25792
rect 5997 25789 6009 25792
rect 6043 25789 6055 25823
rect 5997 25783 6055 25789
rect 6638 25780 6644 25832
rect 6696 25829 6702 25832
rect 6696 25823 6729 25829
rect 6717 25789 6729 25823
rect 6696 25783 6729 25789
rect 6825 25823 6883 25829
rect 6825 25789 6837 25823
rect 6871 25789 6883 25823
rect 6825 25783 6883 25789
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25820 6975 25823
rect 6963 25792 7052 25820
rect 6963 25789 6975 25792
rect 6917 25783 6975 25789
rect 6696 25780 6702 25783
rect 5629 25687 5687 25693
rect 5629 25684 5641 25687
rect 5500 25656 5641 25684
rect 5500 25644 5506 25656
rect 5629 25653 5641 25656
rect 5675 25653 5687 25687
rect 5629 25647 5687 25653
rect 5810 25644 5816 25696
rect 5868 25684 5874 25696
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 5868 25656 6377 25684
rect 5868 25644 5874 25656
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6840 25684 6868 25783
rect 7024 25764 7052 25792
rect 7098 25780 7104 25832
rect 7156 25780 7162 25832
rect 8570 25780 8576 25832
rect 8628 25780 8634 25832
rect 8846 25780 8852 25832
rect 8904 25820 8910 25832
rect 9030 25820 9036 25832
rect 8904 25792 9036 25820
rect 8904 25780 8910 25792
rect 9030 25780 9036 25792
rect 9088 25820 9094 25832
rect 9309 25823 9367 25829
rect 9309 25820 9321 25823
rect 9088 25792 9321 25820
rect 9088 25780 9094 25792
rect 9309 25789 9321 25792
rect 9355 25789 9367 25823
rect 9309 25783 9367 25789
rect 9398 25780 9404 25832
rect 9456 25820 9462 25832
rect 9493 25823 9551 25829
rect 9493 25820 9505 25823
rect 9456 25792 9505 25820
rect 9456 25780 9462 25792
rect 9493 25789 9505 25792
rect 9539 25789 9551 25823
rect 9493 25783 9551 25789
rect 10413 25823 10471 25829
rect 10413 25789 10425 25823
rect 10459 25789 10471 25823
rect 10413 25783 10471 25789
rect 7006 25712 7012 25764
rect 7064 25712 7070 25764
rect 8757 25755 8815 25761
rect 8757 25721 8769 25755
rect 8803 25752 8815 25755
rect 9122 25752 9128 25764
rect 8803 25724 9128 25752
rect 8803 25721 8815 25724
rect 8757 25715 8815 25721
rect 9122 25712 9128 25724
rect 9180 25752 9186 25764
rect 9766 25752 9772 25764
rect 9180 25724 9772 25752
rect 9180 25712 9186 25724
rect 9766 25712 9772 25724
rect 9824 25712 9830 25764
rect 10428 25752 10456 25783
rect 10502 25780 10508 25832
rect 10560 25780 10566 25832
rect 10888 25829 10916 25996
rect 10873 25823 10931 25829
rect 10873 25789 10885 25823
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 10594 25752 10600 25764
rect 10428 25724 10600 25752
rect 10594 25712 10600 25724
rect 10652 25712 10658 25764
rect 10888 25752 10916 25783
rect 11054 25780 11060 25832
rect 11112 25820 11118 25832
rect 11149 25823 11207 25829
rect 11149 25820 11161 25823
rect 11112 25792 11161 25820
rect 11112 25780 11118 25792
rect 11149 25789 11161 25792
rect 11195 25789 11207 25823
rect 11149 25783 11207 25789
rect 11333 25823 11391 25829
rect 11333 25789 11345 25823
rect 11379 25820 11391 25823
rect 11885 25823 11943 25829
rect 11379 25792 11560 25820
rect 11379 25789 11391 25792
rect 11333 25783 11391 25789
rect 11422 25752 11428 25764
rect 10888 25724 11428 25752
rect 11422 25712 11428 25724
rect 11480 25712 11486 25764
rect 8294 25684 8300 25696
rect 6840 25656 8300 25684
rect 6365 25647 6423 25653
rect 8294 25644 8300 25656
rect 8352 25684 8358 25696
rect 8662 25684 8668 25696
rect 8352 25656 8668 25684
rect 8352 25644 8358 25656
rect 8662 25644 8668 25656
rect 8720 25644 8726 25696
rect 9401 25687 9459 25693
rect 9401 25653 9413 25687
rect 9447 25684 9459 25687
rect 9582 25684 9588 25696
rect 9447 25656 9588 25684
rect 9447 25653 9459 25656
rect 9401 25647 9459 25653
rect 9582 25644 9588 25656
rect 9640 25644 9646 25696
rect 10229 25687 10287 25693
rect 10229 25653 10241 25687
rect 10275 25684 10287 25687
rect 10410 25684 10416 25696
rect 10275 25656 10416 25684
rect 10275 25653 10287 25656
rect 10229 25647 10287 25653
rect 10410 25644 10416 25656
rect 10468 25644 10474 25696
rect 11238 25644 11244 25696
rect 11296 25644 11302 25696
rect 11532 25684 11560 25792
rect 11885 25789 11897 25823
rect 11931 25789 11943 25823
rect 11885 25783 11943 25789
rect 11977 25823 12035 25829
rect 11977 25789 11989 25823
rect 12023 25820 12035 25823
rect 12618 25820 12624 25832
rect 12023 25792 12624 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 11900 25752 11928 25783
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 12066 25752 12072 25764
rect 11900 25724 12072 25752
rect 12066 25712 12072 25724
rect 12124 25712 12130 25764
rect 11790 25684 11796 25696
rect 11532 25656 11796 25684
rect 11790 25644 11796 25656
rect 11848 25684 11854 25696
rect 11974 25684 11980 25696
rect 11848 25656 11980 25684
rect 11848 25644 11854 25656
rect 11974 25644 11980 25656
rect 12032 25644 12038 25696
rect 12158 25644 12164 25696
rect 12216 25644 12222 25696
rect 552 25594 12604 25616
rect 552 25542 4322 25594
rect 4374 25542 4386 25594
rect 4438 25542 4450 25594
rect 4502 25542 4514 25594
rect 4566 25542 4578 25594
rect 4630 25542 10722 25594
rect 10774 25542 10786 25594
rect 10838 25542 10850 25594
rect 10902 25542 10914 25594
rect 10966 25542 10978 25594
rect 11030 25542 12604 25594
rect 552 25520 12604 25542
rect 845 25483 903 25489
rect 845 25480 857 25483
rect 492 25452 857 25480
rect 845 25449 857 25452
rect 891 25449 903 25483
rect 845 25443 903 25449
rect 1670 25440 1676 25492
rect 1728 25480 1734 25492
rect 1728 25452 2360 25480
rect 1728 25440 1734 25452
rect 1394 25372 1400 25424
rect 1452 25412 1458 25424
rect 1452 25384 2268 25412
rect 1452 25372 1458 25384
rect 1946 25304 1952 25356
rect 2004 25353 2010 25356
rect 2240 25353 2268 25384
rect 2004 25344 2016 25353
rect 2225 25347 2283 25353
rect 2004 25316 2049 25344
rect 2004 25307 2016 25316
rect 2225 25313 2237 25347
rect 2271 25313 2283 25347
rect 2332 25344 2360 25452
rect 2590 25440 2596 25492
rect 2648 25480 2654 25492
rect 2869 25483 2927 25489
rect 2869 25480 2881 25483
rect 2648 25452 2881 25480
rect 2648 25440 2654 25452
rect 2869 25449 2881 25452
rect 2915 25449 2927 25483
rect 2869 25443 2927 25449
rect 3142 25440 3148 25492
rect 3200 25440 3206 25492
rect 4062 25440 4068 25492
rect 4120 25480 4126 25492
rect 6641 25483 6699 25489
rect 6641 25480 6653 25483
rect 4120 25452 6653 25480
rect 4120 25440 4126 25452
rect 6641 25449 6653 25452
rect 6687 25449 6699 25483
rect 6641 25443 6699 25449
rect 7098 25440 7104 25492
rect 7156 25480 7162 25492
rect 7377 25483 7435 25489
rect 7377 25480 7389 25483
rect 7156 25452 7389 25480
rect 7156 25440 7162 25452
rect 7377 25449 7389 25452
rect 7423 25449 7435 25483
rect 7377 25443 7435 25449
rect 7926 25440 7932 25492
rect 7984 25480 7990 25492
rect 8662 25480 8668 25492
rect 7984 25452 8668 25480
rect 7984 25440 7990 25452
rect 8662 25440 8668 25452
rect 8720 25440 8726 25492
rect 9217 25483 9275 25489
rect 9217 25449 9229 25483
rect 9263 25449 9275 25483
rect 9217 25443 9275 25449
rect 10321 25483 10379 25489
rect 10321 25449 10333 25483
rect 10367 25480 10379 25483
rect 10502 25480 10508 25492
rect 10367 25452 10508 25480
rect 10367 25449 10379 25452
rect 10321 25443 10379 25449
rect 2498 25372 2504 25424
rect 2556 25412 2562 25424
rect 2685 25415 2743 25421
rect 2685 25412 2697 25415
rect 2556 25384 2697 25412
rect 2556 25372 2562 25384
rect 2685 25381 2697 25384
rect 2731 25381 2743 25415
rect 5074 25412 5080 25424
rect 2685 25375 2743 25381
rect 2976 25384 5080 25412
rect 2976 25353 3004 25384
rect 5074 25372 5080 25384
rect 5132 25372 5138 25424
rect 5169 25415 5227 25421
rect 5169 25381 5181 25415
rect 5215 25412 5227 25415
rect 6822 25412 6828 25424
rect 5215 25384 6828 25412
rect 5215 25381 5227 25384
rect 5169 25375 5227 25381
rect 6822 25372 6828 25384
rect 6880 25372 6886 25424
rect 9232 25412 9260 25443
rect 10502 25440 10508 25452
rect 10560 25480 10566 25492
rect 10597 25483 10655 25489
rect 10597 25480 10609 25483
rect 10560 25452 10609 25480
rect 10560 25440 10566 25452
rect 10597 25449 10609 25452
rect 10643 25449 10655 25483
rect 10965 25483 11023 25489
rect 10965 25480 10977 25483
rect 10597 25443 10655 25449
rect 10704 25452 10977 25480
rect 7116 25384 9260 25412
rect 2593 25347 2651 25353
rect 2593 25344 2605 25347
rect 2332 25316 2605 25344
rect 2225 25307 2283 25313
rect 2593 25313 2605 25316
rect 2639 25313 2651 25347
rect 2593 25307 2651 25313
rect 2961 25347 3019 25353
rect 2961 25313 2973 25347
rect 3007 25313 3019 25347
rect 2961 25307 3019 25313
rect 3329 25347 3387 25353
rect 3329 25313 3341 25347
rect 3375 25344 3387 25347
rect 3418 25344 3424 25356
rect 3375 25316 3424 25344
rect 3375 25313 3387 25316
rect 3329 25307 3387 25313
rect 2004 25304 2010 25307
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25276 2375 25279
rect 2406 25276 2412 25288
rect 2363 25248 2412 25276
rect 2363 25245 2375 25248
rect 2317 25239 2375 25245
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 2608 25276 2636 25307
rect 3344 25276 3372 25307
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 3510 25304 3516 25356
rect 3568 25304 3574 25356
rect 4706 25304 4712 25356
rect 4764 25344 4770 25356
rect 4801 25347 4859 25353
rect 4801 25344 4813 25347
rect 4764 25316 4813 25344
rect 4764 25304 4770 25316
rect 4801 25313 4813 25316
rect 4847 25313 4859 25347
rect 4801 25307 4859 25313
rect 4985 25347 5043 25353
rect 4985 25313 4997 25347
rect 5031 25313 5043 25347
rect 4985 25307 5043 25313
rect 2608 25248 3372 25276
rect 5000 25276 5028 25307
rect 6362 25304 6368 25356
rect 6420 25344 6426 25356
rect 6917 25347 6975 25353
rect 6917 25344 6929 25347
rect 6420 25316 6929 25344
rect 6420 25304 6426 25316
rect 6917 25313 6929 25316
rect 6963 25313 6975 25347
rect 6917 25307 6975 25313
rect 7006 25304 7012 25356
rect 7064 25304 7070 25356
rect 7116 25353 7144 25384
rect 9582 25372 9588 25424
rect 9640 25412 9646 25424
rect 9677 25415 9735 25421
rect 9677 25412 9689 25415
rect 9640 25384 9689 25412
rect 9640 25372 9646 25384
rect 9677 25381 9689 25384
rect 9723 25381 9735 25415
rect 9677 25375 9735 25381
rect 10410 25372 10416 25424
rect 10468 25372 10474 25424
rect 7101 25347 7159 25353
rect 7101 25313 7113 25347
rect 7147 25313 7159 25347
rect 7101 25307 7159 25313
rect 7285 25347 7343 25353
rect 7285 25313 7297 25347
rect 7331 25313 7343 25347
rect 7285 25307 7343 25313
rect 7653 25347 7711 25353
rect 7653 25313 7665 25347
rect 7699 25344 7711 25347
rect 7742 25344 7748 25356
rect 7699 25316 7748 25344
rect 7699 25313 7711 25316
rect 7653 25307 7711 25313
rect 5074 25276 5080 25288
rect 5000 25248 5080 25276
rect 5074 25236 5080 25248
rect 5132 25236 5138 25288
rect 5534 25236 5540 25288
rect 5592 25276 5598 25288
rect 6822 25276 6828 25288
rect 5592 25248 6828 25276
rect 5592 25236 5598 25248
rect 6822 25236 6828 25248
rect 6880 25276 6886 25288
rect 7300 25276 7328 25307
rect 7742 25304 7748 25316
rect 7800 25304 7806 25356
rect 7929 25347 7987 25353
rect 7929 25313 7941 25347
rect 7975 25344 7987 25347
rect 8202 25344 8208 25356
rect 7975 25316 8208 25344
rect 7975 25313 7987 25316
rect 7929 25307 7987 25313
rect 8202 25304 8208 25316
rect 8260 25344 8266 25356
rect 8573 25347 8631 25353
rect 8573 25344 8585 25347
rect 8260 25316 8585 25344
rect 8260 25304 8266 25316
rect 8573 25313 8585 25316
rect 8619 25313 8631 25347
rect 8573 25307 8631 25313
rect 8662 25304 8668 25356
rect 8720 25344 8726 25356
rect 9401 25347 9459 25353
rect 9401 25344 9413 25347
rect 8720 25316 9413 25344
rect 8720 25304 8726 25316
rect 9401 25313 9413 25316
rect 9447 25313 9459 25347
rect 9401 25307 9459 25313
rect 9950 25304 9956 25356
rect 10008 25304 10014 25356
rect 10594 25304 10600 25356
rect 10652 25344 10658 25356
rect 10704 25353 10732 25452
rect 10965 25449 10977 25452
rect 11011 25449 11023 25483
rect 10965 25443 11023 25449
rect 10689 25347 10747 25353
rect 10689 25344 10701 25347
rect 10652 25316 10701 25344
rect 10652 25304 10658 25316
rect 10689 25313 10701 25316
rect 10735 25313 10747 25347
rect 10689 25307 10747 25313
rect 11333 25347 11391 25353
rect 11333 25313 11345 25347
rect 11379 25344 11391 25347
rect 11606 25344 11612 25356
rect 11379 25316 11612 25344
rect 11379 25313 11391 25316
rect 11333 25307 11391 25313
rect 11606 25304 11612 25316
rect 11664 25304 11670 25356
rect 11977 25347 12035 25353
rect 11977 25313 11989 25347
rect 12023 25344 12035 25347
rect 12066 25344 12072 25356
rect 12023 25316 12072 25344
rect 12023 25313 12035 25316
rect 11977 25307 12035 25313
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 6880 25248 7328 25276
rect 6880 25236 6886 25248
rect 7374 25236 7380 25288
rect 7432 25236 7438 25288
rect 7834 25276 7840 25288
rect 7668 25248 7840 25276
rect 2501 25211 2559 25217
rect 2501 25177 2513 25211
rect 2547 25208 2559 25211
rect 2866 25208 2872 25220
rect 2547 25180 2872 25208
rect 2547 25177 2559 25180
rect 2501 25171 2559 25177
rect 2866 25168 2872 25180
rect 2924 25208 2930 25220
rect 3050 25208 3056 25220
rect 2924 25180 3056 25208
rect 2924 25168 2930 25180
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 3142 25168 3148 25220
rect 3200 25208 3206 25220
rect 3694 25208 3700 25220
rect 3200 25180 3700 25208
rect 3200 25168 3206 25180
rect 3694 25168 3700 25180
rect 3752 25168 3758 25220
rect 4614 25168 4620 25220
rect 4672 25208 4678 25220
rect 4798 25208 4804 25220
rect 4672 25180 4804 25208
rect 4672 25168 4678 25180
rect 4798 25168 4804 25180
rect 4856 25168 4862 25220
rect 7006 25168 7012 25220
rect 7064 25208 7070 25220
rect 7668 25208 7696 25248
rect 7834 25236 7840 25248
rect 7892 25236 7898 25288
rect 8478 25236 8484 25288
rect 8536 25236 8542 25288
rect 8941 25279 8999 25285
rect 8941 25245 8953 25279
rect 8987 25276 8999 25279
rect 8987 25248 9444 25276
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 7064 25180 7696 25208
rect 8297 25211 8355 25217
rect 7064 25168 7070 25180
rect 8297 25177 8309 25211
rect 8343 25208 8355 25211
rect 9030 25208 9036 25220
rect 8343 25180 9036 25208
rect 8343 25177 8355 25180
rect 8297 25171 8355 25177
rect 9030 25168 9036 25180
rect 9088 25168 9094 25220
rect 9416 25208 9444 25248
rect 9490 25236 9496 25288
rect 9548 25236 9554 25288
rect 9766 25276 9772 25288
rect 9600 25248 9772 25276
rect 9600 25208 9628 25248
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 10045 25279 10103 25285
rect 10045 25245 10057 25279
rect 10091 25276 10103 25279
rect 10502 25276 10508 25288
rect 10091 25248 10508 25276
rect 10091 25245 10103 25248
rect 10045 25239 10103 25245
rect 10502 25236 10508 25248
rect 10560 25236 10566 25288
rect 11238 25236 11244 25288
rect 11296 25236 11302 25288
rect 11698 25236 11704 25288
rect 11756 25276 11762 25288
rect 11885 25279 11943 25285
rect 11885 25276 11897 25279
rect 11756 25248 11897 25276
rect 11756 25236 11762 25248
rect 11885 25245 11897 25248
rect 11931 25276 11943 25279
rect 12618 25276 12624 25288
rect 11931 25248 12624 25276
rect 11931 25245 11943 25248
rect 11885 25239 11943 25245
rect 12618 25236 12624 25248
rect 12676 25236 12682 25288
rect 10413 25211 10471 25217
rect 10413 25208 10425 25211
rect 9416 25180 9628 25208
rect 9692 25180 10425 25208
rect 2314 25100 2320 25152
rect 2372 25140 2378 25152
rect 2409 25143 2467 25149
rect 2409 25140 2421 25143
rect 2372 25112 2421 25140
rect 2372 25100 2378 25112
rect 2409 25109 2421 25112
rect 2455 25109 2467 25143
rect 2409 25103 2467 25109
rect 2685 25143 2743 25149
rect 2685 25109 2697 25143
rect 2731 25140 2743 25143
rect 2774 25140 2780 25152
rect 2731 25112 2780 25140
rect 2731 25109 2743 25112
rect 2685 25103 2743 25109
rect 2774 25100 2780 25112
rect 2832 25100 2838 25152
rect 6546 25100 6552 25152
rect 6604 25140 6610 25152
rect 7190 25140 7196 25152
rect 6604 25112 7196 25140
rect 6604 25100 6610 25112
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 7558 25100 7564 25152
rect 7616 25140 7622 25152
rect 8110 25140 8116 25152
rect 7616 25112 8116 25140
rect 7616 25100 7622 25112
rect 8110 25100 8116 25112
rect 8168 25100 8174 25152
rect 9692 25149 9720 25180
rect 10413 25177 10425 25180
rect 10459 25177 10471 25211
rect 10413 25171 10471 25177
rect 11514 25168 11520 25220
rect 11572 25208 11578 25220
rect 11609 25211 11667 25217
rect 11609 25208 11621 25211
rect 11572 25180 11621 25208
rect 11572 25168 11578 25180
rect 11609 25177 11621 25180
rect 11655 25177 11667 25211
rect 11609 25171 11667 25177
rect 9677 25143 9735 25149
rect 9677 25109 9689 25143
rect 9723 25109 9735 25143
rect 9677 25103 9735 25109
rect 552 25050 12604 25072
rect 552 24998 3662 25050
rect 3714 24998 3726 25050
rect 3778 24998 3790 25050
rect 3842 24998 3854 25050
rect 3906 24998 3918 25050
rect 3970 24998 10062 25050
rect 10114 24998 10126 25050
rect 10178 24998 10190 25050
rect 10242 24998 10254 25050
rect 10306 24998 10318 25050
rect 10370 24998 12604 25050
rect 552 24976 12604 24998
rect 3329 24939 3387 24945
rect 3329 24905 3341 24939
rect 3375 24936 3387 24939
rect 3694 24936 3700 24948
rect 3375 24908 3700 24936
rect 3375 24905 3387 24908
rect 3329 24899 3387 24905
rect 3694 24896 3700 24908
rect 3752 24896 3758 24948
rect 6546 24896 6552 24948
rect 6604 24896 6610 24948
rect 6638 24896 6644 24948
rect 6696 24896 6702 24948
rect 7009 24939 7067 24945
rect 7009 24905 7021 24939
rect 7055 24936 7067 24939
rect 7374 24936 7380 24948
rect 7055 24908 7380 24936
rect 7055 24905 7067 24908
rect 7009 24899 7067 24905
rect 7374 24896 7380 24908
rect 7432 24896 7438 24948
rect 7742 24896 7748 24948
rect 7800 24896 7806 24948
rect 7834 24896 7840 24948
rect 7892 24896 7898 24948
rect 7929 24939 7987 24945
rect 7929 24905 7941 24939
rect 7975 24936 7987 24939
rect 8754 24936 8760 24948
rect 7975 24908 8760 24936
rect 7975 24905 7987 24908
rect 7929 24899 7987 24905
rect 8754 24896 8760 24908
rect 8812 24896 8818 24948
rect 9401 24939 9459 24945
rect 9401 24905 9413 24939
rect 9447 24936 9459 24939
rect 9490 24936 9496 24948
rect 9447 24908 9496 24936
rect 9447 24905 9459 24908
rect 9401 24899 9459 24905
rect 9490 24896 9496 24908
rect 9548 24896 9554 24948
rect 9950 24896 9956 24948
rect 10008 24936 10014 24948
rect 10229 24939 10287 24945
rect 10229 24936 10241 24939
rect 10008 24908 10241 24936
rect 10008 24896 10014 24908
rect 10229 24905 10241 24908
rect 10275 24905 10287 24939
rect 10229 24899 10287 24905
rect 3878 24828 3884 24880
rect 3936 24868 3942 24880
rect 4706 24868 4712 24880
rect 3936 24840 4712 24868
rect 3936 24828 3942 24840
rect 4706 24828 4712 24840
rect 4764 24868 4770 24880
rect 5353 24871 5411 24877
rect 4764 24840 4936 24868
rect 4764 24828 4770 24840
rect 106 24760 112 24812
rect 164 24800 170 24812
rect 658 24800 664 24812
rect 164 24772 664 24800
rect 164 24760 170 24772
rect 658 24760 664 24772
rect 716 24760 722 24812
rect 4246 24800 4252 24812
rect 3895 24772 4252 24800
rect 1302 24692 1308 24744
rect 1360 24732 1366 24744
rect 1486 24732 1492 24744
rect 1360 24704 1492 24732
rect 1360 24692 1366 24704
rect 1486 24692 1492 24704
rect 1544 24692 1550 24744
rect 1673 24735 1731 24741
rect 1673 24701 1685 24735
rect 1719 24701 1731 24735
rect 1673 24695 1731 24701
rect 1026 24624 1032 24676
rect 1084 24624 1090 24676
rect 1118 24624 1124 24676
rect 1176 24664 1182 24676
rect 1688 24664 1716 24695
rect 1762 24692 1768 24744
rect 1820 24692 1826 24744
rect 2130 24692 2136 24744
rect 2188 24692 2194 24744
rect 2314 24692 2320 24744
rect 2372 24732 2378 24744
rect 2409 24735 2467 24741
rect 2409 24732 2421 24735
rect 2372 24704 2421 24732
rect 2372 24692 2378 24704
rect 2409 24701 2421 24704
rect 2455 24701 2467 24735
rect 2409 24695 2467 24701
rect 2593 24735 2651 24741
rect 2593 24701 2605 24735
rect 2639 24732 2651 24735
rect 2774 24732 2780 24744
rect 2639 24704 2780 24732
rect 2639 24701 2651 24704
rect 2593 24695 2651 24701
rect 2774 24692 2780 24704
rect 2832 24692 2838 24744
rect 3513 24735 3571 24741
rect 3513 24701 3525 24735
rect 3559 24701 3571 24735
rect 3513 24695 3571 24701
rect 1176 24636 1716 24664
rect 1176 24624 1182 24636
rect 1854 24624 1860 24676
rect 1912 24664 1918 24676
rect 2501 24667 2559 24673
rect 2501 24664 2513 24667
rect 1912 24636 2513 24664
rect 1912 24624 1918 24636
rect 2501 24633 2513 24636
rect 2547 24633 2559 24667
rect 3528 24664 3556 24695
rect 3602 24692 3608 24744
rect 3660 24732 3666 24744
rect 3895 24741 3923 24772
rect 4246 24760 4252 24772
rect 4304 24800 4310 24812
rect 4304 24772 4844 24800
rect 4304 24760 4310 24772
rect 3880 24735 3938 24741
rect 3880 24732 3892 24735
rect 3660 24704 3892 24732
rect 3660 24692 3666 24704
rect 3880 24701 3892 24704
rect 3926 24701 3938 24735
rect 3880 24695 3938 24701
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 4154 24732 4160 24744
rect 4019 24704 4160 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 4154 24692 4160 24704
rect 4212 24732 4218 24744
rect 4816 24741 4844 24772
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 4212 24704 4445 24732
rect 4212 24692 4218 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 4801 24735 4859 24741
rect 4801 24701 4813 24735
rect 4847 24701 4859 24735
rect 4908 24732 4936 24840
rect 5353 24837 5365 24871
rect 5399 24868 5411 24871
rect 5718 24868 5724 24880
rect 5399 24840 5724 24868
rect 5399 24837 5411 24840
rect 5353 24831 5411 24837
rect 5718 24828 5724 24840
rect 5776 24828 5782 24880
rect 6564 24800 6592 24896
rect 6196 24772 6592 24800
rect 5258 24732 5264 24744
rect 4908 24704 5264 24732
rect 4801 24695 4859 24701
rect 5258 24692 5264 24704
rect 5316 24732 5322 24744
rect 5537 24735 5595 24741
rect 5537 24732 5549 24735
rect 5316 24704 5549 24732
rect 5316 24692 5322 24704
rect 5537 24701 5549 24704
rect 5583 24732 5595 24735
rect 5721 24735 5779 24741
rect 5721 24732 5733 24735
rect 5583 24704 5733 24732
rect 5583 24701 5595 24704
rect 5537 24695 5595 24701
rect 5721 24701 5733 24704
rect 5767 24701 5779 24735
rect 5721 24695 5779 24701
rect 5810 24692 5816 24744
rect 5868 24732 5874 24744
rect 6196 24741 6224 24772
rect 5905 24735 5963 24741
rect 5905 24732 5917 24735
rect 5868 24704 5917 24732
rect 5868 24692 5874 24704
rect 5905 24701 5917 24704
rect 5951 24701 5963 24735
rect 5905 24695 5963 24701
rect 6181 24735 6239 24741
rect 6181 24701 6193 24735
rect 6227 24701 6239 24735
rect 6181 24695 6239 24701
rect 6454 24692 6460 24744
rect 6512 24692 6518 24744
rect 6656 24732 6684 24896
rect 7760 24868 7788 24896
rect 7392 24840 9674 24868
rect 7006 24800 7012 24812
rect 6932 24772 7012 24800
rect 6733 24735 6791 24741
rect 6733 24732 6745 24735
rect 6656 24704 6745 24732
rect 6733 24701 6745 24704
rect 6779 24701 6791 24735
rect 6733 24695 6791 24701
rect 6825 24735 6883 24741
rect 6825 24701 6837 24735
rect 6871 24732 6883 24735
rect 6932 24732 6960 24772
rect 7006 24760 7012 24772
rect 7064 24800 7070 24812
rect 7392 24809 7420 24840
rect 7377 24803 7435 24809
rect 7064 24772 7328 24800
rect 7064 24760 7070 24772
rect 7300 24741 7328 24772
rect 7377 24769 7389 24803
rect 7423 24769 7435 24803
rect 7377 24763 7435 24769
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 7834 24800 7840 24812
rect 7576 24772 7840 24800
rect 6871 24704 6960 24732
rect 7101 24735 7159 24741
rect 6871 24701 6883 24704
rect 6825 24695 6883 24701
rect 7101 24701 7113 24735
rect 7147 24701 7159 24735
rect 7101 24695 7159 24701
rect 7285 24735 7343 24741
rect 7285 24701 7297 24735
rect 7331 24732 7343 24735
rect 7576 24732 7604 24772
rect 7834 24760 7840 24772
rect 7892 24760 7898 24812
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8220 24772 8493 24800
rect 7331 24704 7604 24732
rect 7331 24701 7343 24704
rect 7285 24695 7343 24701
rect 4706 24664 4712 24676
rect 3528 24636 4712 24664
rect 2501 24627 2559 24633
rect 4706 24624 4712 24636
rect 4764 24624 4770 24676
rect 5074 24624 5080 24676
rect 5132 24664 5138 24676
rect 5828 24664 5856 24692
rect 5132 24636 5856 24664
rect 5997 24667 6055 24673
rect 5132 24624 5138 24636
rect 5997 24633 6009 24667
rect 6043 24664 6055 24667
rect 6086 24664 6092 24676
rect 6043 24636 6092 24664
rect 6043 24633 6055 24636
rect 5997 24627 6055 24633
rect 6086 24624 6092 24636
rect 6144 24624 6150 24676
rect 6365 24667 6423 24673
rect 6365 24633 6377 24667
rect 6411 24664 6423 24667
rect 7120 24664 7148 24695
rect 7650 24692 7656 24744
rect 7708 24692 7714 24744
rect 7742 24692 7748 24744
rect 7800 24732 7806 24744
rect 8220 24741 8248 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 8481 24763 8539 24769
rect 9214 24760 9220 24812
rect 9272 24760 9278 24812
rect 9398 24760 9404 24812
rect 9456 24800 9462 24812
rect 9493 24803 9551 24809
rect 9493 24800 9505 24803
rect 9456 24772 9505 24800
rect 9456 24760 9462 24772
rect 9493 24769 9505 24772
rect 9539 24769 9551 24803
rect 9646 24800 9674 24840
rect 9858 24828 9864 24880
rect 9916 24868 9922 24880
rect 10042 24868 10048 24880
rect 9916 24840 10048 24868
rect 9916 24828 9922 24840
rect 10042 24828 10048 24840
rect 10100 24828 10106 24880
rect 11698 24868 11704 24880
rect 11348 24840 11704 24868
rect 10318 24800 10324 24812
rect 9646 24772 10324 24800
rect 9493 24763 9551 24769
rect 10318 24760 10324 24772
rect 10376 24760 10382 24812
rect 10686 24760 10692 24812
rect 10744 24760 10750 24812
rect 11149 24803 11207 24809
rect 11149 24769 11161 24803
rect 11195 24800 11207 24803
rect 11348 24800 11376 24840
rect 11698 24828 11704 24840
rect 11756 24828 11762 24880
rect 11195 24772 11376 24800
rect 11425 24803 11483 24809
rect 11195 24769 11207 24772
rect 11149 24763 11207 24769
rect 11425 24769 11437 24803
rect 11471 24800 11483 24803
rect 11606 24800 11612 24812
rect 11471 24772 11612 24800
rect 11471 24769 11483 24772
rect 11425 24763 11483 24769
rect 11606 24760 11612 24772
rect 11664 24760 11670 24812
rect 12158 24760 12164 24812
rect 12216 24760 12222 24812
rect 8205 24735 8263 24741
rect 7800 24704 8156 24732
rect 7800 24692 7806 24704
rect 6411 24636 7148 24664
rect 6411 24633 6423 24636
rect 6365 24627 6423 24633
rect 7558 24624 7564 24676
rect 7616 24664 7622 24676
rect 7929 24667 7987 24673
rect 7929 24664 7941 24667
rect 7616 24636 7941 24664
rect 7616 24624 7622 24636
rect 7929 24633 7941 24636
rect 7975 24633 7987 24667
rect 8128 24664 8156 24704
rect 8205 24701 8217 24735
rect 8251 24701 8263 24735
rect 8205 24695 8263 24701
rect 8389 24735 8447 24741
rect 8389 24701 8401 24735
rect 8435 24701 8447 24735
rect 8389 24695 8447 24701
rect 8404 24664 8432 24695
rect 8570 24692 8576 24744
rect 8628 24732 8634 24744
rect 8757 24735 8815 24741
rect 8757 24732 8769 24735
rect 8628 24704 8769 24732
rect 8628 24692 8634 24704
rect 8757 24701 8769 24704
rect 8803 24701 8815 24735
rect 8757 24695 8815 24701
rect 8941 24735 8999 24741
rect 8941 24701 8953 24735
rect 8987 24701 8999 24735
rect 8941 24695 8999 24701
rect 8128 24636 8432 24664
rect 8956 24664 8984 24695
rect 9030 24692 9036 24744
rect 9088 24692 9094 24744
rect 9122 24692 9128 24744
rect 9180 24692 9186 24744
rect 9232 24732 9260 24760
rect 9582 24732 9588 24744
rect 9232 24704 9588 24732
rect 9582 24692 9588 24704
rect 9640 24732 9646 24744
rect 9769 24735 9827 24741
rect 9769 24732 9781 24735
rect 9640 24704 9781 24732
rect 9640 24692 9646 24704
rect 9769 24701 9781 24704
rect 9815 24701 9827 24735
rect 9769 24695 9827 24701
rect 9858 24692 9864 24744
rect 9916 24692 9922 24744
rect 9953 24735 10011 24741
rect 9953 24701 9965 24735
rect 9999 24701 10011 24735
rect 10137 24735 10195 24741
rect 10137 24732 10149 24735
rect 9953 24695 10011 24701
rect 10060 24704 10149 24732
rect 9214 24664 9220 24676
rect 8956 24636 9220 24664
rect 7929 24627 7987 24633
rect 9214 24624 9220 24636
rect 9272 24664 9278 24676
rect 9968 24664 9996 24695
rect 9272 24636 9996 24664
rect 9272 24624 9278 24636
rect 1486 24556 1492 24608
rect 1544 24596 1550 24608
rect 2225 24599 2283 24605
rect 2225 24596 2237 24599
rect 1544 24568 2237 24596
rect 1544 24556 1550 24568
rect 2225 24565 2237 24568
rect 2271 24565 2283 24599
rect 2225 24559 2283 24565
rect 3605 24599 3663 24605
rect 3605 24565 3617 24599
rect 3651 24596 3663 24599
rect 3786 24596 3792 24608
rect 3651 24568 3792 24596
rect 3651 24565 3663 24568
rect 3605 24559 3663 24565
rect 3786 24556 3792 24568
rect 3844 24556 3850 24608
rect 5813 24599 5871 24605
rect 5813 24565 5825 24599
rect 5859 24596 5871 24599
rect 8018 24596 8024 24608
rect 5859 24568 8024 24596
rect 5859 24565 5871 24568
rect 5813 24559 5871 24565
rect 8018 24556 8024 24568
rect 8076 24556 8082 24608
rect 8113 24599 8171 24605
rect 8113 24565 8125 24599
rect 8159 24596 8171 24599
rect 8202 24596 8208 24608
rect 8159 24568 8208 24596
rect 8159 24565 8171 24568
rect 8113 24559 8171 24565
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 8938 24556 8944 24608
rect 8996 24596 9002 24608
rect 9858 24596 9864 24608
rect 8996 24568 9864 24596
rect 8996 24556 9002 24568
rect 9858 24556 9864 24568
rect 9916 24596 9922 24608
rect 10060 24596 10088 24704
rect 10137 24701 10149 24704
rect 10183 24701 10195 24735
rect 10137 24695 10195 24701
rect 10597 24735 10655 24741
rect 10597 24701 10609 24735
rect 10643 24732 10655 24735
rect 11057 24735 11115 24741
rect 11057 24732 11069 24735
rect 10643 24704 11069 24732
rect 10643 24701 10655 24704
rect 10597 24695 10655 24701
rect 11057 24701 11069 24704
rect 11103 24732 11115 24735
rect 11330 24732 11336 24744
rect 11103 24704 11336 24732
rect 11103 24701 11115 24704
rect 11057 24695 11115 24701
rect 11330 24692 11336 24704
rect 11388 24692 11394 24744
rect 11514 24692 11520 24744
rect 11572 24732 11578 24744
rect 11885 24735 11943 24741
rect 11885 24732 11897 24735
rect 11572 24704 11897 24732
rect 11572 24692 11578 24704
rect 11885 24701 11897 24704
rect 11931 24701 11943 24735
rect 11885 24695 11943 24701
rect 11974 24692 11980 24744
rect 12032 24692 12038 24744
rect 12069 24735 12127 24741
rect 12069 24701 12081 24735
rect 12115 24732 12127 24735
rect 12342 24732 12348 24744
rect 12115 24704 12348 24732
rect 12115 24701 12127 24704
rect 12069 24695 12127 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 9916 24568 10088 24596
rect 9916 24556 9922 24568
rect 11698 24556 11704 24608
rect 11756 24556 11762 24608
rect 552 24506 12604 24528
rect 552 24454 4322 24506
rect 4374 24454 4386 24506
rect 4438 24454 4450 24506
rect 4502 24454 4514 24506
rect 4566 24454 4578 24506
rect 4630 24454 10722 24506
rect 10774 24454 10786 24506
rect 10838 24454 10850 24506
rect 10902 24454 10914 24506
rect 10966 24454 10978 24506
rect 11030 24454 12604 24506
rect 552 24432 12604 24454
rect 750 24352 756 24404
rect 808 24392 814 24404
rect 934 24392 940 24404
rect 808 24364 940 24392
rect 808 24352 814 24364
rect 934 24352 940 24364
rect 992 24392 998 24404
rect 2409 24395 2467 24401
rect 2409 24392 2421 24395
rect 992 24364 2421 24392
rect 992 24352 998 24364
rect 2409 24361 2421 24364
rect 2455 24361 2467 24395
rect 2409 24355 2467 24361
rect 3605 24395 3663 24401
rect 3605 24361 3617 24395
rect 3651 24361 3663 24395
rect 3605 24355 3663 24361
rect 1394 24324 1400 24336
rect 860 24296 1400 24324
rect 860 24265 888 24296
rect 1394 24284 1400 24296
rect 1452 24324 1458 24336
rect 1452 24296 2820 24324
rect 1452 24284 1458 24296
rect 2792 24268 2820 24296
rect 3510 24284 3516 24336
rect 3568 24324 3574 24336
rect 3620 24324 3648 24355
rect 4154 24352 4160 24404
rect 4212 24392 4218 24404
rect 4614 24392 4620 24404
rect 4212 24364 4620 24392
rect 4212 24352 4218 24364
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 4801 24395 4859 24401
rect 4801 24361 4813 24395
rect 4847 24392 4859 24395
rect 5074 24392 5080 24404
rect 4847 24364 5080 24392
rect 4847 24361 4859 24364
rect 4801 24355 4859 24361
rect 5074 24352 5080 24364
rect 5132 24352 5138 24404
rect 7006 24392 7012 24404
rect 5828 24364 7012 24392
rect 4985 24327 5043 24333
rect 4985 24324 4997 24327
rect 3568 24296 4997 24324
rect 3568 24284 3574 24296
rect 845 24259 903 24265
rect 845 24225 857 24259
rect 891 24225 903 24259
rect 845 24219 903 24225
rect 1112 24259 1170 24265
rect 1112 24225 1124 24259
rect 1158 24256 1170 24259
rect 1486 24256 1492 24268
rect 1158 24228 1492 24256
rect 1158 24225 1170 24228
rect 1112 24219 1170 24225
rect 1486 24216 1492 24228
rect 1544 24256 1550 24268
rect 1946 24256 1952 24268
rect 1544 24228 1952 24256
rect 1544 24216 1550 24228
rect 1946 24216 1952 24228
rect 2004 24216 2010 24268
rect 2593 24259 2651 24265
rect 2593 24225 2605 24259
rect 2639 24225 2651 24259
rect 2593 24219 2651 24225
rect 2608 24188 2636 24219
rect 2774 24216 2780 24268
rect 2832 24216 2838 24268
rect 3329 24259 3387 24265
rect 3329 24225 3341 24259
rect 3375 24256 3387 24259
rect 3602 24256 3608 24268
rect 3375 24228 3608 24256
rect 3375 24225 3387 24228
rect 3329 24219 3387 24225
rect 3602 24216 3608 24228
rect 3660 24216 3666 24268
rect 3694 24216 3700 24268
rect 3752 24216 3758 24268
rect 3786 24216 3792 24268
rect 3844 24216 3850 24268
rect 3988 24265 4016 24296
rect 4985 24293 4997 24296
rect 5031 24324 5043 24327
rect 5031 24296 5488 24324
rect 5031 24293 5043 24296
rect 4985 24287 5043 24293
rect 3973 24259 4031 24265
rect 3973 24225 3985 24259
rect 4019 24225 4031 24259
rect 3973 24219 4031 24225
rect 4062 24216 4068 24268
rect 4120 24256 4126 24268
rect 4157 24259 4215 24265
rect 4157 24256 4169 24259
rect 4120 24228 4169 24256
rect 4120 24216 4126 24228
rect 4157 24225 4169 24228
rect 4203 24225 4215 24259
rect 4157 24219 4215 24225
rect 4246 24216 4252 24268
rect 4304 24256 4310 24268
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 4304 24228 4353 24256
rect 4304 24216 4310 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 5169 24259 5227 24265
rect 5169 24225 5181 24259
rect 5215 24256 5227 24259
rect 5350 24256 5356 24268
rect 5215 24228 5356 24256
rect 5215 24225 5227 24228
rect 5169 24219 5227 24225
rect 5350 24216 5356 24228
rect 5408 24216 5414 24268
rect 5460 24265 5488 24296
rect 5445 24259 5503 24265
rect 5445 24225 5457 24259
rect 5491 24225 5503 24259
rect 5445 24219 5503 24225
rect 5537 24259 5595 24265
rect 5537 24225 5549 24259
rect 5583 24225 5595 24259
rect 5537 24219 5595 24225
rect 3513 24191 3571 24197
rect 2608 24160 2774 24188
rect 2746 24120 2774 24160
rect 3513 24157 3525 24191
rect 3559 24157 3571 24191
rect 3804 24188 3832 24216
rect 5552 24188 5580 24219
rect 5626 24216 5632 24268
rect 5684 24256 5690 24268
rect 5828 24265 5856 24364
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 7558 24352 7564 24404
rect 7616 24352 7622 24404
rect 7650 24352 7656 24404
rect 7708 24392 7714 24404
rect 7926 24392 7932 24404
rect 7708 24364 7932 24392
rect 7708 24352 7714 24364
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 8389 24395 8447 24401
rect 8389 24361 8401 24395
rect 8435 24392 8447 24395
rect 8478 24392 8484 24404
rect 8435 24364 8484 24392
rect 8435 24361 8447 24364
rect 8389 24355 8447 24361
rect 8478 24352 8484 24364
rect 8536 24352 8542 24404
rect 9214 24352 9220 24404
rect 9272 24352 9278 24404
rect 9398 24352 9404 24404
rect 9456 24392 9462 24404
rect 11882 24392 11888 24404
rect 9456 24364 11888 24392
rect 9456 24352 9462 24364
rect 11882 24352 11888 24364
rect 11940 24392 11946 24404
rect 12434 24392 12440 24404
rect 11940 24364 12440 24392
rect 11940 24352 11946 24364
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 6733 24327 6791 24333
rect 6733 24324 6745 24327
rect 5920 24296 6745 24324
rect 5813 24259 5871 24265
rect 5813 24256 5825 24259
rect 5684 24228 5825 24256
rect 5684 24216 5690 24228
rect 5813 24225 5825 24228
rect 5859 24225 5871 24259
rect 5813 24219 5871 24225
rect 5920 24188 5948 24296
rect 6472 24268 6500 24296
rect 6733 24293 6745 24296
rect 6779 24293 6791 24327
rect 6733 24287 6791 24293
rect 6917 24327 6975 24333
rect 6917 24293 6929 24327
rect 6963 24324 6975 24327
rect 6963 24296 7696 24324
rect 6963 24293 6975 24296
rect 6917 24287 6975 24293
rect 5997 24259 6055 24265
rect 5997 24225 6009 24259
rect 6043 24225 6055 24259
rect 5997 24219 6055 24225
rect 3804 24160 4200 24188
rect 5552 24160 5948 24188
rect 3513 24151 3571 24157
rect 3421 24123 3479 24129
rect 3421 24120 3433 24123
rect 2746 24092 3433 24120
rect 3421 24089 3433 24092
rect 3467 24089 3479 24123
rect 3528 24120 3556 24151
rect 4172 24132 4200 24160
rect 3878 24120 3884 24132
rect 3528 24092 3884 24120
rect 3421 24083 3479 24089
rect 3878 24080 3884 24092
rect 3936 24080 3942 24132
rect 4154 24080 4160 24132
rect 4212 24080 4218 24132
rect 4614 24080 4620 24132
rect 4672 24080 4678 24132
rect 5718 24080 5724 24132
rect 5776 24120 5782 24132
rect 6012 24120 6040 24219
rect 6270 24216 6276 24268
rect 6328 24216 6334 24268
rect 6454 24216 6460 24268
rect 6512 24216 6518 24268
rect 6546 24216 6552 24268
rect 6604 24216 6610 24268
rect 6638 24216 6644 24268
rect 6696 24256 6702 24268
rect 7009 24259 7067 24265
rect 7009 24256 7021 24259
rect 6696 24228 7021 24256
rect 6696 24216 6702 24228
rect 7009 24225 7021 24228
rect 7055 24225 7067 24259
rect 7009 24219 7067 24225
rect 7193 24259 7251 24265
rect 7193 24225 7205 24259
rect 7239 24225 7251 24259
rect 7193 24219 7251 24225
rect 6086 24148 6092 24200
rect 6144 24188 6150 24200
rect 6181 24191 6239 24197
rect 6181 24188 6193 24191
rect 6144 24160 6193 24188
rect 6144 24148 6150 24160
rect 6181 24157 6193 24160
rect 6227 24157 6239 24191
rect 6564 24188 6592 24216
rect 7208 24188 7236 24219
rect 7282 24216 7288 24268
rect 7340 24216 7346 24268
rect 7377 24259 7435 24265
rect 7377 24225 7389 24259
rect 7423 24258 7435 24259
rect 7466 24258 7472 24268
rect 7423 24230 7472 24258
rect 7423 24225 7435 24230
rect 7377 24219 7435 24225
rect 7466 24216 7472 24230
rect 7524 24216 7530 24268
rect 7668 24265 7696 24296
rect 8018 24284 8024 24336
rect 8076 24324 8082 24336
rect 8076 24296 9720 24324
rect 8076 24284 8082 24296
rect 7653 24259 7711 24265
rect 7653 24225 7665 24259
rect 7699 24225 7711 24259
rect 7653 24219 7711 24225
rect 7834 24216 7840 24268
rect 7892 24216 7898 24268
rect 8202 24216 8208 24268
rect 8260 24216 8266 24268
rect 8481 24259 8539 24265
rect 8481 24225 8493 24259
rect 8527 24225 8539 24259
rect 8481 24219 8539 24225
rect 6564 24160 7236 24188
rect 6181 24151 6239 24157
rect 5776 24092 6040 24120
rect 6196 24120 6224 24151
rect 7926 24148 7932 24200
rect 7984 24148 7990 24200
rect 8018 24148 8024 24200
rect 8076 24188 8082 24200
rect 8496 24188 8524 24219
rect 8570 24216 8576 24268
rect 8628 24256 8634 24268
rect 9125 24259 9183 24265
rect 9125 24256 9137 24259
rect 8628 24228 9137 24256
rect 8628 24216 8634 24228
rect 9125 24225 9137 24228
rect 9171 24225 9183 24259
rect 9125 24219 9183 24225
rect 8076 24160 8524 24188
rect 9140 24188 9168 24219
rect 9306 24216 9312 24268
rect 9364 24216 9370 24268
rect 9692 24265 9720 24296
rect 10594 24284 10600 24336
rect 10652 24324 10658 24336
rect 11238 24324 11244 24336
rect 10652 24296 11244 24324
rect 10652 24284 10658 24296
rect 9677 24259 9735 24265
rect 9677 24225 9689 24259
rect 9723 24225 9735 24259
rect 9677 24219 9735 24225
rect 9950 24216 9956 24268
rect 10008 24256 10014 24268
rect 10229 24259 10287 24265
rect 10229 24256 10241 24259
rect 10008 24228 10241 24256
rect 10008 24216 10014 24228
rect 10229 24225 10241 24228
rect 10275 24225 10287 24259
rect 10229 24219 10287 24225
rect 10318 24216 10324 24268
rect 10376 24216 10382 24268
rect 10413 24259 10471 24265
rect 10413 24225 10425 24259
rect 10459 24256 10471 24259
rect 11054 24256 11060 24268
rect 10459 24228 11060 24256
rect 10459 24225 10471 24228
rect 10413 24219 10471 24225
rect 11054 24216 11060 24228
rect 11112 24216 11118 24268
rect 11164 24265 11192 24296
rect 11238 24284 11244 24296
rect 11296 24284 11302 24336
rect 11149 24259 11207 24265
rect 11149 24225 11161 24259
rect 11195 24225 11207 24259
rect 11149 24219 11207 24225
rect 11606 24216 11612 24268
rect 11664 24216 11670 24268
rect 11793 24259 11851 24265
rect 11793 24225 11805 24259
rect 11839 24256 11851 24259
rect 12066 24256 12072 24268
rect 11839 24228 12072 24256
rect 11839 24225 11851 24228
rect 11793 24219 11851 24225
rect 12066 24216 12072 24228
rect 12124 24216 12130 24268
rect 9582 24188 9588 24200
rect 9140 24160 9588 24188
rect 8076 24148 8082 24160
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 7006 24120 7012 24132
rect 6196 24092 7012 24120
rect 5776 24080 5782 24092
rect 7006 24080 7012 24092
rect 7064 24080 7070 24132
rect 7466 24080 7472 24132
rect 7524 24120 7530 24132
rect 8573 24123 8631 24129
rect 8573 24120 8585 24123
rect 7524 24092 8585 24120
rect 7524 24080 7530 24092
rect 8573 24089 8585 24092
rect 8619 24089 8631 24123
rect 8573 24083 8631 24089
rect 9490 24080 9496 24132
rect 9548 24120 9554 24132
rect 10045 24123 10103 24129
rect 10045 24120 10057 24123
rect 9548 24092 10057 24120
rect 9548 24080 9554 24092
rect 10045 24089 10057 24092
rect 10091 24089 10103 24123
rect 10336 24120 10364 24216
rect 10505 24191 10563 24197
rect 10505 24157 10517 24191
rect 10551 24188 10563 24191
rect 10965 24191 11023 24197
rect 10965 24188 10977 24191
rect 10551 24160 10977 24188
rect 10551 24157 10563 24160
rect 10505 24151 10563 24157
rect 10965 24157 10977 24160
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 11330 24148 11336 24200
rect 11388 24148 11394 24200
rect 11701 24191 11759 24197
rect 11701 24157 11713 24191
rect 11747 24157 11759 24191
rect 11701 24151 11759 24157
rect 11885 24191 11943 24197
rect 11885 24157 11897 24191
rect 11931 24188 11943 24191
rect 11974 24188 11980 24200
rect 11931 24160 11980 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 10686 24120 10692 24132
rect 10336 24092 10692 24120
rect 10045 24083 10103 24089
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 11716 24120 11744 24151
rect 11974 24148 11980 24160
rect 12032 24148 12038 24200
rect 11716 24092 11928 24120
rect 11900 24064 11928 24092
rect 2222 24012 2228 24064
rect 2280 24012 2286 24064
rect 4062 24012 4068 24064
rect 4120 24012 4126 24064
rect 4522 24012 4528 24064
rect 4580 24052 4586 24064
rect 4890 24052 4896 24064
rect 4580 24024 4896 24052
rect 4580 24012 4586 24024
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 5353 24055 5411 24061
rect 5353 24021 5365 24055
rect 5399 24052 5411 24055
rect 5442 24052 5448 24064
rect 5399 24024 5448 24052
rect 5399 24021 5411 24024
rect 5353 24015 5411 24021
rect 5442 24012 5448 24024
rect 5500 24012 5506 24064
rect 6086 24012 6092 24064
rect 6144 24052 6150 24064
rect 6365 24055 6423 24061
rect 6365 24052 6377 24055
rect 6144 24024 6377 24052
rect 6144 24012 6150 24024
rect 6365 24021 6377 24024
rect 6411 24021 6423 24055
rect 6365 24015 6423 24021
rect 6638 24012 6644 24064
rect 6696 24052 6702 24064
rect 8294 24052 8300 24064
rect 6696 24024 8300 24052
rect 6696 24012 6702 24024
rect 8294 24012 8300 24024
rect 8352 24012 8358 24064
rect 9858 24012 9864 24064
rect 9916 24012 9922 24064
rect 11422 24012 11428 24064
rect 11480 24012 11486 24064
rect 11882 24012 11888 24064
rect 11940 24012 11946 24064
rect 552 23962 12604 23984
rect 552 23910 3662 23962
rect 3714 23910 3726 23962
rect 3778 23910 3790 23962
rect 3842 23910 3854 23962
rect 3906 23910 3918 23962
rect 3970 23910 10062 23962
rect 10114 23910 10126 23962
rect 10178 23910 10190 23962
rect 10242 23910 10254 23962
rect 10306 23910 10318 23962
rect 10370 23910 12604 23962
rect 552 23888 12604 23910
rect 4338 23808 4344 23860
rect 4396 23848 4402 23860
rect 5074 23848 5080 23860
rect 4396 23820 5080 23848
rect 4396 23808 4402 23820
rect 5074 23808 5080 23820
rect 5132 23848 5138 23860
rect 5537 23851 5595 23857
rect 5537 23848 5549 23851
rect 5132 23820 5549 23848
rect 5132 23808 5138 23820
rect 5537 23817 5549 23820
rect 5583 23848 5595 23851
rect 5626 23848 5632 23860
rect 5583 23820 5632 23848
rect 5583 23817 5595 23820
rect 5537 23811 5595 23817
rect 5626 23808 5632 23820
rect 5684 23808 5690 23860
rect 5813 23851 5871 23857
rect 5813 23817 5825 23851
rect 5859 23848 5871 23851
rect 6546 23848 6552 23860
rect 5859 23820 6552 23848
rect 5859 23817 5871 23820
rect 5813 23811 5871 23817
rect 6546 23808 6552 23820
rect 6604 23808 6610 23860
rect 7558 23808 7564 23860
rect 7616 23848 7622 23860
rect 8018 23848 8024 23860
rect 7616 23820 8024 23848
rect 7616 23808 7622 23820
rect 8018 23808 8024 23820
rect 8076 23808 8082 23860
rect 10137 23851 10195 23857
rect 10137 23817 10149 23851
rect 10183 23848 10195 23851
rect 10502 23848 10508 23860
rect 10183 23820 10508 23848
rect 10183 23817 10195 23820
rect 10137 23811 10195 23817
rect 10502 23808 10508 23820
rect 10560 23808 10566 23860
rect 11514 23808 11520 23860
rect 11572 23848 11578 23860
rect 11572 23820 11928 23848
rect 11572 23808 11578 23820
rect 1026 23740 1032 23792
rect 1084 23780 1090 23792
rect 1210 23780 1216 23792
rect 1084 23752 1216 23780
rect 1084 23740 1090 23752
rect 1210 23740 1216 23752
rect 1268 23740 1274 23792
rect 3053 23783 3111 23789
rect 3053 23749 3065 23783
rect 3099 23749 3111 23783
rect 3053 23743 3111 23749
rect 842 23672 848 23724
rect 900 23712 906 23724
rect 1670 23712 1676 23724
rect 900 23684 1676 23712
rect 900 23672 906 23684
rect 1670 23672 1676 23684
rect 1728 23672 1734 23724
rect 3068 23712 3096 23743
rect 4246 23740 4252 23792
rect 4304 23780 4310 23792
rect 4433 23783 4491 23789
rect 4433 23780 4445 23783
rect 4304 23752 4445 23780
rect 4304 23740 4310 23752
rect 4433 23749 4445 23752
rect 4479 23749 4491 23783
rect 4433 23743 4491 23749
rect 4614 23740 4620 23792
rect 4672 23780 4678 23792
rect 4890 23780 4896 23792
rect 4672 23752 4896 23780
rect 4672 23740 4678 23752
rect 4890 23740 4896 23752
rect 4948 23740 4954 23792
rect 5350 23780 5356 23792
rect 5092 23752 5356 23780
rect 3510 23712 3516 23724
rect 3068 23684 3516 23712
rect 3510 23672 3516 23684
rect 3568 23712 3574 23724
rect 3697 23715 3755 23721
rect 3697 23712 3709 23715
rect 3568 23684 3709 23712
rect 3568 23672 3574 23684
rect 3697 23681 3709 23684
rect 3743 23681 3755 23715
rect 3697 23675 3755 23681
rect 3881 23715 3939 23721
rect 3881 23681 3893 23715
rect 3927 23712 3939 23715
rect 4798 23712 4804 23724
rect 3927 23684 4804 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 934 23604 940 23656
rect 992 23644 998 23656
rect 1121 23647 1179 23653
rect 1121 23644 1133 23647
rect 992 23616 1133 23644
rect 992 23604 998 23616
rect 1121 23613 1133 23616
rect 1167 23644 1179 23647
rect 1210 23644 1216 23656
rect 1167 23616 1216 23644
rect 1167 23613 1179 23616
rect 1121 23607 1179 23613
rect 1210 23604 1216 23616
rect 1268 23604 1274 23656
rect 1302 23604 1308 23656
rect 1360 23644 1366 23656
rect 1397 23647 1455 23653
rect 1397 23644 1409 23647
rect 1360 23616 1409 23644
rect 1360 23604 1366 23616
rect 1397 23613 1409 23616
rect 1443 23644 1455 23647
rect 1486 23644 1492 23656
rect 1443 23616 1492 23644
rect 1443 23613 1455 23616
rect 1397 23607 1455 23613
rect 1486 23604 1492 23616
rect 1544 23604 1550 23656
rect 3050 23604 3056 23656
rect 3108 23644 3114 23656
rect 3108 23616 3372 23644
rect 3108 23604 3114 23616
rect 1940 23579 1998 23585
rect 1940 23545 1952 23579
rect 1986 23576 1998 23579
rect 1986 23548 3280 23576
rect 1986 23545 1998 23548
rect 1940 23539 1998 23545
rect 3252 23517 3280 23548
rect 3237 23511 3295 23517
rect 3237 23477 3249 23511
rect 3283 23477 3295 23511
rect 3344 23508 3372 23616
rect 3418 23604 3424 23656
rect 3476 23644 3482 23656
rect 3605 23647 3663 23653
rect 3605 23644 3617 23647
rect 3476 23616 3617 23644
rect 3476 23604 3482 23616
rect 3605 23613 3617 23616
rect 3651 23613 3663 23647
rect 3712 23644 3740 23675
rect 4798 23672 4804 23684
rect 4856 23672 4862 23724
rect 4065 23647 4123 23653
rect 4065 23644 4077 23647
rect 3712 23616 4077 23644
rect 3605 23607 3663 23613
rect 4065 23613 4077 23616
rect 4111 23613 4123 23647
rect 4065 23607 4123 23613
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 4522 23644 4528 23656
rect 4295 23616 4528 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4522 23604 4528 23616
rect 4580 23604 4586 23656
rect 4614 23604 4620 23656
rect 4672 23604 4678 23656
rect 5092 23653 5120 23752
rect 5350 23740 5356 23752
rect 5408 23740 5414 23792
rect 7190 23780 7196 23792
rect 6932 23752 7196 23780
rect 5261 23715 5319 23721
rect 5261 23681 5273 23715
rect 5307 23712 5319 23715
rect 5534 23712 5540 23724
rect 5307 23684 5540 23712
rect 5307 23681 5319 23684
rect 5261 23675 5319 23681
rect 5534 23672 5540 23684
rect 5592 23672 5598 23724
rect 6086 23712 6092 23724
rect 5736 23684 6092 23712
rect 4893 23647 4951 23653
rect 4893 23613 4905 23647
rect 4939 23613 4951 23647
rect 4893 23607 4951 23613
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23613 5135 23647
rect 5077 23607 5135 23613
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23613 5227 23647
rect 5169 23607 5227 23613
rect 4338 23536 4344 23588
rect 4396 23536 4402 23588
rect 4540 23576 4568 23604
rect 4908 23576 4936 23607
rect 4540 23548 4936 23576
rect 4982 23536 4988 23588
rect 5040 23576 5046 23588
rect 5184 23576 5212 23607
rect 5350 23604 5356 23656
rect 5408 23604 5414 23656
rect 5736 23653 5764 23684
rect 6086 23672 6092 23684
rect 6144 23672 6150 23724
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6638 23721 6644 23724
rect 6457 23715 6515 23721
rect 6457 23712 6469 23715
rect 6328 23684 6469 23712
rect 6328 23672 6334 23684
rect 6457 23681 6469 23684
rect 6503 23681 6515 23715
rect 6457 23675 6515 23681
rect 6616 23715 6644 23721
rect 6616 23681 6628 23715
rect 6616 23675 6644 23681
rect 6638 23672 6644 23675
rect 6696 23672 6702 23724
rect 6733 23715 6791 23721
rect 6733 23681 6745 23715
rect 6779 23712 6791 23715
rect 6932 23712 6960 23752
rect 7190 23740 7196 23752
rect 7248 23780 7254 23792
rect 7466 23780 7472 23792
rect 7248 23752 7472 23780
rect 7248 23740 7254 23752
rect 7466 23740 7472 23752
rect 7524 23740 7530 23792
rect 8202 23740 8208 23792
rect 8260 23780 8266 23792
rect 10594 23780 10600 23792
rect 8260 23752 10600 23780
rect 8260 23740 8266 23752
rect 10594 23740 10600 23752
rect 10652 23740 10658 23792
rect 11790 23740 11796 23792
rect 11848 23740 11854 23792
rect 11900 23780 11928 23820
rect 11974 23808 11980 23860
rect 12032 23808 12038 23860
rect 12158 23780 12164 23792
rect 11900 23752 12164 23780
rect 12158 23740 12164 23752
rect 12216 23780 12222 23792
rect 12618 23780 12624 23792
rect 12216 23752 12624 23780
rect 12216 23740 12222 23752
rect 12618 23740 12624 23752
rect 12676 23740 12682 23792
rect 6779 23684 6960 23712
rect 7009 23715 7067 23721
rect 6779 23681 6791 23684
rect 6733 23675 6791 23681
rect 7009 23681 7021 23715
rect 7055 23712 7067 23715
rect 7098 23712 7104 23724
rect 7055 23684 7104 23712
rect 7055 23681 7067 23684
rect 7009 23675 7067 23681
rect 7098 23672 7104 23684
rect 7156 23672 7162 23724
rect 7484 23684 10180 23712
rect 7484 23653 7512 23684
rect 5721 23647 5779 23653
rect 5721 23613 5733 23647
rect 5767 23613 5779 23647
rect 5721 23607 5779 23613
rect 7469 23647 7527 23653
rect 7469 23613 7481 23647
rect 7515 23613 7527 23647
rect 7469 23607 7527 23613
rect 7650 23604 7656 23656
rect 7708 23604 7714 23656
rect 10045 23647 10103 23653
rect 10045 23613 10057 23647
rect 10091 23613 10103 23647
rect 10045 23607 10103 23613
rect 5040 23548 5212 23576
rect 5040 23536 5046 23548
rect 3418 23508 3424 23520
rect 3344 23480 3424 23508
rect 3237 23471 3295 23477
rect 3418 23468 3424 23480
rect 3476 23468 3482 23520
rect 4157 23511 4215 23517
rect 4157 23477 4169 23511
rect 4203 23508 4215 23511
rect 4798 23508 4804 23520
rect 4203 23480 4804 23508
rect 4203 23477 4215 23480
rect 4157 23471 4215 23477
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 5077 23511 5135 23517
rect 5077 23477 5089 23511
rect 5123 23508 5135 23511
rect 5626 23508 5632 23520
rect 5123 23480 5632 23508
rect 5123 23477 5135 23480
rect 5077 23471 5135 23477
rect 5626 23468 5632 23480
rect 5684 23468 5690 23520
rect 10060 23508 10088 23607
rect 10152 23576 10180 23684
rect 11238 23672 11244 23724
rect 11296 23712 11302 23724
rect 11808 23712 11836 23740
rect 11296 23684 12296 23712
rect 11296 23672 11302 23684
rect 10229 23647 10287 23653
rect 10229 23613 10241 23647
rect 10275 23644 10287 23647
rect 10318 23644 10324 23656
rect 10275 23616 10324 23644
rect 10275 23613 10287 23616
rect 10229 23607 10287 23613
rect 10318 23604 10324 23616
rect 10376 23644 10382 23656
rect 10686 23644 10692 23656
rect 10376 23616 10692 23644
rect 10376 23604 10382 23616
rect 10686 23604 10692 23616
rect 10744 23604 10750 23656
rect 11330 23604 11336 23656
rect 11388 23644 11394 23656
rect 11701 23647 11759 23653
rect 11701 23644 11713 23647
rect 11388 23616 11713 23644
rect 11388 23604 11394 23616
rect 11701 23613 11713 23616
rect 11747 23613 11759 23647
rect 11701 23607 11759 23613
rect 11793 23647 11851 23653
rect 11793 23613 11805 23647
rect 11839 23644 11851 23647
rect 12069 23647 12127 23653
rect 12069 23644 12081 23647
rect 11839 23616 12081 23644
rect 11839 23613 11851 23616
rect 11793 23607 11851 23613
rect 12069 23613 12081 23616
rect 12115 23644 12127 23647
rect 12158 23644 12164 23656
rect 12115 23616 12164 23644
rect 12115 23613 12127 23616
rect 12069 23607 12127 23613
rect 11514 23576 11520 23588
rect 10152 23548 11520 23576
rect 11514 23536 11520 23548
rect 11572 23536 11578 23588
rect 11716 23576 11744 23607
rect 12158 23604 12164 23616
rect 12216 23604 12222 23656
rect 12268 23653 12296 23684
rect 12253 23647 12311 23653
rect 12253 23613 12265 23647
rect 12299 23613 12311 23647
rect 12253 23607 12311 23613
rect 11974 23576 11980 23588
rect 11716 23548 11980 23576
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 12526 23576 12532 23588
rect 12084 23548 12532 23576
rect 11054 23508 11060 23520
rect 10060 23480 11060 23508
rect 11054 23468 11060 23480
rect 11112 23508 11118 23520
rect 12084 23508 12112 23548
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 11112 23480 12112 23508
rect 11112 23468 11118 23480
rect 12158 23468 12164 23520
rect 12216 23468 12222 23520
rect 552 23418 12604 23440
rect 552 23366 4322 23418
rect 4374 23366 4386 23418
rect 4438 23366 4450 23418
rect 4502 23366 4514 23418
rect 4566 23366 4578 23418
rect 4630 23366 10722 23418
rect 10774 23366 10786 23418
rect 10838 23366 10850 23418
rect 10902 23366 10914 23418
rect 10966 23366 10978 23418
rect 11030 23366 12604 23418
rect 552 23344 12604 23366
rect 382 23264 388 23316
rect 440 23304 446 23316
rect 1486 23304 1492 23316
rect 440 23276 1492 23304
rect 440 23264 446 23276
rect 1486 23264 1492 23276
rect 1544 23264 1550 23316
rect 1762 23264 1768 23316
rect 1820 23304 1826 23316
rect 2225 23307 2283 23313
rect 2225 23304 2237 23307
rect 1820 23276 2237 23304
rect 1820 23264 1826 23276
rect 2225 23273 2237 23276
rect 2271 23273 2283 23307
rect 5074 23304 5080 23316
rect 2225 23267 2283 23273
rect 4724 23276 5080 23304
rect 2774 23236 2780 23248
rect 860 23208 2780 23236
rect 860 23177 888 23208
rect 2774 23196 2780 23208
rect 2832 23196 2838 23248
rect 3234 23196 3240 23248
rect 3292 23236 3298 23248
rect 4430 23236 4436 23248
rect 3292 23208 4436 23236
rect 3292 23196 3298 23208
rect 4430 23196 4436 23208
rect 4488 23196 4494 23248
rect 845 23171 903 23177
rect 845 23137 857 23171
rect 891 23137 903 23171
rect 845 23131 903 23137
rect 934 23128 940 23180
rect 992 23168 998 23180
rect 1118 23177 1124 23180
rect 1112 23168 1124 23177
rect 992 23140 1124 23168
rect 992 23128 998 23140
rect 1112 23131 1124 23140
rect 1118 23128 1124 23131
rect 1176 23128 1182 23180
rect 2314 23128 2320 23180
rect 2372 23128 2378 23180
rect 2498 23168 2504 23180
rect 2424 23140 2504 23168
rect 2424 22976 2452 23140
rect 2498 23128 2504 23140
rect 2556 23128 2562 23180
rect 4246 23128 4252 23180
rect 4304 23168 4310 23180
rect 4724 23177 4752 23276
rect 5074 23264 5080 23276
rect 5132 23264 5138 23316
rect 6086 23304 6092 23316
rect 5184 23276 6092 23304
rect 5184 23236 5212 23276
rect 6086 23264 6092 23276
rect 6144 23264 6150 23316
rect 7742 23304 7748 23316
rect 6472 23276 7748 23304
rect 5000 23208 5212 23236
rect 4525 23171 4583 23177
rect 4525 23168 4537 23171
rect 4304 23140 4537 23168
rect 4304 23128 4310 23140
rect 4525 23137 4537 23140
rect 4571 23137 4583 23171
rect 4525 23131 4583 23137
rect 4709 23171 4767 23177
rect 4709 23137 4721 23171
rect 4755 23137 4767 23171
rect 4709 23131 4767 23137
rect 4801 23171 4859 23177
rect 4801 23137 4813 23171
rect 4847 23168 4859 23171
rect 5000 23168 5028 23208
rect 5442 23196 5448 23248
rect 5500 23196 5506 23248
rect 5552 23208 6408 23236
rect 4847 23140 5028 23168
rect 4847 23137 4859 23140
rect 4801 23131 4859 23137
rect 5074 23128 5080 23180
rect 5132 23168 5138 23180
rect 5552 23168 5580 23208
rect 5132 23140 5580 23168
rect 5132 23128 5138 23140
rect 5626 23128 5632 23180
rect 5684 23168 5690 23180
rect 6380 23177 6408 23208
rect 5813 23171 5871 23177
rect 5813 23168 5825 23171
rect 5684 23140 5825 23168
rect 5684 23128 5690 23140
rect 5813 23137 5825 23140
rect 5859 23137 5871 23171
rect 5813 23131 5871 23137
rect 5997 23171 6055 23177
rect 5997 23137 6009 23171
rect 6043 23168 6055 23171
rect 6365 23171 6423 23177
rect 6043 23140 6316 23168
rect 6043 23137 6055 23140
rect 5997 23131 6055 23137
rect 4890 23060 4896 23112
rect 4948 23100 4954 23112
rect 5718 23100 5724 23112
rect 4948 23072 5724 23100
rect 4948 23060 4954 23072
rect 5718 23060 5724 23072
rect 5776 23100 5782 23112
rect 6012 23100 6040 23131
rect 5776 23072 6040 23100
rect 5776 23060 5782 23072
rect 6086 23060 6092 23112
rect 6144 23060 6150 23112
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23069 6239 23103
rect 6288 23100 6316 23140
rect 6365 23137 6377 23171
rect 6411 23137 6423 23171
rect 6365 23131 6423 23137
rect 6472 23100 6500 23276
rect 7742 23264 7748 23276
rect 7800 23264 7806 23316
rect 7926 23264 7932 23316
rect 7984 23304 7990 23316
rect 9398 23304 9404 23316
rect 7984 23276 9404 23304
rect 7984 23264 7990 23276
rect 6546 23196 6552 23248
rect 6604 23236 6610 23248
rect 7193 23239 7251 23245
rect 7193 23236 7205 23239
rect 6604 23208 7205 23236
rect 6604 23196 6610 23208
rect 7193 23205 7205 23208
rect 7239 23205 7251 23239
rect 7193 23199 7251 23205
rect 6733 23171 6791 23177
rect 6733 23137 6745 23171
rect 6779 23168 6791 23171
rect 6822 23168 6828 23180
rect 6779 23140 6828 23168
rect 6779 23137 6791 23140
rect 6733 23131 6791 23137
rect 6822 23128 6828 23140
rect 6880 23128 6886 23180
rect 6917 23171 6975 23177
rect 6917 23137 6929 23171
rect 6963 23137 6975 23171
rect 6917 23131 6975 23137
rect 6288 23072 6500 23100
rect 6181 23063 6239 23069
rect 5629 23035 5687 23041
rect 5629 23001 5641 23035
rect 5675 23032 5687 23035
rect 6196 23032 6224 23063
rect 6638 23032 6644 23044
rect 5675 23004 6644 23032
rect 5675 23001 5687 23004
rect 5629 22995 5687 23001
rect 6638 22992 6644 23004
rect 6696 22992 6702 23044
rect 6932 23032 6960 23131
rect 7006 23128 7012 23180
rect 7064 23128 7070 23180
rect 7377 23171 7435 23177
rect 7377 23137 7389 23171
rect 7423 23168 7435 23171
rect 7469 23171 7527 23177
rect 7469 23168 7481 23171
rect 7423 23140 7481 23168
rect 7423 23137 7435 23140
rect 7377 23131 7435 23137
rect 7469 23137 7481 23140
rect 7515 23137 7527 23171
rect 7469 23131 7527 23137
rect 7650 23128 7656 23180
rect 7708 23128 7714 23180
rect 7760 23168 7788 23264
rect 7837 23171 7895 23177
rect 7837 23168 7849 23171
rect 7760 23140 7849 23168
rect 7837 23137 7849 23140
rect 7883 23137 7895 23171
rect 7837 23131 7895 23137
rect 7926 23128 7932 23180
rect 7984 23128 7990 23180
rect 8036 23177 8064 23276
rect 9398 23264 9404 23276
rect 9456 23304 9462 23316
rect 9456 23276 10272 23304
rect 9456 23264 9462 23276
rect 8665 23239 8723 23245
rect 8665 23205 8677 23239
rect 8711 23236 8723 23239
rect 9030 23236 9036 23248
rect 8711 23208 9036 23236
rect 8711 23205 8723 23208
rect 8665 23199 8723 23205
rect 9030 23196 9036 23208
rect 9088 23196 9094 23248
rect 8021 23171 8079 23177
rect 8021 23137 8033 23171
rect 8067 23137 8079 23171
rect 8021 23131 8079 23137
rect 8294 23128 8300 23180
rect 8352 23128 8358 23180
rect 8573 23171 8631 23177
rect 8573 23137 8585 23171
rect 8619 23137 8631 23171
rect 8573 23131 8631 23137
rect 8849 23171 8907 23177
rect 8849 23137 8861 23171
rect 8895 23137 8907 23171
rect 8849 23131 8907 23137
rect 7024 23100 7052 23128
rect 7745 23103 7803 23109
rect 7024 23072 7696 23100
rect 7668 23044 7696 23072
rect 7745 23069 7757 23103
rect 7791 23100 7803 23103
rect 7944 23100 7972 23128
rect 8588 23100 8616 23131
rect 7791 23072 7972 23100
rect 8496 23072 8616 23100
rect 7791 23069 7803 23072
rect 7745 23063 7803 23069
rect 7098 23032 7104 23044
rect 6932 23004 7104 23032
rect 7098 22992 7104 23004
rect 7156 22992 7162 23044
rect 7650 22992 7656 23044
rect 7708 22992 7714 23044
rect 8110 23032 8116 23044
rect 7852 23004 8116 23032
rect 2406 22924 2412 22976
rect 2464 22924 2470 22976
rect 2501 22967 2559 22973
rect 2501 22933 2513 22967
rect 2547 22964 2559 22967
rect 2774 22964 2780 22976
rect 2547 22936 2780 22964
rect 2547 22933 2559 22936
rect 2501 22927 2559 22933
rect 2774 22924 2780 22936
rect 2832 22924 2838 22976
rect 3510 22924 3516 22976
rect 3568 22964 3574 22976
rect 5261 22967 5319 22973
rect 5261 22964 5273 22967
rect 3568 22936 5273 22964
rect 3568 22924 3574 22936
rect 5261 22933 5273 22936
rect 5307 22933 5319 22967
rect 5261 22927 5319 22933
rect 5718 22924 5724 22976
rect 5776 22964 5782 22976
rect 6549 22967 6607 22973
rect 6549 22964 6561 22967
rect 5776 22936 6561 22964
rect 5776 22924 5782 22936
rect 6549 22933 6561 22936
rect 6595 22933 6607 22967
rect 6549 22927 6607 22933
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7006 22964 7012 22976
rect 6963 22936 7012 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7006 22924 7012 22936
rect 7064 22924 7070 22976
rect 7116 22964 7144 22992
rect 7852 22964 7880 23004
rect 8110 22992 8116 23004
rect 8168 23032 8174 23044
rect 8496 23032 8524 23072
rect 8168 23004 8524 23032
rect 8168 22992 8174 23004
rect 8570 22992 8576 23044
rect 8628 23032 8634 23044
rect 8864 23032 8892 23131
rect 9214 23128 9220 23180
rect 9272 23168 9278 23180
rect 9309 23171 9367 23177
rect 9309 23168 9321 23171
rect 9272 23140 9321 23168
rect 9272 23128 9278 23140
rect 9309 23137 9321 23140
rect 9355 23137 9367 23171
rect 9309 23131 9367 23137
rect 9398 23128 9404 23180
rect 9456 23168 9462 23180
rect 10244 23177 10272 23276
rect 11238 23264 11244 23316
rect 11296 23304 11302 23316
rect 11333 23307 11391 23313
rect 11333 23304 11345 23307
rect 11296 23276 11345 23304
rect 11296 23264 11302 23276
rect 11333 23273 11345 23276
rect 11379 23273 11391 23307
rect 11333 23267 11391 23273
rect 11422 23264 11428 23316
rect 11480 23264 11486 23316
rect 11790 23264 11796 23316
rect 11848 23304 11854 23316
rect 12161 23307 12219 23313
rect 12161 23304 12173 23307
rect 11848 23276 12173 23304
rect 11848 23264 11854 23276
rect 12161 23273 12173 23276
rect 12207 23273 12219 23307
rect 12161 23267 12219 23273
rect 11440 23236 11468 23264
rect 11885 23239 11943 23245
rect 11885 23236 11897 23239
rect 10612 23208 11897 23236
rect 10045 23171 10103 23177
rect 10045 23168 10057 23171
rect 9456 23140 10057 23168
rect 9456 23128 9462 23140
rect 10045 23137 10057 23140
rect 10091 23137 10103 23171
rect 10045 23131 10103 23137
rect 10229 23171 10287 23177
rect 10229 23137 10241 23171
rect 10275 23137 10287 23171
rect 10229 23131 10287 23137
rect 10318 23128 10324 23180
rect 10376 23168 10382 23180
rect 10612 23177 10640 23208
rect 11885 23205 11897 23208
rect 11931 23205 11943 23239
rect 11885 23199 11943 23205
rect 10597 23171 10655 23177
rect 10376 23140 10548 23168
rect 10376 23128 10382 23140
rect 9582 23060 9588 23112
rect 9640 23060 9646 23112
rect 10520 23100 10548 23140
rect 10597 23137 10609 23171
rect 10643 23137 10655 23171
rect 10597 23131 10655 23137
rect 10686 23128 10692 23180
rect 10744 23168 10750 23180
rect 10781 23171 10839 23177
rect 10781 23168 10793 23171
rect 10744 23140 10793 23168
rect 10744 23128 10750 23140
rect 10781 23137 10793 23140
rect 10827 23137 10839 23171
rect 10781 23131 10839 23137
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 11149 23171 11207 23177
rect 11149 23168 11161 23171
rect 11020 23140 11161 23168
rect 11020 23128 11026 23140
rect 11149 23137 11161 23140
rect 11195 23137 11207 23171
rect 11149 23131 11207 23137
rect 11425 23171 11483 23177
rect 11425 23137 11437 23171
rect 11471 23137 11483 23171
rect 11425 23131 11483 23137
rect 11238 23100 11244 23112
rect 10520 23072 11244 23100
rect 11238 23060 11244 23072
rect 11296 23100 11302 23112
rect 11440 23100 11468 23131
rect 11514 23128 11520 23180
rect 11572 23128 11578 23180
rect 11701 23171 11759 23177
rect 11701 23137 11713 23171
rect 11747 23168 11759 23171
rect 11790 23168 11796 23180
rect 11747 23140 11796 23168
rect 11747 23137 11759 23140
rect 11701 23131 11759 23137
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 11977 23171 12035 23177
rect 11977 23137 11989 23171
rect 12023 23168 12035 23171
rect 12342 23168 12348 23180
rect 12023 23140 12348 23168
rect 12023 23137 12035 23140
rect 11977 23131 12035 23137
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 11296 23072 11468 23100
rect 11296 23060 11302 23072
rect 8628 23004 8892 23032
rect 9033 23035 9091 23041
rect 8628 22992 8634 23004
rect 9033 23001 9045 23035
rect 9079 23032 9091 23035
rect 9493 23035 9551 23041
rect 9493 23032 9505 23035
rect 9079 23004 9505 23032
rect 9079 23001 9091 23004
rect 9033 22995 9091 23001
rect 9493 23001 9505 23004
rect 9539 23001 9551 23035
rect 9493 22995 9551 23001
rect 10502 22992 10508 23044
rect 10560 23032 10566 23044
rect 10965 23035 11023 23041
rect 10965 23032 10977 23035
rect 10560 23004 10977 23032
rect 10560 22992 10566 23004
rect 10965 23001 10977 23004
rect 11011 23001 11023 23035
rect 10965 22995 11023 23001
rect 7116 22936 7880 22964
rect 7926 22924 7932 22976
rect 7984 22964 7990 22976
rect 8205 22967 8263 22973
rect 8205 22964 8217 22967
rect 7984 22936 8217 22964
rect 7984 22924 7990 22936
rect 8205 22933 8217 22936
rect 8251 22933 8263 22967
rect 8205 22927 8263 22933
rect 8294 22924 8300 22976
rect 8352 22964 8358 22976
rect 8389 22967 8447 22973
rect 8389 22964 8401 22967
rect 8352 22936 8401 22964
rect 8352 22924 8358 22936
rect 8389 22933 8401 22936
rect 8435 22933 8447 22967
rect 8389 22927 8447 22933
rect 8846 22924 8852 22976
rect 8904 22964 8910 22976
rect 9125 22967 9183 22973
rect 9125 22964 9137 22967
rect 8904 22936 9137 22964
rect 8904 22924 8910 22936
rect 9125 22933 9137 22936
rect 9171 22933 9183 22967
rect 9125 22927 9183 22933
rect 9674 22924 9680 22976
rect 9732 22964 9738 22976
rect 10137 22967 10195 22973
rect 10137 22964 10149 22967
rect 9732 22936 10149 22964
rect 9732 22924 9738 22936
rect 10137 22933 10149 22936
rect 10183 22964 10195 22967
rect 10410 22964 10416 22976
rect 10183 22936 10416 22964
rect 10183 22933 10195 22936
rect 10137 22927 10195 22933
rect 10410 22924 10416 22936
rect 10468 22924 10474 22976
rect 10594 22924 10600 22976
rect 10652 22924 10658 22976
rect 11698 22924 11704 22976
rect 11756 22964 11762 22976
rect 12342 22964 12348 22976
rect 11756 22936 12348 22964
rect 11756 22924 11762 22936
rect 12342 22924 12348 22936
rect 12400 22924 12406 22976
rect 552 22874 12604 22896
rect 552 22822 3662 22874
rect 3714 22822 3726 22874
rect 3778 22822 3790 22874
rect 3842 22822 3854 22874
rect 3906 22822 3918 22874
rect 3970 22822 10062 22874
rect 10114 22822 10126 22874
rect 10178 22822 10190 22874
rect 10242 22822 10254 22874
rect 10306 22822 10318 22874
rect 10370 22822 12604 22874
rect 552 22800 12604 22822
rect 2958 22720 2964 22772
rect 3016 22760 3022 22772
rect 3694 22760 3700 22772
rect 3016 22732 3700 22760
rect 3016 22720 3022 22732
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 3789 22763 3847 22769
rect 3789 22729 3801 22763
rect 3835 22760 3847 22763
rect 4062 22760 4068 22772
rect 3835 22732 4068 22760
rect 3835 22729 3847 22732
rect 3789 22723 3847 22729
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 4154 22720 4160 22772
rect 4212 22760 4218 22772
rect 4341 22763 4399 22769
rect 4341 22760 4353 22763
rect 4212 22732 4353 22760
rect 4212 22720 4218 22732
rect 4341 22729 4353 22732
rect 4387 22729 4399 22763
rect 4341 22723 4399 22729
rect 4448 22732 5120 22760
rect 1026 22652 1032 22704
rect 1084 22652 1090 22704
rect 2501 22695 2559 22701
rect 2501 22661 2513 22695
rect 2547 22692 2559 22695
rect 3142 22692 3148 22704
rect 2547 22664 3148 22692
rect 2547 22661 2559 22664
rect 2501 22655 2559 22661
rect 3142 22652 3148 22664
rect 3200 22652 3206 22704
rect 4448 22692 4476 22732
rect 3436 22664 4476 22692
rect 4893 22695 4951 22701
rect 1302 22584 1308 22636
rect 1360 22584 1366 22636
rect 2041 22627 2099 22633
rect 2041 22593 2053 22627
rect 2087 22624 2099 22627
rect 2222 22624 2228 22636
rect 2087 22596 2228 22624
rect 2087 22593 2099 22596
rect 2041 22587 2099 22593
rect 2222 22584 2228 22596
rect 2280 22584 2286 22636
rect 2590 22584 2596 22636
rect 2648 22624 2654 22636
rect 2648 22596 2820 22624
rect 2648 22584 2654 22596
rect 658 22516 664 22568
rect 716 22556 722 22568
rect 1213 22559 1271 22565
rect 1213 22556 1225 22559
rect 716 22528 1225 22556
rect 716 22516 722 22528
rect 1213 22525 1225 22528
rect 1259 22525 1271 22559
rect 1213 22519 1271 22525
rect 1578 22516 1584 22568
rect 1636 22556 1642 22568
rect 1765 22559 1823 22565
rect 1765 22556 1777 22559
rect 1636 22528 1777 22556
rect 1636 22516 1642 22528
rect 1765 22525 1777 22528
rect 1811 22525 1823 22559
rect 1765 22519 1823 22525
rect 1946 22516 1952 22568
rect 2004 22516 2010 22568
rect 2792 22565 2820 22596
rect 2685 22559 2743 22565
rect 2685 22525 2697 22559
rect 2731 22525 2743 22559
rect 2685 22519 2743 22525
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22525 2835 22559
rect 2777 22519 2835 22525
rect 2700 22488 2728 22519
rect 2958 22516 2964 22568
rect 3016 22516 3022 22568
rect 3053 22559 3111 22565
rect 3053 22525 3065 22559
rect 3099 22556 3111 22559
rect 3142 22556 3148 22568
rect 3099 22528 3148 22556
rect 3099 22525 3111 22528
rect 3053 22519 3111 22525
rect 3142 22516 3148 22528
rect 3200 22516 3206 22568
rect 3436 22565 3464 22664
rect 4893 22661 4905 22695
rect 4939 22692 4951 22695
rect 4982 22692 4988 22704
rect 4939 22664 4988 22692
rect 4939 22661 4951 22664
rect 4893 22655 4951 22661
rect 4982 22652 4988 22664
rect 5040 22652 5046 22704
rect 5092 22692 5120 22732
rect 5350 22720 5356 22772
rect 5408 22720 5414 22772
rect 6914 22720 6920 22772
rect 6972 22720 6978 22772
rect 8846 22720 8852 22772
rect 8904 22720 8910 22772
rect 9582 22720 9588 22772
rect 9640 22760 9646 22772
rect 10045 22763 10103 22769
rect 10045 22760 10057 22763
rect 9640 22732 10057 22760
rect 9640 22720 9646 22732
rect 10045 22729 10057 22732
rect 10091 22729 10103 22763
rect 10045 22723 10103 22729
rect 10962 22720 10968 22772
rect 11020 22720 11026 22772
rect 11425 22763 11483 22769
rect 11425 22729 11437 22763
rect 11471 22760 11483 22763
rect 11790 22760 11796 22772
rect 11471 22732 11796 22760
rect 11471 22729 11483 22732
rect 11425 22723 11483 22729
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 5092 22664 5672 22692
rect 3510 22584 3516 22636
rect 3568 22584 3574 22636
rect 4246 22624 4252 22636
rect 4172 22596 4252 22624
rect 4172 22565 4200 22596
rect 4246 22584 4252 22596
rect 4304 22584 4310 22636
rect 5258 22624 5264 22636
rect 4632 22596 5264 22624
rect 3421 22559 3479 22565
rect 3421 22525 3433 22559
rect 3467 22525 3479 22559
rect 3421 22519 3479 22525
rect 4065 22559 4123 22565
rect 4065 22525 4077 22559
rect 4111 22525 4123 22559
rect 4065 22519 4123 22525
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22525 4215 22559
rect 4157 22519 4215 22525
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22556 4491 22559
rect 4632 22556 4660 22596
rect 5258 22584 5264 22596
rect 5316 22584 5322 22636
rect 5644 22565 5672 22664
rect 6638 22652 6644 22704
rect 6696 22692 6702 22704
rect 7558 22692 7564 22704
rect 6696 22664 7564 22692
rect 6696 22652 6702 22664
rect 7558 22652 7564 22664
rect 7616 22652 7622 22704
rect 10594 22692 10600 22704
rect 9140 22664 10600 22692
rect 5718 22584 5724 22636
rect 5776 22584 5782 22636
rect 4479 22528 4660 22556
rect 5629 22559 5687 22565
rect 4479 22525 4491 22528
rect 4433 22519 4491 22525
rect 5629 22525 5641 22559
rect 5675 22556 5687 22559
rect 5675 22528 6316 22556
rect 5675 22525 5687 22528
rect 5629 22519 5687 22525
rect 3881 22491 3939 22497
rect 3881 22488 3893 22491
rect 2700 22460 3893 22488
rect 3881 22457 3893 22460
rect 3927 22457 3939 22491
rect 4080 22488 4108 22519
rect 3881 22451 3939 22457
rect 3988 22460 4108 22488
rect 4525 22491 4583 22497
rect 1026 22380 1032 22432
rect 1084 22420 1090 22432
rect 3988 22420 4016 22460
rect 4525 22457 4537 22491
rect 4571 22457 4583 22491
rect 4525 22451 4583 22457
rect 1084 22392 4016 22420
rect 1084 22380 1090 22392
rect 4062 22380 4068 22432
rect 4120 22420 4126 22432
rect 4540 22420 4568 22451
rect 4614 22448 4620 22500
rect 4672 22488 4678 22500
rect 6181 22491 6239 22497
rect 6181 22488 6193 22491
rect 4672 22460 6193 22488
rect 4672 22448 4678 22460
rect 6181 22457 6193 22460
rect 6227 22457 6239 22491
rect 6288 22488 6316 22528
rect 6362 22516 6368 22568
rect 6420 22556 6426 22568
rect 6730 22556 6736 22568
rect 6420 22528 6736 22556
rect 6420 22516 6426 22528
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 8202 22516 8208 22568
rect 8260 22516 8266 22568
rect 8386 22516 8392 22568
rect 8444 22516 8450 22568
rect 8757 22559 8815 22565
rect 8757 22525 8769 22559
rect 8803 22556 8815 22559
rect 8846 22556 8852 22568
rect 8803 22528 8852 22556
rect 8803 22525 8815 22528
rect 8757 22519 8815 22525
rect 8846 22516 8852 22528
rect 8904 22516 8910 22568
rect 9030 22516 9036 22568
rect 9088 22516 9094 22568
rect 9140 22565 9168 22664
rect 10594 22652 10600 22664
rect 10652 22652 10658 22704
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10134 22624 10140 22636
rect 9907 22596 10140 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10134 22584 10140 22596
rect 10192 22584 10198 22636
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 10870 22624 10876 22636
rect 10735 22596 10876 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 10870 22584 10876 22596
rect 10928 22584 10934 22636
rect 9125 22559 9183 22565
rect 9125 22525 9137 22559
rect 9171 22525 9183 22559
rect 9125 22519 9183 22525
rect 9214 22516 9220 22568
rect 9272 22556 9278 22568
rect 9582 22556 9588 22568
rect 9272 22528 9588 22556
rect 9272 22516 9278 22528
rect 9582 22516 9588 22528
rect 9640 22516 9646 22568
rect 9769 22559 9827 22565
rect 9769 22525 9781 22559
rect 9815 22556 9827 22559
rect 9950 22556 9956 22568
rect 9815 22528 9956 22556
rect 9815 22525 9827 22528
rect 9769 22519 9827 22525
rect 9950 22516 9956 22528
rect 10008 22516 10014 22568
rect 10045 22559 10103 22565
rect 10045 22525 10057 22559
rect 10091 22525 10103 22559
rect 10045 22519 10103 22525
rect 10229 22559 10287 22565
rect 10229 22525 10241 22559
rect 10275 22525 10287 22559
rect 10229 22519 10287 22525
rect 10597 22559 10655 22565
rect 10597 22525 10609 22559
rect 10643 22556 10655 22559
rect 10778 22556 10784 22568
rect 10643 22528 10784 22556
rect 10643 22525 10655 22528
rect 10597 22519 10655 22525
rect 6822 22488 6828 22500
rect 6288 22460 6828 22488
rect 6181 22451 6239 22457
rect 6822 22448 6828 22460
rect 6880 22448 6886 22500
rect 8110 22448 8116 22500
rect 8168 22488 8174 22500
rect 10060 22488 10088 22519
rect 8168 22460 10088 22488
rect 8168 22448 8174 22460
rect 4120 22392 4568 22420
rect 4120 22380 4126 22392
rect 4982 22380 4988 22432
rect 5040 22380 5046 22432
rect 5997 22423 6055 22429
rect 5997 22389 6009 22423
rect 6043 22420 6055 22423
rect 6914 22420 6920 22432
rect 6043 22392 6920 22420
rect 6043 22389 6055 22392
rect 5997 22383 6055 22389
rect 6914 22380 6920 22392
rect 6972 22380 6978 22432
rect 8202 22380 8208 22432
rect 8260 22420 8266 22432
rect 8573 22423 8631 22429
rect 8573 22420 8585 22423
rect 8260 22392 8585 22420
rect 8260 22380 8266 22392
rect 8573 22389 8585 22392
rect 8619 22389 8631 22423
rect 8573 22383 8631 22389
rect 9122 22380 9128 22432
rect 9180 22420 9186 22432
rect 9309 22423 9367 22429
rect 9309 22420 9321 22423
rect 9180 22392 9321 22420
rect 9180 22380 9186 22392
rect 9309 22389 9321 22392
rect 9355 22389 9367 22423
rect 9309 22383 9367 22389
rect 9398 22380 9404 22432
rect 9456 22380 9462 22432
rect 9582 22380 9588 22432
rect 9640 22420 9646 22432
rect 10244 22420 10272 22519
rect 10778 22516 10784 22528
rect 10836 22516 10842 22568
rect 10980 22556 11008 22720
rect 12161 22695 12219 22701
rect 12161 22661 12173 22695
rect 12207 22692 12219 22695
rect 12342 22692 12348 22704
rect 12207 22664 12348 22692
rect 12207 22661 12219 22664
rect 12161 22655 12219 22661
rect 12342 22652 12348 22664
rect 12400 22652 12406 22704
rect 11057 22559 11115 22565
rect 11057 22556 11069 22559
rect 10980 22528 11069 22556
rect 11057 22525 11069 22528
rect 11103 22525 11115 22559
rect 11057 22519 11115 22525
rect 11330 22516 11336 22568
rect 11388 22556 11394 22568
rect 12342 22556 12348 22568
rect 11388 22528 12348 22556
rect 11388 22516 11394 22528
rect 12342 22516 12348 22528
rect 12400 22516 12406 22568
rect 11238 22448 11244 22500
rect 11296 22448 11302 22500
rect 11701 22491 11759 22497
rect 11701 22457 11713 22491
rect 11747 22488 11759 22491
rect 11747 22460 12020 22488
rect 11747 22457 11759 22460
rect 11701 22451 11759 22457
rect 9640 22392 10272 22420
rect 9640 22380 9646 22392
rect 11330 22380 11336 22432
rect 11388 22380 11394 22432
rect 11609 22423 11667 22429
rect 11609 22389 11621 22423
rect 11655 22420 11667 22423
rect 11882 22420 11888 22432
rect 11655 22392 11888 22420
rect 11655 22389 11667 22392
rect 11609 22383 11667 22389
rect 11882 22380 11888 22392
rect 11940 22380 11946 22432
rect 11992 22420 12020 22460
rect 12158 22448 12164 22500
rect 12216 22448 12222 22500
rect 12434 22420 12440 22432
rect 11992 22392 12440 22420
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 552 22330 12604 22352
rect 552 22278 4322 22330
rect 4374 22278 4386 22330
rect 4438 22278 4450 22330
rect 4502 22278 4514 22330
rect 4566 22278 4578 22330
rect 4630 22278 10722 22330
rect 10774 22278 10786 22330
rect 10838 22278 10850 22330
rect 10902 22278 10914 22330
rect 10966 22278 10978 22330
rect 11030 22278 12604 22330
rect 552 22256 12604 22278
rect 3142 22176 3148 22228
rect 3200 22216 3206 22228
rect 5261 22219 5319 22225
rect 5261 22216 5273 22219
rect 3200 22188 5273 22216
rect 3200 22176 3206 22188
rect 5261 22185 5273 22188
rect 5307 22216 5319 22219
rect 8662 22216 8668 22228
rect 5307 22188 8668 22216
rect 5307 22185 5319 22188
rect 5261 22179 5319 22185
rect 8662 22176 8668 22188
rect 8720 22176 8726 22228
rect 9858 22176 9864 22228
rect 9916 22176 9922 22228
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 10008 22188 10548 22216
rect 10008 22176 10014 22188
rect 3234 22108 3240 22160
rect 3292 22108 3298 22160
rect 5718 22148 5724 22160
rect 3620 22120 3832 22148
rect 2406 22040 2412 22092
rect 2464 22080 2470 22092
rect 3620 22089 3648 22120
rect 3605 22083 3663 22089
rect 3605 22080 3617 22083
rect 2464 22052 3617 22080
rect 2464 22040 2470 22052
rect 3605 22049 3617 22052
rect 3651 22049 3663 22083
rect 3605 22043 3663 22049
rect 3694 22040 3700 22092
rect 3752 22040 3758 22092
rect 3804 22080 3832 22120
rect 5276 22120 5724 22148
rect 3804 22052 4016 22080
rect 2682 21972 2688 22024
rect 2740 22012 2746 22024
rect 3988 22012 4016 22052
rect 4062 22040 4068 22092
rect 4120 22040 4126 22092
rect 4246 22040 4252 22092
rect 4304 22040 4310 22092
rect 4525 22083 4583 22089
rect 4525 22049 4537 22083
rect 4571 22049 4583 22083
rect 4525 22043 4583 22049
rect 4540 22012 4568 22043
rect 4890 22040 4896 22092
rect 4948 22040 4954 22092
rect 5169 22083 5227 22089
rect 5276 22083 5304 22120
rect 5718 22108 5724 22120
rect 5776 22108 5782 22160
rect 9398 22148 9404 22160
rect 9048 22120 9404 22148
rect 5169 22049 5181 22083
rect 5215 22055 5304 22083
rect 5445 22083 5503 22089
rect 5215 22049 5227 22055
rect 5169 22043 5227 22049
rect 5445 22049 5457 22083
rect 5491 22080 5503 22083
rect 5810 22080 5816 22092
rect 5491 22052 5816 22080
rect 5491 22049 5503 22052
rect 5445 22043 5503 22049
rect 5810 22040 5816 22052
rect 5868 22040 5874 22092
rect 6730 22040 6736 22092
rect 6788 22089 6794 22092
rect 6788 22083 6837 22089
rect 6788 22049 6791 22083
rect 6825 22049 6837 22083
rect 6788 22043 6837 22049
rect 7576 22052 7972 22080
rect 6788 22040 6794 22043
rect 2740 21984 3924 22012
rect 3988 21984 4568 22012
rect 2740 21972 2746 21984
rect 842 21904 848 21956
rect 900 21944 906 21956
rect 1394 21944 1400 21956
rect 900 21916 1400 21944
rect 900 21904 906 21916
rect 1394 21904 1400 21916
rect 1452 21904 1458 21956
rect 2958 21904 2964 21956
rect 3016 21944 3022 21956
rect 3896 21953 3924 21984
rect 5718 21972 5724 22024
rect 5776 21972 5782 22024
rect 5828 22012 5856 22040
rect 7576 22024 7604 22052
rect 6641 22015 6699 22021
rect 6641 22012 6653 22015
rect 5828 21984 6132 22012
rect 3881 21947 3939 21953
rect 3016 21916 3556 21944
rect 3016 21904 3022 21916
rect 658 21836 664 21888
rect 716 21876 722 21888
rect 1029 21879 1087 21885
rect 1029 21876 1041 21879
rect 716 21848 1041 21876
rect 716 21836 722 21848
rect 1029 21845 1041 21848
rect 1075 21876 1087 21879
rect 1118 21876 1124 21888
rect 1075 21848 1124 21876
rect 1075 21845 1087 21848
rect 1029 21839 1087 21845
rect 1118 21836 1124 21848
rect 1176 21836 1182 21888
rect 1670 21836 1676 21888
rect 1728 21876 1734 21888
rect 1949 21879 2007 21885
rect 1949 21876 1961 21879
rect 1728 21848 1961 21876
rect 1728 21836 1734 21848
rect 1949 21845 1961 21848
rect 1995 21876 2007 21879
rect 2222 21876 2228 21888
rect 1995 21848 2228 21876
rect 1995 21845 2007 21848
rect 1949 21839 2007 21845
rect 2222 21836 2228 21848
rect 2280 21836 2286 21888
rect 3234 21836 3240 21888
rect 3292 21876 3298 21888
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 3292 21848 3433 21876
rect 3292 21836 3298 21848
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 3528 21876 3556 21916
rect 3881 21913 3893 21947
rect 3927 21913 3939 21947
rect 5736 21944 5764 21972
rect 5997 21947 6055 21953
rect 5997 21944 6009 21947
rect 5736 21916 6009 21944
rect 3881 21907 3939 21913
rect 5997 21913 6009 21916
rect 6043 21913 6055 21947
rect 5997 21907 6055 21913
rect 4065 21879 4123 21885
rect 4065 21876 4077 21879
rect 3528 21848 4077 21876
rect 3421 21839 3479 21845
rect 4065 21845 4077 21848
rect 4111 21845 4123 21879
rect 4065 21839 4123 21845
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4341 21879 4399 21885
rect 4341 21876 4353 21879
rect 4212 21848 4353 21876
rect 4212 21836 4218 21848
rect 4341 21845 4353 21848
rect 4387 21845 4399 21879
rect 4341 21839 4399 21845
rect 4709 21879 4767 21885
rect 4709 21845 4721 21879
rect 4755 21876 4767 21879
rect 4890 21876 4896 21888
rect 4755 21848 4896 21876
rect 4755 21845 4767 21848
rect 4709 21839 4767 21845
rect 4890 21836 4896 21848
rect 4948 21836 4954 21888
rect 5629 21879 5687 21885
rect 5629 21845 5641 21879
rect 5675 21876 5687 21879
rect 5718 21876 5724 21888
rect 5675 21848 5724 21876
rect 5675 21845 5687 21848
rect 5629 21839 5687 21845
rect 5718 21836 5724 21848
rect 5776 21836 5782 21888
rect 6104 21876 6132 21984
rect 6196 21984 6653 22012
rect 6196 21956 6224 21984
rect 6641 21981 6653 21984
rect 6687 21981 6699 22015
rect 6641 21975 6699 21981
rect 6917 22015 6975 22021
rect 6917 21981 6929 22015
rect 6963 22012 6975 22015
rect 6963 21984 7144 22012
rect 6963 21981 6975 21984
rect 6917 21975 6975 21981
rect 6178 21904 6184 21956
rect 6236 21904 6242 21956
rect 6638 21876 6644 21888
rect 6104 21848 6644 21876
rect 6638 21836 6644 21848
rect 6696 21836 6702 21888
rect 6730 21836 6736 21888
rect 6788 21876 6794 21888
rect 7116 21876 7144 21984
rect 7190 21972 7196 22024
rect 7248 21972 7254 22024
rect 7558 21972 7564 22024
rect 7616 21972 7622 22024
rect 7653 22015 7711 22021
rect 7653 21981 7665 22015
rect 7699 22012 7711 22015
rect 7742 22012 7748 22024
rect 7699 21984 7748 22012
rect 7699 21981 7711 21984
rect 7653 21975 7711 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 21981 7895 22015
rect 7944 22012 7972 22052
rect 8110 22040 8116 22092
rect 8168 22040 8174 22092
rect 8205 22083 8263 22089
rect 8205 22049 8217 22083
rect 8251 22080 8263 22083
rect 8294 22080 8300 22092
rect 8251 22052 8300 22080
rect 8251 22049 8263 22052
rect 8205 22043 8263 22049
rect 8294 22040 8300 22052
rect 8352 22040 8358 22092
rect 8478 22040 8484 22092
rect 8536 22040 8542 22092
rect 8938 22040 8944 22092
rect 8996 22040 9002 22092
rect 9048 22089 9076 22120
rect 9398 22108 9404 22120
rect 9456 22108 9462 22160
rect 9876 22148 9904 22176
rect 10045 22151 10103 22157
rect 10045 22148 10057 22151
rect 9876 22120 10057 22148
rect 10045 22117 10057 22120
rect 10091 22117 10103 22151
rect 10045 22111 10103 22117
rect 10229 22151 10287 22157
rect 10229 22117 10241 22151
rect 10275 22148 10287 22151
rect 10410 22148 10416 22160
rect 10275 22120 10416 22148
rect 10275 22117 10287 22120
rect 10229 22111 10287 22117
rect 10410 22108 10416 22120
rect 10468 22108 10474 22160
rect 10520 22148 10548 22188
rect 10594 22176 10600 22228
rect 10652 22216 10658 22228
rect 10781 22219 10839 22225
rect 10781 22216 10793 22219
rect 10652 22188 10793 22216
rect 10652 22176 10658 22188
rect 10781 22185 10793 22188
rect 10827 22216 10839 22219
rect 11333 22219 11391 22225
rect 11333 22216 11345 22219
rect 10827 22188 11345 22216
rect 10827 22185 10839 22188
rect 10781 22179 10839 22185
rect 11333 22185 11345 22188
rect 11379 22185 11391 22219
rect 11333 22179 11391 22185
rect 11514 22176 11520 22228
rect 11572 22176 11578 22228
rect 11701 22219 11759 22225
rect 11701 22185 11713 22219
rect 11747 22216 11759 22219
rect 11882 22216 11888 22228
rect 11747 22188 11888 22216
rect 11747 22185 11759 22188
rect 11701 22179 11759 22185
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 12434 22216 12440 22228
rect 11992 22188 12440 22216
rect 11992 22148 12020 22188
rect 12434 22176 12440 22188
rect 12492 22176 12498 22228
rect 12158 22148 12164 22160
rect 10520 22120 10732 22148
rect 10704 22092 10732 22120
rect 11713 22120 12020 22148
rect 12084 22120 12164 22148
rect 9033 22083 9091 22089
rect 9033 22049 9045 22083
rect 9079 22049 9091 22083
rect 9033 22043 9091 22049
rect 9122 22038 9128 22090
rect 9180 22089 9186 22090
rect 9180 22043 9188 22089
rect 9309 22083 9367 22089
rect 9309 22080 9321 22083
rect 9232 22052 9321 22080
rect 9180 22038 9186 22043
rect 9232 22024 9260 22052
rect 9309 22049 9321 22052
rect 9355 22049 9367 22083
rect 9309 22043 9367 22049
rect 9860 22083 9918 22089
rect 9860 22049 9872 22083
rect 9906 22049 9918 22083
rect 9860 22043 9918 22049
rect 8389 22015 8447 22021
rect 8389 22012 8401 22015
rect 7944 21984 8401 22012
rect 7837 21975 7895 21981
rect 8389 21981 8401 21984
rect 8435 21981 8447 22015
rect 8389 21975 8447 21981
rect 7466 21904 7472 21956
rect 7524 21944 7530 21956
rect 7852 21944 7880 21975
rect 9214 21972 9220 22024
rect 9272 21972 9278 22024
rect 9876 22012 9904 22043
rect 9950 22040 9956 22092
rect 10008 22040 10014 22092
rect 10321 22083 10379 22089
rect 10321 22049 10333 22083
rect 10367 22080 10379 22083
rect 10367 22052 10456 22080
rect 10367 22049 10379 22052
rect 10321 22043 10379 22049
rect 9876 21984 10364 22012
rect 7524 21916 7880 21944
rect 7524 21904 7530 21916
rect 6788 21848 7144 21876
rect 6788 21836 6794 21848
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 7929 21879 7987 21885
rect 7929 21876 7941 21879
rect 7432 21848 7941 21876
rect 7432 21836 7438 21848
rect 7929 21845 7941 21848
rect 7975 21845 7987 21879
rect 7929 21839 7987 21845
rect 8110 21836 8116 21888
rect 8168 21876 8174 21888
rect 8665 21879 8723 21885
rect 8665 21876 8677 21879
rect 8168 21848 8677 21876
rect 8168 21836 8174 21848
rect 8665 21845 8677 21848
rect 8711 21845 8723 21879
rect 8665 21839 8723 21845
rect 9769 21879 9827 21885
rect 9769 21845 9781 21879
rect 9815 21876 9827 21879
rect 10042 21876 10048 21888
rect 9815 21848 10048 21876
rect 9815 21845 9827 21848
rect 9769 21839 9827 21845
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10336 21885 10364 21984
rect 10428 21944 10456 22052
rect 10502 22040 10508 22092
rect 10560 22040 10566 22092
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22049 10655 22083
rect 10597 22043 10655 22049
rect 10612 22012 10640 22043
rect 10686 22040 10692 22092
rect 10744 22080 10750 22092
rect 11149 22083 11207 22089
rect 11149 22080 11161 22083
rect 10744 22052 11161 22080
rect 10744 22040 10750 22052
rect 11149 22049 11161 22052
rect 11195 22049 11207 22083
rect 11149 22043 11207 22049
rect 11422 22040 11428 22092
rect 11480 22040 11486 22092
rect 11713 22089 11741 22120
rect 12084 22089 12112 22120
rect 12158 22108 12164 22120
rect 12216 22108 12222 22160
rect 11698 22083 11756 22089
rect 11698 22049 11710 22083
rect 11744 22049 11756 22083
rect 11698 22043 11756 22049
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 12115 22052 12149 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 11330 22012 11336 22024
rect 10612 21984 11336 22012
rect 11330 21972 11336 21984
rect 11388 21972 11394 22024
rect 12161 22015 12219 22021
rect 12161 21981 12173 22015
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 10594 21944 10600 21956
rect 10428 21916 10600 21944
rect 10594 21904 10600 21916
rect 10652 21944 10658 21956
rect 11146 21944 11152 21956
rect 10652 21916 11152 21944
rect 10652 21904 10658 21916
rect 11146 21904 11152 21916
rect 11204 21904 11210 21956
rect 11698 21904 11704 21956
rect 11756 21944 11762 21956
rect 12176 21944 12204 21975
rect 11756 21916 12204 21944
rect 11756 21904 11762 21916
rect 10321 21879 10379 21885
rect 10321 21845 10333 21879
rect 10367 21876 10379 21879
rect 10502 21876 10508 21888
rect 10367 21848 10508 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10962 21836 10968 21888
rect 11020 21836 11026 21888
rect 552 21786 12604 21808
rect 552 21734 3662 21786
rect 3714 21734 3726 21786
rect 3778 21734 3790 21786
rect 3842 21734 3854 21786
rect 3906 21734 3918 21786
rect 3970 21734 10062 21786
rect 10114 21734 10126 21786
rect 10178 21734 10190 21786
rect 10242 21734 10254 21786
rect 10306 21734 10318 21786
rect 10370 21734 12604 21786
rect 552 21712 12604 21734
rect 1486 21632 1492 21684
rect 1544 21672 1550 21684
rect 1544 21644 3372 21672
rect 1544 21632 1550 21644
rect 2774 21564 2780 21616
rect 2832 21604 2838 21616
rect 3344 21604 3372 21644
rect 3418 21632 3424 21684
rect 3476 21672 3482 21684
rect 3881 21675 3939 21681
rect 3881 21672 3893 21675
rect 3476 21644 3893 21672
rect 3476 21632 3482 21644
rect 3881 21641 3893 21644
rect 3927 21641 3939 21675
rect 3881 21635 3939 21641
rect 4433 21675 4491 21681
rect 4433 21641 4445 21675
rect 4479 21672 4491 21675
rect 4479 21644 5212 21672
rect 4479 21641 4491 21644
rect 4433 21635 4491 21641
rect 4154 21604 4160 21616
rect 2832 21576 3280 21604
rect 3344 21576 4160 21604
rect 2832 21564 2838 21576
rect 1210 21496 1216 21548
rect 1268 21536 1274 21548
rect 2869 21539 2927 21545
rect 1268 21508 2820 21536
rect 1268 21496 1274 21508
rect 1302 21428 1308 21480
rect 1360 21468 1366 21480
rect 1397 21471 1455 21477
rect 1397 21468 1409 21471
rect 1360 21440 1409 21468
rect 1360 21428 1366 21440
rect 1397 21437 1409 21440
rect 1443 21437 1455 21471
rect 1397 21431 1455 21437
rect 2133 21471 2191 21477
rect 2133 21437 2145 21471
rect 2179 21468 2191 21471
rect 2222 21468 2228 21480
rect 2179 21440 2228 21468
rect 2179 21437 2191 21440
rect 2133 21431 2191 21437
rect 2222 21428 2228 21440
rect 2280 21428 2286 21480
rect 2498 21428 2504 21480
rect 2556 21468 2562 21480
rect 2593 21471 2651 21477
rect 2593 21468 2605 21471
rect 2556 21440 2605 21468
rect 2556 21428 2562 21440
rect 2593 21437 2605 21440
rect 2639 21437 2651 21471
rect 2792 21468 2820 21508
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 3252 21536 3280 21576
rect 4154 21564 4160 21576
rect 4212 21564 4218 21616
rect 4264 21576 4660 21604
rect 3329 21539 3387 21545
rect 3329 21536 3341 21539
rect 3252 21508 3341 21536
rect 3329 21505 3341 21508
rect 3375 21505 3387 21539
rect 3329 21499 3387 21505
rect 3510 21496 3516 21548
rect 3568 21536 3574 21548
rect 3620 21536 3923 21544
rect 4264 21536 4292 21576
rect 3568 21516 4292 21536
rect 3568 21508 3648 21516
rect 3895 21508 4292 21516
rect 4632 21536 4660 21576
rect 4709 21539 4767 21545
rect 4709 21536 4721 21539
rect 4632 21508 4721 21536
rect 3568 21496 3574 21508
rect 4709 21505 4721 21508
rect 4755 21505 4767 21539
rect 5184 21536 5212 21644
rect 5258 21632 5264 21684
rect 5316 21672 5322 21684
rect 5537 21675 5595 21681
rect 5537 21672 5549 21675
rect 5316 21644 5549 21672
rect 5316 21632 5322 21644
rect 5537 21641 5549 21644
rect 5583 21641 5595 21675
rect 5537 21635 5595 21641
rect 5810 21632 5816 21684
rect 5868 21632 5874 21684
rect 7193 21675 7251 21681
rect 7193 21641 7205 21675
rect 7239 21672 7251 21675
rect 8202 21672 8208 21684
rect 7239 21644 8208 21672
rect 7239 21641 7251 21644
rect 7193 21635 7251 21641
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 8386 21632 8392 21684
rect 8444 21632 8450 21684
rect 10594 21672 10600 21684
rect 9876 21644 10600 21672
rect 5721 21607 5779 21613
rect 5721 21573 5733 21607
rect 5767 21573 5779 21607
rect 5721 21567 5779 21573
rect 5626 21536 5632 21548
rect 5184 21508 5632 21536
rect 4709 21499 4767 21505
rect 5626 21496 5632 21508
rect 5684 21496 5690 21548
rect 5736 21536 5764 21567
rect 6546 21564 6552 21616
rect 6604 21564 6610 21616
rect 6641 21607 6699 21613
rect 6641 21573 6653 21607
rect 6687 21604 6699 21607
rect 7006 21604 7012 21616
rect 6687 21576 7012 21604
rect 6687 21573 6699 21576
rect 6641 21567 6699 21573
rect 7006 21564 7012 21576
rect 7064 21564 7070 21616
rect 7098 21564 7104 21616
rect 7156 21604 7162 21616
rect 7285 21607 7343 21613
rect 7285 21604 7297 21607
rect 7156 21576 7297 21604
rect 7156 21564 7162 21576
rect 7285 21573 7297 21576
rect 7331 21573 7343 21607
rect 9582 21604 9588 21616
rect 7285 21567 7343 21573
rect 7852 21576 9588 21604
rect 5736 21508 6132 21536
rect 3602 21468 3608 21480
rect 2792 21440 3608 21468
rect 2593 21431 2651 21437
rect 3602 21428 3608 21440
rect 3660 21428 3666 21480
rect 3786 21428 3792 21480
rect 3844 21428 3850 21480
rect 3970 21428 3976 21480
rect 4028 21428 4034 21480
rect 4246 21428 4252 21480
rect 4304 21428 4310 21480
rect 4338 21428 4344 21480
rect 4396 21468 4402 21480
rect 4525 21471 4583 21477
rect 4525 21470 4537 21471
rect 4448 21468 4537 21470
rect 4396 21442 4537 21468
rect 4396 21440 4476 21442
rect 4396 21428 4402 21440
rect 4525 21437 4537 21442
rect 4571 21437 4583 21471
rect 4525 21431 4583 21437
rect 4623 21471 4681 21477
rect 4623 21437 4635 21471
rect 4669 21470 4681 21471
rect 4801 21471 4859 21477
rect 4669 21442 4752 21470
rect 4669 21437 4681 21442
rect 4623 21431 4681 21437
rect 1121 21403 1179 21409
rect 1121 21369 1133 21403
rect 1167 21369 1179 21403
rect 1121 21363 1179 21369
rect 1136 21332 1164 21363
rect 3878 21360 3884 21412
rect 3936 21400 3942 21412
rect 4065 21403 4123 21409
rect 4065 21400 4077 21403
rect 3936 21372 4077 21400
rect 3936 21360 3942 21372
rect 4065 21369 4077 21372
rect 4111 21369 4123 21403
rect 4065 21363 4123 21369
rect 1394 21332 1400 21344
rect 1136 21304 1400 21332
rect 1394 21292 1400 21304
rect 1452 21292 1458 21344
rect 2314 21292 2320 21344
rect 2372 21332 2378 21344
rect 2409 21335 2467 21341
rect 2409 21332 2421 21335
rect 2372 21304 2421 21332
rect 2372 21292 2378 21304
rect 2409 21301 2421 21304
rect 2455 21301 2467 21335
rect 2409 21295 2467 21301
rect 2958 21292 2964 21344
rect 3016 21332 3022 21344
rect 4724 21332 4752 21442
rect 4801 21437 4813 21471
rect 4847 21468 4859 21471
rect 4890 21468 4896 21480
rect 4847 21440 4896 21468
rect 4847 21437 4859 21440
rect 4801 21431 4859 21437
rect 4890 21428 4896 21440
rect 4948 21428 4954 21480
rect 5718 21428 5724 21480
rect 5776 21468 5782 21480
rect 6104 21477 6132 21508
rect 6822 21496 6828 21548
rect 6880 21536 6886 21548
rect 6880 21508 7236 21536
rect 6880 21496 6886 21508
rect 5813 21471 5871 21477
rect 5813 21468 5825 21471
rect 5776 21440 5825 21468
rect 5776 21428 5782 21440
rect 5813 21437 5825 21440
rect 5859 21437 5871 21471
rect 5813 21431 5871 21437
rect 6089 21471 6147 21477
rect 6089 21437 6101 21471
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6457 21471 6515 21477
rect 6457 21437 6469 21471
rect 6503 21468 6515 21471
rect 6638 21468 6644 21480
rect 6503 21440 6644 21468
rect 6503 21437 6515 21440
rect 6457 21431 6515 21437
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 6733 21471 6791 21477
rect 6733 21437 6745 21471
rect 6779 21468 6791 21471
rect 6914 21468 6920 21480
rect 6779 21440 6920 21468
rect 6779 21437 6791 21440
rect 6733 21431 6791 21437
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 7101 21471 7159 21477
rect 7101 21437 7113 21471
rect 7147 21437 7159 21471
rect 7208 21468 7236 21508
rect 7374 21496 7380 21548
rect 7432 21496 7438 21548
rect 7852 21477 7880 21576
rect 9582 21564 9588 21576
rect 9640 21564 9646 21616
rect 7926 21496 7932 21548
rect 7984 21496 7990 21548
rect 8205 21539 8263 21545
rect 8205 21505 8217 21539
rect 8251 21536 8263 21539
rect 8754 21536 8760 21548
rect 8251 21508 8760 21536
rect 8251 21505 8263 21508
rect 8205 21499 8263 21505
rect 8754 21496 8760 21508
rect 8812 21496 8818 21548
rect 8864 21508 9628 21536
rect 7837 21471 7895 21477
rect 7837 21468 7849 21471
rect 7208 21440 7849 21468
rect 7101 21431 7159 21437
rect 7837 21437 7849 21440
rect 7883 21437 7895 21471
rect 7944 21468 7972 21496
rect 8573 21471 8631 21477
rect 8573 21468 8585 21471
rect 7944 21440 8585 21468
rect 7837 21431 7895 21437
rect 8573 21437 8585 21440
rect 8619 21437 8631 21471
rect 8573 21431 8631 21437
rect 5350 21360 5356 21412
rect 5408 21360 5414 21412
rect 5534 21360 5540 21412
rect 5592 21409 5598 21412
rect 5592 21403 5611 21409
rect 5599 21369 5611 21403
rect 5592 21363 5611 21369
rect 5592 21360 5598 21363
rect 3016 21304 4752 21332
rect 3016 21292 3022 21304
rect 5994 21292 6000 21344
rect 6052 21292 6058 21344
rect 6270 21292 6276 21344
rect 6328 21292 6334 21344
rect 6656 21332 6684 21428
rect 7116 21400 7144 21431
rect 7374 21400 7380 21412
rect 7116 21372 7380 21400
rect 7374 21360 7380 21372
rect 7432 21360 7438 21412
rect 7852 21400 7880 21431
rect 8662 21428 8668 21480
rect 8720 21428 8726 21480
rect 8864 21477 8892 21508
rect 9600 21480 9628 21508
rect 8849 21471 8907 21477
rect 8849 21437 8861 21471
rect 8895 21437 8907 21471
rect 8849 21431 8907 21437
rect 8941 21471 8999 21477
rect 8941 21437 8953 21471
rect 8987 21437 8999 21471
rect 8941 21431 8999 21437
rect 8478 21400 8484 21412
rect 7852 21372 8484 21400
rect 8478 21360 8484 21372
rect 8536 21360 8542 21412
rect 8956 21332 8984 21431
rect 9582 21428 9588 21480
rect 9640 21428 9646 21480
rect 9674 21428 9680 21480
rect 9732 21428 9738 21480
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21468 9827 21471
rect 9876 21468 9904 21644
rect 10594 21632 10600 21644
rect 10652 21632 10658 21684
rect 10870 21632 10876 21684
rect 10928 21672 10934 21684
rect 11514 21672 11520 21684
rect 10928 21644 11520 21672
rect 10928 21632 10934 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 9950 21564 9956 21616
rect 10008 21564 10014 21616
rect 10042 21564 10048 21616
rect 10100 21564 10106 21616
rect 9815 21440 9904 21468
rect 9968 21468 9996 21564
rect 10502 21536 10508 21548
rect 10244 21508 10508 21536
rect 10244 21477 10272 21508
rect 10502 21496 10508 21508
rect 10560 21496 10566 21548
rect 12710 21536 12716 21548
rect 11900 21508 12716 21536
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9968 21440 10057 21468
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 10045 21437 10057 21440
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 10229 21471 10287 21477
rect 10229 21437 10241 21471
rect 10275 21437 10287 21471
rect 10229 21431 10287 21437
rect 10321 21471 10379 21477
rect 10321 21437 10333 21471
rect 10367 21468 10379 21471
rect 10410 21468 10416 21480
rect 10367 21440 10416 21468
rect 10367 21437 10379 21440
rect 10321 21431 10379 21437
rect 10410 21428 10416 21440
rect 10468 21428 10474 21480
rect 11900 21477 11928 21508
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 11885 21471 11943 21477
rect 11885 21437 11897 21471
rect 11931 21437 11943 21471
rect 11885 21431 11943 21437
rect 12069 21471 12127 21477
rect 12069 21437 12081 21471
rect 12115 21468 12127 21471
rect 12342 21468 12348 21480
rect 12115 21440 12348 21468
rect 12115 21437 12127 21440
rect 12069 21431 12127 21437
rect 9858 21360 9864 21412
rect 9916 21400 9922 21412
rect 9953 21403 10011 21409
rect 9953 21400 9965 21403
rect 9916 21372 9965 21400
rect 9916 21360 9922 21372
rect 9953 21369 9965 21372
rect 9999 21369 10011 21403
rect 9953 21363 10011 21369
rect 10502 21360 10508 21412
rect 10560 21400 10566 21412
rect 12084 21400 12112 21431
rect 12342 21428 12348 21440
rect 12400 21428 12406 21480
rect 10560 21372 12112 21400
rect 10560 21360 10566 21372
rect 6656 21304 8984 21332
rect 9030 21292 9036 21344
rect 9088 21332 9094 21344
rect 10962 21332 10968 21344
rect 9088 21304 10968 21332
rect 9088 21292 9094 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11698 21292 11704 21344
rect 11756 21292 11762 21344
rect 552 21242 12604 21264
rect 552 21190 4322 21242
rect 4374 21190 4386 21242
rect 4438 21190 4450 21242
rect 4502 21190 4514 21242
rect 4566 21190 4578 21242
rect 4630 21190 10722 21242
rect 10774 21190 10786 21242
rect 10838 21190 10850 21242
rect 10902 21190 10914 21242
rect 10966 21190 10978 21242
rect 11030 21190 12604 21242
rect 552 21168 12604 21190
rect 2406 21088 2412 21140
rect 2464 21088 2470 21140
rect 2961 21131 3019 21137
rect 2961 21097 2973 21131
rect 3007 21128 3019 21131
rect 3050 21128 3056 21140
rect 3007 21100 3056 21128
rect 3007 21097 3019 21100
rect 2961 21091 3019 21097
rect 3050 21088 3056 21100
rect 3108 21088 3114 21140
rect 3694 21088 3700 21140
rect 3752 21128 3758 21140
rect 4890 21128 4896 21140
rect 3752 21100 4896 21128
rect 3752 21088 3758 21100
rect 4890 21088 4896 21100
rect 4948 21088 4954 21140
rect 4982 21088 4988 21140
rect 5040 21128 5046 21140
rect 5445 21131 5503 21137
rect 5445 21128 5457 21131
rect 5040 21100 5457 21128
rect 5040 21088 5046 21100
rect 5445 21097 5457 21100
rect 5491 21097 5503 21131
rect 5445 21091 5503 21097
rect 6730 21088 6736 21140
rect 6788 21128 6794 21140
rect 7190 21128 7196 21140
rect 6788 21100 7196 21128
rect 6788 21088 6794 21100
rect 7190 21088 7196 21100
rect 7248 21088 7254 21140
rect 7745 21131 7803 21137
rect 7745 21128 7757 21131
rect 7668 21100 7757 21128
rect 3786 21060 3792 21072
rect 2792 21032 3792 21060
rect 1486 20952 1492 21004
rect 1544 20992 1550 21004
rect 1958 20995 2016 21001
rect 1958 20992 1970 20995
rect 1544 20964 1970 20992
rect 1544 20952 1550 20964
rect 1958 20961 1970 20964
rect 2004 20961 2016 20995
rect 1958 20955 2016 20961
rect 2314 20952 2320 21004
rect 2372 20992 2378 21004
rect 2792 21001 2820 21032
rect 3786 21020 3792 21032
rect 3844 21020 3850 21072
rect 6270 21060 6276 21072
rect 4448 21032 6276 21060
rect 2593 20995 2651 21001
rect 2593 20992 2605 20995
rect 2372 20964 2605 20992
rect 2372 20952 2378 20964
rect 2593 20961 2605 20964
rect 2639 20961 2651 20995
rect 2593 20955 2651 20961
rect 2777 20995 2835 21001
rect 2777 20961 2789 20995
rect 2823 20961 2835 20995
rect 2777 20955 2835 20961
rect 3142 20952 3148 21004
rect 3200 20952 3206 21004
rect 3329 20995 3387 21001
rect 3329 20961 3341 20995
rect 3375 20992 3387 20995
rect 3510 20992 3516 21004
rect 3375 20964 3516 20992
rect 3375 20961 3387 20964
rect 3329 20955 3387 20961
rect 3510 20952 3516 20964
rect 3568 20952 3574 21004
rect 3602 20952 3608 21004
rect 3660 20992 3666 21004
rect 3697 20995 3755 21001
rect 3697 20992 3709 20995
rect 3660 20964 3709 20992
rect 3660 20952 3666 20964
rect 3697 20961 3709 20964
rect 3743 20961 3755 20995
rect 3697 20955 3755 20961
rect 3881 20995 3939 21001
rect 3881 20961 3893 20995
rect 3927 20992 3939 20995
rect 3927 20964 4200 20992
rect 3927 20961 3939 20964
rect 3881 20955 3939 20961
rect 2222 20884 2228 20936
rect 2280 20884 2286 20936
rect 2881 20927 2939 20933
rect 2522 20896 2820 20924
rect 2522 20800 2550 20896
rect 2792 20856 2820 20896
rect 2881 20893 2893 20927
rect 2927 20924 2939 20927
rect 3050 20924 3056 20936
rect 2927 20896 3056 20924
rect 2927 20893 2939 20896
rect 2881 20887 2939 20893
rect 3050 20884 3056 20896
rect 3108 20884 3114 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20924 3479 20927
rect 3786 20924 3792 20936
rect 3467 20896 3792 20924
rect 3467 20893 3479 20896
rect 3421 20887 3479 20893
rect 3786 20884 3792 20896
rect 3844 20884 3850 20936
rect 4065 20859 4123 20865
rect 4065 20856 4077 20859
rect 2792 20828 4077 20856
rect 4065 20825 4077 20828
rect 4111 20825 4123 20859
rect 4172 20856 4200 20964
rect 4246 20952 4252 21004
rect 4304 20952 4310 21004
rect 4448 21001 4476 21032
rect 6270 21020 6276 21032
rect 6328 21020 6334 21072
rect 7668 21060 7696 21100
rect 7745 21097 7757 21100
rect 7791 21097 7803 21131
rect 7745 21091 7803 21097
rect 8938 21088 8944 21140
rect 8996 21128 9002 21140
rect 9950 21128 9956 21140
rect 8996 21100 9956 21128
rect 8996 21088 9002 21100
rect 9950 21088 9956 21100
rect 10008 21088 10014 21140
rect 11517 21131 11575 21137
rect 11517 21097 11529 21131
rect 11563 21097 11575 21131
rect 11517 21091 11575 21097
rect 7208 21032 7696 21060
rect 7208 21004 7236 21032
rect 9766 21020 9772 21072
rect 9824 21060 9830 21072
rect 10042 21060 10048 21072
rect 9824 21032 10048 21060
rect 9824 21020 9830 21032
rect 10042 21020 10048 21032
rect 10100 21020 10106 21072
rect 11532 21060 11560 21091
rect 11348 21032 11560 21060
rect 11348 21004 11376 21032
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 4614 20952 4620 21004
rect 4672 20952 4678 21004
rect 4801 20995 4859 21001
rect 4801 20961 4813 20995
rect 4847 20992 4859 20995
rect 4890 20992 4896 21004
rect 4847 20964 4896 20992
rect 4847 20961 4859 20964
rect 4801 20955 4859 20961
rect 4890 20952 4896 20964
rect 4948 20952 4954 21004
rect 5261 20995 5319 21001
rect 5261 20961 5273 20995
rect 5307 20992 5319 20995
rect 5537 20995 5595 21001
rect 5307 20964 5396 20992
rect 5307 20961 5319 20964
rect 5261 20955 5319 20961
rect 5368 20936 5396 20964
rect 5537 20961 5549 20995
rect 5583 20961 5595 20995
rect 5537 20955 5595 20961
rect 4522 20884 4528 20936
rect 4580 20884 4586 20936
rect 4709 20927 4767 20933
rect 4709 20893 4721 20927
rect 4755 20924 4767 20927
rect 4982 20924 4988 20936
rect 4755 20896 4988 20924
rect 4755 20893 4767 20896
rect 4709 20887 4767 20893
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 5350 20884 5356 20936
rect 5408 20884 5414 20936
rect 5552 20924 5580 20955
rect 5810 20952 5816 21004
rect 5868 20952 5874 21004
rect 6638 20952 6644 21004
rect 6696 20992 6702 21004
rect 6733 20995 6791 21001
rect 6733 20992 6745 20995
rect 6696 20964 6745 20992
rect 6696 20952 6702 20964
rect 6733 20961 6745 20964
rect 6779 20961 6791 20995
rect 6733 20955 6791 20961
rect 6917 20995 6975 21001
rect 6917 20961 6929 20995
rect 6963 20992 6975 20995
rect 7190 20992 7196 21004
rect 6963 20964 7196 20992
rect 6963 20961 6975 20964
rect 6917 20955 6975 20961
rect 7190 20952 7196 20964
rect 7248 20952 7254 21004
rect 7374 20952 7380 21004
rect 7432 20952 7438 21004
rect 7466 20952 7472 21004
rect 7524 20992 7530 21004
rect 8386 20992 8392 21004
rect 7524 20964 8392 20992
rect 7524 20952 7530 20964
rect 8386 20952 8392 20964
rect 8444 20992 8450 21004
rect 10502 20992 10508 21004
rect 8444 20964 10508 20992
rect 8444 20952 8450 20964
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 11057 20995 11115 21001
rect 11057 20961 11069 20995
rect 11103 20992 11115 20995
rect 11146 20992 11152 21004
rect 11103 20964 11152 20992
rect 11103 20961 11115 20964
rect 11057 20955 11115 20961
rect 11146 20952 11152 20964
rect 11204 20952 11210 21004
rect 11241 20995 11299 21001
rect 11241 20961 11253 20995
rect 11287 20961 11299 20995
rect 11241 20955 11299 20961
rect 6270 20924 6276 20936
rect 5552 20896 6276 20924
rect 6270 20884 6276 20896
rect 6328 20924 6334 20936
rect 6822 20924 6828 20936
rect 6328 20896 6828 20924
rect 6328 20884 6334 20896
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 7098 20884 7104 20936
rect 7156 20884 7162 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 7650 20924 7656 20936
rect 7331 20896 7656 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 7742 20884 7748 20936
rect 7800 20884 7806 20936
rect 5368 20856 5396 20884
rect 5997 20859 6055 20865
rect 5997 20856 6009 20859
rect 4172 20828 5212 20856
rect 5368 20828 6009 20856
rect 4065 20819 4123 20825
rect 845 20791 903 20797
rect 845 20757 857 20791
rect 891 20788 903 20791
rect 1210 20788 1216 20800
rect 891 20760 1216 20788
rect 891 20757 903 20760
rect 845 20751 903 20757
rect 1210 20748 1216 20760
rect 1268 20748 1274 20800
rect 2498 20748 2504 20800
rect 2556 20748 2562 20800
rect 3510 20748 3516 20800
rect 3568 20748 3574 20800
rect 4246 20748 4252 20800
rect 4304 20788 4310 20800
rect 5077 20791 5135 20797
rect 5077 20788 5089 20791
rect 4304 20760 5089 20788
rect 4304 20748 4310 20760
rect 5077 20757 5089 20760
rect 5123 20757 5135 20791
rect 5184 20788 5212 20828
rect 5997 20825 6009 20828
rect 6043 20825 6055 20859
rect 5997 20819 6055 20825
rect 7193 20859 7251 20865
rect 7193 20825 7205 20859
rect 7239 20856 7251 20859
rect 8386 20856 8392 20868
rect 7239 20828 8392 20856
rect 7239 20825 7251 20828
rect 7193 20819 7251 20825
rect 8386 20816 8392 20828
rect 8444 20816 8450 20868
rect 11256 20856 11284 20955
rect 11330 20952 11336 21004
rect 11388 20952 11394 21004
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20992 11483 20995
rect 11514 20992 11520 21004
rect 11471 20964 11520 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 11606 20952 11612 21004
rect 11664 20992 11670 21004
rect 12066 20992 12072 21004
rect 11664 20964 12072 20992
rect 11664 20952 11670 20964
rect 12066 20952 12072 20964
rect 12124 20952 12130 21004
rect 11422 20856 11428 20868
rect 11256 20828 11428 20856
rect 11422 20816 11428 20828
rect 11480 20816 11486 20868
rect 6362 20788 6368 20800
rect 5184 20760 6368 20788
rect 5077 20751 5135 20757
rect 6362 20748 6368 20760
rect 6420 20748 6426 20800
rect 6914 20748 6920 20800
rect 6972 20748 6978 20800
rect 7561 20791 7619 20797
rect 7561 20757 7573 20791
rect 7607 20788 7619 20791
rect 8202 20788 8208 20800
rect 7607 20760 8208 20788
rect 7607 20757 7619 20760
rect 7561 20751 7619 20757
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 11054 20748 11060 20800
rect 11112 20788 11118 20800
rect 11149 20791 11207 20797
rect 11149 20788 11161 20791
rect 11112 20760 11161 20788
rect 11112 20748 11118 20760
rect 11149 20757 11161 20760
rect 11195 20757 11207 20791
rect 11149 20751 11207 20757
rect 552 20698 12604 20720
rect 552 20646 3662 20698
rect 3714 20646 3726 20698
rect 3778 20646 3790 20698
rect 3842 20646 3854 20698
rect 3906 20646 3918 20698
rect 3970 20646 10062 20698
rect 10114 20646 10126 20698
rect 10178 20646 10190 20698
rect 10242 20646 10254 20698
rect 10306 20646 10318 20698
rect 10370 20646 12604 20698
rect 552 20624 12604 20646
rect 658 20544 664 20596
rect 716 20584 722 20596
rect 3694 20584 3700 20596
rect 716 20556 3700 20584
rect 716 20544 722 20556
rect 3694 20544 3700 20556
rect 3752 20544 3758 20596
rect 3786 20544 3792 20596
rect 3844 20584 3850 20596
rect 4614 20584 4620 20596
rect 3844 20556 4620 20584
rect 3844 20544 3850 20556
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 5626 20544 5632 20596
rect 5684 20544 5690 20596
rect 5718 20544 5724 20596
rect 5776 20584 5782 20596
rect 6638 20584 6644 20596
rect 5776 20556 6644 20584
rect 5776 20544 5782 20556
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 7190 20544 7196 20596
rect 7248 20584 7254 20596
rect 7558 20584 7564 20596
rect 7248 20556 7564 20584
rect 7248 20544 7254 20556
rect 7558 20544 7564 20556
rect 7616 20544 7622 20596
rect 7653 20587 7711 20593
rect 7653 20553 7665 20587
rect 7699 20584 7711 20587
rect 7742 20584 7748 20596
rect 7699 20556 7748 20584
rect 7699 20553 7711 20556
rect 7653 20547 7711 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 7926 20544 7932 20596
rect 7984 20544 7990 20596
rect 8754 20544 8760 20596
rect 8812 20544 8818 20596
rect 9490 20584 9496 20596
rect 9232 20556 9496 20584
rect 14 20476 20 20528
rect 72 20516 78 20528
rect 72 20488 2176 20516
rect 72 20476 78 20488
rect 750 20408 756 20460
rect 808 20448 814 20460
rect 845 20451 903 20457
rect 845 20448 857 20451
rect 808 20420 857 20448
rect 808 20408 814 20420
rect 845 20417 857 20420
rect 891 20417 903 20451
rect 845 20411 903 20417
rect 1210 20408 1216 20460
rect 1268 20448 1274 20460
rect 1581 20451 1639 20457
rect 1581 20448 1593 20451
rect 1268 20420 1593 20448
rect 1268 20408 1274 20420
rect 1581 20417 1593 20420
rect 1627 20417 1639 20451
rect 2148 20448 2176 20488
rect 2682 20476 2688 20528
rect 2740 20476 2746 20528
rect 3418 20516 3424 20528
rect 3160 20488 3424 20516
rect 2777 20451 2835 20457
rect 2148 20437 2728 20448
rect 2777 20437 2789 20451
rect 2148 20420 2789 20437
rect 1581 20411 1639 20417
rect 2700 20417 2789 20420
rect 2823 20437 2835 20451
rect 3160 20448 3188 20488
rect 3418 20476 3424 20488
rect 3476 20476 3482 20528
rect 3970 20476 3976 20528
rect 4028 20516 4034 20528
rect 4801 20519 4859 20525
rect 4801 20516 4813 20519
rect 4028 20488 4813 20516
rect 4028 20476 4034 20488
rect 4801 20485 4813 20488
rect 4847 20485 4859 20519
rect 4801 20479 4859 20485
rect 2884 20437 3188 20448
rect 2823 20420 3188 20437
rect 2823 20417 2912 20420
rect 2700 20409 2912 20417
rect 3234 20408 3240 20460
rect 3292 20448 3298 20460
rect 3605 20451 3663 20457
rect 3605 20448 3617 20451
rect 3292 20420 3617 20448
rect 3292 20408 3298 20420
rect 3605 20417 3617 20420
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20448 3755 20451
rect 4062 20448 4068 20460
rect 3743 20420 4068 20448
rect 3743 20417 3755 20420
rect 3697 20411 3755 20417
rect 4062 20408 4068 20420
rect 4120 20408 4126 20460
rect 4433 20451 4491 20457
rect 4172 20420 4384 20448
rect 1305 20383 1363 20389
rect 1305 20349 1317 20383
rect 1351 20380 1363 20383
rect 1394 20380 1400 20392
rect 1351 20352 1400 20380
rect 1351 20349 1363 20352
rect 1305 20343 1363 20349
rect 1394 20340 1400 20352
rect 1452 20340 1458 20392
rect 1486 20340 1492 20392
rect 1544 20340 1550 20392
rect 1762 20340 1768 20392
rect 1820 20380 1826 20392
rect 2406 20380 2412 20392
rect 1820 20352 2412 20380
rect 1820 20340 1826 20352
rect 2406 20340 2412 20352
rect 2464 20374 2470 20392
rect 2501 20383 2559 20389
rect 2501 20374 2513 20383
rect 2464 20349 2513 20374
rect 2547 20349 2559 20383
rect 2464 20346 2559 20349
rect 2464 20340 2470 20346
rect 2501 20343 2559 20346
rect 3142 20340 3148 20392
rect 3200 20340 3206 20392
rect 3421 20383 3479 20389
rect 3421 20349 3433 20383
rect 3467 20349 3479 20383
rect 4172 20380 4200 20420
rect 3421 20343 3479 20349
rect 3620 20352 4200 20380
rect 3160 20312 3188 20340
rect 3436 20312 3464 20343
rect 3620 20324 3648 20352
rect 4246 20340 4252 20392
rect 4304 20340 4310 20392
rect 4356 20380 4384 20420
rect 4433 20417 4445 20451
rect 4479 20448 4491 20451
rect 4816 20448 4844 20479
rect 5350 20476 5356 20528
rect 5408 20516 5414 20528
rect 5905 20519 5963 20525
rect 5905 20516 5917 20519
rect 5408 20488 5917 20516
rect 5408 20476 5414 20488
rect 5905 20485 5917 20488
rect 5951 20485 5963 20519
rect 5905 20479 5963 20485
rect 5997 20519 6055 20525
rect 5997 20485 6009 20519
rect 6043 20516 6055 20519
rect 6914 20516 6920 20528
rect 6043 20488 6920 20516
rect 6043 20485 6055 20488
rect 5997 20479 6055 20485
rect 6914 20476 6920 20488
rect 6972 20476 6978 20528
rect 9232 20516 9260 20556
rect 9490 20544 9496 20556
rect 9548 20584 9554 20596
rect 9548 20556 9674 20584
rect 9548 20544 9554 20556
rect 7116 20488 9260 20516
rect 6549 20451 6607 20457
rect 4479 20420 4752 20448
rect 4816 20420 5856 20448
rect 4479 20417 4491 20420
rect 4433 20411 4491 20417
rect 4522 20380 4528 20392
rect 4356 20352 4528 20380
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 4617 20383 4675 20389
rect 4617 20349 4629 20383
rect 4663 20349 4675 20383
rect 4617 20343 4675 20349
rect 2332 20284 3464 20312
rect 1578 20204 1584 20256
rect 1636 20244 1642 20256
rect 2332 20253 2360 20284
rect 3602 20272 3608 20324
rect 3660 20272 3666 20324
rect 3694 20272 3700 20324
rect 3752 20312 3758 20324
rect 4065 20315 4123 20321
rect 4065 20312 4077 20315
rect 3752 20284 4077 20312
rect 3752 20272 3758 20284
rect 4065 20281 4077 20284
rect 4111 20281 4123 20315
rect 4065 20275 4123 20281
rect 4154 20272 4160 20324
rect 4212 20312 4218 20324
rect 4632 20312 4660 20343
rect 4212 20284 4660 20312
rect 4212 20272 4218 20284
rect 2317 20247 2375 20253
rect 2317 20244 2329 20247
rect 1636 20216 2329 20244
rect 1636 20204 1642 20216
rect 2317 20213 2329 20216
rect 2363 20213 2375 20247
rect 2317 20207 2375 20213
rect 3237 20247 3295 20253
rect 3237 20213 3249 20247
rect 3283 20244 3295 20247
rect 3326 20244 3332 20256
rect 3283 20216 3332 20244
rect 3283 20213 3295 20216
rect 3237 20207 3295 20213
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 3970 20204 3976 20256
rect 4028 20244 4034 20256
rect 4614 20244 4620 20256
rect 4028 20216 4620 20244
rect 4028 20204 4034 20216
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 4724 20244 4752 20420
rect 5828 20392 5856 20420
rect 6549 20417 6561 20451
rect 6595 20448 6607 20451
rect 7006 20448 7012 20460
rect 6595 20420 7012 20448
rect 6595 20417 6607 20420
rect 6549 20411 6607 20417
rect 7006 20408 7012 20420
rect 7064 20408 7070 20460
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 6089 20383 6147 20389
rect 6089 20349 6101 20383
rect 6135 20380 6147 20383
rect 6270 20380 6276 20392
rect 6135 20352 6276 20380
rect 6135 20349 6147 20352
rect 6089 20343 6147 20349
rect 6270 20340 6276 20352
rect 6328 20340 6334 20392
rect 6457 20383 6515 20389
rect 6457 20349 6469 20383
rect 6503 20349 6515 20383
rect 6457 20343 6515 20349
rect 5828 20312 5856 20340
rect 6472 20312 6500 20343
rect 6638 20340 6644 20392
rect 6696 20340 6702 20392
rect 6733 20383 6791 20389
rect 6733 20349 6745 20383
rect 6779 20380 6791 20383
rect 6822 20380 6828 20392
rect 6779 20352 6828 20380
rect 6779 20349 6791 20352
rect 6733 20343 6791 20349
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7116 20389 7144 20488
rect 9306 20476 9312 20528
rect 9364 20476 9370 20528
rect 9646 20516 9674 20556
rect 9858 20544 9864 20596
rect 9916 20544 9922 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11241 20587 11299 20593
rect 11241 20584 11253 20587
rect 11204 20556 11253 20584
rect 11204 20544 11210 20556
rect 11241 20553 11253 20556
rect 11287 20553 11299 20587
rect 11241 20547 11299 20553
rect 11701 20519 11759 20525
rect 11701 20516 11713 20519
rect 9646 20488 11713 20516
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20448 7251 20451
rect 7926 20448 7932 20460
rect 7239 20420 7932 20448
rect 7239 20417 7251 20420
rect 7193 20411 7251 20417
rect 7101 20383 7159 20389
rect 7101 20349 7113 20383
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 5828 20284 6500 20312
rect 6914 20272 6920 20324
rect 6972 20312 6978 20324
rect 7208 20312 7236 20411
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 8294 20408 8300 20460
rect 8352 20448 8358 20460
rect 8846 20448 8852 20460
rect 8352 20420 8852 20448
rect 8352 20408 8358 20420
rect 8846 20408 8852 20420
rect 8904 20448 8910 20460
rect 8941 20451 8999 20457
rect 8941 20448 8953 20451
rect 8904 20420 8953 20448
rect 8904 20408 8910 20420
rect 8941 20417 8953 20420
rect 8987 20417 8999 20451
rect 8941 20411 8999 20417
rect 7282 20340 7288 20392
rect 7340 20380 7346 20392
rect 7377 20383 7435 20389
rect 7377 20380 7389 20383
rect 7340 20352 7389 20380
rect 7340 20340 7346 20352
rect 7377 20349 7389 20352
rect 7423 20349 7435 20383
rect 7377 20343 7435 20349
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 6972 20284 7236 20312
rect 6972 20272 6978 20284
rect 6273 20247 6331 20253
rect 6273 20244 6285 20247
rect 4724 20216 6285 20244
rect 6273 20213 6285 20216
rect 6319 20213 6331 20247
rect 6273 20207 6331 20213
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 7484 20244 7512 20343
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 7745 20383 7803 20389
rect 7745 20380 7757 20383
rect 7616 20352 7757 20380
rect 7616 20340 7622 20352
rect 7745 20349 7757 20352
rect 7791 20380 7803 20383
rect 8018 20380 8024 20392
rect 7791 20352 8024 20380
rect 7791 20349 7803 20352
rect 7745 20343 7803 20349
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 8386 20340 8392 20392
rect 8444 20340 8450 20392
rect 8478 20340 8484 20392
rect 8536 20380 8542 20392
rect 8573 20383 8631 20389
rect 8573 20380 8585 20383
rect 8536 20352 8585 20380
rect 8536 20340 8542 20352
rect 8573 20349 8585 20352
rect 8619 20349 8631 20383
rect 8573 20343 8631 20349
rect 8110 20272 8116 20324
rect 8168 20312 8174 20324
rect 8588 20312 8616 20343
rect 8662 20340 8668 20392
rect 8720 20340 8726 20392
rect 8754 20340 8760 20392
rect 8812 20380 8818 20392
rect 9033 20383 9091 20389
rect 9033 20380 9045 20383
rect 8812 20352 9045 20380
rect 8812 20340 8818 20352
rect 9033 20349 9045 20352
rect 9079 20349 9091 20383
rect 9033 20343 9091 20349
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9324 20380 9352 20476
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 10888 20457 10916 20488
rect 11701 20485 11713 20488
rect 11747 20485 11759 20519
rect 11701 20479 11759 20485
rect 10045 20451 10103 20457
rect 10045 20448 10057 20451
rect 9640 20420 10057 20448
rect 9640 20408 9646 20420
rect 10045 20417 10057 20420
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 9498 20383 9556 20389
rect 9498 20380 9510 20383
rect 9180 20352 9225 20380
rect 9324 20352 9510 20380
rect 9180 20340 9186 20352
rect 9498 20349 9510 20352
rect 9544 20349 9556 20383
rect 9498 20343 9556 20349
rect 10137 20383 10195 20389
rect 10137 20349 10149 20383
rect 10183 20380 10195 20383
rect 10502 20380 10508 20392
rect 10183 20352 10508 20380
rect 10183 20349 10195 20352
rect 10137 20343 10195 20349
rect 10502 20340 10508 20352
rect 10560 20340 10566 20392
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11974 20380 11980 20392
rect 11011 20352 11980 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 11974 20340 11980 20352
rect 12032 20380 12038 20392
rect 12342 20380 12348 20392
rect 12032 20352 12348 20380
rect 12032 20340 12038 20352
rect 12342 20340 12348 20352
rect 12400 20340 12406 20392
rect 8168 20284 8616 20312
rect 8168 20272 8174 20284
rect 7248 20216 7512 20244
rect 7248 20204 7254 20216
rect 8478 20204 8484 20256
rect 8536 20204 8542 20256
rect 8588 20244 8616 20284
rect 8941 20315 8999 20321
rect 8941 20281 8953 20315
rect 8987 20312 8999 20315
rect 9309 20315 9367 20321
rect 9309 20312 9321 20315
rect 8987 20284 9321 20312
rect 8987 20281 8999 20284
rect 8941 20275 8999 20281
rect 9309 20281 9321 20284
rect 9355 20281 9367 20315
rect 9309 20275 9367 20281
rect 9398 20272 9404 20324
rect 9456 20312 9462 20324
rect 10410 20312 10416 20324
rect 9456 20284 10416 20312
rect 9456 20272 9462 20284
rect 10410 20272 10416 20284
rect 10468 20272 10474 20324
rect 10686 20272 10692 20324
rect 10744 20312 10750 20324
rect 11517 20315 11575 20321
rect 11517 20312 11529 20315
rect 10744 20284 11529 20312
rect 10744 20272 10750 20284
rect 11517 20281 11529 20284
rect 11563 20281 11575 20315
rect 11517 20275 11575 20281
rect 9214 20244 9220 20256
rect 8588 20216 9220 20244
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9677 20247 9735 20253
rect 9677 20213 9689 20247
rect 9723 20244 9735 20247
rect 9858 20244 9864 20256
rect 9723 20216 9864 20244
rect 9723 20213 9735 20216
rect 9677 20207 9735 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 552 20154 12604 20176
rect 552 20102 4322 20154
rect 4374 20102 4386 20154
rect 4438 20102 4450 20154
rect 4502 20102 4514 20154
rect 4566 20102 4578 20154
rect 4630 20102 10722 20154
rect 10774 20102 10786 20154
rect 10838 20102 10850 20154
rect 10902 20102 10914 20154
rect 10966 20102 10978 20154
rect 11030 20102 12604 20154
rect 552 20080 12604 20102
rect 934 20000 940 20052
rect 992 20000 998 20052
rect 1670 20000 1676 20052
rect 1728 20040 1734 20052
rect 2682 20040 2688 20052
rect 1728 20012 2688 20040
rect 1728 20000 1734 20012
rect 2682 20000 2688 20012
rect 2740 20000 2746 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 2884 20012 3433 20040
rect 2406 19932 2412 19984
rect 2464 19972 2470 19984
rect 2501 19975 2559 19981
rect 2501 19972 2513 19975
rect 2464 19944 2513 19972
rect 2464 19932 2470 19944
rect 2501 19941 2513 19944
rect 2547 19941 2559 19975
rect 2501 19935 2559 19941
rect 1121 19907 1179 19913
rect 1121 19873 1133 19907
rect 1167 19904 1179 19907
rect 1670 19904 1676 19916
rect 1167 19876 1676 19904
rect 1167 19873 1179 19876
rect 1121 19867 1179 19873
rect 1670 19864 1676 19876
rect 1728 19904 1734 19916
rect 2133 19907 2191 19913
rect 2133 19904 2145 19907
rect 1728 19876 2145 19904
rect 1728 19864 1734 19876
rect 2133 19873 2145 19876
rect 2179 19873 2191 19907
rect 2133 19867 2191 19873
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 2884 19904 2912 20012
rect 3421 20009 3433 20012
rect 3467 20040 3479 20043
rect 3510 20040 3516 20052
rect 3467 20012 3516 20040
rect 3467 20009 3479 20012
rect 3421 20003 3479 20009
rect 3510 20000 3516 20012
rect 3568 20040 3574 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 3568 20012 3801 20040
rect 3568 20000 3574 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 3789 20003 3847 20009
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4065 20043 4123 20049
rect 4065 20040 4077 20043
rect 4028 20012 4077 20040
rect 4028 20000 4034 20012
rect 4065 20009 4077 20012
rect 4111 20009 4123 20043
rect 4065 20003 4123 20009
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 5626 20040 5632 20052
rect 4212 20012 4752 20040
rect 4212 20000 4218 20012
rect 4724 19972 4752 20012
rect 5092 20012 5632 20040
rect 5092 19972 5120 20012
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 6362 20040 6368 20052
rect 6104 20012 6368 20040
rect 6104 19972 6132 20012
rect 6362 20000 6368 20012
rect 6420 20040 6426 20052
rect 6917 20043 6975 20049
rect 6420 20012 6714 20040
rect 6420 20000 6426 20012
rect 3252 19944 3648 19972
rect 4724 19944 5120 19972
rect 5568 19944 6132 19972
rect 6181 19975 6239 19981
rect 3252 19913 3280 19944
rect 3620 19916 3648 19944
rect 2823 19876 2912 19904
rect 3237 19907 3295 19913
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 658 19796 664 19848
rect 716 19836 722 19848
rect 1305 19839 1363 19845
rect 1305 19836 1317 19839
rect 716 19808 1317 19836
rect 716 19796 722 19808
rect 1305 19805 1317 19808
rect 1351 19805 1363 19839
rect 1305 19799 1363 19805
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19836 1455 19839
rect 2038 19836 2044 19848
rect 1443 19808 2044 19836
rect 1443 19805 1455 19808
rect 1397 19799 1455 19805
rect 1412 19768 1440 19799
rect 2038 19796 2044 19808
rect 2096 19836 2102 19848
rect 2409 19839 2467 19845
rect 2409 19836 2421 19839
rect 2096 19808 2421 19836
rect 2096 19796 2102 19808
rect 2409 19805 2421 19808
rect 2455 19805 2467 19839
rect 2409 19799 2467 19805
rect 2498 19796 2504 19848
rect 2556 19796 2562 19848
rect 2884 19845 2912 19876
rect 3126 19897 3184 19903
rect 3126 19863 3138 19897
rect 3172 19894 3184 19897
rect 3172 19863 3188 19894
rect 3237 19873 3249 19907
rect 3283 19873 3295 19907
rect 3237 19867 3295 19873
rect 3510 19864 3516 19916
rect 3568 19864 3574 19916
rect 3602 19864 3608 19916
rect 3660 19864 3666 19916
rect 3878 19864 3884 19916
rect 3936 19864 3942 19916
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19904 4031 19907
rect 4062 19904 4068 19916
rect 4019 19876 4068 19904
rect 4019 19873 4031 19876
rect 3973 19867 4031 19873
rect 3126 19857 3188 19863
rect 2869 19839 2927 19845
rect 2869 19805 2881 19839
rect 2915 19805 2927 19839
rect 3160 19836 3188 19857
rect 3988 19836 4016 19867
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 4154 19864 4160 19916
rect 4212 19864 4218 19916
rect 4430 19864 4436 19916
rect 4488 19864 4494 19916
rect 4522 19864 4528 19916
rect 4580 19904 4586 19916
rect 4709 19907 4767 19913
rect 4709 19904 4721 19907
rect 4580 19876 4721 19904
rect 4580 19864 4586 19876
rect 4709 19873 4721 19876
rect 4755 19873 4767 19907
rect 4709 19867 4767 19873
rect 4801 19907 4859 19913
rect 4801 19873 4813 19907
rect 4847 19873 4859 19907
rect 4801 19867 4859 19873
rect 3160 19808 3372 19836
rect 2869 19799 2927 19805
rect 1320 19740 1440 19768
rect 2317 19771 2375 19777
rect 1320 19712 1348 19740
rect 2317 19737 2329 19771
rect 2363 19768 2375 19771
rect 2516 19768 2544 19796
rect 2363 19740 2544 19768
rect 2363 19737 2375 19740
rect 2317 19731 2375 19737
rect 3050 19728 3056 19780
rect 3108 19728 3114 19780
rect 3142 19728 3148 19780
rect 3200 19768 3206 19780
rect 3237 19771 3295 19777
rect 3237 19768 3249 19771
rect 3200 19740 3249 19768
rect 3200 19728 3206 19740
rect 3237 19737 3249 19740
rect 3283 19737 3295 19771
rect 3344 19768 3372 19808
rect 3895 19808 4016 19836
rect 4617 19839 4675 19845
rect 3895 19768 3923 19808
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 4663 19808 4752 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 3344 19740 3923 19768
rect 3237 19731 3295 19737
rect 3970 19728 3976 19780
rect 4028 19768 4034 19780
rect 4028 19740 4660 19768
rect 4028 19728 4034 19740
rect 4632 19712 4660 19740
rect 1302 19660 1308 19712
rect 1360 19660 1366 19712
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 1949 19703 2007 19709
rect 1949 19700 1961 19703
rect 1728 19672 1961 19700
rect 1728 19660 1734 19672
rect 1949 19669 1961 19672
rect 1995 19669 2007 19703
rect 1949 19663 2007 19669
rect 2498 19660 2504 19712
rect 2556 19660 2562 19712
rect 2866 19660 2872 19712
rect 2924 19700 2930 19712
rect 2961 19703 3019 19709
rect 2961 19700 2973 19703
rect 2924 19672 2973 19700
rect 2924 19660 2930 19672
rect 2961 19669 2973 19672
rect 3007 19669 3019 19703
rect 2961 19663 3019 19669
rect 3605 19703 3663 19709
rect 3605 19669 3617 19703
rect 3651 19700 3663 19703
rect 3786 19700 3792 19712
rect 3651 19672 3792 19700
rect 3651 19669 3663 19672
rect 3605 19663 3663 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4154 19660 4160 19712
rect 4212 19700 4218 19712
rect 4249 19703 4307 19709
rect 4249 19700 4261 19703
rect 4212 19672 4261 19700
rect 4212 19660 4218 19672
rect 4249 19669 4261 19672
rect 4295 19669 4307 19703
rect 4249 19663 4307 19669
rect 4614 19660 4620 19712
rect 4672 19660 4678 19712
rect 4724 19700 4752 19808
rect 4816 19828 4844 19867
rect 4890 19864 4896 19916
rect 4948 19904 4954 19916
rect 4985 19907 5043 19913
rect 4985 19904 4997 19907
rect 4948 19876 4997 19904
rect 4948 19864 4954 19876
rect 4985 19873 4997 19876
rect 5031 19873 5043 19907
rect 4985 19867 5043 19873
rect 5353 19907 5411 19913
rect 5353 19873 5365 19907
rect 5399 19904 5411 19907
rect 5442 19904 5448 19916
rect 5399 19876 5448 19904
rect 5399 19873 5411 19876
rect 5353 19867 5411 19873
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 5568 19836 5596 19944
rect 6181 19941 6193 19975
rect 6227 19972 6239 19975
rect 6270 19972 6276 19984
rect 6227 19944 6276 19972
rect 6227 19941 6239 19944
rect 6181 19935 6239 19941
rect 6270 19932 6276 19944
rect 6328 19932 6334 19984
rect 5626 19864 5632 19916
rect 5684 19904 5690 19916
rect 5813 19907 5871 19913
rect 5813 19904 5825 19907
rect 5684 19876 5825 19904
rect 5684 19864 5690 19876
rect 5813 19873 5825 19876
rect 5859 19873 5871 19907
rect 6549 19907 6607 19913
rect 6549 19904 6561 19907
rect 5813 19867 5871 19873
rect 6288 19876 6561 19904
rect 6288 19848 6316 19876
rect 6549 19873 6561 19876
rect 6595 19873 6607 19907
rect 6686 19904 6714 20012
rect 6917 20009 6929 20043
rect 6963 20040 6975 20043
rect 7098 20040 7104 20052
rect 6963 20012 7104 20040
rect 6963 20009 6975 20012
rect 6917 20003 6975 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7466 20000 7472 20052
rect 7524 20000 7530 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 8570 20040 8576 20052
rect 8260 20012 8576 20040
rect 8260 20000 8266 20012
rect 8570 20000 8576 20012
rect 8628 20000 8634 20052
rect 10594 20040 10600 20052
rect 8680 20012 10600 20040
rect 7484 19972 7512 20000
rect 8478 19972 8484 19984
rect 7208 19944 7512 19972
rect 7852 19944 8484 19972
rect 6914 19904 6920 19916
rect 6686 19876 6920 19904
rect 6549 19867 6607 19873
rect 6914 19864 6920 19876
rect 6972 19904 6978 19916
rect 7208 19913 7236 19944
rect 7852 19913 7880 19944
rect 8478 19932 8484 19944
rect 8536 19932 8542 19984
rect 8680 19972 8708 20012
rect 10594 20000 10600 20012
rect 10652 20040 10658 20052
rect 10962 20040 10968 20052
rect 10652 20012 10968 20040
rect 10652 20000 10658 20012
rect 10962 20000 10968 20012
rect 11020 20000 11026 20052
rect 11330 20000 11336 20052
rect 11388 20000 11394 20052
rect 11532 20012 12020 20040
rect 8588 19944 8708 19972
rect 7101 19907 7159 19913
rect 7101 19904 7113 19907
rect 6972 19876 7113 19904
rect 6972 19864 6978 19876
rect 7101 19873 7113 19876
rect 7147 19873 7159 19907
rect 7101 19867 7159 19873
rect 7193 19907 7251 19913
rect 7193 19873 7205 19907
rect 7239 19873 7251 19907
rect 7193 19867 7251 19873
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 7837 19907 7895 19913
rect 7837 19873 7849 19907
rect 7883 19873 7895 19907
rect 7837 19867 7895 19873
rect 5000 19828 5596 19836
rect 4816 19808 5596 19828
rect 4816 19800 5028 19808
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5776 19808 5856 19836
rect 5776 19796 5782 19808
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 4724 19672 5181 19700
rect 5169 19669 5181 19672
rect 5215 19700 5227 19703
rect 5718 19700 5724 19712
rect 5215 19672 5724 19700
rect 5215 19669 5227 19672
rect 5169 19663 5227 19669
rect 5718 19660 5724 19672
rect 5776 19660 5782 19712
rect 5828 19700 5856 19808
rect 6270 19796 6276 19848
rect 6328 19796 6334 19848
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 7377 19839 7435 19845
rect 7377 19836 7389 19839
rect 7340 19808 7389 19836
rect 7340 19796 7346 19808
rect 7377 19805 7389 19808
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 6454 19728 6460 19780
rect 6512 19768 6518 19780
rect 7484 19768 7512 19867
rect 7926 19864 7932 19916
rect 7984 19864 7990 19916
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19873 8079 19907
rect 8021 19867 8079 19873
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19904 8263 19907
rect 8294 19904 8300 19916
rect 8251 19876 8300 19904
rect 8251 19873 8263 19876
rect 8205 19867 8263 19873
rect 8036 19836 8064 19867
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 8588 19836 8616 19944
rect 8846 19932 8852 19984
rect 8904 19972 8910 19984
rect 10689 19975 10747 19981
rect 10689 19972 10701 19975
rect 8904 19944 10088 19972
rect 8904 19932 8910 19944
rect 8665 19907 8723 19913
rect 8665 19873 8677 19907
rect 8711 19904 8723 19907
rect 9122 19904 9128 19916
rect 8711 19876 9128 19904
rect 8711 19873 8723 19876
rect 8665 19867 8723 19873
rect 9122 19864 9128 19876
rect 9180 19904 9186 19916
rect 9180 19876 9260 19904
rect 9180 19864 9186 19876
rect 8036 19808 8616 19836
rect 8754 19796 8760 19848
rect 8812 19796 8818 19848
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19836 8999 19839
rect 9030 19836 9036 19848
rect 8987 19808 9036 19836
rect 8987 19805 8999 19808
rect 8941 19799 8999 19805
rect 9030 19796 9036 19808
rect 9088 19796 9094 19848
rect 9232 19845 9260 19876
rect 9306 19864 9312 19916
rect 9364 19864 9370 19916
rect 10060 19913 10088 19944
rect 10336 19944 10701 19972
rect 10336 19913 10364 19944
rect 10689 19941 10701 19944
rect 10735 19972 10747 19975
rect 10870 19972 10876 19984
rect 10735 19944 10876 19972
rect 10735 19941 10747 19944
rect 10689 19935 10747 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19873 10103 19907
rect 10045 19867 10103 19873
rect 10321 19907 10379 19913
rect 10321 19873 10333 19907
rect 10367 19873 10379 19907
rect 10321 19867 10379 19873
rect 10505 19907 10563 19913
rect 10505 19873 10517 19907
rect 10551 19873 10563 19907
rect 10505 19867 10563 19873
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 9769 19839 9827 19845
rect 9769 19805 9781 19839
rect 9815 19805 9827 19839
rect 10520 19836 10548 19867
rect 10594 19864 10600 19916
rect 10652 19864 10658 19916
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 11054 19904 11060 19916
rect 10827 19876 11060 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 11146 19864 11152 19916
rect 11204 19864 11210 19916
rect 11422 19864 11428 19916
rect 11480 19864 11486 19916
rect 11532 19836 11560 20012
rect 11882 19932 11888 19984
rect 11940 19932 11946 19984
rect 11992 19913 12020 20012
rect 11701 19907 11759 19913
rect 11701 19873 11713 19907
rect 11747 19902 11759 19907
rect 11977 19907 12035 19913
rect 11808 19902 11928 19904
rect 11747 19876 11928 19902
rect 11747 19874 11836 19876
rect 11747 19873 11759 19874
rect 11701 19867 11759 19873
rect 11900 19848 11928 19876
rect 11977 19873 11989 19907
rect 12023 19904 12035 19907
rect 12158 19904 12164 19916
rect 12023 19876 12164 19904
rect 12023 19873 12035 19876
rect 11977 19867 12035 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 10520 19808 11560 19836
rect 9769 19799 9827 19805
rect 7742 19768 7748 19780
rect 6512 19740 7748 19768
rect 6512 19728 6518 19740
rect 7742 19728 7748 19740
rect 7800 19728 7806 19780
rect 8294 19728 8300 19780
rect 8352 19728 8358 19780
rect 8662 19728 8668 19780
rect 8720 19768 8726 19780
rect 9306 19768 9312 19780
rect 8720 19740 9312 19768
rect 8720 19728 8726 19740
rect 9048 19712 9076 19740
rect 9306 19728 9312 19740
rect 9364 19768 9370 19780
rect 9784 19768 9812 19799
rect 11882 19796 11888 19848
rect 11940 19796 11946 19848
rect 9364 19740 9812 19768
rect 9364 19728 9370 19740
rect 10594 19728 10600 19780
rect 10652 19768 10658 19780
rect 11517 19771 11575 19777
rect 11517 19768 11529 19771
rect 10652 19740 11529 19768
rect 10652 19728 10658 19740
rect 11517 19737 11529 19740
rect 11563 19737 11575 19771
rect 11517 19731 11575 19737
rect 6733 19703 6791 19709
rect 6733 19700 6745 19703
rect 5828 19672 6745 19700
rect 6733 19669 6745 19672
rect 6779 19700 6791 19703
rect 6822 19700 6828 19712
rect 6779 19672 6828 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7561 19703 7619 19709
rect 7561 19669 7573 19703
rect 7607 19700 7619 19703
rect 8202 19700 8208 19712
rect 7607 19672 8208 19700
rect 7607 19669 7619 19672
rect 7561 19663 7619 19669
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 9030 19660 9036 19712
rect 9088 19660 9094 19712
rect 9677 19703 9735 19709
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 9861 19703 9919 19709
rect 9861 19700 9873 19703
rect 9723 19672 9873 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 9861 19669 9873 19672
rect 9907 19669 9919 19703
rect 9861 19663 9919 19669
rect 10229 19703 10287 19709
rect 10229 19669 10241 19703
rect 10275 19700 10287 19703
rect 10410 19700 10416 19712
rect 10275 19672 10416 19700
rect 10275 19669 10287 19672
rect 10229 19663 10287 19669
rect 10410 19660 10416 19672
rect 10468 19660 10474 19712
rect 10502 19660 10508 19712
rect 10560 19660 10566 19712
rect 10962 19660 10968 19712
rect 11020 19660 11026 19712
rect 11054 19660 11060 19712
rect 11112 19700 11118 19712
rect 11882 19700 11888 19712
rect 11112 19672 11888 19700
rect 11112 19660 11118 19672
rect 11882 19660 11888 19672
rect 11940 19660 11946 19712
rect 552 19610 12604 19632
rect 552 19558 3662 19610
rect 3714 19558 3726 19610
rect 3778 19558 3790 19610
rect 3842 19558 3854 19610
rect 3906 19558 3918 19610
rect 3970 19558 10062 19610
rect 10114 19558 10126 19610
rect 10178 19558 10190 19610
rect 10242 19558 10254 19610
rect 10306 19558 10318 19610
rect 10370 19558 12604 19610
rect 552 19536 12604 19558
rect 1397 19499 1455 19505
rect 1397 19465 1409 19499
rect 1443 19496 1455 19499
rect 1486 19496 1492 19508
rect 1443 19468 1492 19496
rect 1443 19465 1455 19468
rect 1397 19459 1455 19465
rect 1486 19456 1492 19468
rect 1544 19456 1550 19508
rect 2501 19499 2559 19505
rect 2501 19465 2513 19499
rect 2547 19496 2559 19499
rect 3234 19496 3240 19508
rect 2547 19468 3240 19496
rect 2547 19465 2559 19468
rect 2501 19459 2559 19465
rect 3234 19456 3240 19468
rect 3292 19456 3298 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 5166 19496 5172 19508
rect 4488 19468 5172 19496
rect 4488 19456 4494 19468
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 6638 19456 6644 19508
rect 6696 19496 6702 19508
rect 7469 19499 7527 19505
rect 7469 19496 7481 19499
rect 6696 19468 7481 19496
rect 6696 19456 6702 19468
rect 7469 19465 7481 19468
rect 7515 19465 7527 19499
rect 7469 19459 7527 19465
rect 7745 19499 7803 19505
rect 7745 19465 7757 19499
rect 7791 19496 7803 19499
rect 7926 19496 7932 19508
rect 7791 19468 7932 19496
rect 7791 19465 7803 19468
rect 7745 19459 7803 19465
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 8266 19468 8524 19496
rect 1946 19388 1952 19440
rect 2004 19428 2010 19440
rect 2866 19428 2872 19440
rect 2004 19400 2872 19428
rect 2004 19388 2010 19400
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 4798 19388 4804 19440
rect 4856 19428 4862 19440
rect 5442 19428 5448 19440
rect 4856 19400 5448 19428
rect 4856 19388 4862 19400
rect 5442 19388 5448 19400
rect 5500 19388 5506 19440
rect 7834 19388 7840 19440
rect 7892 19428 7898 19440
rect 8266 19428 8294 19468
rect 7892 19400 8294 19428
rect 7892 19388 7898 19400
rect 8386 19388 8392 19440
rect 8444 19388 8450 19440
rect 1486 19320 1492 19372
rect 1544 19360 1550 19372
rect 3326 19360 3332 19372
rect 1544 19332 3332 19360
rect 1544 19320 1550 19332
rect 3326 19320 3332 19332
rect 3384 19320 3390 19372
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 4706 19360 4712 19372
rect 3752 19332 4712 19360
rect 3752 19320 3758 19332
rect 4706 19320 4712 19332
rect 4764 19320 4770 19372
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 8404 19360 8432 19388
rect 7484 19332 8432 19360
rect 8496 19360 8524 19468
rect 8754 19456 8760 19508
rect 8812 19456 8818 19508
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8904 19468 9413 19496
rect 8904 19456 8910 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 9401 19459 9459 19465
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 10042 19496 10048 19508
rect 9824 19468 10048 19496
rect 9824 19456 9830 19468
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10410 19456 10416 19508
rect 10468 19496 10474 19508
rect 10781 19499 10839 19505
rect 10781 19496 10793 19499
rect 10468 19468 10793 19496
rect 10468 19456 10474 19468
rect 10781 19465 10793 19468
rect 10827 19465 10839 19499
rect 10781 19459 10839 19465
rect 11790 19456 11796 19508
rect 11848 19456 11854 19508
rect 8772 19428 8800 19456
rect 9677 19431 9735 19437
rect 9677 19428 9689 19431
rect 8772 19400 9689 19428
rect 9677 19397 9689 19400
rect 9723 19397 9735 19431
rect 9677 19391 9735 19397
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8496 19332 8769 19360
rect 1578 19252 1584 19304
rect 1636 19252 1642 19304
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 1857 19295 1915 19301
rect 1857 19261 1869 19295
rect 1903 19292 1915 19295
rect 1946 19292 1952 19304
rect 1903 19264 1952 19292
rect 1903 19261 1915 19264
rect 1857 19255 1915 19261
rect 1780 19224 1808 19255
rect 1946 19252 1952 19264
rect 2004 19252 2010 19304
rect 2225 19295 2283 19301
rect 2225 19261 2237 19295
rect 2271 19292 2283 19295
rect 2958 19292 2964 19304
rect 2271 19264 2964 19292
rect 2271 19261 2283 19264
rect 2225 19255 2283 19261
rect 2958 19252 2964 19264
rect 3016 19252 3022 19304
rect 5534 19252 5540 19304
rect 5592 19252 5598 19304
rect 5626 19252 5632 19304
rect 5684 19292 5690 19304
rect 5721 19295 5779 19301
rect 5721 19292 5733 19295
rect 5684 19264 5733 19292
rect 5684 19252 5690 19264
rect 5721 19261 5733 19264
rect 5767 19261 5779 19295
rect 5721 19255 5779 19261
rect 1780 19196 2452 19224
rect 2314 19116 2320 19168
rect 2372 19116 2378 19168
rect 2424 19156 2452 19196
rect 2498 19184 2504 19236
rect 2556 19184 2562 19236
rect 3050 19184 3056 19236
rect 3108 19224 3114 19236
rect 3510 19224 3516 19236
rect 3108 19196 3516 19224
rect 3108 19184 3114 19196
rect 3510 19184 3516 19196
rect 3568 19184 3574 19236
rect 4982 19156 4988 19168
rect 2424 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5736 19156 5764 19255
rect 6454 19252 6460 19304
rect 6512 19252 6518 19304
rect 6546 19252 6552 19304
rect 6604 19301 6610 19304
rect 6604 19295 6632 19301
rect 6620 19261 6632 19295
rect 6604 19255 6632 19261
rect 6604 19252 6610 19255
rect 6730 19252 6736 19304
rect 6788 19252 6794 19304
rect 7484 19301 7512 19332
rect 7469 19295 7527 19301
rect 7469 19261 7481 19295
rect 7515 19261 7527 19295
rect 7469 19255 7527 19261
rect 7650 19252 7656 19304
rect 7708 19252 7714 19304
rect 7926 19252 7932 19304
rect 7984 19252 7990 19304
rect 8110 19252 8116 19304
rect 8168 19252 8174 19304
rect 8220 19301 8248 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 9122 19320 9128 19372
rect 9180 19320 9186 19372
rect 9582 19320 9588 19372
rect 9640 19320 9646 19372
rect 9950 19320 9956 19372
rect 10008 19320 10014 19372
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 8294 19252 8300 19304
rect 8352 19292 8358 19304
rect 8389 19295 8447 19301
rect 8389 19292 8401 19295
rect 8352 19264 8401 19292
rect 8352 19252 8358 19264
rect 8389 19261 8401 19264
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 8570 19252 8576 19304
rect 8628 19252 8634 19304
rect 8665 19295 8723 19301
rect 8665 19261 8677 19295
rect 8711 19261 8723 19295
rect 8665 19255 8723 19261
rect 8941 19295 8999 19301
rect 8941 19261 8953 19295
rect 8987 19261 8999 19295
rect 8941 19255 8999 19261
rect 8680 19168 8708 19255
rect 6638 19156 6644 19168
rect 5736 19128 6644 19156
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 7190 19116 7196 19168
rect 7248 19156 7254 19168
rect 7377 19159 7435 19165
rect 7377 19156 7389 19159
rect 7248 19128 7389 19156
rect 7248 19116 7254 19128
rect 7377 19125 7389 19128
rect 7423 19125 7435 19159
rect 7377 19119 7435 19125
rect 8662 19116 8668 19168
rect 8720 19116 8726 19168
rect 8956 19156 8984 19255
rect 9306 19252 9312 19304
rect 9364 19252 9370 19304
rect 9486 19295 9544 19301
rect 9486 19261 9498 19295
rect 9532 19292 9544 19295
rect 9600 19292 9628 19320
rect 9532 19264 9628 19292
rect 9532 19261 9544 19264
rect 9486 19255 9544 19261
rect 9122 19184 9128 19236
rect 9180 19224 9186 19236
rect 9508 19224 9536 19255
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 9861 19295 9919 19301
rect 9861 19292 9873 19295
rect 9824 19264 9873 19292
rect 9824 19252 9830 19264
rect 9861 19261 9873 19264
rect 9907 19261 9919 19295
rect 9968 19292 9996 19320
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9968 19264 10241 19292
rect 9861 19255 9919 19261
rect 10229 19261 10241 19264
rect 10275 19261 10287 19295
rect 10229 19255 10287 19261
rect 10502 19252 10508 19304
rect 10560 19252 10566 19304
rect 10594 19252 10600 19304
rect 10652 19252 10658 19304
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19292 10931 19295
rect 11238 19292 11244 19304
rect 10919 19264 11244 19292
rect 10919 19261 10931 19264
rect 10873 19255 10931 19261
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 11698 19252 11704 19304
rect 11756 19252 11762 19304
rect 11974 19252 11980 19304
rect 12032 19252 12038 19304
rect 12250 19252 12256 19304
rect 12308 19252 12314 19304
rect 9180 19196 9536 19224
rect 9180 19184 9186 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 9953 19227 10011 19233
rect 9953 19224 9965 19227
rect 9640 19196 9965 19224
rect 9640 19184 9646 19196
rect 9953 19193 9965 19196
rect 9999 19193 10011 19227
rect 9953 19187 10011 19193
rect 10045 19227 10103 19233
rect 10045 19193 10057 19227
rect 10091 19224 10103 19227
rect 10321 19227 10379 19233
rect 10321 19224 10333 19227
rect 10091 19196 10333 19224
rect 10091 19193 10103 19196
rect 10045 19187 10103 19193
rect 10321 19193 10333 19196
rect 10367 19193 10379 19227
rect 10321 19187 10379 19193
rect 11054 19184 11060 19236
rect 11112 19224 11118 19236
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 11112 19196 11161 19224
rect 11112 19184 11118 19196
rect 11149 19193 11161 19196
rect 11195 19193 11207 19227
rect 11149 19187 11207 19193
rect 11517 19227 11575 19233
rect 11517 19193 11529 19227
rect 11563 19224 11575 19227
rect 12268 19224 12296 19252
rect 11563 19196 12296 19224
rect 11563 19193 11575 19196
rect 11517 19187 11575 19193
rect 11606 19156 11612 19168
rect 8956 19128 11612 19156
rect 11606 19116 11612 19128
rect 11664 19116 11670 19168
rect 12161 19159 12219 19165
rect 12161 19125 12173 19159
rect 12207 19156 12219 19159
rect 12250 19156 12256 19168
rect 12207 19128 12256 19156
rect 12207 19125 12219 19128
rect 12161 19119 12219 19125
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 552 19066 12604 19088
rect 552 19014 4322 19066
rect 4374 19014 4386 19066
rect 4438 19014 4450 19066
rect 4502 19014 4514 19066
rect 4566 19014 4578 19066
rect 4630 19014 10722 19066
rect 10774 19014 10786 19066
rect 10838 19014 10850 19066
rect 10902 19014 10914 19066
rect 10966 19014 10978 19066
rect 11030 19014 12604 19066
rect 552 18992 12604 19014
rect 2041 18955 2099 18961
rect 2041 18921 2053 18955
rect 2087 18952 2099 18955
rect 2130 18952 2136 18964
rect 2087 18924 2136 18952
rect 2087 18921 2099 18924
rect 2041 18915 2099 18921
rect 2130 18912 2136 18924
rect 2188 18912 2194 18964
rect 2774 18912 2780 18964
rect 2832 18912 2838 18964
rect 2958 18912 2964 18964
rect 3016 18952 3022 18964
rect 6546 18952 6552 18964
rect 3016 18924 3648 18952
rect 3016 18912 3022 18924
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 2792 18884 2820 18912
rect 3237 18887 3295 18893
rect 1820 18856 2728 18884
rect 2792 18856 3004 18884
rect 1820 18844 1826 18856
rect 1394 18776 1400 18828
rect 1452 18776 1458 18828
rect 1578 18776 1584 18828
rect 1636 18776 1642 18828
rect 2225 18819 2283 18825
rect 2225 18785 2237 18819
rect 2271 18816 2283 18819
rect 2314 18816 2320 18828
rect 2271 18788 2320 18816
rect 2271 18785 2283 18788
rect 2225 18779 2283 18785
rect 2314 18776 2320 18788
rect 2372 18816 2378 18828
rect 2593 18819 2651 18825
rect 2593 18816 2605 18819
rect 2372 18788 2605 18816
rect 2372 18776 2378 18788
rect 2593 18785 2605 18788
rect 2639 18785 2651 18819
rect 2700 18816 2728 18856
rect 2976 18825 3004 18856
rect 3237 18853 3249 18887
rect 3283 18884 3295 18887
rect 3510 18884 3516 18896
rect 3283 18856 3516 18884
rect 3283 18853 3295 18856
rect 3237 18847 3295 18853
rect 3510 18844 3516 18856
rect 3568 18844 3574 18896
rect 3620 18884 3648 18924
rect 5828 18924 6552 18952
rect 4433 18887 4491 18893
rect 4433 18884 4445 18887
rect 3620 18856 4445 18884
rect 2777 18819 2835 18825
rect 2777 18816 2789 18819
rect 2700 18788 2789 18816
rect 2593 18779 2651 18785
rect 2777 18785 2789 18788
rect 2823 18785 2835 18819
rect 2777 18779 2835 18785
rect 2961 18819 3019 18825
rect 2961 18785 2973 18819
rect 3007 18785 3019 18819
rect 2961 18779 3019 18785
rect 3050 18776 3056 18828
rect 3108 18776 3114 18828
rect 3142 18776 3148 18828
rect 3200 18776 3206 18828
rect 3620 18825 3648 18856
rect 4433 18853 4445 18856
rect 4479 18853 4491 18887
rect 4433 18847 4491 18853
rect 5000 18856 5396 18884
rect 3421 18819 3479 18825
rect 3421 18785 3433 18819
rect 3467 18785 3479 18819
rect 3421 18779 3479 18785
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18785 3663 18819
rect 3605 18779 3663 18785
rect 3789 18819 3847 18825
rect 3789 18785 3801 18819
rect 3835 18816 3847 18819
rect 4522 18816 4528 18828
rect 3835 18788 4528 18816
rect 3835 18785 3847 18788
rect 3789 18779 3847 18785
rect 934 18708 940 18760
rect 992 18708 998 18760
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 1688 18680 1716 18711
rect 1946 18708 1952 18760
rect 2004 18748 2010 18760
rect 2130 18748 2136 18760
rect 2004 18720 2136 18748
rect 2004 18708 2010 18720
rect 2130 18708 2136 18720
rect 2188 18748 2194 18760
rect 2501 18751 2559 18757
rect 2501 18748 2513 18751
rect 2188 18720 2513 18748
rect 2188 18708 2194 18720
rect 2501 18717 2513 18720
rect 2547 18748 2559 18751
rect 3436 18748 3464 18779
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 4614 18776 4620 18828
rect 4672 18776 4678 18828
rect 5000 18825 5028 18856
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18785 5043 18819
rect 4985 18779 5043 18785
rect 5169 18819 5227 18825
rect 5169 18785 5181 18819
rect 5215 18816 5227 18819
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 5215 18788 5273 18816
rect 5215 18785 5227 18788
rect 5169 18779 5227 18785
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 3694 18748 3700 18760
rect 2547 18720 3372 18748
rect 3436 18720 3700 18748
rect 2547 18717 2559 18720
rect 2501 18711 2559 18717
rect 492 18652 1716 18680
rect 3344 18680 3372 18720
rect 3694 18708 3700 18720
rect 3752 18748 3758 18760
rect 4338 18748 4344 18760
rect 3752 18720 4344 18748
rect 3752 18708 3758 18720
rect 4338 18708 4344 18720
rect 4396 18708 4402 18760
rect 4801 18751 4859 18757
rect 4801 18717 4813 18751
rect 4847 18717 4859 18751
rect 4801 18711 4859 18717
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 5074 18748 5080 18760
rect 4939 18720 5080 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 3786 18680 3792 18692
rect 3344 18652 3792 18680
rect 492 18408 520 18652
rect 3786 18640 3792 18652
rect 3844 18640 3850 18692
rect 4816 18680 4844 18711
rect 5074 18708 5080 18720
rect 5132 18708 5138 18760
rect 4982 18680 4988 18692
rect 4816 18652 4988 18680
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 2406 18572 2412 18624
rect 2464 18572 2470 18624
rect 3418 18572 3424 18624
rect 3476 18572 3482 18624
rect 3602 18572 3608 18624
rect 3660 18612 3666 18624
rect 3697 18615 3755 18621
rect 3697 18612 3709 18615
rect 3660 18584 3709 18612
rect 3660 18572 3666 18584
rect 3697 18581 3709 18584
rect 3743 18581 3755 18615
rect 5368 18612 5396 18856
rect 5442 18844 5448 18896
rect 5500 18844 5506 18896
rect 5626 18776 5632 18828
rect 5684 18776 5690 18828
rect 5828 18825 5856 18924
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7929 18955 7987 18961
rect 7929 18952 7941 18955
rect 7064 18924 7941 18952
rect 7064 18912 7070 18924
rect 7929 18921 7941 18924
rect 7975 18921 7987 18955
rect 7929 18915 7987 18921
rect 8110 18912 8116 18964
rect 8168 18952 8174 18964
rect 8938 18952 8944 18964
rect 8168 18924 8944 18952
rect 8168 18912 8174 18924
rect 8938 18912 8944 18924
rect 8996 18912 9002 18964
rect 9490 18952 9496 18964
rect 9048 18924 9496 18952
rect 8662 18844 8668 18896
rect 8720 18884 8726 18896
rect 9048 18884 9076 18924
rect 9490 18912 9496 18924
rect 9548 18912 9554 18964
rect 9582 18912 9588 18964
rect 9640 18912 9646 18964
rect 9766 18912 9772 18964
rect 9824 18912 9830 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 9916 18924 10364 18952
rect 9916 18912 9922 18924
rect 8720 18856 9076 18884
rect 8720 18844 8726 18856
rect 9122 18844 9128 18896
rect 9180 18884 9186 18896
rect 9306 18884 9312 18896
rect 9180 18856 9312 18884
rect 9180 18844 9186 18856
rect 9306 18844 9312 18856
rect 9364 18844 9370 18896
rect 9398 18844 9404 18896
rect 9456 18884 9462 18896
rect 10336 18893 10364 18924
rect 12158 18912 12164 18964
rect 12216 18912 12222 18964
rect 10321 18887 10379 18893
rect 9456 18856 9996 18884
rect 9456 18844 9462 18856
rect 5813 18819 5871 18825
rect 5813 18785 5825 18819
rect 5859 18785 5871 18819
rect 5813 18779 5871 18785
rect 6822 18776 6828 18828
rect 6880 18825 6886 18828
rect 6880 18819 6908 18825
rect 6896 18785 6908 18819
rect 6880 18779 6908 18785
rect 6880 18776 6886 18779
rect 7006 18776 7012 18828
rect 7064 18776 7070 18828
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 5534 18708 5540 18760
rect 5592 18748 5598 18760
rect 5997 18751 6055 18757
rect 5997 18748 6009 18751
rect 5592 18720 6009 18748
rect 5592 18708 5598 18720
rect 5997 18717 6009 18720
rect 6043 18717 6055 18751
rect 5997 18711 6055 18717
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6457 18751 6515 18757
rect 6457 18748 6469 18751
rect 6236 18720 6469 18748
rect 6236 18708 6242 18720
rect 6457 18717 6469 18720
rect 6503 18717 6515 18751
rect 6733 18751 6791 18757
rect 6733 18748 6745 18751
rect 6457 18711 6515 18717
rect 6564 18720 6745 18748
rect 6086 18640 6092 18692
rect 6144 18680 6150 18692
rect 6564 18680 6592 18720
rect 6733 18717 6745 18720
rect 6779 18748 6791 18751
rect 7745 18751 7803 18757
rect 7745 18748 7757 18751
rect 6779 18720 7757 18748
rect 6779 18717 6791 18720
rect 6733 18711 6791 18717
rect 7745 18717 7757 18720
rect 7791 18717 7803 18751
rect 7745 18711 7803 18717
rect 6144 18652 6592 18680
rect 6144 18640 6150 18652
rect 7558 18612 7564 18624
rect 5368 18584 7564 18612
rect 3697 18575 3755 18581
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 7650 18572 7656 18624
rect 7708 18572 7714 18624
rect 8128 18612 8156 18779
rect 8202 18776 8208 18828
rect 8260 18816 8266 18828
rect 8297 18819 8355 18825
rect 8297 18816 8309 18819
rect 8260 18788 8309 18816
rect 8260 18776 8266 18788
rect 8297 18785 8309 18788
rect 8343 18785 8355 18819
rect 8297 18779 8355 18785
rect 8386 18776 8392 18828
rect 8444 18776 8450 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 9416 18816 9444 18844
rect 8619 18788 9444 18816
rect 9493 18819 9551 18825
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 9493 18785 9505 18819
rect 9539 18816 9551 18819
rect 9677 18819 9735 18825
rect 9539 18788 9628 18816
rect 9539 18785 9551 18788
rect 9493 18779 9551 18785
rect 9398 18708 9404 18760
rect 9456 18748 9462 18760
rect 9494 18748 9522 18779
rect 9456 18720 9522 18748
rect 9600 18748 9628 18788
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 9858 18816 9864 18828
rect 9723 18788 9864 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 9968 18825 9996 18856
rect 10321 18853 10333 18887
rect 10367 18853 10379 18887
rect 10321 18847 10379 18853
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 10042 18776 10048 18828
rect 10100 18816 10106 18828
rect 10229 18819 10287 18825
rect 10229 18816 10241 18819
rect 10100 18788 10241 18816
rect 10100 18776 10106 18788
rect 10229 18785 10241 18788
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 10410 18776 10416 18828
rect 10468 18816 10474 18828
rect 10505 18819 10563 18825
rect 10505 18816 10517 18819
rect 10468 18788 10517 18816
rect 10468 18776 10474 18788
rect 10505 18785 10517 18788
rect 10551 18785 10563 18819
rect 10505 18779 10563 18785
rect 10594 18776 10600 18828
rect 10652 18776 10658 18828
rect 11606 18776 11612 18828
rect 11664 18776 11670 18828
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 12250 18776 12256 18828
rect 12308 18776 12314 18828
rect 10137 18751 10195 18757
rect 10137 18748 10149 18751
rect 9600 18720 10149 18748
rect 9456 18708 9462 18720
rect 10137 18717 10149 18720
rect 10183 18717 10195 18751
rect 10137 18711 10195 18717
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11517 18751 11575 18757
rect 11517 18748 11529 18751
rect 11112 18720 11529 18748
rect 11112 18708 11118 18720
rect 11517 18717 11529 18720
rect 11563 18717 11575 18751
rect 11517 18711 11575 18717
rect 11974 18708 11980 18760
rect 12032 18708 12038 18760
rect 8205 18683 8263 18689
rect 8205 18649 8217 18683
rect 8251 18680 8263 18683
rect 8251 18652 9628 18680
rect 8251 18649 8263 18652
rect 8205 18643 8263 18649
rect 8757 18615 8815 18621
rect 8757 18612 8769 18615
rect 8128 18584 8769 18612
rect 8757 18581 8769 18584
rect 8803 18612 8815 18615
rect 9030 18612 9036 18624
rect 8803 18584 9036 18612
rect 8803 18581 8815 18584
rect 8757 18575 8815 18581
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 9600 18612 9628 18652
rect 9674 18640 9680 18692
rect 9732 18680 9738 18692
rect 10321 18683 10379 18689
rect 10321 18680 10333 18683
rect 9732 18652 10333 18680
rect 9732 18640 9738 18652
rect 10321 18649 10333 18652
rect 10367 18649 10379 18683
rect 10321 18643 10379 18649
rect 11606 18612 11612 18624
rect 9600 18584 11612 18612
rect 11606 18572 11612 18584
rect 11664 18572 11670 18624
rect 552 18522 12604 18544
rect 552 18470 3662 18522
rect 3714 18470 3726 18522
rect 3778 18470 3790 18522
rect 3842 18470 3854 18522
rect 3906 18470 3918 18522
rect 3970 18470 10062 18522
rect 10114 18470 10126 18522
rect 10178 18470 10190 18522
rect 10242 18470 10254 18522
rect 10306 18470 10318 18522
rect 10370 18470 12604 18522
rect 552 18448 12604 18470
rect 845 18411 903 18417
rect 845 18408 857 18411
rect 492 18380 857 18408
rect 845 18377 857 18380
rect 891 18377 903 18411
rect 845 18371 903 18377
rect 1578 18368 1584 18420
rect 1636 18408 1642 18420
rect 2317 18411 2375 18417
rect 2317 18408 2329 18411
rect 1636 18380 2329 18408
rect 1636 18368 1642 18380
rect 2240 18272 2268 18380
rect 2317 18377 2329 18380
rect 2363 18377 2375 18411
rect 2317 18371 2375 18377
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 3881 18411 3939 18417
rect 3881 18408 3893 18411
rect 2464 18380 3893 18408
rect 2464 18368 2470 18380
rect 3881 18377 3893 18380
rect 3927 18377 3939 18411
rect 3881 18371 3939 18377
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 6178 18408 6184 18420
rect 5868 18380 6184 18408
rect 5868 18368 5874 18380
rect 6178 18368 6184 18380
rect 6236 18368 6242 18420
rect 7561 18411 7619 18417
rect 7561 18377 7573 18411
rect 7607 18408 7619 18411
rect 8294 18408 8300 18420
rect 7607 18380 8300 18408
rect 7607 18377 7619 18380
rect 7561 18371 7619 18377
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8386 18368 8392 18420
rect 8444 18368 8450 18420
rect 10410 18368 10416 18420
rect 10468 18368 10474 18420
rect 11977 18411 12035 18417
rect 11977 18377 11989 18411
rect 12023 18408 12035 18411
rect 12066 18408 12072 18420
rect 12023 18380 12072 18408
rect 12023 18377 12035 18380
rect 11977 18371 12035 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 2590 18300 2596 18352
rect 2648 18340 2654 18352
rect 2685 18343 2743 18349
rect 2685 18340 2697 18343
rect 2648 18312 2697 18340
rect 2648 18300 2654 18312
rect 2685 18309 2697 18312
rect 2731 18309 2743 18343
rect 4246 18340 4252 18352
rect 2685 18303 2743 18309
rect 3712 18312 4252 18340
rect 3050 18272 3056 18284
rect 2148 18244 2268 18272
rect 2976 18244 3056 18272
rect 1969 18207 2027 18213
rect 1969 18173 1981 18207
rect 2015 18204 2027 18207
rect 2148 18204 2176 18244
rect 2015 18176 2176 18204
rect 2015 18173 2027 18176
rect 1969 18167 2027 18173
rect 2222 18164 2228 18216
rect 2280 18164 2286 18216
rect 2314 18164 2320 18216
rect 2372 18204 2378 18216
rect 2501 18207 2559 18213
rect 2501 18204 2513 18207
rect 2372 18176 2513 18204
rect 2372 18164 2378 18176
rect 2501 18173 2513 18176
rect 2547 18173 2559 18207
rect 2777 18207 2835 18213
rect 2777 18204 2789 18207
rect 2501 18167 2559 18173
rect 2700 18176 2789 18204
rect 1302 18096 1308 18148
rect 1360 18136 1366 18148
rect 1578 18136 1584 18148
rect 1360 18108 1584 18136
rect 1360 18096 1366 18108
rect 1578 18096 1584 18108
rect 1636 18096 1642 18148
rect 2130 18096 2136 18148
rect 2188 18136 2194 18148
rect 2700 18136 2728 18176
rect 2777 18173 2789 18176
rect 2823 18204 2835 18207
rect 2866 18204 2872 18216
rect 2823 18176 2872 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 2976 18136 3004 18244
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3513 18275 3571 18281
rect 3513 18272 3525 18275
rect 3160 18244 3525 18272
rect 2188 18108 2728 18136
rect 2792 18108 3004 18136
rect 2188 18096 2194 18108
rect 2792 18080 2820 18108
rect 3050 18096 3056 18148
rect 3108 18136 3114 18148
rect 3160 18136 3188 18244
rect 3513 18241 3525 18244
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 3602 18232 3608 18284
rect 3660 18232 3666 18284
rect 3712 18216 3740 18312
rect 4246 18300 4252 18312
rect 4304 18340 4310 18352
rect 4798 18340 4804 18352
rect 4304 18312 4804 18340
rect 4304 18300 4310 18312
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 9125 18343 9183 18349
rect 9125 18340 9137 18343
rect 5408 18312 9137 18340
rect 5408 18300 5414 18312
rect 9125 18309 9137 18312
rect 9171 18309 9183 18343
rect 9125 18303 9183 18309
rect 9214 18300 9220 18352
rect 9272 18340 9278 18352
rect 9766 18340 9772 18352
rect 9272 18312 9772 18340
rect 9272 18300 9278 18312
rect 9766 18300 9772 18312
rect 9824 18300 9830 18352
rect 11241 18343 11299 18349
rect 11241 18340 11253 18343
rect 11164 18312 11253 18340
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 3329 18207 3387 18213
rect 3329 18204 3341 18207
rect 3108 18108 3188 18136
rect 3252 18176 3341 18204
rect 3108 18096 3114 18108
rect 2774 18028 2780 18080
rect 2832 18028 2838 18080
rect 3252 18068 3280 18176
rect 3329 18173 3341 18176
rect 3375 18173 3387 18207
rect 3329 18167 3387 18173
rect 3421 18207 3479 18213
rect 3421 18173 3433 18207
rect 3467 18204 3479 18207
rect 3694 18204 3700 18216
rect 3467 18176 3700 18204
rect 3467 18173 3479 18176
rect 3421 18167 3479 18173
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 3804 18204 3832 18235
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 4120 18244 4476 18272
rect 4120 18232 4126 18244
rect 4157 18207 4215 18213
rect 4157 18204 4169 18207
rect 3804 18176 4169 18204
rect 4157 18173 4169 18176
rect 4203 18173 4215 18207
rect 4157 18167 4215 18173
rect 4246 18164 4252 18216
rect 4304 18164 4310 18216
rect 4448 18213 4476 18244
rect 7926 18232 7932 18284
rect 7984 18232 7990 18284
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8757 18275 8815 18281
rect 8757 18272 8769 18275
rect 8076 18244 8769 18272
rect 8076 18232 8082 18244
rect 8757 18241 8769 18244
rect 8803 18272 8815 18275
rect 11054 18272 11060 18284
rect 8803 18244 11060 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 4433 18207 4491 18213
rect 4433 18173 4445 18207
rect 4479 18173 4491 18207
rect 4433 18167 4491 18173
rect 5810 18164 5816 18216
rect 5868 18204 5874 18216
rect 6733 18207 6791 18213
rect 6733 18204 6745 18207
rect 5868 18176 6745 18204
rect 5868 18164 5874 18176
rect 6733 18173 6745 18176
rect 6779 18204 6791 18207
rect 7650 18204 7656 18216
rect 6779 18176 7656 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 7837 18207 7895 18213
rect 7837 18204 7849 18207
rect 7800 18176 7849 18204
rect 7800 18164 7806 18176
rect 7837 18173 7849 18176
rect 7883 18173 7895 18207
rect 7944 18204 7972 18232
rect 8573 18207 8631 18213
rect 8573 18204 8585 18207
rect 7944 18176 8585 18204
rect 7837 18167 7895 18173
rect 8573 18173 8585 18176
rect 8619 18173 8631 18207
rect 8573 18167 8631 18173
rect 8662 18164 8668 18216
rect 8720 18164 8726 18216
rect 8849 18207 8907 18213
rect 8849 18173 8861 18207
rect 8895 18204 8907 18207
rect 8938 18204 8944 18216
rect 8895 18176 8944 18204
rect 8895 18173 8907 18176
rect 8849 18167 8907 18173
rect 8938 18164 8944 18176
rect 8996 18164 9002 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9272 18176 9321 18204
rect 9272 18164 9278 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 9398 18164 9404 18216
rect 9456 18164 9462 18216
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18204 10379 18207
rect 10410 18204 10416 18216
rect 10367 18176 10416 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 10410 18164 10416 18176
rect 10468 18164 10474 18216
rect 10502 18164 10508 18216
rect 10560 18164 10566 18216
rect 10980 18213 11008 18244
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 10965 18207 11023 18213
rect 10965 18173 10977 18207
rect 11011 18173 11023 18207
rect 10965 18167 11023 18173
rect 3510 18096 3516 18148
rect 3568 18136 3574 18148
rect 3881 18139 3939 18145
rect 3881 18136 3893 18139
rect 3568 18108 3893 18136
rect 3568 18096 3574 18108
rect 3881 18105 3893 18108
rect 3927 18105 3939 18139
rect 3881 18099 3939 18105
rect 3988 18108 4292 18136
rect 3326 18068 3332 18080
rect 3252 18040 3332 18068
rect 3326 18028 3332 18040
rect 3384 18068 3390 18080
rect 3988 18068 4016 18108
rect 4264 18080 4292 18108
rect 4614 18096 4620 18148
rect 4672 18136 4678 18148
rect 4672 18108 5028 18136
rect 4672 18096 4678 18108
rect 5000 18080 5028 18108
rect 5626 18096 5632 18148
rect 5684 18136 5690 18148
rect 6549 18139 6607 18145
rect 6549 18136 6561 18139
rect 5684 18108 6561 18136
rect 5684 18096 5690 18108
rect 6549 18105 6561 18108
rect 6595 18136 6607 18139
rect 7098 18136 7104 18148
rect 6595 18108 7104 18136
rect 6595 18105 6607 18108
rect 6549 18099 6607 18105
rect 7098 18096 7104 18108
rect 7156 18096 7162 18148
rect 7190 18096 7196 18148
rect 7248 18096 7254 18148
rect 7374 18096 7380 18148
rect 7432 18096 7438 18148
rect 9122 18096 9128 18148
rect 9180 18096 9186 18148
rect 11164 18136 11192 18312
rect 11241 18309 11253 18312
rect 11287 18309 11299 18343
rect 11241 18303 11299 18309
rect 11790 18300 11796 18352
rect 11848 18340 11854 18352
rect 11885 18343 11943 18349
rect 11885 18340 11897 18343
rect 11848 18312 11897 18340
rect 11848 18300 11854 18312
rect 11885 18309 11897 18312
rect 11931 18309 11943 18343
rect 11885 18303 11943 18309
rect 12250 18272 12256 18284
rect 11256 18244 12256 18272
rect 11256 18213 11284 18244
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18173 11299 18207
rect 11241 18167 11299 18173
rect 11698 18164 11704 18216
rect 11756 18164 11762 18216
rect 11974 18164 11980 18216
rect 12032 18164 12038 18216
rect 12434 18136 12440 18148
rect 9646 18108 11100 18136
rect 11164 18108 12440 18136
rect 3384 18040 4016 18068
rect 3384 18028 3390 18040
rect 4062 18028 4068 18080
rect 4120 18028 4126 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4341 18071 4399 18077
rect 4341 18068 4353 18071
rect 4304 18040 4353 18068
rect 4304 18028 4310 18040
rect 4341 18037 4353 18040
rect 4387 18037 4399 18071
rect 4341 18031 4399 18037
rect 4522 18028 4528 18080
rect 4580 18068 4586 18080
rect 4798 18068 4804 18080
rect 4580 18040 4804 18068
rect 4580 18028 4586 18040
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 4982 18028 4988 18080
rect 5040 18068 5046 18080
rect 6454 18068 6460 18080
rect 5040 18040 6460 18068
rect 5040 18028 5046 18040
rect 6454 18028 6460 18040
rect 6512 18028 6518 18080
rect 6914 18028 6920 18080
rect 6972 18028 6978 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7208 18068 7236 18096
rect 7064 18040 7236 18068
rect 7064 18028 7070 18040
rect 8018 18028 8024 18080
rect 8076 18028 8082 18080
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 9646 18068 9674 18108
rect 11072 18077 11100 18108
rect 12434 18096 12440 18108
rect 12492 18096 12498 18148
rect 8444 18040 9674 18068
rect 11057 18071 11115 18077
rect 8444 18028 8450 18040
rect 11057 18037 11069 18071
rect 11103 18068 11115 18071
rect 11514 18068 11520 18080
rect 11103 18040 11520 18068
rect 11103 18037 11115 18040
rect 11057 18031 11115 18037
rect 11514 18028 11520 18040
rect 11572 18028 11578 18080
rect 552 17978 12604 18000
rect 552 17926 4322 17978
rect 4374 17926 4386 17978
rect 4438 17926 4450 17978
rect 4502 17926 4514 17978
rect 4566 17926 4578 17978
rect 4630 17926 10722 17978
rect 10774 17926 10786 17978
rect 10838 17926 10850 17978
rect 10902 17926 10914 17978
rect 10966 17926 10978 17978
rect 11030 17926 12604 17978
rect 552 17904 12604 17926
rect 2961 17867 3019 17873
rect 2961 17833 2973 17867
rect 3007 17864 3019 17867
rect 3142 17864 3148 17876
rect 3007 17836 3148 17864
rect 3007 17833 3019 17836
rect 2961 17827 3019 17833
rect 3142 17824 3148 17836
rect 3200 17824 3206 17876
rect 3234 17824 3240 17876
rect 3292 17864 3298 17876
rect 3418 17864 3424 17876
rect 3292 17836 3424 17864
rect 3292 17824 3298 17836
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 3694 17864 3700 17876
rect 3620 17836 3700 17864
rect 2314 17756 2320 17808
rect 2372 17796 2378 17808
rect 2372 17768 2544 17796
rect 2372 17756 2378 17768
rect 2516 17737 2544 17768
rect 3326 17756 3332 17808
rect 3384 17756 3390 17808
rect 3620 17796 3648 17836
rect 3694 17824 3700 17836
rect 3752 17864 3758 17876
rect 3878 17864 3884 17876
rect 3752 17836 3884 17864
rect 3752 17824 3758 17836
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4246 17864 4252 17876
rect 3988 17836 4252 17864
rect 3988 17796 4016 17836
rect 4246 17824 4252 17836
rect 4304 17824 4310 17876
rect 4430 17824 4436 17876
rect 4488 17864 4494 17876
rect 6270 17864 6276 17876
rect 4488 17836 6276 17864
rect 4488 17824 4494 17836
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 7742 17864 7748 17876
rect 6840 17836 7748 17864
rect 3528 17768 3648 17796
rect 3712 17768 4016 17796
rect 1969 17731 2027 17737
rect 1969 17697 1981 17731
rect 2015 17728 2027 17731
rect 2501 17731 2559 17737
rect 2015 17700 2360 17728
rect 2015 17697 2027 17700
rect 1969 17691 2027 17697
rect 2222 17620 2228 17672
rect 2280 17620 2286 17672
rect 845 17527 903 17533
rect 845 17524 857 17527
rect 492 17496 857 17524
rect 492 17184 520 17496
rect 845 17493 857 17496
rect 891 17493 903 17527
rect 845 17487 903 17493
rect 1302 17484 1308 17536
rect 1360 17524 1366 17536
rect 2332 17533 2360 17700
rect 2501 17697 2513 17731
rect 2547 17697 2559 17731
rect 2501 17691 2559 17697
rect 2590 17688 2596 17740
rect 2648 17688 2654 17740
rect 2777 17731 2835 17737
rect 2777 17697 2789 17731
rect 2823 17728 2835 17731
rect 2866 17728 2872 17740
rect 2823 17700 2872 17728
rect 2823 17697 2835 17700
rect 2777 17691 2835 17697
rect 2866 17688 2872 17700
rect 2924 17688 2930 17740
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 3344 17728 3372 17756
rect 3528 17737 3556 17768
rect 3099 17700 3372 17728
rect 3513 17731 3571 17737
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 3513 17697 3525 17731
rect 3559 17697 3571 17731
rect 3513 17691 3571 17697
rect 3605 17731 3663 17737
rect 3605 17697 3617 17731
rect 3651 17728 3663 17731
rect 3712 17728 3740 17768
rect 4062 17756 4068 17808
rect 4120 17756 4126 17808
rect 4985 17799 5043 17805
rect 4985 17765 4997 17799
rect 5031 17796 5043 17799
rect 5258 17796 5264 17808
rect 5031 17768 5264 17796
rect 5031 17765 5043 17768
rect 4985 17759 5043 17765
rect 5258 17756 5264 17768
rect 5316 17796 5322 17808
rect 5442 17796 5448 17808
rect 5316 17768 5448 17796
rect 5316 17756 5322 17768
rect 5442 17756 5448 17768
rect 5500 17756 5506 17808
rect 5718 17756 5724 17808
rect 5776 17796 5782 17808
rect 6546 17796 6552 17808
rect 5776 17768 6552 17796
rect 5776 17756 5782 17768
rect 3651 17700 3740 17728
rect 3973 17731 4031 17737
rect 3651 17697 3663 17700
rect 3605 17691 3663 17697
rect 3973 17697 3985 17731
rect 4019 17728 4031 17731
rect 4080 17728 4108 17756
rect 4019 17700 4108 17728
rect 4019 17697 4031 17700
rect 3973 17691 4031 17697
rect 4246 17688 4252 17740
rect 4304 17688 4310 17740
rect 4709 17731 4767 17737
rect 4709 17697 4721 17731
rect 4755 17728 4767 17731
rect 4798 17728 4804 17740
rect 4755 17700 4804 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 4798 17688 4804 17700
rect 4856 17688 4862 17740
rect 5169 17731 5227 17737
rect 5169 17697 5181 17731
rect 5215 17697 5227 17731
rect 5169 17691 5227 17697
rect 5353 17731 5411 17737
rect 5353 17697 5365 17731
rect 5399 17728 5411 17731
rect 5813 17731 5871 17737
rect 5813 17728 5825 17731
rect 5399 17700 5825 17728
rect 5399 17697 5411 17700
rect 5353 17691 5411 17697
rect 5813 17697 5825 17700
rect 5859 17697 5871 17731
rect 5813 17691 5871 17697
rect 2608 17536 2636 17688
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3467 17632 3556 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3528 17592 3556 17632
rect 3878 17620 3884 17672
rect 3936 17660 3942 17672
rect 4065 17663 4123 17669
rect 4065 17660 4077 17663
rect 3936 17632 4077 17660
rect 3936 17620 3942 17632
rect 4065 17629 4077 17632
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17660 4215 17663
rect 5184 17660 5212 17691
rect 5994 17688 6000 17740
rect 6052 17688 6058 17740
rect 6196 17737 6224 17768
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 6840 17805 6868 17836
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 7926 17824 7932 17876
rect 7984 17864 7990 17876
rect 7984 17836 8984 17864
rect 7984 17824 7990 17836
rect 6825 17799 6883 17805
rect 6825 17765 6837 17799
rect 6871 17765 6883 17799
rect 6825 17759 6883 17765
rect 6181 17731 6239 17737
rect 6181 17697 6193 17731
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 6365 17731 6423 17737
rect 6365 17697 6377 17731
rect 6411 17728 6423 17731
rect 6454 17728 6460 17740
rect 6411 17700 6460 17728
rect 6411 17697 6423 17700
rect 6365 17691 6423 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6840 17728 6868 17759
rect 7006 17756 7012 17808
rect 7064 17756 7070 17808
rect 7469 17799 7527 17805
rect 7469 17765 7481 17799
rect 7515 17796 7527 17799
rect 7558 17796 7564 17808
rect 7515 17768 7564 17796
rect 7515 17765 7527 17768
rect 7469 17759 7527 17765
rect 7558 17756 7564 17768
rect 7616 17756 7622 17808
rect 8386 17796 8392 17808
rect 7944 17768 8392 17796
rect 6564 17700 6868 17728
rect 7653 17731 7711 17737
rect 4203 17632 4292 17660
rect 5184 17632 5580 17660
rect 4203 17629 4215 17632
rect 4157 17623 4215 17629
rect 4264 17604 4292 17632
rect 5552 17604 5580 17632
rect 6086 17620 6092 17672
rect 6144 17620 6150 17672
rect 6270 17620 6276 17672
rect 6328 17660 6334 17672
rect 6564 17660 6592 17700
rect 7653 17697 7665 17731
rect 7699 17697 7711 17731
rect 7653 17691 7711 17697
rect 6328 17632 6592 17660
rect 6641 17663 6699 17669
rect 6328 17620 6334 17632
rect 6641 17629 6653 17663
rect 6687 17660 6699 17663
rect 7668 17660 7696 17691
rect 7742 17688 7748 17740
rect 7800 17728 7806 17740
rect 7944 17737 7972 17768
rect 8386 17756 8392 17768
rect 8444 17756 8450 17808
rect 8665 17799 8723 17805
rect 8665 17765 8677 17799
rect 8711 17796 8723 17799
rect 8754 17796 8760 17808
rect 8711 17768 8760 17796
rect 8711 17765 8723 17768
rect 8665 17759 8723 17765
rect 8754 17756 8760 17768
rect 8812 17756 8818 17808
rect 7837 17731 7895 17737
rect 7837 17728 7849 17731
rect 7800 17700 7849 17728
rect 7800 17688 7806 17700
rect 7837 17697 7849 17700
rect 7883 17697 7895 17731
rect 7837 17691 7895 17697
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17697 7987 17731
rect 7929 17691 7987 17697
rect 7944 17660 7972 17691
rect 8202 17688 8208 17740
rect 8260 17688 8266 17740
rect 8481 17731 8539 17737
rect 8481 17697 8493 17731
rect 8527 17728 8539 17731
rect 8570 17728 8576 17740
rect 8527 17700 8576 17728
rect 8527 17697 8539 17700
rect 8481 17691 8539 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 8956 17737 8984 17836
rect 9030 17824 9036 17876
rect 9088 17824 9094 17876
rect 9122 17824 9128 17876
rect 9180 17864 9186 17876
rect 9585 17867 9643 17873
rect 9585 17864 9597 17867
rect 9180 17836 9597 17864
rect 9180 17824 9186 17836
rect 9585 17833 9597 17836
rect 9631 17833 9643 17867
rect 9585 17827 9643 17833
rect 9858 17824 9864 17876
rect 9916 17864 9922 17876
rect 10134 17864 10140 17876
rect 9916 17836 10140 17864
rect 9916 17824 9922 17836
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 10594 17824 10600 17876
rect 10652 17864 10658 17876
rect 10781 17867 10839 17873
rect 10781 17864 10793 17867
rect 10652 17836 10793 17864
rect 10652 17824 10658 17836
rect 10781 17833 10793 17836
rect 10827 17833 10839 17867
rect 10781 17827 10839 17833
rect 11514 17824 11520 17876
rect 11572 17864 11578 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 11572 17836 11805 17864
rect 11572 17824 11578 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 11793 17827 11851 17833
rect 9048 17796 9076 17824
rect 9309 17799 9367 17805
rect 9309 17796 9321 17799
rect 9048 17768 9321 17796
rect 9309 17765 9321 17768
rect 9355 17765 9367 17799
rect 9309 17759 9367 17765
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 9824 17768 10640 17796
rect 9824 17756 9830 17768
rect 9122 17737 9128 17740
rect 8941 17731 8999 17737
rect 8941 17697 8953 17731
rect 8987 17697 8999 17731
rect 8941 17691 8999 17697
rect 9089 17731 9128 17737
rect 9089 17697 9101 17731
rect 9089 17691 9128 17697
rect 6687 17632 7696 17660
rect 7760 17632 7972 17660
rect 8021 17663 8079 17669
rect 6687 17629 6699 17632
rect 6641 17623 6699 17629
rect 3528 17564 3924 17592
rect 2317 17527 2375 17533
rect 2317 17524 2329 17527
rect 1360 17496 2329 17524
rect 1360 17484 1366 17496
rect 2317 17493 2329 17496
rect 2363 17493 2375 17527
rect 2317 17487 2375 17493
rect 2590 17484 2596 17536
rect 2648 17484 2654 17536
rect 2682 17484 2688 17536
rect 2740 17484 2746 17536
rect 3142 17484 3148 17536
rect 3200 17484 3206 17536
rect 3234 17484 3240 17536
rect 3292 17524 3298 17536
rect 3789 17527 3847 17533
rect 3789 17524 3801 17527
rect 3292 17496 3801 17524
rect 3292 17484 3298 17496
rect 3789 17493 3801 17496
rect 3835 17493 3847 17527
rect 3896 17524 3924 17564
rect 3970 17552 3976 17604
rect 4028 17592 4034 17604
rect 4246 17592 4252 17604
rect 4028 17564 4252 17592
rect 4028 17552 4034 17564
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 5442 17592 5448 17604
rect 4448 17564 5448 17592
rect 4448 17524 4476 17564
rect 5442 17552 5448 17564
rect 5500 17552 5506 17604
rect 5534 17552 5540 17604
rect 5592 17592 5598 17604
rect 7374 17592 7380 17604
rect 5592 17564 7380 17592
rect 5592 17552 5598 17564
rect 7374 17552 7380 17564
rect 7432 17552 7438 17604
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 7760 17592 7788 17632
rect 8021 17629 8033 17663
rect 8067 17629 8079 17663
rect 8021 17623 8079 17629
rect 7708 17564 7788 17592
rect 7708 17552 7714 17564
rect 7834 17552 7840 17604
rect 7892 17592 7898 17604
rect 8036 17592 8064 17623
rect 8386 17620 8392 17672
rect 8444 17660 8450 17672
rect 8956 17660 8984 17691
rect 9122 17688 9128 17691
rect 9180 17688 9186 17740
rect 9217 17731 9275 17737
rect 9217 17697 9229 17731
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 8444 17632 8984 17660
rect 9232 17660 9260 17691
rect 9398 17688 9404 17740
rect 9456 17737 9462 17740
rect 9456 17728 9464 17737
rect 9456 17700 9501 17728
rect 9456 17691 9464 17700
rect 9456 17688 9462 17691
rect 9582 17688 9588 17740
rect 9640 17728 9646 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9640 17700 9873 17728
rect 9640 17688 9646 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 9861 17691 9919 17697
rect 10134 17688 10140 17740
rect 10192 17688 10198 17740
rect 10612 17737 10640 17768
rect 10597 17731 10655 17737
rect 10597 17697 10609 17731
rect 10643 17697 10655 17731
rect 10597 17691 10655 17697
rect 11330 17688 11336 17740
rect 11388 17688 11394 17740
rect 11701 17731 11759 17737
rect 11701 17697 11713 17731
rect 11747 17728 11759 17731
rect 12526 17728 12532 17740
rect 11747 17700 12532 17728
rect 11747 17697 11759 17700
rect 11701 17691 11759 17697
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 9677 17663 9735 17669
rect 9677 17660 9689 17663
rect 9232 17632 9689 17660
rect 8444 17620 8450 17632
rect 9677 17629 9689 17632
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 9953 17663 10011 17669
rect 9953 17629 9965 17663
rect 9999 17629 10011 17663
rect 9953 17623 10011 17629
rect 10045 17663 10103 17669
rect 10045 17629 10057 17663
rect 10091 17629 10103 17663
rect 10045 17623 10103 17629
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10410 17660 10416 17672
rect 10367 17632 10416 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 7892 17564 8064 17592
rect 8849 17595 8907 17601
rect 7892 17552 7898 17564
rect 8849 17561 8861 17595
rect 8895 17592 8907 17595
rect 9968 17592 9996 17623
rect 8895 17564 9996 17592
rect 10060 17592 10088 17623
rect 10410 17620 10416 17632
rect 10468 17620 10474 17672
rect 11422 17620 11428 17672
rect 11480 17620 11486 17672
rect 10594 17592 10600 17604
rect 10060 17564 10600 17592
rect 8895 17561 8907 17564
rect 8849 17555 8907 17561
rect 10594 17552 10600 17564
rect 10652 17552 10658 17604
rect 10965 17595 11023 17601
rect 10965 17561 10977 17595
rect 11011 17561 11023 17595
rect 10965 17555 11023 17561
rect 3896 17496 4476 17524
rect 3789 17487 3847 17493
rect 4522 17484 4528 17536
rect 4580 17484 4586 17536
rect 4798 17484 4804 17536
rect 4856 17524 4862 17536
rect 5166 17524 5172 17536
rect 4856 17496 5172 17524
rect 4856 17484 4862 17496
rect 5166 17484 5172 17496
rect 5224 17524 5230 17536
rect 6549 17527 6607 17533
rect 6549 17524 6561 17527
rect 5224 17496 6561 17524
rect 5224 17484 5230 17496
rect 6549 17493 6561 17496
rect 6595 17493 6607 17527
rect 6549 17487 6607 17493
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 7156 17496 7205 17524
rect 7156 17484 7162 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 8389 17527 8447 17533
rect 8389 17493 8401 17527
rect 8435 17524 8447 17527
rect 8754 17524 8760 17536
rect 8435 17496 8760 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 9766 17524 9772 17536
rect 9272 17496 9772 17524
rect 9272 17484 9278 17496
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 10413 17527 10471 17533
rect 10413 17493 10425 17527
rect 10459 17524 10471 17527
rect 10502 17524 10508 17536
rect 10459 17496 10508 17524
rect 10459 17493 10471 17496
rect 10413 17487 10471 17493
rect 10502 17484 10508 17496
rect 10560 17524 10566 17536
rect 10980 17524 11008 17555
rect 10560 17496 11008 17524
rect 10560 17484 10566 17496
rect 552 17434 12604 17456
rect 552 17382 3662 17434
rect 3714 17382 3726 17434
rect 3778 17382 3790 17434
rect 3842 17382 3854 17434
rect 3906 17382 3918 17434
rect 3970 17382 10062 17434
rect 10114 17382 10126 17434
rect 10178 17382 10190 17434
rect 10242 17382 10254 17434
rect 10306 17382 10318 17434
rect 10370 17382 12604 17434
rect 552 17360 12604 17382
rect 2501 17323 2559 17329
rect 2501 17289 2513 17323
rect 2547 17320 2559 17323
rect 2682 17320 2688 17332
rect 2547 17292 2688 17320
rect 2547 17289 2559 17292
rect 2501 17283 2559 17289
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 4249 17323 4307 17329
rect 4249 17320 4261 17323
rect 3384 17292 4261 17320
rect 3384 17280 3390 17292
rect 4249 17289 4261 17292
rect 4295 17289 4307 17323
rect 4249 17283 4307 17289
rect 5258 17280 5264 17332
rect 5316 17280 5322 17332
rect 6270 17320 6276 17332
rect 5368 17292 6276 17320
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 2314 17252 2320 17264
rect 1636 17224 2320 17252
rect 1636 17212 1642 17224
rect 2314 17212 2320 17224
rect 2372 17212 2378 17264
rect 2590 17212 2596 17264
rect 2648 17212 2654 17264
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 4430 17252 4436 17264
rect 3936 17224 4436 17252
rect 3936 17212 3942 17224
rect 4430 17212 4436 17224
rect 4488 17212 4494 17264
rect 4982 17212 4988 17264
rect 5040 17212 5046 17264
rect 1213 17187 1271 17193
rect 1213 17184 1225 17187
rect 492 17156 1225 17184
rect 1213 17153 1225 17156
rect 1259 17153 1271 17187
rect 1213 17147 1271 17153
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 4522 17184 4528 17196
rect 2188 17156 2452 17184
rect 2188 17144 2194 17156
rect 1302 17076 1308 17128
rect 1360 17076 1366 17128
rect 1394 17076 1400 17128
rect 1452 17116 1458 17128
rect 1489 17119 1547 17125
rect 1489 17116 1501 17119
rect 1452 17088 1501 17116
rect 1452 17076 1458 17088
rect 1489 17085 1501 17088
rect 1535 17085 1547 17119
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 1489 17079 1547 17085
rect 2056 17088 2237 17116
rect 1946 17008 1952 17060
rect 2004 17008 2010 17060
rect 2056 16980 2084 17088
rect 2225 17085 2237 17088
rect 2271 17085 2283 17119
rect 2424 17116 2452 17156
rect 4172 17156 4528 17184
rect 2501 17119 2559 17125
rect 2501 17116 2513 17119
rect 2424 17088 2513 17116
rect 2225 17079 2283 17085
rect 2501 17085 2513 17088
rect 2547 17116 2559 17119
rect 2593 17119 2651 17125
rect 2593 17116 2605 17119
rect 2547 17088 2605 17116
rect 2547 17085 2559 17088
rect 2501 17079 2559 17085
rect 2593 17085 2605 17088
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3142 17116 3148 17128
rect 2915 17088 3148 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 3142 17076 3148 17088
rect 3200 17076 3206 17128
rect 4172 17125 4200 17156
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 5000 17184 5028 17212
rect 5000 17156 5120 17184
rect 4157 17119 4215 17125
rect 4157 17085 4169 17119
rect 4203 17085 4215 17119
rect 4157 17079 4215 17085
rect 4341 17119 4399 17125
rect 4341 17085 4353 17119
rect 4387 17116 4399 17119
rect 4798 17116 4804 17128
rect 4387 17088 4804 17116
rect 4387 17085 4399 17088
rect 4341 17079 4399 17085
rect 4798 17076 4804 17088
rect 4856 17076 4862 17128
rect 4982 17076 4988 17128
rect 5040 17076 5046 17128
rect 5092 17125 5120 17156
rect 5368 17125 5396 17292
rect 6270 17280 6276 17292
rect 6328 17280 6334 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17320 6423 17323
rect 6454 17320 6460 17332
rect 6411 17292 6460 17320
rect 6411 17289 6423 17292
rect 6365 17283 6423 17289
rect 6454 17280 6460 17292
rect 6512 17280 6518 17332
rect 6549 17323 6607 17329
rect 6549 17289 6561 17323
rect 6595 17320 6607 17323
rect 6638 17320 6644 17332
rect 6595 17292 6644 17320
rect 6595 17289 6607 17292
rect 6549 17283 6607 17289
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7558 17320 7564 17332
rect 7064 17292 7564 17320
rect 7064 17280 7070 17292
rect 7558 17280 7564 17292
rect 7616 17280 7622 17332
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 7892 17292 8524 17320
rect 7892 17280 7898 17292
rect 5445 17255 5503 17261
rect 5445 17221 5457 17255
rect 5491 17252 5503 17255
rect 5491 17224 6316 17252
rect 5491 17221 5503 17224
rect 5445 17215 5503 17221
rect 6288 17184 6316 17224
rect 6932 17224 8432 17252
rect 6932 17184 6960 17224
rect 5644 17156 6224 17184
rect 6288 17156 6960 17184
rect 7009 17187 7067 17193
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5644 17125 5672 17156
rect 5629 17119 5687 17125
rect 5629 17116 5641 17119
rect 5592 17088 5641 17116
rect 5592 17076 5598 17088
rect 5629 17085 5641 17088
rect 5675 17085 5687 17119
rect 5629 17079 5687 17085
rect 5718 17076 5724 17128
rect 5776 17116 5782 17128
rect 5813 17119 5871 17125
rect 5813 17116 5825 17119
rect 5776 17088 5825 17116
rect 5776 17076 5782 17088
rect 5813 17085 5825 17088
rect 5859 17085 5871 17119
rect 5813 17079 5871 17085
rect 5902 17076 5908 17128
rect 5960 17118 5966 17128
rect 6196 17125 6224 17156
rect 7009 17153 7021 17187
rect 7055 17184 7067 17187
rect 7190 17184 7196 17196
rect 7055 17156 7196 17184
rect 7055 17153 7067 17156
rect 7009 17147 7067 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7742 17144 7748 17196
rect 7800 17184 7806 17196
rect 7800 17156 8064 17184
rect 7800 17144 7806 17156
rect 6089 17119 6147 17125
rect 6089 17118 6101 17119
rect 5960 17090 6101 17118
rect 5960 17076 5966 17090
rect 6089 17085 6101 17090
rect 6135 17085 6147 17119
rect 6089 17079 6147 17085
rect 6181 17119 6239 17125
rect 6181 17085 6193 17119
rect 6227 17085 6239 17119
rect 6457 17119 6515 17125
rect 6457 17116 6469 17119
rect 6181 17079 6239 17085
rect 6380 17088 6469 17116
rect 2130 17008 2136 17060
rect 2188 17048 2194 17060
rect 2317 17051 2375 17057
rect 2317 17048 2329 17051
rect 2188 17020 2329 17048
rect 2188 17008 2194 17020
rect 2317 17017 2329 17020
rect 2363 17017 2375 17051
rect 2317 17011 2375 17017
rect 2406 17008 2412 17060
rect 2464 17048 2470 17060
rect 2777 17051 2835 17057
rect 2777 17048 2789 17051
rect 2464 17020 2789 17048
rect 2464 17008 2470 17020
rect 2777 17017 2789 17020
rect 2823 17048 2835 17051
rect 3234 17048 3240 17060
rect 2823 17020 3240 17048
rect 2823 17017 2835 17020
rect 2777 17011 2835 17017
rect 3234 17008 3240 17020
rect 3292 17008 3298 17060
rect 3326 16980 3332 16992
rect 2056 16952 3332 16980
rect 3326 16940 3332 16952
rect 3384 16940 3390 16992
rect 4798 16940 4804 16992
rect 4856 16940 4862 16992
rect 5902 16940 5908 16992
rect 5960 16940 5966 16992
rect 6380 16980 6408 17088
rect 6457 17085 6469 17088
rect 6503 17085 6515 17119
rect 6457 17079 6515 17085
rect 6546 17076 6552 17128
rect 6604 17118 6610 17128
rect 6733 17119 6791 17125
rect 6733 17118 6745 17119
rect 6604 17090 6745 17118
rect 6604 17076 6610 17090
rect 6733 17085 6745 17090
rect 6779 17085 6791 17119
rect 6733 17079 6791 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7101 17119 7159 17125
rect 7101 17085 7113 17119
rect 7147 17116 7159 17119
rect 7374 17116 7380 17128
rect 7147 17088 7380 17116
rect 7147 17085 7159 17088
rect 7101 17079 7159 17085
rect 6546 16980 6552 16992
rect 6380 16952 6552 16980
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 6850 16980 6878 17079
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7650 17076 7656 17128
rect 7708 17076 7714 17128
rect 7837 17119 7895 17125
rect 7837 17085 7849 17119
rect 7883 17085 7895 17119
rect 7837 17079 7895 17085
rect 7190 17008 7196 17060
rect 7248 17048 7254 17060
rect 7852 17048 7880 17079
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 8036 17125 8064 17156
rect 8021 17119 8079 17125
rect 8021 17085 8033 17119
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8202 17076 8208 17128
rect 8260 17076 8266 17128
rect 8404 17125 8432 17224
rect 8496 17184 8524 17292
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 10594 17320 10600 17332
rect 9180 17292 10600 17320
rect 9180 17280 9186 17292
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11054 17280 11060 17332
rect 11112 17320 11118 17332
rect 11112 17292 11836 17320
rect 11112 17280 11118 17292
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9732 17224 10180 17252
rect 9732 17212 9738 17224
rect 10152 17196 10180 17224
rect 10410 17212 10416 17264
rect 10468 17212 10474 17264
rect 11422 17212 11428 17264
rect 11480 17212 11486 17264
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 8496 17156 8769 17184
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 8389 17079 8447 17085
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17085 8631 17119
rect 8573 17079 8631 17085
rect 8665 17119 8723 17125
rect 8665 17085 8677 17119
rect 8711 17116 8723 17119
rect 8846 17116 8852 17128
rect 8711 17088 8852 17116
rect 8711 17085 8723 17088
rect 8665 17079 8723 17085
rect 8588 17048 8616 17079
rect 8846 17076 8852 17088
rect 8904 17076 8910 17128
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17085 8999 17119
rect 8941 17079 8999 17085
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17116 9551 17119
rect 9674 17116 9680 17128
rect 9539 17088 9680 17116
rect 9539 17085 9551 17088
rect 9493 17079 9551 17085
rect 8956 17048 8984 17079
rect 9674 17076 9680 17088
rect 9732 17076 9738 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 9968 17116 9996 17147
rect 10134 17144 10140 17196
rect 10192 17144 10198 17196
rect 11054 17184 11060 17196
rect 10612 17156 11060 17184
rect 9824 17088 9996 17116
rect 10045 17119 10103 17125
rect 9824 17076 9830 17088
rect 10045 17085 10057 17119
rect 10091 17116 10103 17119
rect 10226 17116 10232 17128
rect 10091 17088 10232 17116
rect 10091 17085 10103 17088
rect 10045 17079 10103 17085
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 10612 17125 10640 17156
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11440 17184 11468 17212
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11440 17156 11529 17184
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10781 17119 10839 17125
rect 10781 17085 10793 17119
rect 10827 17116 10839 17119
rect 10827 17088 11376 17116
rect 10827 17085 10839 17088
rect 10781 17079 10839 17085
rect 10689 17051 10747 17057
rect 7248 17020 8616 17048
rect 8680 17020 10364 17048
rect 7248 17008 7254 17020
rect 6696 16952 6878 16980
rect 6696 16940 6702 16952
rect 7466 16940 7472 16992
rect 7524 16940 7530 16992
rect 7650 16940 7656 16992
rect 7708 16980 7714 16992
rect 8680 16980 8708 17020
rect 10336 16992 10364 17020
rect 10689 17017 10701 17051
rect 10735 17048 10747 17051
rect 10873 17051 10931 17057
rect 10873 17048 10885 17051
rect 10735 17020 10885 17048
rect 10735 17017 10747 17020
rect 10689 17011 10747 17017
rect 10873 17017 10885 17020
rect 10919 17048 10931 17051
rect 11238 17048 11244 17060
rect 10919 17020 11244 17048
rect 10919 17017 10931 17020
rect 10873 17011 10931 17017
rect 11238 17008 11244 17020
rect 11296 17008 11302 17060
rect 11348 17048 11376 17088
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11701 17119 11759 17125
rect 11701 17116 11713 17119
rect 11480 17088 11713 17116
rect 11480 17076 11486 17088
rect 11701 17085 11713 17088
rect 11747 17085 11759 17119
rect 11808 17116 11836 17292
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 11808 17088 12081 17116
rect 11701 17079 11759 17085
rect 12069 17085 12081 17088
rect 12115 17085 12127 17119
rect 12069 17079 12127 17085
rect 11885 17051 11943 17057
rect 11885 17048 11897 17051
rect 11348 17020 11897 17048
rect 11885 17017 11897 17020
rect 11931 17048 11943 17051
rect 12158 17048 12164 17060
rect 11931 17020 12164 17048
rect 11931 17017 11943 17020
rect 11885 17011 11943 17017
rect 12158 17008 12164 17020
rect 12216 17008 12222 17060
rect 7708 16952 8708 16980
rect 7708 16940 7714 16952
rect 8846 16940 8852 16992
rect 8904 16980 8910 16992
rect 9125 16983 9183 16989
rect 9125 16980 9137 16983
rect 8904 16952 9137 16980
rect 8904 16940 8910 16952
rect 9125 16949 9137 16952
rect 9171 16949 9183 16983
rect 9125 16943 9183 16949
rect 9306 16940 9312 16992
rect 9364 16940 9370 16992
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 10042 16980 10048 16992
rect 9723 16952 10048 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10318 16940 10324 16992
rect 10376 16940 10382 16992
rect 10410 16940 10416 16992
rect 10468 16980 10474 16992
rect 11149 16983 11207 16989
rect 11149 16980 11161 16983
rect 10468 16952 11161 16980
rect 10468 16940 10474 16952
rect 11149 16949 11161 16952
rect 11195 16949 11207 16983
rect 11149 16943 11207 16949
rect 552 16890 12604 16912
rect 552 16838 4322 16890
rect 4374 16838 4386 16890
rect 4438 16838 4450 16890
rect 4502 16838 4514 16890
rect 4566 16838 4578 16890
rect 4630 16838 10722 16890
rect 10774 16838 10786 16890
rect 10838 16838 10850 16890
rect 10902 16838 10914 16890
rect 10966 16838 10978 16890
rect 11030 16838 12604 16890
rect 552 16816 12604 16838
rect 1762 16736 1768 16788
rect 1820 16776 1826 16788
rect 2406 16776 2412 16788
rect 1820 16748 2412 16776
rect 1820 16736 1826 16748
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2498 16736 2504 16788
rect 2556 16776 2562 16788
rect 2774 16776 2780 16788
rect 2556 16748 2780 16776
rect 2556 16736 2562 16748
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 3789 16779 3847 16785
rect 3789 16745 3801 16779
rect 3835 16776 3847 16779
rect 4062 16776 4068 16788
rect 3835 16748 4068 16776
rect 3835 16745 3847 16748
rect 3789 16739 3847 16745
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4249 16779 4307 16785
rect 4249 16776 4261 16779
rect 4172 16748 4261 16776
rect 934 16668 940 16720
rect 992 16668 998 16720
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 4172 16717 4200 16748
rect 4249 16745 4261 16748
rect 4295 16776 4307 16779
rect 4706 16776 4712 16788
rect 4295 16748 4712 16776
rect 4295 16745 4307 16748
rect 4249 16739 4307 16745
rect 4706 16736 4712 16748
rect 4764 16736 4770 16788
rect 5810 16776 5816 16788
rect 5275 16748 5816 16776
rect 3973 16711 4031 16717
rect 3973 16708 3985 16711
rect 3936 16680 3985 16708
rect 3936 16668 3942 16680
rect 3973 16677 3985 16680
rect 4019 16677 4031 16711
rect 3973 16671 4031 16677
rect 4157 16711 4215 16717
rect 4157 16677 4169 16711
rect 4203 16677 4215 16711
rect 4798 16708 4804 16720
rect 4157 16671 4215 16677
rect 4356 16680 4804 16708
rect 1210 16600 1216 16652
rect 1268 16640 1274 16652
rect 1397 16643 1455 16649
rect 1397 16640 1409 16643
rect 1268 16612 1409 16640
rect 1268 16600 1274 16612
rect 1397 16609 1409 16612
rect 1443 16609 1455 16643
rect 1397 16603 1455 16609
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16640 1639 16643
rect 1762 16640 1768 16652
rect 1627 16612 1768 16640
rect 1627 16609 1639 16612
rect 1581 16603 1639 16609
rect 1762 16600 1768 16612
rect 1820 16600 1826 16652
rect 4356 16640 4384 16680
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 4982 16668 4988 16720
rect 5040 16668 5046 16720
rect 4264 16612 4384 16640
rect 4525 16643 4583 16649
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2130 16572 2136 16584
rect 1719 16544 2136 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 4264 16581 4292 16612
rect 4525 16609 4537 16643
rect 4571 16640 4583 16643
rect 5074 16640 5080 16652
rect 4571 16612 5080 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 5074 16600 5080 16612
rect 5132 16600 5138 16652
rect 5275 16649 5303 16748
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 7834 16776 7840 16788
rect 7392 16748 7840 16776
rect 5626 16668 5632 16720
rect 5684 16668 5690 16720
rect 6454 16668 6460 16720
rect 6512 16708 6518 16720
rect 7392 16708 7420 16748
rect 7834 16736 7840 16748
rect 7892 16736 7898 16788
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7984 16748 8217 16776
rect 7984 16736 7990 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 9582 16776 9588 16788
rect 8803 16748 9588 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 6512 16680 7420 16708
rect 8220 16708 8248 16739
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 9674 16736 9680 16788
rect 9732 16776 9738 16788
rect 9732 16748 9812 16776
rect 9732 16736 9738 16748
rect 9784 16717 9812 16748
rect 10226 16736 10232 16788
rect 10284 16736 10290 16788
rect 10428 16748 10732 16776
rect 9769 16711 9827 16717
rect 8220 16680 9720 16708
rect 6512 16668 6518 16680
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 6273 16643 6331 16649
rect 6273 16609 6285 16643
rect 6319 16609 6331 16643
rect 6273 16603 6331 16609
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4430 16532 4436 16584
rect 4488 16532 4494 16584
rect 4985 16575 5043 16581
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 5368 16572 5396 16603
rect 4985 16535 5043 16541
rect 5092 16544 5396 16572
rect 5629 16575 5687 16581
rect 5000 16436 5028 16535
rect 5092 16516 5120 16544
rect 5629 16541 5641 16575
rect 5675 16572 5687 16575
rect 5902 16572 5908 16584
rect 5675 16544 5908 16572
rect 5675 16541 5687 16544
rect 5629 16535 5687 16541
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 5074 16464 5080 16516
rect 5132 16464 5138 16516
rect 5169 16507 5227 16513
rect 5169 16473 5181 16507
rect 5215 16504 5227 16507
rect 5718 16504 5724 16516
rect 5215 16476 5724 16504
rect 5215 16473 5227 16476
rect 5169 16467 5227 16473
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 6288 16504 6316 16603
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 6641 16643 6699 16649
rect 6641 16640 6653 16643
rect 6420 16612 6653 16640
rect 6420 16600 6426 16612
rect 6641 16609 6653 16612
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 6454 16532 6460 16584
rect 6512 16532 6518 16584
rect 6546 16532 6552 16584
rect 6604 16532 6610 16584
rect 6656 16572 6684 16603
rect 6822 16600 6828 16652
rect 6880 16600 6886 16652
rect 7282 16600 7288 16652
rect 7340 16600 7346 16652
rect 7392 16640 7420 16680
rect 9692 16652 9720 16680
rect 9769 16677 9781 16711
rect 9815 16677 9827 16711
rect 9769 16671 9827 16677
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 10428 16708 10456 16748
rect 10704 16717 10732 16748
rect 11330 16736 11336 16788
rect 11388 16736 11394 16788
rect 10192 16680 10456 16708
rect 10689 16711 10747 16717
rect 10192 16668 10198 16680
rect 10689 16677 10701 16711
rect 10735 16677 10747 16711
rect 10689 16671 10747 16677
rect 7469 16643 7527 16649
rect 7469 16640 7481 16643
rect 7392 16612 7481 16640
rect 7469 16609 7481 16612
rect 7515 16609 7527 16643
rect 7469 16603 7527 16609
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 7742 16640 7748 16652
rect 7699 16612 7748 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 7742 16600 7748 16612
rect 7800 16600 7806 16652
rect 7837 16643 7895 16649
rect 7837 16609 7849 16643
rect 7883 16640 7895 16643
rect 8018 16640 8024 16652
rect 7883 16612 8024 16640
rect 7883 16609 7895 16612
rect 7837 16603 7895 16609
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 8294 16600 8300 16652
rect 8352 16600 8358 16652
rect 8570 16600 8576 16652
rect 8628 16600 8634 16652
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 8720 16612 8769 16640
rect 8720 16600 8726 16612
rect 8757 16609 8769 16612
rect 8803 16609 8815 16643
rect 8757 16603 8815 16609
rect 8849 16643 8907 16649
rect 8849 16609 8861 16643
rect 8895 16609 8907 16643
rect 8849 16603 8907 16609
rect 7006 16572 7012 16584
rect 6656 16544 7012 16572
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7561 16575 7619 16581
rect 7561 16572 7573 16575
rect 7300 16544 7573 16572
rect 7300 16516 7328 16544
rect 7561 16541 7573 16544
rect 7607 16541 7619 16575
rect 7561 16535 7619 16541
rect 8386 16532 8392 16584
rect 8444 16572 8450 16584
rect 8864 16572 8892 16603
rect 8938 16600 8944 16652
rect 8996 16600 9002 16652
rect 9030 16600 9036 16652
rect 9088 16600 9094 16652
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9582 16640 9588 16652
rect 9539 16612 9588 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 9674 16600 9680 16652
rect 9732 16600 9738 16652
rect 10505 16643 10563 16649
rect 10505 16609 10517 16643
rect 10551 16640 10563 16643
rect 10551 16612 10585 16640
rect 10551 16609 10563 16612
rect 10505 16603 10563 16609
rect 8444 16544 8892 16572
rect 9309 16575 9367 16581
rect 8444 16532 8450 16544
rect 9309 16541 9321 16575
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 6638 16504 6644 16516
rect 6013 16476 6224 16504
rect 6288 16476 6644 16504
rect 5258 16436 5264 16448
rect 5000 16408 5264 16436
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 5445 16439 5503 16445
rect 5445 16405 5457 16439
rect 5491 16436 5503 16439
rect 6013 16436 6041 16476
rect 5491 16408 6041 16436
rect 5491 16405 5503 16408
rect 5445 16399 5503 16405
rect 6086 16396 6092 16448
rect 6144 16396 6150 16448
rect 6196 16436 6224 16476
rect 6638 16464 6644 16476
rect 6696 16464 6702 16516
rect 7190 16504 7196 16516
rect 7024 16476 7196 16504
rect 7024 16436 7052 16476
rect 7190 16464 7196 16476
rect 7248 16464 7254 16516
rect 7282 16464 7288 16516
rect 7340 16464 7346 16516
rect 7374 16464 7380 16516
rect 7432 16504 7438 16516
rect 9324 16504 9352 16535
rect 9398 16532 9404 16584
rect 9456 16572 9462 16584
rect 9766 16572 9772 16584
rect 9456 16544 9772 16572
rect 9456 16532 9462 16544
rect 9766 16532 9772 16544
rect 9824 16532 9830 16584
rect 10520 16572 10548 16603
rect 11238 16600 11244 16652
rect 11296 16600 11302 16652
rect 11422 16600 11428 16652
rect 11480 16600 11486 16652
rect 11793 16643 11851 16649
rect 11793 16609 11805 16643
rect 11839 16640 11851 16643
rect 11882 16640 11888 16652
rect 11839 16612 11888 16640
rect 11839 16609 11851 16612
rect 11793 16603 11851 16609
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 11974 16600 11980 16652
rect 12032 16600 12038 16652
rect 12066 16600 12072 16652
rect 12124 16600 12130 16652
rect 12158 16572 12164 16584
rect 9968 16544 12164 16572
rect 9968 16504 9996 16544
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 7432 16476 9996 16504
rect 7432 16464 7438 16476
rect 10042 16464 10048 16516
rect 10100 16504 10106 16516
rect 10321 16507 10379 16513
rect 10321 16504 10333 16507
rect 10100 16476 10333 16504
rect 10100 16464 10106 16476
rect 10321 16473 10333 16476
rect 10367 16473 10379 16507
rect 12342 16504 12348 16516
rect 10321 16467 10379 16473
rect 10428 16476 12348 16504
rect 6196 16408 7052 16436
rect 7101 16439 7159 16445
rect 7101 16405 7113 16439
rect 7147 16436 7159 16439
rect 7650 16436 7656 16448
rect 7147 16408 7656 16436
rect 7147 16405 7159 16408
rect 7101 16399 7159 16405
rect 7650 16396 7656 16408
rect 7708 16396 7714 16448
rect 9582 16396 9588 16448
rect 9640 16436 9646 16448
rect 9766 16436 9772 16448
rect 9640 16408 9772 16436
rect 9640 16396 9646 16408
rect 9766 16396 9772 16408
rect 9824 16436 9830 16448
rect 10134 16436 10140 16448
rect 9824 16408 10140 16436
rect 9824 16396 9830 16408
rect 10134 16396 10140 16408
rect 10192 16396 10198 16448
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 10428 16436 10456 16476
rect 12342 16464 12348 16476
rect 12400 16464 12406 16516
rect 10284 16408 10456 16436
rect 10284 16396 10290 16408
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 552 16346 12604 16368
rect 552 16294 3662 16346
rect 3714 16294 3726 16346
rect 3778 16294 3790 16346
rect 3842 16294 3854 16346
rect 3906 16294 3918 16346
rect 3970 16294 10062 16346
rect 10114 16294 10126 16346
rect 10178 16294 10190 16346
rect 10242 16294 10254 16346
rect 10306 16294 10318 16346
rect 10370 16294 12604 16346
rect 552 16272 12604 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1946 16232 1952 16244
rect 1636 16204 1952 16232
rect 1636 16192 1642 16204
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2225 16235 2283 16241
rect 2225 16232 2237 16235
rect 2188 16204 2237 16232
rect 2188 16192 2194 16204
rect 2225 16201 2237 16204
rect 2271 16201 2283 16235
rect 2225 16195 2283 16201
rect 2774 16192 2780 16244
rect 2832 16192 2838 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6822 16232 6828 16244
rect 6227 16204 6828 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 8021 16235 8079 16241
rect 8021 16201 8033 16235
rect 8067 16232 8079 16235
rect 8202 16232 8208 16244
rect 8067 16204 8208 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8941 16235 8999 16241
rect 8941 16232 8953 16235
rect 8312 16204 8953 16232
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 8312 16164 8340 16204
rect 8941 16201 8953 16204
rect 8987 16201 8999 16235
rect 8941 16195 8999 16201
rect 9674 16192 9680 16244
rect 9732 16232 9738 16244
rect 9769 16235 9827 16241
rect 9769 16232 9781 16235
rect 9732 16204 9781 16232
rect 9732 16192 9738 16204
rect 9769 16201 9781 16204
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 11606 16192 11612 16244
rect 11664 16192 11670 16244
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 12066 16232 12072 16244
rect 12023 16204 12072 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12066 16192 12072 16204
rect 12124 16192 12130 16244
rect 6604 16136 8340 16164
rect 6604 16124 6610 16136
rect 8662 16124 8668 16176
rect 8720 16124 8726 16176
rect 10045 16167 10103 16173
rect 10045 16133 10057 16167
rect 10091 16164 10103 16167
rect 10318 16164 10324 16176
rect 10091 16136 10324 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10318 16124 10324 16136
rect 10376 16124 10382 16176
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 2869 16099 2927 16105
rect 2869 16096 2881 16099
rect 2740 16068 2881 16096
rect 2740 16056 2746 16068
rect 2869 16065 2881 16068
rect 2915 16065 2927 16099
rect 2869 16059 2927 16065
rect 845 16031 903 16037
rect 845 15997 857 16031
rect 891 16028 903 16031
rect 2222 16028 2228 16040
rect 891 16000 2228 16028
rect 891 15997 903 16000
rect 845 15991 903 15997
rect 2222 15988 2228 16000
rect 2280 15988 2286 16040
rect 2498 15988 2504 16040
rect 2556 16028 2562 16040
rect 2593 16031 2651 16037
rect 2593 16028 2605 16031
rect 2556 16000 2605 16028
rect 2556 15988 2562 16000
rect 2593 15997 2605 16000
rect 2639 15997 2651 16031
rect 2593 15991 2651 15997
rect 1112 15963 1170 15969
rect 1112 15929 1124 15963
rect 1158 15960 1170 15963
rect 1762 15960 1768 15972
rect 1158 15932 1768 15960
rect 1158 15929 1170 15932
rect 1112 15923 1170 15929
rect 1762 15920 1768 15932
rect 1820 15920 1826 15972
rect 2406 15852 2412 15904
rect 2464 15852 2470 15904
rect 2884 15892 2912 16059
rect 5074 16056 5080 16108
rect 5132 16096 5138 16108
rect 5902 16096 5908 16108
rect 5132 16068 5908 16096
rect 5132 16056 5138 16068
rect 5902 16056 5908 16068
rect 5960 16096 5966 16108
rect 7742 16096 7748 16108
rect 5960 16068 6592 16096
rect 5960 16056 5966 16068
rect 5810 15988 5816 16040
rect 5868 15988 5874 16040
rect 5997 16031 6055 16037
rect 5997 15997 6009 16031
rect 6043 16028 6055 16031
rect 6270 16028 6276 16040
rect 6043 16000 6276 16028
rect 6043 15997 6055 16000
rect 5997 15991 6055 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 6564 16037 6592 16068
rect 7024 16068 7748 16096
rect 7024 16040 7052 16068
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 8680 16096 8708 16124
rect 8352 16068 9444 16096
rect 8352 16056 8358 16068
rect 6549 16031 6607 16037
rect 6549 15997 6561 16031
rect 6595 15997 6607 16031
rect 6549 15991 6607 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 6914 16028 6920 16040
rect 6871 16000 6920 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 6914 15988 6920 16000
rect 6972 15988 6978 16040
rect 7006 15988 7012 16040
rect 7064 15988 7070 16040
rect 7098 15988 7104 16040
rect 7156 15988 7162 16040
rect 7190 15988 7196 16040
rect 7248 15988 7254 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 7340 16000 7389 16028
rect 7340 15988 7346 16000
rect 7377 15997 7389 16000
rect 7423 15997 7435 16031
rect 7377 15991 7435 15997
rect 7558 15988 7564 16040
rect 7616 16028 7622 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7616 16000 7849 16028
rect 7616 15988 7622 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 8389 16031 8447 16037
rect 8389 16028 8401 16031
rect 8076 16000 8401 16028
rect 8076 15988 8082 16000
rect 8389 15997 8401 16000
rect 8435 15997 8447 16031
rect 8389 15991 8447 15997
rect 8478 15988 8484 16040
rect 8536 15988 8542 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 5718 15920 5724 15972
rect 5776 15960 5782 15972
rect 7653 15963 7711 15969
rect 7653 15960 7665 15963
rect 5776 15932 7665 15960
rect 5776 15920 5782 15932
rect 7653 15929 7665 15932
rect 7699 15929 7711 15963
rect 7653 15923 7711 15929
rect 7926 15920 7932 15972
rect 7984 15960 7990 15972
rect 8680 15960 8708 15991
rect 8754 15988 8760 16040
rect 8812 15988 8818 16040
rect 9306 15988 9312 16040
rect 9364 15988 9370 16040
rect 9416 16037 9444 16068
rect 9582 16056 9588 16108
rect 9640 16096 9646 16108
rect 9640 16068 10456 16096
rect 9640 16056 9646 16068
rect 9401 16031 9459 16037
rect 9401 15997 9413 16031
rect 9447 15997 9459 16031
rect 9401 15991 9459 15997
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10321 16031 10379 16037
rect 10321 16028 10333 16031
rect 9732 16000 10333 16028
rect 9732 15988 9738 16000
rect 10321 15997 10333 16000
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 7984 15932 8708 15960
rect 9324 15960 9352 15988
rect 9953 15963 10011 15969
rect 9324 15932 9720 15960
rect 7984 15920 7990 15932
rect 5810 15892 5816 15904
rect 2884 15864 5816 15892
rect 5810 15852 5816 15864
rect 5868 15852 5874 15904
rect 6638 15852 6644 15904
rect 6696 15852 6702 15904
rect 7558 15852 7564 15904
rect 7616 15852 7622 15904
rect 9309 15895 9367 15901
rect 9309 15861 9321 15895
rect 9355 15892 9367 15895
rect 9398 15892 9404 15904
rect 9355 15864 9404 15892
rect 9355 15861 9367 15864
rect 9309 15855 9367 15861
rect 9398 15852 9404 15864
rect 9456 15852 9462 15904
rect 9582 15852 9588 15904
rect 9640 15852 9646 15904
rect 9692 15892 9720 15932
rect 9953 15929 9965 15963
rect 9999 15929 10011 15963
rect 9953 15923 10011 15929
rect 10045 15963 10103 15969
rect 10045 15929 10057 15963
rect 10091 15960 10103 15963
rect 10428 15960 10456 16068
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 16028 11575 16031
rect 11698 16028 11704 16040
rect 11563 16000 11704 16028
rect 11563 15997 11575 16000
rect 11517 15991 11575 15997
rect 11698 15988 11704 16000
rect 11756 15988 11762 16040
rect 11790 15988 11796 16040
rect 11848 15988 11854 16040
rect 11974 15988 11980 16040
rect 12032 16028 12038 16040
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 12032 16000 12081 16028
rect 12032 15988 12038 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 12069 15991 12127 15997
rect 10091 15932 10456 15960
rect 10091 15929 10103 15932
rect 10045 15923 10103 15929
rect 9748 15895 9806 15901
rect 9748 15892 9760 15895
rect 9692 15864 9760 15892
rect 9748 15861 9760 15864
rect 9794 15861 9806 15895
rect 9968 15892 9996 15923
rect 10134 15892 10140 15904
rect 9968 15864 10140 15892
rect 9748 15855 9806 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10226 15852 10232 15904
rect 10284 15852 10290 15904
rect 11514 15852 11520 15904
rect 11572 15852 11578 15904
rect 552 15802 12604 15824
rect 552 15750 4322 15802
rect 4374 15750 4386 15802
rect 4438 15750 4450 15802
rect 4502 15750 4514 15802
rect 4566 15750 4578 15802
rect 4630 15750 10722 15802
rect 10774 15750 10786 15802
rect 10838 15750 10850 15802
rect 10902 15750 10914 15802
rect 10966 15750 10978 15802
rect 11030 15750 12604 15802
rect 552 15728 12604 15750
rect 1670 15648 1676 15700
rect 1728 15648 1734 15700
rect 1762 15648 1768 15700
rect 1820 15648 1826 15700
rect 3510 15648 3516 15700
rect 3568 15648 3574 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4154 15688 4160 15700
rect 3927 15660 4160 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4154 15648 4160 15660
rect 4212 15648 4218 15700
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 7285 15691 7343 15697
rect 6236 15660 6500 15688
rect 6236 15648 6242 15660
rect 3145 15623 3203 15629
rect 3145 15620 3157 15623
rect 2792 15592 3157 15620
rect 1489 15555 1547 15561
rect 1489 15521 1501 15555
rect 1535 15552 1547 15555
rect 1949 15555 2007 15561
rect 1949 15552 1961 15555
rect 1535 15524 1961 15552
rect 1535 15521 1547 15524
rect 1489 15515 1547 15521
rect 1949 15521 1961 15524
rect 1995 15552 2007 15555
rect 2130 15552 2136 15564
rect 1995 15524 2136 15552
rect 1995 15521 2007 15524
rect 1949 15515 2007 15521
rect 2130 15512 2136 15524
rect 2188 15552 2194 15564
rect 2406 15552 2412 15564
rect 2188 15524 2412 15552
rect 2188 15512 2194 15524
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2498 15512 2504 15564
rect 2556 15512 2562 15564
rect 2682 15512 2688 15564
rect 2740 15512 2746 15564
rect 2792 15561 2820 15592
rect 3145 15589 3157 15592
rect 3191 15620 3203 15623
rect 3602 15620 3608 15632
rect 3191 15592 3608 15620
rect 3191 15589 3203 15592
rect 3145 15583 3203 15589
rect 3602 15580 3608 15592
rect 3660 15580 3666 15632
rect 5994 15580 6000 15632
rect 6052 15620 6058 15632
rect 6052 15592 6224 15620
rect 6052 15580 6058 15592
rect 2777 15555 2835 15561
rect 2777 15521 2789 15555
rect 2823 15521 2835 15555
rect 2777 15515 2835 15521
rect 3329 15555 3387 15561
rect 3329 15521 3341 15555
rect 3375 15552 3387 15555
rect 4246 15552 4252 15564
rect 3375 15524 4252 15552
rect 3375 15521 3387 15524
rect 3329 15515 3387 15521
rect 4246 15512 4252 15524
rect 4304 15552 4310 15564
rect 4614 15552 4620 15564
rect 4304 15524 4620 15552
rect 4304 15512 4310 15524
rect 4614 15512 4620 15524
rect 4672 15512 4678 15564
rect 4985 15555 5043 15561
rect 4985 15521 4997 15555
rect 5031 15552 5043 15555
rect 5074 15552 5080 15564
rect 5031 15524 5080 15552
rect 5031 15521 5043 15524
rect 4985 15515 5043 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 5169 15555 5227 15561
rect 5169 15521 5181 15555
rect 5215 15552 5227 15555
rect 5905 15555 5963 15561
rect 5905 15552 5917 15555
rect 5215 15524 5917 15552
rect 5215 15521 5227 15524
rect 5169 15515 5227 15521
rect 5905 15521 5917 15524
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 6086 15512 6092 15564
rect 6144 15512 6150 15564
rect 6196 15561 6224 15592
rect 6181 15555 6239 15561
rect 6181 15521 6193 15555
rect 6227 15521 6239 15555
rect 6181 15515 6239 15521
rect 6362 15512 6368 15564
rect 6420 15512 6426 15564
rect 6472 15561 6500 15660
rect 7285 15657 7297 15691
rect 7331 15688 7343 15691
rect 7331 15660 8432 15688
rect 7331 15657 7343 15660
rect 7285 15651 7343 15657
rect 8404 15620 8432 15660
rect 8478 15648 8484 15700
rect 8536 15648 8542 15700
rect 8662 15648 8668 15700
rect 8720 15648 8726 15700
rect 10226 15688 10232 15700
rect 8772 15660 10232 15688
rect 8772 15620 8800 15660
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 10781 15691 10839 15697
rect 10781 15657 10793 15691
rect 10827 15688 10839 15691
rect 11054 15688 11060 15700
rect 10827 15660 11060 15688
rect 10827 15657 10839 15660
rect 10781 15651 10839 15657
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11146 15648 11152 15700
rect 11204 15648 11210 15700
rect 11330 15648 11336 15700
rect 11388 15648 11394 15700
rect 11698 15648 11704 15700
rect 11756 15688 11762 15700
rect 12069 15691 12127 15697
rect 12069 15688 12081 15691
rect 11756 15660 12081 15688
rect 11756 15648 11762 15660
rect 12069 15657 12081 15660
rect 12115 15657 12127 15691
rect 12069 15651 12127 15657
rect 9582 15620 9588 15632
rect 7392 15592 8340 15620
rect 8404 15592 8800 15620
rect 9140 15592 9588 15620
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15552 6515 15555
rect 7006 15552 7012 15564
rect 6503 15524 7012 15552
rect 6503 15521 6515 15524
rect 6457 15515 6515 15521
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 7190 15512 7196 15564
rect 7248 15512 7254 15564
rect 7392 15561 7420 15592
rect 7377 15555 7435 15561
rect 7377 15521 7389 15555
rect 7423 15521 7435 15555
rect 7377 15515 7435 15521
rect 7650 15512 7656 15564
rect 7708 15512 7714 15564
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 7834 15552 7840 15564
rect 7791 15524 7840 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 7926 15512 7932 15564
rect 7984 15512 7990 15564
rect 8018 15512 8024 15564
rect 8076 15512 8082 15564
rect 8113 15555 8171 15561
rect 8113 15521 8125 15555
rect 8159 15552 8171 15555
rect 8202 15552 8208 15564
rect 8159 15524 8208 15552
rect 8159 15521 8171 15524
rect 8113 15515 8171 15521
rect 8202 15512 8208 15524
rect 8260 15512 8266 15564
rect 8312 15552 8340 15592
rect 8312 15524 8432 15552
rect 1213 15487 1271 15493
rect 1213 15453 1225 15487
rect 1259 15484 1271 15487
rect 2225 15487 2283 15493
rect 2225 15484 2237 15487
rect 1259 15456 2237 15484
rect 1259 15453 1271 15456
rect 1213 15447 1271 15453
rect 2225 15453 2237 15456
rect 2271 15484 2283 15487
rect 2314 15484 2320 15496
rect 2271 15456 2320 15484
rect 2271 15453 2283 15456
rect 2225 15447 2283 15453
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 3510 15444 3516 15496
rect 3568 15484 3574 15496
rect 3973 15487 4031 15493
rect 3973 15484 3985 15487
rect 3568 15456 3985 15484
rect 3568 15444 3574 15456
rect 3973 15453 3985 15456
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 7024 15484 7052 15512
rect 8036 15484 8064 15512
rect 7024 15456 8064 15484
rect 8404 15484 8432 15524
rect 8570 15512 8576 15564
rect 8628 15561 8634 15564
rect 8628 15555 8664 15561
rect 8652 15521 8664 15555
rect 8628 15515 8664 15521
rect 8628 15512 8634 15515
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 9140 15561 9168 15592
rect 9582 15580 9588 15592
rect 9640 15580 9646 15632
rect 9766 15580 9772 15632
rect 9824 15580 9830 15632
rect 10686 15620 10692 15632
rect 10152 15592 10692 15620
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8996 15524 9045 15552
rect 8996 15512 9002 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 9033 15515 9091 15521
rect 9125 15555 9183 15561
rect 9125 15521 9137 15555
rect 9171 15521 9183 15555
rect 9125 15515 9183 15521
rect 9217 15555 9275 15561
rect 9217 15521 9229 15555
rect 9263 15521 9275 15555
rect 9217 15515 9275 15521
rect 8754 15484 8760 15496
rect 8404 15456 8760 15484
rect 8754 15444 8760 15456
rect 8812 15484 8818 15496
rect 9232 15484 9260 15515
rect 9398 15512 9404 15564
rect 9456 15512 9462 15564
rect 8812 15456 9260 15484
rect 9585 15487 9643 15493
rect 8812 15444 8818 15456
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 9674 15484 9680 15496
rect 9631 15456 9680 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9674 15444 9680 15456
rect 9732 15444 9738 15496
rect 9784 15484 9812 15580
rect 10152 15561 10180 15592
rect 10686 15580 10692 15592
rect 10744 15620 10750 15632
rect 10965 15623 11023 15629
rect 10965 15620 10977 15623
rect 10744 15592 10977 15620
rect 10744 15580 10750 15592
rect 10965 15589 10977 15592
rect 11011 15620 11023 15623
rect 11164 15620 11192 15648
rect 11011 15592 12296 15620
rect 11011 15589 11023 15592
rect 10965 15583 11023 15589
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 11149 15555 11207 15561
rect 11149 15521 11161 15555
rect 11195 15521 11207 15555
rect 11149 15515 11207 15521
rect 9861 15487 9919 15493
rect 9861 15484 9873 15487
rect 9784 15456 9873 15484
rect 9861 15453 9873 15456
rect 9907 15453 9919 15487
rect 9861 15447 9919 15453
rect 2133 15419 2191 15425
rect 2133 15385 2145 15419
rect 2179 15416 2191 15419
rect 2406 15416 2412 15428
rect 2179 15388 2412 15416
rect 2179 15385 2191 15388
rect 2133 15379 2191 15385
rect 2406 15376 2412 15388
rect 2464 15376 2470 15428
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 7469 15419 7527 15425
rect 7469 15416 7481 15419
rect 5592 15388 7481 15416
rect 5592 15376 5598 15388
rect 7469 15385 7481 15388
rect 7515 15385 7527 15419
rect 7469 15379 7527 15385
rect 8297 15419 8355 15425
rect 8297 15385 8309 15419
rect 8343 15416 8355 15419
rect 8570 15416 8576 15428
rect 8343 15388 8576 15416
rect 8343 15385 8355 15388
rect 8297 15379 8355 15385
rect 8570 15376 8576 15388
rect 8628 15416 8634 15428
rect 8628 15388 9628 15416
rect 8628 15376 8634 15388
rect 9600 15360 9628 15388
rect 9876 15360 9904 15447
rect 9950 15444 9956 15496
rect 10008 15484 10014 15496
rect 10318 15484 10324 15496
rect 10008 15456 10324 15484
rect 10008 15444 10014 15456
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10226 15376 10232 15428
rect 10284 15416 10290 15428
rect 10962 15416 10968 15428
rect 10284 15388 10968 15416
rect 10284 15376 10290 15388
rect 10962 15376 10968 15388
rect 11020 15376 11026 15428
rect 11164 15416 11192 15515
rect 11514 15512 11520 15564
rect 11572 15552 11578 15564
rect 12268 15561 12296 15592
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 11572 15524 11621 15552
rect 11572 15512 11578 15524
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15521 12127 15555
rect 12069 15515 12127 15521
rect 12253 15555 12311 15561
rect 12253 15521 12265 15555
rect 12299 15521 12311 15555
rect 12253 15515 12311 15521
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15484 11759 15487
rect 11790 15484 11796 15496
rect 11747 15456 11796 15484
rect 11747 15453 11759 15456
rect 11701 15447 11759 15453
rect 11790 15444 11796 15456
rect 11848 15444 11854 15496
rect 12084 15484 12112 15515
rect 12342 15484 12348 15496
rect 11900 15456 12348 15484
rect 11606 15416 11612 15428
rect 11164 15388 11612 15416
rect 11606 15376 11612 15388
rect 11664 15416 11670 15428
rect 11900 15416 11928 15456
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 11664 15388 11928 15416
rect 11977 15419 12035 15425
rect 11664 15376 11670 15388
rect 11977 15385 11989 15419
rect 12023 15416 12035 15419
rect 12066 15416 12072 15428
rect 12023 15388 12072 15416
rect 12023 15385 12035 15388
rect 11977 15379 12035 15385
rect 12066 15376 12072 15388
rect 12124 15376 12130 15428
rect 1305 15351 1363 15357
rect 1305 15317 1317 15351
rect 1351 15348 1363 15351
rect 2038 15348 2044 15360
rect 1351 15320 2044 15348
rect 1351 15317 1363 15320
rect 1305 15311 1363 15317
rect 2038 15308 2044 15320
rect 2096 15308 2102 15360
rect 2317 15351 2375 15357
rect 2317 15317 2329 15351
rect 2363 15348 2375 15351
rect 2682 15348 2688 15360
rect 2363 15320 2688 15348
rect 2363 15317 2375 15320
rect 2317 15311 2375 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 2774 15308 2780 15360
rect 2832 15348 2838 15360
rect 2961 15351 3019 15357
rect 2961 15348 2973 15351
rect 2832 15320 2973 15348
rect 2832 15308 2838 15320
rect 2961 15317 2973 15320
rect 3007 15317 3019 15351
rect 2961 15311 3019 15317
rect 4522 15308 4528 15360
rect 4580 15348 4586 15360
rect 5077 15351 5135 15357
rect 5077 15348 5089 15351
rect 4580 15320 5089 15348
rect 4580 15308 4586 15320
rect 5077 15317 5089 15320
rect 5123 15317 5135 15351
rect 5077 15311 5135 15317
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 9398 15348 9404 15360
rect 7248 15320 9404 15348
rect 7248 15308 7254 15320
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 552 15258 12604 15280
rect 552 15206 3662 15258
rect 3714 15206 3726 15258
rect 3778 15206 3790 15258
rect 3842 15206 3854 15258
rect 3906 15206 3918 15258
rect 3970 15206 10062 15258
rect 10114 15206 10126 15258
rect 10178 15206 10190 15258
rect 10242 15206 10254 15258
rect 10306 15206 10318 15258
rect 10370 15206 12604 15258
rect 552 15184 12604 15206
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2096 15116 2268 15144
rect 2096 15104 2102 15116
rect 2240 15076 2268 15116
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 4249 15147 4307 15153
rect 4249 15144 4261 15147
rect 2464 15116 4261 15144
rect 2464 15104 2470 15116
rect 4249 15113 4261 15116
rect 4295 15113 4307 15147
rect 5534 15144 5540 15156
rect 4249 15107 4307 15113
rect 4356 15116 5540 15144
rect 3237 15079 3295 15085
rect 2240 15048 2636 15076
rect 2222 14968 2228 15020
rect 2280 14968 2286 15020
rect 2608 15008 2636 15048
rect 3237 15045 3249 15079
rect 3283 15076 3295 15079
rect 3418 15076 3424 15088
rect 3283 15048 3424 15076
rect 3283 15045 3295 15048
rect 3237 15039 3295 15045
rect 3418 15036 3424 15048
rect 3476 15036 3482 15088
rect 3881 15079 3939 15085
rect 3881 15045 3893 15079
rect 3927 15045 3939 15079
rect 4356 15076 4384 15116
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 5810 15104 5816 15156
rect 5868 15104 5874 15156
rect 8386 15144 8392 15156
rect 7484 15116 8392 15144
rect 3881 15039 3939 15045
rect 4080 15048 4384 15076
rect 4801 15079 4859 15085
rect 3896 15008 3924 15039
rect 2608 14980 3924 15008
rect 3142 14900 3148 14952
rect 3200 14940 3206 14952
rect 3513 14943 3571 14949
rect 3200 14912 3464 14940
rect 3200 14900 3206 14912
rect 1946 14832 1952 14884
rect 2004 14881 2010 14884
rect 2004 14872 2016 14881
rect 2004 14844 2049 14872
rect 2004 14835 2016 14844
rect 2004 14832 2010 14835
rect 2590 14832 2596 14884
rect 2648 14872 2654 14884
rect 3237 14875 3295 14881
rect 3237 14872 3249 14875
rect 2648 14844 3249 14872
rect 2648 14832 2654 14844
rect 3237 14841 3249 14844
rect 3283 14841 3295 14875
rect 3436 14872 3464 14912
rect 3513 14909 3525 14943
rect 3559 14940 3571 14943
rect 4080 14940 4108 15048
rect 4801 15045 4813 15079
rect 4847 15045 4859 15079
rect 4801 15039 4859 15045
rect 4816 15008 4844 15039
rect 5074 15036 5080 15088
rect 5132 15076 5138 15088
rect 5629 15079 5687 15085
rect 5629 15076 5641 15079
rect 5132 15048 5641 15076
rect 5132 15036 5138 15048
rect 5629 15045 5641 15048
rect 5675 15045 5687 15079
rect 5629 15039 5687 15045
rect 5828 15008 5856 15104
rect 6178 15036 6184 15088
rect 6236 15076 6242 15088
rect 7484 15076 7512 15116
rect 8386 15104 8392 15116
rect 8444 15104 8450 15156
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 9401 15147 9459 15153
rect 9401 15144 9413 15147
rect 8720 15116 9413 15144
rect 8720 15104 8726 15116
rect 9401 15113 9413 15116
rect 9447 15113 9459 15147
rect 11882 15144 11888 15156
rect 9401 15107 9459 15113
rect 9494 15116 11888 15144
rect 6236 15048 7512 15076
rect 6236 15036 6242 15048
rect 4264 14980 4844 15008
rect 5275 14980 5856 15008
rect 4264 14952 4292 14980
rect 3559 14912 4108 14940
rect 3559 14909 3571 14912
rect 3513 14903 3571 14909
rect 4154 14900 4160 14952
rect 4212 14900 4218 14952
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4522 14900 4528 14952
rect 4580 14900 4586 14952
rect 4614 14900 4620 14952
rect 4672 14940 4678 14952
rect 4672 14912 4936 14940
rect 4672 14900 4678 14912
rect 3881 14875 3939 14881
rect 3436 14844 3556 14872
rect 3237 14835 3295 14841
rect 845 14807 903 14813
rect 845 14804 857 14807
rect 492 14776 857 14804
rect 492 14532 520 14776
rect 845 14773 857 14776
rect 891 14773 903 14807
rect 845 14767 903 14773
rect 2774 14764 2780 14816
rect 2832 14804 2838 14816
rect 3421 14807 3479 14813
rect 3421 14804 3433 14807
rect 2832 14776 3433 14804
rect 2832 14764 2838 14776
rect 3421 14773 3433 14776
rect 3467 14773 3479 14807
rect 3528 14804 3556 14844
rect 3881 14841 3893 14875
rect 3927 14872 3939 14875
rect 4264 14872 4292 14900
rect 4798 14872 4804 14884
rect 3927 14844 4292 14872
rect 4448 14844 4804 14872
rect 3927 14841 3939 14844
rect 3881 14835 3939 14841
rect 4448 14813 4476 14844
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 4908 14872 4936 14912
rect 5074 14900 5080 14952
rect 5132 14900 5138 14952
rect 5275 14949 5303 14980
rect 6086 14968 6092 15020
rect 6144 14968 6150 15020
rect 6730 14968 6736 15020
rect 6788 15008 6794 15020
rect 7484 15017 7512 15048
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 9494 15076 9522 15116
rect 11882 15104 11888 15116
rect 11940 15104 11946 15156
rect 7708 15048 8708 15076
rect 7708 15036 7714 15048
rect 7469 15011 7527 15017
rect 6788 14980 7328 15008
rect 6788 14968 6794 14980
rect 7300 14952 7328 14980
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 7561 15011 7619 15017
rect 7561 14977 7573 15011
rect 7607 15008 7619 15011
rect 7834 15008 7840 15020
rect 7607 14980 7840 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 7834 14968 7840 14980
rect 7892 14968 7898 15020
rect 8386 14968 8392 15020
rect 8444 14968 8450 15020
rect 8680 15017 8708 15048
rect 9140 15048 9522 15076
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 5261 14943 5319 14949
rect 5261 14909 5273 14943
rect 5307 14909 5319 14943
rect 5261 14903 5319 14909
rect 5445 14943 5503 14949
rect 5445 14909 5457 14943
rect 5491 14940 5503 14943
rect 5534 14940 5540 14952
rect 5491 14912 5540 14940
rect 5491 14909 5503 14912
rect 5445 14903 5503 14909
rect 5460 14872 5488 14903
rect 5534 14900 5540 14912
rect 5592 14900 5598 14952
rect 5721 14943 5779 14949
rect 5721 14909 5733 14943
rect 5767 14909 5779 14943
rect 5721 14903 5779 14909
rect 6181 14943 6239 14949
rect 6181 14909 6193 14943
rect 6227 14940 6239 14943
rect 7190 14940 7196 14952
rect 6227 14912 7196 14940
rect 6227 14909 6239 14912
rect 6181 14903 6239 14909
rect 4908 14844 5488 14872
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3528 14776 4077 14804
rect 3421 14767 3479 14773
rect 4065 14773 4077 14776
rect 4111 14804 4123 14807
rect 4433 14807 4491 14813
rect 4433 14804 4445 14807
rect 4111 14776 4445 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 4433 14773 4445 14776
rect 4479 14773 4491 14807
rect 4433 14767 4491 14773
rect 4985 14807 5043 14813
rect 4985 14773 4997 14807
rect 5031 14804 5043 14807
rect 5074 14804 5080 14816
rect 5031 14776 5080 14804
rect 5031 14773 5043 14776
rect 4985 14767 5043 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 5736 14804 5764 14903
rect 7190 14900 7196 14912
rect 7248 14900 7254 14952
rect 7282 14900 7288 14952
rect 7340 14900 7346 14952
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14909 7435 14943
rect 7377 14903 7435 14909
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 9140 14940 9168 15048
rect 9858 15036 9864 15088
rect 9916 15076 9922 15088
rect 10505 15079 10563 15085
rect 9916 15048 10180 15076
rect 9916 15036 9922 15048
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9769 15011 9827 15017
rect 9272 14980 9628 15008
rect 9272 14968 9278 14980
rect 9600 14949 9628 14980
rect 9769 14977 9781 15011
rect 9815 15008 9827 15011
rect 9950 15008 9956 15020
rect 9815 14980 9956 15008
rect 9815 14977 9827 14980
rect 9769 14971 9827 14977
rect 9950 14968 9956 14980
rect 10008 14968 10014 15020
rect 10152 15017 10180 15048
rect 10505 15045 10517 15079
rect 10551 15076 10563 15079
rect 10686 15076 10692 15088
rect 10551 15048 10692 15076
rect 10551 15045 10563 15048
rect 10505 15039 10563 15045
rect 10686 15036 10692 15048
rect 10744 15036 10750 15088
rect 11790 15076 11796 15088
rect 11256 15048 11796 15076
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 14977 10195 15011
rect 10137 14971 10195 14977
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 10643 14980 10916 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 9140 14912 9321 14940
rect 8757 14903 8815 14909
rect 9309 14909 9321 14912
rect 9355 14909 9367 14943
rect 9309 14903 9367 14909
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 5902 14832 5908 14884
rect 5960 14872 5966 14884
rect 6638 14872 6644 14884
rect 5960 14844 6644 14872
rect 5960 14832 5966 14844
rect 6638 14832 6644 14844
rect 6696 14872 6702 14884
rect 7392 14872 7420 14903
rect 6696 14844 7420 14872
rect 7929 14875 7987 14881
rect 6696 14832 6702 14844
rect 7929 14841 7941 14875
rect 7975 14872 7987 14875
rect 8294 14872 8300 14884
rect 7975 14844 8300 14872
rect 7975 14841 7987 14844
rect 7929 14835 7987 14841
rect 8294 14832 8300 14844
rect 8352 14832 8358 14884
rect 5408 14776 5764 14804
rect 5408 14764 5414 14776
rect 6546 14764 6552 14816
rect 6604 14764 6610 14816
rect 6914 14764 6920 14816
rect 6972 14804 6978 14816
rect 7101 14807 7159 14813
rect 7101 14804 7113 14807
rect 6972 14776 7113 14804
rect 6972 14764 6978 14776
rect 7101 14773 7113 14776
rect 7147 14773 7159 14807
rect 7101 14767 7159 14773
rect 7834 14764 7840 14816
rect 7892 14804 7898 14816
rect 8772 14804 8800 14903
rect 9674 14900 9680 14952
rect 9732 14900 9738 14952
rect 9861 14943 9919 14949
rect 9861 14909 9873 14943
rect 9907 14909 9919 14943
rect 9861 14903 9919 14909
rect 9876 14872 9904 14903
rect 10042 14900 10048 14952
rect 10100 14900 10106 14952
rect 10888 14949 10916 14980
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11112 14980 11192 15008
rect 11112 14968 11118 14980
rect 11164 14949 11192 14980
rect 11256 14949 11284 15048
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 10873 14943 10931 14949
rect 10873 14909 10885 14943
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14909 11207 14943
rect 11149 14903 11207 14909
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 11330 14900 11336 14952
rect 11388 14900 11394 14952
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14940 12127 14943
rect 12342 14940 12348 14952
rect 12115 14912 12348 14940
rect 12115 14909 12127 14912
rect 12069 14903 12127 14909
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 11698 14872 11704 14884
rect 9876 14844 11704 14872
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 7892 14776 8800 14804
rect 7892 14764 7898 14776
rect 9122 14764 9128 14816
rect 9180 14764 9186 14816
rect 9766 14764 9772 14816
rect 9824 14804 9830 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 9824 14776 10701 14804
rect 9824 14764 9830 14776
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11146 14804 11152 14816
rect 11103 14776 11152 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11238 14764 11244 14816
rect 11296 14804 11302 14816
rect 11425 14807 11483 14813
rect 11425 14804 11437 14807
rect 11296 14776 11437 14804
rect 11296 14764 11302 14776
rect 11425 14773 11437 14776
rect 11471 14773 11483 14807
rect 11425 14767 11483 14773
rect 11606 14764 11612 14816
rect 11664 14804 11670 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11664 14776 11897 14804
rect 11664 14764 11670 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 11885 14767 11943 14773
rect 552 14714 12604 14736
rect 552 14662 4322 14714
rect 4374 14662 4386 14714
rect 4438 14662 4450 14714
rect 4502 14662 4514 14714
rect 4566 14662 4578 14714
rect 4630 14662 10722 14714
rect 10774 14662 10786 14714
rect 10838 14662 10850 14714
rect 10902 14662 10914 14714
rect 10966 14662 10978 14714
rect 11030 14662 12604 14714
rect 552 14640 12604 14662
rect 2866 14560 2872 14612
rect 2924 14600 2930 14612
rect 3142 14600 3148 14612
rect 2924 14572 3148 14600
rect 2924 14560 2930 14572
rect 3142 14560 3148 14572
rect 3200 14560 3206 14612
rect 4154 14560 4160 14612
rect 4212 14560 4218 14612
rect 4433 14603 4491 14609
rect 4433 14569 4445 14603
rect 4479 14600 4491 14603
rect 4798 14600 4804 14612
rect 4479 14572 4804 14600
rect 4479 14569 4491 14572
rect 4433 14563 4491 14569
rect 4798 14560 4804 14572
rect 4856 14560 4862 14612
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 4908 14572 5825 14600
rect 492 14504 1624 14532
rect 842 14424 848 14476
rect 900 14424 906 14476
rect 1305 14467 1363 14473
rect 1305 14433 1317 14467
rect 1351 14464 1363 14467
rect 1394 14464 1400 14476
rect 1351 14436 1400 14464
rect 1351 14433 1363 14436
rect 1305 14427 1363 14433
rect 1394 14424 1400 14436
rect 1452 14424 1458 14476
rect 1596 14473 1624 14504
rect 2332 14504 3832 14532
rect 1489 14467 1547 14473
rect 1489 14433 1501 14467
rect 1535 14433 1547 14467
rect 1489 14427 1547 14433
rect 1581 14467 1639 14473
rect 1581 14433 1593 14467
rect 1627 14433 1639 14467
rect 1581 14427 1639 14433
rect 1504 14328 1532 14427
rect 2130 14424 2136 14476
rect 2188 14424 2194 14476
rect 2332 14473 2360 14504
rect 2317 14467 2375 14473
rect 2317 14433 2329 14467
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 2682 14424 2688 14476
rect 2740 14424 2746 14476
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 3053 14467 3111 14473
rect 3053 14464 3065 14467
rect 2832 14436 3065 14464
rect 2832 14424 2838 14436
rect 3053 14433 3065 14436
rect 3099 14433 3111 14467
rect 3053 14427 3111 14433
rect 3145 14467 3203 14473
rect 3145 14433 3157 14467
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 1946 14356 1952 14408
rect 2004 14356 2010 14408
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 2409 14399 2467 14405
rect 2409 14396 2421 14399
rect 2280 14368 2421 14396
rect 2280 14356 2286 14368
rect 2409 14365 2421 14368
rect 2455 14396 2467 14399
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2455 14368 2973 14396
rect 2455 14365 2467 14368
rect 2409 14359 2467 14365
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 3160 14396 3188 14427
rect 3234 14424 3240 14476
rect 3292 14464 3298 14476
rect 3329 14467 3387 14473
rect 3329 14464 3341 14467
rect 3292 14436 3341 14464
rect 3292 14424 3298 14436
rect 3329 14433 3341 14436
rect 3375 14433 3387 14467
rect 3329 14427 3387 14433
rect 3418 14424 3424 14476
rect 3476 14424 3482 14476
rect 3602 14424 3608 14476
rect 3660 14424 3666 14476
rect 3694 14396 3700 14408
rect 3160 14368 3700 14396
rect 2961 14359 3019 14365
rect 3694 14356 3700 14368
rect 3752 14356 3758 14408
rect 3804 14396 3832 14504
rect 4172 14464 4200 14560
rect 4246 14492 4252 14544
rect 4304 14492 4310 14544
rect 4525 14467 4583 14473
rect 4172 14436 4476 14464
rect 4448 14396 4476 14436
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 4908 14464 4936 14572
rect 5813 14569 5825 14572
rect 5859 14569 5871 14603
rect 6086 14600 6092 14612
rect 5813 14563 5871 14569
rect 6013 14572 6092 14600
rect 4571 14436 4936 14464
rect 5261 14467 5319 14473
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5534 14464 5540 14476
rect 5307 14436 5540 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 3804 14368 4292 14396
rect 4448 14368 4905 14396
rect 1964 14328 1992 14356
rect 4264 14337 4292 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 5074 14356 5080 14408
rect 5132 14356 5138 14408
rect 5169 14399 5227 14405
rect 5169 14365 5181 14399
rect 5215 14365 5227 14399
rect 5169 14359 5227 14365
rect 2501 14331 2559 14337
rect 2501 14328 2513 14331
rect 1504 14300 2513 14328
rect 2501 14297 2513 14300
rect 2547 14297 2559 14331
rect 2501 14291 2559 14297
rect 2869 14331 2927 14337
rect 2869 14297 2881 14331
rect 2915 14328 2927 14331
rect 3421 14331 3479 14337
rect 3421 14328 3433 14331
rect 2915 14300 3433 14328
rect 2915 14297 2927 14300
rect 2869 14291 2927 14297
rect 3421 14297 3433 14300
rect 3467 14297 3479 14331
rect 3421 14291 3479 14297
rect 4249 14331 4307 14337
rect 4249 14297 4261 14331
rect 4295 14297 4307 14331
rect 4249 14291 4307 14297
rect 1762 14220 1768 14272
rect 1820 14260 1826 14272
rect 1949 14263 2007 14269
rect 1949 14260 1961 14263
rect 1820 14232 1961 14260
rect 1820 14220 1826 14232
rect 1949 14229 1961 14232
rect 1995 14229 2007 14263
rect 1949 14223 2007 14229
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 3329 14263 3387 14269
rect 3329 14260 3341 14263
rect 2648 14232 3341 14260
rect 2648 14220 2654 14232
rect 3329 14229 3341 14232
rect 3375 14260 3387 14263
rect 3602 14260 3608 14272
rect 3375 14232 3608 14260
rect 3375 14229 3387 14232
rect 3329 14223 3387 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3970 14220 3976 14272
rect 4028 14260 4034 14272
rect 4338 14260 4344 14272
rect 4028 14232 4344 14260
rect 4028 14220 4034 14232
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 5184 14260 5212 14359
rect 5350 14356 5356 14408
rect 5408 14356 5414 14408
rect 5460 14396 5488 14436
rect 5534 14424 5540 14436
rect 5592 14424 5598 14476
rect 6013 14473 6041 14572
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 6362 14560 6368 14612
rect 6420 14600 6426 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6420 14572 6469 14600
rect 6420 14560 6426 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 8478 14600 8484 14612
rect 6457 14563 6515 14569
rect 7392 14572 8484 14600
rect 6270 14492 6276 14544
rect 6328 14532 6334 14544
rect 6328 14504 6684 14532
rect 6328 14492 6334 14504
rect 6656 14473 6684 14504
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6090 14467 6148 14473
rect 6090 14433 6102 14467
rect 6136 14466 6148 14467
rect 6641 14467 6699 14473
rect 6136 14464 6224 14466
rect 6136 14438 6592 14464
rect 6136 14433 6148 14438
rect 6196 14436 6592 14438
rect 6090 14427 6148 14433
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5460 14368 6193 14396
rect 6181 14365 6193 14368
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6273 14399 6331 14405
rect 6273 14365 6285 14399
rect 6319 14365 6331 14399
rect 6564 14396 6592 14436
rect 6641 14433 6653 14467
rect 6687 14433 6699 14467
rect 6641 14427 6699 14433
rect 6914 14424 6920 14476
rect 6972 14424 6978 14476
rect 7392 14473 7420 14572
rect 8478 14560 8484 14572
rect 8536 14560 8542 14612
rect 9122 14560 9128 14612
rect 9180 14600 9186 14612
rect 9180 14572 9444 14600
rect 9180 14560 9186 14572
rect 8386 14532 8392 14544
rect 7484 14504 8392 14532
rect 7484 14473 7512 14504
rect 8386 14492 8392 14504
rect 8444 14492 8450 14544
rect 8938 14492 8944 14544
rect 8996 14532 9002 14544
rect 8996 14504 9260 14532
rect 8996 14492 9002 14504
rect 7377 14467 7435 14473
rect 7377 14433 7389 14467
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 7282 14396 7288 14408
rect 6564 14368 7288 14396
rect 6273 14359 6331 14365
rect 5368 14328 5396 14356
rect 6288 14328 6316 14359
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 5368 14300 6316 14328
rect 6730 14288 6736 14340
rect 6788 14288 6794 14340
rect 6822 14288 6828 14340
rect 6880 14288 6886 14340
rect 7392 14328 7420 14427
rect 7650 14424 7656 14476
rect 7708 14424 7714 14476
rect 8110 14424 8116 14476
rect 8168 14424 8174 14476
rect 8478 14424 8484 14476
rect 8536 14424 8542 14476
rect 9232 14473 9260 14504
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14433 8723 14467
rect 8665 14427 8723 14433
rect 9217 14467 9275 14473
rect 9217 14433 9229 14467
rect 9263 14433 9275 14467
rect 9217 14427 9275 14433
rect 7837 14399 7895 14405
rect 7837 14365 7849 14399
rect 7883 14396 7895 14399
rect 8297 14399 8355 14405
rect 8297 14396 8309 14399
rect 7883 14368 8309 14396
rect 7883 14365 7895 14368
rect 7837 14359 7895 14365
rect 8297 14365 8309 14368
rect 8343 14365 8355 14399
rect 8297 14359 8355 14365
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8680 14396 8708 14427
rect 8757 14399 8815 14405
rect 8757 14396 8769 14399
rect 8444 14368 8649 14396
rect 8680 14368 8769 14396
rect 8444 14356 8450 14368
rect 6932 14300 7420 14328
rect 5442 14260 5448 14272
rect 5184 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5718 14220 5724 14272
rect 5776 14260 5782 14272
rect 6932 14260 6960 14300
rect 7926 14288 7932 14340
rect 7984 14288 7990 14340
rect 8621 14328 8649 14368
rect 8757 14365 8769 14368
rect 8803 14365 8815 14399
rect 8757 14359 8815 14365
rect 8938 14356 8944 14408
rect 8996 14356 9002 14408
rect 9030 14356 9036 14408
rect 9088 14356 9094 14408
rect 9125 14399 9183 14405
rect 9125 14365 9137 14399
rect 9171 14396 9183 14399
rect 9306 14396 9312 14408
rect 9171 14368 9312 14396
rect 9171 14365 9183 14368
rect 9125 14359 9183 14365
rect 9306 14356 9312 14368
rect 9364 14356 9370 14408
rect 9416 14328 9444 14572
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 11609 14603 11667 14609
rect 11609 14600 11621 14603
rect 10100 14572 11621 14600
rect 10100 14560 10106 14572
rect 11609 14569 11621 14572
rect 11655 14569 11667 14603
rect 11609 14563 11667 14569
rect 9646 14504 10364 14532
rect 9490 14356 9496 14408
rect 9548 14396 9554 14408
rect 9646 14396 9674 14504
rect 9861 14467 9919 14473
rect 9861 14433 9873 14467
rect 9907 14464 9919 14467
rect 9950 14464 9956 14476
rect 9907 14436 9956 14464
rect 9907 14433 9919 14436
rect 9861 14427 9919 14433
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10336 14473 10364 14504
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10321 14467 10379 14473
rect 10321 14433 10333 14467
rect 10367 14433 10379 14467
rect 10321 14427 10379 14433
rect 9548 14368 9674 14396
rect 9548 14356 9554 14368
rect 9766 14356 9772 14408
rect 9824 14356 9830 14408
rect 10152 14396 10180 14427
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11149 14467 11207 14473
rect 11149 14464 11161 14467
rect 11112 14436 11161 14464
rect 11112 14424 11118 14436
rect 11149 14433 11161 14436
rect 11195 14433 11207 14467
rect 11793 14467 11851 14473
rect 11793 14464 11805 14467
rect 11149 14427 11207 14433
rect 11348 14436 11805 14464
rect 10502 14396 10508 14408
rect 10152 14368 10508 14396
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 11348 14328 11376 14436
rect 11793 14433 11805 14436
rect 11839 14433 11851 14467
rect 11793 14427 11851 14433
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 11977 14467 12035 14473
rect 11977 14464 11989 14467
rect 11940 14436 11989 14464
rect 11940 14424 11946 14436
rect 11977 14433 11989 14436
rect 12023 14433 12035 14467
rect 11977 14427 12035 14433
rect 12066 14424 12072 14476
rect 12124 14424 12130 14476
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 12084 14396 12112 14424
rect 11563 14368 12112 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 8621 14300 11376 14328
rect 5776 14232 6960 14260
rect 5776 14220 5782 14232
rect 7098 14220 7104 14272
rect 7156 14260 7162 14272
rect 8754 14260 8760 14272
rect 7156 14232 8760 14260
rect 7156 14220 7162 14232
rect 8754 14220 8760 14232
rect 8812 14260 8818 14272
rect 9030 14260 9036 14272
rect 8812 14232 9036 14260
rect 8812 14220 8818 14232
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 10321 14263 10379 14269
rect 10321 14229 10333 14263
rect 10367 14260 10379 14263
rect 10502 14260 10508 14272
rect 10367 14232 10508 14260
rect 10367 14229 10379 14232
rect 10321 14223 10379 14229
rect 10502 14220 10508 14232
rect 10560 14220 10566 14272
rect 10594 14220 10600 14272
rect 10652 14220 10658 14272
rect 552 14170 12604 14192
rect 552 14118 3662 14170
rect 3714 14118 3726 14170
rect 3778 14118 3790 14170
rect 3842 14118 3854 14170
rect 3906 14118 3918 14170
rect 3970 14118 10062 14170
rect 10114 14118 10126 14170
rect 10178 14118 10190 14170
rect 10242 14118 10254 14170
rect 10306 14118 10318 14170
rect 10370 14118 12604 14170
rect 552 14096 12604 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 1670 14056 1676 14068
rect 1627 14028 1676 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 1670 14016 1676 14028
rect 1728 14016 1734 14068
rect 2314 14016 2320 14068
rect 2372 14056 2378 14068
rect 2372 14028 2820 14056
rect 2372 14016 2378 14028
rect 1949 13991 2007 13997
rect 1949 13957 1961 13991
rect 1995 13988 2007 13991
rect 2685 13991 2743 13997
rect 2685 13988 2697 13991
rect 1995 13960 2697 13988
rect 1995 13957 2007 13960
rect 1949 13951 2007 13957
rect 2685 13957 2697 13960
rect 2731 13957 2743 13991
rect 2685 13951 2743 13957
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1670 13920 1676 13932
rect 1544 13892 1676 13920
rect 1544 13880 1550 13892
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2406 13920 2412 13932
rect 1780 13892 2412 13920
rect 1780 13861 1808 13892
rect 1765 13855 1823 13861
rect 1765 13821 1777 13855
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 2041 13855 2099 13861
rect 2041 13821 2053 13855
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 2056 13784 2084 13815
rect 2130 13812 2136 13864
rect 2188 13812 2194 13864
rect 2222 13812 2228 13864
rect 2280 13812 2286 13864
rect 2332 13861 2360 13892
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2792 13920 2820 14028
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5537 14059 5595 14065
rect 5537 14056 5549 14059
rect 5132 14028 5549 14056
rect 5132 14016 5138 14028
rect 5537 14025 5549 14028
rect 5583 14025 5595 14059
rect 5537 14019 5595 14025
rect 6086 14016 6092 14068
rect 6144 14016 6150 14068
rect 6822 14016 6828 14068
rect 6880 14016 6886 14068
rect 9766 14016 9772 14068
rect 9824 14056 9830 14068
rect 10137 14059 10195 14065
rect 9824 14028 9996 14056
rect 9824 14016 9830 14028
rect 4798 13948 4804 14000
rect 4856 13988 4862 14000
rect 5718 13988 5724 14000
rect 4856 13960 5724 13988
rect 4856 13948 4862 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 7926 13988 7932 14000
rect 6380 13960 7932 13988
rect 2639 13892 2820 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 2498 13812 2504 13864
rect 2556 13812 2562 13864
rect 2958 13812 2964 13864
rect 3016 13812 3022 13864
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 5040 13824 5181 13852
rect 5040 13812 5046 13824
rect 5169 13821 5181 13824
rect 5215 13821 5227 13855
rect 5169 13815 5227 13821
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 5721 13855 5779 13861
rect 5721 13852 5733 13855
rect 5684 13824 5733 13852
rect 5684 13812 5690 13824
rect 5721 13821 5733 13824
rect 5767 13852 5779 13855
rect 6380 13852 6408 13960
rect 7926 13948 7932 13960
rect 7984 13948 7990 14000
rect 9968 13997 9996 14028
rect 10137 14025 10149 14059
rect 10183 14056 10195 14059
rect 10594 14056 10600 14068
rect 10183 14028 10600 14056
rect 10183 14025 10195 14028
rect 10137 14019 10195 14025
rect 10594 14016 10600 14028
rect 10652 14016 10658 14068
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 12069 14059 12127 14065
rect 12069 14056 12081 14059
rect 11756 14028 12081 14056
rect 11756 14016 11762 14028
rect 12069 14025 12081 14028
rect 12115 14025 12127 14059
rect 12069 14019 12127 14025
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13957 10011 13991
rect 11793 13991 11851 13997
rect 11793 13988 11805 13991
rect 9953 13951 10011 13957
rect 10520 13960 11805 13988
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7558 13920 7564 13932
rect 6512 13892 7564 13920
rect 6512 13880 6518 13892
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 5767 13824 6408 13852
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 6546 13812 6552 13864
rect 6604 13812 6610 13864
rect 6638 13812 6644 13864
rect 6696 13852 6702 13864
rect 6825 13855 6883 13861
rect 6825 13852 6837 13855
rect 6696 13824 6837 13852
rect 6696 13812 6702 13824
rect 6825 13821 6837 13824
rect 6871 13821 6883 13855
rect 6825 13815 6883 13821
rect 9858 13812 9864 13864
rect 9916 13852 9922 13864
rect 10520 13861 10548 13960
rect 11793 13957 11805 13960
rect 11839 13957 11851 13991
rect 11793 13951 11851 13957
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 10505 13855 10563 13861
rect 9916 13824 10456 13852
rect 9916 13812 9922 13824
rect 2240 13784 2268 13812
rect 2056 13756 2268 13784
rect 2590 13744 2596 13796
rect 2648 13784 2654 13796
rect 2685 13787 2743 13793
rect 2685 13784 2697 13787
rect 2648 13756 2697 13784
rect 2648 13744 2654 13756
rect 2685 13753 2697 13756
rect 2731 13753 2743 13787
rect 2685 13747 2743 13753
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13784 2927 13787
rect 3234 13784 3240 13796
rect 2915 13756 3240 13784
rect 2915 13753 2927 13756
rect 2869 13747 2927 13753
rect 2406 13676 2412 13728
rect 2464 13716 2470 13728
rect 2884 13716 2912 13747
rect 3234 13744 3240 13756
rect 3292 13744 3298 13796
rect 3418 13744 3424 13796
rect 3476 13784 3482 13796
rect 4338 13784 4344 13796
rect 3476 13756 4344 13784
rect 3476 13744 3482 13756
rect 4338 13744 4344 13756
rect 4396 13784 4402 13796
rect 5353 13787 5411 13793
rect 5353 13784 5365 13787
rect 4396 13756 5365 13784
rect 4396 13744 4402 13756
rect 5353 13753 5365 13756
rect 5399 13784 5411 13787
rect 5905 13787 5963 13793
rect 5905 13784 5917 13787
rect 5399 13756 5917 13784
rect 5399 13753 5411 13756
rect 5353 13747 5411 13753
rect 5905 13753 5917 13756
rect 5951 13784 5963 13787
rect 7374 13784 7380 13796
rect 5951 13756 7380 13784
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 7374 13744 7380 13756
rect 7432 13784 7438 13796
rect 8938 13784 8944 13796
rect 7432 13756 8944 13784
rect 7432 13744 7438 13756
rect 8938 13744 8944 13756
rect 8996 13784 9002 13796
rect 9398 13784 9404 13796
rect 8996 13756 9404 13784
rect 8996 13744 9002 13756
rect 9398 13744 9404 13756
rect 9456 13744 9462 13796
rect 9677 13787 9735 13793
rect 9677 13753 9689 13787
rect 9723 13784 9735 13787
rect 9950 13784 9956 13796
rect 9723 13756 9956 13784
rect 9723 13753 9735 13756
rect 9677 13747 9735 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10428 13784 10456 13824
rect 10505 13821 10517 13855
rect 10551 13821 10563 13855
rect 10505 13815 10563 13821
rect 10594 13812 10600 13864
rect 10652 13852 10658 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10652 13824 10701 13852
rect 10652 13812 10658 13824
rect 10689 13821 10701 13824
rect 10735 13852 10747 13855
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10735 13824 10793 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13821 10931 13855
rect 11072 13852 11100 13880
rect 10873 13815 10931 13821
rect 10980 13824 11100 13852
rect 11149 13855 11207 13861
rect 10888 13784 10916 13815
rect 10428 13756 10916 13784
rect 2464 13688 2912 13716
rect 2464 13676 2470 13688
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6641 13719 6699 13725
rect 6641 13716 6653 13719
rect 6420 13688 6653 13716
rect 6420 13676 6426 13688
rect 6641 13685 6653 13688
rect 6687 13716 6699 13719
rect 6822 13716 6828 13728
rect 6687 13688 6828 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 10689 13719 10747 13725
rect 10689 13685 10701 13719
rect 10735 13716 10747 13719
rect 10980 13716 11008 13824
rect 11149 13821 11161 13855
rect 11195 13852 11207 13855
rect 11238 13852 11244 13864
rect 11195 13824 11244 13852
rect 11195 13821 11207 13824
rect 11149 13815 11207 13821
rect 11238 13812 11244 13824
rect 11296 13812 11302 13864
rect 11514 13812 11520 13864
rect 11572 13852 11578 13864
rect 11882 13852 11888 13864
rect 11572 13824 11888 13852
rect 11572 13812 11578 13824
rect 11882 13812 11888 13824
rect 11940 13812 11946 13864
rect 12066 13812 12072 13864
rect 12124 13812 12130 13864
rect 11425 13787 11483 13793
rect 11425 13753 11437 13787
rect 11471 13753 11483 13787
rect 11425 13747 11483 13753
rect 10735 13688 11008 13716
rect 10735 13685 10747 13688
rect 10689 13679 10747 13685
rect 11146 13676 11152 13728
rect 11204 13716 11210 13728
rect 11440 13716 11468 13747
rect 11606 13744 11612 13796
rect 11664 13744 11670 13796
rect 11204 13688 11468 13716
rect 11204 13676 11210 13688
rect 552 13626 12604 13648
rect 552 13574 4322 13626
rect 4374 13574 4386 13626
rect 4438 13574 4450 13626
rect 4502 13574 4514 13626
rect 4566 13574 4578 13626
rect 4630 13574 10722 13626
rect 10774 13574 10786 13626
rect 10838 13574 10850 13626
rect 10902 13574 10914 13626
rect 10966 13574 10978 13626
rect 11030 13574 12604 13626
rect 552 13552 12604 13574
rect 2406 13472 2412 13524
rect 2464 13472 2470 13524
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 2958 13512 2964 13524
rect 2823 13484 2964 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 6362 13472 6368 13524
rect 6420 13512 6426 13524
rect 6549 13515 6607 13521
rect 6549 13512 6561 13515
rect 6420 13484 6561 13512
rect 6420 13472 6426 13484
rect 6549 13481 6561 13484
rect 6595 13481 6607 13515
rect 6549 13475 6607 13481
rect 6730 13472 6736 13524
rect 6788 13512 6794 13524
rect 7558 13512 7564 13524
rect 6788 13484 7564 13512
rect 6788 13472 6794 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 8941 13515 8999 13521
rect 8941 13481 8953 13515
rect 8987 13512 8999 13515
rect 9214 13512 9220 13524
rect 8987 13484 9220 13512
rect 8987 13481 8999 13484
rect 8941 13475 8999 13481
rect 2590 13404 2596 13456
rect 2648 13404 2654 13456
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 8570 13444 8576 13456
rect 7340 13416 8576 13444
rect 7340 13404 7346 13416
rect 8570 13404 8576 13416
rect 8628 13404 8634 13456
rect 8956 13444 8984 13475
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 10594 13472 10600 13524
rect 10652 13512 10658 13524
rect 10965 13515 11023 13521
rect 10965 13512 10977 13515
rect 10652 13484 10977 13512
rect 10652 13472 10658 13484
rect 10965 13481 10977 13484
rect 11011 13481 11023 13515
rect 10965 13475 11023 13481
rect 11606 13444 11612 13456
rect 8680 13416 8984 13444
rect 10980 13416 11612 13444
rect 1946 13336 1952 13388
rect 2004 13385 2010 13388
rect 2004 13376 2016 13385
rect 2004 13348 2049 13376
rect 2004 13339 2016 13348
rect 2004 13336 2010 13339
rect 2314 13336 2320 13388
rect 2372 13336 2378 13388
rect 2685 13379 2743 13385
rect 2685 13345 2697 13379
rect 2731 13376 2743 13379
rect 2774 13376 2780 13388
rect 2731 13348 2780 13376
rect 2731 13345 2743 13348
rect 2685 13339 2743 13345
rect 2774 13336 2780 13348
rect 2832 13336 2838 13388
rect 2869 13379 2927 13385
rect 2869 13345 2881 13379
rect 2915 13376 2927 13379
rect 3234 13376 3240 13388
rect 2915 13348 3240 13376
rect 2915 13345 2927 13348
rect 2869 13339 2927 13345
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 3789 13379 3847 13385
rect 3789 13345 3801 13379
rect 3835 13376 3847 13379
rect 4614 13376 4620 13388
rect 3835 13348 4620 13376
rect 3835 13345 3847 13348
rect 3789 13339 3847 13345
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 4798 13336 4804 13388
rect 4856 13336 4862 13388
rect 5534 13336 5540 13388
rect 5592 13376 5598 13388
rect 6457 13379 6515 13385
rect 6457 13376 6469 13379
rect 5592 13348 6469 13376
rect 5592 13336 5598 13348
rect 6457 13345 6469 13348
rect 6503 13345 6515 13379
rect 6457 13339 6515 13345
rect 6638 13336 6644 13388
rect 6696 13376 6702 13388
rect 6733 13379 6791 13385
rect 6733 13376 6745 13379
rect 6696 13348 6745 13376
rect 6696 13336 6702 13348
rect 6733 13345 6745 13348
rect 6779 13345 6791 13379
rect 6733 13339 6791 13345
rect 7098 13336 7104 13388
rect 7156 13376 7162 13388
rect 8680 13376 8708 13416
rect 7156 13348 8708 13376
rect 8849 13379 8907 13385
rect 7156 13336 7162 13348
rect 8849 13345 8861 13379
rect 8895 13345 8907 13379
rect 8849 13339 8907 13345
rect 9125 13379 9183 13385
rect 9125 13345 9137 13379
rect 9171 13376 9183 13379
rect 9398 13376 9404 13388
rect 9171 13348 9404 13376
rect 9171 13345 9183 13348
rect 9125 13339 9183 13345
rect 2222 13268 2228 13320
rect 2280 13268 2286 13320
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 4062 13308 4068 13320
rect 3927 13280 4068 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 4062 13268 4068 13280
rect 4120 13268 4126 13320
rect 8864 13308 8892 13339
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 10594 13336 10600 13388
rect 10652 13376 10658 13388
rect 10980 13385 11008 13416
rect 11606 13404 11612 13416
rect 11664 13404 11670 13456
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10652 13348 10977 13376
rect 10652 13336 10658 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11146 13336 11152 13388
rect 11204 13336 11210 13388
rect 9306 13308 9312 13320
rect 8864 13280 9312 13308
rect 9306 13268 9312 13280
rect 9364 13268 9370 13320
rect 2498 13200 2504 13252
rect 2556 13240 2562 13252
rect 2593 13243 2651 13249
rect 2593 13240 2605 13243
rect 2556 13212 2605 13240
rect 2556 13200 2562 13212
rect 2593 13209 2605 13212
rect 2639 13209 2651 13243
rect 2593 13203 2651 13209
rect 845 13175 903 13181
rect 845 13172 857 13175
rect 492 13144 857 13172
rect 492 12832 520 13144
rect 845 13141 857 13144
rect 891 13141 903 13175
rect 845 13135 903 13141
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4430 13172 4436 13184
rect 4203 13144 4436 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4430 13132 4436 13144
rect 4488 13132 4494 13184
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 4890 13172 4896 13184
rect 4663 13144 4896 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7282 13172 7288 13184
rect 6963 13144 7288 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7282 13132 7288 13144
rect 7340 13132 7346 13184
rect 8110 13132 8116 13184
rect 8168 13172 8174 13184
rect 9125 13175 9183 13181
rect 9125 13172 9137 13175
rect 8168 13144 9137 13172
rect 8168 13132 8174 13144
rect 9125 13141 9137 13144
rect 9171 13141 9183 13175
rect 9125 13135 9183 13141
rect 552 13082 12604 13104
rect 552 13030 3662 13082
rect 3714 13030 3726 13082
rect 3778 13030 3790 13082
rect 3842 13030 3854 13082
rect 3906 13030 3918 13082
rect 3970 13030 10062 13082
rect 10114 13030 10126 13082
rect 10178 13030 10190 13082
rect 10242 13030 10254 13082
rect 10306 13030 10318 13082
rect 10370 13030 12604 13082
rect 552 13008 12604 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 2593 12971 2651 12977
rect 2593 12968 2605 12971
rect 2372 12940 2605 12968
rect 2372 12928 2378 12940
rect 2593 12937 2605 12940
rect 2639 12937 2651 12971
rect 2593 12931 2651 12937
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 6273 12971 6331 12977
rect 6273 12968 6285 12971
rect 3292 12940 6285 12968
rect 3292 12928 3298 12940
rect 6273 12937 6285 12940
rect 6319 12937 6331 12971
rect 6273 12931 6331 12937
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 7742 12968 7748 12980
rect 6604 12940 7748 12968
rect 6604 12928 6610 12940
rect 7742 12928 7748 12940
rect 7800 12968 7806 12980
rect 7926 12968 7932 12980
rect 7800 12940 7932 12968
rect 7800 12928 7806 12940
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9398 12928 9404 12980
rect 9456 12928 9462 12980
rect 9950 12928 9956 12980
rect 10008 12928 10014 12980
rect 2774 12900 2780 12912
rect 2746 12860 2780 12900
rect 2832 12860 2838 12912
rect 5166 12860 5172 12912
rect 5224 12860 5230 12912
rect 5534 12860 5540 12912
rect 5592 12860 5598 12912
rect 6181 12903 6239 12909
rect 5736 12872 6040 12900
rect 1581 12835 1639 12841
rect 1581 12832 1593 12835
rect 492 12804 1593 12832
rect 1581 12801 1593 12804
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2746 12832 2774 12860
rect 2547 12804 2774 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 5184 12832 5212 12860
rect 5261 12835 5319 12841
rect 5261 12832 5273 12835
rect 4672 12804 5028 12832
rect 5184 12804 5273 12832
rect 4672 12792 4678 12804
rect 1305 12767 1363 12773
rect 1305 12733 1317 12767
rect 1351 12764 1363 12767
rect 1394 12764 1400 12776
rect 1351 12736 1400 12764
rect 1351 12733 1363 12736
rect 1305 12727 1363 12733
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 1489 12767 1547 12773
rect 1489 12733 1501 12767
rect 1535 12764 1547 12767
rect 2038 12764 2044 12776
rect 1535 12736 2044 12764
rect 1535 12733 1547 12736
rect 1489 12727 1547 12733
rect 2038 12724 2044 12736
rect 2096 12724 2102 12776
rect 2682 12724 2688 12776
rect 2740 12724 2746 12776
rect 2774 12724 2780 12776
rect 2832 12724 2838 12776
rect 4154 12724 4160 12776
rect 4212 12724 4218 12776
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4304 12736 4353 12764
rect 4304 12724 4310 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 4341 12727 4399 12733
rect 4430 12724 4436 12776
rect 4488 12724 4494 12776
rect 4525 12767 4583 12773
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 4890 12764 4896 12776
rect 4571 12736 4896 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 842 12656 848 12708
rect 900 12656 906 12708
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 4540 12696 4568 12727
rect 4890 12724 4896 12736
rect 4948 12724 4954 12776
rect 5000 12764 5028 12804
rect 5261 12801 5273 12804
rect 5307 12801 5319 12835
rect 5261 12795 5319 12801
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 5000 12736 5181 12764
rect 5169 12733 5181 12736
rect 5215 12764 5227 12767
rect 5626 12764 5632 12776
rect 5215 12736 5632 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 5626 12724 5632 12736
rect 5684 12764 5690 12776
rect 5736 12764 5764 12872
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12801 5963 12835
rect 6012 12832 6040 12872
rect 6181 12869 6193 12903
rect 6227 12900 6239 12903
rect 6822 12900 6828 12912
rect 6227 12872 6828 12900
rect 6227 12869 6239 12872
rect 6181 12863 6239 12869
rect 6822 12860 6828 12872
rect 6880 12860 6886 12912
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 7607 12872 8493 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8481 12869 8493 12872
rect 8527 12869 8539 12903
rect 8481 12863 8539 12869
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 9732 12872 10456 12900
rect 9732 12860 9738 12872
rect 10428 12844 10456 12872
rect 11974 12860 11980 12912
rect 12032 12860 12038 12912
rect 7285 12835 7343 12841
rect 6012 12804 7236 12832
rect 5905 12795 5963 12801
rect 5684 12736 5764 12764
rect 5813 12767 5871 12773
rect 5684 12724 5690 12736
rect 5813 12733 5825 12767
rect 5859 12733 5871 12767
rect 5920 12764 5948 12795
rect 7208 12776 7236 12804
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7466 12832 7472 12844
rect 7331 12804 7472 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7653 12835 7711 12841
rect 7653 12801 7665 12835
rect 7699 12832 7711 12835
rect 7742 12832 7748 12844
rect 7699 12804 7748 12832
rect 7699 12801 7711 12804
rect 7653 12795 7711 12801
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 7944 12804 8524 12832
rect 6454 12764 6460 12776
rect 5920 12736 6460 12764
rect 5813 12727 5871 12733
rect 4028 12668 4568 12696
rect 4028 12656 4034 12668
rect 4798 12588 4804 12640
rect 4856 12588 4862 12640
rect 5828 12628 5856 12727
rect 6454 12724 6460 12736
rect 6512 12724 6518 12776
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 6733 12767 6791 12773
rect 6733 12733 6745 12767
rect 6779 12733 6791 12767
rect 6733 12727 6791 12733
rect 6825 12767 6883 12773
rect 6825 12733 6837 12767
rect 6871 12764 6883 12767
rect 7006 12764 7012 12776
rect 6871 12736 7012 12764
rect 6871 12733 6883 12736
rect 6825 12727 6883 12733
rect 6748 12696 6776 12727
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7190 12724 7196 12776
rect 7248 12724 7254 12776
rect 7484 12764 7512 12792
rect 7944 12776 7972 12804
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7484 12736 7849 12764
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 7926 12724 7932 12776
rect 7984 12724 7990 12776
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 6914 12696 6920 12708
rect 6748 12668 6920 12696
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7024 12696 7052 12724
rect 8220 12696 8248 12727
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 8352 12736 8401 12764
rect 8352 12724 8358 12736
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8496 12764 8524 12804
rect 8662 12792 8668 12844
rect 8720 12792 8726 12844
rect 9490 12792 9496 12844
rect 9548 12832 9554 12844
rect 9585 12835 9643 12841
rect 9585 12832 9597 12835
rect 9548 12804 9597 12832
rect 9548 12792 9554 12804
rect 9585 12801 9597 12804
rect 9631 12801 9643 12835
rect 9585 12795 9643 12801
rect 10410 12792 10416 12844
rect 10468 12792 10474 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 8938 12773 8944 12776
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8496 12736 8769 12764
rect 8389 12727 8447 12733
rect 8757 12733 8769 12736
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 8905 12767 8944 12773
rect 8905 12733 8917 12767
rect 8905 12727 8944 12733
rect 8938 12724 8944 12727
rect 8996 12724 9002 12776
rect 9122 12724 9128 12776
rect 9180 12724 9186 12776
rect 9263 12767 9321 12773
rect 9263 12733 9275 12767
rect 9309 12764 9321 12767
rect 9508 12764 9536 12792
rect 9309 12736 9536 12764
rect 9677 12767 9735 12773
rect 9309 12733 9321 12736
rect 9263 12727 9321 12733
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 11238 12764 11244 12776
rect 9723 12736 11244 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11606 12724 11612 12776
rect 11664 12724 11670 12776
rect 7024 12668 8248 12696
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12696 8723 12699
rect 9033 12699 9091 12705
rect 9033 12696 9045 12699
rect 8711 12668 9045 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 9033 12665 9045 12668
rect 9079 12665 9091 12699
rect 9033 12659 9091 12665
rect 7834 12628 7840 12640
rect 5828 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12628 7898 12640
rect 8938 12628 8944 12640
rect 7892 12600 8944 12628
rect 7892 12588 7898 12600
rect 8938 12588 8944 12600
rect 8996 12588 9002 12640
rect 9140 12628 9168 12724
rect 9766 12628 9772 12640
rect 9140 12600 9772 12628
rect 9766 12588 9772 12600
rect 9824 12588 9830 12640
rect 552 12538 12604 12560
rect 552 12486 4322 12538
rect 4374 12486 4386 12538
rect 4438 12486 4450 12538
rect 4502 12486 4514 12538
rect 4566 12486 4578 12538
rect 4630 12486 10722 12538
rect 10774 12486 10786 12538
rect 10838 12486 10850 12538
rect 10902 12486 10914 12538
rect 10966 12486 10978 12538
rect 11030 12486 12604 12538
rect 552 12464 12604 12486
rect 474 12384 480 12436
rect 532 12424 538 12436
rect 750 12424 756 12436
rect 532 12396 756 12424
rect 532 12384 538 12396
rect 750 12384 756 12396
rect 808 12384 814 12436
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 2866 12424 2872 12436
rect 2740 12396 2872 12424
rect 2740 12384 2746 12396
rect 2866 12384 2872 12396
rect 2924 12384 2930 12436
rect 3050 12384 3056 12436
rect 3108 12384 3114 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 4580 12396 4629 12424
rect 4580 12384 4586 12396
rect 4617 12393 4629 12396
rect 4663 12393 4675 12427
rect 4617 12387 4675 12393
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5997 12427 6055 12433
rect 4764 12396 5488 12424
rect 4764 12384 4770 12396
rect 1394 12316 1400 12368
rect 1452 12316 1458 12368
rect 1578 12316 1584 12368
rect 1636 12356 1642 12368
rect 3418 12356 3424 12368
rect 1636 12328 2084 12356
rect 1636 12316 1642 12328
rect 382 12248 388 12300
rect 440 12288 446 12300
rect 2056 12297 2084 12328
rect 3068 12328 3424 12356
rect 1213 12291 1271 12297
rect 1213 12288 1225 12291
rect 440 12260 1225 12288
rect 440 12248 446 12260
rect 1213 12257 1225 12260
rect 1259 12257 1271 12291
rect 1857 12291 1915 12297
rect 1857 12288 1869 12291
rect 1213 12251 1271 12257
rect 1412 12260 1869 12288
rect 1412 12232 1440 12260
rect 1857 12257 1869 12260
rect 1903 12257 1915 12291
rect 1857 12251 1915 12257
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 2823 12260 3004 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 1394 12180 1400 12232
rect 1452 12180 1458 12232
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2682 12220 2688 12232
rect 2179 12192 2688 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2682 12180 2688 12192
rect 2740 12180 2746 12232
rect 2976 12152 3004 12260
rect 3068 12229 3096 12328
rect 3418 12316 3424 12328
rect 3476 12316 3482 12368
rect 3896 12328 5396 12356
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3896 12288 3924 12328
rect 4356 12300 4384 12328
rect 3375 12260 3924 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4065 12291 4123 12297
rect 4065 12288 4077 12291
rect 4028 12260 4077 12288
rect 4028 12248 4034 12260
rect 4065 12257 4077 12260
rect 4111 12257 4123 12291
rect 4065 12251 4123 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12257 4215 12291
rect 4157 12251 4215 12257
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3142 12180 3148 12232
rect 3200 12220 3206 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3200 12192 3249 12220
rect 3200 12180 3206 12192
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3697 12223 3755 12229
rect 3697 12189 3709 12223
rect 3743 12220 3755 12223
rect 4172 12220 4200 12251
rect 4246 12248 4252 12300
rect 4304 12248 4310 12300
rect 4338 12248 4344 12300
rect 4396 12248 4402 12300
rect 4430 12248 4436 12300
rect 4488 12248 4494 12300
rect 5000 12297 5028 12328
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 4525 12251 4583 12257
rect 4709 12291 4767 12297
rect 4709 12257 4721 12291
rect 4755 12257 4767 12291
rect 4709 12251 4767 12257
rect 4985 12291 5043 12297
rect 4985 12257 4997 12291
rect 5031 12257 5043 12291
rect 4985 12251 5043 12257
rect 3743 12192 4200 12220
rect 3743 12189 3755 12192
rect 3697 12183 3755 12189
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 2976 12124 3801 12152
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4540 12152 4568 12251
rect 4724 12220 4752 12251
rect 5166 12248 5172 12300
rect 5224 12248 5230 12300
rect 4890 12220 4896 12232
rect 4724 12192 4896 12220
rect 4890 12180 4896 12192
rect 4948 12180 4954 12232
rect 5077 12223 5135 12229
rect 5077 12189 5089 12223
rect 5123 12220 5135 12223
rect 5184 12220 5212 12248
rect 5123 12192 5212 12220
rect 5368 12220 5396 12328
rect 5460 12300 5488 12396
rect 5997 12393 6009 12427
rect 6043 12424 6055 12427
rect 6638 12424 6644 12436
rect 6043 12396 6644 12424
rect 6043 12393 6055 12396
rect 5997 12387 6055 12393
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 8202 12424 8208 12436
rect 6748 12396 8208 12424
rect 6748 12356 6776 12396
rect 8202 12384 8208 12396
rect 8260 12424 8266 12436
rect 8260 12396 8340 12424
rect 8260 12384 8266 12396
rect 6472 12328 6776 12356
rect 5442 12248 5448 12300
rect 5500 12248 5506 12300
rect 5626 12248 5632 12300
rect 5684 12248 5690 12300
rect 6181 12291 6239 12297
rect 6181 12257 6193 12291
rect 6227 12257 6239 12291
rect 6181 12251 6239 12257
rect 5644 12220 5672 12248
rect 5368 12192 5672 12220
rect 5123 12189 5135 12192
rect 5077 12183 5135 12189
rect 5537 12155 5595 12161
rect 5537 12152 5549 12155
rect 4212 12124 4568 12152
rect 4632 12124 5549 12152
rect 4212 12112 4218 12124
rect 4632 12096 4660 12124
rect 5537 12121 5549 12124
rect 5583 12121 5595 12155
rect 6196 12152 6224 12251
rect 6362 12248 6368 12300
rect 6420 12248 6426 12300
rect 6472 12297 6500 12328
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 7064 12328 7328 12356
rect 7064 12316 7070 12328
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12257 6515 12291
rect 6457 12251 6515 12257
rect 6549 12291 6607 12297
rect 6549 12257 6561 12291
rect 6595 12257 6607 12291
rect 6549 12251 6607 12257
rect 6380 12220 6408 12248
rect 6564 12220 6592 12251
rect 6730 12248 6736 12300
rect 6788 12248 6794 12300
rect 6822 12248 6828 12300
rect 6880 12248 6886 12300
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 7300 12297 7328 12328
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 7926 12356 7932 12368
rect 7524 12328 7604 12356
rect 7524 12316 7530 12328
rect 7576 12297 7604 12328
rect 7852 12328 7932 12356
rect 7285 12291 7343 12297
rect 7285 12257 7297 12291
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7650 12248 7656 12300
rect 7708 12248 7714 12300
rect 7852 12297 7880 12328
rect 7926 12316 7932 12328
rect 7984 12316 7990 12368
rect 7837 12291 7895 12297
rect 7837 12257 7849 12291
rect 7883 12257 7895 12291
rect 7837 12251 7895 12257
rect 8021 12291 8079 12297
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8110 12288 8116 12300
rect 8067 12260 8116 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8312 12288 8340 12396
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9732 12396 11284 12424
rect 9732 12384 9738 12396
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 8996 12328 9536 12356
rect 8996 12316 9002 12328
rect 8251 12260 8340 12288
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 8386 12248 8392 12300
rect 8444 12248 8450 12300
rect 8846 12248 8852 12300
rect 8904 12288 8910 12300
rect 9508 12297 9536 12328
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 10410 12356 10416 12368
rect 9916 12328 10416 12356
rect 9916 12316 9922 12328
rect 9493 12291 9551 12297
rect 8904 12260 9444 12288
rect 8904 12248 8910 12260
rect 7116 12220 7144 12248
rect 6380 12192 6592 12220
rect 6656 12192 7144 12220
rect 7929 12223 7987 12229
rect 6270 12152 6276 12164
rect 6196 12124 6276 12152
rect 5537 12115 5595 12121
rect 6270 12112 6276 12124
rect 6328 12152 6334 12164
rect 6656 12152 6684 12192
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 6328 12124 6684 12152
rect 6328 12112 6334 12124
rect 7282 12112 7288 12164
rect 7340 12152 7346 12164
rect 7944 12152 7972 12183
rect 8404 12152 8432 12248
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9122 12180 9128 12232
rect 9180 12180 9186 12232
rect 9416 12229 9444 12260
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 9953 12291 10011 12297
rect 9953 12288 9965 12291
rect 9493 12251 9551 12257
rect 9876 12260 9965 12288
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9674 12152 9680 12164
rect 7340 12124 9680 12152
rect 7340 12112 7346 12124
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 9876 12161 9904 12260
rect 9953 12257 9965 12260
rect 9999 12257 10011 12291
rect 9953 12251 10011 12257
rect 10042 12248 10048 12300
rect 10100 12248 10106 12300
rect 10244 12297 10272 12328
rect 10410 12316 10416 12328
rect 10468 12316 10474 12368
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 10229 12251 10287 12257
rect 10778 12248 10784 12300
rect 10836 12288 10842 12300
rect 10962 12288 10968 12300
rect 10836 12260 10968 12288
rect 10836 12248 10842 12260
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11146 12248 11152 12300
rect 11204 12248 11210 12300
rect 11256 12220 11284 12396
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11664 12396 11805 12424
rect 11664 12384 11670 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 11808 12356 11836 12387
rect 11808 12328 12204 12356
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12257 11483 12291
rect 11425 12251 11483 12257
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 10980 12192 11345 12220
rect 10980 12164 11008 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 9861 12155 9919 12161
rect 9861 12121 9873 12155
rect 9907 12121 9919 12155
rect 9861 12115 9919 12121
rect 10962 12112 10968 12164
rect 11020 12112 11026 12164
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11440 12152 11468 12251
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 12176 12297 12204 12328
rect 12069 12291 12127 12297
rect 12069 12288 12081 12291
rect 11756 12260 12081 12288
rect 11756 12248 11762 12260
rect 12069 12257 12081 12260
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 11882 12180 11888 12232
rect 11940 12180 11946 12232
rect 11606 12152 11612 12164
rect 11296 12124 11612 12152
rect 11296 12112 11302 12124
rect 11606 12112 11612 12124
rect 11664 12152 11670 12164
rect 12526 12152 12532 12164
rect 11664 12124 12532 12152
rect 11664 12112 11670 12124
rect 12526 12112 12532 12124
rect 12584 12112 12590 12164
rect 566 12044 572 12096
rect 624 12084 630 12096
rect 1029 12087 1087 12093
rect 1029 12084 1041 12087
rect 624 12056 1041 12084
rect 624 12044 630 12056
rect 1029 12053 1041 12056
rect 1075 12053 1087 12087
rect 1029 12047 1087 12053
rect 2869 12087 2927 12093
rect 2869 12053 2881 12087
rect 2915 12084 2927 12087
rect 3234 12084 3240 12096
rect 2915 12056 3240 12084
rect 2915 12053 2927 12056
rect 2869 12047 2927 12053
rect 3234 12044 3240 12056
rect 3292 12044 3298 12096
rect 4614 12044 4620 12096
rect 4672 12044 4678 12096
rect 5350 12044 5356 12096
rect 5408 12044 5414 12096
rect 5626 12044 5632 12096
rect 5684 12084 5690 12096
rect 5994 12084 6000 12096
rect 5684 12056 6000 12084
rect 5684 12044 5690 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6730 12044 6736 12096
rect 6788 12084 6794 12096
rect 7009 12087 7067 12093
rect 7009 12084 7021 12087
rect 6788 12056 7021 12084
rect 6788 12044 6794 12056
rect 7009 12053 7021 12056
rect 7055 12053 7067 12087
rect 7009 12047 7067 12053
rect 7098 12044 7104 12096
rect 7156 12044 7162 12096
rect 7469 12087 7527 12093
rect 7469 12053 7481 12087
rect 7515 12084 7527 12087
rect 7650 12084 7656 12096
rect 7515 12056 7656 12084
rect 7515 12053 7527 12056
rect 7469 12047 7527 12053
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8386 12044 8392 12096
rect 8444 12044 8450 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 10318 12084 10324 12096
rect 9272 12056 10324 12084
rect 9272 12044 9278 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10410 12044 10416 12096
rect 10468 12044 10474 12096
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10652 12056 11069 12084
rect 10652 12044 10658 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11057 12047 11115 12053
rect 11330 12044 11336 12096
rect 11388 12084 11394 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11388 12056 11989 12084
rect 11388 12044 11394 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 11977 12047 12035 12053
rect 552 11994 12604 12016
rect 552 11942 3662 11994
rect 3714 11942 3726 11994
rect 3778 11942 3790 11994
rect 3842 11942 3854 11994
rect 3906 11942 3918 11994
rect 3970 11942 10062 11994
rect 10114 11942 10126 11994
rect 10178 11942 10190 11994
rect 10242 11942 10254 11994
rect 10306 11942 10318 11994
rect 10370 11942 12604 11994
rect 552 11920 12604 11942
rect 1026 11840 1032 11892
rect 1084 11880 1090 11892
rect 1084 11852 2268 11880
rect 1084 11840 1090 11852
rect 2240 11812 2268 11852
rect 2682 11840 2688 11892
rect 2740 11840 2746 11892
rect 2866 11840 2872 11892
rect 2924 11880 2930 11892
rect 6273 11883 6331 11889
rect 2924 11852 6224 11880
rect 2924 11840 2930 11852
rect 5442 11812 5448 11824
rect 2240 11784 2774 11812
rect 2746 11744 2774 11784
rect 4264 11784 5448 11812
rect 4154 11744 4160 11756
rect 2746 11716 4160 11744
rect 4154 11704 4160 11716
rect 4212 11704 4218 11756
rect 1118 11636 1124 11688
rect 1176 11676 1182 11688
rect 1213 11679 1271 11685
rect 1213 11676 1225 11679
rect 1176 11648 1225 11676
rect 1176 11636 1182 11648
rect 1213 11645 1225 11648
rect 1259 11645 1271 11679
rect 1213 11639 1271 11645
rect 1305 11679 1363 11685
rect 1305 11645 1317 11679
rect 1351 11676 1363 11679
rect 3973 11679 4031 11685
rect 1351 11648 2268 11676
rect 1351 11645 1363 11648
rect 1305 11639 1363 11645
rect 2240 11620 2268 11648
rect 3973 11645 3985 11679
rect 4019 11676 4031 11679
rect 4264 11676 4292 11784
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5813 11815 5871 11821
rect 5813 11781 5825 11815
rect 5859 11812 5871 11815
rect 5994 11812 6000 11824
rect 5859 11784 6000 11812
rect 5859 11781 5871 11784
rect 5813 11775 5871 11781
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 6196 11812 6224 11852
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 6362 11880 6368 11892
rect 6319 11852 6368 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 6362 11840 6368 11852
rect 6420 11840 6426 11892
rect 7650 11840 7656 11892
rect 7708 11840 7714 11892
rect 8481 11883 8539 11889
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 8570 11880 8576 11892
rect 8527 11852 8576 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 8849 11883 8907 11889
rect 8849 11880 8861 11883
rect 8720 11852 8861 11880
rect 8720 11840 8726 11852
rect 8849 11849 8861 11852
rect 8895 11849 8907 11883
rect 8849 11843 8907 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 9858 11880 9864 11892
rect 9815 11852 9864 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11425 11883 11483 11889
rect 11425 11880 11437 11883
rect 11204 11852 11437 11880
rect 11204 11840 11210 11852
rect 11425 11849 11437 11852
rect 11471 11849 11483 11883
rect 11425 11843 11483 11849
rect 11701 11883 11759 11889
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 11882 11880 11888 11892
rect 11747 11852 11888 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 6196 11784 8524 11812
rect 8496 11756 8524 11784
rect 9582 11772 9588 11824
rect 9640 11772 9646 11824
rect 10962 11772 10968 11824
rect 11020 11812 11026 11824
rect 11020 11784 11284 11812
rect 11020 11772 11026 11784
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4709 11747 4767 11753
rect 4709 11744 4721 11747
rect 4387 11716 4721 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4709 11713 4721 11716
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11744 5595 11747
rect 6641 11747 6699 11753
rect 6641 11744 6653 11747
rect 5583 11716 5856 11744
rect 5583 11713 5595 11716
rect 5537 11707 5595 11713
rect 5828 11688 5856 11716
rect 5920 11716 6653 11744
rect 4019 11648 4292 11676
rect 4019 11645 4031 11648
rect 3973 11639 4031 11645
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 4801 11679 4859 11685
rect 4801 11676 4813 11679
rect 4724 11648 4813 11676
rect 4724 11620 4752 11648
rect 4801 11645 4813 11648
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 5074 11676 5080 11688
rect 4939 11648 5080 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 5074 11636 5080 11648
rect 5132 11636 5138 11688
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 5626 11676 5632 11688
rect 5500 11648 5632 11676
rect 5500 11636 5506 11648
rect 5626 11636 5632 11648
rect 5684 11636 5690 11688
rect 5810 11636 5816 11688
rect 5868 11636 5874 11688
rect 1578 11617 1584 11620
rect 1572 11608 1584 11617
rect 1539 11580 1584 11608
rect 1572 11571 1584 11580
rect 1578 11568 1584 11571
rect 1636 11568 1642 11620
rect 2222 11568 2228 11620
rect 2280 11568 2286 11620
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4338 11608 4344 11620
rect 4203 11580 4344 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4338 11568 4344 11580
rect 4396 11568 4402 11620
rect 4706 11568 4712 11620
rect 4764 11568 4770 11620
rect 4982 11568 4988 11620
rect 5040 11608 5046 11620
rect 5920 11608 5948 11716
rect 6641 11713 6653 11716
rect 6687 11744 6699 11747
rect 8202 11744 8208 11756
rect 6687 11716 8208 11744
rect 6687 11713 6699 11716
rect 6641 11707 6699 11713
rect 5994 11636 6000 11688
rect 6052 11676 6058 11688
rect 6457 11679 6515 11685
rect 6457 11676 6469 11679
rect 6052 11648 6469 11676
rect 6052 11636 6058 11648
rect 6457 11645 6469 11648
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 6730 11636 6736 11688
rect 6788 11636 6794 11688
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 5040 11580 5948 11608
rect 5040 11568 5046 11580
rect 6362 11568 6368 11620
rect 6420 11608 6426 11620
rect 6932 11608 6960 11639
rect 7006 11636 7012 11688
rect 7064 11636 7070 11688
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11645 7159 11679
rect 7101 11639 7159 11645
rect 7285 11679 7343 11685
rect 7285 11645 7297 11679
rect 7331 11676 7343 11679
rect 7466 11676 7472 11688
rect 7331 11648 7472 11676
rect 7331 11645 7343 11648
rect 7285 11639 7343 11645
rect 6420 11580 6960 11608
rect 7116 11608 7144 11639
rect 7466 11636 7472 11648
rect 7524 11636 7530 11688
rect 7852 11685 7880 11716
rect 8202 11704 8208 11716
rect 8260 11744 8266 11756
rect 8260 11716 8340 11744
rect 8260 11704 8266 11716
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 8018 11636 8024 11688
rect 8076 11676 8082 11688
rect 8113 11679 8171 11685
rect 8113 11676 8125 11679
rect 8076 11648 8125 11676
rect 8076 11636 8082 11648
rect 8113 11645 8125 11648
rect 8159 11645 8171 11679
rect 8113 11639 8171 11645
rect 8202 11608 8208 11620
rect 7116 11580 8208 11608
rect 6420 11568 6426 11580
rect 8202 11568 8208 11580
rect 8260 11568 8266 11620
rect 8312 11608 8340 11716
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8478 11704 8484 11756
rect 8536 11704 8542 11756
rect 9600 11744 9628 11772
rect 10410 11744 10416 11756
rect 8680 11716 9628 11744
rect 10060 11716 10416 11744
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 8680 11685 8708 11716
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8757 11679 8815 11685
rect 8757 11645 8769 11679
rect 8803 11676 8815 11679
rect 8846 11676 8852 11688
rect 8803 11648 8852 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 8941 11679 8999 11685
rect 8941 11645 8953 11679
rect 8987 11676 8999 11679
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 8987 11648 9413 11676
rect 8987 11645 8999 11648
rect 8941 11639 8999 11645
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9401 11639 9459 11645
rect 8956 11608 8984 11639
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9548 11648 9597 11676
rect 9548 11636 9554 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9861 11679 9919 11685
rect 9861 11676 9873 11679
rect 9732 11648 9873 11676
rect 9732 11636 9738 11648
rect 9861 11645 9873 11648
rect 9907 11645 9919 11679
rect 9861 11639 9919 11645
rect 9950 11636 9956 11688
rect 10008 11636 10014 11688
rect 10060 11685 10088 11716
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 11256 11744 11284 11784
rect 11256 11716 11836 11744
rect 10045 11679 10103 11685
rect 10045 11645 10057 11679
rect 10091 11645 10103 11679
rect 10045 11639 10103 11645
rect 10226 11636 10232 11688
rect 10284 11676 10290 11688
rect 10686 11676 10692 11688
rect 10284 11648 10692 11676
rect 10284 11636 10290 11648
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11146 11676 11152 11688
rect 10919 11648 11152 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 11146 11636 11152 11648
rect 11204 11636 11210 11688
rect 11532 11685 11560 11716
rect 11333 11679 11391 11685
rect 11333 11645 11345 11679
rect 11379 11676 11391 11679
rect 11517 11679 11575 11685
rect 11379 11648 11468 11676
rect 11379 11645 11391 11648
rect 11333 11639 11391 11645
rect 8312 11580 8984 11608
rect 9968 11608 9996 11636
rect 10597 11611 10655 11617
rect 10597 11608 10609 11611
rect 9968 11580 10609 11608
rect 10597 11577 10609 11580
rect 10643 11577 10655 11611
rect 11440 11608 11468 11648
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 11808 11685 11836 11716
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 11698 11608 11704 11620
rect 11440 11580 11704 11608
rect 10597 11571 10655 11577
rect 11698 11568 11704 11580
rect 11756 11568 11762 11620
rect 1026 11500 1032 11552
rect 1084 11500 1090 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4433 11543 4491 11549
rect 4433 11540 4445 11543
rect 4304 11512 4445 11540
rect 4304 11500 4310 11512
rect 4433 11509 4445 11512
rect 4479 11509 4491 11543
rect 4433 11503 4491 11509
rect 7006 11500 7012 11552
rect 7064 11540 7070 11552
rect 7469 11543 7527 11549
rect 7469 11540 7481 11543
rect 7064 11512 7481 11540
rect 7064 11500 7070 11512
rect 7469 11509 7481 11512
rect 7515 11509 7527 11543
rect 7469 11503 7527 11509
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8021 11543 8079 11549
rect 8021 11540 8033 11543
rect 7892 11512 8033 11540
rect 7892 11500 7898 11512
rect 8021 11509 8033 11512
rect 8067 11540 8079 11543
rect 8110 11540 8116 11552
rect 8067 11512 8116 11540
rect 8067 11509 8079 11512
rect 8021 11503 8079 11509
rect 8110 11500 8116 11512
rect 8168 11500 8174 11552
rect 9953 11543 10011 11549
rect 9953 11509 9965 11543
rect 9999 11540 10011 11543
rect 10042 11540 10048 11552
rect 9999 11512 10048 11540
rect 9999 11509 10011 11512
rect 9953 11503 10011 11509
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10413 11543 10471 11549
rect 10413 11540 10425 11543
rect 10376 11512 10425 11540
rect 10376 11500 10382 11512
rect 10413 11509 10425 11512
rect 10459 11509 10471 11543
rect 10413 11503 10471 11509
rect 11238 11500 11244 11552
rect 11296 11500 11302 11552
rect 552 11450 12604 11472
rect 552 11398 4322 11450
rect 4374 11398 4386 11450
rect 4438 11398 4450 11450
rect 4502 11398 4514 11450
rect 4566 11398 4578 11450
rect 4630 11398 10722 11450
rect 10774 11398 10786 11450
rect 10838 11398 10850 11450
rect 10902 11398 10914 11450
rect 10966 11398 10978 11450
rect 11030 11398 12604 11450
rect 552 11376 12604 11398
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4764 11308 5273 11336
rect 4764 11296 4770 11308
rect 5261 11305 5273 11308
rect 5307 11336 5319 11339
rect 6638 11336 6644 11348
rect 5307 11308 6644 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 6914 11296 6920 11348
rect 6972 11296 6978 11348
rect 7098 11296 7104 11348
rect 7156 11336 7162 11348
rect 7282 11336 7288 11348
rect 7156 11308 7288 11336
rect 7156 11296 7162 11308
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7929 11339 7987 11345
rect 7929 11336 7941 11339
rect 7432 11308 7941 11336
rect 7432 11296 7438 11308
rect 7929 11305 7941 11308
rect 7975 11305 7987 11339
rect 7929 11299 7987 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8846 11336 8852 11348
rect 8260 11308 8852 11336
rect 8260 11296 8266 11308
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 8938 11296 8944 11348
rect 8996 11336 9002 11348
rect 9401 11339 9459 11345
rect 9401 11336 9413 11339
rect 8996 11308 9413 11336
rect 8996 11296 9002 11308
rect 9401 11305 9413 11308
rect 9447 11305 9459 11339
rect 9401 11299 9459 11305
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 10686 11336 10692 11348
rect 10284 11308 10692 11336
rect 10284 11296 10290 11308
rect 10686 11296 10692 11308
rect 10744 11296 10750 11348
rect 1670 11228 1676 11280
rect 1728 11268 1734 11280
rect 1728 11240 2360 11268
rect 1728 11228 1734 11240
rect 2332 11212 2360 11240
rect 5626 11228 5632 11280
rect 5684 11268 5690 11280
rect 5684 11240 6316 11268
rect 5684 11228 5690 11240
rect 1946 11160 1952 11212
rect 2004 11209 2010 11212
rect 2004 11200 2016 11209
rect 2004 11172 2049 11200
rect 2004 11163 2016 11172
rect 2004 11160 2010 11163
rect 2314 11160 2320 11212
rect 2372 11160 2378 11212
rect 5074 11160 5080 11212
rect 5132 11160 5138 11212
rect 5350 11160 5356 11212
rect 5408 11160 5414 11212
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6086 11160 6092 11212
rect 6144 11160 6150 11212
rect 6288 11209 6316 11240
rect 7466 11228 7472 11280
rect 7524 11268 7530 11280
rect 9582 11268 9588 11280
rect 7524 11240 9588 11268
rect 7524 11228 7530 11240
rect 9582 11228 9588 11240
rect 9640 11268 9646 11280
rect 10962 11268 10968 11280
rect 9640 11240 10272 11268
rect 9640 11228 9646 11240
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11169 6331 11203
rect 6273 11163 6331 11169
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11200 6423 11203
rect 6546 11200 6552 11212
rect 6411 11172 6552 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6546 11160 6552 11172
rect 6604 11200 6610 11212
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6604 11172 6837 11200
rect 6604 11160 6610 11172
rect 6825 11169 6837 11172
rect 6871 11200 6883 11203
rect 6914 11200 6920 11212
rect 6871 11172 6920 11200
rect 6871 11169 6883 11172
rect 6825 11163 6883 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7006 11160 7012 11212
rect 7064 11160 7070 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 7926 11200 7932 11212
rect 7883 11172 7932 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 8021 11203 8079 11209
rect 8021 11169 8033 11203
rect 8067 11200 8079 11203
rect 8110 11200 8116 11212
rect 8067 11172 8116 11200
rect 8067 11169 8079 11172
rect 8021 11163 8079 11169
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 9766 11160 9772 11212
rect 9824 11160 9830 11212
rect 10042 11160 10048 11212
rect 10100 11160 10106 11212
rect 10244 11209 10272 11240
rect 10336 11240 10968 11268
rect 10336 11209 10364 11240
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10410 11160 10416 11212
rect 10468 11160 10474 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 12158 11200 12164 11212
rect 11379 11172 12164 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 2222 11092 2228 11144
rect 2280 11092 2286 11144
rect 6012 11132 6040 11160
rect 7374 11132 7380 11144
rect 6012 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 9582 11092 9588 11144
rect 9640 11092 9646 11144
rect 9674 11092 9680 11144
rect 9732 11092 9738 11144
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 10689 11135 10747 11141
rect 10689 11132 10701 11135
rect 9907 11104 10701 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 10689 11101 10701 11104
rect 10735 11101 10747 11135
rect 10689 11095 10747 11101
rect 10870 11092 10876 11144
rect 10928 11132 10934 11144
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 10928 11104 11253 11132
rect 10928 11092 10934 11104
rect 11241 11101 11253 11104
rect 11287 11101 11299 11135
rect 11241 11095 11299 11101
rect 845 11067 903 11073
rect 845 11033 857 11067
rect 891 11064 903 11067
rect 891 11036 1348 11064
rect 891 11033 903 11036
rect 845 11027 903 11033
rect 1320 10996 1348 11036
rect 2498 11024 2504 11076
rect 2556 11024 2562 11076
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4764 11036 4905 11064
rect 4764 11024 4770 11036
rect 4893 11033 4905 11036
rect 4939 11033 4951 11067
rect 4893 11027 4951 11033
rect 7650 11024 7656 11076
rect 7708 11064 7714 11076
rect 10318 11064 10324 11076
rect 7708 11036 10324 11064
rect 7708 11024 7714 11036
rect 10318 11024 10324 11036
rect 10376 11064 10382 11076
rect 11348 11064 11376 11163
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 10376 11036 11376 11064
rect 10376 11024 10382 11036
rect 1578 10996 1584 11008
rect 1320 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 5534 10956 5540 11008
rect 5592 10996 5598 11008
rect 5813 10999 5871 11005
rect 5813 10996 5825 10999
rect 5592 10968 5825 10996
rect 5592 10956 5598 10968
rect 5813 10965 5825 10968
rect 5859 10965 5871 10999
rect 5813 10959 5871 10965
rect 10965 10999 11023 11005
rect 10965 10965 10977 10999
rect 11011 10996 11023 10999
rect 11238 10996 11244 11008
rect 11011 10968 11244 10996
rect 11011 10965 11023 10968
rect 10965 10959 11023 10965
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 552 10906 12604 10928
rect 552 10854 3662 10906
rect 3714 10854 3726 10906
rect 3778 10854 3790 10906
rect 3842 10854 3854 10906
rect 3906 10854 3918 10906
rect 3970 10854 10062 10906
rect 10114 10854 10126 10906
rect 10178 10854 10190 10906
rect 10242 10854 10254 10906
rect 10306 10854 10318 10906
rect 10370 10854 12604 10906
rect 552 10832 12604 10854
rect 2314 10752 2320 10804
rect 2372 10752 2378 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 3099 10764 3525 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 3970 10752 3976 10804
rect 4028 10792 4034 10804
rect 4154 10792 4160 10804
rect 4028 10764 4160 10792
rect 4028 10752 4034 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 5718 10752 5724 10804
rect 5776 10792 5782 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 5776 10764 6377 10792
rect 5776 10752 5782 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 9493 10795 9551 10801
rect 8168 10764 9444 10792
rect 8168 10752 8174 10764
rect 3326 10684 3332 10736
rect 3384 10724 3390 10736
rect 3881 10727 3939 10733
rect 3881 10724 3893 10727
rect 3384 10696 3893 10724
rect 3384 10684 3390 10696
rect 3881 10693 3893 10696
rect 3927 10693 3939 10727
rect 6914 10724 6920 10736
rect 3881 10687 3939 10693
rect 3989 10696 6920 10724
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1029 10659 1087 10665
rect 1029 10656 1041 10659
rect 992 10628 1041 10656
rect 992 10616 998 10628
rect 1029 10625 1041 10628
rect 1075 10625 1087 10659
rect 1029 10619 1087 10625
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 1765 10659 1823 10665
rect 1765 10656 1777 10659
rect 1636 10628 1777 10656
rect 1636 10616 1642 10628
rect 1765 10625 1777 10628
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 3989 10656 4017 10696
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 9122 10684 9128 10736
rect 9180 10684 9186 10736
rect 9416 10724 9444 10764
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 9582 10792 9588 10804
rect 9539 10764 9588 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9582 10752 9588 10764
rect 9640 10752 9646 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10045 10795 10103 10801
rect 10045 10792 10057 10795
rect 9732 10764 10057 10792
rect 9732 10752 9738 10764
rect 10045 10761 10057 10764
rect 10091 10761 10103 10795
rect 10045 10755 10103 10761
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 11020 10764 11805 10792
rect 11020 10752 11026 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 11974 10724 11980 10736
rect 9416 10696 11980 10724
rect 11974 10684 11980 10696
rect 12032 10684 12038 10736
rect 3651 10628 4017 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4120 10628 4476 10656
rect 4120 10616 4126 10628
rect 1394 10548 1400 10600
rect 1452 10588 1458 10600
rect 1489 10591 1547 10597
rect 1489 10588 1501 10591
rect 1452 10560 1501 10588
rect 1452 10548 1458 10560
rect 1489 10557 1501 10560
rect 1535 10557 1547 10591
rect 1489 10551 1547 10557
rect 1673 10591 1731 10597
rect 1673 10557 1685 10591
rect 1719 10588 1731 10591
rect 1946 10588 1952 10600
rect 1719 10560 1952 10588
rect 1719 10557 1731 10560
rect 1673 10551 1731 10557
rect 1946 10548 1952 10560
rect 2004 10548 2010 10600
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 2958 10588 2964 10600
rect 2823 10560 2964 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3510 10548 3516 10600
rect 3568 10548 3574 10600
rect 4154 10548 4160 10600
rect 4212 10548 4218 10600
rect 4448 10597 4476 10628
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6089 10659 6147 10665
rect 6089 10656 6101 10659
rect 5960 10628 6101 10656
rect 5960 10616 5966 10628
rect 6089 10625 6101 10628
rect 6135 10625 6147 10659
rect 6089 10619 6147 10625
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10656 6331 10659
rect 6454 10656 6460 10668
rect 6319 10628 6460 10656
rect 6319 10625 6331 10628
rect 6273 10619 6331 10625
rect 6454 10616 6460 10628
rect 6512 10656 6518 10668
rect 7561 10659 7619 10665
rect 7561 10656 7573 10659
rect 6512 10628 7573 10656
rect 6512 10616 6518 10628
rect 7561 10625 7573 10628
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 7834 10616 7840 10668
rect 7892 10656 7898 10668
rect 9582 10656 9588 10668
rect 7892 10628 9588 10656
rect 7892 10616 7898 10628
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11238 10656 11244 10668
rect 11011 10628 11244 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 4249 10591 4307 10597
rect 4249 10557 4261 10591
rect 4295 10588 4307 10591
rect 4433 10591 4491 10597
rect 4295 10560 4384 10588
rect 4295 10557 4307 10560
rect 4249 10551 4307 10557
rect 658 10480 664 10532
rect 716 10520 722 10532
rect 2869 10523 2927 10529
rect 2869 10520 2881 10523
rect 716 10492 2881 10520
rect 716 10480 722 10492
rect 2792 10464 2820 10492
rect 2869 10489 2881 10492
rect 2915 10489 2927 10523
rect 2869 10483 2927 10489
rect 3053 10523 3111 10529
rect 3053 10489 3065 10523
rect 3099 10520 3111 10523
rect 3142 10520 3148 10532
rect 3099 10492 3148 10520
rect 3099 10489 3111 10492
rect 3053 10483 3111 10489
rect 3142 10480 3148 10492
rect 3200 10480 3206 10532
rect 2774 10412 2780 10464
rect 2832 10412 2838 10464
rect 3973 10455 4031 10461
rect 3973 10421 3985 10455
rect 4019 10452 4031 10455
rect 4062 10452 4068 10464
rect 4019 10424 4068 10452
rect 4019 10421 4031 10424
rect 3973 10415 4031 10421
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 4356 10452 4384 10560
rect 4433 10557 4445 10591
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10588 4583 10591
rect 4890 10588 4896 10600
rect 4571 10560 4896 10588
rect 4571 10557 4583 10560
rect 4525 10551 4583 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5350 10588 5356 10600
rect 5224 10560 5356 10588
rect 5224 10548 5230 10560
rect 5350 10548 5356 10560
rect 5408 10548 5414 10600
rect 5997 10591 6055 10597
rect 5997 10557 6009 10591
rect 6043 10588 6055 10591
rect 6196 10588 6224 10616
rect 6043 10560 6224 10588
rect 6043 10557 6055 10560
rect 5997 10551 6055 10557
rect 6546 10548 6552 10600
rect 6604 10548 6610 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 4908 10520 4936 10548
rect 6086 10520 6092 10532
rect 4908 10492 6092 10520
rect 6086 10480 6092 10492
rect 6144 10520 6150 10532
rect 6656 10520 6684 10551
rect 6144 10492 6684 10520
rect 6840 10520 6868 10551
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 7469 10591 7527 10597
rect 7469 10588 7481 10591
rect 7432 10560 7481 10588
rect 7432 10548 7438 10560
rect 7469 10557 7481 10560
rect 7515 10557 7527 10591
rect 7469 10551 7527 10557
rect 7650 10548 7656 10600
rect 7708 10548 7714 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9692 10560 9965 10588
rect 7098 10520 7104 10532
rect 6840 10492 7104 10520
rect 6144 10480 6150 10492
rect 7098 10480 7104 10492
rect 7156 10480 7162 10532
rect 7193 10523 7251 10529
rect 7193 10489 7205 10523
rect 7239 10520 7251 10523
rect 7668 10520 7696 10548
rect 9692 10532 9720 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10137 10591 10195 10597
rect 10137 10557 10149 10591
rect 10183 10588 10195 10591
rect 10502 10588 10508 10600
rect 10183 10560 10508 10588
rect 10183 10557 10195 10560
rect 10137 10551 10195 10557
rect 7239 10492 7696 10520
rect 8757 10523 8815 10529
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 8757 10489 8769 10523
rect 8803 10520 8815 10523
rect 8846 10520 8852 10532
rect 8803 10492 8852 10520
rect 8803 10489 8815 10492
rect 8757 10483 8815 10489
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 9674 10480 9680 10532
rect 9732 10480 9738 10532
rect 9858 10480 9864 10532
rect 9916 10520 9922 10532
rect 10152 10520 10180 10551
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10594 10548 10600 10600
rect 10652 10588 10658 10600
rect 10873 10591 10931 10597
rect 10873 10588 10885 10591
rect 10652 10560 10885 10588
rect 10652 10548 10658 10560
rect 10873 10557 10885 10560
rect 10919 10557 10931 10591
rect 10873 10551 10931 10557
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11333 10591 11391 10597
rect 11333 10588 11345 10591
rect 11112 10560 11345 10588
rect 11112 10548 11118 10560
rect 11333 10557 11345 10560
rect 11379 10557 11391 10591
rect 11333 10551 11391 10557
rect 11609 10591 11667 10597
rect 11609 10557 11621 10591
rect 11655 10588 11667 10591
rect 11790 10588 11796 10600
rect 11655 10560 11796 10588
rect 11655 10557 11667 10560
rect 11609 10551 11667 10557
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 9916 10492 10180 10520
rect 9916 10480 9922 10492
rect 4982 10452 4988 10464
rect 4356 10424 4988 10452
rect 4982 10412 4988 10424
rect 5040 10452 5046 10464
rect 5166 10452 5172 10464
rect 5040 10424 5172 10452
rect 5040 10412 5046 10424
rect 5166 10412 5172 10424
rect 5224 10412 5230 10464
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5592 10424 6285 10452
rect 5592 10412 5598 10424
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6273 10415 6331 10421
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6972 10424 7021 10452
rect 6972 10412 6978 10424
rect 7009 10421 7021 10424
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 9217 10455 9275 10461
rect 9217 10421 9229 10455
rect 9263 10452 9275 10455
rect 9398 10452 9404 10464
rect 9263 10424 9404 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 10870 10452 10876 10464
rect 10560 10424 10876 10452
rect 10560 10412 10566 10424
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11146 10412 11152 10464
rect 11204 10452 11210 10464
rect 11241 10455 11299 10461
rect 11241 10452 11253 10455
rect 11204 10424 11253 10452
rect 11204 10412 11210 10424
rect 11241 10421 11253 10424
rect 11287 10452 11299 10455
rect 11425 10455 11483 10461
rect 11425 10452 11437 10455
rect 11287 10424 11437 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11425 10421 11437 10424
rect 11471 10421 11483 10455
rect 11425 10415 11483 10421
rect 552 10362 12604 10384
rect 552 10310 4322 10362
rect 4374 10310 4386 10362
rect 4438 10310 4450 10362
rect 4502 10310 4514 10362
rect 4566 10310 4578 10362
rect 4630 10310 10722 10362
rect 10774 10310 10786 10362
rect 10838 10310 10850 10362
rect 10902 10310 10914 10362
rect 10966 10310 10978 10362
rect 11030 10310 12604 10362
rect 552 10288 12604 10310
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 4614 10248 4620 10260
rect 3108 10220 4620 10248
rect 3108 10208 3114 10220
rect 1854 10140 1860 10192
rect 1912 10180 1918 10192
rect 1958 10183 2016 10189
rect 1958 10180 1970 10183
rect 1912 10152 1970 10180
rect 1912 10140 1918 10152
rect 1958 10149 1970 10152
rect 2004 10149 2016 10183
rect 1958 10143 2016 10149
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3329 10115 3387 10121
rect 3329 10112 3341 10115
rect 3016 10084 3341 10112
rect 3016 10072 3022 10084
rect 3329 10081 3341 10084
rect 3375 10112 3387 10115
rect 3602 10112 3608 10124
rect 3375 10084 3608 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 3697 10115 3755 10121
rect 3697 10081 3709 10115
rect 3743 10112 3755 10115
rect 3988 10112 4016 10220
rect 4614 10208 4620 10220
rect 4672 10248 4678 10260
rect 5258 10248 5264 10260
rect 4672 10220 5264 10248
rect 4672 10208 4678 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 8570 10248 8576 10260
rect 8251 10220 8576 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 9125 10251 9183 10257
rect 9125 10217 9137 10251
rect 9171 10248 9183 10251
rect 9585 10251 9643 10257
rect 9585 10248 9597 10251
rect 9171 10220 9597 10248
rect 9171 10217 9183 10220
rect 9125 10211 9183 10217
rect 9585 10217 9597 10220
rect 9631 10248 9643 10251
rect 9674 10248 9680 10260
rect 9631 10220 9680 10248
rect 9631 10217 9643 10220
rect 9585 10211 9643 10217
rect 9674 10208 9680 10220
rect 9732 10208 9738 10260
rect 4890 10180 4896 10192
rect 4540 10152 4896 10180
rect 4540 10121 4568 10152
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 5077 10183 5135 10189
rect 5077 10149 5089 10183
rect 5123 10180 5135 10183
rect 5166 10180 5172 10192
rect 5123 10152 5172 10180
rect 5123 10149 5135 10152
rect 5077 10143 5135 10149
rect 5166 10140 5172 10152
rect 5224 10140 5230 10192
rect 7926 10180 7932 10192
rect 7852 10152 7932 10180
rect 3743 10084 4016 10112
rect 4525 10115 4583 10121
rect 3743 10081 3755 10084
rect 3697 10075 3755 10081
rect 4525 10081 4537 10115
rect 4571 10081 4583 10115
rect 4525 10075 4583 10081
rect 4614 10072 4620 10124
rect 4672 10072 4678 10124
rect 4798 10072 4804 10124
rect 4856 10072 4862 10124
rect 4982 10072 4988 10124
rect 5040 10072 5046 10124
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10112 5319 10115
rect 6270 10112 6276 10124
rect 5307 10084 6276 10112
rect 5307 10081 5319 10084
rect 5261 10075 5319 10081
rect 2222 10004 2228 10056
rect 2280 10004 2286 10056
rect 3970 10004 3976 10056
rect 4028 10004 4034 10056
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4338 10044 4344 10056
rect 4212 10016 4344 10044
rect 4212 10004 4218 10016
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4709 10047 4767 10053
rect 4709 10013 4721 10047
rect 4755 10013 4767 10047
rect 4709 10007 4767 10013
rect 3326 9936 3332 9988
rect 3384 9976 3390 9988
rect 3988 9976 4016 10004
rect 3384 9948 4016 9976
rect 4724 9976 4752 10007
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5276 10044 5304 10075
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 7558 10072 7564 10124
rect 7616 10072 7622 10124
rect 7852 10121 7880 10152
rect 7926 10140 7932 10152
rect 7984 10180 7990 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 7984 10152 9229 10180
rect 7984 10140 7990 10152
rect 9217 10149 9229 10152
rect 9263 10149 9275 10183
rect 9858 10180 9864 10192
rect 9217 10143 9275 10149
rect 9692 10152 9864 10180
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8297 10115 8355 10121
rect 8297 10081 8309 10115
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 4948 10016 5304 10044
rect 4948 10004 4954 10016
rect 7650 10004 7656 10056
rect 7708 10044 7714 10056
rect 7745 10047 7803 10053
rect 7745 10044 7757 10047
rect 7708 10016 7757 10044
rect 7708 10004 7714 10016
rect 7745 10013 7757 10016
rect 7791 10013 7803 10047
rect 7745 10007 7803 10013
rect 4798 9976 4804 9988
rect 4724 9948 4804 9976
rect 3384 9936 3390 9948
rect 4798 9936 4804 9948
rect 4856 9936 4862 9988
rect 6822 9936 6828 9988
rect 6880 9976 6886 9988
rect 8312 9976 8340 10075
rect 8478 10072 8484 10124
rect 8536 10072 8542 10124
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 8846 10112 8852 10124
rect 8803 10084 8852 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 8846 10072 8852 10084
rect 8904 10072 8910 10124
rect 9398 10072 9404 10124
rect 9456 10072 9462 10124
rect 9692 10121 9720 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 11422 10140 11428 10192
rect 11480 10180 11486 10192
rect 11517 10183 11575 10189
rect 11517 10180 11529 10183
rect 11480 10152 11529 10180
rect 11480 10140 11486 10152
rect 11517 10149 11529 10152
rect 11563 10180 11575 10183
rect 11563 10152 11928 10180
rect 11563 10149 11575 10152
rect 11517 10143 11575 10149
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9769 10115 9827 10121
rect 9769 10081 9781 10115
rect 9815 10112 9827 10115
rect 9953 10115 10011 10121
rect 9815 10084 9904 10112
rect 9815 10081 9827 10084
rect 9769 10075 9827 10081
rect 9876 10056 9904 10084
rect 9953 10081 9965 10115
rect 9999 10112 10011 10115
rect 10778 10112 10784 10124
rect 9999 10084 10784 10112
rect 9999 10081 10011 10084
rect 9953 10075 10011 10081
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11054 10112 11060 10124
rect 11011 10084 11060 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11146 10072 11152 10124
rect 11204 10072 11210 10124
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10112 11759 10115
rect 11790 10112 11796 10124
rect 11747 10084 11796 10112
rect 11747 10081 11759 10084
rect 11701 10075 11759 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 11900 10121 11928 10152
rect 11885 10115 11943 10121
rect 11885 10081 11897 10115
rect 11931 10081 11943 10115
rect 11885 10075 11943 10081
rect 11974 10072 11980 10124
rect 12032 10072 12038 10124
rect 8386 10004 8392 10056
rect 8444 10004 8450 10056
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10044 8723 10047
rect 9122 10044 9128 10056
rect 8711 10016 9128 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 10502 10044 10508 10056
rect 9916 10016 10508 10044
rect 9916 10004 9922 10016
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10044 12219 10047
rect 12250 10044 12256 10056
rect 12207 10016 12256 10044
rect 12207 10013 12219 10016
rect 12161 10007 12219 10013
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 6880 9948 8340 9976
rect 6880 9936 6886 9948
rect 10410 9936 10416 9988
rect 10468 9976 10474 9988
rect 10965 9979 11023 9985
rect 10965 9976 10977 9979
rect 10468 9948 10977 9976
rect 10468 9936 10474 9948
rect 10965 9945 10977 9948
rect 11011 9945 11023 9979
rect 10965 9939 11023 9945
rect 845 9911 903 9917
rect 845 9877 857 9911
rect 891 9908 903 9911
rect 1946 9908 1952 9920
rect 891 9880 1952 9908
rect 891 9877 903 9880
rect 845 9871 903 9877
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4341 9911 4399 9917
rect 4341 9908 4353 9911
rect 4212 9880 4353 9908
rect 4212 9868 4218 9880
rect 4341 9877 4353 9880
rect 4387 9877 4399 9911
rect 4341 9871 4399 9877
rect 5074 9868 5080 9920
rect 5132 9908 5138 9920
rect 5445 9911 5503 9917
rect 5445 9908 5457 9911
rect 5132 9880 5457 9908
rect 5132 9868 5138 9880
rect 5445 9877 5457 9880
rect 5491 9908 5503 9911
rect 5810 9908 5816 9920
rect 5491 9880 5816 9908
rect 5491 9877 5503 9880
rect 5445 9871 5503 9877
rect 5810 9868 5816 9880
rect 5868 9868 5874 9920
rect 6270 9868 6276 9920
rect 6328 9868 6334 9920
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 9769 9911 9827 9917
rect 9769 9908 9781 9911
rect 9732 9880 9781 9908
rect 9732 9868 9738 9880
rect 9769 9877 9781 9880
rect 9815 9877 9827 9911
rect 9769 9871 9827 9877
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 552 9818 12604 9840
rect 552 9766 3662 9818
rect 3714 9766 3726 9818
rect 3778 9766 3790 9818
rect 3842 9766 3854 9818
rect 3906 9766 3918 9818
rect 3970 9766 10062 9818
rect 10114 9766 10126 9818
rect 10178 9766 10190 9818
rect 10242 9766 10254 9818
rect 10306 9766 10318 9818
rect 10370 9766 12604 9818
rect 552 9744 12604 9766
rect 3142 9664 3148 9716
rect 3200 9704 3206 9716
rect 3602 9704 3608 9716
rect 3200 9676 3608 9704
rect 3200 9664 3206 9676
rect 3602 9664 3608 9676
rect 3660 9664 3666 9716
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4338 9704 4344 9716
rect 4028 9676 4344 9704
rect 4028 9664 4034 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 6472 9676 6776 9704
rect 750 9596 756 9648
rect 808 9636 814 9648
rect 3237 9639 3295 9645
rect 3237 9636 3249 9639
rect 808 9608 3249 9636
rect 808 9596 814 9608
rect 3237 9605 3249 9608
rect 3283 9605 3295 9639
rect 3237 9599 3295 9605
rect 3418 9596 3424 9648
rect 3476 9636 3482 9648
rect 3881 9639 3939 9645
rect 3881 9636 3893 9639
rect 3476 9608 3893 9636
rect 3476 9596 3482 9608
rect 3881 9605 3893 9608
rect 3927 9605 3939 9639
rect 3881 9599 3939 9605
rect 4062 9596 4068 9648
rect 4120 9596 4126 9648
rect 5350 9596 5356 9648
rect 5408 9636 5414 9648
rect 6472 9636 6500 9676
rect 5408 9608 6500 9636
rect 5408 9596 5414 9608
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6641 9639 6699 9645
rect 6641 9636 6653 9639
rect 6604 9608 6653 9636
rect 6604 9596 6610 9608
rect 6641 9605 6653 9608
rect 6687 9605 6699 9639
rect 6748 9636 6776 9676
rect 7576 9676 7757 9704
rect 7006 9636 7012 9648
rect 6748 9608 7012 9636
rect 6641 9599 6699 9605
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 7576 9636 7604 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 8846 9664 8852 9716
rect 8904 9664 8910 9716
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10778 9704 10784 9716
rect 10551 9676 10784 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 12253 9707 12311 9713
rect 12253 9704 12265 9707
rect 11848 9676 12265 9704
rect 11848 9664 11854 9676
rect 12253 9673 12265 9676
rect 12299 9673 12311 9707
rect 12253 9667 12311 9673
rect 7116 9608 7604 9636
rect 1210 9528 1216 9580
rect 1268 9528 1274 9580
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2406 9528 2412 9580
rect 2464 9528 2470 9580
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4080 9568 4108 9596
rect 3743 9540 4108 9568
rect 4801 9571 4859 9577
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 4982 9568 4988 9580
rect 4847 9540 4988 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5534 9568 5540 9580
rect 5491 9540 5540 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 5721 9571 5779 9577
rect 5721 9537 5733 9571
rect 5767 9568 5779 9571
rect 6917 9571 6975 9577
rect 6917 9568 6929 9571
rect 5767 9540 6929 9568
rect 5767 9537 5779 9540
rect 5721 9531 5779 9537
rect 6656 9512 6684 9540
rect 6917 9537 6929 9540
rect 6963 9537 6975 9571
rect 6917 9531 6975 9537
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 1673 9503 1731 9509
rect 1673 9500 1685 9503
rect 1452 9472 1685 9500
rect 1452 9460 1458 9472
rect 1673 9469 1685 9472
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 1854 9460 1860 9512
rect 1912 9460 1918 9512
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9469 2559 9503
rect 2501 9463 2559 9469
rect 842 9392 848 9444
rect 900 9432 906 9444
rect 2516 9432 2544 9463
rect 3418 9460 3424 9512
rect 3476 9460 3482 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 3513 9463 3571 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3970 9500 3976 9512
rect 3651 9472 3976 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3528 9432 3556 9463
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4065 9503 4123 9509
rect 4065 9469 4077 9503
rect 4111 9502 4123 9503
rect 4154 9502 4160 9512
rect 4111 9474 4160 9502
rect 4111 9469 4123 9474
rect 4065 9463 4123 9469
rect 4154 9460 4160 9474
rect 4212 9460 4218 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 4709 9503 4767 9509
rect 4387 9472 4660 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 3878 9432 3884 9444
rect 900 9404 3464 9432
rect 3528 9404 3884 9432
rect 900 9392 906 9404
rect 2866 9324 2872 9376
rect 2924 9324 2930 9376
rect 3436 9364 3464 9404
rect 3878 9392 3884 9404
rect 3936 9392 3942 9444
rect 4632 9432 4660 9472
rect 4709 9469 4721 9503
rect 4755 9500 4767 9503
rect 5166 9500 5172 9512
rect 4755 9472 5172 9500
rect 4755 9469 4767 9472
rect 4709 9463 4767 9469
rect 5166 9460 5172 9472
rect 5224 9460 5230 9512
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5902 9500 5908 9512
rect 5399 9472 5908 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 4982 9432 4988 9444
rect 4632 9404 4988 9432
rect 4982 9392 4988 9404
rect 5040 9392 5046 9444
rect 3786 9364 3792 9376
rect 3436 9336 3792 9364
rect 3786 9324 3792 9336
rect 3844 9324 3850 9376
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4249 9367 4307 9373
rect 4249 9364 4261 9367
rect 4120 9336 4261 9364
rect 4120 9324 4126 9336
rect 4249 9333 4261 9336
rect 4295 9364 4307 9367
rect 4890 9364 4896 9376
rect 4295 9336 4896 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5077 9367 5135 9373
rect 5077 9333 5089 9367
rect 5123 9364 5135 9367
rect 5368 9364 5396 9463
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 6270 9460 6276 9512
rect 6328 9460 6334 9512
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 6730 9460 6736 9512
rect 6788 9500 6794 9512
rect 7009 9503 7067 9509
rect 7009 9500 7021 9503
rect 6788 9472 7021 9500
rect 6788 9460 6794 9472
rect 7009 9469 7021 9472
rect 7055 9500 7067 9503
rect 7116 9500 7144 9608
rect 7650 9596 7656 9648
rect 7708 9596 7714 9648
rect 9646 9608 10640 9636
rect 7576 9540 8064 9568
rect 7055 9472 7144 9500
rect 7055 9469 7067 9472
rect 7009 9463 7067 9469
rect 7282 9460 7288 9512
rect 7340 9460 7346 9512
rect 7439 9503 7497 9509
rect 7439 9469 7451 9503
rect 7485 9500 7497 9503
rect 7576 9500 7604 9540
rect 8036 9509 8064 9540
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 8260 9540 8493 9568
rect 8260 9528 8266 9540
rect 8481 9537 8493 9540
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9568 9367 9571
rect 9490 9568 9496 9580
rect 9355 9540 9496 9568
rect 9355 9537 9367 9540
rect 9309 9531 9367 9537
rect 9490 9528 9496 9540
rect 9548 9528 9554 9580
rect 8021 9503 8079 9509
rect 7485 9472 7604 9500
rect 7668 9472 7972 9500
rect 7485 9469 7497 9472
rect 7439 9463 7497 9469
rect 6288 9432 6316 9460
rect 7668 9432 7696 9472
rect 6288 9404 7696 9432
rect 7745 9435 7803 9441
rect 7745 9401 7757 9435
rect 7791 9401 7803 9435
rect 7944 9432 7972 9472
rect 8021 9469 8033 9503
rect 8067 9500 8079 9503
rect 8386 9500 8392 9512
rect 8067 9472 8392 9500
rect 8067 9469 8079 9472
rect 8021 9463 8079 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8573 9503 8631 9509
rect 8573 9469 8585 9503
rect 8619 9500 8631 9503
rect 9646 9500 9674 9608
rect 10134 9528 10140 9580
rect 10192 9568 10198 9580
rect 10502 9568 10508 9580
rect 10192 9540 10508 9568
rect 10192 9528 10198 9540
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 10612 9568 10640 9608
rect 10612 9540 11008 9568
rect 9950 9500 9956 9512
rect 8619 9472 9956 9500
rect 8619 9469 8631 9472
rect 8573 9463 8631 9469
rect 9950 9460 9956 9472
rect 10008 9460 10014 9512
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 10594 9500 10600 9512
rect 10100 9472 10600 9500
rect 10100 9460 10106 9472
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10873 9503 10931 9509
rect 10873 9469 10885 9503
rect 10919 9469 10931 9503
rect 10980 9500 11008 9540
rect 11698 9500 11704 9512
rect 10980 9472 11704 9500
rect 10873 9463 10931 9469
rect 10888 9432 10916 9463
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 7944 9404 10916 9432
rect 11140 9435 11198 9441
rect 7745 9395 7803 9401
rect 5123 9336 5396 9364
rect 5123 9333 5135 9336
rect 5077 9327 5135 9333
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7760 9364 7788 9395
rect 10612 9376 10640 9404
rect 11140 9401 11152 9435
rect 11186 9432 11198 9435
rect 12158 9432 12164 9444
rect 11186 9404 12164 9432
rect 11186 9401 11198 9404
rect 11140 9395 11198 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 7340 9336 7788 9364
rect 7340 9324 7346 9336
rect 7926 9324 7932 9376
rect 7984 9324 7990 9376
rect 10594 9324 10600 9376
rect 10652 9324 10658 9376
rect 552 9274 12604 9296
rect 552 9222 4322 9274
rect 4374 9222 4386 9274
rect 4438 9222 4450 9274
rect 4502 9222 4514 9274
rect 4566 9222 4578 9274
rect 4630 9222 10722 9274
rect 10774 9222 10786 9274
rect 10838 9222 10850 9274
rect 10902 9222 10914 9274
rect 10966 9222 10978 9274
rect 11030 9222 12604 9274
rect 552 9200 12604 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 1360 9132 2774 9160
rect 1360 9120 1366 9132
rect 2746 9092 2774 9132
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 3476 9132 3893 9160
rect 3476 9120 3482 9132
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 3970 9120 3976 9172
rect 4028 9160 4034 9172
rect 4341 9163 4399 9169
rect 4341 9160 4353 9163
rect 4028 9132 4353 9160
rect 4028 9120 4034 9132
rect 4341 9129 4353 9132
rect 4387 9129 4399 9163
rect 4341 9123 4399 9129
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 6822 9160 6828 9172
rect 6687 9132 6828 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 6917 9163 6975 9169
rect 6917 9129 6929 9163
rect 6963 9160 6975 9163
rect 7282 9160 7288 9172
rect 6963 9132 7288 9160
rect 6963 9129 6975 9132
rect 6917 9123 6975 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 9122 9120 9128 9172
rect 9180 9120 9186 9172
rect 9493 9163 9551 9169
rect 9493 9129 9505 9163
rect 9539 9160 9551 9163
rect 11606 9160 11612 9172
rect 9539 9132 11612 9160
rect 9539 9129 9551 9132
rect 9493 9123 9551 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 12158 9120 12164 9172
rect 12216 9120 12222 9172
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 2746 9064 3801 9092
rect 3789 9061 3801 9064
rect 3835 9092 3847 9095
rect 7558 9092 7564 9104
rect 3835 9064 7564 9092
rect 3835 9061 3847 9064
rect 3789 9055 3847 9061
rect 7558 9052 7564 9064
rect 7616 9052 7622 9104
rect 8478 9092 8484 9104
rect 7668 9064 8484 9092
rect 1857 9027 1915 9033
rect 1857 8993 1869 9027
rect 1903 9024 1915 9027
rect 2222 9024 2228 9036
rect 1903 8996 2228 9024
rect 1903 8993 1915 8996
rect 1857 8987 1915 8993
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 4249 9027 4307 9033
rect 4249 9024 4261 9027
rect 2924 8996 4261 9024
rect 2924 8984 2930 8996
rect 4249 8993 4261 8996
rect 4295 8993 4307 9027
rect 4249 8987 4307 8993
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 4157 8959 4215 8965
rect 4157 8956 4169 8959
rect 3200 8928 4169 8956
rect 3200 8916 3206 8928
rect 4157 8925 4169 8928
rect 4203 8925 4215 8959
rect 4264 8956 4292 8987
rect 4341 8959 4399 8965
rect 4341 8956 4353 8959
rect 4264 8928 4353 8956
rect 4157 8919 4215 8925
rect 4341 8925 4353 8928
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4172 8888 4200 8919
rect 4632 8888 4660 8987
rect 4172 8860 4660 8888
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2317 8823 2375 8829
rect 2317 8820 2329 8823
rect 2280 8792 2329 8820
rect 2280 8780 2286 8792
rect 2317 8789 2329 8792
rect 2363 8789 2375 8823
rect 2317 8783 2375 8789
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4212 8792 4537 8820
rect 4212 8780 4218 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4525 8783 4583 8789
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 4724 8820 4752 8987
rect 4890 8984 4896 9036
rect 4948 8984 4954 9036
rect 5629 9027 5687 9033
rect 5629 8993 5641 9027
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5644 8956 5672 8987
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6273 9027 6331 9033
rect 6273 9024 6285 9027
rect 5960 8996 6285 9024
rect 5960 8984 5966 8996
rect 6273 8993 6285 8996
rect 6319 8993 6331 9027
rect 6273 8987 6331 8993
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 6549 9027 6607 9033
rect 6549 9024 6561 9027
rect 6512 8996 6561 9024
rect 6512 8984 6518 8996
rect 6549 8993 6561 8996
rect 6595 8993 6607 9027
rect 6549 8987 6607 8993
rect 6733 9027 6791 9033
rect 6733 8993 6745 9027
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5644 8928 5825 8956
rect 5813 8925 5825 8928
rect 5859 8925 5871 8959
rect 6748 8956 6776 8987
rect 6822 8984 6828 9036
rect 6880 8984 6886 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 7668 9024 7696 9064
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 8754 9052 8760 9104
rect 8812 9052 8818 9104
rect 9674 9092 9680 9104
rect 9324 9064 9680 9092
rect 9324 9033 9352 9064
rect 9674 9052 9680 9064
rect 9732 9052 9738 9104
rect 9769 9095 9827 9101
rect 9769 9061 9781 9095
rect 9815 9092 9827 9095
rect 10042 9092 10048 9104
rect 9815 9064 10048 9092
rect 9815 9061 9827 9064
rect 9769 9055 9827 9061
rect 7055 8996 7696 9024
rect 7929 9027 7987 9033
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7929 8993 7941 9027
rect 7975 9024 7987 9027
rect 9309 9027 9367 9033
rect 7975 8996 8524 9024
rect 7975 8993 7987 8996
rect 7929 8987 7987 8993
rect 6914 8956 6920 8968
rect 6748 8928 6920 8956
rect 5813 8919 5871 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8067 8928 8432 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 5552 8888 5580 8916
rect 5905 8891 5963 8897
rect 5905 8888 5917 8891
rect 5552 8860 5917 8888
rect 5905 8857 5917 8860
rect 5951 8857 5963 8891
rect 7208 8888 7236 8919
rect 7282 8888 7288 8900
rect 7208 8860 7288 8888
rect 5905 8851 5963 8857
rect 7282 8848 7288 8860
rect 7340 8888 7346 8900
rect 8202 8888 8208 8900
rect 7340 8860 8208 8888
rect 7340 8848 7346 8860
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 4672 8792 4752 8820
rect 4672 8780 4678 8792
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 5537 8823 5595 8829
rect 5537 8789 5549 8823
rect 5583 8820 5595 8823
rect 6362 8820 6368 8832
rect 5583 8792 6368 8820
rect 5583 8789 5595 8792
rect 5537 8783 5595 8789
rect 6362 8780 6368 8792
rect 6420 8780 6426 8832
rect 8294 8780 8300 8832
rect 8352 8780 8358 8832
rect 8404 8820 8432 8928
rect 8496 8897 8524 8996
rect 9309 8993 9321 9027
rect 9355 8993 9367 9027
rect 9309 8987 9367 8993
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9585 9027 9643 9033
rect 9585 9024 9597 9027
rect 9548 8996 9597 9024
rect 9548 8984 9554 8996
rect 9585 8993 9597 8996
rect 9631 8993 9643 9027
rect 9585 8987 9643 8993
rect 9784 8956 9812 9055
rect 10042 9052 10048 9064
rect 10100 9092 10106 9104
rect 12434 9092 12440 9104
rect 10100 9064 10548 9092
rect 10100 9052 10106 9064
rect 9950 8984 9956 9036
rect 10008 8984 10014 9036
rect 10410 8984 10416 9036
rect 10468 8984 10474 9036
rect 9508 8928 9812 8956
rect 10520 8956 10548 9064
rect 10612 9064 12440 9092
rect 10612 9033 10640 9064
rect 10597 9027 10655 9033
rect 10597 8993 10609 9027
rect 10643 8993 10655 9027
rect 11149 9027 11207 9033
rect 11149 9024 11161 9027
rect 10597 8987 10655 8993
rect 10704 8996 11161 9024
rect 10704 8968 10732 8996
rect 11149 8993 11161 8996
rect 11195 8993 11207 9027
rect 11149 8987 11207 8993
rect 10520 8928 10640 8956
rect 9508 8900 9536 8928
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 9030 8888 9036 8900
rect 8527 8860 9036 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 9030 8848 9036 8860
rect 9088 8848 9094 8900
rect 9490 8848 9496 8900
rect 9548 8848 9554 8900
rect 10042 8888 10048 8900
rect 9692 8860 10048 8888
rect 8754 8820 8760 8832
rect 8404 8792 8760 8820
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9692 8820 9720 8860
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 10137 8891 10195 8897
rect 10137 8857 10149 8891
rect 10183 8888 10195 8891
rect 10502 8888 10508 8900
rect 10183 8860 10508 8888
rect 10183 8857 10195 8860
rect 10137 8851 10195 8857
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 10612 8888 10640 8928
rect 10686 8916 10692 8968
rect 10744 8916 10750 8968
rect 11256 8965 11284 9064
rect 12434 9052 12440 9064
rect 12492 9052 12498 9104
rect 11422 8984 11428 9036
rect 11480 9024 11486 9036
rect 11609 9027 11667 9033
rect 11609 9024 11621 9027
rect 11480 8996 11621 9024
rect 11480 8984 11486 8996
rect 11609 8993 11621 8996
rect 11655 8993 11667 9027
rect 11609 8987 11667 8993
rect 11793 9027 11851 9033
rect 11793 8993 11805 9027
rect 11839 9024 11851 9027
rect 11974 9024 11980 9036
rect 11839 8996 11980 9024
rect 11839 8993 11851 8996
rect 11793 8987 11851 8993
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12066 8984 12072 9036
rect 12124 8984 12130 9036
rect 12253 9027 12311 9033
rect 12253 8993 12265 9027
rect 12299 8993 12311 9027
rect 12253 8987 12311 8993
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 12268 8956 12296 8987
rect 11241 8919 11299 8925
rect 11992 8928 12296 8956
rect 10962 8888 10968 8900
rect 10612 8860 10968 8888
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 11517 8891 11575 8897
rect 11517 8888 11529 8891
rect 11112 8860 11529 8888
rect 11112 8848 11118 8860
rect 11517 8857 11529 8860
rect 11563 8857 11575 8891
rect 11517 8851 11575 8857
rect 9640 8792 9720 8820
rect 9640 8780 9646 8792
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10229 8823 10287 8829
rect 10229 8820 10241 8823
rect 10008 8792 10241 8820
rect 10008 8780 10014 8792
rect 10229 8789 10241 8792
rect 10275 8789 10287 8823
rect 10229 8783 10287 8789
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 11992 8829 12020 8928
rect 11977 8823 12035 8829
rect 11977 8820 11989 8823
rect 11756 8792 11989 8820
rect 11756 8780 11762 8792
rect 11977 8789 11989 8792
rect 12023 8789 12035 8823
rect 11977 8783 12035 8789
rect 552 8730 12604 8752
rect 552 8678 3662 8730
rect 3714 8678 3726 8730
rect 3778 8678 3790 8730
rect 3842 8678 3854 8730
rect 3906 8678 3918 8730
rect 3970 8678 10062 8730
rect 10114 8678 10126 8730
rect 10178 8678 10190 8730
rect 10242 8678 10254 8730
rect 10306 8678 10318 8730
rect 10370 8678 12604 8730
rect 552 8656 12604 8678
rect 2409 8619 2467 8625
rect 2409 8585 2421 8619
rect 2455 8616 2467 8619
rect 3142 8616 3148 8628
rect 2455 8588 3148 8616
rect 2455 8585 2467 8588
rect 2409 8579 2467 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 3234 8576 3240 8628
rect 3292 8576 3298 8628
rect 5534 8576 5540 8628
rect 5592 8576 5598 8628
rect 6638 8576 6644 8628
rect 6696 8576 6702 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8478 8616 8484 8628
rect 7791 8588 8484 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 10597 8619 10655 8625
rect 8588 8588 9628 8616
rect 3053 8551 3111 8557
rect 3053 8517 3065 8551
rect 3099 8548 3111 8551
rect 4341 8551 4399 8557
rect 4341 8548 4353 8551
rect 3099 8520 4353 8548
rect 3099 8517 3111 8520
rect 3053 8511 3111 8517
rect 4341 8517 4353 8520
rect 4387 8548 4399 8551
rect 4890 8548 4896 8560
rect 4387 8520 4896 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 4890 8508 4896 8520
rect 4948 8508 4954 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 5184 8520 6561 8548
rect 2590 8440 2596 8492
rect 2648 8440 2654 8492
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 4798 8480 4804 8492
rect 3927 8452 4804 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 4798 8440 4804 8452
rect 4856 8440 4862 8492
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 1581 8415 1639 8421
rect 1581 8412 1593 8415
rect 1452 8384 1593 8412
rect 1452 8372 1458 8384
rect 1581 8381 1593 8384
rect 1627 8381 1639 8415
rect 1581 8375 1639 8381
rect 1762 8372 1768 8424
rect 1820 8372 1826 8424
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 2225 8415 2283 8421
rect 2225 8381 2237 8415
rect 2271 8412 2283 8415
rect 2314 8412 2320 8424
rect 2271 8384 2320 8412
rect 2271 8381 2283 8384
rect 2225 8375 2283 8381
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 2409 8415 2467 8421
rect 2409 8381 2421 8415
rect 2455 8412 2467 8415
rect 2498 8412 2504 8424
rect 2455 8384 2504 8412
rect 2455 8381 2467 8384
rect 2409 8375 2467 8381
rect 2498 8372 2504 8384
rect 2556 8372 2562 8424
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 3326 8412 3332 8424
rect 2731 8384 3332 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 3602 8412 3608 8424
rect 3559 8384 3608 8412
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8412 3847 8415
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3835 8384 3985 8412
rect 3835 8381 3847 8384
rect 3789 8375 3847 8381
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4062 8372 4068 8424
rect 4120 8412 4126 8424
rect 4157 8415 4215 8421
rect 4157 8412 4169 8415
rect 4120 8384 4169 8412
rect 4120 8372 4126 8384
rect 4157 8381 4169 8384
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 1118 8304 1124 8356
rect 1176 8304 1182 8356
rect 2516 8344 2544 8372
rect 3050 8344 3056 8356
rect 2516 8316 3056 8344
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 4448 8344 4476 8375
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 4890 8412 4896 8424
rect 4580 8384 4896 8412
rect 4580 8372 4586 8384
rect 4890 8372 4896 8384
rect 4948 8372 4954 8424
rect 5184 8421 5212 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 5718 8480 5724 8492
rect 5276 8452 5724 8480
rect 5276 8421 5304 8452
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6457 8483 6515 8489
rect 6457 8480 6469 8483
rect 6380 8452 6469 8480
rect 6380 8424 6408 8452
rect 6457 8449 6469 8452
rect 6503 8449 6515 8483
rect 6457 8443 6515 8449
rect 4985 8415 5043 8421
rect 4985 8381 4997 8415
rect 5031 8381 5043 8415
rect 4985 8375 5043 8381
rect 5169 8415 5227 8421
rect 5169 8381 5181 8415
rect 5215 8381 5227 8415
rect 5169 8375 5227 8381
rect 5261 8415 5319 8421
rect 5261 8381 5273 8415
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 4614 8344 4620 8356
rect 4448 8316 4620 8344
rect 4614 8304 4620 8316
rect 4672 8344 4678 8356
rect 4798 8344 4804 8356
rect 4672 8316 4804 8344
rect 4672 8304 4678 8316
rect 4798 8304 4804 8316
rect 4856 8304 4862 8356
rect 5000 8344 5028 8375
rect 5350 8372 5356 8424
rect 5408 8372 5414 8424
rect 5813 8415 5871 8421
rect 5813 8381 5825 8415
rect 5859 8412 5871 8415
rect 5997 8415 6055 8421
rect 5859 8384 5948 8412
rect 5859 8381 5871 8384
rect 5813 8375 5871 8381
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5000 8316 5212 8344
rect 5184 8276 5212 8316
rect 5368 8316 5641 8344
rect 5368 8276 5396 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 5629 8307 5687 8313
rect 5184 8248 5396 8276
rect 5920 8276 5948 8384
rect 5997 8381 6009 8415
rect 6043 8381 6055 8415
rect 5997 8375 6055 8381
rect 6012 8344 6040 8375
rect 6086 8372 6092 8424
rect 6144 8372 6150 8424
rect 6178 8372 6184 8424
rect 6236 8372 6242 8424
rect 6362 8372 6368 8424
rect 6420 8372 6426 8424
rect 6656 8344 6684 8576
rect 8588 8548 8616 8588
rect 8496 8520 8616 8548
rect 7006 8440 7012 8492
rect 7064 8480 7070 8492
rect 7558 8480 7564 8492
rect 7064 8452 7564 8480
rect 7064 8440 7070 8452
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 6730 8372 6736 8424
rect 6788 8372 6794 8424
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7469 8415 7527 8421
rect 7469 8412 7481 8415
rect 7340 8384 7481 8412
rect 7340 8372 7346 8384
rect 7469 8381 7481 8384
rect 7515 8381 7527 8415
rect 7469 8375 7527 8381
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8294 8412 8300 8424
rect 7791 8384 8300 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 6012 8316 6684 8344
rect 6748 8276 6776 8372
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 8496 8344 8524 8520
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 9490 8548 9496 8560
rect 8720 8520 9496 8548
rect 8720 8508 8726 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 9600 8548 9628 8588
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 10686 8616 10692 8628
rect 10643 8588 10692 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11241 8619 11299 8625
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11330 8616 11336 8628
rect 11287 8588 11336 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11330 8576 11336 8588
rect 11388 8576 11394 8628
rect 11606 8576 11612 8628
rect 11664 8576 11670 8628
rect 9858 8548 9864 8560
rect 9600 8520 9864 8548
rect 9858 8508 9864 8520
rect 9916 8548 9922 8560
rect 11425 8551 11483 8557
rect 9916 8520 10824 8548
rect 9916 8508 9922 8520
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 8904 8452 9352 8480
rect 8904 8440 8910 8452
rect 9030 8372 9036 8424
rect 9088 8372 9094 8424
rect 9324 8421 9352 8452
rect 10410 8440 10416 8492
rect 10468 8480 10474 8492
rect 10796 8480 10824 8520
rect 11425 8517 11437 8551
rect 11471 8548 11483 8551
rect 12158 8548 12164 8560
rect 11471 8520 12164 8548
rect 11471 8517 11483 8520
rect 11425 8511 11483 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 11330 8480 11336 8492
rect 10468 8452 10732 8480
rect 10468 8440 10474 8452
rect 9217 8415 9275 8421
rect 9217 8381 9229 8415
rect 9263 8381 9275 8415
rect 9217 8375 9275 8381
rect 9309 8415 9367 8421
rect 9309 8381 9321 8415
rect 9355 8381 9367 8415
rect 9309 8375 9367 8381
rect 7607 8316 8524 8344
rect 9232 8344 9260 8375
rect 9490 8372 9496 8424
rect 9548 8372 9554 8424
rect 10502 8372 10508 8424
rect 10560 8372 10566 8424
rect 10704 8421 10732 8452
rect 10796 8452 11336 8480
rect 10796 8421 10824 8452
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8381 10747 8415
rect 10689 8375 10747 8381
rect 10781 8415 10839 8421
rect 10781 8381 10793 8415
rect 10827 8381 10839 8415
rect 10781 8375 10839 8381
rect 9398 8344 9404 8356
rect 9232 8316 9404 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 9398 8304 9404 8316
rect 9456 8304 9462 8356
rect 5920 8248 6776 8276
rect 9214 8236 9220 8288
rect 9272 8236 9278 8288
rect 10704 8276 10732 8375
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 11974 8412 11980 8424
rect 11716 8384 11980 8412
rect 11057 8347 11115 8353
rect 11057 8313 11069 8347
rect 11103 8344 11115 8347
rect 11606 8344 11612 8356
rect 11103 8316 11612 8344
rect 11103 8313 11115 8316
rect 11057 8307 11115 8313
rect 11606 8304 11612 8316
rect 11664 8304 11670 8356
rect 10781 8279 10839 8285
rect 10781 8276 10793 8279
rect 10704 8248 10793 8276
rect 10781 8245 10793 8248
rect 10827 8245 10839 8279
rect 10781 8239 10839 8245
rect 11267 8279 11325 8285
rect 11267 8245 11279 8279
rect 11313 8276 11325 8279
rect 11716 8276 11744 8384
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 11882 8304 11888 8356
rect 11940 8304 11946 8356
rect 11313 8248 11744 8276
rect 11313 8245 11325 8248
rect 11267 8239 11325 8245
rect 552 8186 12604 8208
rect 552 8134 4322 8186
rect 4374 8134 4386 8186
rect 4438 8134 4450 8186
rect 4502 8134 4514 8186
rect 4566 8134 4578 8186
rect 4630 8134 10722 8186
rect 10774 8134 10786 8186
rect 10838 8134 10850 8186
rect 10902 8134 10914 8186
rect 10966 8134 10978 8186
rect 11030 8134 12604 8186
rect 552 8112 12604 8134
rect 845 8075 903 8081
rect 845 8041 857 8075
rect 891 8072 903 8075
rect 1854 8072 1860 8084
rect 891 8044 1860 8072
rect 891 8041 903 8044
rect 845 8035 903 8041
rect 1854 8032 1860 8044
rect 1912 8032 1918 8084
rect 2317 8075 2375 8081
rect 2317 8041 2329 8075
rect 2363 8072 2375 8075
rect 2406 8072 2412 8084
rect 2363 8044 2412 8072
rect 2363 8041 2375 8044
rect 2317 8035 2375 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 3973 8075 4031 8081
rect 3973 8072 3985 8075
rect 3660 8044 3985 8072
rect 3660 8032 3666 8044
rect 3973 8041 3985 8044
rect 4019 8072 4031 8075
rect 4430 8072 4436 8084
rect 4019 8044 4436 8072
rect 4019 8041 4031 8044
rect 3973 8035 4031 8041
rect 4430 8032 4436 8044
rect 4488 8072 4494 8084
rect 5074 8072 5080 8084
rect 4488 8044 5080 8072
rect 4488 8032 4494 8044
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5350 8072 5356 8084
rect 5307 8044 5356 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 6178 8032 6184 8084
rect 6236 8032 6242 8084
rect 7374 8072 7380 8084
rect 7116 8044 7380 8072
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 1958 8007 2016 8013
rect 1958 8004 1970 8007
rect 1820 7976 1970 8004
rect 1820 7964 1826 7976
rect 1958 7973 1970 7976
rect 2004 7973 2016 8007
rect 1958 7967 2016 7973
rect 4801 8007 4859 8013
rect 4801 7973 4813 8007
rect 4847 8004 4859 8007
rect 4847 7976 4935 8004
rect 4847 7973 4859 7976
rect 4801 7967 4859 7973
rect 2593 7939 2651 7945
rect 2593 7905 2605 7939
rect 2639 7936 2651 7939
rect 2682 7936 2688 7948
rect 2639 7908 2688 7936
rect 2639 7905 2651 7908
rect 2593 7899 2651 7905
rect 2682 7896 2688 7908
rect 2740 7896 2746 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 3050 7936 3056 7948
rect 2832 7908 3056 7936
rect 2832 7896 2838 7908
rect 3050 7896 3056 7908
rect 3108 7936 3114 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 3108 7908 3157 7936
rect 3108 7896 3114 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 3145 7899 3203 7905
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4522 7936 4528 7948
rect 4295 7908 4528 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 4709 7939 4767 7945
rect 4709 7905 4721 7939
rect 4755 7905 4767 7939
rect 4907 7936 4935 7976
rect 4995 7939 5053 7945
rect 4907 7908 4937 7936
rect 4709 7899 4767 7905
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2406 7868 2412 7880
rect 2363 7840 2412 7868
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2866 7828 2872 7880
rect 2924 7868 2930 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 2924 7840 3249 7868
rect 2924 7828 2930 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 3237 7831 3295 7837
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4157 7871 4215 7877
rect 4157 7868 4169 7871
rect 3384 7840 4169 7868
rect 3384 7828 3390 7840
rect 4157 7837 4169 7840
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 4724 7800 4752 7899
rect 4488 7772 4752 7800
rect 4909 7800 4937 7908
rect 4995 7905 5007 7939
rect 5041 7936 5053 7939
rect 5350 7936 5356 7948
rect 5041 7908 5356 7936
rect 5041 7905 5053 7908
rect 4995 7899 5053 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 5445 7939 5503 7945
rect 5445 7905 5457 7939
rect 5491 7905 5503 7939
rect 5445 7899 5503 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7936 5687 7939
rect 5902 7936 5908 7948
rect 5675 7908 5908 7936
rect 5675 7905 5687 7908
rect 5629 7899 5687 7905
rect 5460 7868 5488 7899
rect 5902 7896 5908 7908
rect 5960 7936 5966 7948
rect 5997 7939 6055 7945
rect 5997 7936 6009 7939
rect 5960 7908 6009 7936
rect 5960 7896 5966 7908
rect 5997 7905 6009 7908
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 7006 7896 7012 7948
rect 7064 7936 7070 7948
rect 7116 7945 7144 8044
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9030 8072 9036 8084
rect 8803 8044 9036 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 9490 8032 9496 8084
rect 9548 8032 9554 8084
rect 8018 7964 8024 8016
rect 8076 8004 8082 8016
rect 8573 8007 8631 8013
rect 8573 8004 8585 8007
rect 8076 7976 8585 8004
rect 8076 7964 8082 7976
rect 8573 7973 8585 7976
rect 8619 8004 8631 8007
rect 8846 8004 8852 8016
rect 8619 7976 8852 8004
rect 8619 7973 8631 7976
rect 8573 7967 8631 7973
rect 8846 7964 8852 7976
rect 8904 8004 8910 8016
rect 10137 8007 10195 8013
rect 10137 8004 10149 8007
rect 8904 7976 10149 8004
rect 8904 7964 8910 7976
rect 10137 7973 10149 7976
rect 10183 7973 10195 8007
rect 10137 7967 10195 7973
rect 10318 7964 10324 8016
rect 10376 7964 10382 8016
rect 11885 8007 11943 8013
rect 11885 7973 11897 8007
rect 11931 7973 11943 8007
rect 11885 7967 11943 7973
rect 7101 7939 7159 7945
rect 7101 7936 7113 7939
rect 7064 7908 7113 7936
rect 7064 7896 7070 7908
rect 7101 7905 7113 7908
rect 7147 7905 7159 7939
rect 7101 7899 7159 7905
rect 7282 7896 7288 7948
rect 7340 7896 7346 7948
rect 7374 7896 7380 7948
rect 7432 7896 7438 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8662 7936 8668 7948
rect 8435 7908 8668 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 9033 7939 9091 7945
rect 9033 7905 9045 7939
rect 9079 7936 9091 7939
rect 9214 7936 9220 7948
rect 9079 7908 9220 7936
rect 9079 7905 9091 7908
rect 9033 7899 9091 7905
rect 9214 7896 9220 7908
rect 9272 7896 9278 7948
rect 9858 7896 9864 7948
rect 9916 7896 9922 7948
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7936 11207 7939
rect 11238 7936 11244 7948
rect 11195 7908 11244 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 11238 7896 11244 7908
rect 11296 7896 11302 7948
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 11698 7896 11704 7948
rect 11756 7896 11762 7948
rect 11900 7936 11928 7967
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11900 7908 11989 7936
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 12158 7896 12164 7948
rect 12216 7896 12222 7948
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5460 7840 5825 7868
rect 5166 7800 5172 7812
rect 4909 7772 5172 7800
rect 4488 7760 4494 7772
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 2774 7732 2780 7744
rect 2547 7704 2780 7732
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 4614 7692 4620 7744
rect 4672 7692 4678 7744
rect 4985 7735 5043 7741
rect 4985 7701 4997 7735
rect 5031 7732 5043 7735
rect 5460 7732 5488 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 9122 7828 9128 7880
rect 9180 7828 9186 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9447 7840 9781 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 9769 7831 9827 7837
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7868 11943 7871
rect 12250 7868 12256 7880
rect 11931 7840 12256 7868
rect 11931 7837 11943 7840
rect 11885 7831 11943 7837
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 6638 7760 6644 7812
rect 6696 7800 6702 7812
rect 7190 7800 7196 7812
rect 6696 7772 7196 7800
rect 6696 7760 6702 7772
rect 7190 7760 7196 7772
rect 7248 7760 7254 7812
rect 5626 7732 5632 7744
rect 5031 7704 5632 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 6914 7692 6920 7744
rect 6972 7692 6978 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10318 7732 10324 7744
rect 9548 7704 10324 7732
rect 9548 7692 9554 7704
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 11974 7692 11980 7744
rect 12032 7692 12038 7744
rect 552 7642 12604 7664
rect 552 7590 3662 7642
rect 3714 7590 3726 7642
rect 3778 7590 3790 7642
rect 3842 7590 3854 7642
rect 3906 7590 3918 7642
rect 3970 7590 10062 7642
rect 10114 7590 10126 7642
rect 10178 7590 10190 7642
rect 10242 7590 10254 7642
rect 10306 7590 10318 7642
rect 10370 7590 12604 7642
rect 552 7568 12604 7590
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 2774 7488 2780 7540
rect 2832 7488 2838 7540
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4580 7500 6592 7528
rect 4580 7488 4586 7500
rect 3050 7420 3056 7472
rect 3108 7460 3114 7472
rect 4893 7463 4951 7469
rect 4893 7460 4905 7463
rect 3108 7432 4905 7460
rect 3108 7420 3114 7432
rect 4893 7429 4905 7432
rect 4939 7429 4951 7463
rect 4893 7423 4951 7429
rect 5077 7463 5135 7469
rect 5077 7429 5089 7463
rect 5123 7460 5135 7463
rect 5350 7460 5356 7472
rect 5123 7432 5356 7460
rect 5123 7429 5135 7432
rect 5077 7423 5135 7429
rect 5350 7420 5356 7432
rect 5408 7420 5414 7472
rect 5537 7463 5595 7469
rect 5537 7429 5549 7463
rect 5583 7460 5595 7463
rect 6086 7460 6092 7472
rect 5583 7432 6092 7460
rect 5583 7429 5595 7432
rect 5537 7423 5595 7429
rect 6086 7420 6092 7432
rect 6144 7420 6150 7472
rect 2516 7364 2820 7392
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 2222 7324 2228 7336
rect 1544 7296 2228 7324
rect 1544 7284 1550 7296
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2314 7284 2320 7336
rect 2372 7284 2378 7336
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2516 7333 2544 7364
rect 2792 7333 2820 7364
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3142 7392 3148 7404
rect 2924 7364 3148 7392
rect 2924 7352 2930 7364
rect 3142 7352 3148 7364
rect 3200 7392 3206 7404
rect 4617 7395 4675 7401
rect 4617 7392 4629 7395
rect 3200 7364 4629 7392
rect 3200 7352 3206 7364
rect 4617 7361 4629 7364
rect 4663 7361 4675 7395
rect 5902 7392 5908 7404
rect 4617 7355 4675 7361
rect 5276 7364 5908 7392
rect 2501 7327 2559 7333
rect 2501 7324 2513 7327
rect 2464 7296 2513 7324
rect 2464 7284 2470 7296
rect 2501 7293 2513 7296
rect 2547 7293 2559 7327
rect 2501 7287 2559 7293
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7293 2651 7327
rect 2593 7287 2651 7293
rect 2777 7327 2835 7333
rect 2777 7293 2789 7327
rect 2823 7324 2835 7327
rect 2958 7324 2964 7336
rect 2823 7296 2964 7324
rect 2823 7293 2835 7296
rect 2777 7287 2835 7293
rect 1980 7259 2038 7265
rect 1980 7225 1992 7259
rect 2026 7256 2038 7259
rect 2130 7256 2136 7268
rect 2026 7228 2136 7256
rect 2026 7225 2038 7228
rect 1980 7219 2038 7225
rect 2130 7216 2136 7228
rect 2188 7216 2194 7268
rect 2332 7256 2360 7284
rect 2608 7256 2636 7287
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 5276 7324 5304 7364
rect 5552 7333 5580 7364
rect 4632 7296 5304 7324
rect 5353 7327 5411 7333
rect 4632 7268 4660 7296
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5353 7287 5411 7293
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7293 5595 7327
rect 5537 7287 5595 7293
rect 2332 7228 2636 7256
rect 4614 7216 4620 7268
rect 4672 7216 4678 7268
rect 5368 7256 5396 7287
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5828 7333 5856 7364
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 6564 7336 6592 7500
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 7285 7531 7343 7537
rect 7285 7528 7297 7531
rect 7156 7500 7297 7528
rect 7156 7488 7162 7500
rect 7285 7497 7297 7500
rect 7331 7497 7343 7531
rect 7285 7491 7343 7497
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 9858 7528 9864 7540
rect 8987 7500 9864 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 11882 7488 11888 7540
rect 11940 7528 11946 7540
rect 12253 7531 12311 7537
rect 12253 7528 12265 7531
rect 11940 7500 12265 7528
rect 11940 7488 11946 7500
rect 12253 7497 12265 7500
rect 12299 7497 12311 7531
rect 12253 7491 12311 7497
rect 9122 7420 9128 7472
rect 9180 7420 9186 7472
rect 7466 7392 7472 7404
rect 6840 7364 7472 7392
rect 5813 7327 5871 7333
rect 5813 7293 5825 7327
rect 5859 7293 5871 7327
rect 5813 7287 5871 7293
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 6052 7296 6377 7324
rect 6052 7284 6058 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6546 7284 6552 7336
rect 6604 7284 6610 7336
rect 6638 7284 6644 7336
rect 6696 7284 6702 7336
rect 6840 7333 6868 7364
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7392 8263 7395
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 8251 7364 8677 7392
rect 8251 7361 8263 7364
rect 8205 7355 8263 7361
rect 8665 7361 8677 7364
rect 8711 7392 8723 7395
rect 8846 7392 8852 7404
rect 8711 7364 8852 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 6825 7327 6883 7333
rect 6825 7293 6837 7327
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6914 7284 6920 7336
rect 6972 7284 6978 7336
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7324 7067 7327
rect 7190 7324 7196 7336
rect 7055 7296 7196 7324
rect 7055 7293 7067 7296
rect 7009 7287 7067 7293
rect 7190 7284 7196 7296
rect 7248 7284 7254 7336
rect 7837 7327 7895 7333
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7944 7324 7972 7355
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 9214 7392 9220 7404
rect 9048 7364 9220 7392
rect 8478 7324 8484 7336
rect 7944 7296 8484 7324
rect 7837 7287 7895 7293
rect 5644 7256 5672 7284
rect 5368 7228 5672 7256
rect 5718 7216 5724 7268
rect 5776 7216 5782 7268
rect 7852 7256 7880 7287
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8570 7284 8576 7336
rect 8628 7284 8634 7336
rect 9048 7333 9076 7364
rect 9214 7352 9220 7364
rect 9272 7352 9278 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9398 7392 9404 7404
rect 9355 7364 9404 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 10594 7352 10600 7404
rect 10652 7392 10658 7404
rect 10873 7395 10931 7401
rect 10873 7392 10885 7395
rect 10652 7364 10885 7392
rect 10652 7352 10658 7364
rect 10873 7361 10885 7364
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 11140 7327 11198 7333
rect 11140 7293 11152 7327
rect 11186 7324 11198 7327
rect 11974 7324 11980 7336
rect 11186 7296 11980 7324
rect 11186 7293 11198 7296
rect 11140 7287 11198 7293
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 8018 7256 8024 7268
rect 6472 7228 8024 7256
rect 845 7191 903 7197
rect 845 7157 857 7191
rect 891 7188 903 7191
rect 1670 7188 1676 7200
rect 891 7160 1676 7188
rect 891 7157 903 7160
rect 845 7151 903 7157
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 6472 7188 6500 7228
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 5224 7160 6500 7188
rect 6549 7191 6607 7197
rect 5224 7148 5230 7160
rect 6549 7157 6561 7191
rect 6595 7188 6607 7191
rect 6914 7188 6920 7200
rect 6595 7160 6920 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 9306 7148 9312 7200
rect 9364 7148 9370 7200
rect 552 7098 12604 7120
rect 552 7046 4322 7098
rect 4374 7046 4386 7098
rect 4438 7046 4450 7098
rect 4502 7046 4514 7098
rect 4566 7046 4578 7098
rect 4630 7046 10722 7098
rect 10774 7046 10786 7098
rect 10838 7046 10850 7098
rect 10902 7046 10914 7098
rect 10966 7046 10978 7098
rect 11030 7046 12604 7098
rect 552 7024 12604 7046
rect 1946 6944 1952 6996
rect 2004 6984 2010 6996
rect 2406 6984 2412 6996
rect 2004 6956 2412 6984
rect 2004 6944 2010 6956
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 4890 6984 4896 6996
rect 4448 6956 4896 6984
rect 2130 6916 2136 6928
rect 1596 6888 2136 6916
rect 1394 6808 1400 6860
rect 1452 6808 1458 6860
rect 1596 6857 1624 6888
rect 2130 6876 2136 6888
rect 2188 6876 2194 6928
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6817 1639 6851
rect 1581 6811 1639 6817
rect 1670 6808 1676 6860
rect 1728 6808 1734 6860
rect 2314 6808 2320 6860
rect 2372 6808 2378 6860
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6817 3111 6851
rect 3053 6811 3111 6817
rect 3973 6851 4031 6857
rect 3973 6817 3985 6851
rect 4019 6817 4031 6851
rect 3973 6811 4031 6817
rect 4065 6851 4123 6857
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6848 4215 6851
rect 4246 6848 4252 6860
rect 4203 6820 4252 6848
rect 4203 6817 4215 6820
rect 4157 6811 4215 6817
rect 934 6740 940 6792
rect 992 6740 998 6792
rect 2038 6740 2044 6792
rect 2096 6740 2102 6792
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 3068 6780 3096 6811
rect 2188 6752 3096 6780
rect 2188 6740 2194 6752
rect 3510 6740 3516 6792
rect 3568 6780 3574 6792
rect 3697 6783 3755 6789
rect 3697 6780 3709 6783
rect 3568 6752 3709 6780
rect 3568 6740 3574 6752
rect 3697 6749 3709 6752
rect 3743 6749 3755 6783
rect 3697 6743 3755 6749
rect 1854 6672 1860 6724
rect 1912 6712 1918 6724
rect 2225 6715 2283 6721
rect 2225 6712 2237 6715
rect 1912 6684 2237 6712
rect 1912 6672 1918 6684
rect 2225 6681 2237 6684
rect 2271 6681 2283 6715
rect 2225 6675 2283 6681
rect 1026 6604 1032 6656
rect 1084 6644 1090 6656
rect 2133 6647 2191 6653
rect 2133 6644 2145 6647
rect 1084 6616 2145 6644
rect 1084 6604 1090 6616
rect 2133 6613 2145 6616
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3050 6644 3056 6656
rect 3007 6616 3056 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3988 6644 4016 6811
rect 4080 6712 4108 6811
rect 4246 6808 4252 6820
rect 4304 6808 4310 6860
rect 4448 6857 4476 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7340 6956 7573 6984
rect 7340 6944 7346 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 8076 6956 8340 6984
rect 8076 6944 8082 6956
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6848 4399 6851
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4387 6820 4445 6848
rect 4387 6817 4399 6820
rect 4341 6811 4399 6817
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4614 6808 4620 6860
rect 4672 6808 4678 6860
rect 4706 6808 4712 6860
rect 4764 6808 4770 6860
rect 4801 6851 4859 6857
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 4890 6848 4896 6860
rect 4847 6820 4896 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5166 6808 5172 6860
rect 5224 6848 5230 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5224 6820 5365 6848
rect 5224 6808 5230 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5537 6851 5595 6857
rect 5537 6817 5549 6851
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5077 6783 5135 6789
rect 5077 6749 5089 6783
rect 5123 6780 5135 6783
rect 5442 6780 5448 6792
rect 5123 6752 5448 6780
rect 5123 6749 5135 6752
rect 5077 6743 5135 6749
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5552 6780 5580 6811
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 5736 6820 5948 6848
rect 5736 6780 5764 6820
rect 5920 6792 5948 6820
rect 6086 6808 6092 6860
rect 6144 6808 6150 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 6595 6820 7205 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7193 6817 7205 6820
rect 7239 6848 7251 6851
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7239 6820 7665 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 7834 6808 7840 6860
rect 7892 6808 7898 6860
rect 8312 6857 8340 6956
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8628 6956 8953 6984
rect 8628 6944 8634 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 10689 6987 10747 6993
rect 10689 6953 10701 6987
rect 10735 6984 10747 6987
rect 11238 6984 11244 6996
rect 10735 6956 11244 6984
rect 10735 6953 10747 6956
rect 10689 6947 10747 6953
rect 11238 6944 11244 6956
rect 11296 6944 11302 6996
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 8904 6888 9076 6916
rect 8904 6876 8910 6888
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6817 8355 6851
rect 8297 6811 8355 6817
rect 5552 6752 5764 6780
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 5960 6752 6285 6780
rect 5960 6740 5966 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6457 6783 6515 6789
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6822 6780 6828 6792
rect 6503 6752 6828 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 6914 6740 6920 6792
rect 6972 6740 6978 6792
rect 7006 6740 7012 6792
rect 7064 6780 7070 6792
rect 7101 6783 7159 6789
rect 7101 6780 7113 6783
rect 7064 6752 7113 6780
rect 7064 6740 7070 6752
rect 7101 6749 7113 6752
rect 7147 6749 7159 6783
rect 8128 6780 8156 6811
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 9048 6857 9076 6888
rect 9692 6888 9904 6916
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6848 8723 6851
rect 8757 6851 8815 6857
rect 8757 6848 8769 6851
rect 8711 6820 8769 6848
rect 8711 6817 8723 6820
rect 8665 6811 8723 6817
rect 8757 6817 8769 6820
rect 8803 6817 8815 6851
rect 8757 6811 8815 6817
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6817 9091 6851
rect 9033 6811 9091 6817
rect 9582 6808 9588 6860
rect 9640 6848 9646 6860
rect 9692 6848 9720 6888
rect 9640 6820 9720 6848
rect 9640 6808 9646 6820
rect 8846 6780 8852 6792
rect 8128 6752 8852 6780
rect 7101 6743 7159 6749
rect 8846 6740 8852 6752
rect 8904 6740 8910 6792
rect 4154 6712 4160 6724
rect 4080 6684 4160 6712
rect 4154 6672 4160 6684
rect 4212 6672 4218 6724
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 4798 6712 4804 6724
rect 4580 6684 4804 6712
rect 4580 6672 4586 6684
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5169 6715 5227 6721
rect 5169 6681 5181 6715
rect 5215 6712 5227 6715
rect 5997 6715 6055 6721
rect 5997 6712 6009 6715
rect 5215 6684 6009 6712
rect 5215 6681 5227 6684
rect 5169 6675 5227 6681
rect 5997 6681 6009 6684
rect 6043 6681 6055 6715
rect 5997 6675 6055 6681
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 9692 6712 9720 6820
rect 9766 6808 9772 6860
rect 9824 6808 9830 6860
rect 9876 6848 9904 6888
rect 10704 6888 11376 6916
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9876 6820 10057 6848
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10229 6851 10287 6857
rect 10229 6817 10241 6851
rect 10275 6848 10287 6851
rect 10505 6851 10563 6857
rect 10505 6848 10517 6851
rect 10275 6820 10517 6848
rect 10275 6817 10287 6820
rect 10229 6811 10287 6817
rect 10505 6817 10517 6820
rect 10551 6817 10563 6851
rect 10505 6811 10563 6817
rect 9861 6783 9919 6789
rect 9861 6749 9873 6783
rect 9907 6780 9919 6783
rect 10704 6780 10732 6888
rect 11348 6860 11376 6888
rect 10781 6851 10839 6857
rect 10781 6817 10793 6851
rect 10827 6848 10839 6851
rect 10827 6820 11008 6848
rect 10827 6817 10839 6820
rect 10781 6811 10839 6817
rect 10980 6789 11008 6820
rect 11330 6808 11336 6860
rect 11388 6808 11394 6860
rect 9907 6752 10732 6780
rect 10965 6783 11023 6789
rect 9907 6749 9919 6752
rect 9861 6743 9919 6749
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11054 6780 11060 6792
rect 11011 6752 11060 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 11241 6783 11299 6789
rect 11241 6749 11253 6783
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11256 6712 11284 6743
rect 8536 6684 11284 6712
rect 8536 6672 8542 6684
rect 4614 6644 4620 6656
rect 3988 6616 4620 6644
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5905 6647 5963 6653
rect 5905 6644 5917 6647
rect 5316 6616 5917 6644
rect 5316 6604 5322 6616
rect 5905 6613 5917 6616
rect 5951 6613 5963 6647
rect 5905 6607 5963 6613
rect 8754 6604 8760 6656
rect 8812 6604 8818 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10321 6647 10379 6653
rect 10321 6644 10333 6647
rect 9824 6616 10333 6644
rect 9824 6604 9830 6616
rect 10321 6613 10333 6616
rect 10367 6613 10379 6647
rect 10321 6607 10379 6613
rect 552 6554 12604 6576
rect 552 6502 3662 6554
rect 3714 6502 3726 6554
rect 3778 6502 3790 6554
rect 3842 6502 3854 6554
rect 3906 6502 3918 6554
rect 3970 6502 10062 6554
rect 10114 6502 10126 6554
rect 10178 6502 10190 6554
rect 10242 6502 10254 6554
rect 10306 6502 10318 6554
rect 10370 6502 12604 6554
rect 552 6480 12604 6502
rect 474 6400 480 6452
rect 532 6440 538 6452
rect 532 6412 2176 6440
rect 532 6400 538 6412
rect 845 6239 903 6245
rect 845 6205 857 6239
rect 891 6205 903 6239
rect 845 6199 903 6205
rect 860 6100 888 6199
rect 1026 6196 1032 6248
rect 1084 6196 1090 6248
rect 1121 6239 1179 6245
rect 1121 6205 1133 6239
rect 1167 6236 1179 6239
rect 1167 6208 1532 6236
rect 1167 6205 1179 6208
rect 1121 6199 1179 6205
rect 1504 6180 1532 6208
rect 937 6171 995 6177
rect 937 6137 949 6171
rect 983 6168 995 6171
rect 1366 6171 1424 6177
rect 1366 6168 1378 6171
rect 983 6140 1378 6168
rect 983 6137 995 6140
rect 937 6131 995 6137
rect 1366 6137 1378 6140
rect 1412 6137 1424 6171
rect 1366 6131 1424 6137
rect 1486 6128 1492 6180
rect 1544 6128 1550 6180
rect 2148 6168 2176 6412
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2501 6443 2559 6449
rect 2501 6440 2513 6443
rect 2372 6412 2513 6440
rect 2372 6400 2378 6412
rect 2501 6409 2513 6412
rect 2547 6409 2559 6443
rect 2501 6403 2559 6409
rect 3053 6443 3111 6449
rect 3053 6409 3065 6443
rect 3099 6440 3111 6443
rect 4522 6440 4528 6452
rect 3099 6412 4528 6440
rect 3099 6409 3111 6412
rect 3053 6403 3111 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4617 6443 4675 6449
rect 4617 6409 4629 6443
rect 4663 6440 4675 6443
rect 4706 6440 4712 6452
rect 4663 6412 4712 6440
rect 4663 6409 4675 6412
rect 4617 6403 4675 6409
rect 4706 6400 4712 6412
rect 4764 6400 4770 6452
rect 4890 6400 4896 6452
rect 4948 6400 4954 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 6086 6440 6092 6452
rect 5675 6412 6092 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 6822 6400 6828 6452
rect 6880 6400 6886 6452
rect 7006 6400 7012 6452
rect 7064 6400 7070 6452
rect 7190 6400 7196 6452
rect 7248 6400 7254 6452
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 7892 6412 9505 6440
rect 7892 6400 7898 6412
rect 9493 6409 9505 6412
rect 9539 6440 9551 6443
rect 10134 6440 10140 6452
rect 9539 6412 10140 6440
rect 9539 6409 9551 6412
rect 9493 6403 9551 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10244 6412 10701 6440
rect 5258 6372 5264 6384
rect 3712 6344 5264 6372
rect 3510 6264 3516 6316
rect 3568 6264 3574 6316
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2866 6236 2872 6248
rect 2823 6208 2872 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 2866 6196 2872 6208
rect 2924 6196 2930 6248
rect 3050 6196 3056 6248
rect 3108 6196 3114 6248
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3602 6236 3608 6248
rect 3467 6208 3608 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 3712 6168 3740 6344
rect 5258 6332 5264 6344
rect 5316 6332 5322 6384
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6304 3847 6307
rect 3835 6276 4752 6304
rect 3835 6273 3847 6276
rect 3789 6267 3847 6273
rect 4264 6245 4292 6276
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 4249 6239 4307 6245
rect 4249 6205 4261 6239
rect 4295 6205 4307 6239
rect 4249 6199 4307 6205
rect 2148 6140 3740 6168
rect 4172 6168 4200 6199
rect 4430 6196 4436 6248
rect 4488 6196 4494 6248
rect 4724 6245 4752 6276
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 4709 6199 4767 6205
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 4908 6168 4936 6199
rect 5534 6196 5540 6248
rect 5592 6236 5598 6248
rect 5629 6239 5687 6245
rect 5629 6236 5641 6239
rect 5592 6208 5641 6236
rect 5592 6196 5598 6208
rect 5629 6205 5641 6208
rect 5675 6205 5687 6239
rect 5629 6199 5687 6205
rect 5813 6239 5871 6245
rect 5813 6205 5825 6239
rect 5859 6236 5871 6239
rect 5902 6236 5908 6248
rect 5859 6208 5908 6236
rect 5859 6205 5871 6208
rect 5813 6199 5871 6205
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 5994 6196 6000 6248
rect 6052 6236 6058 6248
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6052 6208 6469 6236
rect 6052 6196 6058 6208
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6604 6208 6653 6236
rect 6604 6196 6610 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6840 6236 6868 6400
rect 10244 6304 10272 6412
rect 10689 6409 10701 6412
rect 10735 6440 10747 6443
rect 11146 6440 11152 6452
rect 10735 6412 11152 6440
rect 10735 6409 10747 6412
rect 10689 6403 10747 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 9784 6276 10272 6304
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6840 6208 6929 6236
rect 6641 6199 6699 6205
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7101 6239 7159 6245
rect 7101 6236 7113 6239
rect 7064 6208 7113 6236
rect 7064 6196 7070 6208
rect 7101 6205 7113 6208
rect 7147 6205 7159 6239
rect 7101 6199 7159 6205
rect 7190 6196 7196 6248
rect 7248 6196 7254 6248
rect 7282 6196 7288 6248
rect 7340 6236 7346 6248
rect 7377 6239 7435 6245
rect 7377 6236 7389 6239
rect 7340 6208 7389 6236
rect 7340 6196 7346 6208
rect 7377 6205 7389 6208
rect 7423 6205 7435 6239
rect 7377 6199 7435 6205
rect 9674 6196 9680 6248
rect 9732 6196 9738 6248
rect 9784 6245 9812 6276
rect 10318 6264 10324 6316
rect 10376 6264 10382 6316
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 9950 6196 9956 6248
rect 10008 6236 10014 6248
rect 10229 6239 10287 6245
rect 10008 6230 10180 6236
rect 10229 6230 10241 6239
rect 10008 6208 10241 6230
rect 10008 6196 10014 6208
rect 10152 6205 10241 6208
rect 10275 6205 10287 6239
rect 10152 6202 10287 6205
rect 10229 6199 10287 6202
rect 4172 6140 4936 6168
rect 9493 6171 9551 6177
rect 4264 6112 4292 6140
rect 9493 6137 9505 6171
rect 9539 6168 9551 6171
rect 10410 6168 10416 6180
rect 9539 6140 10416 6168
rect 9539 6137 9551 6140
rect 9493 6131 9551 6137
rect 10410 6128 10416 6140
rect 10468 6168 10474 6180
rect 10657 6171 10715 6177
rect 10657 6168 10669 6171
rect 10468 6140 10669 6168
rect 10468 6128 10474 6140
rect 10657 6137 10669 6140
rect 10703 6137 10715 6171
rect 10657 6131 10715 6137
rect 10870 6128 10876 6180
rect 10928 6128 10934 6180
rect 492 6072 888 6100
rect 492 5896 520 6072
rect 2682 6060 2688 6112
rect 2740 6100 2746 6112
rect 2869 6103 2927 6109
rect 2869 6100 2881 6103
rect 2740 6072 2881 6100
rect 2740 6060 2746 6072
rect 2869 6069 2881 6072
rect 2915 6100 2927 6103
rect 3602 6100 3608 6112
rect 2915 6072 3608 6100
rect 2915 6069 2927 6072
rect 2869 6063 2927 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 4246 6060 4252 6112
rect 4304 6060 4310 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 4798 6100 4804 6112
rect 4488 6072 4804 6100
rect 4488 6060 4494 6072
rect 4798 6060 4804 6072
rect 4856 6100 4862 6112
rect 5166 6100 5172 6112
rect 4856 6072 5172 6100
rect 4856 6060 4862 6072
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 9861 6103 9919 6109
rect 9861 6100 9873 6103
rect 9640 6072 9873 6100
rect 9640 6060 9646 6072
rect 9861 6069 9873 6072
rect 9907 6069 9919 6103
rect 9861 6063 9919 6069
rect 10318 6060 10324 6112
rect 10376 6100 10382 6112
rect 10505 6103 10563 6109
rect 10505 6100 10517 6103
rect 10376 6072 10517 6100
rect 10376 6060 10382 6072
rect 10505 6069 10517 6072
rect 10551 6069 10563 6103
rect 10505 6063 10563 6069
rect 552 6010 12604 6032
rect 552 5958 4322 6010
rect 4374 5958 4386 6010
rect 4438 5958 4450 6010
rect 4502 5958 4514 6010
rect 4566 5958 4578 6010
rect 4630 5958 10722 6010
rect 10774 5958 10786 6010
rect 10838 5958 10850 6010
rect 10902 5958 10914 6010
rect 10966 5958 10978 6010
rect 11030 5958 12604 6010
rect 552 5936 12604 5958
rect 1673 5899 1731 5905
rect 1673 5896 1685 5899
rect 492 5868 1685 5896
rect 1673 5865 1685 5868
rect 1719 5865 1731 5899
rect 1673 5859 1731 5865
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 2961 5899 3019 5905
rect 2372 5868 2636 5896
rect 2372 5856 2378 5868
rect 2332 5828 2360 5856
rect 2608 5837 2636 5868
rect 2961 5865 2973 5899
rect 3007 5896 3019 5899
rect 3007 5868 3464 5896
rect 3007 5865 3019 5868
rect 2961 5859 3019 5865
rect 2056 5800 2360 5828
rect 2593 5831 2651 5837
rect 1854 5720 1860 5772
rect 1912 5720 1918 5772
rect 2056 5769 2084 5800
rect 2593 5797 2605 5831
rect 2639 5797 2651 5831
rect 2593 5791 2651 5797
rect 2682 5788 2688 5840
rect 2740 5788 2746 5840
rect 3053 5831 3111 5837
rect 3053 5828 3065 5831
rect 2792 5800 3065 5828
rect 2041 5763 2099 5769
rect 2041 5729 2053 5763
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 2133 5763 2191 5769
rect 2133 5729 2145 5763
rect 2179 5729 2191 5763
rect 2133 5723 2191 5729
rect 2317 5763 2375 5769
rect 2317 5729 2329 5763
rect 2363 5729 2375 5763
rect 2317 5723 2375 5729
rect 2148 5556 2176 5723
rect 2332 5692 2360 5723
rect 2406 5720 2412 5772
rect 2464 5760 2470 5772
rect 2501 5763 2559 5769
rect 2501 5760 2513 5763
rect 2464 5732 2513 5760
rect 2464 5720 2470 5732
rect 2501 5729 2513 5732
rect 2547 5729 2559 5763
rect 2501 5723 2559 5729
rect 2792 5692 2820 5800
rect 3053 5797 3065 5800
rect 3099 5828 3111 5831
rect 3142 5828 3148 5840
rect 3099 5800 3148 5828
rect 3099 5797 3111 5800
rect 3053 5791 3111 5797
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 3436 5828 3464 5868
rect 3510 5856 3516 5908
rect 3568 5856 3574 5908
rect 3602 5856 3608 5908
rect 3660 5896 3666 5908
rect 5166 5896 5172 5908
rect 3660 5868 5172 5896
rect 3660 5856 3666 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 9677 5899 9735 5905
rect 9677 5865 9689 5899
rect 9723 5865 9735 5899
rect 9677 5859 9735 5865
rect 4062 5828 4068 5840
rect 3436 5800 4068 5828
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 9692 5828 9720 5859
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 10410 5896 10416 5908
rect 10060 5868 10416 5896
rect 10060 5828 10088 5868
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 9692 5800 10088 5828
rect 10134 5788 10140 5840
rect 10192 5788 10198 5840
rect 10318 5788 10324 5840
rect 10376 5788 10382 5840
rect 2866 5720 2872 5772
rect 2924 5720 2930 5772
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3007 5732 3096 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3068 5704 3096 5732
rect 3234 5720 3240 5772
rect 3292 5720 3298 5772
rect 3418 5720 3424 5772
rect 3476 5720 3482 5772
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5758 3571 5763
rect 3559 5730 3648 5758
rect 3559 5729 3571 5730
rect 3513 5723 3571 5729
rect 2332 5664 2820 5692
rect 3050 5652 3056 5704
rect 3108 5652 3114 5704
rect 2222 5584 2228 5636
rect 2280 5624 2286 5636
rect 3620 5624 3648 5730
rect 3694 5720 3700 5772
rect 3752 5720 3758 5772
rect 9122 5720 9128 5772
rect 9180 5760 9186 5772
rect 9309 5763 9367 5769
rect 9309 5760 9321 5763
rect 9180 5732 9321 5760
rect 9180 5720 9186 5732
rect 9309 5729 9321 5732
rect 9355 5729 9367 5763
rect 9309 5723 9367 5729
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8846 5692 8852 5704
rect 8076 5664 8852 5692
rect 8076 5652 8082 5664
rect 8846 5652 8852 5664
rect 8904 5692 8910 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8904 5664 9229 5692
rect 8904 5652 8910 5664
rect 9217 5661 9229 5664
rect 9263 5692 9275 5695
rect 9490 5692 9496 5704
rect 9263 5664 9496 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9490 5652 9496 5664
rect 9548 5652 9554 5704
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 9858 5692 9864 5704
rect 9732 5664 9864 5692
rect 9732 5652 9738 5664
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 2280 5596 3648 5624
rect 2280 5584 2286 5596
rect 2314 5556 2320 5568
rect 2148 5528 2320 5556
rect 2314 5516 2320 5528
rect 2372 5556 2378 5568
rect 2866 5556 2872 5568
rect 2372 5528 2872 5556
rect 2372 5516 2378 5528
rect 2866 5516 2872 5528
rect 2924 5556 2930 5568
rect 3234 5556 3240 5568
rect 2924 5528 3240 5556
rect 2924 5516 2930 5528
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 10226 5556 10232 5568
rect 9916 5528 10232 5556
rect 9916 5516 9922 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 552 5466 12604 5488
rect 552 5414 3662 5466
rect 3714 5414 3726 5466
rect 3778 5414 3790 5466
rect 3842 5414 3854 5466
rect 3906 5414 3918 5466
rect 3970 5414 10062 5466
rect 10114 5414 10126 5466
rect 10178 5414 10190 5466
rect 10242 5414 10254 5466
rect 10306 5414 10318 5466
rect 10370 5414 12604 5466
rect 552 5392 12604 5414
rect 2774 5312 2780 5364
rect 2832 5312 2838 5364
rect 4154 5312 4160 5364
rect 4212 5312 4218 5364
rect 4706 5312 4712 5364
rect 4764 5312 4770 5364
rect 5166 5312 5172 5364
rect 5224 5312 5230 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 5644 5324 8033 5352
rect 2958 5284 2964 5296
rect 2516 5256 2964 5284
rect 2314 5108 2320 5160
rect 2372 5108 2378 5160
rect 2516 5157 2544 5256
rect 2958 5244 2964 5256
rect 3016 5244 3022 5296
rect 3973 5287 4031 5293
rect 3973 5253 3985 5287
rect 4019 5284 4031 5287
rect 4246 5284 4252 5296
rect 4019 5256 4252 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 4246 5244 4252 5256
rect 4304 5244 4310 5296
rect 4798 5284 4804 5296
rect 4356 5256 4804 5284
rect 3694 5216 3700 5228
rect 3068 5188 3700 5216
rect 3068 5157 3096 5188
rect 3694 5176 3700 5188
rect 3752 5176 3758 5228
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 2593 5151 2651 5157
rect 2593 5117 2605 5151
rect 2639 5117 2651 5151
rect 2593 5111 2651 5117
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 2409 5083 2467 5089
rect 2409 5049 2421 5083
rect 2455 5080 2467 5083
rect 2608 5080 2636 5111
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 4356 5157 4384 5256
rect 4798 5244 4804 5256
rect 4856 5284 4862 5296
rect 5258 5284 5264 5296
rect 4856 5256 5264 5284
rect 4856 5244 4862 5256
rect 5258 5244 5264 5256
rect 5316 5244 5322 5296
rect 5644 5284 5672 5324
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 8021 5315 8079 5321
rect 11333 5355 11391 5361
rect 11333 5321 11345 5355
rect 11379 5352 11391 5355
rect 11606 5352 11612 5364
rect 11379 5324 11612 5352
rect 11379 5321 11391 5324
rect 11333 5315 11391 5321
rect 11606 5312 11612 5324
rect 11664 5352 11670 5364
rect 12158 5352 12164 5364
rect 11664 5324 12164 5352
rect 11664 5312 11670 5324
rect 12158 5312 12164 5324
rect 12216 5312 12222 5364
rect 5552 5256 5672 5284
rect 6917 5287 6975 5293
rect 3605 5151 3663 5157
rect 3605 5148 3617 5151
rect 3476 5120 3617 5148
rect 3476 5108 3482 5120
rect 3605 5117 3617 5120
rect 3651 5117 3663 5151
rect 3605 5111 3663 5117
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4709 5151 4767 5157
rect 4709 5148 4721 5151
rect 4663 5120 4721 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 4709 5117 4721 5120
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 4893 5151 4951 5157
rect 4893 5117 4905 5151
rect 4939 5117 4951 5151
rect 4893 5111 4951 5117
rect 3326 5080 3332 5092
rect 2455 5052 3332 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 3326 5040 3332 5052
rect 3384 5040 3390 5092
rect 4908 5080 4936 5111
rect 4982 5108 4988 5160
rect 5040 5148 5046 5160
rect 5353 5151 5411 5157
rect 5353 5148 5365 5151
rect 5040 5120 5365 5148
rect 5040 5108 5046 5120
rect 5353 5117 5365 5120
rect 5399 5117 5411 5151
rect 5353 5111 5411 5117
rect 5442 5108 5448 5160
rect 5500 5148 5506 5160
rect 5552 5157 5580 5256
rect 6917 5253 6929 5287
rect 6963 5284 6975 5287
rect 7650 5284 7656 5296
rect 6963 5256 7656 5284
rect 6963 5253 6975 5256
rect 6917 5247 6975 5253
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 7745 5287 7803 5293
rect 7745 5253 7757 5287
rect 7791 5253 7803 5287
rect 7745 5247 7803 5253
rect 7929 5287 7987 5293
rect 7929 5253 7941 5287
rect 7975 5284 7987 5287
rect 7975 5256 8708 5284
rect 7975 5253 7987 5256
rect 7929 5247 7987 5253
rect 7760 5216 7788 5247
rect 7116 5188 7788 5216
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5500 5120 5549 5148
rect 5500 5108 5506 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 5718 5148 5724 5160
rect 5675 5120 5724 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 5718 5108 5724 5120
rect 5776 5108 5782 5160
rect 5994 5108 6000 5160
rect 6052 5148 6058 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 6052 5120 6101 5148
rect 6052 5108 6058 5120
rect 6089 5117 6101 5120
rect 6135 5148 6147 5151
rect 6822 5148 6828 5160
rect 6135 5120 6828 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 6822 5108 6828 5120
rect 6880 5108 6886 5160
rect 7116 5157 7144 5188
rect 8110 5176 8116 5228
rect 8168 5176 8174 5228
rect 8680 5225 8708 5256
rect 8846 5244 8852 5296
rect 8904 5284 8910 5296
rect 9033 5287 9091 5293
rect 9033 5284 9045 5287
rect 8904 5256 9045 5284
rect 8904 5244 8910 5256
rect 9033 5253 9045 5256
rect 9079 5253 9091 5287
rect 9033 5247 9091 5253
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 8754 5216 8760 5228
rect 8711 5188 8760 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11330 5216 11336 5228
rect 11195 5188 11336 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11330 5176 11336 5188
rect 11388 5216 11394 5228
rect 12250 5216 12256 5228
rect 11388 5188 12256 5216
rect 11388 5176 11394 5188
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5117 7159 5151
rect 7101 5111 7159 5117
rect 7282 5108 7288 5160
rect 7340 5108 7346 5160
rect 7374 5108 7380 5160
rect 7432 5108 7438 5160
rect 7466 5108 7472 5160
rect 7524 5108 7530 5160
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 8573 5151 8631 5157
rect 8573 5148 8585 5151
rect 7892 5120 8585 5148
rect 7892 5108 7898 5120
rect 8573 5117 8585 5120
rect 8619 5117 8631 5151
rect 9306 5148 9312 5160
rect 8573 5111 8631 5117
rect 8680 5120 9312 5148
rect 4540 5052 4936 5080
rect 2961 5015 3019 5021
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 3142 5012 3148 5024
rect 3007 4984 3148 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 3142 4972 3148 4984
rect 3200 4972 3206 5024
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 4540 5021 4568 5052
rect 5258 5040 5264 5092
rect 5316 5080 5322 5092
rect 5316 5052 5856 5080
rect 5316 5040 5322 5052
rect 4525 5015 4583 5021
rect 4525 5012 4537 5015
rect 4304 4984 4537 5012
rect 4304 4972 4310 4984
rect 4525 4981 4537 4984
rect 4571 4981 4583 5015
rect 4525 4975 4583 4981
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 5828 5012 5856 5052
rect 5902 5040 5908 5092
rect 5960 5040 5966 5092
rect 7392 5080 7420 5108
rect 7561 5083 7619 5089
rect 7561 5080 7573 5083
rect 7392 5052 7573 5080
rect 7561 5049 7573 5052
rect 7607 5049 7619 5083
rect 7561 5043 7619 5049
rect 7745 5083 7803 5089
rect 7745 5049 7757 5083
rect 7791 5049 7803 5083
rect 7745 5043 7803 5049
rect 7098 5012 7104 5024
rect 5828 4984 7104 5012
rect 7098 4972 7104 4984
rect 7156 5012 7162 5024
rect 7760 5012 7788 5043
rect 8294 5040 8300 5092
rect 8352 5080 8358 5092
rect 8680 5080 8708 5120
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 11054 5108 11060 5160
rect 11112 5148 11118 5160
rect 11422 5148 11428 5160
rect 11112 5120 11428 5148
rect 11112 5108 11118 5120
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 8352 5052 8708 5080
rect 8352 5040 8358 5052
rect 9030 5040 9036 5092
rect 9088 5040 9094 5092
rect 11514 5040 11520 5092
rect 11572 5040 11578 5092
rect 11701 5083 11759 5089
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12250 5080 12256 5092
rect 11747 5052 12256 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 12250 5040 12256 5052
rect 12308 5040 12314 5092
rect 7156 4984 7788 5012
rect 7156 4972 7162 4984
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8720 4984 8953 5012
rect 8720 4972 8726 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 9214 4972 9220 5024
rect 9272 4972 9278 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11238 5012 11244 5024
rect 11195 4984 11244 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 552 4922 12604 4944
rect 552 4870 4322 4922
rect 4374 4870 4386 4922
rect 4438 4870 4450 4922
rect 4502 4870 4514 4922
rect 4566 4870 4578 4922
rect 4630 4870 10722 4922
rect 10774 4870 10786 4922
rect 10838 4870 10850 4922
rect 10902 4870 10914 4922
rect 10966 4870 10978 4922
rect 11030 4870 12604 4922
rect 552 4848 12604 4870
rect 3142 4768 3148 4820
rect 3200 4768 3206 4820
rect 3418 4768 3424 4820
rect 3476 4768 3482 4820
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 3752 4780 4261 4808
rect 3752 4768 3758 4780
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 4540 4780 6132 4808
rect 2866 4700 2872 4752
rect 2924 4740 2930 4752
rect 2961 4743 3019 4749
rect 2961 4740 2973 4743
rect 2924 4712 2973 4740
rect 2924 4700 2930 4712
rect 2961 4709 2973 4712
rect 3007 4709 3019 4743
rect 2961 4703 3019 4709
rect 2777 4675 2835 4681
rect 2777 4641 2789 4675
rect 2823 4641 2835 4675
rect 3160 4672 3188 4768
rect 3237 4675 3295 4681
rect 3237 4672 3249 4675
rect 3160 4644 3249 4672
rect 2777 4635 2835 4641
rect 3237 4641 3249 4644
rect 3283 4641 3295 4675
rect 3237 4635 3295 4641
rect 2792 4604 2820 4635
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 4540 4681 4568 4780
rect 6104 4752 6132 4780
rect 6454 4768 6460 4820
rect 6512 4808 6518 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 6512 4780 6561 4808
rect 6512 4768 6518 4780
rect 6549 4777 6561 4780
rect 6595 4777 6607 4811
rect 6549 4771 6607 4777
rect 7653 4811 7711 4817
rect 7653 4777 7665 4811
rect 7699 4808 7711 4811
rect 7834 4808 7840 4820
rect 7699 4780 7840 4808
rect 7699 4777 7711 4780
rect 7653 4771 7711 4777
rect 7834 4768 7840 4780
rect 7892 4768 7898 4820
rect 8846 4808 8852 4820
rect 7944 4780 8852 4808
rect 5718 4740 5724 4752
rect 4908 4712 5724 4740
rect 4908 4681 4936 4712
rect 5718 4700 5724 4712
rect 5776 4700 5782 4752
rect 6086 4700 6092 4752
rect 6144 4740 6150 4752
rect 7944 4740 7972 4780
rect 8846 4768 8852 4780
rect 8904 4768 8910 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9398 4808 9404 4820
rect 9079 4780 9404 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 11133 4811 11191 4817
rect 11133 4777 11145 4811
rect 11179 4808 11191 4811
rect 11606 4808 11612 4820
rect 11179 4780 11612 4808
rect 11179 4777 11191 4780
rect 11133 4771 11191 4777
rect 11606 4768 11612 4780
rect 11664 4768 11670 4820
rect 8570 4740 8576 4752
rect 6144 4712 7972 4740
rect 8036 4712 8576 4740
rect 6144 4700 6150 4712
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 3384 4644 3433 4672
rect 3384 4632 3390 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 3421 4635 3479 4641
rect 4525 4675 4583 4681
rect 4525 4641 4537 4675
rect 4571 4641 4583 4675
rect 4525 4635 4583 4641
rect 4892 4675 4950 4681
rect 4892 4641 4904 4675
rect 4938 4641 4950 4675
rect 4892 4635 4950 4641
rect 4982 4632 4988 4684
rect 5040 4632 5046 4684
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 5442 4672 5448 4684
rect 5307 4644 5448 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6181 4635 6239 4641
rect 2958 4604 2964 4616
rect 2792 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4604 4675 4607
rect 5169 4607 5227 4613
rect 5169 4604 5181 4607
rect 4663 4576 5181 4604
rect 4663 4573 4675 4576
rect 4617 4567 4675 4573
rect 5169 4573 5181 4576
rect 5215 4573 5227 4607
rect 5169 4567 5227 4573
rect 4264 4536 4292 4567
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 5868 4576 6101 4604
rect 5868 4564 5874 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 5258 4536 5264 4548
rect 4264 4508 5264 4536
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 5629 4539 5687 4545
rect 5629 4505 5641 4539
rect 5675 4536 5687 4539
rect 6196 4536 6224 4635
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 6822 4632 6828 4684
rect 6880 4632 6886 4684
rect 8036 4681 8064 4712
rect 8570 4700 8576 4712
rect 8628 4740 8634 4752
rect 9214 4740 9220 4752
rect 8628 4712 9220 4740
rect 8628 4700 8634 4712
rect 9214 4700 9220 4712
rect 9272 4700 9278 4752
rect 9306 4700 9312 4752
rect 9364 4740 9370 4752
rect 9585 4743 9643 4749
rect 9585 4740 9597 4743
rect 9364 4712 9597 4740
rect 9364 4700 9370 4712
rect 9585 4709 9597 4712
rect 9631 4740 9643 4743
rect 9674 4740 9680 4752
rect 9631 4712 9680 4740
rect 9631 4709 9643 4712
rect 9585 4703 9643 4709
rect 9674 4700 9680 4712
rect 9732 4740 9738 4752
rect 11333 4743 11391 4749
rect 11333 4740 11345 4743
rect 9732 4712 11345 4740
rect 9732 4700 9738 4712
rect 11333 4709 11345 4712
rect 11379 4740 11391 4743
rect 11514 4740 11520 4752
rect 11379 4712 11520 4740
rect 11379 4709 11391 4712
rect 11333 4703 11391 4709
rect 11514 4700 11520 4712
rect 11572 4700 11578 4752
rect 7285 4675 7343 4681
rect 7285 4641 7297 4675
rect 7331 4641 7343 4675
rect 7285 4635 7343 4641
rect 8021 4675 8079 4681
rect 8021 4641 8033 4675
rect 8067 4641 8079 4675
rect 8021 4635 8079 4641
rect 5675 4508 6224 4536
rect 7300 4536 7328 4635
rect 8662 4632 8668 4684
rect 8720 4632 8726 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 9490 4672 9496 4684
rect 9447 4644 9496 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 10597 4675 10655 4681
rect 10597 4641 10609 4675
rect 10643 4641 10655 4675
rect 10597 4635 10655 4641
rect 10781 4675 10839 4681
rect 10781 4641 10793 4675
rect 10827 4672 10839 4675
rect 11238 4672 11244 4684
rect 10827 4644 11244 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 7926 4604 7932 4616
rect 7423 4576 7932 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8573 4607 8631 4613
rect 8573 4604 8585 4607
rect 8404 4576 8585 4604
rect 8404 4545 8432 4576
rect 8573 4573 8585 4576
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 8389 4539 8447 4545
rect 7300 4508 7603 4536
rect 5675 4505 5687 4508
rect 5629 4499 5687 4505
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 7009 4471 7067 4477
rect 7009 4437 7021 4471
rect 7055 4468 7067 4471
rect 7466 4468 7472 4480
rect 7055 4440 7472 4468
rect 7055 4437 7067 4440
rect 7009 4431 7067 4437
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 7575 4468 7603 4508
rect 8389 4505 8401 4539
rect 8435 4505 8447 4539
rect 10612 4536 10640 4635
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 11606 4632 11612 4684
rect 11664 4632 11670 4684
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12342 4672 12348 4684
rect 12207 4644 12348 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 11146 4604 11152 4616
rect 10735 4576 11152 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11422 4564 11428 4616
rect 11480 4604 11486 4616
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 11480 4576 11805 4604
rect 11480 4564 11486 4576
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 11808 4536 11836 4567
rect 11977 4539 12035 4545
rect 11977 4536 11989 4539
rect 10612 4508 11468 4536
rect 11808 4508 11989 4536
rect 8389 4499 8447 4505
rect 8754 4468 8760 4480
rect 7575 4440 8760 4468
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9769 4471 9827 4477
rect 9769 4468 9781 4471
rect 9732 4440 9781 4468
rect 9732 4428 9738 4440
rect 9769 4437 9781 4440
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 10410 4428 10416 4480
rect 10468 4468 10474 4480
rect 10965 4471 11023 4477
rect 10965 4468 10977 4471
rect 10468 4440 10977 4468
rect 10468 4428 10474 4440
rect 10965 4437 10977 4440
rect 11011 4437 11023 4471
rect 10965 4431 11023 4437
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11440 4477 11468 4508
rect 11977 4505 11989 4508
rect 12023 4505 12035 4539
rect 11977 4499 12035 4505
rect 11158 4471 11216 4477
rect 11158 4468 11170 4471
rect 11112 4440 11170 4468
rect 11112 4428 11118 4440
rect 11158 4437 11170 4440
rect 11204 4437 11216 4471
rect 11158 4431 11216 4437
rect 11425 4471 11483 4477
rect 11425 4437 11437 4471
rect 11471 4468 11483 4471
rect 11698 4468 11704 4480
rect 11471 4440 11704 4468
rect 11471 4437 11483 4440
rect 11425 4431 11483 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 552 4378 12604 4400
rect 552 4326 3662 4378
rect 3714 4326 3726 4378
rect 3778 4326 3790 4378
rect 3842 4326 3854 4378
rect 3906 4326 3918 4378
rect 3970 4326 10062 4378
rect 10114 4326 10126 4378
rect 10178 4326 10190 4378
rect 10242 4326 10254 4378
rect 10306 4326 10318 4378
rect 10370 4326 12604 4378
rect 552 4304 12604 4326
rect 2777 4267 2835 4273
rect 2777 4233 2789 4267
rect 2823 4264 2835 4267
rect 2866 4264 2872 4276
rect 2823 4236 2872 4264
rect 2823 4233 2835 4236
rect 2777 4227 2835 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4341 4267 4399 4273
rect 4341 4264 4353 4267
rect 4304 4236 4353 4264
rect 4304 4224 4310 4236
rect 4341 4233 4353 4236
rect 4387 4233 4399 4267
rect 4341 4227 4399 4233
rect 4982 4224 4988 4276
rect 5040 4264 5046 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 5040 4236 5273 4264
rect 5040 4224 5046 4236
rect 5261 4233 5273 4236
rect 5307 4233 5319 4267
rect 5261 4227 5319 4233
rect 5810 4224 5816 4276
rect 5868 4224 5874 4276
rect 7285 4267 7343 4273
rect 7285 4233 7297 4267
rect 7331 4264 7343 4267
rect 7374 4264 7380 4276
rect 7331 4236 7380 4264
rect 7331 4233 7343 4236
rect 7285 4227 7343 4233
rect 7374 4224 7380 4236
rect 7432 4224 7438 4276
rect 8110 4224 8116 4276
rect 8168 4224 8174 4276
rect 8386 4224 8392 4276
rect 8444 4224 8450 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 8757 4267 8815 4273
rect 8757 4264 8769 4267
rect 8536 4236 8769 4264
rect 8536 4224 8542 4236
rect 8757 4233 8769 4236
rect 8803 4264 8815 4267
rect 9030 4264 9036 4276
rect 8803 4236 9036 4264
rect 8803 4233 8815 4236
rect 8757 4227 8815 4233
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 12253 4267 12311 4273
rect 9416 4236 10272 4264
rect 6089 4199 6147 4205
rect 6089 4196 6101 4199
rect 2746 4168 4292 4196
rect 2746 4140 2774 4168
rect 2682 4088 2688 4140
rect 2740 4100 2774 4140
rect 2740 4088 2746 4100
rect 4154 4088 4160 4140
rect 4212 4088 4218 4140
rect 1394 4020 1400 4072
rect 1452 4020 1458 4072
rect 4065 4063 4123 4069
rect 4065 4029 4077 4063
rect 4111 4029 4123 4063
rect 4264 4060 4292 4168
rect 5276 4168 6101 4196
rect 5276 4140 5304 4168
rect 6089 4165 6101 4168
rect 6135 4165 6147 4199
rect 6089 4159 6147 4165
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 8404 4196 8432 4224
rect 9416 4196 9444 4236
rect 6604 4168 8248 4196
rect 8404 4168 9444 4196
rect 6604 4156 6610 4168
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4632 4100 4905 4128
rect 4632 4069 4660 4100
rect 4893 4097 4905 4100
rect 4939 4128 4951 4131
rect 5166 4128 5172 4140
rect 4939 4100 5172 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4128 5687 4131
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5675 4100 6009 4128
rect 5675 4097 5687 4100
rect 5629 4091 5687 4097
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 7006 4088 7012 4140
rect 7064 4088 7070 4140
rect 8220 4072 8248 4168
rect 9766 4156 9772 4208
rect 9824 4156 9830 4208
rect 10244 4205 10272 4236
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12342 4264 12348 4276
rect 12299 4236 12348 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12342 4224 12348 4236
rect 12400 4224 12406 4276
rect 10229 4199 10287 4205
rect 10229 4165 10241 4199
rect 10275 4165 10287 4199
rect 10229 4159 10287 4165
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4128 8447 4131
rect 8754 4128 8760 4140
rect 8435 4100 8760 4128
rect 8435 4097 8447 4100
rect 8389 4091 8447 4097
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 9784 4128 9812 4156
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9508 4100 9873 4128
rect 4617 4063 4675 4069
rect 4617 4060 4629 4063
rect 4264 4032 4629 4060
rect 4065 4023 4123 4029
rect 4617 4029 4629 4032
rect 4663 4029 4675 4063
rect 4617 4023 4675 4029
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 4982 4060 4988 4072
rect 4847 4032 4988 4060
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 1670 4001 1676 4004
rect 1664 3955 1676 4001
rect 1670 3952 1676 3955
rect 1728 3952 1734 4004
rect 4080 3936 4108 4023
rect 4982 4020 4988 4032
rect 5040 4020 5046 4072
rect 5077 4063 5135 4069
rect 5077 4029 5089 4063
rect 5123 4060 5135 4063
rect 5442 4060 5448 4072
rect 5123 4032 5448 4060
rect 5123 4029 5135 4032
rect 5077 4023 5135 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4060 5595 4063
rect 6086 4060 6092 4072
rect 5583 4032 6092 4060
rect 5583 4029 5595 4032
rect 5537 4023 5595 4029
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 4430 3952 4436 4004
rect 4488 3992 4494 4004
rect 4709 3995 4767 4001
rect 4709 3992 4721 3995
rect 4488 3964 4721 3992
rect 4488 3952 4494 3964
rect 4709 3961 4721 3964
rect 4755 3992 4767 3995
rect 6457 3995 6515 4001
rect 6457 3992 6469 3995
rect 4755 3964 6469 3992
rect 4755 3961 4767 3964
rect 4709 3955 4767 3961
rect 6457 3961 6469 3964
rect 6503 3961 6515 3995
rect 6932 3992 6960 4023
rect 7466 4020 7472 4072
rect 7524 4060 7530 4072
rect 7561 4063 7619 4069
rect 7561 4060 7573 4063
rect 7524 4032 7573 4060
rect 7524 4020 7530 4032
rect 7561 4029 7573 4032
rect 7607 4029 7619 4063
rect 7561 4023 7619 4029
rect 7834 4020 7840 4072
rect 7892 4020 7898 4072
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8202 4020 8208 4072
rect 8260 4020 8266 4072
rect 8573 4063 8631 4069
rect 8573 4029 8585 4063
rect 8619 4060 8631 4063
rect 8938 4060 8944 4072
rect 8619 4032 8944 4060
rect 8619 4029 8631 4032
rect 8573 4023 8631 4029
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9508 4069 9536 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 9493 4063 9551 4069
rect 9493 4029 9505 4063
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 9766 4020 9772 4072
rect 9824 4020 9830 4072
rect 10152 4060 10180 4091
rect 10502 4088 10508 4140
rect 10560 4088 10566 4140
rect 10686 4088 10692 4140
rect 10744 4128 10750 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10744 4100 10885 4128
rect 10744 4088 10750 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 11146 4069 11152 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10152 4032 10609 4060
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 11140 4060 11152 4069
rect 11107 4032 11152 4060
rect 10597 4023 10655 4029
rect 11140 4023 11152 4032
rect 11146 4020 11152 4023
rect 11204 4020 11210 4072
rect 7745 3995 7803 4001
rect 7745 3992 7757 3995
rect 6932 3964 7757 3992
rect 6457 3955 6515 3961
rect 7745 3961 7757 3964
rect 7791 3992 7803 3995
rect 9033 3995 9091 4001
rect 9033 3992 9045 3995
rect 7791 3964 9045 3992
rect 7791 3961 7803 3964
rect 7745 3955 7803 3961
rect 9033 3961 9045 3964
rect 9079 3961 9091 3995
rect 9033 3955 9091 3961
rect 9401 3995 9459 4001
rect 9401 3961 9413 3995
rect 9447 3992 9459 3995
rect 9674 3992 9680 4004
rect 9447 3964 9680 3992
rect 9447 3961 9459 3964
rect 9401 3955 9459 3961
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 7377 3927 7435 3933
rect 7377 3924 7389 3927
rect 4120 3896 7389 3924
rect 4120 3884 4126 3896
rect 7377 3893 7389 3896
rect 7423 3893 7435 3927
rect 7377 3887 7435 3893
rect 552 3834 12604 3856
rect 552 3782 4322 3834
rect 4374 3782 4386 3834
rect 4438 3782 4450 3834
rect 4502 3782 4514 3834
rect 4566 3782 4578 3834
rect 4630 3782 10722 3834
rect 10774 3782 10786 3834
rect 10838 3782 10850 3834
rect 10902 3782 10914 3834
rect 10966 3782 10978 3834
rect 11030 3782 12604 3834
rect 552 3760 12604 3782
rect 1670 3680 1676 3732
rect 1728 3680 1734 3732
rect 2406 3720 2412 3732
rect 1780 3692 2412 3720
rect 1213 3655 1271 3661
rect 1213 3621 1225 3655
rect 1259 3621 1271 3655
rect 1213 3615 1271 3621
rect 1429 3655 1487 3661
rect 1429 3621 1441 3655
rect 1475 3652 1487 3655
rect 1780 3652 1808 3692
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2682 3680 2688 3732
rect 2740 3680 2746 3732
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 5169 3723 5227 3729
rect 5169 3720 5181 3723
rect 4212 3692 5181 3720
rect 4212 3680 4218 3692
rect 5169 3689 5181 3692
rect 5215 3689 5227 3723
rect 5169 3683 5227 3689
rect 5258 3680 5264 3732
rect 5316 3680 5322 3732
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 6822 3720 6828 3732
rect 5500 3692 6828 3720
rect 5500 3680 5506 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7285 3723 7343 3729
rect 7285 3720 7297 3723
rect 7064 3692 7297 3720
rect 7064 3680 7070 3692
rect 7285 3689 7297 3692
rect 7331 3689 7343 3723
rect 7285 3683 7343 3689
rect 8570 3680 8576 3732
rect 8628 3680 8634 3732
rect 9214 3680 9220 3732
rect 9272 3720 9278 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 9272 3692 9597 3720
rect 9272 3680 9278 3692
rect 9585 3689 9597 3692
rect 9631 3689 9643 3723
rect 9585 3683 9643 3689
rect 1475 3624 1808 3652
rect 1857 3655 1915 3661
rect 1475 3621 1487 3624
rect 1429 3615 1487 3621
rect 1857 3621 1869 3655
rect 1903 3652 1915 3655
rect 2317 3655 2375 3661
rect 2317 3652 2329 3655
rect 1903 3624 2329 3652
rect 1903 3621 1915 3624
rect 1857 3615 1915 3621
rect 2317 3621 2329 3624
rect 2363 3621 2375 3655
rect 2866 3652 2872 3664
rect 2317 3615 2375 3621
rect 2516 3624 2872 3652
rect 1228 3584 1256 3615
rect 2516 3593 2544 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 3513 3655 3571 3661
rect 3513 3621 3525 3655
rect 3559 3652 3571 3655
rect 3559 3624 4844 3652
rect 3559 3621 3571 3624
rect 3513 3615 3571 3621
rect 2501 3587 2559 3593
rect 2501 3584 2513 3587
rect 1228 3556 2513 3584
rect 2501 3553 2513 3556
rect 2547 3553 2559 3587
rect 2501 3547 2559 3553
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 1854 3476 1860 3528
rect 1912 3516 1918 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 1912 3488 2237 3516
rect 1912 3476 1918 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2225 3479 2283 3485
rect 2406 3476 2412 3528
rect 2464 3516 2470 3528
rect 2792 3516 2820 3547
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 4448 3593 4476 3624
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 3292 3556 3341 3584
rect 3292 3544 3298 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3329 3547 3387 3553
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 4249 3587 4307 3593
rect 4249 3584 4261 3587
rect 3835 3556 4261 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 4249 3553 4261 3556
rect 4295 3553 4307 3587
rect 4249 3547 4307 3553
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3553 4491 3587
rect 4433 3547 4491 3553
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 2464 3488 2820 3516
rect 3145 3519 3203 3525
rect 2464 3476 2470 3488
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 1872 3448 1900 3476
rect 2700 3460 2728 3488
rect 3145 3485 3157 3519
rect 3191 3516 3203 3519
rect 3418 3516 3424 3528
rect 3191 3488 3424 3516
rect 3191 3485 3203 3488
rect 3145 3479 3203 3485
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3510 3476 3516 3528
rect 3568 3516 3574 3528
rect 3697 3519 3755 3525
rect 3697 3516 3709 3519
rect 3568 3488 3709 3516
rect 3568 3476 3574 3488
rect 3697 3485 3709 3488
rect 3743 3485 3755 3519
rect 3697 3479 3755 3485
rect 4062 3476 4068 3528
rect 4120 3516 4126 3528
rect 4632 3516 4660 3547
rect 4706 3544 4712 3596
rect 4764 3544 4770 3596
rect 4816 3593 4844 3624
rect 4982 3612 4988 3664
rect 5040 3652 5046 3664
rect 5040 3624 5396 3652
rect 5040 3612 5046 3624
rect 5368 3596 5396 3624
rect 6730 3612 6736 3664
rect 6788 3652 6794 3664
rect 7193 3655 7251 3661
rect 6788 3624 7052 3652
rect 6788 3612 6794 3624
rect 4801 3587 4859 3593
rect 4801 3553 4813 3587
rect 4847 3553 4859 3587
rect 4801 3547 4859 3553
rect 4894 3587 4952 3593
rect 4894 3553 4906 3587
rect 4940 3553 4952 3587
rect 4894 3547 4952 3553
rect 4120 3488 4660 3516
rect 4724 3516 4752 3544
rect 4908 3516 4936 3547
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 5224 3556 5273 3584
rect 5224 3544 5230 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 5350 3544 5356 3596
rect 5408 3584 5414 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 5408 3556 5457 3584
rect 5408 3544 5414 3556
rect 5445 3553 5457 3556
rect 5491 3553 5503 3587
rect 5445 3547 5503 3553
rect 6822 3544 6828 3596
rect 6880 3544 6886 3596
rect 7024 3593 7052 3624
rect 7193 3621 7205 3655
rect 7239 3652 7251 3655
rect 7834 3652 7840 3664
rect 7239 3624 7840 3652
rect 7239 3621 7251 3624
rect 7193 3615 7251 3621
rect 7009 3587 7067 3593
rect 7009 3553 7021 3587
rect 7055 3584 7067 3587
rect 7374 3584 7380 3596
rect 7055 3556 7380 3584
rect 7055 3553 7067 3556
rect 7009 3547 7067 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7576 3593 7604 3624
rect 7834 3612 7840 3624
rect 7892 3612 7898 3664
rect 7560 3587 7618 3593
rect 7560 3584 7572 3587
rect 7539 3556 7572 3584
rect 7560 3553 7572 3556
rect 7606 3553 7618 3587
rect 7560 3547 7618 3553
rect 7653 3587 7711 3593
rect 7653 3553 7665 3587
rect 7699 3553 7711 3587
rect 7653 3547 7711 3553
rect 4724 3488 4936 3516
rect 4120 3476 4126 3488
rect 7466 3476 7472 3528
rect 7524 3516 7530 3528
rect 7668 3516 7696 3547
rect 8478 3544 8484 3596
rect 8536 3544 8542 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3553 8723 3587
rect 8665 3547 8723 3553
rect 7524 3488 7696 3516
rect 8680 3516 8708 3547
rect 8754 3544 8760 3596
rect 8812 3544 8818 3596
rect 8938 3544 8944 3596
rect 8996 3544 9002 3596
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9306 3584 9312 3596
rect 9088 3556 9312 3584
rect 9088 3544 9094 3556
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9401 3587 9459 3593
rect 9401 3553 9413 3587
rect 9447 3584 9459 3587
rect 9490 3584 9496 3596
rect 9447 3556 9496 3584
rect 9447 3553 9459 3556
rect 9401 3547 9459 3553
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 9600 3584 9628 3683
rect 9766 3680 9772 3732
rect 9824 3720 9830 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9824 3692 10057 3720
rect 9824 3680 9830 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 11333 3655 11391 3661
rect 11333 3621 11345 3655
rect 11379 3652 11391 3655
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11379 3624 11621 3652
rect 11379 3621 11391 3624
rect 11333 3615 11391 3621
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 11698 3612 11704 3664
rect 11756 3652 11762 3664
rect 11977 3655 12035 3661
rect 11977 3652 11989 3655
rect 11756 3624 11989 3652
rect 11756 3612 11762 3624
rect 11977 3621 11989 3624
rect 12023 3621 12035 3655
rect 11977 3615 12035 3621
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9600 3556 9689 3584
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 9824 3556 9869 3584
rect 9824 3544 9830 3556
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11514 3584 11520 3596
rect 11296 3556 11520 3584
rect 11296 3544 11302 3556
rect 11514 3544 11520 3556
rect 11572 3584 11578 3596
rect 11793 3587 11851 3593
rect 11793 3584 11805 3587
rect 11572 3556 11805 3584
rect 11572 3544 11578 3556
rect 11793 3553 11805 3556
rect 11839 3553 11851 3587
rect 11793 3547 11851 3553
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8680 3488 8861 3516
rect 7524 3476 7530 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 8849 3479 8907 3485
rect 1627 3420 1900 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2682 3408 2688 3460
rect 2740 3408 2746 3460
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 10428 3448 10456 3544
rect 10965 3451 11023 3457
rect 10965 3448 10977 3451
rect 9732 3420 10977 3448
rect 9732 3408 9738 3420
rect 10965 3417 10977 3420
rect 11011 3417 11023 3451
rect 10965 3411 11023 3417
rect 1397 3383 1455 3389
rect 1397 3349 1409 3383
rect 1443 3380 1455 3383
rect 1486 3380 1492 3392
rect 1443 3352 1492 3380
rect 1443 3349 1455 3352
rect 1397 3343 1455 3349
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 1857 3383 1915 3389
rect 1857 3349 1869 3383
rect 1903 3380 1915 3383
rect 2038 3380 2044 3392
rect 1903 3352 2044 3380
rect 1903 3349 1915 3352
rect 1857 3343 1915 3349
rect 2038 3340 2044 3352
rect 2096 3340 2102 3392
rect 4065 3383 4123 3389
rect 4065 3349 4077 3383
rect 4111 3380 4123 3383
rect 4890 3380 4896 3392
rect 4111 3352 4896 3380
rect 4111 3349 4123 3352
rect 4065 3343 4123 3349
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 9582 3340 9588 3392
rect 9640 3380 9646 3392
rect 9766 3380 9772 3392
rect 9640 3352 9772 3380
rect 9640 3340 9646 3352
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 11330 3340 11336 3392
rect 11388 3340 11394 3392
rect 11514 3340 11520 3392
rect 11572 3340 11578 3392
rect 552 3290 12604 3312
rect 552 3238 3662 3290
rect 3714 3238 3726 3290
rect 3778 3238 3790 3290
rect 3842 3238 3854 3290
rect 3906 3238 3918 3290
rect 3970 3238 10062 3290
rect 10114 3238 10126 3290
rect 10178 3238 10190 3290
rect 10242 3238 10254 3290
rect 10306 3238 10318 3290
rect 10370 3238 12604 3290
rect 552 3216 12604 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 2498 3176 2504 3188
rect 1544 3148 2504 3176
rect 1544 3136 1550 3148
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 4525 3179 4583 3185
rect 4525 3145 4537 3179
rect 4571 3176 4583 3179
rect 4706 3176 4712 3188
rect 4571 3148 4712 3176
rect 4571 3145 4583 3148
rect 4525 3139 4583 3145
rect 4706 3136 4712 3148
rect 4764 3136 4770 3188
rect 12250 3136 12256 3188
rect 12308 3136 12314 3188
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2372 3012 2421 3040
rect 2372 3000 2378 3012
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 2869 3043 2927 3049
rect 2869 3009 2881 3043
rect 2915 3040 2927 3043
rect 3142 3040 3148 3052
rect 2915 3012 3148 3040
rect 2915 3009 2927 3012
rect 2869 3003 2927 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10652 3012 10885 3040
rect 10652 3000 10658 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 1872 2904 1900 2935
rect 2498 2932 2504 2984
rect 2556 2932 2562 2984
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 4154 2972 4160 2984
rect 3292 2944 4160 2972
rect 3292 2932 3298 2944
rect 4154 2932 4160 2944
rect 4212 2932 4218 2984
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 6549 2975 6607 2981
rect 6549 2972 6561 2975
rect 6420 2944 6561 2972
rect 6420 2932 6426 2944
rect 6549 2941 6561 2944
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6733 2975 6791 2981
rect 6733 2972 6745 2975
rect 6696 2944 6745 2972
rect 6696 2932 6702 2944
rect 6733 2941 6745 2944
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 11140 2975 11198 2981
rect 11140 2941 11152 2975
rect 11186 2972 11198 2975
rect 11514 2972 11520 2984
rect 11186 2944 11520 2972
rect 11186 2941 11198 2944
rect 11140 2935 11198 2941
rect 11514 2932 11520 2944
rect 11572 2932 11578 2984
rect 2866 2904 2872 2916
rect 1872 2876 2872 2904
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 3418 2864 3424 2916
rect 3476 2904 3482 2916
rect 4246 2904 4252 2916
rect 3476 2876 4252 2904
rect 3476 2864 3482 2876
rect 4246 2864 4252 2876
rect 4304 2904 4310 2916
rect 4341 2907 4399 2913
rect 4341 2904 4353 2907
rect 4304 2876 4353 2904
rect 4304 2864 4310 2876
rect 4341 2873 4353 2876
rect 4387 2873 4399 2907
rect 4341 2867 4399 2873
rect 6641 2839 6699 2845
rect 6641 2805 6653 2839
rect 6687 2836 6699 2839
rect 6730 2836 6736 2848
rect 6687 2808 6736 2836
rect 6687 2805 6699 2808
rect 6641 2799 6699 2805
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 552 2746 12604 2768
rect 552 2694 4322 2746
rect 4374 2694 4386 2746
rect 4438 2694 4450 2746
rect 4502 2694 4514 2746
rect 4566 2694 4578 2746
rect 4630 2694 10722 2746
rect 10774 2694 10786 2746
rect 10838 2694 10850 2746
rect 10902 2694 10914 2746
rect 10966 2694 10978 2746
rect 11030 2694 12604 2746
rect 552 2672 12604 2694
rect 3510 2592 3516 2644
rect 3568 2592 3574 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7282 2632 7288 2644
rect 6871 2604 7288 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7453 2635 7511 2641
rect 7453 2601 7465 2635
rect 7499 2632 7511 2635
rect 9490 2632 9496 2644
rect 7499 2604 9496 2632
rect 7499 2601 7511 2604
rect 7453 2595 7511 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10321 2635 10379 2641
rect 10321 2601 10333 2635
rect 10367 2632 10379 2635
rect 10502 2632 10508 2644
rect 10367 2604 10508 2632
rect 10367 2601 10379 2604
rect 10321 2595 10379 2601
rect 10502 2592 10508 2604
rect 10560 2592 10566 2644
rect 4246 2524 4252 2576
rect 4304 2564 4310 2576
rect 5997 2567 6055 2573
rect 5997 2564 6009 2567
rect 4304 2536 6009 2564
rect 4304 2524 4310 2536
rect 5997 2533 6009 2536
rect 6043 2564 6055 2567
rect 7650 2564 7656 2576
rect 6043 2536 7656 2564
rect 6043 2533 6055 2536
rect 5997 2527 6055 2533
rect 7650 2524 7656 2536
rect 7708 2564 7714 2576
rect 8754 2564 8760 2576
rect 7708 2536 8760 2564
rect 7708 2524 7714 2536
rect 8754 2524 8760 2536
rect 8812 2524 8818 2576
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 9766 2564 9772 2576
rect 9263 2536 9772 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 10686 2564 10692 2576
rect 9968 2536 10692 2564
rect 2498 2456 2504 2508
rect 2556 2456 2562 2508
rect 3142 2456 3148 2508
rect 3200 2456 3206 2508
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5810 2496 5816 2508
rect 5500 2468 5816 2496
rect 5500 2456 5506 2468
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6454 2456 6460 2508
rect 6512 2456 6518 2508
rect 7009 2499 7067 2505
rect 7009 2465 7021 2499
rect 7055 2465 7067 2499
rect 7009 2459 7067 2465
rect 7193 2499 7251 2505
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7282 2496 7288 2508
rect 7239 2468 7288 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2280 2400 2421 2428
rect 2280 2388 2286 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 2409 2391 2467 2397
rect 2884 2400 3065 2428
rect 2884 2369 2912 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 2869 2363 2927 2369
rect 2869 2329 2881 2363
rect 2915 2329 2927 2363
rect 7024 2360 7052 2459
rect 7282 2456 7288 2468
rect 7340 2456 7346 2508
rect 8021 2499 8079 2505
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8202 2496 8208 2508
rect 8067 2468 8208 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8570 2456 8576 2508
rect 8628 2496 8634 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8628 2468 8677 2496
rect 8628 2456 8634 2468
rect 8665 2465 8677 2468
rect 8711 2465 8723 2499
rect 8665 2459 8723 2465
rect 8849 2499 8907 2505
rect 8849 2465 8861 2499
rect 8895 2465 8907 2499
rect 8849 2459 8907 2465
rect 7742 2388 7748 2440
rect 7800 2388 7806 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8864 2428 8892 2459
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 9125 2499 9183 2505
rect 9125 2496 9137 2499
rect 8996 2468 9137 2496
rect 8996 2456 9002 2468
rect 9125 2465 9137 2468
rect 9171 2465 9183 2499
rect 9125 2459 9183 2465
rect 9309 2499 9367 2505
rect 9309 2465 9321 2499
rect 9355 2465 9367 2499
rect 9309 2459 9367 2465
rect 9493 2499 9551 2505
rect 9493 2465 9505 2499
rect 9539 2496 9551 2499
rect 9674 2496 9680 2508
rect 9539 2468 9680 2496
rect 9539 2465 9551 2468
rect 9493 2459 9551 2465
rect 9324 2428 9352 2459
rect 9674 2456 9680 2468
rect 9732 2496 9738 2508
rect 9968 2505 9996 2536
rect 10686 2524 10692 2536
rect 10744 2524 10750 2576
rect 9953 2499 10011 2505
rect 9732 2468 9812 2496
rect 9732 2456 9738 2468
rect 8168 2400 8892 2428
rect 9140 2400 9352 2428
rect 8168 2388 8174 2400
rect 9140 2372 9168 2400
rect 7285 2363 7343 2369
rect 7285 2360 7297 2363
rect 2869 2323 2927 2329
rect 6104 2332 6500 2360
rect 2682 2252 2688 2304
rect 2740 2292 2746 2304
rect 6104 2292 6132 2332
rect 2740 2264 6132 2292
rect 6181 2295 6239 2301
rect 2740 2252 2746 2264
rect 6181 2261 6193 2295
rect 6227 2292 6239 2295
rect 6270 2292 6276 2304
rect 6227 2264 6276 2292
rect 6227 2261 6239 2264
rect 6181 2255 6239 2261
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 6472 2292 6500 2332
rect 7024 2332 7297 2360
rect 7024 2292 7052 2332
rect 7285 2329 7297 2332
rect 7331 2329 7343 2363
rect 7285 2323 7343 2329
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 9122 2360 9128 2372
rect 8536 2332 9128 2360
rect 8536 2320 8542 2332
rect 9122 2320 9128 2332
rect 9180 2320 9186 2372
rect 9784 2360 9812 2468
rect 9953 2465 9965 2499
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 10410 2456 10416 2508
rect 10468 2496 10474 2508
rect 10597 2499 10655 2505
rect 10597 2496 10609 2499
rect 10468 2468 10609 2496
rect 10468 2456 10474 2468
rect 10597 2465 10609 2468
rect 10643 2465 10655 2499
rect 10597 2459 10655 2465
rect 10042 2388 10048 2440
rect 10100 2428 10106 2440
rect 10502 2428 10508 2440
rect 10100 2400 10508 2428
rect 10100 2388 10106 2400
rect 10502 2388 10508 2400
rect 10560 2388 10566 2440
rect 10413 2363 10471 2369
rect 10413 2360 10425 2363
rect 9784 2332 10425 2360
rect 10413 2329 10425 2332
rect 10459 2329 10471 2363
rect 10413 2323 10471 2329
rect 6472 2264 7052 2292
rect 7190 2252 7196 2304
rect 7248 2252 7254 2304
rect 7466 2252 7472 2304
rect 7524 2252 7530 2304
rect 8662 2252 8668 2304
rect 8720 2252 8726 2304
rect 9140 2292 9168 2320
rect 9585 2295 9643 2301
rect 9585 2292 9597 2295
rect 9140 2264 9597 2292
rect 9585 2261 9597 2264
rect 9631 2292 9643 2295
rect 10778 2292 10784 2304
rect 9631 2264 10784 2292
rect 9631 2261 9643 2264
rect 9585 2255 9643 2261
rect 10778 2252 10784 2264
rect 10836 2252 10842 2304
rect 552 2202 12604 2224
rect 552 2150 3662 2202
rect 3714 2150 3726 2202
rect 3778 2150 3790 2202
rect 3842 2150 3854 2202
rect 3906 2150 3918 2202
rect 3970 2150 10062 2202
rect 10114 2150 10126 2202
rect 10178 2150 10190 2202
rect 10242 2150 10254 2202
rect 10306 2150 10318 2202
rect 10370 2150 12604 2202
rect 552 2128 12604 2150
rect 2498 2048 2504 2100
rect 2556 2088 2562 2100
rect 3237 2091 3295 2097
rect 3237 2088 3249 2091
rect 2556 2060 3249 2088
rect 2556 2048 2562 2060
rect 3237 2057 3249 2060
rect 3283 2057 3295 2091
rect 3237 2051 3295 2057
rect 3326 2048 3332 2100
rect 3384 2088 3390 2100
rect 3973 2091 4031 2097
rect 3973 2088 3985 2091
rect 3384 2060 3985 2088
rect 3384 2048 3390 2060
rect 3973 2057 3985 2060
rect 4019 2088 4031 2091
rect 5166 2088 5172 2100
rect 4019 2060 5172 2088
rect 4019 2057 4031 2060
rect 3973 2051 4031 2057
rect 5166 2048 5172 2060
rect 5224 2048 5230 2100
rect 7466 2088 7472 2100
rect 5644 2060 7472 2088
rect 2590 1980 2596 2032
rect 2648 1980 2654 2032
rect 4893 2023 4951 2029
rect 4893 1989 4905 2023
rect 4939 2020 4951 2023
rect 4939 1992 5120 2020
rect 4939 1989 4951 1992
rect 4893 1983 4951 1989
rect 2038 1912 2044 1964
rect 2096 1952 2102 1964
rect 2498 1952 2504 1964
rect 2096 1924 2504 1952
rect 2096 1912 2102 1924
rect 2498 1912 2504 1924
rect 2556 1912 2562 1964
rect 3510 1912 3516 1964
rect 3568 1952 3574 1964
rect 3697 1955 3755 1961
rect 3697 1952 3709 1955
rect 3568 1924 3709 1952
rect 3568 1912 3574 1924
rect 3697 1921 3709 1924
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 5092 1961 5120 1992
rect 5534 1980 5540 2032
rect 5592 1980 5598 2032
rect 5644 1961 5672 2060
rect 7466 2048 7472 2060
rect 7524 2048 7530 2100
rect 7742 2048 7748 2100
rect 7800 2088 7806 2100
rect 8205 2091 8263 2097
rect 8205 2088 8217 2091
rect 7800 2060 8217 2088
rect 7800 2048 7806 2060
rect 8205 2057 8217 2060
rect 8251 2057 8263 2091
rect 8205 2051 8263 2057
rect 9769 2091 9827 2097
rect 9769 2057 9781 2091
rect 9815 2088 9827 2091
rect 10410 2088 10416 2100
rect 9815 2060 10416 2088
rect 9815 2057 9827 2060
rect 9769 2051 9827 2057
rect 10410 2048 10416 2060
rect 10468 2048 10474 2100
rect 9398 1980 9404 2032
rect 9456 2020 9462 2032
rect 9456 1992 11008 2020
rect 9456 1980 9462 1992
rect 4433 1955 4491 1961
rect 4433 1952 4445 1955
rect 4212 1924 4445 1952
rect 4212 1912 4218 1924
rect 4433 1921 4445 1924
rect 4479 1921 4491 1955
rect 4433 1915 4491 1921
rect 5077 1955 5135 1961
rect 5077 1921 5089 1955
rect 5123 1921 5135 1955
rect 5077 1915 5135 1921
rect 5629 1955 5687 1961
rect 5629 1921 5641 1955
rect 5675 1921 5687 1955
rect 10594 1952 10600 1964
rect 5629 1915 5687 1921
rect 9416 1924 10600 1952
rect 2225 1887 2283 1893
rect 2225 1853 2237 1887
rect 2271 1853 2283 1887
rect 2225 1847 2283 1853
rect 2317 1887 2375 1893
rect 2317 1853 2329 1887
rect 2363 1884 2375 1887
rect 2682 1884 2688 1896
rect 2363 1856 2688 1884
rect 2363 1853 2375 1856
rect 2317 1847 2375 1853
rect 2240 1748 2268 1847
rect 2682 1844 2688 1856
rect 2740 1884 2746 1896
rect 2869 1887 2927 1893
rect 2869 1884 2881 1887
rect 2740 1856 2881 1884
rect 2740 1844 2746 1856
rect 2869 1853 2881 1856
rect 2915 1853 2927 1887
rect 2869 1847 2927 1853
rect 3418 1844 3424 1896
rect 3476 1844 3482 1896
rect 3602 1844 3608 1896
rect 3660 1844 3666 1896
rect 3786 1844 3792 1896
rect 3844 1884 3850 1896
rect 4525 1887 4583 1893
rect 4525 1884 4537 1887
rect 3844 1856 4537 1884
rect 3844 1844 3850 1856
rect 4525 1853 4537 1856
rect 4571 1853 4583 1887
rect 4525 1847 4583 1853
rect 2501 1819 2559 1825
rect 2501 1785 2513 1819
rect 2547 1816 2559 1819
rect 2593 1819 2651 1825
rect 2593 1816 2605 1819
rect 2547 1788 2605 1816
rect 2547 1785 2559 1788
rect 2501 1779 2559 1785
rect 2593 1785 2605 1788
rect 2639 1785 2651 1819
rect 4540 1816 4568 1847
rect 5166 1844 5172 1896
rect 5224 1844 5230 1896
rect 5810 1844 5816 1896
rect 5868 1844 5874 1896
rect 5997 1887 6055 1893
rect 5997 1853 6009 1887
rect 6043 1884 6055 1887
rect 6273 1887 6331 1893
rect 6273 1884 6285 1887
rect 6043 1856 6285 1884
rect 6043 1853 6055 1856
rect 5997 1847 6055 1853
rect 6273 1853 6285 1856
rect 6319 1884 6331 1887
rect 6362 1884 6368 1896
rect 6319 1856 6368 1884
rect 6319 1853 6331 1856
rect 6273 1847 6331 1853
rect 6362 1844 6368 1856
rect 6420 1844 6426 1896
rect 6549 1887 6607 1893
rect 6549 1853 6561 1887
rect 6595 1853 6607 1887
rect 6549 1847 6607 1853
rect 5902 1816 5908 1828
rect 4540 1788 5908 1816
rect 2593 1779 2651 1785
rect 5902 1776 5908 1788
rect 5960 1776 5966 1828
rect 2777 1751 2835 1757
rect 2777 1748 2789 1751
rect 2240 1720 2789 1748
rect 2777 1717 2789 1720
rect 2823 1748 2835 1751
rect 3326 1748 3332 1760
rect 2823 1720 3332 1748
rect 2823 1717 2835 1720
rect 2777 1711 2835 1717
rect 3326 1708 3332 1720
rect 3384 1708 3390 1760
rect 4890 1708 4896 1760
rect 4948 1748 4954 1760
rect 6089 1751 6147 1757
rect 6089 1748 6101 1751
rect 4948 1720 6101 1748
rect 4948 1708 4954 1720
rect 6089 1717 6101 1720
rect 6135 1717 6147 1751
rect 6564 1748 6592 1847
rect 6638 1844 6644 1896
rect 6696 1884 6702 1896
rect 6733 1887 6791 1893
rect 6733 1884 6745 1887
rect 6696 1856 6745 1884
rect 6696 1844 6702 1856
rect 6733 1853 6745 1856
rect 6779 1853 6791 1887
rect 6733 1847 6791 1853
rect 6825 1887 6883 1893
rect 6825 1853 6837 1887
rect 6871 1884 6883 1887
rect 8389 1887 8447 1893
rect 8389 1884 8401 1887
rect 6871 1856 8401 1884
rect 6871 1853 6883 1856
rect 6825 1847 6883 1853
rect 8389 1853 8401 1856
rect 8435 1884 8447 1887
rect 9416 1884 9444 1924
rect 10594 1912 10600 1924
rect 10652 1912 10658 1964
rect 8435 1856 9444 1884
rect 8435 1853 8447 1856
rect 8389 1847 8447 1853
rect 9490 1844 9496 1896
rect 9548 1884 9554 1896
rect 10045 1887 10103 1893
rect 10045 1884 10057 1887
rect 9548 1856 10057 1884
rect 9548 1844 9554 1856
rect 10045 1853 10057 1856
rect 10091 1853 10103 1887
rect 10045 1847 10103 1853
rect 10321 1887 10379 1893
rect 10321 1853 10333 1887
rect 10367 1853 10379 1887
rect 10321 1847 10379 1853
rect 7092 1819 7150 1825
rect 7092 1785 7104 1819
rect 7138 1816 7150 1819
rect 7190 1816 7196 1828
rect 7138 1788 7196 1816
rect 7138 1785 7150 1788
rect 7092 1779 7150 1785
rect 7190 1776 7196 1788
rect 7248 1776 7254 1828
rect 7466 1776 7472 1828
rect 7524 1816 7530 1828
rect 8478 1816 8484 1828
rect 7524 1788 8484 1816
rect 7524 1776 7530 1788
rect 8478 1776 8484 1788
rect 8536 1776 8542 1828
rect 8662 1825 8668 1828
rect 8656 1816 8668 1825
rect 8623 1788 8668 1816
rect 8656 1779 8668 1788
rect 8662 1776 8668 1779
rect 8720 1776 8726 1828
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 9950 1816 9956 1828
rect 9732 1788 9956 1816
rect 9732 1776 9738 1788
rect 9950 1776 9956 1788
rect 10008 1816 10014 1828
rect 10336 1816 10364 1847
rect 10410 1844 10416 1896
rect 10468 1884 10474 1896
rect 10505 1887 10563 1893
rect 10505 1884 10517 1887
rect 10468 1856 10517 1884
rect 10468 1844 10474 1856
rect 10505 1853 10517 1856
rect 10551 1853 10563 1887
rect 10505 1847 10563 1853
rect 10008 1788 10364 1816
rect 10520 1816 10548 1847
rect 10778 1844 10784 1896
rect 10836 1844 10842 1896
rect 10980 1893 11008 1992
rect 10965 1887 11023 1893
rect 10965 1853 10977 1887
rect 11011 1884 11023 1887
rect 11057 1887 11115 1893
rect 11057 1884 11069 1887
rect 11011 1856 11069 1884
rect 11011 1853 11023 1856
rect 10965 1847 11023 1853
rect 11057 1853 11069 1856
rect 11103 1853 11115 1887
rect 11057 1847 11115 1853
rect 11238 1844 11244 1896
rect 11296 1844 11302 1896
rect 11149 1819 11207 1825
rect 11149 1816 11161 1819
rect 10520 1788 11161 1816
rect 10008 1776 10014 1788
rect 11149 1785 11161 1788
rect 11195 1785 11207 1819
rect 11149 1779 11207 1785
rect 6822 1748 6828 1760
rect 6564 1720 6828 1748
rect 6089 1711 6147 1717
rect 6822 1708 6828 1720
rect 6880 1748 6886 1760
rect 9861 1751 9919 1757
rect 9861 1748 9873 1751
rect 6880 1720 9873 1748
rect 6880 1708 6886 1720
rect 9861 1717 9873 1720
rect 9907 1717 9919 1751
rect 9861 1711 9919 1717
rect 10410 1708 10416 1760
rect 10468 1748 10474 1760
rect 10597 1751 10655 1757
rect 10597 1748 10609 1751
rect 10468 1720 10609 1748
rect 10468 1708 10474 1720
rect 10597 1717 10609 1720
rect 10643 1717 10655 1751
rect 10597 1711 10655 1717
rect 552 1658 12604 1680
rect 552 1606 4322 1658
rect 4374 1606 4386 1658
rect 4438 1606 4450 1658
rect 4502 1606 4514 1658
rect 4566 1606 4578 1658
rect 4630 1606 10722 1658
rect 10774 1606 10786 1658
rect 10838 1606 10850 1658
rect 10902 1606 10914 1658
rect 10966 1606 10978 1658
rect 11030 1606 12604 1658
rect 552 1584 12604 1606
rect 3145 1547 3203 1553
rect 3145 1513 3157 1547
rect 3191 1544 3203 1547
rect 3786 1544 3792 1556
rect 3191 1516 3792 1544
rect 3191 1513 3203 1516
rect 3145 1507 3203 1513
rect 3786 1504 3792 1516
rect 3844 1504 3850 1556
rect 5166 1504 5172 1556
rect 5224 1544 5230 1556
rect 5261 1547 5319 1553
rect 5261 1544 5273 1547
rect 5224 1516 5273 1544
rect 5224 1504 5230 1516
rect 5261 1513 5273 1516
rect 5307 1513 5319 1547
rect 5261 1507 5319 1513
rect 7282 1504 7288 1556
rect 7340 1544 7346 1556
rect 7377 1547 7435 1553
rect 7377 1544 7389 1547
rect 7340 1516 7389 1544
rect 7340 1504 7346 1516
rect 7377 1513 7389 1516
rect 7423 1513 7435 1547
rect 7377 1507 7435 1513
rect 7558 1504 7564 1556
rect 7616 1544 7622 1556
rect 8110 1544 8116 1556
rect 7616 1516 8116 1544
rect 7616 1504 7622 1516
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 8294 1504 8300 1556
rect 8352 1544 8358 1556
rect 8389 1547 8447 1553
rect 8389 1544 8401 1547
rect 8352 1516 8401 1544
rect 8352 1504 8358 1516
rect 8389 1513 8401 1516
rect 8435 1513 8447 1547
rect 8389 1507 8447 1513
rect 8570 1504 8576 1556
rect 8628 1504 8634 1556
rect 9309 1547 9367 1553
rect 8671 1516 9076 1544
rect 2032 1479 2090 1485
rect 2032 1445 2044 1479
rect 2078 1476 2090 1479
rect 2590 1476 2596 1488
rect 2078 1448 2596 1476
rect 2078 1445 2090 1448
rect 2032 1439 2090 1445
rect 2590 1436 2596 1448
rect 2648 1436 2654 1488
rect 4264 1448 5672 1476
rect 4264 1420 4292 1448
rect 3510 1368 3516 1420
rect 3568 1408 3574 1420
rect 3605 1411 3663 1417
rect 3605 1408 3617 1411
rect 3568 1380 3617 1408
rect 3568 1368 3574 1380
rect 3605 1377 3617 1380
rect 3651 1377 3663 1411
rect 3605 1371 3663 1377
rect 4246 1368 4252 1420
rect 4304 1368 4310 1420
rect 4890 1368 4896 1420
rect 4948 1368 4954 1420
rect 5442 1368 5448 1420
rect 5500 1398 5506 1420
rect 5644 1417 5672 1448
rect 6546 1436 6552 1488
rect 6604 1476 6610 1488
rect 8671 1476 8699 1516
rect 6604 1448 8699 1476
rect 6604 1436 6610 1448
rect 5629 1411 5687 1417
rect 5500 1370 5535 1398
rect 5629 1377 5641 1411
rect 5675 1377 5687 1411
rect 5629 1371 5687 1377
rect 5997 1411 6055 1417
rect 5997 1377 6009 1411
rect 6043 1377 6055 1411
rect 5997 1371 6055 1377
rect 6273 1411 6331 1417
rect 6273 1377 6285 1411
rect 6319 1408 6331 1411
rect 6454 1408 6460 1420
rect 6319 1380 6460 1408
rect 6319 1377 6331 1380
rect 6273 1371 6331 1377
rect 5500 1368 5506 1370
rect 5445 1367 5457 1368
rect 5491 1367 5503 1368
rect 5445 1361 5503 1367
rect 1394 1300 1400 1352
rect 1452 1340 1458 1352
rect 1765 1343 1823 1349
rect 1765 1340 1777 1343
rect 1452 1312 1777 1340
rect 1452 1300 1458 1312
rect 1765 1309 1777 1312
rect 1811 1309 1823 1343
rect 1765 1303 1823 1309
rect 3697 1343 3755 1349
rect 3697 1309 3709 1343
rect 3743 1309 3755 1343
rect 3697 1303 3755 1309
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 3712 1272 3740 1303
rect 4062 1300 4068 1352
rect 4120 1340 4126 1352
rect 4157 1343 4215 1349
rect 4157 1340 4169 1343
rect 4120 1312 4169 1340
rect 4120 1300 4126 1312
rect 4157 1309 4169 1312
rect 4203 1309 4215 1343
rect 4157 1303 4215 1309
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1340 4675 1343
rect 4801 1343 4859 1349
rect 4801 1340 4813 1343
rect 4663 1312 4813 1340
rect 4663 1309 4675 1312
rect 4617 1303 4675 1309
rect 4801 1309 4813 1312
rect 4847 1309 4859 1343
rect 6012 1340 6040 1371
rect 6454 1368 6460 1380
rect 6512 1368 6518 1420
rect 4801 1303 4859 1309
rect 5920 1312 6040 1340
rect 6181 1343 6239 1349
rect 5813 1275 5871 1281
rect 5813 1272 5825 1275
rect 3660 1244 5825 1272
rect 3660 1232 3666 1244
rect 5813 1241 5825 1244
rect 5859 1241 5871 1275
rect 5813 1235 5871 1241
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1204 4031 1207
rect 4798 1204 4804 1216
rect 4019 1176 4804 1204
rect 4019 1173 4031 1176
rect 3973 1167 4031 1173
rect 4798 1164 4804 1176
rect 4856 1164 4862 1216
rect 5537 1207 5595 1213
rect 5537 1173 5549 1207
rect 5583 1204 5595 1207
rect 5920 1204 5948 1312
rect 6181 1309 6193 1343
rect 6227 1340 6239 1343
rect 6656 1340 6684 1448
rect 8938 1436 8944 1488
rect 8996 1436 9002 1488
rect 9048 1476 9076 1516
rect 9309 1513 9321 1547
rect 9355 1544 9367 1547
rect 9490 1544 9496 1556
rect 9355 1516 9496 1544
rect 9355 1513 9367 1516
rect 9309 1507 9367 1513
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 10410 1504 10416 1556
rect 10468 1504 10474 1556
rect 10594 1504 10600 1556
rect 10652 1504 10658 1556
rect 10428 1476 10456 1504
rect 9048 1448 10272 1476
rect 10428 1448 10824 1476
rect 6730 1368 6736 1420
rect 6788 1368 6794 1420
rect 7558 1368 7564 1420
rect 7616 1368 7622 1420
rect 7650 1368 7656 1420
rect 7708 1408 7714 1420
rect 7929 1411 7987 1417
rect 7708 1380 7880 1408
rect 7708 1368 7714 1380
rect 6227 1312 6684 1340
rect 6227 1309 6239 1312
rect 6181 1303 6239 1309
rect 6822 1300 6828 1352
rect 6880 1300 6886 1352
rect 7374 1300 7380 1352
rect 7432 1300 7438 1352
rect 7466 1300 7472 1352
rect 7524 1340 7530 1352
rect 7745 1343 7803 1349
rect 7745 1340 7757 1343
rect 7524 1312 7757 1340
rect 7524 1300 7530 1312
rect 7745 1309 7757 1312
rect 7791 1309 7803 1343
rect 7745 1303 7803 1309
rect 6086 1204 6092 1216
rect 5583 1176 6092 1204
rect 5583 1173 5595 1176
rect 5537 1167 5595 1173
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 7006 1164 7012 1216
rect 7064 1164 7070 1216
rect 7392 1204 7420 1300
rect 7852 1272 7880 1380
rect 7929 1377 7941 1411
rect 7975 1377 7987 1411
rect 7929 1371 7987 1377
rect 7944 1340 7972 1371
rect 8202 1368 8208 1420
rect 8260 1368 8266 1420
rect 8478 1368 8484 1420
rect 8536 1408 8542 1420
rect 8849 1411 8907 1417
rect 8849 1408 8861 1411
rect 8536 1380 8861 1408
rect 8536 1368 8542 1380
rect 8849 1377 8861 1380
rect 8895 1377 8907 1411
rect 8956 1408 8984 1436
rect 9125 1411 9183 1417
rect 9125 1408 9137 1411
rect 8956 1380 9137 1408
rect 8849 1371 8907 1377
rect 9125 1377 9137 1380
rect 9171 1408 9183 1411
rect 9398 1408 9404 1420
rect 9171 1380 9404 1408
rect 9171 1377 9183 1380
rect 9125 1371 9183 1377
rect 9398 1368 9404 1380
rect 9456 1368 9462 1420
rect 9582 1368 9588 1420
rect 9640 1368 9646 1420
rect 9766 1368 9772 1420
rect 9824 1408 9830 1420
rect 10244 1417 10272 1448
rect 10045 1411 10103 1417
rect 10045 1408 10057 1411
rect 9824 1380 10057 1408
rect 9824 1368 9830 1380
rect 10045 1377 10057 1380
rect 10091 1377 10103 1411
rect 10045 1371 10103 1377
rect 10229 1411 10287 1417
rect 10229 1377 10241 1411
rect 10275 1377 10287 1411
rect 10229 1371 10287 1377
rect 8386 1340 8392 1352
rect 7944 1312 8392 1340
rect 8386 1300 8392 1312
rect 8444 1300 8450 1352
rect 8573 1343 8631 1349
rect 8573 1309 8585 1343
rect 8619 1309 8631 1343
rect 8573 1303 8631 1309
rect 8941 1343 8999 1349
rect 8941 1309 8953 1343
rect 8987 1340 8999 1343
rect 9030 1340 9036 1352
rect 8987 1312 9036 1340
rect 8987 1309 8999 1312
rect 8941 1303 8999 1309
rect 8294 1272 8300 1284
rect 7852 1244 8300 1272
rect 8294 1232 8300 1244
rect 8352 1232 8358 1284
rect 8588 1204 8616 1303
rect 9030 1300 9036 1312
rect 9088 1300 9094 1352
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 10060 1340 10088 1371
rect 10502 1368 10508 1420
rect 10560 1368 10566 1420
rect 10796 1417 10824 1448
rect 10597 1411 10655 1417
rect 10597 1377 10609 1411
rect 10643 1377 10655 1411
rect 10597 1371 10655 1377
rect 10781 1411 10839 1417
rect 10781 1377 10793 1411
rect 10827 1377 10839 1411
rect 10781 1371 10839 1377
rect 10612 1340 10640 1371
rect 10060 1312 10640 1340
rect 8754 1232 8760 1284
rect 8812 1272 8818 1284
rect 9306 1272 9312 1284
rect 8812 1244 9312 1272
rect 8812 1232 8818 1244
rect 9306 1232 9312 1244
rect 9364 1232 9370 1284
rect 11422 1272 11428 1284
rect 9646 1244 11428 1272
rect 9646 1204 9674 1244
rect 11422 1232 11428 1244
rect 11480 1232 11486 1284
rect 7392 1176 9674 1204
rect 9858 1164 9864 1216
rect 9916 1164 9922 1216
rect 552 1114 12604 1136
rect 552 1062 3662 1114
rect 3714 1062 3726 1114
rect 3778 1062 3790 1114
rect 3842 1062 3854 1114
rect 3906 1062 3918 1114
rect 3970 1062 10062 1114
rect 10114 1062 10126 1114
rect 10178 1062 10190 1114
rect 10242 1062 10254 1114
rect 10306 1062 10318 1114
rect 10370 1062 12604 1114
rect 552 1040 12604 1062
rect 3510 960 3516 1012
rect 3568 1000 3574 1012
rect 3789 1003 3847 1009
rect 3789 1000 3801 1003
rect 3568 972 3801 1000
rect 3568 960 3574 972
rect 3789 969 3801 972
rect 3835 969 3847 1003
rect 3789 963 3847 969
rect 6181 1003 6239 1009
rect 6181 969 6193 1003
rect 6227 1000 6239 1003
rect 6454 1000 6460 1012
rect 6227 972 6460 1000
rect 6227 969 6239 972
rect 6181 963 6239 969
rect 6454 960 6460 972
rect 6512 960 6518 1012
rect 6638 960 6644 1012
rect 6696 960 6702 1012
rect 9582 960 9588 1012
rect 9640 960 9646 1012
rect 3418 824 3424 876
rect 3476 864 3482 876
rect 4065 867 4123 873
rect 4065 864 4077 867
rect 3476 836 4077 864
rect 3476 824 3482 836
rect 2774 756 2780 808
rect 2832 796 2838 808
rect 3896 805 3924 836
rect 4065 833 4077 836
rect 4111 833 4123 867
rect 4065 827 4123 833
rect 5534 824 5540 876
rect 5592 864 5598 876
rect 5592 836 6684 864
rect 5592 824 5598 836
rect 3237 799 3295 805
rect 3237 796 3249 799
rect 2832 768 3249 796
rect 2832 756 2838 768
rect 3237 765 3249 768
rect 3283 796 3295 799
rect 3605 799 3663 805
rect 3283 768 3556 796
rect 3283 765 3295 768
rect 3237 759 3295 765
rect 3326 688 3332 740
rect 3384 728 3390 740
rect 3421 731 3479 737
rect 3421 728 3433 731
rect 3384 700 3433 728
rect 3384 688 3390 700
rect 3421 697 3433 700
rect 3467 697 3479 731
rect 3528 728 3556 768
rect 3605 765 3617 799
rect 3651 796 3663 799
rect 3697 799 3755 805
rect 3697 796 3709 799
rect 3651 768 3709 796
rect 3651 765 3663 768
rect 3605 759 3663 765
rect 3697 765 3709 768
rect 3743 765 3755 799
rect 3697 759 3755 765
rect 3881 799 3939 805
rect 3881 765 3893 799
rect 3927 765 3939 799
rect 3881 759 3939 765
rect 3970 756 3976 808
rect 4028 756 4034 808
rect 4157 799 4215 805
rect 4157 765 4169 799
rect 4203 765 4215 799
rect 4157 759 4215 765
rect 4062 728 4068 740
rect 3528 700 4068 728
rect 3421 691 3479 697
rect 3436 660 3464 691
rect 4062 688 4068 700
rect 4120 728 4126 740
rect 4172 728 4200 759
rect 6086 756 6092 808
rect 6144 756 6150 808
rect 6270 756 6276 808
rect 6328 756 6334 808
rect 6656 805 6684 836
rect 6641 799 6699 805
rect 6641 765 6653 799
rect 6687 765 6699 799
rect 6641 759 6699 765
rect 6825 799 6883 805
rect 6825 765 6837 799
rect 6871 796 6883 799
rect 7466 796 7472 808
rect 6871 768 7472 796
rect 6871 765 6883 768
rect 6825 759 6883 765
rect 7466 756 7472 768
rect 7524 756 7530 808
rect 9401 799 9459 805
rect 9401 765 9413 799
rect 9447 796 9459 799
rect 9490 796 9496 808
rect 9447 768 9496 796
rect 9447 765 9459 768
rect 9401 759 9459 765
rect 9490 756 9496 768
rect 9548 756 9554 808
rect 9585 799 9643 805
rect 9585 765 9597 799
rect 9631 796 9643 799
rect 10410 796 10416 808
rect 9631 768 10416 796
rect 9631 765 9643 768
rect 9585 759 9643 765
rect 10410 756 10416 768
rect 10468 756 10474 808
rect 4120 700 4200 728
rect 4120 688 4126 700
rect 3970 660 3976 672
rect 3436 632 3976 660
rect 3970 620 3976 632
rect 4028 620 4034 672
rect 552 570 12604 592
rect 552 518 4322 570
rect 4374 518 4386 570
rect 4438 518 4450 570
rect 4502 518 4514 570
rect 4566 518 4578 570
rect 4630 518 10722 570
rect 10774 518 10786 570
rect 10838 518 10850 570
rect 10902 518 10914 570
rect 10966 518 10978 570
rect 11030 518 12604 570
rect 552 496 12604 518
<< via1 >>
rect 7196 43324 7248 43376
rect 10048 43324 10100 43376
rect 2964 43120 3016 43172
rect 8668 43120 8720 43172
rect 7472 43052 7524 43104
rect 9956 43052 10008 43104
rect 4322 42950 4374 43002
rect 4386 42950 4438 43002
rect 4450 42950 4502 43002
rect 4514 42950 4566 43002
rect 4578 42950 4630 43002
rect 10722 42950 10774 43002
rect 10786 42950 10838 43002
rect 10850 42950 10902 43002
rect 10914 42950 10966 43002
rect 10978 42950 11030 43002
rect 8300 42848 8352 42900
rect 6644 42780 6696 42832
rect 20 42712 72 42764
rect 1308 42712 1360 42764
rect 1492 42755 1544 42764
rect 1492 42721 1526 42755
rect 1526 42721 1544 42755
rect 1492 42712 1544 42721
rect 4252 42712 4304 42764
rect 5356 42712 5408 42764
rect 6184 42712 6236 42764
rect 6276 42712 6328 42764
rect 7748 42780 7800 42832
rect 7472 42755 7524 42764
rect 7472 42721 7476 42755
rect 7476 42721 7510 42755
rect 7510 42721 7524 42755
rect 7472 42712 7524 42721
rect 7932 42755 7984 42764
rect 7932 42721 7941 42755
rect 7941 42721 7975 42755
rect 7975 42721 7984 42755
rect 7932 42712 7984 42721
rect 8024 42755 8076 42764
rect 8024 42721 8033 42755
rect 8033 42721 8067 42755
rect 8067 42721 8076 42755
rect 8024 42712 8076 42721
rect 3148 42576 3200 42628
rect 4896 42644 4948 42696
rect 5264 42644 5316 42696
rect 7288 42644 7340 42696
rect 8116 42644 8168 42696
rect 8300 42644 8352 42696
rect 8484 42755 8536 42764
rect 8484 42721 8494 42755
rect 8494 42721 8528 42755
rect 8528 42721 8536 42755
rect 8484 42712 8536 42721
rect 8668 42755 8720 42764
rect 8668 42721 8677 42755
rect 8677 42721 8711 42755
rect 8711 42721 8720 42755
rect 8668 42712 8720 42721
rect 9036 42780 9088 42832
rect 10048 42755 10100 42764
rect 10048 42721 10057 42755
rect 10057 42721 10091 42755
rect 10091 42721 10100 42755
rect 10048 42712 10100 42721
rect 10784 42712 10836 42764
rect 11152 42712 11204 42764
rect 11704 42780 11756 42832
rect 9680 42687 9732 42696
rect 9680 42653 9689 42687
rect 9689 42653 9723 42687
rect 9723 42653 9732 42687
rect 9680 42644 9732 42653
rect 9772 42644 9824 42696
rect 940 42551 992 42560
rect 940 42517 949 42551
rect 949 42517 983 42551
rect 983 42517 992 42551
rect 940 42508 992 42517
rect 2596 42551 2648 42560
rect 2596 42517 2605 42551
rect 2605 42517 2639 42551
rect 2639 42517 2648 42551
rect 2596 42508 2648 42517
rect 2872 42551 2924 42560
rect 2872 42517 2881 42551
rect 2881 42517 2915 42551
rect 2915 42517 2924 42551
rect 2872 42508 2924 42517
rect 4068 42508 4120 42560
rect 5632 42551 5684 42560
rect 5632 42517 5641 42551
rect 5641 42517 5675 42551
rect 5675 42517 5684 42551
rect 5632 42508 5684 42517
rect 5816 42551 5868 42560
rect 5816 42517 5825 42551
rect 5825 42517 5859 42551
rect 5859 42517 5868 42551
rect 5816 42508 5868 42517
rect 6552 42551 6604 42560
rect 6552 42517 6561 42551
rect 6561 42517 6595 42551
rect 6595 42517 6604 42551
rect 6552 42508 6604 42517
rect 9404 42576 9456 42628
rect 10876 42576 10928 42628
rect 8208 42551 8260 42560
rect 8208 42517 8217 42551
rect 8217 42517 8251 42551
rect 8251 42517 8260 42551
rect 8208 42508 8260 42517
rect 8392 42508 8444 42560
rect 9128 42508 9180 42560
rect 10968 42508 11020 42560
rect 11244 42619 11296 42628
rect 11244 42585 11253 42619
rect 11253 42585 11287 42619
rect 11287 42585 11296 42619
rect 11244 42576 11296 42585
rect 12072 42712 12124 42764
rect 12164 42644 12216 42696
rect 11796 42551 11848 42560
rect 11796 42517 11805 42551
rect 11805 42517 11839 42551
rect 11839 42517 11848 42551
rect 11796 42508 11848 42517
rect 11888 42508 11940 42560
rect 12440 42508 12492 42560
rect 3662 42406 3714 42458
rect 3726 42406 3778 42458
rect 3790 42406 3842 42458
rect 3854 42406 3906 42458
rect 3918 42406 3970 42458
rect 10062 42406 10114 42458
rect 10126 42406 10178 42458
rect 10190 42406 10242 42458
rect 10254 42406 10306 42458
rect 10318 42406 10370 42458
rect 848 42143 900 42152
rect 848 42109 857 42143
rect 857 42109 891 42143
rect 891 42109 900 42143
rect 848 42100 900 42109
rect 1032 42143 1084 42152
rect 1032 42109 1039 42143
rect 1039 42109 1084 42143
rect 1032 42100 1084 42109
rect 2964 42347 3016 42356
rect 2964 42313 2973 42347
rect 2973 42313 3007 42347
rect 3007 42313 3016 42347
rect 2964 42304 3016 42313
rect 4160 42304 4212 42356
rect 5264 42347 5316 42356
rect 5264 42313 5273 42347
rect 5273 42313 5307 42347
rect 5307 42313 5316 42347
rect 5264 42304 5316 42313
rect 5356 42304 5408 42356
rect 5724 42304 5776 42356
rect 6920 42304 6972 42356
rect 8392 42304 8444 42356
rect 9128 42304 9180 42356
rect 3792 42236 3844 42288
rect 7840 42279 7892 42288
rect 7840 42245 7845 42279
rect 7845 42245 7879 42279
rect 7879 42245 7892 42279
rect 1216 42075 1268 42084
rect 1216 42041 1225 42075
rect 1225 42041 1259 42075
rect 1259 42041 1268 42075
rect 1216 42032 1268 42041
rect 1584 42143 1636 42152
rect 1584 42109 1593 42143
rect 1593 42109 1627 42143
rect 1627 42109 1636 42143
rect 1584 42100 1636 42109
rect 2136 42100 2188 42152
rect 3976 42100 4028 42152
rect 4252 42168 4304 42220
rect 7840 42236 7892 42245
rect 4160 42143 4212 42152
rect 4160 42109 4170 42143
rect 4170 42109 4204 42143
rect 4204 42109 4212 42143
rect 4160 42100 4212 42109
rect 4344 42143 4396 42152
rect 4344 42109 4353 42143
rect 4353 42109 4387 42143
rect 4387 42109 4396 42143
rect 4344 42100 4396 42109
rect 1860 42075 1912 42084
rect 1860 42041 1894 42075
rect 1894 42041 1912 42075
rect 1860 42032 1912 42041
rect 3148 42032 3200 42084
rect 2872 41964 2924 42016
rect 4160 41964 4212 42016
rect 4804 42143 4856 42152
rect 4804 42109 4813 42143
rect 4813 42109 4847 42143
rect 4847 42109 4856 42143
rect 4804 42100 4856 42109
rect 5080 42143 5132 42152
rect 5080 42109 5089 42143
rect 5089 42109 5123 42143
rect 5123 42109 5132 42143
rect 5080 42100 5132 42109
rect 5172 42100 5224 42152
rect 5264 42032 5316 42084
rect 6552 42100 6604 42152
rect 6828 42032 6880 42084
rect 5448 41964 5500 42016
rect 6460 41964 6512 42016
rect 7196 42100 7248 42152
rect 7472 42100 7524 42152
rect 7748 42143 7800 42152
rect 7748 42109 7757 42143
rect 7757 42109 7791 42143
rect 7791 42109 7800 42143
rect 7748 42100 7800 42109
rect 7932 42143 7984 42152
rect 7932 42109 7941 42143
rect 7941 42109 7975 42143
rect 7975 42109 7984 42143
rect 7932 42100 7984 42109
rect 8116 42100 8168 42152
rect 8392 42100 8444 42152
rect 8760 42100 8812 42152
rect 9220 42100 9272 42152
rect 9772 42236 9824 42288
rect 10876 42279 10928 42288
rect 10876 42245 10885 42279
rect 10885 42245 10919 42279
rect 10919 42245 10928 42279
rect 10876 42236 10928 42245
rect 9956 42100 10008 42152
rect 10600 42100 10652 42152
rect 12256 42143 12308 42152
rect 12256 42109 12265 42143
rect 12265 42109 12299 42143
rect 12299 42109 12308 42143
rect 12256 42100 12308 42109
rect 7012 42032 7064 42084
rect 8024 42032 8076 42084
rect 8852 42075 8904 42084
rect 8852 42041 8861 42075
rect 8861 42041 8895 42075
rect 8895 42041 8904 42075
rect 8852 42032 8904 42041
rect 8944 42075 8996 42084
rect 8944 42041 8953 42075
rect 8953 42041 8987 42075
rect 8987 42041 8996 42075
rect 8944 42032 8996 42041
rect 7564 41964 7616 42016
rect 8116 42007 8168 42016
rect 8116 41973 8125 42007
rect 8125 41973 8159 42007
rect 8159 41973 8168 42007
rect 8116 41964 8168 41973
rect 8484 41964 8536 42016
rect 10416 42075 10468 42084
rect 10416 42041 10425 42075
rect 10425 42041 10459 42075
rect 10459 42041 10468 42075
rect 10416 42032 10468 42041
rect 10784 42032 10836 42084
rect 11520 42032 11572 42084
rect 9864 42007 9916 42016
rect 9864 41973 9873 42007
rect 9873 41973 9907 42007
rect 9907 41973 9916 42007
rect 9864 41964 9916 41973
rect 10048 42007 10100 42016
rect 10048 41973 10057 42007
rect 10057 41973 10091 42007
rect 10091 41973 10100 42007
rect 10048 41964 10100 41973
rect 10508 42007 10560 42016
rect 10508 41973 10517 42007
rect 10517 41973 10551 42007
rect 10551 41973 10560 42007
rect 10508 41964 10560 41973
rect 4322 41862 4374 41914
rect 4386 41862 4438 41914
rect 4450 41862 4502 41914
rect 4514 41862 4566 41914
rect 4578 41862 4630 41914
rect 10722 41862 10774 41914
rect 10786 41862 10838 41914
rect 10850 41862 10902 41914
rect 10914 41862 10966 41914
rect 10978 41862 11030 41914
rect 1032 41760 1084 41812
rect 1860 41760 1912 41812
rect 2596 41760 2648 41812
rect 4804 41760 4856 41812
rect 5632 41692 5684 41744
rect 6736 41692 6788 41744
rect 1032 41624 1084 41676
rect 1308 41624 1360 41676
rect 2320 41624 2372 41676
rect 2504 41667 2556 41676
rect 2504 41633 2538 41667
rect 2538 41633 2556 41667
rect 2504 41624 2556 41633
rect 2872 41624 2924 41676
rect 4160 41667 4212 41676
rect 4160 41633 4169 41667
rect 4169 41633 4203 41667
rect 4203 41633 4212 41667
rect 4160 41624 4212 41633
rect 5908 41624 5960 41676
rect 6000 41667 6052 41676
rect 6000 41633 6009 41667
rect 6009 41633 6043 41667
rect 6043 41633 6052 41667
rect 6000 41624 6052 41633
rect 7380 41692 7432 41744
rect 8484 41692 8536 41744
rect 9220 41803 9272 41812
rect 9220 41769 9229 41803
rect 9229 41769 9263 41803
rect 9263 41769 9272 41803
rect 9220 41760 9272 41769
rect 10784 41760 10836 41812
rect 11796 41760 11848 41812
rect 1492 41488 1544 41540
rect 3332 41556 3384 41608
rect 3792 41556 3844 41608
rect 4252 41599 4304 41608
rect 4252 41565 4261 41599
rect 4261 41565 4295 41599
rect 4295 41565 4304 41599
rect 4252 41556 4304 41565
rect 5724 41556 5776 41608
rect 8116 41624 8168 41676
rect 8668 41624 8720 41676
rect 10876 41692 10928 41744
rect 11060 41692 11112 41744
rect 6184 41556 6236 41608
rect 7196 41556 7248 41608
rect 1860 41420 1912 41472
rect 3976 41488 4028 41540
rect 3516 41420 3568 41472
rect 6368 41488 6420 41540
rect 9036 41488 9088 41540
rect 5632 41463 5684 41472
rect 5632 41429 5641 41463
rect 5641 41429 5675 41463
rect 5675 41429 5684 41463
rect 5632 41420 5684 41429
rect 7104 41420 7156 41472
rect 7196 41420 7248 41472
rect 8668 41420 8720 41472
rect 9404 41463 9456 41472
rect 9404 41429 9413 41463
rect 9413 41429 9447 41463
rect 9447 41429 9456 41463
rect 9404 41420 9456 41429
rect 10048 41420 10100 41472
rect 10600 41420 10652 41472
rect 11060 41556 11112 41608
rect 11520 41556 11572 41608
rect 10968 41463 11020 41472
rect 10968 41429 10977 41463
rect 10977 41429 11011 41463
rect 11011 41429 11020 41463
rect 10968 41420 11020 41429
rect 11520 41420 11572 41472
rect 12532 41420 12584 41472
rect 3662 41318 3714 41370
rect 3726 41318 3778 41370
rect 3790 41318 3842 41370
rect 3854 41318 3906 41370
rect 3918 41318 3970 41370
rect 10062 41318 10114 41370
rect 10126 41318 10178 41370
rect 10190 41318 10242 41370
rect 10254 41318 10306 41370
rect 10318 41318 10370 41370
rect 1216 41216 1268 41268
rect 2688 41216 2740 41268
rect 5080 41216 5132 41268
rect 6920 41216 6972 41268
rect 6644 41148 6696 41200
rect 6736 41148 6788 41200
rect 7748 41148 7800 41200
rect 8024 41191 8076 41200
rect 8024 41157 8033 41191
rect 8033 41157 8067 41191
rect 8067 41157 8076 41191
rect 8024 41148 8076 41157
rect 1124 41080 1176 41132
rect 1308 41080 1360 41132
rect 11520 41216 11572 41268
rect 1492 41012 1544 41064
rect 1768 41012 1820 41064
rect 2320 41012 2372 41064
rect 4252 41012 4304 41064
rect 5080 41012 5132 41064
rect 5908 41012 5960 41064
rect 6644 41012 6696 41064
rect 1400 40944 1452 40996
rect 3056 40987 3108 40996
rect 3056 40953 3065 40987
rect 3065 40953 3099 40987
rect 3099 40953 3108 40987
rect 3056 40944 3108 40953
rect 2136 40876 2188 40928
rect 2596 40876 2648 40928
rect 3424 40919 3476 40928
rect 3424 40885 3433 40919
rect 3433 40885 3467 40919
rect 3467 40885 3476 40919
rect 3424 40876 3476 40885
rect 4068 40944 4120 40996
rect 5816 40944 5868 40996
rect 6092 40944 6144 40996
rect 7196 41012 7248 41064
rect 7380 41012 7432 41064
rect 7472 41055 7524 41064
rect 7472 41021 7481 41055
rect 7481 41021 7515 41055
rect 7515 41021 7524 41055
rect 7472 41012 7524 41021
rect 7840 41080 7892 41132
rect 8116 41080 8168 41132
rect 7932 41012 7984 41064
rect 5172 40876 5224 40928
rect 5540 40876 5592 40928
rect 6000 40876 6052 40928
rect 6184 40876 6236 40928
rect 6828 40876 6880 40928
rect 7380 40876 7432 40928
rect 8944 41012 8996 41064
rect 8392 40987 8444 40996
rect 8392 40953 8401 40987
rect 8401 40953 8435 40987
rect 8435 40953 8444 40987
rect 8392 40944 8444 40953
rect 8852 40944 8904 40996
rect 8300 40876 8352 40928
rect 8484 40876 8536 40928
rect 9128 40876 9180 40928
rect 9312 41055 9364 41064
rect 9312 41021 9321 41055
rect 9321 41021 9355 41055
rect 9355 41021 9364 41055
rect 9312 41012 9364 41021
rect 12624 41080 12676 41132
rect 10508 41012 10560 41064
rect 10968 41012 11020 41064
rect 11152 41012 11204 41064
rect 12164 41055 12216 41064
rect 12164 41021 12173 41055
rect 12173 41021 12207 41055
rect 12207 41021 12216 41055
rect 12164 41012 12216 41021
rect 9956 40987 10008 40996
rect 9956 40953 9965 40987
rect 9965 40953 9999 40987
rect 9999 40953 10008 40987
rect 9956 40944 10008 40953
rect 10048 40944 10100 40996
rect 11796 40944 11848 40996
rect 11152 40876 11204 40928
rect 4322 40774 4374 40826
rect 4386 40774 4438 40826
rect 4450 40774 4502 40826
rect 4514 40774 4566 40826
rect 4578 40774 4630 40826
rect 10722 40774 10774 40826
rect 10786 40774 10838 40826
rect 10850 40774 10902 40826
rect 10914 40774 10966 40826
rect 10978 40774 11030 40826
rect 1216 40715 1268 40724
rect 1216 40681 1225 40715
rect 1225 40681 1259 40715
rect 1259 40681 1268 40715
rect 1216 40672 1268 40681
rect 1400 40672 1452 40724
rect 2504 40672 2556 40724
rect 4160 40672 4212 40724
rect 3240 40604 3292 40656
rect 3516 40604 3568 40656
rect 1308 40536 1360 40588
rect 2320 40579 2372 40588
rect 2320 40545 2329 40579
rect 2329 40545 2363 40579
rect 2363 40545 2372 40579
rect 2320 40536 2372 40545
rect 2412 40536 2464 40588
rect 4160 40579 4212 40588
rect 4160 40545 4169 40579
rect 4169 40545 4203 40579
rect 4203 40545 4212 40579
rect 4160 40536 4212 40545
rect 4252 40579 4304 40588
rect 4252 40545 4261 40579
rect 4261 40545 4295 40579
rect 4295 40545 4304 40579
rect 4252 40536 4304 40545
rect 2136 40511 2188 40520
rect 2136 40477 2145 40511
rect 2145 40477 2179 40511
rect 2179 40477 2188 40511
rect 2136 40468 2188 40477
rect 3332 40468 3384 40520
rect 4528 40579 4580 40588
rect 4528 40545 4537 40579
rect 4537 40545 4571 40579
rect 4571 40545 4580 40579
rect 4988 40604 5040 40656
rect 8668 40672 8720 40724
rect 11520 40672 11572 40724
rect 5540 40604 5592 40656
rect 4528 40536 4580 40545
rect 1492 40400 1544 40452
rect 1768 40443 1820 40452
rect 1768 40409 1777 40443
rect 1777 40409 1811 40443
rect 1811 40409 1820 40443
rect 1768 40400 1820 40409
rect 2228 40332 2280 40384
rect 4252 40400 4304 40452
rect 4620 40468 4672 40520
rect 5264 40579 5316 40588
rect 5264 40545 5278 40579
rect 5278 40545 5312 40579
rect 5312 40545 5316 40579
rect 5264 40536 5316 40545
rect 5448 40536 5500 40588
rect 6184 40536 6236 40588
rect 6828 40604 6880 40656
rect 7104 40604 7156 40656
rect 6644 40579 6696 40588
rect 6644 40545 6653 40579
rect 6653 40545 6687 40579
rect 6687 40545 6696 40579
rect 6644 40536 6696 40545
rect 7380 40579 7432 40588
rect 7380 40545 7389 40579
rect 7389 40545 7423 40579
rect 7423 40545 7432 40579
rect 7380 40536 7432 40545
rect 7656 40604 7708 40656
rect 8024 40604 8076 40656
rect 8208 40604 8260 40656
rect 9864 40604 9916 40656
rect 7472 40468 7524 40520
rect 9128 40579 9180 40588
rect 9128 40545 9137 40579
rect 9137 40545 9171 40579
rect 9171 40545 9180 40579
rect 9128 40536 9180 40545
rect 9220 40536 9272 40588
rect 9588 40579 9640 40588
rect 9588 40545 9597 40579
rect 9597 40545 9631 40579
rect 9631 40545 9640 40579
rect 9588 40536 9640 40545
rect 9772 40536 9824 40588
rect 12532 40604 12584 40656
rect 11428 40579 11480 40588
rect 11428 40545 11437 40579
rect 11437 40545 11471 40579
rect 11471 40545 11480 40579
rect 11428 40536 11480 40545
rect 8760 40468 8812 40520
rect 11336 40468 11388 40520
rect 11704 40468 11756 40520
rect 7656 40400 7708 40452
rect 8392 40400 8444 40452
rect 10692 40400 10744 40452
rect 11244 40400 11296 40452
rect 12348 40536 12400 40588
rect 4436 40332 4488 40384
rect 4988 40332 5040 40384
rect 5908 40375 5960 40384
rect 5908 40341 5917 40375
rect 5917 40341 5951 40375
rect 5951 40341 5960 40375
rect 5908 40332 5960 40341
rect 7288 40375 7340 40384
rect 7288 40341 7297 40375
rect 7297 40341 7331 40375
rect 7331 40341 7340 40375
rect 7288 40332 7340 40341
rect 7472 40375 7524 40384
rect 7472 40341 7481 40375
rect 7481 40341 7515 40375
rect 7515 40341 7524 40375
rect 7472 40332 7524 40341
rect 7932 40332 7984 40384
rect 9220 40332 9272 40384
rect 11888 40375 11940 40384
rect 11888 40341 11897 40375
rect 11897 40341 11931 40375
rect 11931 40341 11940 40375
rect 11888 40332 11940 40341
rect 12072 40332 12124 40384
rect 3662 40230 3714 40282
rect 3726 40230 3778 40282
rect 3790 40230 3842 40282
rect 3854 40230 3906 40282
rect 3918 40230 3970 40282
rect 10062 40230 10114 40282
rect 10126 40230 10178 40282
rect 10190 40230 10242 40282
rect 10254 40230 10306 40282
rect 10318 40230 10370 40282
rect 1768 40128 1820 40180
rect 2136 40171 2188 40180
rect 2136 40137 2145 40171
rect 2145 40137 2179 40171
rect 2179 40137 2188 40171
rect 2136 40128 2188 40137
rect 2412 40128 2464 40180
rect 2504 40171 2556 40180
rect 2504 40137 2513 40171
rect 2513 40137 2547 40171
rect 2547 40137 2556 40171
rect 2504 40128 2556 40137
rect 3056 40128 3108 40180
rect 3700 40128 3752 40180
rect 6644 40128 6696 40180
rect 7656 40128 7708 40180
rect 8208 40128 8260 40180
rect 9128 40171 9180 40180
rect 9128 40137 9137 40171
rect 9137 40137 9171 40171
rect 9171 40137 9180 40171
rect 9128 40128 9180 40137
rect 10508 40128 10560 40180
rect 10692 40128 10744 40180
rect 2044 40060 2096 40112
rect 1032 39924 1084 39976
rect 1216 39967 1268 39976
rect 1216 39933 1225 39967
rect 1225 39933 1259 39967
rect 1259 39933 1268 39967
rect 1216 39924 1268 39933
rect 1952 39992 2004 40044
rect 940 39831 992 39840
rect 940 39797 949 39831
rect 949 39797 983 39831
rect 983 39797 992 39831
rect 940 39788 992 39797
rect 1124 39788 1176 39840
rect 1492 39788 1544 39840
rect 2412 39992 2464 40044
rect 4160 40060 4212 40112
rect 4988 40060 5040 40112
rect 7380 40060 7432 40112
rect 11060 40060 11112 40112
rect 2688 39967 2740 39976
rect 2688 39933 2697 39967
rect 2697 39933 2740 39967
rect 2688 39924 2740 39933
rect 2964 39967 3016 39976
rect 2964 39933 2973 39967
rect 2973 39933 3007 39967
rect 3007 39933 3016 39967
rect 2964 39924 3016 39933
rect 4160 39924 4212 39976
rect 4528 39992 4580 40044
rect 4344 39967 4396 39976
rect 4344 39933 4353 39967
rect 4353 39933 4387 39967
rect 4387 39933 4396 39967
rect 4344 39924 4396 39933
rect 4436 39967 4488 39976
rect 4436 39933 4446 39967
rect 4446 39933 4480 39967
rect 4480 39933 4488 39967
rect 4436 39924 4488 39933
rect 4620 39967 4672 39976
rect 4620 39933 4629 39967
rect 4629 39933 4663 39967
rect 4663 39933 4672 39967
rect 4620 39924 4672 39933
rect 4896 39924 4948 39976
rect 5080 40035 5132 40044
rect 5080 40001 5089 40035
rect 5089 40001 5123 40035
rect 5123 40001 5132 40035
rect 5080 39992 5132 40001
rect 7288 39992 7340 40044
rect 10416 39992 10468 40044
rect 2044 39856 2096 39908
rect 3148 39856 3200 39908
rect 2964 39788 3016 39840
rect 3700 39899 3752 39908
rect 3700 39865 3709 39899
rect 3709 39865 3743 39899
rect 3743 39865 3752 39899
rect 3700 39856 3752 39865
rect 4528 39788 4580 39840
rect 5908 39924 5960 39976
rect 7012 39924 7064 39976
rect 7472 39924 7524 39976
rect 7564 39967 7616 39976
rect 7564 39933 7573 39967
rect 7573 39933 7607 39967
rect 7607 39933 7616 39967
rect 7564 39924 7616 39933
rect 4804 39788 4856 39840
rect 4988 39831 5040 39840
rect 4988 39797 4997 39831
rect 4997 39797 5031 39831
rect 5031 39797 5040 39831
rect 4988 39788 5040 39797
rect 6184 39856 6236 39908
rect 5356 39788 5408 39840
rect 6368 39788 6420 39840
rect 7196 39788 7248 39840
rect 7656 39788 7708 39840
rect 7748 39788 7800 39840
rect 8668 39967 8720 39976
rect 8668 39933 8677 39967
rect 8677 39933 8711 39967
rect 8711 39933 8720 39967
rect 8668 39924 8720 39933
rect 8944 39924 8996 39976
rect 9220 39967 9272 39976
rect 9220 39933 9229 39967
rect 9229 39933 9263 39967
rect 9263 39933 9272 39967
rect 9220 39924 9272 39933
rect 9680 39924 9732 39976
rect 9312 39856 9364 39908
rect 10140 39899 10192 39908
rect 10140 39865 10149 39899
rect 10149 39865 10183 39899
rect 10183 39865 10192 39899
rect 10140 39856 10192 39865
rect 10232 39856 10284 39908
rect 9680 39831 9732 39840
rect 9680 39797 9705 39831
rect 9705 39797 9732 39831
rect 9680 39788 9732 39797
rect 9864 39831 9916 39840
rect 9864 39797 9873 39831
rect 9873 39797 9907 39831
rect 9907 39797 9916 39831
rect 9864 39788 9916 39797
rect 10048 39831 10100 39840
rect 10048 39797 10057 39831
rect 10057 39797 10091 39831
rect 10091 39797 10100 39831
rect 10048 39788 10100 39797
rect 11244 39992 11296 40044
rect 12256 40035 12308 40044
rect 12256 40001 12265 40035
rect 12265 40001 12299 40035
rect 12299 40001 12308 40035
rect 12256 39992 12308 40001
rect 11060 39856 11112 39908
rect 11612 39856 11664 39908
rect 11888 39856 11940 39908
rect 10876 39831 10928 39840
rect 10876 39797 10885 39831
rect 10885 39797 10919 39831
rect 10919 39797 10928 39831
rect 10876 39788 10928 39797
rect 11244 39788 11296 39840
rect 12072 39788 12124 39840
rect 4322 39686 4374 39738
rect 4386 39686 4438 39738
rect 4450 39686 4502 39738
rect 4514 39686 4566 39738
rect 4578 39686 4630 39738
rect 10722 39686 10774 39738
rect 10786 39686 10838 39738
rect 10850 39686 10902 39738
rect 10914 39686 10966 39738
rect 10978 39686 11030 39738
rect 2780 39584 2832 39636
rect 4712 39584 4764 39636
rect 4988 39584 5040 39636
rect 1492 39448 1544 39500
rect 1860 39491 1912 39500
rect 1860 39457 1869 39491
rect 1869 39457 1903 39491
rect 1903 39457 1912 39491
rect 1860 39448 1912 39457
rect 2412 39516 2464 39568
rect 2320 39491 2372 39500
rect 2320 39457 2329 39491
rect 2329 39457 2363 39491
rect 2363 39457 2372 39491
rect 2320 39448 2372 39457
rect 5080 39516 5132 39568
rect 664 39380 716 39432
rect 1400 39355 1452 39364
rect 1400 39321 1409 39355
rect 1409 39321 1443 39355
rect 1443 39321 1452 39355
rect 1400 39312 1452 39321
rect 1768 39380 1820 39432
rect 3056 39448 3108 39500
rect 4252 39448 4304 39500
rect 4712 39448 4764 39500
rect 6184 39448 6236 39500
rect 7748 39448 7800 39500
rect 3424 39380 3476 39432
rect 5908 39423 5960 39432
rect 5908 39389 5917 39423
rect 5917 39389 5951 39423
rect 5951 39389 5960 39423
rect 5908 39380 5960 39389
rect 7564 39380 7616 39432
rect 7840 39423 7892 39432
rect 7840 39389 7849 39423
rect 7849 39389 7883 39423
rect 7883 39389 7892 39423
rect 7840 39380 7892 39389
rect 8852 39448 8904 39500
rect 10232 39584 10284 39636
rect 11152 39584 11204 39636
rect 9864 39516 9916 39568
rect 4068 39312 4120 39364
rect 8576 39312 8628 39364
rect 940 39287 992 39296
rect 940 39253 949 39287
rect 949 39253 983 39287
rect 983 39253 992 39287
rect 940 39244 992 39253
rect 1952 39244 2004 39296
rect 3056 39244 3108 39296
rect 4252 39244 4304 39296
rect 6644 39244 6696 39296
rect 7196 39244 7248 39296
rect 7748 39244 7800 39296
rect 8208 39244 8260 39296
rect 8944 39244 8996 39296
rect 9404 39448 9456 39500
rect 9956 39448 10008 39500
rect 10324 39448 10376 39500
rect 12072 39516 12124 39568
rect 10692 39355 10744 39364
rect 10692 39321 10701 39355
rect 10701 39321 10735 39355
rect 10735 39321 10744 39355
rect 10692 39312 10744 39321
rect 11244 39312 11296 39364
rect 11428 39312 11480 39364
rect 11612 39380 11664 39432
rect 11796 39312 11848 39364
rect 12440 39312 12492 39364
rect 10968 39287 11020 39296
rect 10968 39253 10977 39287
rect 10977 39253 11011 39287
rect 11011 39253 11020 39287
rect 10968 39244 11020 39253
rect 12348 39244 12400 39296
rect 3662 39142 3714 39194
rect 3726 39142 3778 39194
rect 3790 39142 3842 39194
rect 3854 39142 3906 39194
rect 3918 39142 3970 39194
rect 10062 39142 10114 39194
rect 10126 39142 10178 39194
rect 10190 39142 10242 39194
rect 10254 39142 10306 39194
rect 10318 39142 10370 39194
rect 3332 39040 3384 39092
rect 3516 39040 3568 39092
rect 940 38972 992 39024
rect 480 38836 532 38888
rect 3884 39015 3936 39024
rect 3884 38981 3893 39015
rect 3893 38981 3927 39015
rect 3927 38981 3936 39015
rect 3884 38972 3936 38981
rect 7196 39015 7248 39024
rect 7196 38981 7205 39015
rect 7205 38981 7239 39015
rect 7239 38981 7248 39015
rect 7196 38972 7248 38981
rect 7380 38972 7432 39024
rect 9864 39040 9916 39092
rect 9956 39083 10008 39092
rect 9956 39049 9965 39083
rect 9965 39049 9999 39083
rect 9999 39049 10008 39083
rect 9956 39040 10008 39049
rect 10968 39040 11020 39092
rect 8300 38972 8352 39024
rect 9588 39015 9640 39024
rect 9588 38981 9597 39015
rect 9597 38981 9631 39015
rect 9631 38981 9640 39015
rect 9588 38972 9640 38981
rect 10048 38972 10100 39024
rect 10600 38972 10652 39024
rect 1400 38879 1452 38888
rect 1400 38845 1409 38879
rect 1409 38845 1443 38879
rect 1443 38845 1452 38879
rect 1400 38836 1452 38845
rect 2688 38904 2740 38956
rect 1952 38811 2004 38820
rect 1952 38777 1986 38811
rect 1986 38777 2004 38811
rect 1952 38768 2004 38777
rect 2780 38836 2832 38888
rect 2136 38768 2188 38820
rect 480 38700 532 38752
rect 1124 38700 1176 38752
rect 3516 38743 3568 38752
rect 3516 38709 3525 38743
rect 3525 38709 3559 38743
rect 3559 38709 3568 38743
rect 3516 38700 3568 38709
rect 4160 38904 4212 38956
rect 5080 38904 5132 38956
rect 5816 38879 5868 38888
rect 5816 38845 5825 38879
rect 5825 38845 5859 38879
rect 5859 38845 5868 38879
rect 5816 38836 5868 38845
rect 7656 38904 7708 38956
rect 8668 38947 8720 38956
rect 8668 38913 8677 38947
rect 8677 38913 8711 38947
rect 8711 38913 8720 38947
rect 8668 38904 8720 38913
rect 9496 38904 9548 38956
rect 7748 38836 7800 38888
rect 8024 38836 8076 38888
rect 8760 38836 8812 38888
rect 4160 38811 4212 38820
rect 4160 38777 4169 38811
rect 4169 38777 4203 38811
rect 4203 38777 4212 38811
rect 4160 38768 4212 38777
rect 6092 38811 6144 38820
rect 6092 38777 6126 38811
rect 6126 38777 6144 38811
rect 5080 38700 5132 38752
rect 6092 38768 6144 38777
rect 7564 38768 7616 38820
rect 9772 38836 9824 38888
rect 10324 38836 10376 38888
rect 9036 38811 9088 38820
rect 9036 38777 9045 38811
rect 9045 38777 9079 38811
rect 9079 38777 9088 38811
rect 9036 38768 9088 38777
rect 11888 38768 11940 38820
rect 7196 38700 7248 38752
rect 7380 38700 7432 38752
rect 7656 38700 7708 38752
rect 7748 38700 7800 38752
rect 8024 38700 8076 38752
rect 8944 38700 8996 38752
rect 9312 38743 9364 38752
rect 9312 38709 9321 38743
rect 9321 38709 9355 38743
rect 9355 38709 9364 38743
rect 9312 38700 9364 38709
rect 9404 38700 9456 38752
rect 10140 38743 10192 38752
rect 10140 38709 10149 38743
rect 10149 38709 10183 38743
rect 10183 38709 10192 38743
rect 10140 38700 10192 38709
rect 10416 38700 10468 38752
rect 11980 38700 12032 38752
rect 12256 38700 12308 38752
rect 4322 38598 4374 38650
rect 4386 38598 4438 38650
rect 4450 38598 4502 38650
rect 4514 38598 4566 38650
rect 4578 38598 4630 38650
rect 10722 38598 10774 38650
rect 10786 38598 10838 38650
rect 10850 38598 10902 38650
rect 10914 38598 10966 38650
rect 10978 38598 11030 38650
rect 1400 38496 1452 38548
rect 2228 38496 2280 38548
rect 2320 38496 2372 38548
rect 296 38428 348 38480
rect 1676 38428 1728 38480
rect 1492 38360 1544 38412
rect 1952 38360 2004 38412
rect 4160 38496 4212 38548
rect 4344 38496 4396 38548
rect 4896 38496 4948 38548
rect 5264 38496 5316 38548
rect 2136 38360 2188 38412
rect 940 38335 992 38344
rect 940 38301 949 38335
rect 949 38301 983 38335
rect 983 38301 992 38335
rect 940 38292 992 38301
rect 3700 38403 3752 38412
rect 3700 38369 3709 38403
rect 3709 38369 3743 38403
rect 3743 38369 3752 38403
rect 3700 38360 3752 38369
rect 3792 38403 3844 38412
rect 3792 38369 3801 38403
rect 3801 38369 3835 38403
rect 3835 38369 3844 38403
rect 3792 38360 3844 38369
rect 4068 38403 4120 38412
rect 4068 38369 4102 38403
rect 4102 38369 4120 38403
rect 4068 38360 4120 38369
rect 4436 38360 4488 38412
rect 5356 38428 5408 38480
rect 6460 38428 6512 38480
rect 9036 38496 9088 38548
rect 9312 38496 9364 38548
rect 10232 38496 10284 38548
rect 10508 38496 10560 38548
rect 10416 38471 10468 38480
rect 4804 38292 4856 38344
rect 3424 38267 3476 38276
rect 3424 38233 3433 38267
rect 3433 38233 3467 38267
rect 3467 38233 3476 38267
rect 3424 38224 3476 38233
rect 5540 38403 5592 38412
rect 5540 38369 5549 38403
rect 5549 38369 5583 38403
rect 5583 38369 5592 38403
rect 5540 38360 5592 38369
rect 5816 38403 5868 38412
rect 5816 38369 5825 38403
rect 5825 38369 5859 38403
rect 5859 38369 5868 38403
rect 5816 38360 5868 38369
rect 7932 38360 7984 38412
rect 9036 38403 9088 38412
rect 5632 38292 5684 38344
rect 7104 38292 7156 38344
rect 7840 38292 7892 38344
rect 8300 38292 8352 38344
rect 9036 38369 9045 38403
rect 9045 38369 9079 38403
rect 9079 38369 9088 38403
rect 9036 38360 9088 38369
rect 8668 38292 8720 38344
rect 9588 38403 9640 38412
rect 9588 38369 9597 38403
rect 9597 38369 9631 38403
rect 9631 38369 9640 38403
rect 9588 38360 9640 38369
rect 9772 38403 9824 38412
rect 9772 38369 9781 38403
rect 9781 38369 9815 38403
rect 9815 38369 9824 38403
rect 9772 38360 9824 38369
rect 9864 38360 9916 38412
rect 10048 38360 10100 38412
rect 10416 38437 10425 38471
rect 10425 38437 10459 38471
rect 10459 38437 10468 38471
rect 10416 38428 10468 38437
rect 10600 38471 10652 38480
rect 10600 38437 10625 38471
rect 10625 38437 10652 38471
rect 10600 38428 10652 38437
rect 10968 38471 11020 38480
rect 10968 38437 10977 38471
rect 10977 38437 11011 38471
rect 11011 38437 11020 38471
rect 10968 38428 11020 38437
rect 11152 38496 11204 38548
rect 11704 38496 11756 38548
rect 11244 38403 11296 38412
rect 11244 38369 11253 38403
rect 11253 38369 11287 38403
rect 11287 38369 11296 38403
rect 11244 38360 11296 38369
rect 5816 38224 5868 38276
rect 7748 38224 7800 38276
rect 8576 38224 8628 38276
rect 3240 38156 3292 38208
rect 7104 38156 7156 38208
rect 7656 38156 7708 38208
rect 8668 38199 8720 38208
rect 8668 38165 8677 38199
rect 8677 38165 8711 38199
rect 8711 38165 8720 38199
rect 8668 38156 8720 38165
rect 8760 38156 8812 38208
rect 9404 38156 9456 38208
rect 10508 38156 10560 38208
rect 11428 38292 11480 38344
rect 12072 38403 12124 38412
rect 12072 38369 12081 38403
rect 12081 38369 12115 38403
rect 12115 38369 12124 38403
rect 12072 38360 12124 38369
rect 12716 38292 12768 38344
rect 10692 38224 10744 38276
rect 10784 38199 10836 38208
rect 10784 38165 10793 38199
rect 10793 38165 10827 38199
rect 10827 38165 10836 38199
rect 10784 38156 10836 38165
rect 11152 38224 11204 38276
rect 11796 38224 11848 38276
rect 3662 38054 3714 38106
rect 3726 38054 3778 38106
rect 3790 38054 3842 38106
rect 3854 38054 3906 38106
rect 3918 38054 3970 38106
rect 10062 38054 10114 38106
rect 10126 38054 10178 38106
rect 10190 38054 10242 38106
rect 10254 38054 10306 38106
rect 10318 38054 10370 38106
rect 1032 37952 1084 38004
rect 2044 37952 2096 38004
rect 3976 37952 4028 38004
rect 4712 37952 4764 38004
rect 5264 37952 5316 38004
rect 5356 37952 5408 38004
rect 6828 37952 6880 38004
rect 7104 37952 7156 38004
rect 2872 37884 2924 37936
rect 2596 37859 2648 37868
rect 2596 37825 2605 37859
rect 2605 37825 2639 37859
rect 2639 37825 2648 37859
rect 2596 37816 2648 37825
rect 3332 37816 3384 37868
rect 4528 37884 4580 37936
rect 5448 37884 5500 37936
rect 6092 37884 6144 37936
rect 11244 37952 11296 38004
rect 11796 37952 11848 38004
rect 12624 37884 12676 37936
rect 1584 37748 1636 37800
rect 2504 37748 2556 37800
rect 1124 37723 1176 37732
rect 1124 37689 1158 37723
rect 1158 37689 1176 37723
rect 1124 37680 1176 37689
rect 1676 37680 1728 37732
rect 3792 37748 3844 37800
rect 3976 37748 4028 37800
rect 4252 37791 4304 37800
rect 4252 37757 4262 37791
rect 4262 37757 4296 37791
rect 4296 37757 4304 37791
rect 4252 37748 4304 37757
rect 4804 37748 4856 37800
rect 5356 37748 5408 37800
rect 6644 37748 6696 37800
rect 6920 37748 6972 37800
rect 3056 37680 3108 37732
rect 1216 37612 1268 37664
rect 1860 37612 1912 37664
rect 2228 37655 2280 37664
rect 2228 37621 2237 37655
rect 2237 37621 2271 37655
rect 2271 37621 2280 37655
rect 2228 37612 2280 37621
rect 2872 37612 2924 37664
rect 3516 37612 3568 37664
rect 3700 37655 3752 37664
rect 3700 37621 3709 37655
rect 3709 37621 3743 37655
rect 3743 37621 3752 37655
rect 3700 37612 3752 37621
rect 4436 37723 4488 37732
rect 4436 37689 4445 37723
rect 4445 37689 4479 37723
rect 4479 37689 4488 37723
rect 4436 37680 4488 37689
rect 4528 37723 4580 37732
rect 4528 37689 4537 37723
rect 4537 37689 4571 37723
rect 4571 37689 4580 37723
rect 4528 37680 4580 37689
rect 5540 37680 5592 37732
rect 7104 37680 7156 37732
rect 7196 37680 7248 37732
rect 4620 37612 4672 37664
rect 5724 37612 5776 37664
rect 5908 37612 5960 37664
rect 7840 37655 7892 37664
rect 7840 37621 7849 37655
rect 7849 37621 7883 37655
rect 7883 37621 7892 37655
rect 7840 37612 7892 37621
rect 8208 37791 8260 37800
rect 8208 37757 8217 37791
rect 8217 37757 8251 37791
rect 8251 37757 8260 37791
rect 8208 37748 8260 37757
rect 8484 37748 8536 37800
rect 8576 37791 8628 37800
rect 8576 37757 8585 37791
rect 8585 37757 8619 37791
rect 8619 37757 8628 37791
rect 8576 37748 8628 37757
rect 8668 37748 8720 37800
rect 8944 37748 8996 37800
rect 10784 37816 10836 37868
rect 9220 37748 9272 37800
rect 9588 37791 9640 37800
rect 9588 37757 9597 37791
rect 9597 37757 9631 37791
rect 9631 37757 9640 37791
rect 9588 37748 9640 37757
rect 11796 37791 11848 37800
rect 11796 37757 11805 37791
rect 11805 37757 11839 37791
rect 11839 37757 11848 37791
rect 11796 37748 11848 37757
rect 9312 37680 9364 37732
rect 12072 37748 12124 37800
rect 9220 37612 9272 37664
rect 10416 37612 10468 37664
rect 4322 37510 4374 37562
rect 4386 37510 4438 37562
rect 4450 37510 4502 37562
rect 4514 37510 4566 37562
rect 4578 37510 4630 37562
rect 10722 37510 10774 37562
rect 10786 37510 10838 37562
rect 10850 37510 10902 37562
rect 10914 37510 10966 37562
rect 10978 37510 11030 37562
rect 848 37408 900 37460
rect 1032 37315 1084 37324
rect 1032 37281 1041 37315
rect 1041 37281 1075 37315
rect 1075 37281 1084 37315
rect 1032 37272 1084 37281
rect 5908 37408 5960 37460
rect 1492 37340 1544 37392
rect 1216 37315 1268 37324
rect 1216 37281 1225 37315
rect 1225 37281 1259 37315
rect 1259 37281 1268 37315
rect 1216 37272 1268 37281
rect 1400 37315 1452 37324
rect 1400 37281 1409 37315
rect 1409 37281 1443 37315
rect 1443 37281 1452 37315
rect 1400 37272 1452 37281
rect 1584 37272 1636 37324
rect 1768 37272 1820 37324
rect 2228 37272 2280 37324
rect 3608 37315 3660 37324
rect 3608 37281 3617 37315
rect 3617 37281 3651 37315
rect 3651 37281 3660 37315
rect 3608 37272 3660 37281
rect 3792 37315 3844 37324
rect 3792 37281 3801 37315
rect 3801 37281 3835 37315
rect 3835 37281 3844 37315
rect 3792 37272 3844 37281
rect 1676 37136 1728 37188
rect 2688 37136 2740 37188
rect 4160 37204 4212 37256
rect 5080 37315 5132 37324
rect 5080 37281 5089 37315
rect 5089 37281 5123 37315
rect 5123 37281 5132 37315
rect 5080 37272 5132 37281
rect 6828 37340 6880 37392
rect 5540 37315 5592 37324
rect 5540 37281 5549 37315
rect 5549 37281 5583 37315
rect 5583 37281 5592 37315
rect 5540 37272 5592 37281
rect 6460 37315 6512 37324
rect 6460 37281 6469 37315
rect 6469 37281 6503 37315
rect 6503 37281 6512 37315
rect 6460 37272 6512 37281
rect 6552 37272 6604 37324
rect 6920 37315 6972 37324
rect 6920 37281 6929 37315
rect 6929 37281 6963 37315
rect 6963 37281 6972 37315
rect 6920 37272 6972 37281
rect 4436 37136 4488 37188
rect 4804 37204 4856 37256
rect 7196 37451 7248 37460
rect 7196 37417 7205 37451
rect 7205 37417 7239 37451
rect 7239 37417 7248 37451
rect 7196 37408 7248 37417
rect 7840 37408 7892 37460
rect 8852 37451 8904 37460
rect 8852 37417 8861 37451
rect 8861 37417 8895 37451
rect 8895 37417 8904 37451
rect 8852 37408 8904 37417
rect 9588 37408 9640 37460
rect 10876 37408 10928 37460
rect 11152 37408 11204 37460
rect 7656 37383 7708 37392
rect 7656 37349 7665 37383
rect 7665 37349 7699 37383
rect 7699 37349 7708 37383
rect 7656 37340 7708 37349
rect 8116 37204 8168 37256
rect 8300 37315 8352 37324
rect 8300 37281 8309 37315
rect 8309 37281 8343 37315
rect 8343 37281 8352 37315
rect 8300 37272 8352 37281
rect 9680 37340 9732 37392
rect 11244 37340 11296 37392
rect 11796 37340 11848 37392
rect 8760 37315 8812 37324
rect 8760 37281 8769 37315
rect 8769 37281 8803 37315
rect 8803 37281 8812 37315
rect 8760 37272 8812 37281
rect 8852 37272 8904 37324
rect 9588 37272 9640 37324
rect 10324 37272 10376 37324
rect 3056 37111 3108 37120
rect 3056 37077 3065 37111
rect 3065 37077 3099 37111
rect 3099 37077 3108 37111
rect 3056 37068 3108 37077
rect 3332 37068 3384 37120
rect 5540 37136 5592 37188
rect 7288 37136 7340 37188
rect 7656 37136 7708 37188
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 8392 37136 8444 37188
rect 9036 37136 9088 37188
rect 11244 37247 11296 37256
rect 11244 37213 11253 37247
rect 11253 37213 11287 37247
rect 11287 37213 11296 37247
rect 11244 37204 11296 37213
rect 11428 37204 11480 37256
rect 11704 37315 11756 37324
rect 11704 37281 11713 37315
rect 11713 37281 11747 37315
rect 11747 37281 11756 37315
rect 11704 37272 11756 37281
rect 11980 37315 12032 37324
rect 11980 37281 11989 37315
rect 11989 37281 12023 37315
rect 12023 37281 12032 37315
rect 11980 37272 12032 37281
rect 12532 37204 12584 37256
rect 11704 37136 11756 37188
rect 8576 37068 8628 37120
rect 9128 37068 9180 37120
rect 9404 37068 9456 37120
rect 9772 37068 9824 37120
rect 11152 37111 11204 37120
rect 11152 37077 11161 37111
rect 11161 37077 11195 37111
rect 11195 37077 11204 37111
rect 11152 37068 11204 37077
rect 12716 37068 12768 37120
rect 3662 36966 3714 37018
rect 3726 36966 3778 37018
rect 3790 36966 3842 37018
rect 3854 36966 3906 37018
rect 3918 36966 3970 37018
rect 10062 36966 10114 37018
rect 10126 36966 10178 37018
rect 10190 36966 10242 37018
rect 10254 36966 10306 37018
rect 10318 36966 10370 37018
rect 1400 36864 1452 36916
rect 3148 36864 3200 36916
rect 3240 36907 3292 36916
rect 3240 36873 3249 36907
rect 3249 36873 3283 36907
rect 3283 36873 3292 36907
rect 3240 36864 3292 36873
rect 3884 36864 3936 36916
rect 3056 36796 3108 36848
rect 3516 36796 3568 36848
rect 1584 36728 1636 36780
rect 2780 36728 2832 36780
rect 3148 36728 3200 36780
rect 204 36660 256 36712
rect 1124 36660 1176 36712
rect 1768 36660 1820 36712
rect 7656 36864 7708 36916
rect 8300 36864 8352 36916
rect 8576 36864 8628 36916
rect 8668 36864 8720 36916
rect 8760 36907 8812 36916
rect 8760 36873 8769 36907
rect 8769 36873 8803 36907
rect 8803 36873 8812 36907
rect 8760 36864 8812 36873
rect 9220 36864 9272 36916
rect 4896 36796 4948 36848
rect 6736 36796 6788 36848
rect 7104 36796 7156 36848
rect 8392 36796 8444 36848
rect 5448 36728 5500 36780
rect 6092 36728 6144 36780
rect 6552 36728 6604 36780
rect 4988 36660 5040 36712
rect 3056 36635 3108 36644
rect 3056 36601 3065 36635
rect 3065 36601 3099 36635
rect 3099 36601 3108 36635
rect 3056 36592 3108 36601
rect 4252 36592 4304 36644
rect 4344 36635 4396 36644
rect 4344 36601 4384 36635
rect 4384 36601 4396 36635
rect 4344 36592 4396 36601
rect 5080 36592 5132 36644
rect 5632 36592 5684 36644
rect 7012 36660 7064 36712
rect 7288 36703 7340 36712
rect 7288 36669 7297 36703
rect 7297 36669 7331 36703
rect 7331 36669 7340 36703
rect 7288 36660 7340 36669
rect 7472 36703 7524 36712
rect 7472 36669 7481 36703
rect 7481 36669 7515 36703
rect 7515 36669 7524 36703
rect 7472 36660 7524 36669
rect 7748 36660 7800 36712
rect 7840 36660 7892 36712
rect 8760 36728 8812 36780
rect 7104 36592 7156 36644
rect 8392 36592 8444 36644
rect 388 36524 440 36576
rect 3792 36524 3844 36576
rect 4528 36524 4580 36576
rect 4712 36524 4764 36576
rect 5908 36567 5960 36576
rect 5908 36533 5917 36567
rect 5917 36533 5951 36567
rect 5951 36533 5960 36567
rect 5908 36524 5960 36533
rect 6276 36524 6328 36576
rect 6736 36567 6788 36576
rect 6736 36533 6745 36567
rect 6745 36533 6779 36567
rect 6779 36533 6788 36567
rect 6736 36524 6788 36533
rect 7288 36524 7340 36576
rect 7656 36567 7708 36576
rect 7656 36533 7665 36567
rect 7665 36533 7699 36567
rect 7699 36533 7708 36567
rect 7656 36524 7708 36533
rect 7748 36524 7800 36576
rect 8664 36635 8716 36678
rect 8664 36626 8677 36635
rect 8677 36626 8711 36635
rect 8711 36626 8716 36635
rect 8944 36796 8996 36848
rect 9128 36796 9180 36848
rect 9036 36771 9088 36780
rect 9036 36737 9045 36771
rect 9045 36737 9079 36771
rect 9079 36737 9088 36771
rect 9036 36728 9088 36737
rect 11244 36864 11296 36916
rect 11796 36864 11848 36916
rect 9680 36796 9732 36848
rect 10324 36771 10376 36780
rect 10324 36737 10333 36771
rect 10333 36737 10367 36771
rect 10367 36737 10376 36771
rect 10324 36728 10376 36737
rect 10600 36728 10652 36780
rect 10876 36771 10928 36780
rect 10876 36737 10885 36771
rect 10885 36737 10919 36771
rect 10919 36737 10928 36771
rect 10876 36728 10928 36737
rect 9036 36592 9088 36644
rect 9404 36703 9456 36712
rect 9404 36669 9413 36703
rect 9413 36669 9447 36703
rect 9447 36669 9456 36703
rect 9404 36660 9456 36669
rect 10416 36660 10468 36712
rect 11980 36660 12032 36712
rect 9404 36524 9456 36576
rect 9496 36524 9548 36576
rect 9772 36567 9824 36576
rect 9772 36533 9781 36567
rect 9781 36533 9815 36567
rect 9815 36533 9824 36567
rect 9772 36524 9824 36533
rect 9864 36524 9916 36576
rect 9956 36524 10008 36576
rect 10416 36524 10468 36576
rect 11152 36635 11204 36644
rect 11152 36601 11186 36635
rect 11186 36601 11204 36635
rect 11152 36592 11204 36601
rect 11244 36524 11296 36576
rect 12072 36524 12124 36576
rect 4322 36422 4374 36474
rect 4386 36422 4438 36474
rect 4450 36422 4502 36474
rect 4514 36422 4566 36474
rect 4578 36422 4630 36474
rect 10722 36422 10774 36474
rect 10786 36422 10838 36474
rect 10850 36422 10902 36474
rect 10914 36422 10966 36474
rect 10978 36422 11030 36474
rect 3516 36320 3568 36372
rect 4804 36320 4856 36372
rect 6276 36363 6328 36372
rect 6276 36329 6285 36363
rect 6285 36329 6319 36363
rect 6319 36329 6328 36363
rect 6276 36320 6328 36329
rect 6644 36320 6696 36372
rect 5908 36252 5960 36304
rect 6736 36252 6788 36304
rect 112 36184 164 36236
rect 296 36184 348 36236
rect 1032 36184 1084 36236
rect 1492 36184 1544 36236
rect 1584 36227 1636 36236
rect 1584 36193 1593 36227
rect 1593 36193 1627 36227
rect 1627 36193 1636 36227
rect 1584 36184 1636 36193
rect 3516 36184 3568 36236
rect 4160 36184 4212 36236
rect 4252 36227 4304 36236
rect 4252 36193 4261 36227
rect 4261 36193 4295 36227
rect 4295 36193 4304 36227
rect 4252 36184 4304 36193
rect 4344 36184 4396 36236
rect 5632 36184 5684 36236
rect 6552 36184 6604 36236
rect 6644 36227 6696 36236
rect 6644 36193 6653 36227
rect 6653 36193 6687 36227
rect 6687 36193 6696 36227
rect 6644 36184 6696 36193
rect 7012 36252 7064 36304
rect 8024 36252 8076 36304
rect 8208 36252 8260 36304
rect 756 36116 808 36168
rect 3976 36116 4028 36168
rect 6368 36159 6420 36168
rect 6368 36125 6377 36159
rect 6377 36125 6411 36159
rect 6411 36125 6420 36159
rect 6368 36116 6420 36125
rect 6460 36116 6512 36168
rect 1952 36048 2004 36100
rect 3792 36048 3844 36100
rect 4160 36048 4212 36100
rect 5816 36048 5868 36100
rect 7380 36184 7432 36236
rect 7012 36116 7064 36168
rect 7840 36184 7892 36236
rect 7932 36116 7984 36168
rect 7840 36048 7892 36100
rect 8208 36048 8260 36100
rect 8760 36252 8812 36304
rect 8944 36252 8996 36304
rect 10324 36320 10376 36372
rect 10416 36320 10468 36372
rect 10692 36320 10744 36372
rect 11152 36320 11204 36372
rect 12164 36320 12216 36372
rect 9404 36184 9456 36236
rect 10232 36252 10284 36304
rect 10140 36184 10192 36236
rect 10416 36227 10468 36236
rect 10416 36193 10425 36227
rect 10425 36193 10459 36227
rect 10459 36193 10468 36227
rect 10416 36184 10468 36193
rect 8576 36116 8628 36168
rect 9312 36116 9364 36168
rect 9680 36159 9732 36168
rect 9680 36125 9689 36159
rect 9689 36125 9723 36159
rect 9723 36125 9732 36159
rect 9680 36116 9732 36125
rect 10048 36116 10100 36168
rect 10140 36048 10192 36100
rect 10968 36116 11020 36168
rect 11152 36048 11204 36100
rect 940 36023 992 36032
rect 940 35989 949 36023
rect 949 35989 983 36023
rect 983 35989 992 36023
rect 940 35980 992 35989
rect 3424 35980 3476 36032
rect 3884 35980 3936 36032
rect 5448 35980 5500 36032
rect 6460 35980 6512 36032
rect 7380 35980 7432 36032
rect 8116 35980 8168 36032
rect 8392 36023 8444 36032
rect 8392 35989 8401 36023
rect 8401 35989 8435 36023
rect 8435 35989 8444 36023
rect 8392 35980 8444 35989
rect 8484 35980 8536 36032
rect 8852 36023 8904 36032
rect 8852 35989 8861 36023
rect 8861 35989 8895 36023
rect 8895 35989 8904 36023
rect 8852 35980 8904 35989
rect 9128 35980 9180 36032
rect 10324 35980 10376 36032
rect 10508 35980 10560 36032
rect 11888 36227 11940 36236
rect 11888 36193 11897 36227
rect 11897 36193 11931 36227
rect 11931 36193 11940 36227
rect 11888 36184 11940 36193
rect 11980 36227 12032 36236
rect 11980 36193 11989 36227
rect 11989 36193 12023 36227
rect 12023 36193 12032 36227
rect 11980 36184 12032 36193
rect 12072 36116 12124 36168
rect 11704 36048 11756 36100
rect 12716 36048 12768 36100
rect 12164 35980 12216 36032
rect 12624 35980 12676 36032
rect 3662 35878 3714 35930
rect 3726 35878 3778 35930
rect 3790 35878 3842 35930
rect 3854 35878 3906 35930
rect 3918 35878 3970 35930
rect 10062 35878 10114 35930
rect 10126 35878 10178 35930
rect 10190 35878 10242 35930
rect 10254 35878 10306 35930
rect 10318 35878 10370 35930
rect 1032 35776 1084 35828
rect 1584 35819 1636 35828
rect 1584 35785 1593 35819
rect 1593 35785 1627 35819
rect 1627 35785 1636 35819
rect 1584 35776 1636 35785
rect 2412 35776 2464 35828
rect 2688 35776 2740 35828
rect 6368 35776 6420 35828
rect 6736 35776 6788 35828
rect 7104 35776 7156 35828
rect 8392 35776 8444 35828
rect 9680 35819 9732 35828
rect 9680 35785 9689 35819
rect 9689 35785 9723 35819
rect 9723 35785 9732 35819
rect 9680 35776 9732 35785
rect 9956 35776 10008 35828
rect 10416 35819 10468 35828
rect 10416 35785 10425 35819
rect 10425 35785 10459 35819
rect 10459 35785 10468 35819
rect 10416 35776 10468 35785
rect 3056 35708 3108 35760
rect 3792 35708 3844 35760
rect 4068 35708 4120 35760
rect 1952 35640 2004 35692
rect 2504 35640 2556 35692
rect 2688 35640 2740 35692
rect 3884 35683 3936 35692
rect 3884 35649 3893 35683
rect 3893 35649 3927 35683
rect 3927 35649 3936 35683
rect 3884 35640 3936 35649
rect 3976 35640 4028 35692
rect 6184 35708 6236 35760
rect 1768 35572 1820 35624
rect 2780 35572 2832 35624
rect 3056 35547 3108 35556
rect 3056 35513 3065 35547
rect 3065 35513 3099 35547
rect 3099 35513 3108 35547
rect 3056 35504 3108 35513
rect 5724 35572 5776 35624
rect 6184 35615 6236 35624
rect 6184 35581 6193 35615
rect 6193 35581 6227 35615
rect 6227 35581 6236 35615
rect 6184 35572 6236 35581
rect 6460 35615 6512 35624
rect 6460 35581 6469 35615
rect 6469 35581 6503 35615
rect 6503 35581 6512 35615
rect 6460 35572 6512 35581
rect 6644 35572 6696 35624
rect 7288 35708 7340 35760
rect 7472 35751 7524 35760
rect 7472 35717 7481 35751
rect 7481 35717 7515 35751
rect 7515 35717 7524 35751
rect 7472 35708 7524 35717
rect 9312 35751 9364 35760
rect 9312 35717 9321 35751
rect 9321 35717 9355 35751
rect 9355 35717 9364 35751
rect 9312 35708 9364 35717
rect 7196 35572 7248 35624
rect 8760 35572 8812 35624
rect 9128 35615 9180 35624
rect 9128 35581 9137 35615
rect 9137 35581 9171 35615
rect 9171 35581 9180 35615
rect 9128 35572 9180 35581
rect 11520 35776 11572 35828
rect 11888 35776 11940 35828
rect 10876 35751 10928 35760
rect 10876 35717 10885 35751
rect 10885 35717 10919 35751
rect 10919 35717 10928 35751
rect 10876 35708 10928 35717
rect 9496 35572 9548 35624
rect 9680 35615 9732 35624
rect 9680 35581 9689 35615
rect 9689 35581 9723 35615
rect 9723 35581 9732 35615
rect 9680 35572 9732 35581
rect 3240 35479 3292 35488
rect 3240 35445 3249 35479
rect 3249 35445 3283 35479
rect 3283 35445 3292 35479
rect 3240 35436 3292 35445
rect 3608 35479 3660 35488
rect 3608 35445 3617 35479
rect 3617 35445 3651 35479
rect 3651 35445 3660 35479
rect 3608 35436 3660 35445
rect 4344 35436 4396 35488
rect 4712 35504 4764 35556
rect 4988 35504 5040 35556
rect 5632 35504 5684 35556
rect 6000 35436 6052 35488
rect 6184 35436 6236 35488
rect 7288 35547 7340 35556
rect 7288 35513 7297 35547
rect 7297 35513 7331 35547
rect 7331 35513 7340 35547
rect 7288 35504 7340 35513
rect 8116 35547 8168 35556
rect 8116 35513 8125 35547
rect 8125 35513 8159 35547
rect 8159 35513 8168 35547
rect 8116 35504 8168 35513
rect 8208 35504 8260 35556
rect 8576 35547 8628 35556
rect 8576 35513 8585 35547
rect 8585 35513 8619 35547
rect 8619 35513 8628 35547
rect 8576 35504 8628 35513
rect 8852 35504 8904 35556
rect 10232 35640 10284 35692
rect 10324 35640 10376 35692
rect 9864 35572 9916 35624
rect 10140 35572 10192 35624
rect 10600 35572 10652 35624
rect 10048 35504 10100 35556
rect 10508 35504 10560 35556
rect 8668 35436 8720 35488
rect 9312 35436 9364 35488
rect 10876 35436 10928 35488
rect 11888 35436 11940 35488
rect 12072 35436 12124 35488
rect 4322 35334 4374 35386
rect 4386 35334 4438 35386
rect 4450 35334 4502 35386
rect 4514 35334 4566 35386
rect 4578 35334 4630 35386
rect 10722 35334 10774 35386
rect 10786 35334 10838 35386
rect 10850 35334 10902 35386
rect 10914 35334 10966 35386
rect 10978 35334 11030 35386
rect 664 35232 716 35284
rect 1124 35232 1176 35284
rect 1492 35232 1544 35284
rect 2780 35232 2832 35284
rect 4068 35275 4120 35284
rect 4068 35241 4077 35275
rect 4077 35241 4111 35275
rect 4111 35241 4120 35275
rect 4068 35232 4120 35241
rect 4160 35232 4212 35284
rect 4344 35232 4396 35284
rect 4712 35232 4764 35284
rect 1032 35139 1084 35148
rect 1032 35105 1041 35139
rect 1041 35105 1075 35139
rect 1075 35105 1084 35139
rect 1032 35096 1084 35105
rect 1492 35096 1544 35148
rect 2136 35164 2188 35216
rect 3240 35164 3292 35216
rect 1768 35139 1820 35148
rect 1768 35105 1777 35139
rect 1777 35105 1811 35139
rect 1811 35105 1820 35139
rect 1768 35096 1820 35105
rect 1952 35096 2004 35148
rect 4252 35164 4304 35216
rect 1216 35028 1268 35080
rect 3884 35096 3936 35148
rect 3792 35028 3844 35080
rect 4896 35096 4948 35148
rect 4344 35028 4396 35080
rect 6000 35275 6052 35284
rect 6000 35241 6009 35275
rect 6009 35241 6043 35275
rect 6043 35241 6052 35275
rect 6000 35232 6052 35241
rect 6460 35232 6512 35284
rect 6736 35232 6788 35284
rect 5540 35139 5592 35148
rect 5540 35105 5549 35139
rect 5549 35105 5583 35139
rect 5583 35105 5592 35139
rect 5540 35096 5592 35105
rect 5816 35139 5868 35148
rect 5816 35105 5825 35139
rect 5825 35105 5859 35139
rect 5859 35105 5868 35139
rect 5816 35096 5868 35105
rect 6276 35164 6328 35216
rect 6552 35164 6604 35216
rect 9496 35232 9548 35284
rect 9680 35232 9732 35284
rect 1124 34892 1176 34944
rect 5448 34960 5500 35012
rect 4712 34892 4764 34944
rect 4988 34892 5040 34944
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 5632 35028 5684 35080
rect 6552 35028 6604 35080
rect 6920 35096 6972 35148
rect 7104 35139 7156 35148
rect 7104 35105 7113 35139
rect 7113 35105 7147 35139
rect 7147 35105 7156 35139
rect 7104 35096 7156 35105
rect 7472 35139 7524 35148
rect 7472 35105 7481 35139
rect 7481 35105 7515 35139
rect 7515 35105 7524 35139
rect 7472 35096 7524 35105
rect 7564 35096 7616 35148
rect 8484 35139 8536 35148
rect 8484 35105 8493 35139
rect 8493 35105 8527 35139
rect 8527 35105 8536 35139
rect 8484 35096 8536 35105
rect 9312 35096 9364 35148
rect 9404 35096 9456 35148
rect 9956 35164 10008 35216
rect 10140 35164 10192 35216
rect 10416 35164 10468 35216
rect 11796 35232 11848 35284
rect 12164 35232 12216 35284
rect 11152 35139 11204 35148
rect 11152 35105 11161 35139
rect 11161 35105 11195 35139
rect 11195 35105 11204 35139
rect 11152 35096 11204 35105
rect 11980 35164 12032 35216
rect 12256 35207 12308 35216
rect 12256 35173 12265 35207
rect 12265 35173 12299 35207
rect 12299 35173 12308 35207
rect 12256 35164 12308 35173
rect 11428 35139 11480 35148
rect 11428 35105 11437 35139
rect 11437 35105 11471 35139
rect 11471 35105 11480 35139
rect 11428 35096 11480 35105
rect 7380 35028 7432 35080
rect 9680 35071 9732 35080
rect 6644 34960 6696 35012
rect 6736 34960 6788 35012
rect 7472 34960 7524 35012
rect 7748 34960 7800 35012
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 9680 35028 9732 35037
rect 8852 34960 8904 35012
rect 9864 35028 9916 35080
rect 6368 34892 6420 34944
rect 6920 34892 6972 34944
rect 7288 34935 7340 34944
rect 7288 34901 7297 34935
rect 7297 34901 7331 34935
rect 7331 34901 7340 34935
rect 7288 34892 7340 34901
rect 7932 34935 7984 34944
rect 7932 34901 7941 34935
rect 7941 34901 7975 34935
rect 7975 34901 7984 34935
rect 7932 34892 7984 34901
rect 9312 34892 9364 34944
rect 9864 34892 9916 34944
rect 11888 35028 11940 35080
rect 11980 34960 12032 35012
rect 11336 34892 11388 34944
rect 3662 34790 3714 34842
rect 3726 34790 3778 34842
rect 3790 34790 3842 34842
rect 3854 34790 3906 34842
rect 3918 34790 3970 34842
rect 10062 34790 10114 34842
rect 10126 34790 10178 34842
rect 10190 34790 10242 34842
rect 10254 34790 10306 34842
rect 10318 34790 10370 34842
rect 1216 34688 1268 34740
rect 1400 34688 1452 34740
rect 2044 34688 2096 34740
rect 2596 34688 2648 34740
rect 3424 34688 3476 34740
rect 3700 34688 3752 34740
rect 2412 34620 2464 34672
rect 388 34484 440 34536
rect 1584 34484 1636 34536
rect 2228 34484 2280 34536
rect 4712 34620 4764 34672
rect 3056 34552 3108 34604
rect 3792 34595 3844 34604
rect 3792 34561 3801 34595
rect 3801 34561 3835 34595
rect 3835 34561 3844 34595
rect 3792 34552 3844 34561
rect 1768 34416 1820 34468
rect 3516 34416 3568 34468
rect 4252 34552 4304 34604
rect 5356 34688 5408 34740
rect 5816 34731 5868 34740
rect 5816 34697 5825 34731
rect 5825 34697 5859 34731
rect 5859 34697 5868 34731
rect 5816 34688 5868 34697
rect 7104 34688 7156 34740
rect 10140 34688 10192 34740
rect 6000 34620 6052 34672
rect 5540 34552 5592 34604
rect 5908 34552 5960 34604
rect 4068 34416 4120 34468
rect 572 34348 624 34400
rect 1860 34348 1912 34400
rect 3240 34391 3292 34400
rect 3240 34357 3249 34391
rect 3249 34357 3283 34391
rect 3283 34357 3292 34391
rect 3240 34348 3292 34357
rect 3424 34348 3476 34400
rect 3700 34391 3752 34400
rect 3700 34357 3709 34391
rect 3709 34357 3743 34391
rect 3743 34357 3752 34391
rect 3700 34348 3752 34357
rect 4160 34348 4212 34400
rect 4712 34391 4764 34400
rect 4712 34357 4721 34391
rect 4721 34357 4755 34391
rect 4755 34357 4764 34391
rect 4712 34348 4764 34357
rect 6368 34527 6420 34536
rect 6368 34493 6377 34527
rect 6377 34493 6411 34527
rect 6411 34493 6420 34527
rect 6368 34484 6420 34493
rect 6460 34527 6512 34536
rect 6460 34493 6469 34527
rect 6469 34493 6503 34527
rect 6503 34493 6512 34527
rect 6460 34484 6512 34493
rect 8852 34552 8904 34604
rect 5540 34416 5592 34468
rect 6736 34416 6788 34468
rect 6920 34416 6972 34468
rect 7380 34527 7432 34536
rect 7380 34493 7389 34527
rect 7389 34493 7423 34527
rect 7423 34493 7432 34527
rect 7380 34484 7432 34493
rect 7656 34527 7708 34536
rect 7656 34493 7665 34527
rect 7665 34493 7699 34527
rect 7699 34493 7708 34527
rect 7656 34484 7708 34493
rect 8208 34527 8260 34536
rect 8208 34493 8217 34527
rect 8217 34493 8251 34527
rect 8251 34493 8260 34527
rect 8208 34484 8260 34493
rect 7748 34416 7800 34468
rect 8024 34416 8076 34468
rect 8760 34484 8812 34536
rect 8944 34527 8996 34536
rect 8944 34493 8953 34527
rect 8953 34493 8987 34527
rect 8987 34493 8996 34527
rect 8944 34484 8996 34493
rect 9036 34527 9088 34536
rect 9036 34493 9045 34527
rect 9045 34493 9079 34527
rect 9079 34493 9088 34527
rect 9036 34484 9088 34493
rect 9772 34484 9824 34536
rect 10508 34663 10560 34672
rect 10508 34629 10517 34663
rect 10517 34629 10551 34663
rect 10551 34629 10560 34663
rect 10508 34620 10560 34629
rect 9404 34416 9456 34468
rect 9496 34416 9548 34468
rect 9956 34416 10008 34468
rect 10416 34416 10468 34468
rect 11980 34527 12032 34536
rect 11980 34493 11998 34527
rect 11998 34493 12032 34527
rect 11980 34484 12032 34493
rect 12256 34527 12308 34536
rect 12256 34493 12265 34527
rect 12265 34493 12299 34527
rect 12299 34493 12308 34527
rect 12256 34484 12308 34493
rect 6092 34348 6144 34400
rect 6368 34348 6420 34400
rect 7012 34348 7064 34400
rect 7840 34348 7892 34400
rect 9680 34348 9732 34400
rect 10600 34348 10652 34400
rect 11612 34416 11664 34468
rect 11152 34348 11204 34400
rect 11796 34348 11848 34400
rect 11980 34348 12032 34400
rect 4322 34246 4374 34298
rect 4386 34246 4438 34298
rect 4450 34246 4502 34298
rect 4514 34246 4566 34298
rect 4578 34246 4630 34298
rect 10722 34246 10774 34298
rect 10786 34246 10838 34298
rect 10850 34246 10902 34298
rect 10914 34246 10966 34298
rect 10978 34246 11030 34298
rect 3332 34144 3384 34196
rect 3608 34187 3660 34196
rect 3608 34153 3617 34187
rect 3617 34153 3651 34187
rect 3651 34153 3660 34187
rect 3608 34144 3660 34153
rect 848 34076 900 34128
rect 1216 34076 1268 34128
rect 1032 34051 1084 34060
rect 1032 34017 1041 34051
rect 1041 34017 1075 34051
rect 1075 34017 1084 34051
rect 1032 34008 1084 34017
rect 1492 34008 1544 34060
rect 1952 34008 2004 34060
rect 2228 34051 2280 34060
rect 2228 34017 2237 34051
rect 2237 34017 2271 34051
rect 2271 34017 2280 34051
rect 2228 34008 2280 34017
rect 3240 34076 3292 34128
rect 6276 34144 6328 34196
rect 6644 34144 6696 34196
rect 7564 34144 7616 34196
rect 7656 34144 7708 34196
rect 9680 34144 9732 34196
rect 3424 34008 3476 34060
rect 3976 34008 4028 34060
rect 4528 34051 4580 34060
rect 4528 34017 4562 34051
rect 4562 34017 4580 34051
rect 4528 34008 4580 34017
rect 9036 34076 9088 34128
rect 6092 34008 6144 34060
rect 7380 34008 7432 34060
rect 20 33940 72 33992
rect 848 33940 900 33992
rect 5632 33940 5684 33992
rect 2412 33804 2464 33856
rect 4252 33872 4304 33924
rect 3976 33847 4028 33856
rect 3976 33813 3985 33847
rect 3985 33813 4019 33847
rect 4019 33813 4028 33847
rect 3976 33804 4028 33813
rect 4068 33804 4120 33856
rect 8116 34051 8168 34060
rect 8116 34017 8125 34051
rect 8125 34017 8159 34051
rect 8159 34017 8168 34051
rect 8116 34008 8168 34017
rect 8024 33940 8076 33992
rect 8392 34051 8444 34060
rect 8392 34017 8401 34051
rect 8401 34017 8435 34051
rect 8435 34017 8444 34051
rect 8392 34008 8444 34017
rect 10048 34076 10100 34128
rect 9496 34008 9548 34060
rect 9588 34051 9640 34060
rect 9588 34017 9597 34051
rect 9597 34017 9631 34051
rect 9631 34017 9640 34051
rect 9588 34008 9640 34017
rect 9680 34051 9732 34060
rect 9680 34017 9689 34051
rect 9689 34017 9723 34051
rect 9723 34017 9732 34051
rect 9680 34008 9732 34017
rect 9772 34051 9824 34060
rect 9772 34017 9781 34051
rect 9781 34017 9815 34051
rect 9815 34017 9824 34051
rect 9772 34008 9824 34017
rect 9864 34051 9916 34060
rect 9864 34017 9873 34051
rect 9873 34017 9907 34051
rect 9907 34017 9916 34051
rect 9864 34008 9916 34017
rect 11244 34144 11296 34196
rect 11428 34187 11480 34196
rect 11428 34153 11437 34187
rect 11437 34153 11471 34187
rect 11471 34153 11480 34187
rect 11428 34144 11480 34153
rect 10416 34051 10468 34060
rect 10416 34017 10425 34051
rect 10425 34017 10459 34051
rect 10459 34017 10468 34051
rect 10416 34008 10468 34017
rect 11152 34008 11204 34060
rect 11888 34119 11940 34128
rect 11888 34085 11897 34119
rect 11897 34085 11931 34119
rect 11931 34085 11940 34119
rect 11888 34076 11940 34085
rect 10600 33983 10652 33992
rect 10600 33949 10609 33983
rect 10609 33949 10643 33983
rect 10643 33949 10652 33983
rect 10600 33940 10652 33949
rect 10784 33940 10836 33992
rect 11336 33940 11388 33992
rect 8484 33872 8536 33924
rect 9404 33915 9456 33924
rect 9404 33881 9413 33915
rect 9413 33881 9447 33915
rect 9447 33881 9456 33915
rect 9404 33872 9456 33881
rect 10140 33915 10192 33924
rect 10140 33881 10149 33915
rect 10149 33881 10183 33915
rect 10183 33881 10192 33915
rect 10140 33872 10192 33881
rect 11060 33915 11112 33924
rect 11060 33881 11069 33915
rect 11069 33881 11103 33915
rect 11103 33881 11112 33915
rect 11060 33872 11112 33881
rect 11152 33872 11204 33924
rect 7380 33847 7432 33856
rect 7380 33813 7389 33847
rect 7389 33813 7423 33847
rect 7423 33813 7432 33847
rect 7380 33804 7432 33813
rect 7748 33804 7800 33856
rect 9864 33804 9916 33856
rect 11428 33804 11480 33856
rect 11704 33847 11756 33856
rect 11704 33813 11713 33847
rect 11713 33813 11747 33847
rect 11747 33813 11756 33847
rect 11704 33804 11756 33813
rect 11796 33804 11848 33856
rect 3662 33702 3714 33754
rect 3726 33702 3778 33754
rect 3790 33702 3842 33754
rect 3854 33702 3906 33754
rect 3918 33702 3970 33754
rect 10062 33702 10114 33754
rect 10126 33702 10178 33754
rect 10190 33702 10242 33754
rect 10254 33702 10306 33754
rect 10318 33702 10370 33754
rect 2044 33600 2096 33652
rect 2872 33600 2924 33652
rect 4068 33600 4120 33652
rect 5816 33600 5868 33652
rect 6644 33532 6696 33584
rect 2228 33507 2280 33516
rect 2228 33473 2237 33507
rect 2237 33473 2271 33507
rect 2271 33473 2280 33507
rect 2228 33464 2280 33473
rect 2504 33507 2556 33516
rect 2504 33473 2513 33507
rect 2513 33473 2547 33507
rect 2547 33473 2556 33507
rect 2504 33464 2556 33473
rect 2320 33396 2372 33448
rect 3056 33396 3108 33448
rect 1952 33371 2004 33380
rect 1952 33337 1970 33371
rect 1970 33337 2004 33371
rect 1952 33328 2004 33337
rect 1492 33260 1544 33312
rect 3148 33328 3200 33380
rect 3516 33464 3568 33516
rect 5448 33507 5500 33516
rect 5448 33473 5457 33507
rect 5457 33473 5491 33507
rect 5491 33473 5500 33507
rect 5448 33464 5500 33473
rect 3700 33439 3752 33448
rect 3700 33405 3709 33439
rect 3709 33405 3743 33439
rect 3743 33405 3752 33439
rect 3700 33396 3752 33405
rect 5264 33396 5316 33448
rect 4160 33328 4212 33380
rect 6000 33464 6052 33516
rect 6276 33464 6328 33516
rect 7104 33464 7156 33516
rect 6368 33396 6420 33448
rect 6644 33396 6696 33448
rect 7932 33600 7984 33652
rect 10140 33600 10192 33652
rect 11888 33643 11940 33652
rect 11888 33609 11897 33643
rect 11897 33609 11931 33643
rect 11931 33609 11940 33643
rect 11888 33600 11940 33609
rect 2596 33303 2648 33312
rect 2596 33269 2605 33303
rect 2605 33269 2639 33303
rect 2639 33269 2648 33303
rect 2596 33260 2648 33269
rect 3056 33303 3108 33312
rect 3056 33269 3065 33303
rect 3065 33269 3099 33303
rect 3099 33269 3108 33303
rect 3056 33260 3108 33269
rect 4252 33260 4304 33312
rect 5264 33260 5316 33312
rect 5356 33260 5408 33312
rect 7656 33396 7708 33448
rect 7932 33439 7984 33448
rect 7932 33405 7941 33439
rect 7941 33405 7975 33439
rect 7975 33405 7984 33439
rect 7932 33396 7984 33405
rect 8392 33396 8444 33448
rect 8484 33328 8536 33380
rect 10508 33439 10560 33448
rect 10508 33405 10517 33439
rect 10517 33405 10551 33439
rect 10551 33405 10560 33439
rect 10508 33396 10560 33405
rect 12532 33396 12584 33448
rect 9680 33328 9732 33380
rect 9956 33371 10008 33380
rect 9956 33337 9965 33371
rect 9965 33337 9999 33371
rect 9999 33337 10008 33371
rect 9956 33328 10008 33337
rect 10232 33328 10284 33380
rect 11980 33371 12032 33380
rect 11980 33337 11989 33371
rect 11989 33337 12023 33371
rect 12023 33337 12032 33371
rect 11980 33328 12032 33337
rect 7380 33260 7432 33312
rect 7564 33260 7616 33312
rect 8668 33260 8720 33312
rect 12164 33303 12216 33312
rect 12164 33269 12173 33303
rect 12173 33269 12207 33303
rect 12207 33269 12216 33303
rect 12164 33260 12216 33269
rect 4322 33158 4374 33210
rect 4386 33158 4438 33210
rect 4450 33158 4502 33210
rect 4514 33158 4566 33210
rect 4578 33158 4630 33210
rect 10722 33158 10774 33210
rect 10786 33158 10838 33210
rect 10850 33158 10902 33210
rect 10914 33158 10966 33210
rect 10978 33158 11030 33210
rect 2872 33056 2924 33108
rect 4896 33099 4948 33108
rect 4896 33065 4905 33099
rect 4905 33065 4939 33099
rect 4939 33065 4948 33099
rect 4896 33056 4948 33065
rect 6460 33056 6512 33108
rect 7012 33056 7064 33108
rect 7104 33056 7156 33108
rect 1124 33031 1176 33040
rect 1124 32997 1133 33031
rect 1133 32997 1167 33031
rect 1167 32997 1176 33031
rect 1124 32988 1176 32997
rect 2228 32988 2280 33040
rect 1216 32920 1268 32972
rect 2504 32920 2556 32972
rect 3056 32988 3108 33040
rect 3424 32988 3476 33040
rect 7288 33099 7340 33108
rect 7288 33065 7297 33099
rect 7297 33065 7331 33099
rect 7331 33065 7340 33099
rect 7288 33056 7340 33065
rect 7932 33056 7984 33108
rect 8484 33099 8536 33108
rect 8484 33065 8493 33099
rect 8493 33065 8527 33099
rect 8527 33065 8536 33099
rect 8484 33056 8536 33065
rect 9312 33056 9364 33108
rect 9772 33056 9824 33108
rect 10508 33056 10560 33108
rect 4896 32963 4948 32972
rect 4896 32929 4905 32963
rect 4905 32929 4939 32963
rect 4939 32929 4948 32963
rect 4896 32920 4948 32929
rect 1492 32852 1544 32904
rect 2688 32895 2740 32904
rect 2688 32861 2697 32895
rect 2697 32861 2731 32895
rect 2731 32861 2740 32895
rect 2688 32852 2740 32861
rect 1492 32716 1544 32768
rect 3700 32784 3752 32836
rect 4436 32784 4488 32836
rect 3424 32716 3476 32768
rect 4988 32852 5040 32904
rect 5356 32963 5408 32972
rect 5356 32929 5365 32963
rect 5365 32929 5399 32963
rect 5399 32929 5408 32963
rect 5356 32920 5408 32929
rect 5816 32963 5868 32972
rect 5816 32929 5825 32963
rect 5825 32929 5859 32963
rect 5859 32929 5868 32963
rect 5816 32920 5868 32929
rect 6184 32920 6236 32972
rect 6460 32920 6512 32972
rect 6644 32963 6696 32972
rect 6644 32929 6653 32963
rect 6653 32929 6687 32963
rect 6687 32929 6696 32963
rect 6644 32920 6696 32929
rect 6828 32963 6880 32972
rect 6828 32929 6837 32963
rect 6837 32929 6871 32963
rect 6871 32929 6880 32963
rect 6828 32920 6880 32929
rect 6920 32920 6972 32972
rect 7288 32920 7340 32972
rect 5448 32852 5500 32904
rect 5540 32852 5592 32904
rect 8116 32963 8168 32972
rect 8116 32929 8125 32963
rect 8125 32929 8159 32963
rect 8159 32929 8168 32963
rect 8116 32920 8168 32929
rect 7656 32852 7708 32904
rect 8668 32963 8720 32972
rect 8668 32929 8677 32963
rect 8677 32929 8711 32963
rect 8711 32929 8720 32963
rect 8668 32920 8720 32929
rect 8760 32920 8812 32972
rect 5356 32784 5408 32836
rect 6920 32784 6972 32836
rect 7472 32784 7524 32836
rect 7932 32784 7984 32836
rect 9128 32784 9180 32836
rect 6092 32759 6144 32768
rect 6092 32725 6101 32759
rect 6101 32725 6135 32759
rect 6135 32725 6144 32759
rect 6092 32716 6144 32725
rect 6736 32716 6788 32768
rect 7104 32716 7156 32768
rect 8392 32716 8444 32768
rect 8944 32759 8996 32768
rect 8944 32725 8953 32759
rect 8953 32725 8987 32759
rect 8987 32725 8996 32759
rect 8944 32716 8996 32725
rect 9864 32988 9916 33040
rect 10692 32988 10744 33040
rect 10876 33056 10928 33108
rect 12716 33056 12768 33108
rect 9588 32920 9640 32972
rect 12256 32988 12308 33040
rect 11336 32920 11388 32972
rect 11888 32920 11940 32972
rect 11152 32852 11204 32904
rect 12164 32852 12216 32904
rect 11704 32784 11756 32836
rect 9312 32716 9364 32768
rect 9496 32716 9548 32768
rect 10140 32716 10192 32768
rect 11336 32716 11388 32768
rect 3662 32614 3714 32666
rect 3726 32614 3778 32666
rect 3790 32614 3842 32666
rect 3854 32614 3906 32666
rect 3918 32614 3970 32666
rect 10062 32614 10114 32666
rect 10126 32614 10178 32666
rect 10190 32614 10242 32666
rect 10254 32614 10306 32666
rect 10318 32614 10370 32666
rect 1124 32512 1176 32564
rect 2136 32512 2188 32564
rect 2504 32512 2556 32564
rect 1492 32487 1544 32496
rect 1492 32453 1501 32487
rect 1501 32453 1535 32487
rect 1535 32453 1544 32487
rect 1492 32444 1544 32453
rect 4896 32512 4948 32564
rect 5540 32512 5592 32564
rect 6092 32512 6144 32564
rect 6644 32555 6696 32564
rect 6644 32521 6653 32555
rect 6653 32521 6687 32555
rect 6687 32521 6696 32555
rect 6644 32512 6696 32521
rect 6828 32512 6880 32564
rect 7104 32512 7156 32564
rect 7932 32512 7984 32564
rect 4252 32376 4304 32428
rect 1216 32351 1268 32360
rect 1216 32317 1225 32351
rect 1225 32317 1259 32351
rect 1259 32317 1268 32351
rect 1216 32308 1268 32317
rect 3332 32308 3384 32360
rect 1032 32215 1084 32224
rect 1032 32181 1041 32215
rect 1041 32181 1075 32215
rect 1075 32181 1084 32215
rect 1032 32172 1084 32181
rect 1400 32172 1452 32224
rect 2412 32240 2464 32292
rect 3608 32308 3660 32360
rect 4068 32308 4120 32360
rect 4436 32351 4488 32360
rect 4436 32317 4445 32351
rect 4445 32317 4479 32351
rect 4479 32317 4488 32351
rect 4436 32308 4488 32317
rect 5356 32444 5408 32496
rect 4988 32376 5040 32428
rect 6276 32444 6328 32496
rect 7012 32444 7064 32496
rect 6184 32376 6236 32428
rect 6276 32308 6328 32360
rect 3240 32172 3292 32224
rect 3792 32172 3844 32224
rect 4160 32215 4212 32224
rect 4160 32181 4169 32215
rect 4169 32181 4203 32215
rect 4203 32181 4212 32215
rect 4160 32172 4212 32181
rect 4252 32172 4304 32224
rect 5080 32172 5132 32224
rect 6184 32240 6236 32292
rect 6460 32419 6512 32428
rect 6460 32385 6469 32419
rect 6469 32385 6503 32419
rect 6503 32385 6512 32419
rect 6460 32376 6512 32385
rect 6828 32308 6880 32360
rect 7564 32351 7616 32360
rect 7564 32317 7573 32351
rect 7573 32317 7607 32351
rect 7607 32317 7616 32351
rect 7564 32308 7616 32317
rect 7840 32419 7892 32428
rect 7840 32385 7849 32419
rect 7849 32385 7883 32419
rect 7883 32385 7892 32419
rect 7840 32376 7892 32385
rect 8300 32444 8352 32496
rect 8576 32444 8628 32496
rect 8760 32444 8812 32496
rect 9588 32512 9640 32564
rect 10600 32512 10652 32564
rect 9404 32487 9456 32496
rect 9404 32453 9413 32487
rect 9413 32453 9447 32487
rect 9447 32453 9456 32487
rect 9404 32444 9456 32453
rect 7012 32240 7064 32292
rect 5908 32172 5960 32224
rect 6552 32172 6604 32224
rect 7288 32172 7340 32224
rect 7472 32172 7524 32224
rect 7840 32240 7892 32292
rect 7932 32172 7984 32224
rect 8944 32376 8996 32428
rect 9680 32444 9732 32496
rect 10232 32444 10284 32496
rect 9864 32419 9916 32428
rect 9864 32385 9873 32419
rect 9873 32385 9907 32419
rect 9907 32385 9916 32419
rect 9864 32376 9916 32385
rect 9128 32240 9180 32292
rect 9680 32351 9732 32360
rect 9680 32317 9689 32351
rect 9689 32317 9723 32351
rect 9723 32317 9732 32351
rect 9680 32308 9732 32317
rect 11796 32376 11848 32428
rect 10232 32308 10284 32360
rect 12256 32351 12308 32360
rect 12256 32317 12265 32351
rect 12265 32317 12299 32351
rect 12299 32317 12308 32351
rect 12256 32308 12308 32317
rect 10600 32240 10652 32292
rect 10140 32172 10192 32224
rect 11520 32172 11572 32224
rect 11888 32172 11940 32224
rect 12164 32172 12216 32224
rect 4322 32070 4374 32122
rect 4386 32070 4438 32122
rect 4450 32070 4502 32122
rect 4514 32070 4566 32122
rect 4578 32070 4630 32122
rect 10722 32070 10774 32122
rect 10786 32070 10838 32122
rect 10850 32070 10902 32122
rect 10914 32070 10966 32122
rect 10978 32070 11030 32122
rect 572 31968 624 32020
rect 388 31832 440 31884
rect 572 31832 624 31884
rect 848 31900 900 31952
rect 1032 31900 1084 31952
rect 1676 31968 1728 32020
rect 2044 31968 2096 32020
rect 2320 31943 2372 31952
rect 2320 31909 2329 31943
rect 2329 31909 2363 31943
rect 2363 31909 2372 31943
rect 2320 31900 2372 31909
rect 2412 31900 2464 31952
rect 1216 31832 1268 31884
rect 1952 31832 2004 31884
rect 2136 31832 2188 31884
rect 2228 31875 2280 31884
rect 2228 31841 2237 31875
rect 2237 31841 2271 31875
rect 2271 31841 2280 31875
rect 2228 31832 2280 31841
rect 2596 31875 2648 31884
rect 2596 31841 2605 31875
rect 2605 31841 2639 31875
rect 2639 31841 2648 31875
rect 2596 31832 2648 31841
rect 2872 31875 2924 31884
rect 2872 31841 2881 31875
rect 2881 31841 2915 31875
rect 2915 31841 2924 31875
rect 2872 31832 2924 31841
rect 5448 31968 5500 32020
rect 5908 31968 5960 32020
rect 6644 31968 6696 32020
rect 7012 31968 7064 32020
rect 3792 31900 3844 31952
rect 756 31764 808 31816
rect 1492 31764 1544 31816
rect 2504 31764 2556 31816
rect 3240 31807 3292 31816
rect 3240 31773 3249 31807
rect 3249 31773 3283 31807
rect 3283 31773 3292 31807
rect 3240 31764 3292 31773
rect 3424 31764 3476 31816
rect 4620 31832 4672 31884
rect 4988 31832 5040 31884
rect 5080 31875 5132 31884
rect 5080 31841 5089 31875
rect 5089 31841 5123 31875
rect 5123 31841 5132 31875
rect 5080 31832 5132 31841
rect 6092 31900 6144 31952
rect 6368 31900 6420 31952
rect 6736 31900 6788 31952
rect 5448 31875 5500 31884
rect 5448 31841 5457 31875
rect 5457 31841 5491 31875
rect 5491 31841 5500 31875
rect 5448 31832 5500 31841
rect 5540 31875 5592 31884
rect 5540 31841 5549 31875
rect 5549 31841 5583 31875
rect 5583 31841 5592 31875
rect 5540 31832 5592 31841
rect 6000 31832 6052 31884
rect 6276 31875 6328 31884
rect 6276 31841 6285 31875
rect 6285 31841 6319 31875
rect 6319 31841 6328 31875
rect 6276 31832 6328 31841
rect 5356 31807 5408 31816
rect 5356 31773 5365 31807
rect 5365 31773 5399 31807
rect 5399 31773 5408 31807
rect 5356 31764 5408 31773
rect 6368 31807 6420 31816
rect 6368 31773 6377 31807
rect 6377 31773 6411 31807
rect 6411 31773 6420 31807
rect 6368 31764 6420 31773
rect 6460 31764 6512 31816
rect 6644 31875 6696 31884
rect 6644 31841 6653 31875
rect 6653 31841 6687 31875
rect 6687 31841 6696 31875
rect 6644 31832 6696 31841
rect 7564 31900 7616 31952
rect 7932 31968 7984 32020
rect 8116 31968 8168 32020
rect 8208 31968 8260 32020
rect 8484 31968 8536 32020
rect 8576 31968 8628 32020
rect 8392 31900 8444 31952
rect 8300 31875 8352 31884
rect 1216 31628 1268 31680
rect 2780 31628 2832 31680
rect 4160 31696 4212 31748
rect 4712 31696 4764 31748
rect 5448 31696 5500 31748
rect 7012 31696 7064 31748
rect 7932 31764 7984 31816
rect 8300 31841 8309 31875
rect 8309 31841 8343 31875
rect 8343 31841 8352 31875
rect 8300 31832 8352 31841
rect 8576 31875 8628 31884
rect 8576 31841 8585 31875
rect 8585 31841 8619 31875
rect 8619 31841 8628 31875
rect 8576 31832 8628 31841
rect 8760 31900 8812 31952
rect 8944 31900 8996 31952
rect 9496 31968 9548 32020
rect 8944 31764 8996 31816
rect 9128 31832 9180 31884
rect 10876 31900 10928 31952
rect 9404 31832 9456 31884
rect 10968 31875 11020 31884
rect 10968 31841 10977 31875
rect 10977 31841 11011 31875
rect 11011 31841 11020 31875
rect 10968 31832 11020 31841
rect 11612 31832 11664 31884
rect 11796 31832 11848 31884
rect 8760 31696 8812 31748
rect 10876 31696 10928 31748
rect 4068 31671 4120 31680
rect 4068 31637 4077 31671
rect 4077 31637 4111 31671
rect 4111 31637 4120 31671
rect 4068 31628 4120 31637
rect 4436 31671 4488 31680
rect 4436 31637 4445 31671
rect 4445 31637 4479 31671
rect 4479 31637 4488 31671
rect 4436 31628 4488 31637
rect 5908 31628 5960 31680
rect 7104 31628 7156 31680
rect 7288 31628 7340 31680
rect 7564 31628 7616 31680
rect 7932 31628 7984 31680
rect 8208 31628 8260 31680
rect 8300 31628 8352 31680
rect 10692 31671 10744 31680
rect 10692 31637 10701 31671
rect 10701 31637 10735 31671
rect 10735 31637 10744 31671
rect 10692 31628 10744 31637
rect 11152 31671 11204 31680
rect 11152 31637 11161 31671
rect 11161 31637 11195 31671
rect 11195 31637 11204 31671
rect 11152 31628 11204 31637
rect 11520 31696 11572 31748
rect 12532 31764 12584 31816
rect 12348 31696 12400 31748
rect 12256 31628 12308 31680
rect 3662 31526 3714 31578
rect 3726 31526 3778 31578
rect 3790 31526 3842 31578
rect 3854 31526 3906 31578
rect 3918 31526 3970 31578
rect 10062 31526 10114 31578
rect 10126 31526 10178 31578
rect 10190 31526 10242 31578
rect 10254 31526 10306 31578
rect 10318 31526 10370 31578
rect 1492 31424 1544 31476
rect 2228 31424 2280 31476
rect 3240 31424 3292 31476
rect 3424 31467 3476 31476
rect 3424 31433 3433 31467
rect 3433 31433 3467 31467
rect 3467 31433 3476 31467
rect 3424 31424 3476 31433
rect 5356 31424 5408 31476
rect 5816 31424 5868 31476
rect 6920 31424 6972 31476
rect 8944 31424 8996 31476
rect 10140 31424 10192 31476
rect 10416 31467 10468 31476
rect 10416 31433 10425 31467
rect 10425 31433 10459 31467
rect 10459 31433 10468 31467
rect 10416 31424 10468 31433
rect 1952 31263 2004 31272
rect 1952 31229 1970 31263
rect 1970 31229 2004 31263
rect 1952 31220 2004 31229
rect 1676 31152 1728 31204
rect 2228 31263 2280 31272
rect 2228 31229 2237 31263
rect 2237 31229 2271 31263
rect 2271 31229 2280 31263
rect 2688 31356 2740 31408
rect 5540 31356 5592 31408
rect 3148 31288 3200 31340
rect 2228 31220 2280 31229
rect 2688 31263 2740 31272
rect 2688 31229 2697 31263
rect 2697 31229 2731 31263
rect 2731 31229 2740 31263
rect 2688 31220 2740 31229
rect 3332 31220 3384 31272
rect 1492 31084 1544 31136
rect 2504 31152 2556 31204
rect 3148 31152 3200 31204
rect 3792 31263 3844 31272
rect 3792 31229 3801 31263
rect 3801 31229 3835 31263
rect 3835 31229 3844 31263
rect 3792 31220 3844 31229
rect 4528 31220 4580 31272
rect 5816 31288 5868 31340
rect 6000 31288 6052 31340
rect 7196 31356 7248 31408
rect 4436 31152 4488 31204
rect 5816 31152 5868 31204
rect 3056 31084 3108 31136
rect 4620 31084 4672 31136
rect 5264 31084 5316 31136
rect 6460 31263 6512 31272
rect 6460 31229 6469 31263
rect 6469 31229 6503 31263
rect 6503 31229 6512 31263
rect 6460 31220 6512 31229
rect 6552 31263 6604 31272
rect 6552 31229 6561 31263
rect 6561 31229 6595 31263
rect 6595 31229 6604 31263
rect 6552 31220 6604 31229
rect 6736 31220 6788 31272
rect 6920 31220 6972 31272
rect 7196 31220 7248 31272
rect 7288 31263 7340 31272
rect 7288 31229 7297 31263
rect 7297 31229 7331 31263
rect 7331 31229 7340 31263
rect 7288 31220 7340 31229
rect 7656 31220 7708 31272
rect 8116 31220 8168 31272
rect 10876 31331 10928 31340
rect 10876 31297 10885 31331
rect 10885 31297 10919 31331
rect 10919 31297 10928 31331
rect 10876 31288 10928 31297
rect 9128 31220 9180 31272
rect 9772 31220 9824 31272
rect 11152 31263 11204 31272
rect 11152 31229 11186 31263
rect 11186 31229 11204 31263
rect 11152 31220 11204 31229
rect 7564 31152 7616 31204
rect 8300 31152 8352 31204
rect 8944 31152 8996 31204
rect 9588 31152 9640 31204
rect 7012 31084 7064 31136
rect 7656 31084 7708 31136
rect 7840 31127 7892 31136
rect 7840 31093 7849 31127
rect 7849 31093 7883 31127
rect 7883 31093 7892 31127
rect 7840 31084 7892 31093
rect 9128 31084 9180 31136
rect 11152 31084 11204 31136
rect 11428 31084 11480 31136
rect 4322 30982 4374 31034
rect 4386 30982 4438 31034
rect 4450 30982 4502 31034
rect 4514 30982 4566 31034
rect 4578 30982 4630 31034
rect 10722 30982 10774 31034
rect 10786 30982 10838 31034
rect 10850 30982 10902 31034
rect 10914 30982 10966 31034
rect 10978 30982 11030 31034
rect 2780 30880 2832 30932
rect 940 30812 992 30864
rect 2596 30812 2648 30864
rect 1400 30744 1452 30796
rect 2412 30744 2464 30796
rect 3148 30744 3200 30796
rect 3516 30880 3568 30932
rect 4436 30880 4488 30932
rect 4712 30880 4764 30932
rect 5172 30880 5224 30932
rect 5356 30880 5408 30932
rect 4068 30812 4120 30864
rect 6460 30880 6512 30932
rect 7104 30880 7156 30932
rect 7840 30880 7892 30932
rect 8576 30880 8628 30932
rect 9588 30923 9640 30932
rect 9588 30889 9597 30923
rect 9597 30889 9631 30923
rect 9631 30889 9640 30923
rect 9588 30880 9640 30889
rect 3516 30787 3568 30796
rect 3516 30753 3525 30787
rect 3525 30753 3559 30787
rect 3559 30753 3568 30787
rect 3516 30744 3568 30753
rect 2228 30719 2280 30728
rect 2228 30685 2237 30719
rect 2237 30685 2271 30719
rect 2271 30685 2280 30719
rect 3792 30744 3844 30796
rect 5356 30787 5408 30796
rect 5356 30753 5365 30787
rect 5365 30753 5399 30787
rect 5399 30753 5408 30787
rect 5356 30744 5408 30753
rect 2228 30676 2280 30685
rect 5264 30676 5316 30728
rect 6368 30744 6420 30796
rect 6460 30787 6512 30796
rect 6460 30753 6469 30787
rect 6469 30753 6503 30787
rect 6503 30753 6512 30787
rect 6460 30744 6512 30753
rect 7012 30787 7064 30796
rect 7012 30753 7021 30787
rect 7021 30753 7055 30787
rect 7055 30753 7064 30787
rect 7012 30744 7064 30753
rect 8668 30812 8720 30864
rect 7472 30787 7524 30796
rect 7472 30753 7481 30787
rect 7481 30753 7515 30787
rect 7515 30753 7524 30787
rect 7472 30744 7524 30753
rect 7656 30787 7708 30796
rect 7656 30753 7665 30787
rect 7665 30753 7699 30787
rect 7699 30753 7708 30787
rect 7656 30744 7708 30753
rect 7840 30787 7892 30796
rect 7840 30753 7849 30787
rect 7849 30753 7883 30787
rect 7883 30753 7892 30787
rect 7840 30744 7892 30753
rect 8116 30787 8168 30796
rect 8116 30753 8125 30787
rect 8125 30753 8159 30787
rect 8159 30753 8168 30787
rect 8116 30744 8168 30753
rect 8208 30787 8260 30796
rect 8208 30753 8217 30787
rect 8217 30753 8251 30787
rect 8251 30753 8260 30787
rect 8208 30744 8260 30753
rect 6000 30608 6052 30660
rect 7288 30676 7340 30728
rect 7564 30676 7616 30728
rect 8668 30676 8720 30728
rect 8852 30812 8904 30864
rect 9312 30855 9364 30864
rect 9312 30821 9321 30855
rect 9321 30821 9355 30855
rect 9355 30821 9364 30855
rect 9312 30812 9364 30821
rect 9128 30787 9180 30796
rect 9128 30753 9137 30787
rect 9137 30753 9171 30787
rect 9171 30753 9180 30787
rect 9128 30744 9180 30753
rect 10232 30812 10284 30864
rect 10600 30880 10652 30932
rect 11612 30880 11664 30932
rect 10692 30812 10744 30864
rect 10048 30787 10100 30796
rect 10048 30753 10057 30787
rect 10057 30753 10091 30787
rect 10091 30753 10100 30787
rect 10048 30744 10100 30753
rect 10140 30787 10192 30796
rect 10140 30753 10150 30787
rect 10150 30753 10184 30787
rect 10184 30753 10192 30787
rect 10140 30744 10192 30753
rect 11704 30812 11756 30864
rect 11336 30744 11388 30796
rect 11612 30744 11664 30796
rect 20 30540 72 30592
rect 572 30540 624 30592
rect 848 30583 900 30592
rect 848 30549 857 30583
rect 857 30549 891 30583
rect 891 30549 900 30583
rect 848 30540 900 30549
rect 1860 30540 1912 30592
rect 2872 30540 2924 30592
rect 4620 30540 4672 30592
rect 4712 30540 4764 30592
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 5724 30540 5776 30592
rect 7472 30608 7524 30660
rect 7656 30608 7708 30660
rect 7840 30608 7892 30660
rect 9404 30676 9456 30728
rect 9864 30676 9916 30728
rect 10968 30676 11020 30728
rect 8944 30608 8996 30660
rect 9588 30608 9640 30660
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 11888 30719 11940 30728
rect 11888 30685 11897 30719
rect 11897 30685 11931 30719
rect 11931 30685 11940 30719
rect 11888 30676 11940 30685
rect 12348 30676 12400 30728
rect 12624 30676 12676 30728
rect 8300 30540 8352 30592
rect 10416 30540 10468 30592
rect 11704 30540 11756 30592
rect 11888 30540 11940 30592
rect 3662 30438 3714 30490
rect 3726 30438 3778 30490
rect 3790 30438 3842 30490
rect 3854 30438 3906 30490
rect 3918 30438 3970 30490
rect 10062 30438 10114 30490
rect 10126 30438 10178 30490
rect 10190 30438 10242 30490
rect 10254 30438 10306 30490
rect 10318 30438 10370 30490
rect 572 30268 624 30320
rect 664 30268 716 30320
rect 1124 30268 1176 30320
rect 1952 30336 2004 30388
rect 848 30132 900 30184
rect 1400 30132 1452 30184
rect 1124 30064 1176 30116
rect 2412 30268 2464 30320
rect 3792 30336 3844 30388
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 3240 30200 3292 30252
rect 5632 30336 5684 30388
rect 6000 30336 6052 30388
rect 6552 30336 6604 30388
rect 6736 30379 6788 30388
rect 6736 30345 6745 30379
rect 6745 30345 6779 30379
rect 6779 30345 6788 30379
rect 6736 30336 6788 30345
rect 7012 30336 7064 30388
rect 7196 30336 7248 30388
rect 7840 30336 7892 30388
rect 9496 30336 9548 30388
rect 4160 30268 4212 30320
rect 4712 30268 4764 30320
rect 2320 30132 2372 30184
rect 2412 30175 2464 30184
rect 2412 30141 2421 30175
rect 2421 30141 2455 30175
rect 2455 30141 2464 30175
rect 2412 30132 2464 30141
rect 2596 30132 2648 30184
rect 3332 30132 3384 30184
rect 2688 30107 2740 30116
rect 2688 30073 2697 30107
rect 2697 30073 2731 30107
rect 2731 30073 2740 30107
rect 2688 30064 2740 30073
rect 2780 30064 2832 30116
rect 1400 29996 1452 30048
rect 3424 29996 3476 30048
rect 3700 30175 3752 30184
rect 3700 30141 3709 30175
rect 3709 30141 3743 30175
rect 3743 30141 3752 30175
rect 3700 30132 3752 30141
rect 4160 30132 4212 30184
rect 4436 30132 4488 30184
rect 4988 30132 5040 30184
rect 5540 30132 5592 30184
rect 5816 30268 5868 30320
rect 6920 30268 6972 30320
rect 8760 30311 8812 30320
rect 8760 30277 8769 30311
rect 8769 30277 8803 30311
rect 8803 30277 8812 30311
rect 8760 30268 8812 30277
rect 5724 30132 5776 30184
rect 6736 30200 6788 30252
rect 3976 30064 4028 30116
rect 6276 30175 6328 30184
rect 6276 30141 6285 30175
rect 6285 30141 6319 30175
rect 6319 30141 6328 30175
rect 6276 30132 6328 30141
rect 6644 30132 6696 30184
rect 7104 30175 7156 30184
rect 7104 30141 7113 30175
rect 7113 30141 7147 30175
rect 7147 30141 7156 30175
rect 7104 30132 7156 30141
rect 7288 30175 7340 30184
rect 7288 30141 7297 30175
rect 7297 30141 7331 30175
rect 7331 30141 7340 30175
rect 7932 30200 7984 30252
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 9496 30200 9548 30252
rect 10232 30311 10284 30320
rect 10232 30277 10241 30311
rect 10241 30277 10275 30311
rect 10275 30277 10284 30311
rect 10232 30268 10284 30277
rect 10784 30336 10836 30388
rect 11612 30336 11664 30388
rect 10600 30268 10652 30320
rect 7288 30132 7340 30141
rect 3884 29996 3936 30048
rect 4528 29996 4580 30048
rect 4620 29996 4672 30048
rect 4804 30039 4856 30048
rect 4804 30005 4813 30039
rect 4813 30005 4847 30039
rect 4847 30005 4856 30039
rect 4804 29996 4856 30005
rect 6920 30064 6972 30116
rect 7012 30064 7064 30116
rect 7840 30132 7892 30184
rect 8116 30175 8168 30184
rect 8116 30141 8125 30175
rect 8125 30141 8159 30175
rect 8159 30141 8168 30175
rect 8116 30132 8168 30141
rect 5540 29996 5592 30048
rect 8484 30132 8536 30184
rect 8300 30064 8352 30116
rect 8852 30175 8904 30184
rect 8852 30141 8861 30175
rect 8861 30141 8895 30175
rect 8895 30141 8904 30175
rect 8852 30132 8904 30141
rect 8944 30175 8996 30184
rect 8944 30141 8953 30175
rect 8953 30141 8987 30175
rect 8987 30141 8996 30175
rect 8944 30132 8996 30141
rect 9220 30132 9272 30184
rect 9956 30132 10008 30184
rect 12256 30243 12308 30252
rect 12256 30209 12265 30243
rect 12265 30209 12299 30243
rect 12299 30209 12308 30243
rect 12256 30200 12308 30209
rect 8852 29996 8904 30048
rect 9220 29996 9272 30048
rect 10232 30064 10284 30116
rect 9956 30039 10008 30048
rect 9956 30005 9965 30039
rect 9965 30005 9999 30039
rect 9999 30005 10008 30039
rect 9956 29996 10008 30005
rect 10324 29996 10376 30048
rect 11704 30132 11756 30184
rect 11520 30064 11572 30116
rect 12256 29996 12308 30048
rect 4322 29894 4374 29946
rect 4386 29894 4438 29946
rect 4450 29894 4502 29946
rect 4514 29894 4566 29946
rect 4578 29894 4630 29946
rect 10722 29894 10774 29946
rect 10786 29894 10838 29946
rect 10850 29894 10902 29946
rect 10914 29894 10966 29946
rect 10978 29894 11030 29946
rect 480 29792 532 29844
rect 1492 29835 1544 29844
rect 1492 29801 1501 29835
rect 1501 29801 1535 29835
rect 1535 29801 1544 29835
rect 1492 29792 1544 29801
rect 1768 29835 1820 29844
rect 1768 29801 1777 29835
rect 1777 29801 1811 29835
rect 1811 29801 1820 29835
rect 1768 29792 1820 29801
rect 2136 29792 2188 29844
rect 2320 29792 2372 29844
rect 2412 29792 2464 29844
rect 3516 29792 3568 29844
rect 3792 29792 3844 29844
rect 1676 29767 1728 29776
rect 1676 29733 1685 29767
rect 1685 29733 1719 29767
rect 1719 29733 1728 29767
rect 1676 29724 1728 29733
rect 2688 29724 2740 29776
rect 4160 29792 4212 29844
rect 4988 29835 5040 29844
rect 4988 29801 4997 29835
rect 4997 29801 5031 29835
rect 5031 29801 5040 29835
rect 4988 29792 5040 29801
rect 5448 29792 5500 29844
rect 5724 29792 5776 29844
rect 6092 29792 6144 29844
rect 7104 29792 7156 29844
rect 7656 29792 7708 29844
rect 8116 29792 8168 29844
rect 9404 29792 9456 29844
rect 10140 29792 10192 29844
rect 10324 29792 10376 29844
rect 10508 29792 10560 29844
rect 11888 29835 11940 29844
rect 1032 29656 1084 29708
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 1768 29588 1820 29640
rect 2412 29699 2464 29708
rect 2412 29665 2421 29699
rect 2421 29665 2455 29699
rect 2455 29665 2464 29699
rect 2412 29656 2464 29665
rect 2504 29656 2556 29708
rect 3148 29699 3200 29708
rect 2688 29631 2740 29640
rect 2688 29597 2697 29631
rect 2697 29597 2731 29631
rect 2731 29597 2740 29631
rect 2688 29588 2740 29597
rect 3148 29665 3157 29699
rect 3157 29665 3191 29699
rect 3191 29665 3200 29699
rect 3148 29656 3200 29665
rect 4068 29724 4120 29776
rect 3608 29656 3660 29708
rect 3424 29631 3476 29640
rect 3424 29597 3433 29631
rect 3433 29597 3467 29631
rect 3467 29597 3476 29631
rect 3424 29588 3476 29597
rect 4252 29699 4304 29708
rect 4252 29665 4261 29699
rect 4261 29665 4295 29699
rect 4295 29665 4304 29699
rect 4252 29656 4304 29665
rect 5356 29656 5408 29708
rect 1860 29520 1912 29572
rect 2320 29520 2372 29572
rect 388 29452 440 29504
rect 3976 29588 4028 29640
rect 5080 29588 5132 29640
rect 5816 29699 5868 29708
rect 5816 29665 5825 29699
rect 5825 29665 5859 29699
rect 5859 29665 5868 29699
rect 5816 29656 5868 29665
rect 5908 29656 5960 29708
rect 6092 29656 6144 29708
rect 6184 29599 6236 29651
rect 7380 29724 7432 29776
rect 8944 29724 8996 29776
rect 6552 29656 6604 29708
rect 7748 29656 7800 29708
rect 7932 29656 7984 29708
rect 8116 29656 8168 29708
rect 8484 29656 8536 29708
rect 9220 29699 9272 29708
rect 9220 29665 9229 29699
rect 9229 29665 9263 29699
rect 9263 29665 9272 29699
rect 9220 29656 9272 29665
rect 9680 29656 9732 29708
rect 10600 29699 10652 29708
rect 10600 29665 10609 29699
rect 10609 29665 10643 29699
rect 10643 29665 10652 29699
rect 10600 29656 10652 29665
rect 6920 29588 6972 29640
rect 4804 29520 4856 29572
rect 5264 29520 5316 29572
rect 7380 29588 7432 29640
rect 2872 29452 2924 29504
rect 4160 29452 4212 29504
rect 4620 29452 4672 29504
rect 5356 29495 5408 29504
rect 5356 29461 5365 29495
rect 5365 29461 5399 29495
rect 5399 29461 5408 29495
rect 5356 29452 5408 29461
rect 5632 29452 5684 29504
rect 6092 29452 6144 29504
rect 7564 29520 7616 29572
rect 7840 29520 7892 29572
rect 10232 29588 10284 29640
rect 11060 29656 11112 29708
rect 11888 29801 11915 29835
rect 11915 29801 11940 29835
rect 11888 29792 11940 29801
rect 11704 29724 11756 29776
rect 11612 29699 11664 29708
rect 11612 29665 11621 29699
rect 11621 29665 11655 29699
rect 11655 29665 11664 29699
rect 11612 29656 11664 29665
rect 12256 29588 12308 29640
rect 6552 29495 6604 29504
rect 6552 29461 6561 29495
rect 6561 29461 6595 29495
rect 6595 29461 6604 29495
rect 6552 29452 6604 29461
rect 8208 29452 8260 29504
rect 11336 29520 11388 29572
rect 10784 29452 10836 29504
rect 11612 29452 11664 29504
rect 3662 29350 3714 29402
rect 3726 29350 3778 29402
rect 3790 29350 3842 29402
rect 3854 29350 3906 29402
rect 3918 29350 3970 29402
rect 10062 29350 10114 29402
rect 10126 29350 10178 29402
rect 10190 29350 10242 29402
rect 10254 29350 10306 29402
rect 10318 29350 10370 29402
rect 2320 29291 2372 29300
rect 2320 29257 2329 29291
rect 2329 29257 2363 29291
rect 2363 29257 2372 29291
rect 2320 29248 2372 29257
rect 2872 29248 2924 29300
rect 5080 29248 5132 29300
rect 8760 29248 8812 29300
rect 1584 29180 1636 29232
rect 1860 29180 1912 29232
rect 1952 29180 2004 29232
rect 940 29112 992 29164
rect 1584 29044 1636 29096
rect 1952 29044 2004 29096
rect 2504 29087 2556 29096
rect 2504 29053 2513 29087
rect 2513 29053 2547 29087
rect 2547 29053 2556 29087
rect 2504 29044 2556 29053
rect 2596 29044 2648 29096
rect 2964 29044 3016 29096
rect 3424 29044 3476 29096
rect 5540 29180 5592 29232
rect 4804 29155 4856 29164
rect 4804 29121 4813 29155
rect 4813 29121 4847 29155
rect 4847 29121 4856 29155
rect 4804 29112 4856 29121
rect 5632 29112 5684 29164
rect 6000 29112 6052 29164
rect 3700 29087 3752 29096
rect 3700 29053 3709 29087
rect 3709 29053 3743 29087
rect 3743 29053 3752 29087
rect 3700 29044 3752 29053
rect 3976 29044 4028 29096
rect 4712 29044 4764 29096
rect 5172 29044 5224 29096
rect 5724 29044 5776 29096
rect 1032 29019 1084 29028
rect 1032 28985 1041 29019
rect 1041 28985 1075 29019
rect 1075 28985 1084 29019
rect 1032 28976 1084 28985
rect 2688 29019 2740 29028
rect 2688 28985 2697 29019
rect 2697 28985 2731 29019
rect 2731 28985 2740 29019
rect 2688 28976 2740 28985
rect 3424 28908 3476 28960
rect 3884 28908 3936 28960
rect 3976 28908 4028 28960
rect 5448 28976 5500 29028
rect 4252 28908 4304 28960
rect 5632 28908 5684 28960
rect 5724 28908 5776 28960
rect 6368 29044 6420 29096
rect 6644 29044 6696 29096
rect 6920 29044 6972 29096
rect 8484 29180 8536 29232
rect 9036 29112 9088 29164
rect 9496 29155 9548 29164
rect 9496 29121 9505 29155
rect 9505 29121 9539 29155
rect 9539 29121 9548 29155
rect 9496 29112 9548 29121
rect 9680 29112 9732 29164
rect 10968 29248 11020 29300
rect 11060 29291 11112 29300
rect 11060 29257 11069 29291
rect 11069 29257 11103 29291
rect 11103 29257 11112 29291
rect 11060 29248 11112 29257
rect 11336 29248 11388 29300
rect 11520 29291 11572 29300
rect 11520 29257 11529 29291
rect 11529 29257 11563 29291
rect 11563 29257 11572 29291
rect 11520 29248 11572 29257
rect 11980 29248 12032 29300
rect 10508 29180 10560 29232
rect 8668 29044 8720 29096
rect 8760 29087 8812 29096
rect 8760 29053 8769 29087
rect 8769 29053 8803 29087
rect 8803 29053 8812 29087
rect 8760 29044 8812 29053
rect 6828 29019 6880 29028
rect 6828 28985 6837 29019
rect 6837 28985 6871 29019
rect 6871 28985 6880 29019
rect 6828 28976 6880 28985
rect 7104 28976 7156 29028
rect 8024 28976 8076 29028
rect 10416 29087 10468 29096
rect 10416 29053 10425 29087
rect 10425 29053 10459 29087
rect 10459 29053 10468 29087
rect 10416 29044 10468 29053
rect 10600 29087 10652 29096
rect 10600 29053 10609 29087
rect 10609 29053 10643 29087
rect 10643 29053 10652 29087
rect 10600 29044 10652 29053
rect 10784 29155 10836 29164
rect 10784 29121 10793 29155
rect 10793 29121 10827 29155
rect 10827 29121 10836 29155
rect 10784 29112 10836 29121
rect 7288 28908 7340 28960
rect 7472 28908 7524 28960
rect 7564 28951 7616 28960
rect 7564 28917 7573 28951
rect 7573 28917 7607 28951
rect 7607 28917 7616 28951
rect 7564 28908 7616 28917
rect 7840 28908 7892 28960
rect 8208 28908 8260 28960
rect 8484 28908 8536 28960
rect 8852 28908 8904 28960
rect 9312 28908 9364 28960
rect 9864 28908 9916 28960
rect 10048 28976 10100 29028
rect 10508 28976 10560 29028
rect 11244 29087 11296 29096
rect 11244 29053 11253 29087
rect 11253 29053 11287 29087
rect 11287 29053 11296 29087
rect 11244 29044 11296 29053
rect 11428 29087 11480 29096
rect 11428 29053 11437 29087
rect 11437 29053 11471 29087
rect 11471 29053 11480 29087
rect 11428 29044 11480 29053
rect 12716 29180 12768 29232
rect 12532 29112 12584 29164
rect 11612 29044 11664 29096
rect 11796 28976 11848 29028
rect 4322 28806 4374 28858
rect 4386 28806 4438 28858
rect 4450 28806 4502 28858
rect 4514 28806 4566 28858
rect 4578 28806 4630 28858
rect 10722 28806 10774 28858
rect 10786 28806 10838 28858
rect 10850 28806 10902 28858
rect 10914 28806 10966 28858
rect 10978 28806 11030 28858
rect 2688 28704 2740 28756
rect 4252 28747 4304 28756
rect 4252 28713 4261 28747
rect 4261 28713 4295 28747
rect 4295 28713 4304 28747
rect 4252 28704 4304 28713
rect 5540 28704 5592 28756
rect 5908 28704 5960 28756
rect 7564 28704 7616 28756
rect 2320 28679 2372 28688
rect 2320 28645 2329 28679
rect 2329 28645 2363 28679
rect 2363 28645 2372 28679
rect 2320 28636 2372 28645
rect 296 28568 348 28620
rect 3148 28636 3200 28688
rect 3976 28636 4028 28688
rect 4712 28636 4764 28688
rect 848 28543 900 28552
rect 848 28509 857 28543
rect 857 28509 891 28543
rect 891 28509 900 28543
rect 848 28500 900 28509
rect 1860 28500 1912 28552
rect 2872 28364 2924 28416
rect 3240 28568 3292 28620
rect 3792 28611 3844 28620
rect 3792 28577 3801 28611
rect 3801 28577 3835 28611
rect 3835 28577 3844 28611
rect 3792 28568 3844 28577
rect 3884 28611 3936 28620
rect 3884 28577 3893 28611
rect 3893 28577 3927 28611
rect 3927 28577 3936 28611
rect 3884 28568 3936 28577
rect 3240 28432 3292 28484
rect 3976 28500 4028 28552
rect 5172 28636 5224 28688
rect 5724 28636 5776 28688
rect 6276 28636 6328 28688
rect 5816 28568 5868 28620
rect 4528 28500 4580 28552
rect 6000 28568 6052 28620
rect 6644 28568 6696 28620
rect 7472 28568 7524 28620
rect 7748 28636 7800 28688
rect 7840 28568 7892 28620
rect 8208 28611 8260 28620
rect 8208 28577 8217 28611
rect 8217 28577 8251 28611
rect 8251 28577 8260 28611
rect 8208 28568 8260 28577
rect 6552 28500 6604 28552
rect 6368 28432 6420 28484
rect 7840 28475 7892 28484
rect 7840 28441 7849 28475
rect 7849 28441 7883 28475
rect 7883 28441 7892 28475
rect 7840 28432 7892 28441
rect 8668 28747 8720 28756
rect 8668 28713 8677 28747
rect 8677 28713 8711 28747
rect 8711 28713 8720 28747
rect 8668 28704 8720 28713
rect 9588 28704 9640 28756
rect 8852 28679 8904 28688
rect 8852 28645 8861 28679
rect 8861 28645 8895 28679
rect 8895 28645 8904 28679
rect 8852 28636 8904 28645
rect 8944 28636 8996 28688
rect 11704 28704 11756 28756
rect 11980 28704 12032 28756
rect 12072 28704 12124 28756
rect 8760 28568 8812 28620
rect 9128 28611 9180 28620
rect 9128 28577 9137 28611
rect 9137 28577 9171 28611
rect 9171 28577 9180 28611
rect 9128 28568 9180 28577
rect 9312 28611 9364 28620
rect 9312 28577 9321 28611
rect 9321 28577 9355 28611
rect 9355 28577 9364 28611
rect 9312 28568 9364 28577
rect 9680 28568 9732 28620
rect 9864 28611 9916 28620
rect 9864 28577 9873 28611
rect 9873 28577 9907 28611
rect 9907 28577 9916 28611
rect 9864 28568 9916 28577
rect 9772 28500 9824 28552
rect 9680 28432 9732 28484
rect 11244 28611 11296 28620
rect 11244 28577 11253 28611
rect 11253 28577 11287 28611
rect 11287 28577 11296 28611
rect 11244 28568 11296 28577
rect 12072 28611 12124 28620
rect 12072 28577 12081 28611
rect 12081 28577 12115 28611
rect 12115 28577 12124 28611
rect 12072 28568 12124 28577
rect 12440 28568 12492 28620
rect 11888 28500 11940 28552
rect 12072 28432 12124 28484
rect 5908 28364 5960 28416
rect 6276 28364 6328 28416
rect 8576 28364 8628 28416
rect 9220 28364 9272 28416
rect 9956 28364 10008 28416
rect 10416 28364 10468 28416
rect 11336 28407 11388 28416
rect 11336 28373 11345 28407
rect 11345 28373 11379 28407
rect 11379 28373 11388 28407
rect 11336 28364 11388 28373
rect 11428 28364 11480 28416
rect 3662 28262 3714 28314
rect 3726 28262 3778 28314
rect 3790 28262 3842 28314
rect 3854 28262 3906 28314
rect 3918 28262 3970 28314
rect 10062 28262 10114 28314
rect 10126 28262 10178 28314
rect 10190 28262 10242 28314
rect 10254 28262 10306 28314
rect 10318 28262 10370 28314
rect 940 28160 992 28212
rect 2596 28203 2648 28212
rect 2596 28169 2605 28203
rect 2605 28169 2639 28203
rect 2639 28169 2648 28203
rect 2596 28160 2648 28169
rect 4436 28203 4488 28212
rect 4436 28169 4445 28203
rect 4445 28169 4479 28203
rect 4479 28169 4488 28203
rect 4436 28160 4488 28169
rect 6184 28203 6236 28212
rect 6184 28169 6193 28203
rect 6193 28169 6227 28203
rect 6227 28169 6236 28203
rect 6184 28160 6236 28169
rect 7840 28160 7892 28212
rect 7932 28203 7984 28212
rect 7932 28169 7941 28203
rect 7941 28169 7975 28203
rect 7975 28169 7984 28203
rect 7932 28160 7984 28169
rect 9036 28160 9088 28212
rect 9220 28203 9272 28212
rect 9220 28169 9229 28203
rect 9229 28169 9263 28203
rect 9263 28169 9272 28203
rect 9220 28160 9272 28169
rect 10600 28160 10652 28212
rect 11704 28160 11756 28212
rect 4160 28092 4212 28144
rect 2228 28067 2280 28076
rect 1400 27956 1452 28008
rect 2228 28033 2237 28067
rect 2237 28033 2271 28067
rect 2271 28033 2280 28067
rect 2228 28024 2280 28033
rect 3424 28024 3476 28076
rect 1952 27931 2004 27940
rect 1952 27897 1970 27931
rect 1970 27897 2004 27931
rect 3056 27999 3108 28008
rect 3056 27965 3065 27999
rect 3065 27965 3099 27999
rect 3099 27965 3108 27999
rect 3056 27956 3108 27965
rect 4160 27956 4212 28008
rect 4620 28024 4672 28076
rect 6644 28067 6696 28076
rect 6644 28033 6653 28067
rect 6653 28033 6687 28067
rect 6687 28033 6696 28067
rect 6644 28024 6696 28033
rect 6828 28092 6880 28144
rect 1952 27888 2004 27897
rect 3148 27888 3200 27940
rect 4068 27888 4120 27940
rect 3056 27820 3108 27872
rect 4436 27999 4488 28008
rect 4436 27965 4445 27999
rect 4445 27965 4479 27999
rect 4479 27965 4488 27999
rect 4436 27956 4488 27965
rect 5172 27956 5224 28008
rect 5540 27956 5592 28008
rect 5816 27956 5868 28008
rect 4344 27888 4396 27940
rect 5264 27888 5316 27940
rect 4620 27820 4672 27872
rect 5816 27863 5868 27872
rect 5816 27829 5825 27863
rect 5825 27829 5859 27863
rect 5859 27829 5868 27863
rect 5816 27820 5868 27829
rect 5908 27820 5960 27872
rect 7104 27956 7156 28008
rect 11152 28092 11204 28144
rect 7288 28024 7340 28076
rect 7840 28024 7892 28076
rect 8300 27956 8352 28008
rect 11428 28067 11480 28076
rect 11428 28033 11437 28067
rect 11437 28033 11471 28067
rect 11471 28033 11480 28067
rect 11428 28024 11480 28033
rect 7932 27888 7984 27940
rect 8024 27931 8076 27940
rect 8024 27897 8033 27931
rect 8033 27897 8067 27931
rect 8067 27897 8076 27931
rect 8024 27888 8076 27897
rect 8392 27931 8444 27940
rect 8392 27897 8401 27931
rect 8401 27897 8435 27931
rect 8435 27897 8444 27931
rect 8392 27888 8444 27897
rect 8576 27931 8628 27940
rect 8576 27897 8585 27931
rect 8585 27897 8619 27931
rect 8619 27897 8628 27931
rect 8576 27888 8628 27897
rect 9220 27956 9272 28008
rect 7196 27820 7248 27872
rect 7288 27863 7340 27872
rect 7288 27829 7297 27863
rect 7297 27829 7331 27863
rect 7331 27829 7340 27863
rect 7288 27820 7340 27829
rect 8760 27863 8812 27872
rect 8760 27829 8769 27863
rect 8769 27829 8803 27863
rect 8803 27829 8812 27863
rect 8760 27820 8812 27829
rect 9036 27820 9088 27872
rect 9864 27999 9916 28008
rect 9864 27965 9873 27999
rect 9873 27965 9907 27999
rect 9907 27965 9916 27999
rect 9864 27956 9916 27965
rect 10416 27999 10468 28008
rect 10416 27965 10425 27999
rect 10425 27965 10459 27999
rect 10459 27965 10468 27999
rect 10416 27956 10468 27965
rect 10508 27956 10560 28008
rect 11244 27956 11296 28008
rect 11336 27999 11388 28008
rect 11336 27965 11345 27999
rect 11345 27965 11379 27999
rect 11379 27965 11388 27999
rect 11336 27956 11388 27965
rect 11888 27999 11940 28008
rect 11888 27965 11897 27999
rect 11897 27965 11931 27999
rect 11931 27965 11940 27999
rect 11888 27956 11940 27965
rect 12072 27999 12124 28008
rect 12072 27965 12081 27999
rect 12081 27965 12115 27999
rect 12115 27965 12124 27999
rect 12072 27956 12124 27965
rect 9588 27820 9640 27872
rect 10600 27820 10652 27872
rect 11796 27820 11848 27872
rect 12256 27863 12308 27872
rect 12256 27829 12265 27863
rect 12265 27829 12299 27863
rect 12299 27829 12308 27863
rect 12256 27820 12308 27829
rect 4322 27718 4374 27770
rect 4386 27718 4438 27770
rect 4450 27718 4502 27770
rect 4514 27718 4566 27770
rect 4578 27718 4630 27770
rect 10722 27718 10774 27770
rect 10786 27718 10838 27770
rect 10850 27718 10902 27770
rect 10914 27718 10966 27770
rect 10978 27718 11030 27770
rect 2504 27616 2556 27668
rect 3424 27616 3476 27668
rect 4344 27616 4396 27668
rect 4804 27616 4856 27668
rect 5264 27616 5316 27668
rect 5724 27616 5776 27668
rect 6460 27616 6512 27668
rect 7012 27616 7064 27668
rect 1768 27523 1820 27532
rect 1768 27489 1777 27523
rect 1777 27489 1811 27523
rect 1811 27489 1820 27523
rect 1768 27480 1820 27489
rect 4160 27548 4212 27600
rect 8760 27616 8812 27668
rect 9312 27616 9364 27668
rect 8668 27548 8720 27600
rect 8944 27548 8996 27600
rect 2688 27480 2740 27532
rect 3056 27523 3108 27532
rect 3056 27489 3065 27523
rect 3065 27489 3099 27523
rect 3099 27489 3108 27523
rect 3056 27480 3108 27489
rect 3148 27523 3200 27532
rect 3148 27489 3157 27523
rect 3157 27489 3191 27523
rect 3191 27489 3200 27523
rect 3424 27523 3476 27532
rect 3148 27480 3200 27489
rect 3424 27489 3433 27523
rect 3433 27489 3467 27523
rect 3467 27489 3476 27523
rect 3424 27480 3476 27489
rect 4344 27523 4396 27532
rect 4344 27489 4353 27523
rect 4353 27489 4387 27523
rect 4387 27489 4396 27523
rect 4344 27480 4396 27489
rect 4896 27480 4948 27532
rect 5080 27523 5132 27532
rect 5080 27489 5089 27523
rect 5089 27489 5123 27523
rect 5123 27489 5132 27523
rect 5080 27480 5132 27489
rect 5172 27523 5224 27532
rect 5172 27489 5181 27523
rect 5181 27489 5215 27523
rect 5215 27489 5224 27523
rect 5172 27480 5224 27489
rect 5356 27523 5408 27532
rect 5356 27489 5365 27523
rect 5365 27489 5399 27523
rect 5399 27489 5408 27523
rect 5356 27480 5408 27489
rect 6092 27523 6144 27532
rect 6092 27489 6101 27523
rect 6101 27489 6135 27523
rect 6135 27489 6144 27523
rect 6092 27480 6144 27489
rect 6828 27523 6880 27532
rect 6828 27489 6837 27523
rect 6837 27489 6871 27523
rect 6871 27489 6880 27523
rect 6828 27480 6880 27489
rect 7012 27523 7064 27532
rect 7012 27489 7021 27523
rect 7021 27489 7055 27523
rect 7055 27489 7064 27523
rect 7012 27480 7064 27489
rect 7288 27480 7340 27532
rect 4620 27344 4672 27396
rect 4896 27387 4948 27396
rect 4896 27353 4905 27387
rect 4905 27353 4939 27387
rect 4939 27353 4948 27387
rect 4896 27344 4948 27353
rect 5448 27344 5500 27396
rect 7564 27455 7616 27464
rect 7564 27421 7573 27455
rect 7573 27421 7607 27455
rect 7607 27421 7616 27455
rect 7564 27412 7616 27421
rect 7748 27412 7800 27464
rect 8116 27480 8168 27532
rect 8208 27480 8260 27532
rect 9496 27616 9548 27668
rect 9588 27616 9640 27668
rect 10232 27616 10284 27668
rect 10600 27548 10652 27600
rect 9680 27523 9732 27532
rect 9680 27489 9689 27523
rect 9689 27489 9723 27523
rect 9723 27489 9732 27523
rect 11888 27616 11940 27668
rect 9680 27480 9732 27489
rect 9220 27412 9272 27464
rect 9312 27344 9364 27396
rect 10416 27344 10468 27396
rect 11152 27523 11204 27532
rect 11152 27489 11161 27523
rect 11161 27489 11195 27523
rect 11195 27489 11204 27523
rect 11152 27480 11204 27489
rect 11244 27480 11296 27532
rect 11704 27480 11756 27532
rect 11888 27523 11940 27532
rect 11888 27489 11897 27523
rect 11897 27489 11931 27523
rect 11931 27489 11940 27523
rect 11888 27480 11940 27489
rect 11060 27412 11112 27464
rect 11520 27455 11572 27464
rect 11520 27421 11529 27455
rect 11529 27421 11563 27455
rect 11563 27421 11572 27455
rect 11520 27412 11572 27421
rect 11612 27412 11664 27464
rect 1492 27276 1544 27328
rect 2044 27276 2096 27328
rect 4344 27276 4396 27328
rect 5172 27276 5224 27328
rect 6184 27319 6236 27328
rect 6184 27285 6193 27319
rect 6193 27285 6227 27319
rect 6227 27285 6236 27319
rect 6184 27276 6236 27285
rect 7012 27276 7064 27328
rect 7104 27276 7156 27328
rect 8576 27276 8628 27328
rect 11704 27319 11756 27328
rect 11704 27285 11713 27319
rect 11713 27285 11747 27319
rect 11747 27285 11756 27319
rect 11704 27276 11756 27285
rect 3662 27174 3714 27226
rect 3726 27174 3778 27226
rect 3790 27174 3842 27226
rect 3854 27174 3906 27226
rect 3918 27174 3970 27226
rect 10062 27174 10114 27226
rect 10126 27174 10178 27226
rect 10190 27174 10242 27226
rect 10254 27174 10306 27226
rect 10318 27174 10370 27226
rect 1768 27072 1820 27124
rect 2136 27072 2188 27124
rect 6092 27072 6144 27124
rect 7288 27072 7340 27124
rect 7564 27072 7616 27124
rect 7748 27115 7800 27124
rect 7748 27081 7757 27115
rect 7757 27081 7791 27115
rect 7791 27081 7800 27115
rect 7748 27072 7800 27081
rect 9128 27072 9180 27124
rect 10508 27072 10560 27124
rect 12072 27072 12124 27124
rect 664 27004 716 27056
rect 1676 27004 1728 27056
rect 4712 27004 4764 27056
rect 4988 27004 5040 27056
rect 6184 27004 6236 27056
rect 1860 26936 1912 26988
rect 4160 26979 4212 26988
rect 4160 26945 4169 26979
rect 4169 26945 4203 26979
rect 4203 26945 4212 26979
rect 4160 26936 4212 26945
rect 1492 26911 1544 26920
rect 1492 26877 1501 26911
rect 1501 26877 1535 26911
rect 1535 26877 1544 26911
rect 1492 26868 1544 26877
rect 480 26800 532 26852
rect 1308 26732 1360 26784
rect 4804 26868 4856 26920
rect 5632 26936 5684 26988
rect 6368 26936 6420 26988
rect 6000 26911 6052 26920
rect 6000 26877 6009 26911
rect 6009 26877 6043 26911
rect 6043 26877 6052 26911
rect 6000 26868 6052 26877
rect 6184 26911 6236 26920
rect 6184 26877 6193 26911
rect 6193 26877 6227 26911
rect 6227 26877 6236 26911
rect 6184 26868 6236 26877
rect 6828 27004 6880 27056
rect 7196 27004 7248 27056
rect 8944 27004 8996 27056
rect 7012 26936 7064 26988
rect 6828 26868 6880 26920
rect 7104 26911 7156 26920
rect 7104 26877 7113 26911
rect 7113 26877 7147 26911
rect 7147 26877 7156 26911
rect 7104 26868 7156 26877
rect 7380 26911 7432 26920
rect 7380 26877 7389 26911
rect 7389 26877 7423 26911
rect 7423 26877 7432 26911
rect 7380 26868 7432 26877
rect 7472 26911 7524 26920
rect 7472 26877 7481 26911
rect 7481 26877 7515 26911
rect 7515 26877 7524 26911
rect 7472 26868 7524 26877
rect 7748 26936 7800 26988
rect 8024 26868 8076 26920
rect 4804 26732 4856 26784
rect 5356 26732 5408 26784
rect 6368 26732 6420 26784
rect 6644 26732 6696 26784
rect 7564 26800 7616 26852
rect 8392 26911 8444 26920
rect 8392 26877 8401 26911
rect 8401 26877 8435 26911
rect 8435 26877 8444 26911
rect 8392 26868 8444 26877
rect 8668 26868 8720 26920
rect 8852 26868 8904 26920
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 9220 26868 9272 26920
rect 9772 26979 9824 26988
rect 9772 26945 9781 26979
rect 9781 26945 9815 26979
rect 9815 26945 9824 26979
rect 9772 26936 9824 26945
rect 8484 26800 8536 26852
rect 7932 26732 7984 26784
rect 9404 26732 9456 26784
rect 9772 26800 9824 26852
rect 11612 26936 11664 26988
rect 11704 26979 11756 26988
rect 11704 26945 11713 26979
rect 11713 26945 11747 26979
rect 11747 26945 11756 26979
rect 11704 26936 11756 26945
rect 11060 26911 11112 26920
rect 11060 26877 11069 26911
rect 11069 26877 11103 26911
rect 11103 26877 11112 26911
rect 11060 26868 11112 26877
rect 11152 26868 11204 26920
rect 10508 26800 10560 26852
rect 11796 26911 11848 26920
rect 11796 26877 11805 26911
rect 11805 26877 11839 26911
rect 11839 26877 11848 26911
rect 11796 26868 11848 26877
rect 12348 26800 12400 26852
rect 11336 26732 11388 26784
rect 4322 26630 4374 26682
rect 4386 26630 4438 26682
rect 4450 26630 4502 26682
rect 4514 26630 4566 26682
rect 4578 26630 4630 26682
rect 10722 26630 10774 26682
rect 10786 26630 10838 26682
rect 10850 26630 10902 26682
rect 10914 26630 10966 26682
rect 10978 26630 11030 26682
rect 1308 26528 1360 26580
rect 1400 26460 1452 26512
rect 1492 26392 1544 26444
rect 2136 26324 2188 26376
rect 2320 26460 2372 26512
rect 2504 26392 2556 26444
rect 2596 26435 2648 26444
rect 2596 26401 2605 26435
rect 2605 26401 2639 26435
rect 2639 26401 2648 26435
rect 2596 26392 2648 26401
rect 5816 26528 5868 26580
rect 6184 26528 6236 26580
rect 7380 26528 7432 26580
rect 8944 26571 8996 26580
rect 8944 26537 8953 26571
rect 8953 26537 8987 26571
rect 8987 26537 8996 26571
rect 8944 26528 8996 26537
rect 9220 26528 9272 26580
rect 2964 26503 3016 26512
rect 2964 26469 2973 26503
rect 2973 26469 3007 26503
rect 3007 26469 3016 26503
rect 2964 26460 3016 26469
rect 4160 26460 4212 26512
rect 4712 26392 4764 26444
rect 6644 26460 6696 26512
rect 10508 26528 10560 26580
rect 11888 26528 11940 26580
rect 2780 26299 2832 26308
rect 2780 26265 2789 26299
rect 2789 26265 2823 26299
rect 2823 26265 2832 26299
rect 2780 26256 2832 26265
rect 3240 26256 3292 26308
rect 3516 26256 3568 26308
rect 5356 26435 5408 26444
rect 5356 26401 5365 26435
rect 5365 26401 5399 26435
rect 5399 26401 5408 26435
rect 5356 26392 5408 26401
rect 5448 26367 5500 26376
rect 5448 26333 5457 26367
rect 5457 26333 5491 26367
rect 5491 26333 5500 26367
rect 5448 26324 5500 26333
rect 5540 26367 5592 26376
rect 5540 26333 5549 26367
rect 5549 26333 5583 26367
rect 5583 26333 5592 26367
rect 5540 26324 5592 26333
rect 6368 26392 6420 26444
rect 7104 26324 7156 26376
rect 7288 26324 7340 26376
rect 6368 26256 6420 26308
rect 1492 26188 1544 26240
rect 1860 26188 1912 26240
rect 2412 26188 2464 26240
rect 4252 26188 4304 26240
rect 4528 26231 4580 26240
rect 4528 26197 4537 26231
rect 4537 26197 4571 26231
rect 4571 26197 4580 26231
rect 4528 26188 4580 26197
rect 5080 26231 5132 26240
rect 5080 26197 5089 26231
rect 5089 26197 5123 26231
rect 5123 26197 5132 26231
rect 5080 26188 5132 26197
rect 6644 26188 6696 26240
rect 6828 26188 6880 26240
rect 7012 26188 7064 26240
rect 7288 26231 7340 26240
rect 7288 26197 7297 26231
rect 7297 26197 7331 26231
rect 7331 26197 7340 26231
rect 7288 26188 7340 26197
rect 7748 26392 7800 26444
rect 7932 26435 7984 26444
rect 7932 26401 7941 26435
rect 7941 26401 7975 26435
rect 7975 26401 7984 26435
rect 7932 26392 7984 26401
rect 8208 26435 8260 26444
rect 8208 26401 8217 26435
rect 8217 26401 8251 26435
rect 8251 26401 8260 26435
rect 8208 26392 8260 26401
rect 7656 26256 7708 26308
rect 7748 26256 7800 26308
rect 8300 26188 8352 26240
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 8760 26435 8812 26444
rect 8760 26401 8769 26435
rect 8769 26401 8803 26435
rect 8803 26401 8812 26435
rect 8760 26392 8812 26401
rect 9128 26392 9180 26444
rect 9404 26435 9456 26444
rect 9404 26401 9413 26435
rect 9413 26401 9447 26435
rect 9447 26401 9456 26435
rect 9404 26392 9456 26401
rect 8852 26324 8904 26376
rect 8944 26188 8996 26240
rect 3662 26086 3714 26138
rect 3726 26086 3778 26138
rect 3790 26086 3842 26138
rect 3854 26086 3906 26138
rect 3918 26086 3970 26138
rect 10062 26086 10114 26138
rect 10126 26086 10178 26138
rect 10190 26086 10242 26138
rect 10254 26086 10306 26138
rect 10318 26086 10370 26138
rect 2412 26027 2464 26036
rect 2412 25993 2421 26027
rect 2421 25993 2455 26027
rect 2455 25993 2464 26027
rect 2412 25984 2464 25993
rect 2596 26027 2648 26036
rect 2596 25993 2605 26027
rect 2605 25993 2639 26027
rect 2639 25993 2648 26027
rect 2596 25984 2648 25993
rect 4068 25984 4120 26036
rect 4988 25984 5040 26036
rect 5632 25984 5684 26036
rect 6000 25984 6052 26036
rect 6828 25984 6880 26036
rect 3148 25916 3200 25968
rect 1032 25891 1084 25900
rect 1032 25857 1041 25891
rect 1041 25857 1075 25891
rect 1075 25857 1084 25891
rect 1032 25848 1084 25857
rect 1492 25823 1544 25832
rect 1492 25789 1501 25823
rect 1501 25789 1535 25823
rect 1535 25789 1544 25823
rect 1492 25780 1544 25789
rect 1952 25848 2004 25900
rect 2596 25848 2648 25900
rect 2872 25780 2924 25832
rect 2964 25823 3016 25832
rect 2964 25789 2973 25823
rect 2973 25789 3007 25823
rect 3007 25789 3016 25823
rect 2964 25780 3016 25789
rect 3148 25780 3200 25832
rect 5540 25848 5592 25900
rect 7288 25916 7340 25968
rect 10416 25984 10468 26036
rect 9864 25848 9916 25900
rect 3424 25780 3476 25832
rect 3700 25823 3752 25832
rect 3700 25789 3709 25823
rect 3709 25789 3743 25823
rect 3743 25789 3752 25823
rect 3700 25780 3752 25789
rect 3976 25823 4028 25832
rect 3976 25789 3985 25823
rect 3985 25789 4019 25823
rect 4019 25789 4028 25823
rect 3976 25780 4028 25789
rect 4160 25823 4212 25832
rect 4160 25789 4169 25823
rect 4169 25789 4203 25823
rect 4203 25789 4212 25823
rect 4160 25780 4212 25789
rect 4252 25780 4304 25832
rect 4712 25780 4764 25832
rect 3516 25712 3568 25764
rect 5540 25712 5592 25764
rect 3424 25644 3476 25696
rect 5172 25644 5224 25696
rect 5448 25644 5500 25696
rect 6644 25823 6696 25832
rect 6644 25789 6683 25823
rect 6683 25789 6696 25823
rect 6644 25780 6696 25789
rect 5816 25644 5868 25696
rect 7104 25823 7156 25832
rect 7104 25789 7113 25823
rect 7113 25789 7147 25823
rect 7147 25789 7156 25823
rect 7104 25780 7156 25789
rect 8576 25823 8628 25832
rect 8576 25789 8585 25823
rect 8585 25789 8619 25823
rect 8619 25789 8628 25823
rect 8576 25780 8628 25789
rect 8852 25780 8904 25832
rect 9036 25780 9088 25832
rect 9404 25780 9456 25832
rect 7012 25712 7064 25764
rect 9128 25712 9180 25764
rect 9772 25712 9824 25764
rect 10508 25823 10560 25832
rect 10508 25789 10517 25823
rect 10517 25789 10551 25823
rect 10551 25789 10560 25823
rect 10508 25780 10560 25789
rect 10600 25712 10652 25764
rect 11060 25780 11112 25832
rect 11428 25712 11480 25764
rect 8300 25644 8352 25696
rect 8668 25644 8720 25696
rect 9588 25644 9640 25696
rect 10416 25644 10468 25696
rect 11244 25687 11296 25696
rect 11244 25653 11253 25687
rect 11253 25653 11287 25687
rect 11287 25653 11296 25687
rect 11244 25644 11296 25653
rect 12624 25780 12676 25832
rect 12072 25712 12124 25764
rect 11796 25644 11848 25696
rect 11980 25644 12032 25696
rect 12164 25687 12216 25696
rect 12164 25653 12173 25687
rect 12173 25653 12207 25687
rect 12207 25653 12216 25687
rect 12164 25644 12216 25653
rect 4322 25542 4374 25594
rect 4386 25542 4438 25594
rect 4450 25542 4502 25594
rect 4514 25542 4566 25594
rect 4578 25542 4630 25594
rect 10722 25542 10774 25594
rect 10786 25542 10838 25594
rect 10850 25542 10902 25594
rect 10914 25542 10966 25594
rect 10978 25542 11030 25594
rect 1676 25440 1728 25492
rect 1400 25372 1452 25424
rect 1952 25347 2004 25356
rect 1952 25313 1970 25347
rect 1970 25313 2004 25347
rect 1952 25304 2004 25313
rect 2596 25440 2648 25492
rect 3148 25483 3200 25492
rect 3148 25449 3157 25483
rect 3157 25449 3191 25483
rect 3191 25449 3200 25483
rect 3148 25440 3200 25449
rect 4068 25440 4120 25492
rect 7104 25440 7156 25492
rect 7932 25440 7984 25492
rect 8668 25440 8720 25492
rect 2504 25372 2556 25424
rect 5080 25372 5132 25424
rect 6828 25372 6880 25424
rect 10508 25440 10560 25492
rect 2412 25236 2464 25288
rect 3424 25304 3476 25356
rect 3516 25347 3568 25356
rect 3516 25313 3525 25347
rect 3525 25313 3559 25347
rect 3559 25313 3568 25347
rect 3516 25304 3568 25313
rect 4712 25304 4764 25356
rect 6368 25304 6420 25356
rect 7012 25347 7064 25356
rect 7012 25313 7021 25347
rect 7021 25313 7055 25347
rect 7055 25313 7064 25347
rect 7012 25304 7064 25313
rect 9588 25372 9640 25424
rect 10416 25415 10468 25424
rect 10416 25381 10425 25415
rect 10425 25381 10459 25415
rect 10459 25381 10468 25415
rect 10416 25372 10468 25381
rect 5080 25236 5132 25288
rect 5540 25236 5592 25288
rect 6828 25236 6880 25288
rect 7748 25304 7800 25356
rect 8208 25304 8260 25356
rect 8668 25304 8720 25356
rect 9956 25347 10008 25356
rect 9956 25313 9965 25347
rect 9965 25313 9999 25347
rect 9999 25313 10008 25347
rect 9956 25304 10008 25313
rect 10600 25304 10652 25356
rect 11612 25304 11664 25356
rect 12072 25304 12124 25356
rect 7380 25279 7432 25288
rect 7380 25245 7389 25279
rect 7389 25245 7423 25279
rect 7423 25245 7432 25279
rect 7380 25236 7432 25245
rect 7840 25279 7892 25288
rect 2872 25168 2924 25220
rect 3056 25168 3108 25220
rect 3148 25168 3200 25220
rect 3700 25168 3752 25220
rect 4620 25168 4672 25220
rect 4804 25168 4856 25220
rect 7012 25168 7064 25220
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 8484 25279 8536 25288
rect 8484 25245 8493 25279
rect 8493 25245 8527 25279
rect 8527 25245 8536 25279
rect 8484 25236 8536 25245
rect 9036 25168 9088 25220
rect 9496 25279 9548 25288
rect 9496 25245 9505 25279
rect 9505 25245 9539 25279
rect 9539 25245 9548 25279
rect 9496 25236 9548 25245
rect 9772 25236 9824 25288
rect 10508 25236 10560 25288
rect 11244 25279 11296 25288
rect 11244 25245 11253 25279
rect 11253 25245 11287 25279
rect 11287 25245 11296 25279
rect 11244 25236 11296 25245
rect 11704 25236 11756 25288
rect 12624 25236 12676 25288
rect 2320 25100 2372 25152
rect 2780 25100 2832 25152
rect 6552 25100 6604 25152
rect 7196 25100 7248 25152
rect 7564 25143 7616 25152
rect 7564 25109 7573 25143
rect 7573 25109 7607 25143
rect 7607 25109 7616 25143
rect 7564 25100 7616 25109
rect 8116 25100 8168 25152
rect 11520 25168 11572 25220
rect 3662 24998 3714 25050
rect 3726 24998 3778 25050
rect 3790 24998 3842 25050
rect 3854 24998 3906 25050
rect 3918 24998 3970 25050
rect 10062 24998 10114 25050
rect 10126 24998 10178 25050
rect 10190 24998 10242 25050
rect 10254 24998 10306 25050
rect 10318 24998 10370 25050
rect 3700 24896 3752 24948
rect 6552 24939 6604 24948
rect 6552 24905 6561 24939
rect 6561 24905 6595 24939
rect 6595 24905 6604 24939
rect 6552 24896 6604 24905
rect 6644 24896 6696 24948
rect 7380 24896 7432 24948
rect 7748 24896 7800 24948
rect 7840 24939 7892 24948
rect 7840 24905 7849 24939
rect 7849 24905 7883 24939
rect 7883 24905 7892 24939
rect 7840 24896 7892 24905
rect 8760 24896 8812 24948
rect 9496 24896 9548 24948
rect 9956 24896 10008 24948
rect 3884 24828 3936 24880
rect 4712 24828 4764 24880
rect 112 24760 164 24812
rect 664 24760 716 24812
rect 1308 24692 1360 24744
rect 1492 24735 1544 24744
rect 1492 24701 1501 24735
rect 1501 24701 1535 24735
rect 1535 24701 1544 24735
rect 1492 24692 1544 24701
rect 1032 24667 1084 24676
rect 1032 24633 1041 24667
rect 1041 24633 1075 24667
rect 1075 24633 1084 24667
rect 1032 24624 1084 24633
rect 1124 24624 1176 24676
rect 1768 24735 1820 24744
rect 1768 24701 1777 24735
rect 1777 24701 1811 24735
rect 1811 24701 1820 24735
rect 1768 24692 1820 24701
rect 2136 24735 2188 24744
rect 2136 24701 2145 24735
rect 2145 24701 2179 24735
rect 2179 24701 2188 24735
rect 2136 24692 2188 24701
rect 2320 24735 2372 24744
rect 2320 24701 2329 24735
rect 2329 24701 2363 24735
rect 2363 24701 2372 24735
rect 2320 24692 2372 24701
rect 2780 24692 2832 24744
rect 1860 24624 1912 24676
rect 3608 24692 3660 24744
rect 4252 24760 4304 24812
rect 4160 24692 4212 24744
rect 5724 24828 5776 24880
rect 5264 24692 5316 24744
rect 5816 24692 5868 24744
rect 6460 24735 6512 24744
rect 6460 24701 6469 24735
rect 6469 24701 6503 24735
rect 6503 24701 6512 24735
rect 6460 24692 6512 24701
rect 7012 24760 7064 24812
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 7840 24760 7892 24812
rect 4712 24624 4764 24676
rect 5080 24624 5132 24676
rect 6092 24624 6144 24676
rect 7656 24735 7708 24744
rect 7656 24701 7665 24735
rect 7665 24701 7699 24735
rect 7699 24701 7708 24735
rect 7656 24692 7708 24701
rect 7748 24692 7800 24744
rect 9220 24760 9272 24812
rect 9404 24760 9456 24812
rect 9864 24828 9916 24880
rect 10048 24828 10100 24880
rect 10324 24760 10376 24812
rect 10692 24803 10744 24812
rect 10692 24769 10701 24803
rect 10701 24769 10735 24803
rect 10735 24769 10744 24803
rect 10692 24760 10744 24769
rect 11704 24828 11756 24880
rect 11612 24760 11664 24812
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 7564 24624 7616 24676
rect 8576 24692 8628 24744
rect 9036 24735 9088 24744
rect 9036 24701 9045 24735
rect 9045 24701 9079 24735
rect 9079 24701 9088 24735
rect 9036 24692 9088 24701
rect 9128 24735 9180 24744
rect 9128 24701 9137 24735
rect 9137 24701 9171 24735
rect 9171 24701 9180 24735
rect 9128 24692 9180 24701
rect 9588 24692 9640 24744
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 9220 24624 9272 24676
rect 1492 24556 1544 24608
rect 3792 24556 3844 24608
rect 8024 24556 8076 24608
rect 8208 24556 8260 24608
rect 8944 24556 8996 24608
rect 9864 24556 9916 24608
rect 11336 24692 11388 24744
rect 11520 24692 11572 24744
rect 11980 24735 12032 24744
rect 11980 24701 11989 24735
rect 11989 24701 12023 24735
rect 12023 24701 12032 24735
rect 11980 24692 12032 24701
rect 12348 24692 12400 24744
rect 11704 24599 11756 24608
rect 11704 24565 11713 24599
rect 11713 24565 11747 24599
rect 11747 24565 11756 24599
rect 11704 24556 11756 24565
rect 4322 24454 4374 24506
rect 4386 24454 4438 24506
rect 4450 24454 4502 24506
rect 4514 24454 4566 24506
rect 4578 24454 4630 24506
rect 10722 24454 10774 24506
rect 10786 24454 10838 24506
rect 10850 24454 10902 24506
rect 10914 24454 10966 24506
rect 10978 24454 11030 24506
rect 756 24352 808 24404
rect 940 24352 992 24404
rect 1400 24284 1452 24336
rect 3516 24284 3568 24336
rect 4160 24352 4212 24404
rect 4620 24352 4672 24404
rect 5080 24352 5132 24404
rect 1492 24216 1544 24268
rect 1952 24216 2004 24268
rect 2780 24259 2832 24268
rect 2780 24225 2789 24259
rect 2789 24225 2823 24259
rect 2823 24225 2832 24259
rect 2780 24216 2832 24225
rect 3608 24216 3660 24268
rect 3700 24259 3752 24268
rect 3700 24225 3709 24259
rect 3709 24225 3743 24259
rect 3743 24225 3752 24259
rect 3700 24216 3752 24225
rect 3792 24259 3844 24268
rect 3792 24225 3801 24259
rect 3801 24225 3835 24259
rect 3835 24225 3844 24259
rect 3792 24216 3844 24225
rect 4068 24216 4120 24268
rect 4252 24216 4304 24268
rect 5356 24216 5408 24268
rect 5632 24216 5684 24268
rect 7012 24352 7064 24404
rect 7564 24395 7616 24404
rect 7564 24361 7573 24395
rect 7573 24361 7607 24395
rect 7607 24361 7616 24395
rect 7564 24352 7616 24361
rect 7656 24352 7708 24404
rect 7932 24352 7984 24404
rect 8484 24352 8536 24404
rect 9220 24395 9272 24404
rect 9220 24361 9229 24395
rect 9229 24361 9263 24395
rect 9263 24361 9272 24395
rect 9220 24352 9272 24361
rect 9404 24352 9456 24404
rect 11888 24352 11940 24404
rect 12440 24352 12492 24404
rect 3884 24080 3936 24132
rect 4160 24080 4212 24132
rect 4620 24123 4672 24132
rect 4620 24089 4629 24123
rect 4629 24089 4663 24123
rect 4663 24089 4672 24123
rect 4620 24080 4672 24089
rect 5724 24080 5776 24132
rect 6276 24259 6328 24268
rect 6276 24225 6285 24259
rect 6285 24225 6319 24259
rect 6319 24225 6328 24259
rect 6276 24216 6328 24225
rect 6460 24259 6512 24268
rect 6460 24225 6469 24259
rect 6469 24225 6503 24259
rect 6503 24225 6512 24259
rect 6460 24216 6512 24225
rect 6552 24259 6604 24268
rect 6552 24225 6561 24259
rect 6561 24225 6595 24259
rect 6595 24225 6604 24259
rect 6552 24216 6604 24225
rect 6644 24216 6696 24268
rect 6092 24148 6144 24200
rect 7288 24259 7340 24268
rect 7288 24225 7297 24259
rect 7297 24225 7331 24259
rect 7331 24225 7340 24259
rect 7288 24216 7340 24225
rect 7472 24216 7524 24268
rect 8024 24284 8076 24336
rect 7840 24259 7892 24268
rect 7840 24225 7849 24259
rect 7849 24225 7883 24259
rect 7883 24225 7892 24259
rect 7840 24216 7892 24225
rect 8208 24259 8260 24268
rect 8208 24225 8217 24259
rect 8217 24225 8251 24259
rect 8251 24225 8260 24259
rect 8208 24216 8260 24225
rect 7932 24191 7984 24200
rect 7932 24157 7941 24191
rect 7941 24157 7975 24191
rect 7975 24157 7984 24191
rect 7932 24148 7984 24157
rect 8024 24191 8076 24200
rect 8024 24157 8033 24191
rect 8033 24157 8067 24191
rect 8067 24157 8076 24191
rect 8576 24216 8628 24268
rect 9312 24259 9364 24268
rect 9312 24225 9321 24259
rect 9321 24225 9355 24259
rect 9355 24225 9364 24259
rect 9312 24216 9364 24225
rect 10600 24284 10652 24336
rect 9956 24216 10008 24268
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 11060 24216 11112 24268
rect 11244 24284 11296 24336
rect 11612 24259 11664 24268
rect 11612 24225 11621 24259
rect 11621 24225 11655 24259
rect 11655 24225 11664 24259
rect 11612 24216 11664 24225
rect 12072 24216 12124 24268
rect 8024 24148 8076 24157
rect 9588 24148 9640 24200
rect 7012 24080 7064 24132
rect 7472 24080 7524 24132
rect 9496 24080 9548 24132
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 10692 24080 10744 24132
rect 11980 24148 12032 24200
rect 2228 24055 2280 24064
rect 2228 24021 2237 24055
rect 2237 24021 2271 24055
rect 2271 24021 2280 24055
rect 2228 24012 2280 24021
rect 4068 24055 4120 24064
rect 4068 24021 4077 24055
rect 4077 24021 4111 24055
rect 4111 24021 4120 24055
rect 4068 24012 4120 24021
rect 4528 24012 4580 24064
rect 4896 24012 4948 24064
rect 5448 24012 5500 24064
rect 6092 24012 6144 24064
rect 6644 24012 6696 24064
rect 8300 24012 8352 24064
rect 9864 24055 9916 24064
rect 9864 24021 9873 24055
rect 9873 24021 9907 24055
rect 9907 24021 9916 24055
rect 9864 24012 9916 24021
rect 11428 24055 11480 24064
rect 11428 24021 11437 24055
rect 11437 24021 11471 24055
rect 11471 24021 11480 24055
rect 11428 24012 11480 24021
rect 11888 24012 11940 24064
rect 3662 23910 3714 23962
rect 3726 23910 3778 23962
rect 3790 23910 3842 23962
rect 3854 23910 3906 23962
rect 3918 23910 3970 23962
rect 10062 23910 10114 23962
rect 10126 23910 10178 23962
rect 10190 23910 10242 23962
rect 10254 23910 10306 23962
rect 10318 23910 10370 23962
rect 4344 23808 4396 23860
rect 5080 23808 5132 23860
rect 5632 23808 5684 23860
rect 6552 23808 6604 23860
rect 7564 23808 7616 23860
rect 8024 23808 8076 23860
rect 10508 23808 10560 23860
rect 11520 23808 11572 23860
rect 1032 23740 1084 23792
rect 1216 23740 1268 23792
rect 848 23672 900 23724
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 4252 23740 4304 23792
rect 4620 23740 4672 23792
rect 4896 23740 4948 23792
rect 3516 23672 3568 23724
rect 940 23604 992 23656
rect 1216 23604 1268 23656
rect 1308 23604 1360 23656
rect 1492 23604 1544 23656
rect 3056 23604 3108 23656
rect 3424 23604 3476 23656
rect 4804 23672 4856 23724
rect 4528 23647 4580 23656
rect 4528 23613 4537 23647
rect 4537 23613 4571 23647
rect 4571 23613 4580 23647
rect 4528 23604 4580 23613
rect 4620 23647 4672 23656
rect 4620 23613 4629 23647
rect 4629 23613 4663 23647
rect 4663 23613 4672 23647
rect 4620 23604 4672 23613
rect 5356 23740 5408 23792
rect 5540 23672 5592 23724
rect 4344 23579 4396 23588
rect 4344 23545 4353 23579
rect 4353 23545 4387 23579
rect 4387 23545 4396 23579
rect 4344 23536 4396 23545
rect 4988 23536 5040 23588
rect 5356 23647 5408 23656
rect 5356 23613 5365 23647
rect 5365 23613 5399 23647
rect 5399 23613 5408 23647
rect 5356 23604 5408 23613
rect 6092 23672 6144 23724
rect 6276 23672 6328 23724
rect 6644 23715 6696 23724
rect 6644 23681 6662 23715
rect 6662 23681 6696 23715
rect 6644 23672 6696 23681
rect 7196 23740 7248 23792
rect 7472 23740 7524 23792
rect 8208 23740 8260 23792
rect 10600 23740 10652 23792
rect 11796 23740 11848 23792
rect 11980 23851 12032 23860
rect 11980 23817 11989 23851
rect 11989 23817 12023 23851
rect 12023 23817 12032 23851
rect 11980 23808 12032 23817
rect 12164 23740 12216 23792
rect 12624 23740 12676 23792
rect 7104 23672 7156 23724
rect 7656 23647 7708 23656
rect 7656 23613 7665 23647
rect 7665 23613 7699 23647
rect 7699 23613 7708 23647
rect 7656 23604 7708 23613
rect 3424 23468 3476 23520
rect 4804 23468 4856 23520
rect 5632 23468 5684 23520
rect 11244 23672 11296 23724
rect 10324 23604 10376 23656
rect 10692 23604 10744 23656
rect 11336 23604 11388 23656
rect 11520 23536 11572 23588
rect 12164 23604 12216 23656
rect 11980 23536 12032 23588
rect 11060 23468 11112 23520
rect 12532 23536 12584 23588
rect 12164 23511 12216 23520
rect 12164 23477 12173 23511
rect 12173 23477 12207 23511
rect 12207 23477 12216 23511
rect 12164 23468 12216 23477
rect 4322 23366 4374 23418
rect 4386 23366 4438 23418
rect 4450 23366 4502 23418
rect 4514 23366 4566 23418
rect 4578 23366 4630 23418
rect 10722 23366 10774 23418
rect 10786 23366 10838 23418
rect 10850 23366 10902 23418
rect 10914 23366 10966 23418
rect 10978 23366 11030 23418
rect 388 23264 440 23316
rect 1492 23264 1544 23316
rect 1768 23264 1820 23316
rect 2780 23239 2832 23248
rect 2780 23205 2789 23239
rect 2789 23205 2823 23239
rect 2823 23205 2832 23239
rect 2780 23196 2832 23205
rect 3240 23196 3292 23248
rect 4436 23239 4488 23248
rect 4436 23205 4445 23239
rect 4445 23205 4479 23239
rect 4479 23205 4488 23239
rect 4436 23196 4488 23205
rect 940 23128 992 23180
rect 1124 23171 1176 23180
rect 1124 23137 1158 23171
rect 1158 23137 1176 23171
rect 1124 23128 1176 23137
rect 2320 23171 2372 23180
rect 2320 23137 2329 23171
rect 2329 23137 2363 23171
rect 2363 23137 2372 23171
rect 2320 23128 2372 23137
rect 2504 23128 2556 23180
rect 4252 23128 4304 23180
rect 5080 23264 5132 23316
rect 6092 23264 6144 23316
rect 5448 23239 5500 23248
rect 5448 23205 5457 23239
rect 5457 23205 5491 23239
rect 5491 23205 5500 23239
rect 5448 23196 5500 23205
rect 5080 23171 5132 23180
rect 5080 23137 5089 23171
rect 5089 23137 5123 23171
rect 5123 23137 5132 23171
rect 5080 23128 5132 23137
rect 5632 23128 5684 23180
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 5724 23060 5776 23112
rect 6092 23103 6144 23112
rect 6092 23069 6101 23103
rect 6101 23069 6135 23103
rect 6135 23069 6144 23103
rect 6092 23060 6144 23069
rect 7748 23264 7800 23316
rect 7932 23264 7984 23316
rect 6552 23196 6604 23248
rect 6828 23128 6880 23180
rect 6644 22992 6696 23044
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 7656 23171 7708 23180
rect 7656 23137 7665 23171
rect 7665 23137 7699 23171
rect 7699 23137 7708 23171
rect 7656 23128 7708 23137
rect 7932 23128 7984 23180
rect 9404 23264 9456 23316
rect 9036 23196 9088 23248
rect 8300 23171 8352 23180
rect 8300 23137 8309 23171
rect 8309 23137 8343 23171
rect 8343 23137 8352 23171
rect 8300 23128 8352 23137
rect 7104 22992 7156 23044
rect 7656 22992 7708 23044
rect 2412 22924 2464 22976
rect 2780 22924 2832 22976
rect 3516 22924 3568 22976
rect 5724 22924 5776 22976
rect 7012 22924 7064 22976
rect 8116 22992 8168 23044
rect 8576 22992 8628 23044
rect 9220 23128 9272 23180
rect 9404 23128 9456 23180
rect 11244 23264 11296 23316
rect 11428 23264 11480 23316
rect 11796 23264 11848 23316
rect 10324 23128 10376 23180
rect 9588 23103 9640 23112
rect 9588 23069 9597 23103
rect 9597 23069 9631 23103
rect 9631 23069 9640 23103
rect 9588 23060 9640 23069
rect 10692 23128 10744 23180
rect 10968 23128 11020 23180
rect 11244 23060 11296 23112
rect 11520 23171 11572 23180
rect 11520 23137 11529 23171
rect 11529 23137 11563 23171
rect 11563 23137 11572 23171
rect 11520 23128 11572 23137
rect 11796 23128 11848 23180
rect 12348 23128 12400 23180
rect 10508 22992 10560 23044
rect 7932 22924 7984 22976
rect 8300 22924 8352 22976
rect 8852 22924 8904 22976
rect 9680 22924 9732 22976
rect 10416 22924 10468 22976
rect 10600 22967 10652 22976
rect 10600 22933 10609 22967
rect 10609 22933 10643 22967
rect 10643 22933 10652 22967
rect 10600 22924 10652 22933
rect 11704 22924 11756 22976
rect 12348 22924 12400 22976
rect 3662 22822 3714 22874
rect 3726 22822 3778 22874
rect 3790 22822 3842 22874
rect 3854 22822 3906 22874
rect 3918 22822 3970 22874
rect 10062 22822 10114 22874
rect 10126 22822 10178 22874
rect 10190 22822 10242 22874
rect 10254 22822 10306 22874
rect 10318 22822 10370 22874
rect 2964 22720 3016 22772
rect 3700 22720 3752 22772
rect 4068 22720 4120 22772
rect 4160 22720 4212 22772
rect 1032 22695 1084 22704
rect 1032 22661 1041 22695
rect 1041 22661 1075 22695
rect 1075 22661 1084 22695
rect 1032 22652 1084 22661
rect 3148 22652 3200 22704
rect 1308 22627 1360 22636
rect 1308 22593 1317 22627
rect 1317 22593 1351 22627
rect 1351 22593 1360 22627
rect 1308 22584 1360 22593
rect 2228 22584 2280 22636
rect 2596 22584 2648 22636
rect 664 22516 716 22568
rect 1584 22516 1636 22568
rect 1952 22559 2004 22568
rect 1952 22525 1961 22559
rect 1961 22525 1995 22559
rect 1995 22525 2004 22559
rect 1952 22516 2004 22525
rect 2964 22559 3016 22568
rect 2964 22525 2973 22559
rect 2973 22525 3007 22559
rect 3007 22525 3016 22559
rect 2964 22516 3016 22525
rect 3148 22516 3200 22568
rect 4988 22652 5040 22704
rect 5356 22763 5408 22772
rect 5356 22729 5365 22763
rect 5365 22729 5399 22763
rect 5399 22729 5408 22763
rect 5356 22720 5408 22729
rect 6920 22763 6972 22772
rect 6920 22729 6929 22763
rect 6929 22729 6963 22763
rect 6963 22729 6972 22763
rect 6920 22720 6972 22729
rect 8852 22763 8904 22772
rect 8852 22729 8861 22763
rect 8861 22729 8895 22763
rect 8895 22729 8904 22763
rect 8852 22720 8904 22729
rect 9588 22720 9640 22772
rect 10968 22763 11020 22772
rect 10968 22729 10977 22763
rect 10977 22729 11011 22763
rect 11011 22729 11020 22763
rect 10968 22720 11020 22729
rect 11796 22720 11848 22772
rect 3516 22627 3568 22636
rect 3516 22593 3525 22627
rect 3525 22593 3559 22627
rect 3559 22593 3568 22627
rect 3516 22584 3568 22593
rect 4252 22584 4304 22636
rect 5264 22584 5316 22636
rect 6644 22652 6696 22704
rect 7564 22652 7616 22704
rect 5724 22627 5776 22636
rect 5724 22593 5733 22627
rect 5733 22593 5767 22627
rect 5767 22593 5776 22627
rect 5724 22584 5776 22593
rect 1032 22380 1084 22432
rect 4068 22380 4120 22432
rect 4620 22448 4672 22500
rect 6368 22559 6420 22568
rect 6368 22525 6377 22559
rect 6377 22525 6411 22559
rect 6411 22525 6420 22559
rect 6368 22516 6420 22525
rect 6736 22516 6788 22568
rect 8208 22559 8260 22568
rect 8208 22525 8217 22559
rect 8217 22525 8251 22559
rect 8251 22525 8260 22559
rect 8208 22516 8260 22525
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 8852 22516 8904 22568
rect 9036 22559 9088 22568
rect 9036 22525 9045 22559
rect 9045 22525 9079 22559
rect 9079 22525 9088 22559
rect 9036 22516 9088 22525
rect 10600 22652 10652 22704
rect 10140 22584 10192 22636
rect 10876 22584 10928 22636
rect 9220 22516 9272 22568
rect 9588 22516 9640 22568
rect 9956 22516 10008 22568
rect 6828 22448 6880 22500
rect 8116 22448 8168 22500
rect 4988 22423 5040 22432
rect 4988 22389 4997 22423
rect 4997 22389 5031 22423
rect 5031 22389 5040 22423
rect 4988 22380 5040 22389
rect 6920 22380 6972 22432
rect 8208 22380 8260 22432
rect 9128 22380 9180 22432
rect 9404 22423 9456 22432
rect 9404 22389 9413 22423
rect 9413 22389 9447 22423
rect 9447 22389 9456 22423
rect 9404 22380 9456 22389
rect 9588 22380 9640 22432
rect 10784 22516 10836 22568
rect 12348 22652 12400 22704
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 12348 22516 12400 22568
rect 11244 22491 11296 22500
rect 11244 22457 11253 22491
rect 11253 22457 11287 22491
rect 11287 22457 11296 22491
rect 11244 22448 11296 22457
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 11888 22380 11940 22432
rect 12164 22491 12216 22500
rect 12164 22457 12173 22491
rect 12173 22457 12207 22491
rect 12207 22457 12216 22491
rect 12164 22448 12216 22457
rect 12440 22380 12492 22432
rect 4322 22278 4374 22330
rect 4386 22278 4438 22330
rect 4450 22278 4502 22330
rect 4514 22278 4566 22330
rect 4578 22278 4630 22330
rect 10722 22278 10774 22330
rect 10786 22278 10838 22330
rect 10850 22278 10902 22330
rect 10914 22278 10966 22330
rect 10978 22278 11030 22330
rect 3148 22176 3200 22228
rect 8668 22176 8720 22228
rect 9864 22176 9916 22228
rect 9956 22176 10008 22228
rect 3240 22151 3292 22160
rect 3240 22117 3249 22151
rect 3249 22117 3283 22151
rect 3283 22117 3292 22151
rect 3240 22108 3292 22117
rect 2412 22040 2464 22092
rect 3700 22083 3752 22092
rect 3700 22049 3709 22083
rect 3709 22049 3743 22083
rect 3743 22049 3752 22083
rect 3700 22040 3752 22049
rect 2688 21972 2740 22024
rect 4068 22083 4120 22092
rect 4068 22049 4077 22083
rect 4077 22049 4111 22083
rect 4111 22049 4120 22083
rect 4068 22040 4120 22049
rect 4252 22083 4304 22092
rect 4252 22049 4261 22083
rect 4261 22049 4295 22083
rect 4295 22049 4304 22083
rect 4252 22040 4304 22049
rect 4896 22083 4948 22092
rect 4896 22049 4905 22083
rect 4905 22049 4939 22083
rect 4939 22049 4948 22083
rect 4896 22040 4948 22049
rect 5724 22108 5776 22160
rect 5816 22040 5868 22092
rect 6736 22040 6788 22092
rect 848 21904 900 21956
rect 1400 21904 1452 21956
rect 2964 21904 3016 21956
rect 5724 21972 5776 22024
rect 664 21836 716 21888
rect 1124 21836 1176 21888
rect 1676 21836 1728 21888
rect 2228 21836 2280 21888
rect 3240 21836 3292 21888
rect 4160 21836 4212 21888
rect 4896 21836 4948 21888
rect 5724 21836 5776 21888
rect 6184 21904 6236 21956
rect 6644 21836 6696 21888
rect 6736 21836 6788 21888
rect 7196 22015 7248 22024
rect 7196 21981 7205 22015
rect 7205 21981 7239 22015
rect 7239 21981 7248 22015
rect 7196 21972 7248 21981
rect 7564 21972 7616 22024
rect 7748 21972 7800 22024
rect 8116 22083 8168 22092
rect 8116 22049 8125 22083
rect 8125 22049 8159 22083
rect 8159 22049 8168 22083
rect 8116 22040 8168 22049
rect 8300 22040 8352 22092
rect 8484 22083 8536 22092
rect 8484 22049 8493 22083
rect 8493 22049 8527 22083
rect 8527 22049 8536 22083
rect 8484 22040 8536 22049
rect 8944 22083 8996 22092
rect 8944 22049 8953 22083
rect 8953 22049 8987 22083
rect 8987 22049 8996 22083
rect 8944 22040 8996 22049
rect 9404 22108 9456 22160
rect 10416 22108 10468 22160
rect 10600 22176 10652 22228
rect 11520 22219 11572 22228
rect 11520 22185 11529 22219
rect 11529 22185 11563 22219
rect 11563 22185 11572 22219
rect 11520 22176 11572 22185
rect 11888 22176 11940 22228
rect 12440 22176 12492 22228
rect 9128 22083 9180 22090
rect 9128 22049 9142 22083
rect 9142 22049 9176 22083
rect 9176 22049 9180 22083
rect 9128 22038 9180 22049
rect 7472 21904 7524 21956
rect 9220 21972 9272 22024
rect 9956 22083 10008 22092
rect 9956 22049 9965 22083
rect 9965 22049 9999 22083
rect 9999 22049 10008 22083
rect 9956 22040 10008 22049
rect 7380 21836 7432 21888
rect 8116 21836 8168 21888
rect 10048 21836 10100 21888
rect 10508 22083 10560 22092
rect 10508 22049 10517 22083
rect 10517 22049 10551 22083
rect 10551 22049 10560 22083
rect 10508 22040 10560 22049
rect 10692 22040 10744 22092
rect 11428 22083 11480 22092
rect 11428 22049 11437 22083
rect 11437 22049 11471 22083
rect 11471 22049 11480 22083
rect 11428 22040 11480 22049
rect 12164 22108 12216 22160
rect 11336 21972 11388 22024
rect 10600 21904 10652 21956
rect 11152 21904 11204 21956
rect 11704 21904 11756 21956
rect 10508 21836 10560 21888
rect 10968 21879 11020 21888
rect 10968 21845 10977 21879
rect 10977 21845 11011 21879
rect 11011 21845 11020 21879
rect 10968 21836 11020 21845
rect 3662 21734 3714 21786
rect 3726 21734 3778 21786
rect 3790 21734 3842 21786
rect 3854 21734 3906 21786
rect 3918 21734 3970 21786
rect 10062 21734 10114 21786
rect 10126 21734 10178 21786
rect 10190 21734 10242 21786
rect 10254 21734 10306 21786
rect 10318 21734 10370 21786
rect 1492 21632 1544 21684
rect 2780 21607 2832 21616
rect 2780 21573 2789 21607
rect 2789 21573 2823 21607
rect 2823 21573 2832 21607
rect 3424 21632 3476 21684
rect 2780 21564 2832 21573
rect 1216 21496 1268 21548
rect 1308 21428 1360 21480
rect 2228 21428 2280 21480
rect 2504 21428 2556 21480
rect 2964 21496 3016 21548
rect 4160 21564 4212 21616
rect 3516 21496 3568 21548
rect 5264 21632 5316 21684
rect 5816 21675 5868 21684
rect 5816 21641 5825 21675
rect 5825 21641 5859 21675
rect 5859 21641 5868 21675
rect 5816 21632 5868 21641
rect 8208 21632 8260 21684
rect 8392 21675 8444 21684
rect 8392 21641 8401 21675
rect 8401 21641 8435 21675
rect 8435 21641 8444 21675
rect 8392 21632 8444 21641
rect 5632 21496 5684 21548
rect 6552 21607 6604 21616
rect 6552 21573 6561 21607
rect 6561 21573 6595 21607
rect 6595 21573 6604 21607
rect 6552 21564 6604 21573
rect 7012 21564 7064 21616
rect 7104 21564 7156 21616
rect 3608 21471 3660 21480
rect 3608 21437 3617 21471
rect 3617 21437 3651 21471
rect 3651 21437 3660 21471
rect 3608 21428 3660 21437
rect 3792 21471 3844 21480
rect 3792 21437 3801 21471
rect 3801 21437 3835 21471
rect 3835 21437 3844 21471
rect 3792 21428 3844 21437
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 4252 21471 4304 21480
rect 4252 21437 4261 21471
rect 4261 21437 4295 21471
rect 4295 21437 4304 21471
rect 4252 21428 4304 21437
rect 4344 21428 4396 21480
rect 3884 21360 3936 21412
rect 1400 21292 1452 21344
rect 2320 21292 2372 21344
rect 2964 21292 3016 21344
rect 4896 21428 4948 21480
rect 5724 21428 5776 21480
rect 6828 21496 6880 21548
rect 6644 21428 6696 21480
rect 6920 21428 6972 21480
rect 7380 21539 7432 21548
rect 7380 21505 7389 21539
rect 7389 21505 7423 21539
rect 7423 21505 7432 21539
rect 7380 21496 7432 21505
rect 9588 21564 9640 21616
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 8760 21496 8812 21548
rect 5356 21403 5408 21412
rect 5356 21369 5365 21403
rect 5365 21369 5399 21403
rect 5399 21369 5408 21403
rect 5356 21360 5408 21369
rect 5540 21403 5592 21412
rect 5540 21369 5565 21403
rect 5565 21369 5592 21403
rect 5540 21360 5592 21369
rect 6000 21335 6052 21344
rect 6000 21301 6009 21335
rect 6009 21301 6043 21335
rect 6043 21301 6052 21335
rect 6000 21292 6052 21301
rect 6276 21335 6328 21344
rect 6276 21301 6285 21335
rect 6285 21301 6319 21335
rect 6319 21301 6328 21335
rect 6276 21292 6328 21301
rect 7380 21360 7432 21412
rect 8668 21471 8720 21480
rect 8668 21437 8677 21471
rect 8677 21437 8711 21471
rect 8711 21437 8720 21471
rect 8668 21428 8720 21437
rect 8484 21360 8536 21412
rect 9588 21428 9640 21480
rect 9680 21471 9732 21480
rect 9680 21437 9689 21471
rect 9689 21437 9723 21471
rect 9723 21437 9732 21471
rect 9680 21428 9732 21437
rect 10600 21632 10652 21684
rect 10876 21632 10928 21684
rect 11520 21632 11572 21684
rect 9956 21607 10008 21616
rect 9956 21573 9965 21607
rect 9965 21573 9999 21607
rect 9999 21573 10008 21607
rect 9956 21564 10008 21573
rect 10048 21607 10100 21616
rect 10048 21573 10057 21607
rect 10057 21573 10091 21607
rect 10091 21573 10100 21607
rect 10048 21564 10100 21573
rect 10508 21496 10560 21548
rect 10416 21428 10468 21480
rect 12716 21496 12768 21548
rect 9864 21360 9916 21412
rect 10508 21360 10560 21412
rect 12348 21428 12400 21480
rect 9036 21292 9088 21344
rect 10968 21292 11020 21344
rect 11704 21335 11756 21344
rect 11704 21301 11713 21335
rect 11713 21301 11747 21335
rect 11747 21301 11756 21335
rect 11704 21292 11756 21301
rect 4322 21190 4374 21242
rect 4386 21190 4438 21242
rect 4450 21190 4502 21242
rect 4514 21190 4566 21242
rect 4578 21190 4630 21242
rect 10722 21190 10774 21242
rect 10786 21190 10838 21242
rect 10850 21190 10902 21242
rect 10914 21190 10966 21242
rect 10978 21190 11030 21242
rect 2412 21131 2464 21140
rect 2412 21097 2421 21131
rect 2421 21097 2455 21131
rect 2455 21097 2464 21131
rect 2412 21088 2464 21097
rect 3056 21088 3108 21140
rect 3700 21088 3752 21140
rect 4896 21088 4948 21140
rect 4988 21088 5040 21140
rect 6736 21088 6788 21140
rect 7196 21088 7248 21140
rect 1492 20952 1544 21004
rect 2320 20952 2372 21004
rect 3792 21020 3844 21072
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 3516 20952 3568 21004
rect 3608 20952 3660 21004
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 3056 20884 3108 20936
rect 3792 20884 3844 20936
rect 4252 20995 4304 21004
rect 4252 20961 4261 20995
rect 4261 20961 4295 20995
rect 4295 20961 4304 20995
rect 4252 20952 4304 20961
rect 6276 21020 6328 21072
rect 8944 21088 8996 21140
rect 9956 21088 10008 21140
rect 9772 21020 9824 21072
rect 10048 21020 10100 21072
rect 4620 20995 4672 21004
rect 4620 20961 4629 20995
rect 4629 20961 4663 20995
rect 4663 20961 4672 20995
rect 4620 20952 4672 20961
rect 4896 20952 4948 21004
rect 4528 20927 4580 20936
rect 4528 20893 4537 20927
rect 4537 20893 4571 20927
rect 4571 20893 4580 20927
rect 4528 20884 4580 20893
rect 4988 20884 5040 20936
rect 5356 20884 5408 20936
rect 5816 20995 5868 21004
rect 5816 20961 5825 20995
rect 5825 20961 5859 20995
rect 5859 20961 5868 20995
rect 5816 20952 5868 20961
rect 6644 20952 6696 21004
rect 7196 20952 7248 21004
rect 7380 20995 7432 21004
rect 7380 20961 7389 20995
rect 7389 20961 7423 20995
rect 7423 20961 7432 20995
rect 7380 20952 7432 20961
rect 7472 20995 7524 21004
rect 7472 20961 7481 20995
rect 7481 20961 7515 20995
rect 7515 20961 7524 20995
rect 7472 20952 7524 20961
rect 8392 20952 8444 21004
rect 10508 20952 10560 21004
rect 11152 20952 11204 21004
rect 6276 20884 6328 20936
rect 6828 20884 6880 20936
rect 7104 20927 7156 20936
rect 7104 20893 7113 20927
rect 7113 20893 7147 20927
rect 7147 20893 7156 20927
rect 7104 20884 7156 20893
rect 7656 20884 7708 20936
rect 7748 20927 7800 20936
rect 7748 20893 7757 20927
rect 7757 20893 7791 20927
rect 7791 20893 7800 20927
rect 7748 20884 7800 20893
rect 1216 20748 1268 20800
rect 2504 20748 2556 20800
rect 3516 20791 3568 20800
rect 3516 20757 3525 20791
rect 3525 20757 3559 20791
rect 3559 20757 3568 20791
rect 3516 20748 3568 20757
rect 4252 20748 4304 20800
rect 8392 20816 8444 20868
rect 11336 20995 11388 21004
rect 11336 20961 11345 20995
rect 11345 20961 11379 20995
rect 11379 20961 11388 20995
rect 11336 20952 11388 20961
rect 11520 20952 11572 21004
rect 11612 20995 11664 21004
rect 11612 20961 11621 20995
rect 11621 20961 11655 20995
rect 11655 20961 11664 20995
rect 11612 20952 11664 20961
rect 12072 20952 12124 21004
rect 11428 20816 11480 20868
rect 6368 20748 6420 20800
rect 6920 20791 6972 20800
rect 6920 20757 6929 20791
rect 6929 20757 6963 20791
rect 6963 20757 6972 20791
rect 6920 20748 6972 20757
rect 8208 20748 8260 20800
rect 11060 20748 11112 20800
rect 3662 20646 3714 20698
rect 3726 20646 3778 20698
rect 3790 20646 3842 20698
rect 3854 20646 3906 20698
rect 3918 20646 3970 20698
rect 10062 20646 10114 20698
rect 10126 20646 10178 20698
rect 10190 20646 10242 20698
rect 10254 20646 10306 20698
rect 10318 20646 10370 20698
rect 664 20544 716 20596
rect 3700 20544 3752 20596
rect 3792 20544 3844 20596
rect 4620 20544 4672 20596
rect 5632 20587 5684 20596
rect 5632 20553 5641 20587
rect 5641 20553 5675 20587
rect 5675 20553 5684 20587
rect 5632 20544 5684 20553
rect 5724 20544 5776 20596
rect 6644 20544 6696 20596
rect 7196 20544 7248 20596
rect 7564 20544 7616 20596
rect 7748 20544 7800 20596
rect 7932 20587 7984 20596
rect 7932 20553 7941 20587
rect 7941 20553 7975 20587
rect 7975 20553 7984 20587
rect 7932 20544 7984 20553
rect 8760 20587 8812 20596
rect 8760 20553 8769 20587
rect 8769 20553 8803 20587
rect 8803 20553 8812 20587
rect 8760 20544 8812 20553
rect 20 20476 72 20528
rect 756 20408 808 20460
rect 1216 20408 1268 20460
rect 2688 20519 2740 20528
rect 2688 20485 2697 20519
rect 2697 20485 2731 20519
rect 2731 20485 2740 20519
rect 2688 20476 2740 20485
rect 3424 20476 3476 20528
rect 3976 20476 4028 20528
rect 3240 20408 3292 20460
rect 4068 20408 4120 20460
rect 1400 20340 1452 20392
rect 1492 20383 1544 20392
rect 1492 20349 1501 20383
rect 1501 20349 1535 20383
rect 1535 20349 1544 20383
rect 1492 20340 1544 20349
rect 1768 20340 1820 20392
rect 2412 20340 2464 20392
rect 3148 20340 3200 20392
rect 4252 20383 4304 20392
rect 4252 20349 4261 20383
rect 4261 20349 4295 20383
rect 4295 20349 4304 20383
rect 4252 20340 4304 20349
rect 5356 20476 5408 20528
rect 6920 20476 6972 20528
rect 9496 20544 9548 20596
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 1584 20204 1636 20256
rect 3608 20272 3660 20324
rect 3700 20272 3752 20324
rect 4160 20272 4212 20324
rect 3332 20204 3384 20256
rect 3976 20204 4028 20256
rect 4620 20204 4672 20256
rect 7012 20408 7064 20460
rect 5816 20383 5868 20392
rect 5816 20349 5825 20383
rect 5825 20349 5859 20383
rect 5859 20349 5868 20383
rect 5816 20340 5868 20349
rect 6276 20340 6328 20392
rect 6644 20383 6696 20392
rect 6644 20349 6653 20383
rect 6653 20349 6687 20383
rect 6687 20349 6696 20383
rect 6644 20340 6696 20349
rect 6828 20340 6880 20392
rect 9312 20476 9364 20528
rect 9864 20587 9916 20596
rect 9864 20553 9873 20587
rect 9873 20553 9907 20587
rect 9907 20553 9916 20587
rect 9864 20544 9916 20553
rect 11152 20544 11204 20596
rect 6920 20272 6972 20324
rect 7932 20408 7984 20460
rect 8300 20408 8352 20460
rect 8852 20408 8904 20460
rect 7288 20340 7340 20392
rect 7196 20204 7248 20256
rect 7564 20340 7616 20392
rect 8024 20340 8076 20392
rect 8392 20383 8444 20392
rect 8392 20349 8401 20383
rect 8401 20349 8435 20383
rect 8435 20349 8444 20383
rect 8392 20340 8444 20349
rect 8484 20340 8536 20392
rect 8116 20272 8168 20324
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 8760 20340 8812 20392
rect 9128 20383 9180 20392
rect 9128 20349 9138 20383
rect 9138 20349 9172 20383
rect 9172 20349 9180 20383
rect 9588 20408 9640 20460
rect 9128 20340 9180 20349
rect 10508 20340 10560 20392
rect 11980 20340 12032 20392
rect 12348 20340 12400 20392
rect 8484 20247 8536 20256
rect 8484 20213 8493 20247
rect 8493 20213 8527 20247
rect 8527 20213 8536 20247
rect 8484 20204 8536 20213
rect 9404 20315 9456 20324
rect 9404 20281 9413 20315
rect 9413 20281 9447 20315
rect 9447 20281 9456 20315
rect 9404 20272 9456 20281
rect 10416 20272 10468 20324
rect 10692 20272 10744 20324
rect 9220 20204 9272 20256
rect 9864 20204 9916 20256
rect 4322 20102 4374 20154
rect 4386 20102 4438 20154
rect 4450 20102 4502 20154
rect 4514 20102 4566 20154
rect 4578 20102 4630 20154
rect 10722 20102 10774 20154
rect 10786 20102 10838 20154
rect 10850 20102 10902 20154
rect 10914 20102 10966 20154
rect 10978 20102 11030 20154
rect 940 20043 992 20052
rect 940 20009 949 20043
rect 949 20009 983 20043
rect 983 20009 992 20043
rect 940 20000 992 20009
rect 1676 20000 1728 20052
rect 2688 20043 2740 20052
rect 2688 20009 2697 20043
rect 2697 20009 2731 20043
rect 2731 20009 2740 20043
rect 2688 20000 2740 20009
rect 2412 19932 2464 19984
rect 1676 19864 1728 19916
rect 3516 20000 3568 20052
rect 3976 20000 4028 20052
rect 4160 20000 4212 20052
rect 5632 20000 5684 20052
rect 6368 20000 6420 20052
rect 664 19796 716 19848
rect 2044 19796 2096 19848
rect 2504 19796 2556 19848
rect 3516 19907 3568 19916
rect 3516 19873 3525 19907
rect 3525 19873 3559 19907
rect 3559 19873 3568 19907
rect 3516 19864 3568 19873
rect 3608 19907 3660 19916
rect 3608 19873 3617 19907
rect 3617 19873 3651 19907
rect 3651 19873 3660 19907
rect 3608 19864 3660 19873
rect 3884 19907 3936 19916
rect 3884 19873 3893 19907
rect 3893 19873 3927 19907
rect 3927 19873 3936 19907
rect 3884 19864 3936 19873
rect 4068 19864 4120 19916
rect 4160 19907 4212 19916
rect 4160 19873 4169 19907
rect 4169 19873 4203 19907
rect 4203 19873 4212 19907
rect 4160 19864 4212 19873
rect 4436 19907 4488 19916
rect 4436 19873 4445 19907
rect 4445 19873 4479 19907
rect 4479 19873 4488 19907
rect 4436 19864 4488 19873
rect 4528 19864 4580 19916
rect 3056 19771 3108 19780
rect 3056 19737 3065 19771
rect 3065 19737 3099 19771
rect 3099 19737 3108 19771
rect 3056 19728 3108 19737
rect 3148 19728 3200 19780
rect 3976 19728 4028 19780
rect 1308 19660 1360 19712
rect 1676 19660 1728 19712
rect 2504 19703 2556 19712
rect 2504 19669 2513 19703
rect 2513 19669 2547 19703
rect 2547 19669 2556 19703
rect 2504 19660 2556 19669
rect 2872 19660 2924 19712
rect 3792 19660 3844 19712
rect 4160 19660 4212 19712
rect 4620 19660 4672 19712
rect 4896 19864 4948 19916
rect 5448 19864 5500 19916
rect 6276 19932 6328 19984
rect 5632 19864 5684 19916
rect 7104 20000 7156 20052
rect 7472 20000 7524 20052
rect 8208 20000 8260 20052
rect 8576 20000 8628 20052
rect 6920 19864 6972 19916
rect 8484 19932 8536 19984
rect 10600 20000 10652 20052
rect 10968 20000 11020 20052
rect 11336 20043 11388 20052
rect 11336 20009 11345 20043
rect 11345 20009 11379 20043
rect 11379 20009 11388 20043
rect 11336 20000 11388 20009
rect 5724 19796 5776 19848
rect 5724 19660 5776 19712
rect 6276 19796 6328 19848
rect 7288 19796 7340 19848
rect 6460 19728 6512 19780
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 8300 19864 8352 19916
rect 8852 19932 8904 19984
rect 9128 19864 9180 19916
rect 8760 19839 8812 19848
rect 8760 19805 8769 19839
rect 8769 19805 8803 19839
rect 8803 19805 8812 19839
rect 8760 19796 8812 19805
rect 9036 19796 9088 19848
rect 9312 19907 9364 19916
rect 9312 19873 9321 19907
rect 9321 19873 9355 19907
rect 9355 19873 9364 19907
rect 9312 19864 9364 19873
rect 10876 19932 10928 19984
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 11060 19864 11112 19916
rect 11152 19907 11204 19916
rect 11152 19873 11161 19907
rect 11161 19873 11195 19907
rect 11195 19873 11204 19907
rect 11152 19864 11204 19873
rect 11428 19907 11480 19916
rect 11428 19873 11437 19907
rect 11437 19873 11471 19907
rect 11471 19873 11480 19907
rect 11428 19864 11480 19873
rect 11888 19975 11940 19984
rect 11888 19941 11897 19975
rect 11897 19941 11931 19975
rect 11931 19941 11940 19975
rect 11888 19932 11940 19941
rect 12164 19864 12216 19916
rect 7748 19728 7800 19780
rect 8300 19771 8352 19780
rect 8300 19737 8309 19771
rect 8309 19737 8343 19771
rect 8343 19737 8352 19771
rect 8300 19728 8352 19737
rect 8668 19728 8720 19780
rect 9312 19728 9364 19780
rect 11888 19796 11940 19848
rect 10600 19728 10652 19780
rect 6828 19660 6880 19712
rect 8208 19660 8260 19712
rect 9036 19660 9088 19712
rect 10416 19660 10468 19712
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 10968 19703 11020 19712
rect 10968 19669 10977 19703
rect 10977 19669 11011 19703
rect 11011 19669 11020 19703
rect 10968 19660 11020 19669
rect 11060 19660 11112 19712
rect 11888 19660 11940 19712
rect 3662 19558 3714 19610
rect 3726 19558 3778 19610
rect 3790 19558 3842 19610
rect 3854 19558 3906 19610
rect 3918 19558 3970 19610
rect 10062 19558 10114 19610
rect 10126 19558 10178 19610
rect 10190 19558 10242 19610
rect 10254 19558 10306 19610
rect 10318 19558 10370 19610
rect 1492 19456 1544 19508
rect 3240 19456 3292 19508
rect 4436 19456 4488 19508
rect 5172 19456 5224 19508
rect 6644 19456 6696 19508
rect 7932 19456 7984 19508
rect 1952 19388 2004 19440
rect 2872 19388 2924 19440
rect 4804 19388 4856 19440
rect 5448 19388 5500 19440
rect 7840 19388 7892 19440
rect 8392 19388 8444 19440
rect 1492 19320 1544 19372
rect 3332 19320 3384 19372
rect 3700 19320 3752 19372
rect 4712 19320 4764 19372
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 8760 19456 8812 19508
rect 8852 19456 8904 19508
rect 9772 19456 9824 19508
rect 10048 19456 10100 19508
rect 10416 19456 10468 19508
rect 11796 19499 11848 19508
rect 11796 19465 11805 19499
rect 11805 19465 11839 19499
rect 11839 19465 11848 19499
rect 11796 19456 11848 19465
rect 1584 19295 1636 19304
rect 1584 19261 1593 19295
rect 1593 19261 1627 19295
rect 1627 19261 1636 19295
rect 1584 19252 1636 19261
rect 1952 19252 2004 19304
rect 2964 19252 3016 19304
rect 5540 19295 5592 19304
rect 5540 19261 5549 19295
rect 5549 19261 5583 19295
rect 5583 19261 5592 19295
rect 5540 19252 5592 19261
rect 5632 19252 5684 19304
rect 2320 19159 2372 19168
rect 2320 19125 2329 19159
rect 2329 19125 2363 19159
rect 2363 19125 2372 19159
rect 2320 19116 2372 19125
rect 2504 19227 2556 19236
rect 2504 19193 2513 19227
rect 2513 19193 2547 19227
rect 2547 19193 2556 19227
rect 2504 19184 2556 19193
rect 3056 19184 3108 19236
rect 3516 19184 3568 19236
rect 4988 19116 5040 19168
rect 6460 19295 6512 19304
rect 6460 19261 6469 19295
rect 6469 19261 6503 19295
rect 6503 19261 6512 19295
rect 6460 19252 6512 19261
rect 6552 19295 6604 19304
rect 6552 19261 6586 19295
rect 6586 19261 6604 19295
rect 6552 19252 6604 19261
rect 6736 19295 6788 19304
rect 6736 19261 6745 19295
rect 6745 19261 6779 19295
rect 6779 19261 6788 19295
rect 6736 19252 6788 19261
rect 7656 19295 7708 19304
rect 7656 19261 7665 19295
rect 7665 19261 7699 19295
rect 7699 19261 7708 19295
rect 7656 19252 7708 19261
rect 7932 19295 7984 19304
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 8116 19295 8168 19304
rect 8116 19261 8125 19295
rect 8125 19261 8159 19295
rect 8159 19261 8168 19295
rect 8116 19252 8168 19261
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 9588 19320 9640 19372
rect 9956 19320 10008 19372
rect 8300 19252 8352 19304
rect 8576 19295 8628 19304
rect 8576 19261 8585 19295
rect 8585 19261 8619 19295
rect 8619 19261 8628 19295
rect 8576 19252 8628 19261
rect 6644 19116 6696 19168
rect 7196 19116 7248 19168
rect 8668 19116 8720 19168
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 9128 19184 9180 19236
rect 9772 19252 9824 19304
rect 10508 19295 10560 19304
rect 10508 19261 10517 19295
rect 10517 19261 10551 19295
rect 10551 19261 10560 19295
rect 10508 19252 10560 19261
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 11244 19252 11296 19304
rect 11704 19295 11756 19304
rect 11704 19261 11713 19295
rect 11713 19261 11747 19295
rect 11747 19261 11756 19295
rect 11704 19252 11756 19261
rect 11980 19295 12032 19304
rect 11980 19261 11989 19295
rect 11989 19261 12023 19295
rect 12023 19261 12032 19295
rect 11980 19252 12032 19261
rect 12256 19252 12308 19304
rect 9588 19184 9640 19236
rect 11060 19184 11112 19236
rect 11612 19116 11664 19168
rect 12256 19116 12308 19168
rect 4322 19014 4374 19066
rect 4386 19014 4438 19066
rect 4450 19014 4502 19066
rect 4514 19014 4566 19066
rect 4578 19014 4630 19066
rect 10722 19014 10774 19066
rect 10786 19014 10838 19066
rect 10850 19014 10902 19066
rect 10914 19014 10966 19066
rect 10978 19014 11030 19066
rect 2136 18912 2188 18964
rect 2780 18912 2832 18964
rect 2964 18912 3016 18964
rect 1768 18844 1820 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 1584 18819 1636 18828
rect 1584 18785 1593 18819
rect 1593 18785 1627 18819
rect 1627 18785 1636 18819
rect 1584 18776 1636 18785
rect 2320 18776 2372 18828
rect 3516 18844 3568 18896
rect 3056 18819 3108 18828
rect 3056 18785 3065 18819
rect 3065 18785 3099 18819
rect 3099 18785 3108 18819
rect 3056 18776 3108 18785
rect 3148 18819 3200 18828
rect 3148 18785 3157 18819
rect 3157 18785 3191 18819
rect 3191 18785 3200 18819
rect 3148 18776 3200 18785
rect 940 18751 992 18760
rect 940 18717 949 18751
rect 949 18717 983 18751
rect 983 18717 992 18751
rect 940 18708 992 18717
rect 1952 18708 2004 18760
rect 2136 18708 2188 18760
rect 4528 18776 4580 18828
rect 4620 18819 4672 18828
rect 4620 18785 4629 18819
rect 4629 18785 4663 18819
rect 4663 18785 4672 18819
rect 4620 18776 4672 18785
rect 3700 18708 3752 18760
rect 4344 18708 4396 18760
rect 3792 18640 3844 18692
rect 5080 18708 5132 18760
rect 4988 18640 5040 18692
rect 2412 18615 2464 18624
rect 2412 18581 2421 18615
rect 2421 18581 2455 18615
rect 2455 18581 2464 18615
rect 2412 18572 2464 18581
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 3608 18572 3660 18624
rect 5448 18887 5500 18896
rect 5448 18853 5457 18887
rect 5457 18853 5491 18887
rect 5491 18853 5500 18887
rect 5448 18844 5500 18853
rect 5632 18819 5684 18828
rect 5632 18785 5641 18819
rect 5641 18785 5675 18819
rect 5675 18785 5684 18819
rect 5632 18776 5684 18785
rect 6552 18912 6604 18964
rect 7012 18912 7064 18964
rect 8116 18912 8168 18964
rect 8944 18912 8996 18964
rect 8668 18844 8720 18896
rect 9496 18912 9548 18964
rect 9588 18955 9640 18964
rect 9588 18921 9597 18955
rect 9597 18921 9631 18955
rect 9631 18921 9640 18955
rect 9588 18912 9640 18921
rect 9772 18955 9824 18964
rect 9772 18921 9781 18955
rect 9781 18921 9815 18955
rect 9815 18921 9824 18955
rect 9772 18912 9824 18921
rect 9864 18912 9916 18964
rect 9128 18844 9180 18896
rect 9312 18844 9364 18896
rect 9404 18844 9456 18896
rect 12164 18955 12216 18964
rect 12164 18921 12173 18955
rect 12173 18921 12207 18955
rect 12207 18921 12216 18955
rect 12164 18912 12216 18921
rect 6828 18819 6880 18828
rect 6828 18785 6862 18819
rect 6862 18785 6880 18819
rect 6828 18776 6880 18785
rect 7012 18819 7064 18828
rect 7012 18785 7021 18819
rect 7021 18785 7055 18819
rect 7055 18785 7064 18819
rect 7012 18776 7064 18785
rect 5540 18708 5592 18760
rect 6184 18708 6236 18760
rect 6092 18640 6144 18692
rect 7564 18572 7616 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 8208 18776 8260 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 9404 18708 9456 18760
rect 9864 18776 9916 18828
rect 10048 18776 10100 18828
rect 10416 18776 10468 18828
rect 10600 18819 10652 18828
rect 10600 18785 10609 18819
rect 10609 18785 10643 18819
rect 10643 18785 10652 18819
rect 10600 18776 10652 18785
rect 11612 18819 11664 18828
rect 11612 18785 11621 18819
rect 11621 18785 11655 18819
rect 11655 18785 11664 18819
rect 11612 18776 11664 18785
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 11060 18708 11112 18760
rect 11980 18751 12032 18760
rect 11980 18717 11989 18751
rect 11989 18717 12023 18751
rect 12023 18717 12032 18751
rect 11980 18708 12032 18717
rect 9036 18572 9088 18624
rect 9680 18640 9732 18692
rect 11612 18572 11664 18624
rect 3662 18470 3714 18522
rect 3726 18470 3778 18522
rect 3790 18470 3842 18522
rect 3854 18470 3906 18522
rect 3918 18470 3970 18522
rect 10062 18470 10114 18522
rect 10126 18470 10178 18522
rect 10190 18470 10242 18522
rect 10254 18470 10306 18522
rect 10318 18470 10370 18522
rect 1584 18368 1636 18420
rect 2412 18368 2464 18420
rect 5816 18368 5868 18420
rect 6184 18368 6236 18420
rect 8300 18368 8352 18420
rect 8392 18411 8444 18420
rect 8392 18377 8401 18411
rect 8401 18377 8435 18411
rect 8435 18377 8444 18411
rect 8392 18368 8444 18377
rect 10416 18411 10468 18420
rect 10416 18377 10425 18411
rect 10425 18377 10459 18411
rect 10459 18377 10468 18411
rect 10416 18368 10468 18377
rect 12072 18368 12124 18420
rect 2596 18300 2648 18352
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2320 18164 2372 18216
rect 1308 18096 1360 18148
rect 1584 18096 1636 18148
rect 2136 18096 2188 18148
rect 2872 18164 2924 18216
rect 3056 18232 3108 18284
rect 3056 18096 3108 18148
rect 3608 18275 3660 18284
rect 3608 18241 3617 18275
rect 3617 18241 3651 18275
rect 3651 18241 3660 18275
rect 3608 18232 3660 18241
rect 4252 18300 4304 18352
rect 4804 18300 4856 18352
rect 5356 18300 5408 18352
rect 9220 18300 9272 18352
rect 9772 18300 9824 18352
rect 2780 18028 2832 18080
rect 3700 18164 3752 18216
rect 4068 18232 4120 18284
rect 4252 18207 4304 18216
rect 4252 18173 4261 18207
rect 4261 18173 4295 18207
rect 4295 18173 4304 18207
rect 4252 18164 4304 18173
rect 7932 18232 7984 18284
rect 8024 18232 8076 18284
rect 5816 18164 5868 18216
rect 7656 18207 7708 18216
rect 7656 18173 7665 18207
rect 7665 18173 7699 18207
rect 7699 18173 7708 18207
rect 7656 18164 7708 18173
rect 7748 18164 7800 18216
rect 8668 18207 8720 18216
rect 8668 18173 8677 18207
rect 8677 18173 8711 18207
rect 8711 18173 8720 18207
rect 8668 18164 8720 18173
rect 8944 18164 8996 18216
rect 9220 18164 9272 18216
rect 9404 18207 9456 18216
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 10416 18164 10468 18216
rect 10508 18207 10560 18216
rect 10508 18173 10517 18207
rect 10517 18173 10551 18207
rect 10551 18173 10560 18207
rect 10508 18164 10560 18173
rect 11060 18232 11112 18284
rect 3516 18096 3568 18148
rect 3332 18028 3384 18080
rect 4620 18096 4672 18148
rect 5632 18096 5684 18148
rect 7104 18096 7156 18148
rect 7196 18139 7248 18148
rect 7196 18105 7205 18139
rect 7205 18105 7239 18139
rect 7239 18105 7248 18139
rect 7196 18096 7248 18105
rect 7380 18139 7432 18148
rect 7380 18105 7389 18139
rect 7389 18105 7423 18139
rect 7423 18105 7432 18139
rect 7380 18096 7432 18105
rect 9128 18139 9180 18148
rect 9128 18105 9137 18139
rect 9137 18105 9171 18139
rect 9171 18105 9180 18139
rect 9128 18096 9180 18105
rect 11796 18300 11848 18352
rect 12256 18232 12308 18284
rect 11704 18207 11756 18216
rect 11704 18173 11713 18207
rect 11713 18173 11747 18207
rect 11747 18173 11756 18207
rect 11704 18164 11756 18173
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 4068 18071 4120 18080
rect 4068 18037 4077 18071
rect 4077 18037 4111 18071
rect 4111 18037 4120 18071
rect 4068 18028 4120 18037
rect 4252 18028 4304 18080
rect 4528 18028 4580 18080
rect 4804 18028 4856 18080
rect 4988 18028 5040 18080
rect 6460 18028 6512 18080
rect 6920 18071 6972 18080
rect 6920 18037 6929 18071
rect 6929 18037 6963 18071
rect 6963 18037 6972 18071
rect 6920 18028 6972 18037
rect 7012 18028 7064 18080
rect 8024 18071 8076 18080
rect 8024 18037 8033 18071
rect 8033 18037 8067 18071
rect 8067 18037 8076 18071
rect 8024 18028 8076 18037
rect 8392 18028 8444 18080
rect 12440 18096 12492 18148
rect 11520 18028 11572 18080
rect 4322 17926 4374 17978
rect 4386 17926 4438 17978
rect 4450 17926 4502 17978
rect 4514 17926 4566 17978
rect 4578 17926 4630 17978
rect 10722 17926 10774 17978
rect 10786 17926 10838 17978
rect 10850 17926 10902 17978
rect 10914 17926 10966 17978
rect 10978 17926 11030 17978
rect 3148 17824 3200 17876
rect 3240 17824 3292 17876
rect 3424 17824 3476 17876
rect 2320 17756 2372 17808
rect 3332 17756 3384 17808
rect 3700 17824 3752 17876
rect 3884 17824 3936 17876
rect 4252 17824 4304 17876
rect 4436 17824 4488 17876
rect 6276 17824 6328 17876
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 2228 17620 2280 17629
rect 1308 17484 1360 17536
rect 2596 17688 2648 17740
rect 2872 17688 2924 17740
rect 4068 17756 4120 17808
rect 5264 17756 5316 17808
rect 5448 17756 5500 17808
rect 5724 17756 5776 17808
rect 4252 17731 4304 17740
rect 4252 17697 4261 17731
rect 4261 17697 4295 17731
rect 4295 17697 4304 17731
rect 4252 17688 4304 17697
rect 4804 17688 4856 17740
rect 3332 17663 3384 17672
rect 3332 17629 3341 17663
rect 3341 17629 3375 17663
rect 3375 17629 3384 17663
rect 3332 17620 3384 17629
rect 3884 17620 3936 17672
rect 6000 17731 6052 17740
rect 6000 17697 6009 17731
rect 6009 17697 6043 17731
rect 6043 17697 6052 17731
rect 6000 17688 6052 17697
rect 6552 17756 6604 17808
rect 7748 17824 7800 17876
rect 7932 17824 7984 17876
rect 6460 17688 6512 17740
rect 7012 17799 7064 17808
rect 7012 17765 7021 17799
rect 7021 17765 7055 17799
rect 7055 17765 7064 17799
rect 7012 17756 7064 17765
rect 7564 17756 7616 17808
rect 6092 17663 6144 17672
rect 6092 17629 6101 17663
rect 6101 17629 6135 17663
rect 6135 17629 6144 17663
rect 6092 17620 6144 17629
rect 6276 17620 6328 17672
rect 7748 17688 7800 17740
rect 8392 17756 8444 17808
rect 8760 17756 8812 17808
rect 8208 17731 8260 17740
rect 8208 17697 8217 17731
rect 8217 17697 8251 17731
rect 8251 17697 8260 17731
rect 8208 17688 8260 17697
rect 8576 17688 8628 17740
rect 9036 17824 9088 17876
rect 9128 17824 9180 17876
rect 9864 17824 9916 17876
rect 10140 17824 10192 17876
rect 10600 17824 10652 17876
rect 11520 17824 11572 17876
rect 9772 17756 9824 17808
rect 9128 17731 9180 17740
rect 9128 17697 9135 17731
rect 9135 17697 9180 17731
rect 2596 17484 2648 17536
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 3240 17484 3292 17536
rect 3976 17552 4028 17604
rect 4252 17552 4304 17604
rect 5448 17552 5500 17604
rect 5540 17552 5592 17604
rect 7380 17552 7432 17604
rect 7656 17552 7708 17604
rect 7840 17552 7892 17604
rect 8392 17620 8444 17672
rect 9128 17688 9180 17697
rect 9404 17731 9456 17740
rect 9404 17697 9418 17731
rect 9418 17697 9452 17731
rect 9452 17697 9456 17731
rect 9404 17688 9456 17697
rect 9588 17688 9640 17740
rect 10140 17731 10192 17740
rect 10140 17697 10149 17731
rect 10149 17697 10183 17731
rect 10183 17697 10192 17731
rect 10140 17688 10192 17697
rect 11336 17731 11388 17740
rect 11336 17697 11345 17731
rect 11345 17697 11379 17731
rect 11379 17697 11388 17731
rect 11336 17688 11388 17697
rect 12532 17688 12584 17740
rect 10416 17620 10468 17672
rect 11428 17663 11480 17672
rect 11428 17629 11437 17663
rect 11437 17629 11471 17663
rect 11471 17629 11480 17663
rect 11428 17620 11480 17629
rect 10600 17552 10652 17604
rect 4528 17527 4580 17536
rect 4528 17493 4537 17527
rect 4537 17493 4571 17527
rect 4571 17493 4580 17527
rect 4528 17484 4580 17493
rect 4804 17484 4856 17536
rect 5172 17484 5224 17536
rect 7104 17484 7156 17536
rect 8760 17484 8812 17536
rect 9220 17484 9272 17536
rect 9772 17484 9824 17536
rect 10508 17484 10560 17536
rect 3662 17382 3714 17434
rect 3726 17382 3778 17434
rect 3790 17382 3842 17434
rect 3854 17382 3906 17434
rect 3918 17382 3970 17434
rect 10062 17382 10114 17434
rect 10126 17382 10178 17434
rect 10190 17382 10242 17434
rect 10254 17382 10306 17434
rect 10318 17382 10370 17434
rect 2688 17280 2740 17332
rect 3332 17280 3384 17332
rect 5264 17323 5316 17332
rect 5264 17289 5273 17323
rect 5273 17289 5307 17323
rect 5307 17289 5316 17323
rect 5264 17280 5316 17289
rect 1584 17212 1636 17264
rect 2320 17212 2372 17264
rect 2596 17255 2648 17264
rect 2596 17221 2605 17255
rect 2605 17221 2639 17255
rect 2639 17221 2648 17255
rect 2596 17212 2648 17221
rect 3884 17212 3936 17264
rect 4436 17212 4488 17264
rect 4988 17212 5040 17264
rect 2136 17144 2188 17196
rect 1308 17119 1360 17128
rect 1308 17085 1317 17119
rect 1317 17085 1351 17119
rect 1351 17085 1360 17119
rect 1308 17076 1360 17085
rect 1400 17076 1452 17128
rect 1952 17051 2004 17060
rect 1952 17017 1961 17051
rect 1961 17017 1995 17051
rect 1995 17017 2004 17051
rect 1952 17008 2004 17017
rect 3148 17076 3200 17128
rect 4528 17144 4580 17196
rect 4804 17076 4856 17128
rect 4988 17119 5040 17128
rect 4988 17085 4997 17119
rect 4997 17085 5031 17119
rect 5031 17085 5040 17119
rect 4988 17076 5040 17085
rect 6276 17280 6328 17332
rect 6460 17280 6512 17332
rect 6644 17280 6696 17332
rect 7012 17280 7064 17332
rect 7564 17280 7616 17332
rect 7840 17280 7892 17332
rect 5540 17076 5592 17128
rect 5724 17076 5776 17128
rect 5908 17076 5960 17128
rect 7196 17144 7248 17196
rect 7748 17144 7800 17196
rect 2136 17008 2188 17060
rect 2412 17008 2464 17060
rect 3240 17008 3292 17060
rect 3332 16940 3384 16992
rect 4804 16983 4856 16992
rect 4804 16949 4813 16983
rect 4813 16949 4847 16983
rect 4847 16949 4856 16983
rect 4804 16940 4856 16949
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 6552 17076 6604 17128
rect 6552 16940 6604 16992
rect 6644 16940 6696 16992
rect 7380 17076 7432 17128
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 7196 17008 7248 17060
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 9128 17280 9180 17332
rect 10600 17280 10652 17332
rect 11060 17280 11112 17332
rect 9680 17212 9732 17264
rect 10416 17255 10468 17264
rect 10416 17221 10425 17255
rect 10425 17221 10459 17255
rect 10459 17221 10468 17255
rect 10416 17212 10468 17221
rect 11428 17212 11480 17264
rect 8852 17076 8904 17128
rect 9680 17076 9732 17128
rect 9772 17119 9824 17128
rect 9772 17085 9781 17119
rect 9781 17085 9815 17119
rect 9815 17085 9824 17119
rect 10140 17144 10192 17196
rect 9772 17076 9824 17085
rect 10232 17076 10284 17128
rect 11060 17144 11112 17196
rect 7472 16983 7524 16992
rect 7472 16949 7481 16983
rect 7481 16949 7515 16983
rect 7515 16949 7524 16983
rect 7472 16940 7524 16949
rect 7656 16940 7708 16992
rect 11244 17008 11296 17060
rect 11428 17119 11480 17128
rect 11428 17085 11437 17119
rect 11437 17085 11471 17119
rect 11471 17085 11480 17119
rect 11428 17076 11480 17085
rect 12164 17008 12216 17060
rect 8852 16940 8904 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 10048 16940 10100 16992
rect 10324 16940 10376 16992
rect 10416 16940 10468 16992
rect 4322 16838 4374 16890
rect 4386 16838 4438 16890
rect 4450 16838 4502 16890
rect 4514 16838 4566 16890
rect 4578 16838 4630 16890
rect 10722 16838 10774 16890
rect 10786 16838 10838 16890
rect 10850 16838 10902 16890
rect 10914 16838 10966 16890
rect 10978 16838 11030 16890
rect 1768 16736 1820 16788
rect 2412 16736 2464 16788
rect 2504 16736 2556 16788
rect 2780 16736 2832 16788
rect 4068 16736 4120 16788
rect 940 16711 992 16720
rect 940 16677 949 16711
rect 949 16677 983 16711
rect 983 16677 992 16711
rect 940 16668 992 16677
rect 3884 16668 3936 16720
rect 4712 16736 4764 16788
rect 1216 16600 1268 16652
rect 1768 16600 1820 16652
rect 4804 16668 4856 16720
rect 4988 16711 5040 16720
rect 4988 16677 4997 16711
rect 4997 16677 5031 16711
rect 5031 16677 5040 16711
rect 4988 16668 5040 16677
rect 2136 16532 2188 16584
rect 5080 16600 5132 16652
rect 5816 16736 5868 16788
rect 5632 16711 5684 16720
rect 5632 16677 5641 16711
rect 5641 16677 5675 16711
rect 5675 16677 5684 16711
rect 5632 16668 5684 16677
rect 6460 16668 6512 16720
rect 7840 16736 7892 16788
rect 7932 16736 7984 16788
rect 9588 16736 9640 16788
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 10232 16779 10284 16788
rect 10232 16745 10241 16779
rect 10241 16745 10275 16779
rect 10275 16745 10284 16779
rect 10232 16736 10284 16745
rect 4436 16575 4488 16584
rect 4436 16541 4445 16575
rect 4445 16541 4479 16575
rect 4479 16541 4488 16575
rect 4436 16532 4488 16541
rect 5908 16532 5960 16584
rect 5080 16464 5132 16516
rect 5724 16464 5776 16516
rect 6368 16600 6420 16652
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 6828 16643 6880 16652
rect 6828 16609 6837 16643
rect 6837 16609 6871 16643
rect 6871 16609 6880 16643
rect 6828 16600 6880 16609
rect 7288 16643 7340 16652
rect 7288 16609 7297 16643
rect 7297 16609 7331 16643
rect 7331 16609 7340 16643
rect 7288 16600 7340 16609
rect 10140 16668 10192 16720
rect 11336 16779 11388 16788
rect 11336 16745 11345 16779
rect 11345 16745 11379 16779
rect 11379 16745 11388 16779
rect 11336 16736 11388 16745
rect 7748 16600 7800 16652
rect 8024 16600 8076 16652
rect 8300 16643 8352 16652
rect 8300 16609 8309 16643
rect 8309 16609 8343 16643
rect 8343 16609 8352 16643
rect 8300 16600 8352 16609
rect 8576 16643 8628 16652
rect 8576 16609 8585 16643
rect 8585 16609 8619 16643
rect 8619 16609 8628 16643
rect 8576 16600 8628 16609
rect 8668 16600 8720 16652
rect 7012 16532 7064 16584
rect 8392 16532 8444 16584
rect 8944 16643 8996 16652
rect 8944 16609 8953 16643
rect 8953 16609 8987 16643
rect 8987 16609 8996 16643
rect 8944 16600 8996 16609
rect 9036 16643 9088 16652
rect 9036 16609 9045 16643
rect 9045 16609 9079 16643
rect 9079 16609 9088 16643
rect 9036 16600 9088 16609
rect 9588 16600 9640 16652
rect 9680 16600 9732 16652
rect 5264 16396 5316 16448
rect 6092 16439 6144 16448
rect 6092 16405 6101 16439
rect 6101 16405 6135 16439
rect 6135 16405 6144 16439
rect 6092 16396 6144 16405
rect 6644 16464 6696 16516
rect 7196 16464 7248 16516
rect 7288 16464 7340 16516
rect 7380 16464 7432 16516
rect 9404 16532 9456 16584
rect 9772 16532 9824 16584
rect 11244 16643 11296 16652
rect 11244 16609 11253 16643
rect 11253 16609 11287 16643
rect 11287 16609 11296 16643
rect 11244 16600 11296 16609
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 11888 16600 11940 16652
rect 11980 16643 12032 16652
rect 11980 16609 11989 16643
rect 11989 16609 12023 16643
rect 12023 16609 12032 16643
rect 11980 16600 12032 16609
rect 12072 16643 12124 16652
rect 12072 16609 12081 16643
rect 12081 16609 12115 16643
rect 12115 16609 12124 16643
rect 12072 16600 12124 16609
rect 12164 16532 12216 16584
rect 10048 16507 10100 16516
rect 10048 16473 10057 16507
rect 10057 16473 10091 16507
rect 10091 16473 10100 16507
rect 10048 16464 10100 16473
rect 7656 16396 7708 16448
rect 9588 16396 9640 16448
rect 9772 16396 9824 16448
rect 10140 16396 10192 16448
rect 10232 16396 10284 16448
rect 12348 16464 12400 16516
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 3662 16294 3714 16346
rect 3726 16294 3778 16346
rect 3790 16294 3842 16346
rect 3854 16294 3906 16346
rect 3918 16294 3970 16346
rect 10062 16294 10114 16346
rect 10126 16294 10178 16346
rect 10190 16294 10242 16346
rect 10254 16294 10306 16346
rect 10318 16294 10370 16346
rect 1584 16192 1636 16244
rect 1952 16192 2004 16244
rect 2136 16192 2188 16244
rect 2780 16235 2832 16244
rect 2780 16201 2789 16235
rect 2789 16201 2823 16235
rect 2823 16201 2832 16235
rect 2780 16192 2832 16201
rect 6828 16192 6880 16244
rect 8208 16192 8260 16244
rect 6552 16124 6604 16176
rect 9680 16192 9732 16244
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 12072 16192 12124 16244
rect 8668 16124 8720 16176
rect 10324 16124 10376 16176
rect 2688 16056 2740 16108
rect 2228 15988 2280 16040
rect 2504 15988 2556 16040
rect 1768 15920 1820 15972
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 5080 16056 5132 16108
rect 5908 16056 5960 16108
rect 5816 16031 5868 16040
rect 5816 15997 5825 16031
rect 5825 15997 5859 16031
rect 5859 15997 5868 16031
rect 5816 15988 5868 15997
rect 6276 15988 6328 16040
rect 7748 16056 7800 16108
rect 8300 16056 8352 16108
rect 6920 15988 6972 16040
rect 7012 16031 7064 16040
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7104 16031 7156 16040
rect 7104 15997 7113 16031
rect 7113 15997 7147 16031
rect 7147 15997 7156 16031
rect 7104 15988 7156 15997
rect 7196 16031 7248 16040
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 7288 15988 7340 16040
rect 7564 15988 7616 16040
rect 8024 15988 8076 16040
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 5724 15920 5776 15972
rect 7932 15920 7984 15972
rect 8760 16031 8812 16040
rect 8760 15997 8769 16031
rect 8769 15997 8803 16031
rect 8803 15997 8812 16031
rect 8760 15988 8812 15997
rect 9312 15988 9364 16040
rect 9588 16056 9640 16108
rect 9680 15988 9732 16040
rect 5816 15852 5868 15904
rect 6644 15895 6696 15904
rect 6644 15861 6653 15895
rect 6653 15861 6687 15895
rect 6687 15861 6696 15895
rect 6644 15852 6696 15861
rect 7564 15895 7616 15904
rect 7564 15861 7573 15895
rect 7573 15861 7607 15895
rect 7607 15861 7616 15895
rect 7564 15852 7616 15861
rect 9404 15852 9456 15904
rect 9588 15895 9640 15904
rect 9588 15861 9597 15895
rect 9597 15861 9631 15895
rect 9631 15861 9640 15895
rect 9588 15852 9640 15861
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 11704 15988 11756 16040
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 11980 15988 12032 16040
rect 10140 15852 10192 15904
rect 10232 15895 10284 15904
rect 10232 15861 10241 15895
rect 10241 15861 10275 15895
rect 10275 15861 10284 15895
rect 10232 15852 10284 15861
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 4322 15750 4374 15802
rect 4386 15750 4438 15802
rect 4450 15750 4502 15802
rect 4514 15750 4566 15802
rect 4578 15750 4630 15802
rect 10722 15750 10774 15802
rect 10786 15750 10838 15802
rect 10850 15750 10902 15802
rect 10914 15750 10966 15802
rect 10978 15750 11030 15802
rect 1676 15691 1728 15700
rect 1676 15657 1685 15691
rect 1685 15657 1719 15691
rect 1719 15657 1728 15691
rect 1676 15648 1728 15657
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 3516 15691 3568 15700
rect 3516 15657 3525 15691
rect 3525 15657 3559 15691
rect 3559 15657 3568 15691
rect 3516 15648 3568 15657
rect 4160 15648 4212 15700
rect 6184 15648 6236 15700
rect 2136 15512 2188 15564
rect 2412 15512 2464 15564
rect 2504 15555 2556 15564
rect 2504 15521 2513 15555
rect 2513 15521 2547 15555
rect 2547 15521 2556 15555
rect 2504 15512 2556 15521
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 3608 15580 3660 15632
rect 6000 15580 6052 15632
rect 4252 15512 4304 15564
rect 4620 15512 4672 15564
rect 5080 15512 5132 15564
rect 6092 15555 6144 15564
rect 6092 15521 6101 15555
rect 6101 15521 6135 15555
rect 6135 15521 6144 15555
rect 6092 15512 6144 15521
rect 6368 15555 6420 15564
rect 6368 15521 6377 15555
rect 6377 15521 6411 15555
rect 6411 15521 6420 15555
rect 6368 15512 6420 15521
rect 8484 15691 8536 15700
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 8668 15691 8720 15700
rect 8668 15657 8677 15691
rect 8677 15657 8711 15691
rect 8711 15657 8720 15691
rect 8668 15648 8720 15657
rect 10232 15648 10284 15700
rect 11060 15648 11112 15700
rect 11152 15648 11204 15700
rect 11336 15691 11388 15700
rect 11336 15657 11345 15691
rect 11345 15657 11379 15691
rect 11379 15657 11388 15691
rect 11336 15648 11388 15657
rect 11704 15648 11756 15700
rect 7012 15512 7064 15564
rect 7196 15555 7248 15564
rect 7196 15521 7205 15555
rect 7205 15521 7239 15555
rect 7239 15521 7248 15555
rect 7196 15512 7248 15521
rect 7656 15555 7708 15564
rect 7656 15521 7665 15555
rect 7665 15521 7699 15555
rect 7699 15521 7708 15555
rect 7656 15512 7708 15521
rect 7840 15512 7892 15564
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 8024 15555 8076 15564
rect 8024 15521 8033 15555
rect 8033 15521 8067 15555
rect 8067 15521 8076 15555
rect 8024 15512 8076 15521
rect 8208 15512 8260 15564
rect 2320 15444 2372 15496
rect 3516 15444 3568 15496
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 8576 15555 8628 15564
rect 8576 15521 8618 15555
rect 8618 15521 8628 15555
rect 8576 15512 8628 15521
rect 8944 15512 8996 15564
rect 9588 15580 9640 15632
rect 9772 15580 9824 15632
rect 8760 15444 8812 15496
rect 9404 15555 9456 15564
rect 9404 15521 9413 15555
rect 9413 15521 9447 15555
rect 9447 15521 9456 15555
rect 9404 15512 9456 15521
rect 9680 15444 9732 15496
rect 10692 15580 10744 15632
rect 2412 15376 2464 15428
rect 5540 15376 5592 15428
rect 8576 15376 8628 15428
rect 9956 15444 10008 15496
rect 10324 15444 10376 15496
rect 10232 15376 10284 15428
rect 10968 15376 11020 15428
rect 11520 15512 11572 15564
rect 11796 15444 11848 15496
rect 11612 15376 11664 15428
rect 12348 15444 12400 15496
rect 12072 15376 12124 15428
rect 2044 15308 2096 15360
rect 2688 15308 2740 15360
rect 2780 15308 2832 15360
rect 4528 15308 4580 15360
rect 7196 15308 7248 15360
rect 9404 15308 9456 15360
rect 9588 15308 9640 15360
rect 9864 15308 9916 15360
rect 3662 15206 3714 15258
rect 3726 15206 3778 15258
rect 3790 15206 3842 15258
rect 3854 15206 3906 15258
rect 3918 15206 3970 15258
rect 10062 15206 10114 15258
rect 10126 15206 10178 15258
rect 10190 15206 10242 15258
rect 10254 15206 10306 15258
rect 10318 15206 10370 15258
rect 2044 15104 2096 15156
rect 2412 15104 2464 15156
rect 2228 15011 2280 15020
rect 2228 14977 2237 15011
rect 2237 14977 2271 15011
rect 2271 14977 2280 15011
rect 2228 14968 2280 14977
rect 3424 15036 3476 15088
rect 5540 15104 5592 15156
rect 5816 15104 5868 15156
rect 3148 14900 3200 14952
rect 1952 14875 2004 14884
rect 1952 14841 1970 14875
rect 1970 14841 2004 14875
rect 1952 14832 2004 14841
rect 2596 14832 2648 14884
rect 5080 15036 5132 15088
rect 6184 15036 6236 15088
rect 8392 15104 8444 15156
rect 8668 15104 8720 15156
rect 4160 14943 4212 14952
rect 4160 14909 4169 14943
rect 4169 14909 4203 14943
rect 4203 14909 4212 14943
rect 4160 14900 4212 14909
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4528 14943 4580 14952
rect 4528 14909 4537 14943
rect 4537 14909 4571 14943
rect 4571 14909 4580 14943
rect 4528 14900 4580 14909
rect 4620 14900 4672 14952
rect 2780 14764 2832 14816
rect 4804 14875 4856 14884
rect 4804 14841 4813 14875
rect 4813 14841 4847 14875
rect 4847 14841 4856 14875
rect 4804 14832 4856 14841
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 6092 15011 6144 15020
rect 6092 14977 6101 15011
rect 6101 14977 6135 15011
rect 6135 14977 6144 15011
rect 6092 14968 6144 14977
rect 6736 14968 6788 15020
rect 7656 15036 7708 15088
rect 11888 15104 11940 15156
rect 7840 14968 7892 15020
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 5540 14900 5592 14952
rect 5080 14764 5132 14816
rect 5356 14807 5408 14816
rect 5356 14773 5365 14807
rect 5365 14773 5399 14807
rect 5399 14773 5408 14807
rect 7196 14900 7248 14952
rect 7288 14943 7340 14952
rect 7288 14909 7297 14943
rect 7297 14909 7331 14943
rect 7331 14909 7340 14943
rect 7288 14900 7340 14909
rect 9864 15036 9916 15088
rect 9220 14968 9272 15020
rect 9956 14968 10008 15020
rect 10692 15036 10744 15088
rect 5908 14832 5960 14884
rect 6644 14832 6696 14884
rect 8300 14832 8352 14884
rect 5356 14764 5408 14773
rect 6552 14807 6604 14816
rect 6552 14773 6561 14807
rect 6561 14773 6595 14807
rect 6595 14773 6604 14807
rect 6552 14764 6604 14773
rect 6920 14764 6972 14816
rect 7840 14807 7892 14816
rect 7840 14773 7849 14807
rect 7849 14773 7883 14807
rect 7883 14773 7892 14807
rect 9680 14943 9732 14952
rect 9680 14909 9689 14943
rect 9689 14909 9723 14943
rect 9723 14909 9732 14943
rect 9680 14900 9732 14909
rect 10048 14943 10100 14952
rect 10048 14909 10057 14943
rect 10057 14909 10091 14943
rect 10091 14909 10100 14943
rect 10048 14900 10100 14909
rect 11060 14968 11112 15020
rect 11796 15036 11848 15088
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 11336 14943 11388 14952
rect 11336 14909 11345 14943
rect 11345 14909 11379 14943
rect 11379 14909 11388 14943
rect 11336 14900 11388 14909
rect 12348 14900 12400 14952
rect 11704 14832 11756 14884
rect 7840 14764 7892 14773
rect 9128 14807 9180 14816
rect 9128 14773 9137 14807
rect 9137 14773 9171 14807
rect 9171 14773 9180 14807
rect 9128 14764 9180 14773
rect 9772 14764 9824 14816
rect 11152 14764 11204 14816
rect 11244 14764 11296 14816
rect 11612 14764 11664 14816
rect 4322 14662 4374 14714
rect 4386 14662 4438 14714
rect 4450 14662 4502 14714
rect 4514 14662 4566 14714
rect 4578 14662 4630 14714
rect 10722 14662 10774 14714
rect 10786 14662 10838 14714
rect 10850 14662 10902 14714
rect 10914 14662 10966 14714
rect 10978 14662 11030 14714
rect 2872 14560 2924 14612
rect 3148 14560 3200 14612
rect 4160 14560 4212 14612
rect 4804 14560 4856 14612
rect 848 14467 900 14476
rect 848 14433 857 14467
rect 857 14433 891 14467
rect 891 14433 900 14467
rect 848 14424 900 14433
rect 1400 14424 1452 14476
rect 2136 14467 2188 14476
rect 2136 14433 2145 14467
rect 2145 14433 2179 14467
rect 2179 14433 2188 14467
rect 2136 14424 2188 14433
rect 2688 14467 2740 14476
rect 2688 14433 2697 14467
rect 2697 14433 2731 14467
rect 2731 14433 2740 14467
rect 2688 14424 2740 14433
rect 2780 14424 2832 14476
rect 1952 14356 2004 14408
rect 2228 14356 2280 14408
rect 3240 14424 3292 14476
rect 3424 14467 3476 14476
rect 3424 14433 3433 14467
rect 3433 14433 3467 14467
rect 3467 14433 3476 14467
rect 3424 14424 3476 14433
rect 3608 14467 3660 14476
rect 3608 14433 3617 14467
rect 3617 14433 3651 14467
rect 3651 14433 3660 14467
rect 3608 14424 3660 14433
rect 3700 14356 3752 14408
rect 4252 14535 4304 14544
rect 4252 14501 4261 14535
rect 4261 14501 4295 14535
rect 4295 14501 4304 14535
rect 4252 14492 4304 14501
rect 5080 14399 5132 14408
rect 5080 14365 5089 14399
rect 5089 14365 5123 14399
rect 5123 14365 5132 14399
rect 5080 14356 5132 14365
rect 1768 14220 1820 14272
rect 2596 14220 2648 14272
rect 3608 14220 3660 14272
rect 3976 14220 4028 14272
rect 4344 14220 4396 14272
rect 5356 14399 5408 14408
rect 5356 14365 5365 14399
rect 5365 14365 5399 14399
rect 5399 14365 5408 14399
rect 5356 14356 5408 14365
rect 5540 14424 5592 14476
rect 6092 14560 6144 14612
rect 6368 14560 6420 14612
rect 6276 14492 6328 14544
rect 6920 14467 6972 14476
rect 6920 14433 6929 14467
rect 6929 14433 6963 14467
rect 6963 14433 6972 14467
rect 6920 14424 6972 14433
rect 8484 14560 8536 14612
rect 9128 14560 9180 14612
rect 8392 14492 8444 14544
rect 8944 14492 8996 14544
rect 7288 14356 7340 14408
rect 6736 14331 6788 14340
rect 6736 14297 6745 14331
rect 6745 14297 6779 14331
rect 6779 14297 6788 14331
rect 6736 14288 6788 14297
rect 6828 14331 6880 14340
rect 6828 14297 6837 14331
rect 6837 14297 6871 14331
rect 6871 14297 6880 14331
rect 6828 14288 6880 14297
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 8116 14467 8168 14476
rect 8116 14433 8125 14467
rect 8125 14433 8159 14467
rect 8159 14433 8168 14467
rect 8116 14424 8168 14433
rect 8484 14467 8536 14476
rect 8484 14433 8493 14467
rect 8493 14433 8527 14467
rect 8527 14433 8536 14467
rect 8484 14424 8536 14433
rect 8392 14399 8444 14408
rect 8392 14365 8401 14399
rect 8401 14365 8435 14399
rect 8435 14365 8444 14399
rect 8392 14356 8444 14365
rect 5448 14220 5500 14272
rect 5724 14220 5776 14272
rect 7932 14331 7984 14340
rect 7932 14297 7941 14331
rect 7941 14297 7975 14331
rect 7975 14297 7984 14331
rect 7932 14288 7984 14297
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 9036 14399 9088 14408
rect 9036 14365 9045 14399
rect 9045 14365 9079 14399
rect 9079 14365 9088 14399
rect 9036 14356 9088 14365
rect 9312 14356 9364 14408
rect 10048 14560 10100 14612
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9956 14424 10008 14476
rect 9496 14356 9548 14365
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 9772 14356 9824 14365
rect 11060 14424 11112 14476
rect 10508 14356 10560 14408
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 11888 14424 11940 14476
rect 12072 14467 12124 14476
rect 12072 14433 12081 14467
rect 12081 14433 12115 14467
rect 12115 14433 12124 14467
rect 12072 14424 12124 14433
rect 7104 14220 7156 14272
rect 8760 14220 8812 14272
rect 9036 14220 9088 14272
rect 10508 14220 10560 14272
rect 10600 14263 10652 14272
rect 10600 14229 10609 14263
rect 10609 14229 10643 14263
rect 10643 14229 10652 14263
rect 10600 14220 10652 14229
rect 3662 14118 3714 14170
rect 3726 14118 3778 14170
rect 3790 14118 3842 14170
rect 3854 14118 3906 14170
rect 3918 14118 3970 14170
rect 10062 14118 10114 14170
rect 10126 14118 10178 14170
rect 10190 14118 10242 14170
rect 10254 14118 10306 14170
rect 10318 14118 10370 14170
rect 1676 14016 1728 14068
rect 2320 14016 2372 14068
rect 1492 13880 1544 13932
rect 1676 13880 1728 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2228 13812 2280 13864
rect 2412 13880 2464 13932
rect 5080 14016 5132 14068
rect 6092 14059 6144 14068
rect 6092 14025 6101 14059
rect 6101 14025 6135 14059
rect 6135 14025 6144 14059
rect 6092 14016 6144 14025
rect 6828 14059 6880 14068
rect 6828 14025 6837 14059
rect 6837 14025 6871 14059
rect 6871 14025 6880 14059
rect 6828 14016 6880 14025
rect 9772 14016 9824 14068
rect 4804 13948 4856 14000
rect 5724 13948 5776 14000
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 4988 13812 5040 13864
rect 5632 13812 5684 13864
rect 7932 13948 7984 14000
rect 10600 14016 10652 14068
rect 11704 14016 11756 14068
rect 6460 13880 6512 13932
rect 7564 13880 7616 13932
rect 6552 13855 6604 13864
rect 6552 13821 6561 13855
rect 6561 13821 6595 13855
rect 6595 13821 6604 13855
rect 6552 13812 6604 13821
rect 6644 13812 6696 13864
rect 9864 13812 9916 13864
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 2596 13744 2648 13796
rect 2412 13676 2464 13728
rect 3240 13744 3292 13796
rect 3424 13744 3476 13796
rect 4344 13744 4396 13796
rect 7380 13744 7432 13796
rect 8944 13744 8996 13796
rect 9404 13744 9456 13796
rect 9956 13744 10008 13796
rect 10600 13812 10652 13864
rect 6368 13676 6420 13728
rect 6828 13676 6880 13728
rect 11244 13812 11296 13864
rect 11520 13812 11572 13864
rect 11888 13855 11940 13864
rect 11888 13821 11897 13855
rect 11897 13821 11931 13855
rect 11931 13821 11940 13855
rect 11888 13812 11940 13821
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 11152 13676 11204 13728
rect 11612 13787 11664 13796
rect 11612 13753 11621 13787
rect 11621 13753 11655 13787
rect 11655 13753 11664 13787
rect 11612 13744 11664 13753
rect 4322 13574 4374 13626
rect 4386 13574 4438 13626
rect 4450 13574 4502 13626
rect 4514 13574 4566 13626
rect 4578 13574 4630 13626
rect 10722 13574 10774 13626
rect 10786 13574 10838 13626
rect 10850 13574 10902 13626
rect 10914 13574 10966 13626
rect 10978 13574 11030 13626
rect 2412 13515 2464 13524
rect 2412 13481 2421 13515
rect 2421 13481 2455 13515
rect 2455 13481 2464 13515
rect 2412 13472 2464 13481
rect 2964 13472 3016 13524
rect 6368 13472 6420 13524
rect 6736 13472 6788 13524
rect 7564 13472 7616 13524
rect 2596 13447 2648 13456
rect 2596 13413 2605 13447
rect 2605 13413 2639 13447
rect 2639 13413 2648 13447
rect 2596 13404 2648 13413
rect 7288 13404 7340 13456
rect 8576 13404 8628 13456
rect 9220 13472 9272 13524
rect 10600 13472 10652 13524
rect 1952 13379 2004 13388
rect 1952 13345 1970 13379
rect 1970 13345 2004 13379
rect 1952 13336 2004 13345
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 2780 13336 2832 13388
rect 3240 13336 3292 13388
rect 4620 13336 4672 13388
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 5540 13336 5592 13388
rect 6644 13336 6696 13388
rect 7104 13336 7156 13388
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 4068 13268 4120 13320
rect 9404 13336 9456 13388
rect 10600 13336 10652 13388
rect 11612 13404 11664 13456
rect 11152 13379 11204 13388
rect 11152 13345 11161 13379
rect 11161 13345 11195 13379
rect 11195 13345 11204 13379
rect 11152 13336 11204 13345
rect 9312 13268 9364 13320
rect 2504 13200 2556 13252
rect 4436 13132 4488 13184
rect 4896 13132 4948 13184
rect 7288 13132 7340 13184
rect 8116 13132 8168 13184
rect 3662 13030 3714 13082
rect 3726 13030 3778 13082
rect 3790 13030 3842 13082
rect 3854 13030 3906 13082
rect 3918 13030 3970 13082
rect 10062 13030 10114 13082
rect 10126 13030 10178 13082
rect 10190 13030 10242 13082
rect 10254 13030 10306 13082
rect 10318 13030 10370 13082
rect 2320 12928 2372 12980
rect 3240 12928 3292 12980
rect 6552 12928 6604 12980
rect 7748 12928 7800 12980
rect 7932 12928 7984 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 2780 12860 2832 12912
rect 5172 12860 5224 12912
rect 5540 12903 5592 12912
rect 5540 12869 5549 12903
rect 5549 12869 5583 12903
rect 5583 12869 5592 12903
rect 5540 12860 5592 12869
rect 4620 12792 4672 12844
rect 1400 12724 1452 12776
rect 2044 12724 2096 12776
rect 2688 12767 2740 12776
rect 2688 12733 2697 12767
rect 2697 12733 2731 12767
rect 2731 12733 2740 12767
rect 2688 12724 2740 12733
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 4160 12767 4212 12776
rect 4160 12733 4169 12767
rect 4169 12733 4203 12767
rect 4203 12733 4212 12767
rect 4160 12724 4212 12733
rect 4252 12724 4304 12776
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 848 12699 900 12708
rect 848 12665 857 12699
rect 857 12665 891 12699
rect 891 12665 900 12699
rect 848 12656 900 12665
rect 3976 12656 4028 12708
rect 4896 12724 4948 12776
rect 5632 12724 5684 12776
rect 6828 12860 6880 12912
rect 9680 12860 9732 12912
rect 11980 12903 12032 12912
rect 11980 12869 11989 12903
rect 11989 12869 12023 12903
rect 12023 12869 12032 12903
rect 11980 12860 12032 12869
rect 7472 12792 7524 12844
rect 7748 12792 7800 12844
rect 6460 12767 6512 12776
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 6460 12733 6469 12767
rect 6469 12733 6503 12767
rect 6503 12733 6512 12767
rect 6460 12724 6512 12733
rect 6552 12767 6604 12776
rect 6552 12733 6561 12767
rect 6561 12733 6595 12767
rect 6595 12733 6604 12767
rect 6552 12724 6604 12733
rect 7012 12724 7064 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 7932 12767 7984 12776
rect 7932 12733 7941 12767
rect 7941 12733 7975 12767
rect 7975 12733 7984 12767
rect 7932 12724 7984 12733
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 6920 12656 6972 12708
rect 8300 12724 8352 12776
rect 8668 12835 8720 12844
rect 8668 12801 8677 12835
rect 8677 12801 8711 12835
rect 8711 12801 8720 12835
rect 8668 12792 8720 12801
rect 9496 12792 9548 12844
rect 10416 12792 10468 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 8944 12767 8996 12776
rect 8944 12733 8951 12767
rect 8951 12733 8996 12767
rect 8944 12724 8996 12733
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 11244 12724 11296 12776
rect 11612 12767 11664 12776
rect 11612 12733 11621 12767
rect 11621 12733 11655 12767
rect 11655 12733 11664 12767
rect 11612 12724 11664 12733
rect 7840 12588 7892 12640
rect 8944 12588 8996 12640
rect 9772 12588 9824 12640
rect 4322 12486 4374 12538
rect 4386 12486 4438 12538
rect 4450 12486 4502 12538
rect 4514 12486 4566 12538
rect 4578 12486 4630 12538
rect 10722 12486 10774 12538
rect 10786 12486 10838 12538
rect 10850 12486 10902 12538
rect 10914 12486 10966 12538
rect 10978 12486 11030 12538
rect 480 12384 532 12436
rect 756 12384 808 12436
rect 2688 12384 2740 12436
rect 2872 12384 2924 12436
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 4528 12384 4580 12436
rect 4712 12384 4764 12436
rect 1400 12359 1452 12368
rect 1400 12325 1409 12359
rect 1409 12325 1443 12359
rect 1443 12325 1452 12359
rect 1400 12316 1452 12325
rect 1584 12316 1636 12368
rect 388 12248 440 12300
rect 1400 12180 1452 12232
rect 2688 12180 2740 12232
rect 3424 12316 3476 12368
rect 3976 12248 4028 12300
rect 3148 12180 3200 12232
rect 4252 12291 4304 12300
rect 4252 12257 4261 12291
rect 4261 12257 4295 12291
rect 4295 12257 4304 12291
rect 4252 12248 4304 12257
rect 4344 12248 4396 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 4160 12112 4212 12164
rect 5172 12248 5224 12300
rect 4896 12180 4948 12232
rect 6644 12384 6696 12436
rect 8208 12384 8260 12436
rect 5448 12291 5500 12300
rect 5448 12257 5457 12291
rect 5457 12257 5491 12291
rect 5491 12257 5500 12291
rect 5448 12248 5500 12257
rect 5632 12291 5684 12300
rect 5632 12257 5641 12291
rect 5641 12257 5675 12291
rect 5675 12257 5684 12291
rect 5632 12248 5684 12257
rect 6368 12291 6420 12300
rect 6368 12257 6377 12291
rect 6377 12257 6411 12291
rect 6411 12257 6420 12291
rect 6368 12248 6420 12257
rect 7012 12316 7064 12368
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 7104 12248 7156 12300
rect 7472 12316 7524 12368
rect 7656 12291 7708 12300
rect 7656 12257 7665 12291
rect 7665 12257 7699 12291
rect 7699 12257 7708 12291
rect 7656 12248 7708 12257
rect 7932 12316 7984 12368
rect 8116 12248 8168 12300
rect 9680 12384 9732 12436
rect 8944 12316 8996 12368
rect 8392 12248 8444 12300
rect 8852 12291 8904 12300
rect 8852 12257 8861 12291
rect 8861 12257 8895 12291
rect 8895 12257 8904 12291
rect 9864 12316 9916 12368
rect 8852 12248 8904 12257
rect 6276 12112 6328 12164
rect 7288 12112 7340 12164
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9680 12112 9732 12164
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10416 12316 10468 12368
rect 10784 12248 10836 12300
rect 10968 12291 11020 12300
rect 10968 12257 10977 12291
rect 10977 12257 11011 12291
rect 11011 12257 11020 12291
rect 10968 12248 11020 12257
rect 11152 12291 11204 12300
rect 11152 12257 11161 12291
rect 11161 12257 11195 12291
rect 11195 12257 11204 12291
rect 11152 12248 11204 12257
rect 11612 12384 11664 12436
rect 10968 12112 11020 12164
rect 11244 12112 11296 12164
rect 11704 12248 11756 12300
rect 11888 12223 11940 12232
rect 11888 12189 11897 12223
rect 11897 12189 11931 12223
rect 11931 12189 11940 12223
rect 11888 12180 11940 12189
rect 11612 12112 11664 12164
rect 12532 12112 12584 12164
rect 572 12044 624 12096
rect 3240 12044 3292 12096
rect 4620 12044 4672 12096
rect 5356 12087 5408 12096
rect 5356 12053 5365 12087
rect 5365 12053 5399 12087
rect 5399 12053 5408 12087
rect 5356 12044 5408 12053
rect 5632 12044 5684 12096
rect 6000 12044 6052 12096
rect 6736 12044 6788 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 7656 12044 7708 12096
rect 8392 12087 8444 12096
rect 8392 12053 8401 12087
rect 8401 12053 8435 12087
rect 8435 12053 8444 12087
rect 8392 12044 8444 12053
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9220 12044 9272 12096
rect 10324 12044 10376 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 10600 12044 10652 12096
rect 11336 12044 11388 12096
rect 3662 11942 3714 11994
rect 3726 11942 3778 11994
rect 3790 11942 3842 11994
rect 3854 11942 3906 11994
rect 3918 11942 3970 11994
rect 10062 11942 10114 11994
rect 10126 11942 10178 11994
rect 10190 11942 10242 11994
rect 10254 11942 10306 11994
rect 10318 11942 10370 11994
rect 1032 11840 1084 11892
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 2872 11840 2924 11892
rect 4160 11704 4212 11756
rect 1124 11636 1176 11688
rect 5448 11772 5500 11824
rect 6000 11772 6052 11824
rect 6368 11840 6420 11892
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 8576 11840 8628 11892
rect 8668 11840 8720 11892
rect 9864 11840 9916 11892
rect 11152 11840 11204 11892
rect 11888 11840 11940 11892
rect 9588 11772 9640 11824
rect 10968 11772 11020 11824
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 5080 11636 5132 11688
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 5448 11636 5500 11645
rect 5632 11636 5684 11688
rect 5816 11636 5868 11688
rect 1584 11611 1636 11620
rect 1584 11577 1618 11611
rect 1618 11577 1636 11611
rect 1584 11568 1636 11577
rect 2228 11568 2280 11620
rect 4344 11568 4396 11620
rect 4712 11568 4764 11620
rect 4988 11568 5040 11620
rect 6000 11636 6052 11688
rect 6736 11679 6788 11688
rect 6736 11645 6745 11679
rect 6745 11645 6779 11679
rect 6779 11645 6788 11679
rect 6736 11636 6788 11645
rect 6368 11568 6420 11620
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 7472 11636 7524 11688
rect 8208 11704 8260 11756
rect 8024 11636 8076 11688
rect 8208 11568 8260 11620
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 8484 11704 8536 11756
rect 8576 11679 8628 11688
rect 8576 11645 8585 11679
rect 8585 11645 8619 11679
rect 8619 11645 8628 11679
rect 8576 11636 8628 11645
rect 8852 11636 8904 11688
rect 9496 11636 9548 11688
rect 9680 11636 9732 11688
rect 9956 11636 10008 11688
rect 10416 11704 10468 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10232 11679 10284 11688
rect 10232 11645 10241 11679
rect 10241 11645 10275 11679
rect 10275 11645 10284 11679
rect 10232 11636 10284 11645
rect 10692 11636 10744 11688
rect 11152 11636 11204 11688
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 11704 11568 11756 11620
rect 1032 11543 1084 11552
rect 1032 11509 1041 11543
rect 1041 11509 1075 11543
rect 1075 11509 1084 11543
rect 1032 11500 1084 11509
rect 4252 11500 4304 11552
rect 7012 11500 7064 11552
rect 7840 11500 7892 11552
rect 8116 11500 8168 11552
rect 10048 11500 10100 11552
rect 10324 11500 10376 11552
rect 11244 11543 11296 11552
rect 11244 11509 11253 11543
rect 11253 11509 11287 11543
rect 11287 11509 11296 11543
rect 11244 11500 11296 11509
rect 4322 11398 4374 11450
rect 4386 11398 4438 11450
rect 4450 11398 4502 11450
rect 4514 11398 4566 11450
rect 4578 11398 4630 11450
rect 10722 11398 10774 11450
rect 10786 11398 10838 11450
rect 10850 11398 10902 11450
rect 10914 11398 10966 11450
rect 10978 11398 11030 11450
rect 4712 11296 4764 11348
rect 6644 11296 6696 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7104 11296 7156 11348
rect 7288 11296 7340 11348
rect 7380 11296 7432 11348
rect 8208 11296 8260 11348
rect 8852 11296 8904 11348
rect 8944 11296 8996 11348
rect 10232 11296 10284 11348
rect 10692 11296 10744 11348
rect 1676 11228 1728 11280
rect 5632 11228 5684 11280
rect 1952 11203 2004 11212
rect 1952 11169 1970 11203
rect 1970 11169 2004 11203
rect 1952 11160 2004 11169
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 5080 11203 5132 11212
rect 5080 11169 5089 11203
rect 5089 11169 5123 11203
rect 5123 11169 5132 11203
rect 5080 11160 5132 11169
rect 5356 11203 5408 11212
rect 5356 11169 5365 11203
rect 5365 11169 5399 11203
rect 5399 11169 5408 11203
rect 5356 11160 5408 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 6092 11203 6144 11212
rect 6092 11169 6101 11203
rect 6101 11169 6135 11203
rect 6135 11169 6144 11203
rect 6092 11160 6144 11169
rect 7472 11228 7524 11280
rect 9588 11228 9640 11280
rect 6552 11160 6604 11212
rect 6920 11160 6972 11212
rect 7012 11203 7064 11212
rect 7012 11169 7021 11203
rect 7021 11169 7055 11203
rect 7055 11169 7064 11203
rect 7012 11160 7064 11169
rect 7932 11160 7984 11212
rect 8116 11160 8168 11212
rect 9772 11203 9824 11212
rect 9772 11169 9781 11203
rect 9781 11169 9815 11203
rect 9815 11169 9824 11203
rect 9772 11160 9824 11169
rect 10048 11203 10100 11212
rect 10048 11169 10057 11203
rect 10057 11169 10091 11203
rect 10091 11169 10100 11203
rect 10048 11160 10100 11169
rect 10968 11228 11020 11280
rect 10416 11203 10468 11212
rect 10416 11169 10425 11203
rect 10425 11169 10459 11203
rect 10459 11169 10468 11203
rect 10416 11160 10468 11169
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 7380 11092 7432 11144
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 9680 11135 9732 11144
rect 9680 11101 9689 11135
rect 9689 11101 9723 11135
rect 9723 11101 9732 11135
rect 9680 11092 9732 11101
rect 10876 11092 10928 11144
rect 2504 11067 2556 11076
rect 2504 11033 2513 11067
rect 2513 11033 2547 11067
rect 2547 11033 2556 11067
rect 2504 11024 2556 11033
rect 4712 11024 4764 11076
rect 7656 11024 7708 11076
rect 10324 11024 10376 11076
rect 12164 11160 12216 11212
rect 1584 10956 1636 11008
rect 5540 10956 5592 11008
rect 11244 10956 11296 11008
rect 3662 10854 3714 10906
rect 3726 10854 3778 10906
rect 3790 10854 3842 10906
rect 3854 10854 3906 10906
rect 3918 10854 3970 10906
rect 10062 10854 10114 10906
rect 10126 10854 10178 10906
rect 10190 10854 10242 10906
rect 10254 10854 10306 10906
rect 10318 10854 10370 10906
rect 2320 10795 2372 10804
rect 2320 10761 2329 10795
rect 2329 10761 2363 10795
rect 2363 10761 2372 10795
rect 2320 10752 2372 10761
rect 3976 10752 4028 10804
rect 4160 10752 4212 10804
rect 5724 10752 5776 10804
rect 8116 10752 8168 10804
rect 3332 10684 3384 10736
rect 940 10616 992 10668
rect 1584 10616 1636 10668
rect 6920 10684 6972 10736
rect 9128 10727 9180 10736
rect 9128 10693 9137 10727
rect 9137 10693 9171 10727
rect 9171 10693 9180 10727
rect 9128 10684 9180 10693
rect 9588 10752 9640 10804
rect 9680 10752 9732 10804
rect 10968 10752 11020 10804
rect 11980 10684 12032 10736
rect 4068 10616 4120 10668
rect 1400 10548 1452 10600
rect 1952 10548 2004 10600
rect 2964 10548 3016 10600
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 5908 10616 5960 10668
rect 6184 10616 6236 10668
rect 6460 10616 6512 10668
rect 7840 10616 7892 10668
rect 9588 10616 9640 10668
rect 11244 10616 11296 10668
rect 664 10480 716 10532
rect 3148 10480 3200 10532
rect 2780 10412 2832 10464
rect 4068 10412 4120 10464
rect 4896 10548 4948 10600
rect 5172 10548 5224 10600
rect 5356 10548 5408 10600
rect 6552 10591 6604 10600
rect 6552 10557 6561 10591
rect 6561 10557 6595 10591
rect 6595 10557 6604 10591
rect 6552 10548 6604 10557
rect 6092 10480 6144 10532
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7380 10591 7432 10600
rect 7380 10557 7389 10591
rect 7389 10557 7423 10591
rect 7423 10557 7432 10591
rect 7380 10548 7432 10557
rect 7656 10591 7708 10600
rect 7656 10557 7665 10591
rect 7665 10557 7699 10591
rect 7699 10557 7708 10591
rect 7656 10548 7708 10557
rect 7104 10480 7156 10532
rect 8852 10480 8904 10532
rect 9680 10523 9732 10532
rect 9680 10489 9689 10523
rect 9689 10489 9723 10523
rect 9723 10489 9732 10523
rect 9680 10480 9732 10489
rect 9864 10523 9916 10532
rect 9864 10489 9873 10523
rect 9873 10489 9907 10523
rect 9907 10489 9916 10523
rect 10508 10548 10560 10600
rect 10600 10548 10652 10600
rect 11060 10548 11112 10600
rect 11796 10548 11848 10600
rect 9864 10480 9916 10489
rect 4988 10412 5040 10464
rect 5172 10412 5224 10464
rect 5540 10412 5592 10464
rect 6920 10412 6972 10464
rect 9404 10412 9456 10464
rect 10508 10412 10560 10464
rect 10876 10412 10928 10464
rect 11152 10412 11204 10464
rect 4322 10310 4374 10362
rect 4386 10310 4438 10362
rect 4450 10310 4502 10362
rect 4514 10310 4566 10362
rect 4578 10310 4630 10362
rect 10722 10310 10774 10362
rect 10786 10310 10838 10362
rect 10850 10310 10902 10362
rect 10914 10310 10966 10362
rect 10978 10310 11030 10362
rect 3056 10208 3108 10260
rect 1860 10140 1912 10192
rect 2964 10072 3016 10124
rect 3608 10072 3660 10124
rect 4620 10208 4672 10260
rect 5264 10208 5316 10260
rect 8576 10208 8628 10260
rect 9680 10208 9732 10260
rect 4896 10140 4948 10192
rect 5172 10140 5224 10192
rect 4620 10115 4672 10124
rect 4620 10081 4629 10115
rect 4629 10081 4663 10115
rect 4663 10081 4672 10115
rect 4620 10072 4672 10081
rect 4804 10115 4856 10124
rect 4804 10081 4813 10115
rect 4813 10081 4847 10115
rect 4847 10081 4856 10115
rect 4804 10072 4856 10081
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 3976 10047 4028 10056
rect 3976 10013 3985 10047
rect 3985 10013 4019 10047
rect 4019 10013 4028 10047
rect 3976 10004 4028 10013
rect 4160 10004 4212 10056
rect 4344 10004 4396 10056
rect 3332 9936 3384 9988
rect 4896 10004 4948 10056
rect 6276 10072 6328 10124
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 7932 10140 7984 10192
rect 7656 10004 7708 10056
rect 4804 9936 4856 9988
rect 6828 9936 6880 9988
rect 8484 10115 8536 10124
rect 8484 10081 8493 10115
rect 8493 10081 8527 10115
rect 8527 10081 8536 10115
rect 8484 10072 8536 10081
rect 8852 10072 8904 10124
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 9864 10140 9916 10192
rect 11428 10140 11480 10192
rect 10784 10072 10836 10124
rect 11060 10072 11112 10124
rect 11152 10115 11204 10124
rect 11152 10081 11161 10115
rect 11161 10081 11195 10115
rect 11195 10081 11204 10115
rect 11152 10072 11204 10081
rect 11796 10072 11848 10124
rect 11980 10115 12032 10124
rect 11980 10081 11989 10115
rect 11989 10081 12023 10115
rect 12023 10081 12032 10115
rect 11980 10072 12032 10081
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9128 10004 9180 10056
rect 9864 10004 9916 10056
rect 10508 10004 10560 10056
rect 12256 10004 12308 10056
rect 10416 9936 10468 9988
rect 1952 9868 2004 9920
rect 4160 9868 4212 9920
rect 5080 9868 5132 9920
rect 5816 9868 5868 9920
rect 6276 9911 6328 9920
rect 6276 9877 6285 9911
rect 6285 9877 6319 9911
rect 6319 9877 6328 9911
rect 6276 9868 6328 9877
rect 9680 9868 9732 9920
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 3662 9766 3714 9818
rect 3726 9766 3778 9818
rect 3790 9766 3842 9818
rect 3854 9766 3906 9818
rect 3918 9766 3970 9818
rect 10062 9766 10114 9818
rect 10126 9766 10178 9818
rect 10190 9766 10242 9818
rect 10254 9766 10306 9818
rect 10318 9766 10370 9818
rect 3148 9664 3200 9716
rect 3608 9664 3660 9716
rect 3976 9664 4028 9716
rect 4344 9664 4396 9716
rect 756 9596 808 9648
rect 3424 9596 3476 9648
rect 4068 9596 4120 9648
rect 5356 9596 5408 9648
rect 6552 9596 6604 9648
rect 7012 9596 7064 9648
rect 8852 9707 8904 9716
rect 8852 9673 8861 9707
rect 8861 9673 8895 9707
rect 8895 9673 8904 9707
rect 8852 9664 8904 9673
rect 10784 9664 10836 9716
rect 11796 9664 11848 9716
rect 1216 9571 1268 9580
rect 1216 9537 1225 9571
rect 1225 9537 1259 9571
rect 1259 9537 1268 9571
rect 1216 9528 1268 9537
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2412 9571 2464 9580
rect 2412 9537 2421 9571
rect 2421 9537 2455 9571
rect 2455 9537 2464 9571
rect 2412 9528 2464 9537
rect 4988 9528 5040 9580
rect 5540 9528 5592 9580
rect 1400 9460 1452 9512
rect 1860 9503 1912 9512
rect 1860 9469 1869 9503
rect 1869 9469 1903 9503
rect 1903 9469 1912 9503
rect 1860 9460 1912 9469
rect 848 9392 900 9444
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 3976 9460 4028 9512
rect 4160 9460 4212 9512
rect 2872 9367 2924 9376
rect 2872 9333 2881 9367
rect 2881 9333 2915 9367
rect 2915 9333 2924 9367
rect 2872 9324 2924 9333
rect 3884 9392 3936 9444
rect 5172 9460 5224 9512
rect 4988 9392 5040 9444
rect 3792 9324 3844 9376
rect 4068 9324 4120 9376
rect 4896 9324 4948 9376
rect 5908 9460 5960 9512
rect 6276 9503 6328 9512
rect 6276 9469 6285 9503
rect 6285 9469 6319 9503
rect 6319 9469 6328 9503
rect 6276 9460 6328 9469
rect 6644 9460 6696 9512
rect 6736 9460 6788 9512
rect 7656 9639 7708 9648
rect 7656 9605 7665 9639
rect 7665 9605 7699 9639
rect 7699 9605 7708 9639
rect 7656 9596 7708 9605
rect 7288 9503 7340 9512
rect 7288 9469 7297 9503
rect 7297 9469 7331 9503
rect 7331 9469 7340 9503
rect 7288 9460 7340 9469
rect 8208 9528 8260 9580
rect 9496 9528 9548 9580
rect 8392 9460 8444 9512
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10508 9528 10560 9580
rect 9956 9460 10008 9512
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10600 9503 10652 9512
rect 10048 9460 10100 9469
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 11704 9460 11756 9512
rect 7288 9324 7340 9376
rect 12164 9392 12216 9444
rect 7932 9367 7984 9376
rect 7932 9333 7941 9367
rect 7941 9333 7975 9367
rect 7975 9333 7984 9367
rect 7932 9324 7984 9333
rect 10600 9324 10652 9376
rect 4322 9222 4374 9274
rect 4386 9222 4438 9274
rect 4450 9222 4502 9274
rect 4514 9222 4566 9274
rect 4578 9222 4630 9274
rect 10722 9222 10774 9274
rect 10786 9222 10838 9274
rect 10850 9222 10902 9274
rect 10914 9222 10966 9274
rect 10978 9222 11030 9274
rect 1308 9120 1360 9172
rect 3424 9120 3476 9172
rect 3976 9120 4028 9172
rect 6828 9120 6880 9172
rect 7288 9120 7340 9172
rect 9128 9163 9180 9172
rect 9128 9129 9137 9163
rect 9137 9129 9171 9163
rect 9171 9129 9180 9163
rect 9128 9120 9180 9129
rect 11612 9120 11664 9172
rect 12164 9163 12216 9172
rect 12164 9129 12173 9163
rect 12173 9129 12207 9163
rect 12207 9129 12216 9163
rect 12164 9120 12216 9129
rect 7564 9052 7616 9104
rect 2228 8984 2280 9036
rect 2872 8984 2924 9036
rect 3148 8916 3200 8968
rect 2228 8780 2280 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 4620 8780 4672 8832
rect 4896 9027 4948 9036
rect 4896 8993 4905 9027
rect 4905 8993 4939 9027
rect 4939 8993 4948 9027
rect 4896 8984 4948 8993
rect 5540 8916 5592 8968
rect 5908 8984 5960 9036
rect 6460 8984 6512 9036
rect 6828 9027 6880 9036
rect 6828 8993 6837 9027
rect 6837 8993 6871 9027
rect 6871 8993 6880 9027
rect 6828 8984 6880 8993
rect 8484 9052 8536 9104
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 9680 9052 9732 9104
rect 6920 8916 6972 8968
rect 7288 8848 7340 8900
rect 8208 8848 8260 8900
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 6368 8780 6420 8832
rect 8300 8823 8352 8832
rect 8300 8789 8309 8823
rect 8309 8789 8343 8823
rect 8343 8789 8352 8823
rect 8300 8780 8352 8789
rect 9496 8984 9548 9036
rect 10048 9052 10100 9104
rect 9956 9027 10008 9036
rect 9956 8993 9965 9027
rect 9965 8993 9999 9027
rect 9999 8993 10008 9027
rect 9956 8984 10008 8993
rect 10416 9027 10468 9036
rect 10416 8993 10425 9027
rect 10425 8993 10459 9027
rect 10459 8993 10468 9027
rect 10416 8984 10468 8993
rect 9036 8848 9088 8900
rect 9496 8848 9548 8900
rect 8760 8780 8812 8832
rect 9588 8780 9640 8832
rect 10048 8848 10100 8900
rect 10508 8848 10560 8900
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 12440 9052 12492 9104
rect 11428 8984 11480 9036
rect 11980 8984 12032 9036
rect 12072 9027 12124 9036
rect 12072 8993 12081 9027
rect 12081 8993 12115 9027
rect 12115 8993 12124 9027
rect 12072 8984 12124 8993
rect 10968 8848 11020 8900
rect 11060 8848 11112 8900
rect 9956 8780 10008 8832
rect 11704 8780 11756 8832
rect 3662 8678 3714 8730
rect 3726 8678 3778 8730
rect 3790 8678 3842 8730
rect 3854 8678 3906 8730
rect 3918 8678 3970 8730
rect 10062 8678 10114 8730
rect 10126 8678 10178 8730
rect 10190 8678 10242 8730
rect 10254 8678 10306 8730
rect 10318 8678 10370 8730
rect 3148 8576 3200 8628
rect 3240 8619 3292 8628
rect 3240 8585 3249 8619
rect 3249 8585 3283 8619
rect 3283 8585 3292 8619
rect 3240 8576 3292 8585
rect 5540 8619 5592 8628
rect 5540 8585 5549 8619
rect 5549 8585 5583 8619
rect 5583 8585 5592 8619
rect 5540 8576 5592 8585
rect 6644 8619 6696 8628
rect 6644 8585 6653 8619
rect 6653 8585 6687 8619
rect 6687 8585 6696 8619
rect 6644 8576 6696 8585
rect 8484 8576 8536 8628
rect 4896 8508 4948 8560
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 4804 8440 4856 8492
rect 1400 8372 1452 8424
rect 1768 8415 1820 8424
rect 1768 8381 1777 8415
rect 1777 8381 1811 8415
rect 1811 8381 1820 8415
rect 1768 8372 1820 8381
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 2320 8372 2372 8424
rect 2504 8372 2556 8424
rect 3332 8372 3384 8424
rect 3608 8372 3660 8424
rect 4068 8372 4120 8424
rect 1124 8347 1176 8356
rect 1124 8313 1133 8347
rect 1133 8313 1167 8347
rect 1167 8313 1176 8347
rect 1124 8304 1176 8313
rect 3056 8304 3108 8356
rect 4528 8372 4580 8424
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 5724 8440 5776 8492
rect 4620 8304 4672 8356
rect 4804 8304 4856 8356
rect 5356 8415 5408 8424
rect 5356 8381 5365 8415
rect 5365 8381 5399 8415
rect 5399 8381 5408 8415
rect 5356 8372 5408 8381
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 7012 8440 7064 8492
rect 7564 8440 7616 8492
rect 6736 8415 6788 8424
rect 6736 8381 6745 8415
rect 6745 8381 6779 8415
rect 6779 8381 6788 8415
rect 6736 8372 6788 8381
rect 7288 8372 7340 8424
rect 8300 8372 8352 8424
rect 8668 8508 8720 8560
rect 9496 8508 9548 8560
rect 10692 8576 10744 8628
rect 11336 8576 11388 8628
rect 11612 8619 11664 8628
rect 11612 8585 11621 8619
rect 11621 8585 11655 8619
rect 11655 8585 11664 8619
rect 11612 8576 11664 8585
rect 9864 8508 9916 8560
rect 8852 8440 8904 8492
rect 9036 8415 9088 8424
rect 9036 8381 9045 8415
rect 9045 8381 9079 8415
rect 9079 8381 9088 8415
rect 9036 8372 9088 8381
rect 10416 8440 10468 8492
rect 12164 8508 12216 8560
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11336 8440 11388 8492
rect 9404 8347 9456 8356
rect 9404 8313 9413 8347
rect 9413 8313 9447 8347
rect 9447 8313 9456 8347
rect 9404 8304 9456 8313
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 11612 8304 11664 8356
rect 11980 8372 12032 8424
rect 11888 8347 11940 8356
rect 11888 8313 11897 8347
rect 11897 8313 11931 8347
rect 11931 8313 11940 8347
rect 11888 8304 11940 8313
rect 4322 8134 4374 8186
rect 4386 8134 4438 8186
rect 4450 8134 4502 8186
rect 4514 8134 4566 8186
rect 4578 8134 4630 8186
rect 10722 8134 10774 8186
rect 10786 8134 10838 8186
rect 10850 8134 10902 8186
rect 10914 8134 10966 8186
rect 10978 8134 11030 8186
rect 1860 8032 1912 8084
rect 2412 8032 2464 8084
rect 3608 8032 3660 8084
rect 4436 8032 4488 8084
rect 5080 8032 5132 8084
rect 5356 8032 5408 8084
rect 6184 8075 6236 8084
rect 6184 8041 6193 8075
rect 6193 8041 6227 8075
rect 6227 8041 6236 8075
rect 6184 8032 6236 8041
rect 1768 7964 1820 8016
rect 2688 7896 2740 7948
rect 2780 7896 2832 7948
rect 3056 7896 3108 7948
rect 4528 7896 4580 7948
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2412 7828 2464 7880
rect 2872 7828 2924 7880
rect 3332 7828 3384 7880
rect 4436 7760 4488 7812
rect 5356 7896 5408 7948
rect 5908 7896 5960 7948
rect 7012 7896 7064 7948
rect 7380 8032 7432 8084
rect 9036 8032 9088 8084
rect 9496 8075 9548 8084
rect 9496 8041 9505 8075
rect 9505 8041 9539 8075
rect 9539 8041 9548 8075
rect 9496 8032 9548 8041
rect 8024 7964 8076 8016
rect 8852 7964 8904 8016
rect 10324 8007 10376 8016
rect 10324 7973 10333 8007
rect 10333 7973 10367 8007
rect 10367 7973 10376 8007
rect 10324 7964 10376 7973
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 7380 7939 7432 7948
rect 7380 7905 7389 7939
rect 7389 7905 7423 7939
rect 7423 7905 7432 7939
rect 7380 7896 7432 7905
rect 8668 7896 8720 7948
rect 9220 7896 9272 7948
rect 9864 7939 9916 7948
rect 9864 7905 9873 7939
rect 9873 7905 9907 7939
rect 9907 7905 9916 7939
rect 9864 7896 9916 7905
rect 11244 7896 11296 7948
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 12164 7939 12216 7948
rect 12164 7905 12173 7939
rect 12173 7905 12207 7939
rect 12207 7905 12216 7939
rect 12164 7896 12216 7905
rect 5172 7760 5224 7812
rect 2780 7692 2832 7744
rect 4620 7735 4672 7744
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 9128 7871 9180 7880
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 12256 7828 12308 7880
rect 6644 7760 6696 7812
rect 7196 7760 7248 7812
rect 5632 7692 5684 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 9496 7692 9548 7744
rect 10324 7692 10376 7744
rect 11980 7735 12032 7744
rect 11980 7701 11989 7735
rect 11989 7701 12023 7735
rect 12023 7701 12032 7735
rect 11980 7692 12032 7701
rect 3662 7590 3714 7642
rect 3726 7590 3778 7642
rect 3790 7590 3842 7642
rect 3854 7590 3906 7642
rect 3918 7590 3970 7642
rect 10062 7590 10114 7642
rect 10126 7590 10178 7642
rect 10190 7590 10242 7642
rect 10254 7590 10306 7642
rect 10318 7590 10370 7642
rect 2412 7531 2464 7540
rect 2412 7497 2421 7531
rect 2421 7497 2455 7531
rect 2455 7497 2464 7531
rect 2412 7488 2464 7497
rect 2780 7531 2832 7540
rect 2780 7497 2789 7531
rect 2789 7497 2823 7531
rect 2823 7497 2832 7531
rect 2780 7488 2832 7497
rect 4528 7488 4580 7540
rect 3056 7420 3108 7472
rect 5356 7420 5408 7472
rect 6092 7420 6144 7472
rect 1492 7284 1544 7336
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2320 7327 2372 7336
rect 2320 7293 2329 7327
rect 2329 7293 2363 7327
rect 2363 7293 2372 7327
rect 2320 7284 2372 7293
rect 2412 7284 2464 7336
rect 2872 7352 2924 7404
rect 3148 7352 3200 7404
rect 2136 7216 2188 7268
rect 2964 7284 3016 7336
rect 4620 7216 4672 7268
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5908 7352 5960 7404
rect 7104 7488 7156 7540
rect 9864 7488 9916 7540
rect 11888 7488 11940 7540
rect 9128 7463 9180 7472
rect 9128 7429 9137 7463
rect 9137 7429 9171 7463
rect 9171 7429 9180 7463
rect 9128 7420 9180 7429
rect 6000 7284 6052 7336
rect 6552 7327 6604 7336
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 6644 7327 6696 7336
rect 6644 7293 6653 7327
rect 6653 7293 6687 7327
rect 6687 7293 6696 7327
rect 6644 7284 6696 7293
rect 7472 7352 7524 7404
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 7196 7284 7248 7336
rect 8852 7352 8904 7404
rect 5724 7259 5776 7268
rect 5724 7225 5733 7259
rect 5733 7225 5767 7259
rect 5767 7225 5776 7259
rect 5724 7216 5776 7225
rect 8484 7284 8536 7336
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 9220 7352 9272 7404
rect 9404 7352 9456 7404
rect 10600 7352 10652 7404
rect 11980 7284 12032 7336
rect 1676 7148 1728 7200
rect 5172 7148 5224 7200
rect 8024 7216 8076 7268
rect 6920 7148 6972 7200
rect 9312 7191 9364 7200
rect 9312 7157 9321 7191
rect 9321 7157 9355 7191
rect 9355 7157 9364 7191
rect 9312 7148 9364 7157
rect 4322 7046 4374 7098
rect 4386 7046 4438 7098
rect 4450 7046 4502 7098
rect 4514 7046 4566 7098
rect 4578 7046 4630 7098
rect 10722 7046 10774 7098
rect 10786 7046 10838 7098
rect 10850 7046 10902 7098
rect 10914 7046 10966 7098
rect 10978 7046 11030 7098
rect 1952 6944 2004 6996
rect 2412 6944 2464 6996
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2136 6876 2188 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 940 6783 992 6792
rect 940 6749 949 6783
rect 949 6749 983 6783
rect 983 6749 992 6783
rect 940 6740 992 6749
rect 2044 6783 2096 6792
rect 2044 6749 2053 6783
rect 2053 6749 2087 6783
rect 2087 6749 2096 6783
rect 2044 6740 2096 6749
rect 2136 6740 2188 6792
rect 3516 6740 3568 6792
rect 1860 6672 1912 6724
rect 1032 6604 1084 6656
rect 3056 6604 3108 6656
rect 4252 6808 4304 6860
rect 4896 6944 4948 6996
rect 7288 6944 7340 6996
rect 8024 6987 8076 6996
rect 8024 6953 8033 6987
rect 8033 6953 8067 6987
rect 8067 6953 8076 6987
rect 8024 6944 8076 6953
rect 4620 6851 4672 6860
rect 4620 6817 4629 6851
rect 4629 6817 4663 6851
rect 4663 6817 4672 6851
rect 4620 6808 4672 6817
rect 4712 6851 4764 6860
rect 4712 6817 4721 6851
rect 4721 6817 4755 6851
rect 4755 6817 4764 6851
rect 4712 6808 4764 6817
rect 4896 6808 4948 6860
rect 5172 6808 5224 6860
rect 5448 6740 5500 6792
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 6092 6851 6144 6860
rect 6092 6817 6101 6851
rect 6101 6817 6135 6851
rect 6135 6817 6144 6851
rect 6092 6808 6144 6817
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8576 6944 8628 6996
rect 11244 6944 11296 6996
rect 8852 6876 8904 6928
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 5908 6740 5960 6792
rect 6828 6740 6880 6792
rect 6920 6783 6972 6792
rect 6920 6749 6929 6783
rect 6929 6749 6963 6783
rect 6963 6749 6972 6783
rect 6920 6740 6972 6749
rect 7012 6740 7064 6792
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 8852 6740 8904 6792
rect 4160 6672 4212 6724
rect 4528 6672 4580 6724
rect 4804 6672 4856 6724
rect 8484 6672 8536 6724
rect 9772 6851 9824 6860
rect 9772 6817 9781 6851
rect 9781 6817 9815 6851
rect 9815 6817 9824 6851
rect 9772 6808 9824 6817
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 11060 6740 11112 6792
rect 4620 6604 4672 6656
rect 5264 6604 5316 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 8760 6604 8812 6613
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 9772 6604 9824 6656
rect 3662 6502 3714 6554
rect 3726 6502 3778 6554
rect 3790 6502 3842 6554
rect 3854 6502 3906 6554
rect 3918 6502 3970 6554
rect 10062 6502 10114 6554
rect 10126 6502 10178 6554
rect 10190 6502 10242 6554
rect 10254 6502 10306 6554
rect 10318 6502 10370 6554
rect 480 6400 532 6452
rect 1032 6239 1084 6248
rect 1032 6205 1041 6239
rect 1041 6205 1075 6239
rect 1075 6205 1084 6239
rect 1032 6196 1084 6205
rect 1492 6128 1544 6180
rect 2320 6400 2372 6452
rect 4528 6400 4580 6452
rect 4712 6400 4764 6452
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 6092 6400 6144 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7012 6443 7064 6452
rect 7012 6409 7021 6443
rect 7021 6409 7055 6443
rect 7055 6409 7064 6443
rect 7012 6400 7064 6409
rect 7196 6443 7248 6452
rect 7196 6409 7205 6443
rect 7205 6409 7239 6443
rect 7239 6409 7248 6443
rect 7196 6400 7248 6409
rect 7840 6400 7892 6452
rect 10140 6400 10192 6452
rect 3516 6307 3568 6316
rect 3516 6273 3525 6307
rect 3525 6273 3559 6307
rect 3559 6273 3568 6307
rect 3516 6264 3568 6273
rect 2872 6196 2924 6248
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 3608 6196 3660 6248
rect 5264 6332 5316 6384
rect 4436 6239 4488 6248
rect 4436 6205 4445 6239
rect 4445 6205 4479 6239
rect 4479 6205 4488 6239
rect 4436 6196 4488 6205
rect 5540 6196 5592 6248
rect 5908 6196 5960 6248
rect 6000 6196 6052 6248
rect 6552 6196 6604 6248
rect 11152 6400 11204 6452
rect 7012 6196 7064 6248
rect 7196 6239 7248 6248
rect 7196 6205 7205 6239
rect 7205 6205 7239 6239
rect 7239 6205 7248 6239
rect 7196 6196 7248 6205
rect 7288 6196 7340 6248
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 10324 6307 10376 6316
rect 10324 6273 10333 6307
rect 10333 6273 10367 6307
rect 10367 6273 10376 6307
rect 10324 6264 10376 6273
rect 9956 6196 10008 6248
rect 10416 6128 10468 6180
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 2688 6060 2740 6112
rect 3608 6060 3660 6112
rect 4252 6060 4304 6112
rect 4436 6060 4488 6112
rect 4804 6060 4856 6112
rect 5172 6060 5224 6112
rect 9588 6060 9640 6112
rect 10324 6060 10376 6112
rect 4322 5958 4374 6010
rect 4386 5958 4438 6010
rect 4450 5958 4502 6010
rect 4514 5958 4566 6010
rect 4578 5958 4630 6010
rect 10722 5958 10774 6010
rect 10786 5958 10838 6010
rect 10850 5958 10902 6010
rect 10914 5958 10966 6010
rect 10978 5958 11030 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 2320 5856 2372 5908
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 2688 5831 2740 5840
rect 2688 5797 2697 5831
rect 2697 5797 2731 5831
rect 2731 5797 2740 5831
rect 2688 5788 2740 5797
rect 2412 5720 2464 5772
rect 3148 5788 3200 5840
rect 3516 5899 3568 5908
rect 3516 5865 3525 5899
rect 3525 5865 3559 5899
rect 3559 5865 3568 5899
rect 3516 5856 3568 5865
rect 3608 5856 3660 5908
rect 5172 5856 5224 5908
rect 4068 5788 4120 5840
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 10416 5856 10468 5908
rect 10140 5831 10192 5840
rect 10140 5797 10149 5831
rect 10149 5797 10183 5831
rect 10183 5797 10192 5831
rect 10140 5788 10192 5797
rect 10324 5831 10376 5840
rect 10324 5797 10333 5831
rect 10333 5797 10367 5831
rect 10367 5797 10376 5831
rect 10324 5788 10376 5797
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3424 5720 3476 5729
rect 3056 5652 3108 5704
rect 2228 5584 2280 5636
rect 3700 5763 3752 5772
rect 3700 5729 3709 5763
rect 3709 5729 3743 5763
rect 3743 5729 3752 5763
rect 3700 5720 3752 5729
rect 9128 5720 9180 5772
rect 8024 5652 8076 5704
rect 8852 5652 8904 5704
rect 9496 5652 9548 5704
rect 9680 5652 9732 5704
rect 9864 5652 9916 5704
rect 2320 5516 2372 5568
rect 2872 5516 2924 5568
rect 3240 5516 3292 5568
rect 9864 5516 9916 5568
rect 10232 5516 10284 5568
rect 3662 5414 3714 5466
rect 3726 5414 3778 5466
rect 3790 5414 3842 5466
rect 3854 5414 3906 5466
rect 3918 5414 3970 5466
rect 10062 5414 10114 5466
rect 10126 5414 10178 5466
rect 10190 5414 10242 5466
rect 10254 5414 10306 5466
rect 10318 5414 10370 5466
rect 2780 5355 2832 5364
rect 2780 5321 2789 5355
rect 2789 5321 2823 5355
rect 2823 5321 2832 5355
rect 2780 5312 2832 5321
rect 4160 5355 4212 5364
rect 4160 5321 4169 5355
rect 4169 5321 4203 5355
rect 4203 5321 4212 5355
rect 4160 5312 4212 5321
rect 4712 5355 4764 5364
rect 4712 5321 4721 5355
rect 4721 5321 4755 5355
rect 4755 5321 4764 5355
rect 4712 5312 4764 5321
rect 5172 5355 5224 5364
rect 5172 5321 5181 5355
rect 5181 5321 5215 5355
rect 5215 5321 5224 5355
rect 5172 5312 5224 5321
rect 2320 5151 2372 5160
rect 2320 5117 2329 5151
rect 2329 5117 2363 5151
rect 2363 5117 2372 5151
rect 2320 5108 2372 5117
rect 2964 5244 3016 5296
rect 4252 5244 4304 5296
rect 3700 5219 3752 5228
rect 3700 5185 3709 5219
rect 3709 5185 3743 5219
rect 3743 5185 3752 5219
rect 3700 5176 3752 5185
rect 3424 5108 3476 5160
rect 4804 5244 4856 5296
rect 5264 5244 5316 5296
rect 11612 5312 11664 5364
rect 12164 5312 12216 5364
rect 4804 5108 4856 5160
rect 3332 5040 3384 5092
rect 4988 5108 5040 5160
rect 5448 5108 5500 5160
rect 7656 5244 7708 5296
rect 5724 5108 5776 5160
rect 6000 5108 6052 5160
rect 6828 5108 6880 5160
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 8852 5244 8904 5296
rect 8760 5176 8812 5228
rect 11336 5176 11388 5228
rect 12256 5176 12308 5228
rect 7288 5151 7340 5160
rect 7288 5117 7297 5151
rect 7297 5117 7331 5151
rect 7331 5117 7340 5151
rect 7288 5108 7340 5117
rect 7380 5151 7432 5160
rect 7380 5117 7389 5151
rect 7389 5117 7423 5151
rect 7423 5117 7432 5151
rect 7380 5108 7432 5117
rect 7472 5151 7524 5160
rect 7472 5117 7481 5151
rect 7481 5117 7515 5151
rect 7515 5117 7524 5151
rect 7472 5108 7524 5117
rect 7840 5151 7892 5160
rect 7840 5117 7849 5151
rect 7849 5117 7883 5151
rect 7883 5117 7892 5151
rect 7840 5108 7892 5117
rect 9312 5151 9364 5160
rect 3148 4972 3200 5024
rect 4252 4972 4304 5024
rect 5264 5040 5316 5092
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 5908 5083 5960 5092
rect 5908 5049 5917 5083
rect 5917 5049 5951 5083
rect 5951 5049 5960 5083
rect 5908 5040 5960 5049
rect 7104 4972 7156 5024
rect 8300 5040 8352 5092
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 11060 5108 11112 5160
rect 11428 5151 11480 5160
rect 11428 5117 11437 5151
rect 11437 5117 11471 5151
rect 11471 5117 11480 5151
rect 11428 5108 11480 5117
rect 9036 5083 9088 5092
rect 9036 5049 9045 5083
rect 9045 5049 9079 5083
rect 9079 5049 9088 5083
rect 9036 5040 9088 5049
rect 11520 5083 11572 5092
rect 11520 5049 11529 5083
rect 11529 5049 11563 5083
rect 11563 5049 11572 5083
rect 11520 5040 11572 5049
rect 12256 5040 12308 5092
rect 8668 4972 8720 5024
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 11244 4972 11296 5024
rect 4322 4870 4374 4922
rect 4386 4870 4438 4922
rect 4450 4870 4502 4922
rect 4514 4870 4566 4922
rect 4578 4870 4630 4922
rect 10722 4870 10774 4922
rect 10786 4870 10838 4922
rect 10850 4870 10902 4922
rect 10914 4870 10966 4922
rect 10978 4870 11030 4922
rect 3148 4811 3200 4820
rect 3148 4777 3157 4811
rect 3157 4777 3191 4811
rect 3191 4777 3200 4811
rect 3148 4768 3200 4777
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3700 4768 3752 4820
rect 2872 4700 2924 4752
rect 3332 4632 3384 4684
rect 6460 4768 6512 4820
rect 7840 4768 7892 4820
rect 5724 4700 5776 4752
rect 6092 4700 6144 4752
rect 8852 4768 8904 4820
rect 9404 4768 9456 4820
rect 11612 4768 11664 4820
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5448 4632 5500 4684
rect 2964 4564 3016 4616
rect 5816 4564 5868 4616
rect 5264 4496 5316 4548
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 6828 4675 6880 4684
rect 6828 4641 6837 4675
rect 6837 4641 6871 4675
rect 6871 4641 6880 4675
rect 6828 4632 6880 4641
rect 8576 4700 8628 4752
rect 9220 4700 9272 4752
rect 9312 4700 9364 4752
rect 9680 4700 9732 4752
rect 11520 4700 11572 4752
rect 8668 4675 8720 4684
rect 8668 4641 8677 4675
rect 8677 4641 8711 4675
rect 8711 4641 8720 4675
rect 8668 4632 8720 4641
rect 9496 4632 9548 4684
rect 7932 4564 7984 4616
rect 8300 4564 8352 4616
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 7472 4428 7524 4480
rect 11244 4632 11296 4684
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 12348 4632 12400 4684
rect 11152 4564 11204 4616
rect 11428 4564 11480 4616
rect 8760 4428 8812 4480
rect 9680 4428 9732 4480
rect 10416 4428 10468 4480
rect 11060 4428 11112 4480
rect 11704 4428 11756 4480
rect 3662 4326 3714 4378
rect 3726 4326 3778 4378
rect 3790 4326 3842 4378
rect 3854 4326 3906 4378
rect 3918 4326 3970 4378
rect 10062 4326 10114 4378
rect 10126 4326 10178 4378
rect 10190 4326 10242 4378
rect 10254 4326 10306 4378
rect 10318 4326 10370 4378
rect 2872 4224 2924 4276
rect 4252 4224 4304 4276
rect 4988 4224 5040 4276
rect 5816 4267 5868 4276
rect 5816 4233 5825 4267
rect 5825 4233 5859 4267
rect 5859 4233 5868 4267
rect 5816 4224 5868 4233
rect 7380 4224 7432 4276
rect 8116 4267 8168 4276
rect 8116 4233 8125 4267
rect 8125 4233 8159 4267
rect 8159 4233 8168 4267
rect 8116 4224 8168 4233
rect 8392 4224 8444 4276
rect 8484 4224 8536 4276
rect 9036 4224 9088 4276
rect 2688 4088 2740 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 1400 4063 1452 4072
rect 1400 4029 1409 4063
rect 1409 4029 1443 4063
rect 1443 4029 1452 4063
rect 1400 4020 1452 4029
rect 6552 4156 6604 4208
rect 5172 4088 5224 4140
rect 5264 4088 5316 4140
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 9772 4156 9824 4208
rect 12348 4224 12400 4276
rect 8760 4088 8812 4140
rect 1676 3995 1728 4004
rect 1676 3961 1710 3995
rect 1710 3961 1728 3995
rect 1676 3952 1728 3961
rect 4988 4020 5040 4072
rect 5448 4020 5500 4072
rect 6092 4020 6144 4072
rect 4436 3952 4488 4004
rect 7472 4020 7524 4072
rect 7840 4063 7892 4072
rect 7840 4029 7849 4063
rect 7849 4029 7883 4063
rect 7883 4029 7892 4063
rect 7840 4020 7892 4029
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 8944 4020 8996 4072
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 10692 4088 10744 4140
rect 11152 4063 11204 4072
rect 11152 4029 11186 4063
rect 11186 4029 11204 4063
rect 11152 4020 11204 4029
rect 9680 3952 9732 4004
rect 4068 3884 4120 3936
rect 4322 3782 4374 3834
rect 4386 3782 4438 3834
rect 4450 3782 4502 3834
rect 4514 3782 4566 3834
rect 4578 3782 4630 3834
rect 10722 3782 10774 3834
rect 10786 3782 10838 3834
rect 10850 3782 10902 3834
rect 10914 3782 10966 3834
rect 10978 3782 11030 3834
rect 1676 3723 1728 3732
rect 1676 3689 1685 3723
rect 1685 3689 1719 3723
rect 1719 3689 1728 3723
rect 1676 3680 1728 3689
rect 2412 3680 2464 3732
rect 2688 3723 2740 3732
rect 2688 3689 2697 3723
rect 2697 3689 2731 3723
rect 2731 3689 2740 3723
rect 2688 3680 2740 3689
rect 4160 3680 4212 3732
rect 5264 3723 5316 3732
rect 5264 3689 5273 3723
rect 5273 3689 5307 3723
rect 5307 3689 5316 3723
rect 5264 3680 5316 3689
rect 5448 3680 5500 3732
rect 6828 3680 6880 3732
rect 7012 3680 7064 3732
rect 8576 3723 8628 3732
rect 8576 3689 8585 3723
rect 8585 3689 8619 3723
rect 8619 3689 8628 3723
rect 8576 3680 8628 3689
rect 9220 3680 9272 3732
rect 2872 3612 2924 3664
rect 1860 3476 1912 3528
rect 2412 3476 2464 3528
rect 3240 3544 3292 3596
rect 3424 3476 3476 3528
rect 3516 3476 3568 3528
rect 4068 3476 4120 3528
rect 4712 3587 4764 3596
rect 4712 3553 4721 3587
rect 4721 3553 4755 3587
rect 4755 3553 4764 3587
rect 4712 3544 4764 3553
rect 4988 3612 5040 3664
rect 6736 3612 6788 3664
rect 5172 3544 5224 3596
rect 5356 3544 5408 3596
rect 6828 3587 6880 3596
rect 6828 3553 6837 3587
rect 6837 3553 6871 3587
rect 6871 3553 6880 3587
rect 6828 3544 6880 3553
rect 7380 3544 7432 3596
rect 7840 3612 7892 3664
rect 7472 3476 7524 3528
rect 8484 3587 8536 3596
rect 8484 3553 8493 3587
rect 8493 3553 8527 3587
rect 8527 3553 8536 3587
rect 8484 3544 8536 3553
rect 8760 3587 8812 3596
rect 8760 3553 8769 3587
rect 8769 3553 8803 3587
rect 8803 3553 8812 3587
rect 8760 3544 8812 3553
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9036 3544 9088 3596
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9496 3544 9548 3596
rect 9772 3680 9824 3732
rect 11704 3612 11756 3664
rect 9772 3587 9824 3596
rect 9772 3553 9782 3587
rect 9782 3553 9816 3587
rect 9816 3553 9824 3587
rect 9772 3544 9824 3553
rect 10416 3544 10468 3596
rect 11244 3544 11296 3596
rect 11520 3544 11572 3596
rect 2688 3408 2740 3460
rect 9680 3408 9732 3460
rect 1492 3340 1544 3392
rect 2044 3340 2096 3392
rect 4896 3340 4948 3392
rect 9588 3340 9640 3392
rect 9772 3340 9824 3392
rect 11336 3383 11388 3392
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 11520 3383 11572 3392
rect 11520 3349 11529 3383
rect 11529 3349 11563 3383
rect 11563 3349 11572 3383
rect 11520 3340 11572 3349
rect 3662 3238 3714 3290
rect 3726 3238 3778 3290
rect 3790 3238 3842 3290
rect 3854 3238 3906 3290
rect 3918 3238 3970 3290
rect 10062 3238 10114 3290
rect 10126 3238 10178 3290
rect 10190 3238 10242 3290
rect 10254 3238 10306 3290
rect 10318 3238 10370 3290
rect 1492 3136 1544 3188
rect 2504 3136 2556 3188
rect 4712 3136 4764 3188
rect 12256 3179 12308 3188
rect 12256 3145 12265 3179
rect 12265 3145 12299 3179
rect 12299 3145 12308 3179
rect 12256 3136 12308 3145
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2320 3000 2372 3052
rect 3148 3000 3200 3052
rect 10600 3000 10652 3052
rect 2504 2975 2556 2984
rect 2504 2941 2513 2975
rect 2513 2941 2547 2975
rect 2547 2941 2556 2975
rect 2504 2932 2556 2941
rect 3240 2932 3292 2984
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 6368 2932 6420 2984
rect 6644 2932 6696 2984
rect 11520 2932 11572 2984
rect 2872 2864 2924 2916
rect 3424 2864 3476 2916
rect 4252 2864 4304 2916
rect 6736 2796 6788 2848
rect 4322 2694 4374 2746
rect 4386 2694 4438 2746
rect 4450 2694 4502 2746
rect 4514 2694 4566 2746
rect 4578 2694 4630 2746
rect 10722 2694 10774 2746
rect 10786 2694 10838 2746
rect 10850 2694 10902 2746
rect 10914 2694 10966 2746
rect 10978 2694 11030 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 7288 2592 7340 2644
rect 9496 2592 9548 2644
rect 10508 2592 10560 2644
rect 4252 2524 4304 2576
rect 7656 2567 7708 2576
rect 7656 2533 7665 2567
rect 7665 2533 7699 2567
rect 7699 2533 7708 2567
rect 7656 2524 7708 2533
rect 8760 2524 8812 2576
rect 9772 2524 9824 2576
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 3148 2499 3200 2508
rect 3148 2465 3157 2499
rect 3157 2465 3191 2499
rect 3191 2465 3200 2499
rect 3148 2456 3200 2465
rect 5448 2456 5500 2508
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6460 2499 6512 2508
rect 6460 2465 6469 2499
rect 6469 2465 6503 2499
rect 6503 2465 6512 2499
rect 6460 2456 6512 2465
rect 2228 2388 2280 2440
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7288 2456 7340 2508
rect 8208 2456 8260 2508
rect 8576 2456 8628 2508
rect 7748 2431 7800 2440
rect 7748 2397 7757 2431
rect 7757 2397 7791 2431
rect 7791 2397 7800 2431
rect 7748 2388 7800 2397
rect 8116 2388 8168 2440
rect 8944 2456 8996 2508
rect 9680 2456 9732 2508
rect 10692 2524 10744 2576
rect 2688 2252 2740 2304
rect 6276 2252 6328 2304
rect 8484 2320 8536 2372
rect 9128 2320 9180 2372
rect 10416 2456 10468 2508
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10508 2388 10560 2440
rect 7196 2295 7248 2304
rect 7196 2261 7205 2295
rect 7205 2261 7239 2295
rect 7239 2261 7248 2295
rect 7196 2252 7248 2261
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 10784 2252 10836 2304
rect 3662 2150 3714 2202
rect 3726 2150 3778 2202
rect 3790 2150 3842 2202
rect 3854 2150 3906 2202
rect 3918 2150 3970 2202
rect 10062 2150 10114 2202
rect 10126 2150 10178 2202
rect 10190 2150 10242 2202
rect 10254 2150 10306 2202
rect 10318 2150 10370 2202
rect 2504 2048 2556 2100
rect 3332 2048 3384 2100
rect 5172 2048 5224 2100
rect 2596 2023 2648 2032
rect 2596 1989 2605 2023
rect 2605 1989 2639 2023
rect 2639 1989 2648 2023
rect 2596 1980 2648 1989
rect 2044 1912 2096 1964
rect 2504 1955 2556 1964
rect 2504 1921 2513 1955
rect 2513 1921 2547 1955
rect 2547 1921 2556 1955
rect 2504 1912 2556 1921
rect 3516 1912 3568 1964
rect 4160 1912 4212 1964
rect 5540 2023 5592 2032
rect 5540 1989 5549 2023
rect 5549 1989 5583 2023
rect 5583 1989 5592 2023
rect 5540 1980 5592 1989
rect 7472 2048 7524 2100
rect 7748 2048 7800 2100
rect 10416 2048 10468 2100
rect 9404 1980 9456 2032
rect 2688 1844 2740 1896
rect 3424 1887 3476 1896
rect 3424 1853 3433 1887
rect 3433 1853 3467 1887
rect 3467 1853 3476 1887
rect 3424 1844 3476 1853
rect 3608 1887 3660 1896
rect 3608 1853 3617 1887
rect 3617 1853 3651 1887
rect 3651 1853 3660 1887
rect 3608 1844 3660 1853
rect 3792 1887 3844 1896
rect 3792 1853 3801 1887
rect 3801 1853 3835 1887
rect 3835 1853 3844 1887
rect 3792 1844 3844 1853
rect 5172 1887 5224 1896
rect 5172 1853 5181 1887
rect 5181 1853 5215 1887
rect 5215 1853 5224 1887
rect 5172 1844 5224 1853
rect 5816 1887 5868 1896
rect 5816 1853 5825 1887
rect 5825 1853 5859 1887
rect 5859 1853 5868 1887
rect 5816 1844 5868 1853
rect 6368 1844 6420 1896
rect 5908 1776 5960 1828
rect 3332 1708 3384 1760
rect 4896 1708 4948 1760
rect 6644 1844 6696 1896
rect 10600 1912 10652 1964
rect 9496 1844 9548 1896
rect 7196 1776 7248 1828
rect 7472 1776 7524 1828
rect 8484 1776 8536 1828
rect 8668 1819 8720 1828
rect 8668 1785 8702 1819
rect 8702 1785 8720 1819
rect 8668 1776 8720 1785
rect 9680 1776 9732 1828
rect 9956 1776 10008 1828
rect 10416 1844 10468 1896
rect 10784 1887 10836 1896
rect 10784 1853 10793 1887
rect 10793 1853 10827 1887
rect 10827 1853 10836 1887
rect 10784 1844 10836 1853
rect 11244 1887 11296 1896
rect 11244 1853 11253 1887
rect 11253 1853 11287 1887
rect 11287 1853 11296 1887
rect 11244 1844 11296 1853
rect 6828 1708 6880 1760
rect 10416 1708 10468 1760
rect 4322 1606 4374 1658
rect 4386 1606 4438 1658
rect 4450 1606 4502 1658
rect 4514 1606 4566 1658
rect 4578 1606 4630 1658
rect 10722 1606 10774 1658
rect 10786 1606 10838 1658
rect 10850 1606 10902 1658
rect 10914 1606 10966 1658
rect 10978 1606 11030 1658
rect 3792 1504 3844 1556
rect 5172 1504 5224 1556
rect 7288 1504 7340 1556
rect 7564 1504 7616 1556
rect 8116 1547 8168 1556
rect 8116 1513 8125 1547
rect 8125 1513 8159 1547
rect 8159 1513 8168 1547
rect 8116 1504 8168 1513
rect 8300 1504 8352 1556
rect 8576 1547 8628 1556
rect 8576 1513 8585 1547
rect 8585 1513 8619 1547
rect 8619 1513 8628 1547
rect 8576 1504 8628 1513
rect 2596 1436 2648 1488
rect 3516 1368 3568 1420
rect 4252 1411 4304 1420
rect 4252 1377 4261 1411
rect 4261 1377 4295 1411
rect 4295 1377 4304 1411
rect 4252 1368 4304 1377
rect 4896 1411 4948 1420
rect 4896 1377 4905 1411
rect 4905 1377 4939 1411
rect 4939 1377 4948 1411
rect 4896 1368 4948 1377
rect 5448 1401 5500 1420
rect 5448 1368 5457 1401
rect 5457 1368 5491 1401
rect 5491 1368 5500 1401
rect 6552 1436 6604 1488
rect 1400 1300 1452 1352
rect 3608 1232 3660 1284
rect 4068 1300 4120 1352
rect 6460 1368 6512 1420
rect 4804 1164 4856 1216
rect 8944 1436 8996 1488
rect 9496 1504 9548 1556
rect 10416 1547 10468 1556
rect 10416 1513 10425 1547
rect 10425 1513 10459 1547
rect 10459 1513 10468 1547
rect 10416 1504 10468 1513
rect 10600 1547 10652 1556
rect 10600 1513 10609 1547
rect 10609 1513 10643 1547
rect 10643 1513 10652 1547
rect 10600 1504 10652 1513
rect 6736 1411 6788 1420
rect 6736 1377 6745 1411
rect 6745 1377 6779 1411
rect 6779 1377 6788 1411
rect 6736 1368 6788 1377
rect 7564 1411 7616 1420
rect 7564 1377 7573 1411
rect 7573 1377 7607 1411
rect 7607 1377 7616 1411
rect 7564 1368 7616 1377
rect 7656 1411 7708 1420
rect 7656 1377 7665 1411
rect 7665 1377 7699 1411
rect 7699 1377 7708 1411
rect 7656 1368 7708 1377
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 7472 1300 7524 1352
rect 6092 1164 6144 1216
rect 7012 1207 7064 1216
rect 7012 1173 7021 1207
rect 7021 1173 7055 1207
rect 7055 1173 7064 1207
rect 7012 1164 7064 1173
rect 8208 1411 8260 1420
rect 8208 1377 8217 1411
rect 8217 1377 8251 1411
rect 8251 1377 8260 1411
rect 8208 1368 8260 1377
rect 8484 1368 8536 1420
rect 9404 1368 9456 1420
rect 9588 1411 9640 1420
rect 9588 1377 9597 1411
rect 9597 1377 9631 1411
rect 9631 1377 9640 1411
rect 9588 1368 9640 1377
rect 9772 1368 9824 1420
rect 8392 1300 8444 1352
rect 8300 1232 8352 1284
rect 9036 1300 9088 1352
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 10508 1411 10560 1420
rect 10508 1377 10517 1411
rect 10517 1377 10551 1411
rect 10551 1377 10560 1411
rect 10508 1368 10560 1377
rect 8760 1275 8812 1284
rect 8760 1241 8769 1275
rect 8769 1241 8803 1275
rect 8803 1241 8812 1275
rect 8760 1232 8812 1241
rect 9312 1232 9364 1284
rect 11428 1232 11480 1284
rect 9864 1207 9916 1216
rect 9864 1173 9873 1207
rect 9873 1173 9907 1207
rect 9907 1173 9916 1207
rect 9864 1164 9916 1173
rect 3662 1062 3714 1114
rect 3726 1062 3778 1114
rect 3790 1062 3842 1114
rect 3854 1062 3906 1114
rect 3918 1062 3970 1114
rect 10062 1062 10114 1114
rect 10126 1062 10178 1114
rect 10190 1062 10242 1114
rect 10254 1062 10306 1114
rect 10318 1062 10370 1114
rect 3516 960 3568 1012
rect 6460 960 6512 1012
rect 6644 1003 6696 1012
rect 6644 969 6653 1003
rect 6653 969 6687 1003
rect 6687 969 6696 1003
rect 6644 960 6696 969
rect 9588 1003 9640 1012
rect 9588 969 9597 1003
rect 9597 969 9631 1003
rect 9631 969 9640 1003
rect 9588 960 9640 969
rect 3424 824 3476 876
rect 2780 756 2832 808
rect 5540 824 5592 876
rect 3332 688 3384 740
rect 3976 799 4028 808
rect 3976 765 3985 799
rect 3985 765 4019 799
rect 4019 765 4028 799
rect 3976 756 4028 765
rect 4068 688 4120 740
rect 6092 799 6144 808
rect 6092 765 6101 799
rect 6101 765 6135 799
rect 6135 765 6144 799
rect 6092 756 6144 765
rect 6276 799 6328 808
rect 6276 765 6285 799
rect 6285 765 6319 799
rect 6319 765 6328 799
rect 6276 756 6328 765
rect 7472 756 7524 808
rect 9496 756 9548 808
rect 10416 756 10468 808
rect 3976 620 4028 672
rect 4322 518 4374 570
rect 4386 518 4438 570
rect 4450 518 4502 570
rect 4514 518 4566 570
rect 4578 518 4630 570
rect 10722 518 10774 570
rect 10786 518 10838 570
rect 10850 518 10902 570
rect 10914 518 10966 570
rect 10978 518 11030 570
<< metal2 >>
rect 1674 43500 1730 43900
rect 2226 43616 2282 43900
rect 2226 43500 2282 43560
rect 2778 43500 2834 43900
rect 4434 43500 4490 43900
rect 4986 43616 5042 43900
rect 4986 43500 5042 43560
rect 5538 43500 5594 43900
rect 6090 43616 6146 43900
rect 6090 43500 6146 43560
rect 6642 43500 6698 43900
rect 7194 43602 7250 43900
rect 7746 43616 7802 43900
rect 7194 43574 7512 43602
rect 7194 43500 7250 43574
rect 20 42764 72 42770
rect 20 42706 72 42712
rect 1308 42764 1360 42770
rect 1308 42706 1360 42712
rect 1492 42764 1544 42770
rect 1492 42706 1544 42712
rect 32 33998 60 42706
rect 846 42664 902 42673
rect 846 42599 902 42608
rect 860 42158 888 42599
rect 940 42560 992 42566
rect 940 42502 992 42508
rect 848 42152 900 42158
rect 848 42094 900 42100
rect 952 41449 980 42502
rect 1032 42152 1084 42158
rect 1032 42094 1084 42100
rect 1044 41818 1072 42094
rect 1216 42084 1268 42090
rect 1216 42026 1268 42032
rect 1032 41812 1084 41818
rect 1032 41754 1084 41760
rect 1032 41676 1084 41682
rect 1084 41636 1164 41664
rect 1032 41618 1084 41624
rect 938 41440 994 41449
rect 938 41375 994 41384
rect 386 41168 442 41177
rect 1136 41138 1164 41636
rect 1228 41274 1256 42026
rect 1320 41682 1348 42706
rect 1308 41676 1360 41682
rect 1308 41618 1360 41624
rect 1216 41268 1268 41274
rect 1216 41210 1268 41216
rect 1320 41138 1348 41618
rect 1504 41546 1532 42706
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1492 41540 1544 41546
rect 1492 41482 1544 41488
rect 386 41103 442 41112
rect 1124 41132 1176 41138
rect 400 38593 428 41103
rect 1124 41074 1176 41080
rect 1308 41132 1360 41138
rect 1308 41074 1360 41080
rect 570 40896 626 40905
rect 570 40831 626 40840
rect 478 39944 534 39953
rect 478 39879 534 39888
rect 492 38894 520 39879
rect 480 38888 532 38894
rect 480 38830 532 38836
rect 480 38752 532 38758
rect 480 38694 532 38700
rect 386 38584 442 38593
rect 386 38519 442 38528
rect 296 38480 348 38486
rect 296 38422 348 38428
rect 204 36712 256 36718
rect 204 36654 256 36660
rect 112 36236 164 36242
rect 112 36178 164 36184
rect 20 33992 72 33998
rect 20 33934 72 33940
rect 20 30592 72 30598
rect 20 30534 72 30540
rect 32 20534 60 30534
rect 124 24818 152 36178
rect 216 27713 244 36654
rect 308 36242 336 38422
rect 388 36576 440 36582
rect 388 36518 440 36524
rect 296 36236 348 36242
rect 296 36178 348 36184
rect 400 34649 428 36518
rect 492 34921 520 38694
rect 478 34912 534 34921
rect 478 34847 534 34856
rect 584 34762 612 40831
rect 846 40488 902 40497
rect 846 40423 902 40432
rect 664 39432 716 39438
rect 664 39374 716 39380
rect 754 39400 810 39409
rect 676 35290 704 39374
rect 754 39335 810 39344
rect 768 36174 796 39335
rect 860 37466 888 40423
rect 1032 39976 1084 39982
rect 1032 39918 1084 39924
rect 940 39840 992 39846
rect 940 39782 992 39788
rect 952 39545 980 39782
rect 938 39536 994 39545
rect 938 39471 994 39480
rect 940 39296 992 39302
rect 938 39264 940 39273
rect 992 39264 994 39273
rect 938 39199 994 39208
rect 938 39128 994 39137
rect 938 39063 994 39072
rect 952 39030 980 39063
rect 940 39024 992 39030
rect 940 38966 992 38972
rect 940 38344 992 38350
rect 940 38286 992 38292
rect 848 37460 900 37466
rect 848 37402 900 37408
rect 952 36825 980 38286
rect 1044 38010 1072 39918
rect 1136 39846 1164 41074
rect 1504 41070 1532 41482
rect 1492 41064 1544 41070
rect 1492 41006 1544 41012
rect 1400 40996 1452 41002
rect 1400 40938 1452 40944
rect 1412 40730 1440 40938
rect 1216 40724 1268 40730
rect 1216 40666 1268 40672
rect 1400 40724 1452 40730
rect 1400 40666 1452 40672
rect 1228 40633 1256 40666
rect 1214 40624 1270 40633
rect 1214 40559 1270 40568
rect 1308 40588 1360 40594
rect 1308 40530 1360 40536
rect 1216 39976 1268 39982
rect 1216 39918 1268 39924
rect 1124 39840 1176 39846
rect 1124 39782 1176 39788
rect 1136 39681 1164 39782
rect 1122 39672 1178 39681
rect 1122 39607 1178 39616
rect 1136 38758 1164 39607
rect 1228 39001 1256 39918
rect 1214 38992 1270 39001
rect 1214 38927 1270 38936
rect 1320 38842 1348 40530
rect 1492 40452 1544 40458
rect 1492 40394 1544 40400
rect 1398 40080 1454 40089
rect 1398 40015 1454 40024
rect 1412 39370 1440 40015
rect 1504 39846 1532 40394
rect 1492 39840 1544 39846
rect 1492 39782 1544 39788
rect 1492 39500 1544 39506
rect 1492 39442 1544 39448
rect 1400 39364 1452 39370
rect 1400 39306 1452 39312
rect 1400 38888 1452 38894
rect 1228 38814 1348 38842
rect 1398 38856 1400 38865
rect 1452 38856 1454 38865
rect 1124 38752 1176 38758
rect 1124 38694 1176 38700
rect 1032 38004 1084 38010
rect 1032 37946 1084 37952
rect 1030 37904 1086 37913
rect 1030 37839 1086 37848
rect 1044 37330 1072 37839
rect 1124 37732 1176 37738
rect 1124 37674 1176 37680
rect 1136 37641 1164 37674
rect 1228 37670 1256 38814
rect 1398 38791 1454 38800
rect 1504 38706 1532 39442
rect 1320 38678 1532 38706
rect 1216 37664 1268 37670
rect 1122 37632 1178 37641
rect 1216 37606 1268 37612
rect 1122 37567 1178 37576
rect 1032 37324 1084 37330
rect 1032 37266 1084 37272
rect 1216 37324 1268 37330
rect 1216 37266 1268 37272
rect 1122 36952 1178 36961
rect 1122 36887 1178 36896
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1136 36718 1164 36887
rect 1228 36825 1256 37266
rect 1214 36816 1270 36825
rect 1214 36751 1270 36760
rect 1124 36712 1176 36718
rect 1124 36654 1176 36660
rect 1122 36544 1178 36553
rect 1122 36479 1178 36488
rect 846 36272 902 36281
rect 846 36207 902 36216
rect 1032 36236 1084 36242
rect 756 36168 808 36174
rect 756 36110 808 36116
rect 664 35284 716 35290
rect 664 35226 716 35232
rect 492 34734 612 34762
rect 386 34640 442 34649
rect 386 34575 442 34584
rect 388 34536 440 34542
rect 388 34478 440 34484
rect 400 31890 428 34478
rect 388 31884 440 31890
rect 388 31826 440 31832
rect 386 31104 442 31113
rect 386 31039 442 31048
rect 400 29510 428 31039
rect 492 29850 520 34734
rect 572 34400 624 34406
rect 572 34342 624 34348
rect 584 32026 612 34342
rect 768 32065 796 36110
rect 860 34134 888 36207
rect 1032 36178 1084 36184
rect 940 36032 992 36038
rect 940 35974 992 35980
rect 952 34377 980 35974
rect 1044 35834 1072 36178
rect 1032 35828 1084 35834
rect 1032 35770 1084 35776
rect 1030 35592 1086 35601
rect 1030 35527 1086 35536
rect 1044 35154 1072 35527
rect 1136 35290 1164 36479
rect 1124 35284 1176 35290
rect 1124 35226 1176 35232
rect 1228 35170 1256 36751
rect 1032 35148 1084 35154
rect 1032 35090 1084 35096
rect 1136 35142 1256 35170
rect 1136 35034 1164 35142
rect 1044 35006 1164 35034
rect 1216 35080 1268 35086
rect 1216 35022 1268 35028
rect 938 34368 994 34377
rect 938 34303 994 34312
rect 848 34128 900 34134
rect 848 34070 900 34076
rect 1044 34066 1072 35006
rect 1124 34944 1176 34950
rect 1124 34886 1176 34892
rect 1032 34060 1084 34066
rect 1032 34002 1084 34008
rect 848 33992 900 33998
rect 848 33934 900 33940
rect 754 32056 810 32065
rect 572 32020 624 32026
rect 754 31991 810 32000
rect 572 31962 624 31968
rect 860 31958 888 33934
rect 1136 33046 1164 34886
rect 1228 34746 1256 35022
rect 1216 34740 1268 34746
rect 1216 34682 1268 34688
rect 1216 34128 1268 34134
rect 1216 34070 1268 34076
rect 1124 33040 1176 33046
rect 1124 32982 1176 32988
rect 1228 32978 1256 34070
rect 1216 32972 1268 32978
rect 1216 32914 1268 32920
rect 1124 32564 1176 32570
rect 1124 32506 1176 32512
rect 1032 32224 1084 32230
rect 1032 32166 1084 32172
rect 1044 32042 1072 32166
rect 952 32014 1072 32042
rect 848 31952 900 31958
rect 848 31894 900 31900
rect 572 31884 624 31890
rect 572 31826 624 31832
rect 584 30598 612 31826
rect 756 31816 808 31822
rect 662 31784 718 31793
rect 756 31758 808 31764
rect 662 31719 718 31728
rect 572 30592 624 30598
rect 572 30534 624 30540
rect 676 30410 704 31719
rect 584 30382 704 30410
rect 584 30326 612 30382
rect 572 30320 624 30326
rect 572 30262 624 30268
rect 664 30320 716 30326
rect 664 30262 716 30268
rect 480 29844 532 29850
rect 480 29786 532 29792
rect 388 29504 440 29510
rect 388 29446 440 29452
rect 296 28620 348 28626
rect 296 28562 348 28568
rect 202 27704 258 27713
rect 202 27639 258 27648
rect 112 24812 164 24818
rect 112 24754 164 24760
rect 308 22094 336 28562
rect 400 23322 428 29446
rect 480 26852 532 26858
rect 480 26794 532 26800
rect 492 23769 520 26794
rect 584 26058 612 30262
rect 676 27062 704 30262
rect 768 28393 796 31758
rect 860 31385 888 31894
rect 846 31376 902 31385
rect 846 31311 902 31320
rect 952 30870 980 32014
rect 1032 31952 1084 31958
rect 1032 31894 1084 31900
rect 940 30864 992 30870
rect 940 30806 992 30812
rect 848 30592 900 30598
rect 848 30534 900 30540
rect 860 30190 888 30534
rect 848 30184 900 30190
rect 848 30126 900 30132
rect 1044 29714 1072 31894
rect 1136 30326 1164 32506
rect 1216 32360 1268 32366
rect 1216 32302 1268 32308
rect 1228 31890 1256 32302
rect 1216 31884 1268 31890
rect 1216 31826 1268 31832
rect 1228 31793 1256 31826
rect 1214 31784 1270 31793
rect 1214 31719 1270 31728
rect 1216 31680 1268 31686
rect 1216 31622 1268 31628
rect 1124 30320 1176 30326
rect 1124 30262 1176 30268
rect 1124 30116 1176 30122
rect 1124 30058 1176 30064
rect 1032 29708 1084 29714
rect 1032 29650 1084 29656
rect 940 29164 992 29170
rect 940 29106 992 29112
rect 848 28552 900 28558
rect 848 28494 900 28500
rect 754 28384 810 28393
rect 754 28319 810 28328
rect 664 27056 716 27062
rect 664 26998 716 27004
rect 584 26030 796 26058
rect 570 25120 626 25129
rect 570 25055 626 25064
rect 478 23760 534 23769
rect 478 23695 534 23704
rect 388 23316 440 23322
rect 388 23258 440 23264
rect 308 22066 520 22094
rect 386 21992 442 22001
rect 386 21927 442 21936
rect 20 20528 72 20534
rect 20 20470 72 20476
rect 400 12306 428 21927
rect 492 15337 520 22066
rect 478 15328 534 15337
rect 478 15263 534 15272
rect 480 12436 532 12442
rect 480 12378 532 12384
rect 388 12300 440 12306
rect 388 12242 440 12248
rect 386 7168 442 7177
rect 386 7103 442 7112
rect 400 4729 428 7103
rect 492 6458 520 12378
rect 584 12186 612 25055
rect 664 24812 716 24818
rect 664 24754 716 24760
rect 676 22574 704 24754
rect 768 24410 796 26030
rect 756 24404 808 24410
rect 756 24346 808 24352
rect 754 24304 810 24313
rect 754 24239 810 24248
rect 664 22568 716 22574
rect 664 22510 716 22516
rect 676 21894 704 22510
rect 664 21888 716 21894
rect 664 21830 716 21836
rect 664 20596 716 20602
rect 664 20538 716 20544
rect 676 19854 704 20538
rect 768 20466 796 24239
rect 860 23730 888 28494
rect 952 28218 980 29106
rect 1032 29028 1084 29034
rect 1032 28970 1084 28976
rect 1044 28665 1072 28970
rect 1030 28656 1086 28665
rect 1030 28591 1086 28600
rect 1030 28384 1086 28393
rect 1030 28319 1086 28328
rect 940 28212 992 28218
rect 940 28154 992 28160
rect 1044 25906 1072 28319
rect 1136 28121 1164 30058
rect 1122 28112 1178 28121
rect 1122 28047 1178 28056
rect 1032 25900 1084 25906
rect 1032 25842 1084 25848
rect 1032 24676 1084 24682
rect 1032 24618 1084 24624
rect 1124 24676 1176 24682
rect 1124 24618 1176 24624
rect 940 24404 992 24410
rect 940 24346 992 24352
rect 848 23724 900 23730
rect 848 23666 900 23672
rect 952 23662 980 24346
rect 1044 24041 1072 24618
rect 1030 24032 1086 24041
rect 1030 23967 1086 23976
rect 1032 23792 1084 23798
rect 1032 23734 1084 23740
rect 940 23656 992 23662
rect 940 23598 992 23604
rect 940 23180 992 23186
rect 940 23122 992 23128
rect 848 21956 900 21962
rect 848 21898 900 21904
rect 756 20460 808 20466
rect 756 20402 808 20408
rect 664 19848 716 19854
rect 664 19790 716 19796
rect 860 19292 888 21898
rect 952 20058 980 23122
rect 1044 22794 1072 23734
rect 1136 23186 1164 24618
rect 1228 23798 1256 31622
rect 1320 28914 1348 38678
rect 1400 38548 1452 38554
rect 1400 38490 1452 38496
rect 1412 37330 1440 38490
rect 1492 38412 1544 38418
rect 1492 38354 1544 38360
rect 1504 37505 1532 38354
rect 1596 37806 1624 42094
rect 1688 38486 1716 43500
rect 2596 42560 2648 42566
rect 2596 42502 2648 42508
rect 2136 42152 2188 42158
rect 2136 42094 2188 42100
rect 1860 42084 1912 42090
rect 1860 42026 1912 42032
rect 1872 41818 1900 42026
rect 1860 41812 1912 41818
rect 1860 41754 1912 41760
rect 2042 41712 2098 41721
rect 2042 41647 2098 41656
rect 1860 41472 1912 41478
rect 1860 41414 1912 41420
rect 1768 41064 1820 41070
rect 1768 41006 1820 41012
rect 1780 40458 1808 41006
rect 1768 40452 1820 40458
rect 1768 40394 1820 40400
rect 1768 40180 1820 40186
rect 1768 40122 1820 40128
rect 1780 39438 1808 40122
rect 1872 39506 1900 41414
rect 2056 40118 2084 41647
rect 2148 40934 2176 42094
rect 2608 41818 2636 42502
rect 2596 41812 2648 41818
rect 2596 41754 2648 41760
rect 2320 41676 2372 41682
rect 2320 41618 2372 41624
rect 2504 41676 2556 41682
rect 2504 41618 2556 41624
rect 2332 41070 2360 41618
rect 2320 41064 2372 41070
rect 2320 41006 2372 41012
rect 2136 40928 2188 40934
rect 2136 40870 2188 40876
rect 2332 40594 2360 41006
rect 2516 40730 2544 41618
rect 2608 41177 2636 41754
rect 2688 41268 2740 41274
rect 2688 41210 2740 41216
rect 2594 41168 2650 41177
rect 2594 41103 2650 41112
rect 2596 40928 2648 40934
rect 2596 40870 2648 40876
rect 2504 40724 2556 40730
rect 2504 40666 2556 40672
rect 2502 40624 2558 40633
rect 2320 40588 2372 40594
rect 2320 40530 2372 40536
rect 2412 40588 2464 40594
rect 2502 40559 2558 40568
rect 2412 40530 2464 40536
rect 2136 40520 2188 40526
rect 2136 40462 2188 40468
rect 2148 40186 2176 40462
rect 2228 40384 2280 40390
rect 2228 40326 2280 40332
rect 2136 40180 2188 40186
rect 2136 40122 2188 40128
rect 2044 40112 2096 40118
rect 2044 40054 2096 40060
rect 1952 40044 2004 40050
rect 1952 39986 2004 39992
rect 1860 39500 1912 39506
rect 1860 39442 1912 39448
rect 1768 39432 1820 39438
rect 1768 39374 1820 39380
rect 1676 38480 1728 38486
rect 1676 38422 1728 38428
rect 1584 37800 1636 37806
rect 1780 37777 1808 39374
rect 1872 38865 1900 39442
rect 1964 39409 1992 39986
rect 2044 39908 2096 39914
rect 2044 39850 2096 39856
rect 2056 39681 2084 39850
rect 2042 39672 2098 39681
rect 2042 39607 2098 39616
rect 1950 39400 2006 39409
rect 1950 39335 2006 39344
rect 1952 39296 2004 39302
rect 1952 39238 2004 39244
rect 1858 38856 1914 38865
rect 1964 38826 1992 39238
rect 1858 38791 1914 38800
rect 1952 38820 2004 38826
rect 1952 38762 2004 38768
rect 1952 38412 2004 38418
rect 1952 38354 2004 38360
rect 1584 37742 1636 37748
rect 1766 37768 1822 37777
rect 1490 37496 1546 37505
rect 1490 37431 1546 37440
rect 1492 37392 1544 37398
rect 1492 37334 1544 37340
rect 1400 37324 1452 37330
rect 1400 37266 1452 37272
rect 1504 37097 1532 37334
rect 1596 37330 1624 37742
rect 1676 37732 1728 37738
rect 1766 37703 1822 37712
rect 1676 37674 1728 37680
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1490 37088 1546 37097
rect 1490 37023 1546 37032
rect 1400 36916 1452 36922
rect 1400 36858 1452 36864
rect 1412 34746 1440 36858
rect 1596 36786 1624 37266
rect 1688 37194 1716 37674
rect 1780 37330 1808 37703
rect 1860 37664 1912 37670
rect 1860 37606 1912 37612
rect 1768 37324 1820 37330
rect 1768 37266 1820 37272
rect 1676 37188 1728 37194
rect 1676 37130 1728 37136
rect 1766 37088 1822 37097
rect 1766 37023 1822 37032
rect 1584 36780 1636 36786
rect 1584 36722 1636 36728
rect 1596 36242 1624 36722
rect 1780 36718 1808 37023
rect 1768 36712 1820 36718
rect 1768 36654 1820 36660
rect 1492 36236 1544 36242
rect 1492 36178 1544 36184
rect 1584 36236 1636 36242
rect 1584 36178 1636 36184
rect 1504 35290 1532 36178
rect 1596 35834 1624 36178
rect 1674 35864 1730 35873
rect 1584 35828 1636 35834
rect 1674 35799 1730 35808
rect 1584 35770 1636 35776
rect 1492 35284 1544 35290
rect 1492 35226 1544 35232
rect 1492 35148 1544 35154
rect 1492 35090 1544 35096
rect 1400 34740 1452 34746
rect 1400 34682 1452 34688
rect 1504 34066 1532 35090
rect 1596 34542 1624 35770
rect 1584 34536 1636 34542
rect 1584 34478 1636 34484
rect 1492 34060 1544 34066
rect 1412 34020 1492 34048
rect 1412 32348 1440 34020
rect 1492 34002 1544 34008
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1504 32910 1532 33254
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1492 32768 1544 32774
rect 1492 32710 1544 32716
rect 1504 32502 1532 32710
rect 1492 32496 1544 32502
rect 1492 32438 1544 32444
rect 1412 32320 1624 32348
rect 1400 32224 1452 32230
rect 1400 32166 1452 32172
rect 1412 30977 1440 32166
rect 1492 31816 1544 31822
rect 1492 31758 1544 31764
rect 1504 31482 1532 31758
rect 1492 31476 1544 31482
rect 1492 31418 1544 31424
rect 1492 31136 1544 31142
rect 1492 31078 1544 31084
rect 1398 30968 1454 30977
rect 1398 30903 1454 30912
rect 1400 30796 1452 30802
rect 1400 30738 1452 30744
rect 1412 30190 1440 30738
rect 1400 30184 1452 30190
rect 1400 30126 1452 30132
rect 1400 30048 1452 30054
rect 1400 29990 1452 29996
rect 1412 29714 1440 29990
rect 1504 29850 1532 31078
rect 1492 29844 1544 29850
rect 1492 29786 1544 29792
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1596 29238 1624 32320
rect 1688 32026 1716 35799
rect 1780 35630 1808 36654
rect 1768 35624 1820 35630
rect 1768 35566 1820 35572
rect 1768 35148 1820 35154
rect 1768 35090 1820 35096
rect 1780 35057 1808 35090
rect 1766 35048 1822 35057
rect 1766 34983 1822 34992
rect 1780 34474 1808 34983
rect 1768 34468 1820 34474
rect 1768 34410 1820 34416
rect 1872 34406 1900 37606
rect 1964 37233 1992 38354
rect 2056 38185 2084 39607
rect 2136 38820 2188 38826
rect 2136 38762 2188 38768
rect 2148 38418 2176 38762
rect 2240 38554 2268 40326
rect 2332 39506 2360 40530
rect 2424 40186 2452 40530
rect 2516 40186 2544 40559
rect 2412 40180 2464 40186
rect 2412 40122 2464 40128
rect 2504 40180 2556 40186
rect 2504 40122 2556 40128
rect 2502 40080 2558 40089
rect 2412 40044 2464 40050
rect 2502 40015 2558 40024
rect 2412 39986 2464 39992
rect 2424 39574 2452 39986
rect 2412 39568 2464 39574
rect 2412 39510 2464 39516
rect 2320 39500 2372 39506
rect 2320 39442 2372 39448
rect 2332 39273 2360 39442
rect 2318 39264 2374 39273
rect 2318 39199 2374 39208
rect 2332 38554 2360 39199
rect 2516 38654 2544 40015
rect 2424 38626 2544 38654
rect 2228 38548 2280 38554
rect 2228 38490 2280 38496
rect 2320 38548 2372 38554
rect 2320 38490 2372 38496
rect 2136 38412 2188 38418
rect 2136 38354 2188 38360
rect 2042 38176 2098 38185
rect 2042 38111 2098 38120
rect 2044 38004 2096 38010
rect 2044 37946 2096 37952
rect 1950 37224 2006 37233
rect 1950 37159 2006 37168
rect 1952 36100 2004 36106
rect 1952 36042 2004 36048
rect 1964 35698 1992 36042
rect 2056 35737 2084 37946
rect 2424 37754 2452 38626
rect 2608 38026 2636 40870
rect 2700 39982 2728 41210
rect 2688 39976 2740 39982
rect 2792 39953 2820 43500
rect 4448 43194 4476 43500
rect 2964 43172 3016 43178
rect 2964 43114 3016 43120
rect 4264 43166 4476 43194
rect 2872 42560 2924 42566
rect 2872 42502 2924 42508
rect 2884 42106 2912 42502
rect 2976 42362 3004 43114
rect 4264 42770 4292 43166
rect 4322 43004 4630 43013
rect 4322 43002 4328 43004
rect 4384 43002 4408 43004
rect 4464 43002 4488 43004
rect 4544 43002 4568 43004
rect 4624 43002 4630 43004
rect 4384 42950 4386 43002
rect 4566 42950 4568 43002
rect 4322 42948 4328 42950
rect 4384 42948 4408 42950
rect 4464 42948 4488 42950
rect 4544 42948 4568 42950
rect 4624 42948 4630 42950
rect 4322 42939 4630 42948
rect 4252 42764 4304 42770
rect 4252 42706 4304 42712
rect 5356 42764 5408 42770
rect 5356 42706 5408 42712
rect 4896 42696 4948 42702
rect 4250 42664 4306 42673
rect 3148 42628 3200 42634
rect 4896 42638 4948 42644
rect 5264 42696 5316 42702
rect 5264 42638 5316 42644
rect 4250 42599 4306 42608
rect 3148 42570 3200 42576
rect 2964 42356 3016 42362
rect 2964 42298 3016 42304
rect 2884 42078 3004 42106
rect 3160 42090 3188 42570
rect 4068 42560 4120 42566
rect 4068 42502 4120 42508
rect 4158 42528 4214 42537
rect 3662 42460 3970 42469
rect 3662 42458 3668 42460
rect 3724 42458 3748 42460
rect 3804 42458 3828 42460
rect 3884 42458 3908 42460
rect 3964 42458 3970 42460
rect 3724 42406 3726 42458
rect 3906 42406 3908 42458
rect 3662 42404 3668 42406
rect 3724 42404 3748 42406
rect 3804 42404 3828 42406
rect 3884 42404 3908 42406
rect 3964 42404 3970 42406
rect 3662 42395 3970 42404
rect 3792 42288 3844 42294
rect 3792 42230 3844 42236
rect 2872 42016 2924 42022
rect 2872 41958 2924 41964
rect 2884 41682 2912 41958
rect 2872 41676 2924 41682
rect 2872 41618 2924 41624
rect 2976 40633 3004 42078
rect 3148 42084 3200 42090
rect 3148 42026 3200 42032
rect 3056 40996 3108 41002
rect 3056 40938 3108 40944
rect 2962 40624 3018 40633
rect 2962 40559 3018 40568
rect 2976 40202 3004 40559
rect 3068 40225 3096 40938
rect 2884 40174 3004 40202
rect 3054 40216 3110 40225
rect 2884 40089 2912 40174
rect 3054 40151 3056 40160
rect 3108 40151 3110 40160
rect 3056 40122 3108 40128
rect 2870 40080 2926 40089
rect 2870 40015 2926 40024
rect 2964 39976 3016 39982
rect 2688 39918 2740 39924
rect 2778 39944 2834 39953
rect 2700 38962 2728 39918
rect 2778 39879 2834 39888
rect 2884 39924 2964 39930
rect 2884 39918 3016 39924
rect 2884 39902 3004 39918
rect 3160 39914 3188 42026
rect 3804 41614 3832 42230
rect 3976 42152 4028 42158
rect 3976 42094 4028 42100
rect 3332 41608 3384 41614
rect 3332 41550 3384 41556
rect 3792 41608 3844 41614
rect 3792 41550 3844 41556
rect 3344 40769 3372 41550
rect 3988 41546 4016 42094
rect 3976 41540 4028 41546
rect 3976 41482 4028 41488
rect 3516 41472 3568 41478
rect 3516 41414 3568 41420
rect 3424 40928 3476 40934
rect 3424 40870 3476 40876
rect 3330 40760 3386 40769
rect 3330 40695 3386 40704
rect 3240 40656 3292 40662
rect 3240 40598 3292 40604
rect 3148 39908 3200 39914
rect 2884 39794 2912 39902
rect 3148 39850 3200 39856
rect 2792 39766 2912 39794
rect 2964 39840 3016 39846
rect 2964 39782 3016 39788
rect 2792 39642 2820 39766
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 2688 38956 2740 38962
rect 2688 38898 2740 38904
rect 2792 38894 2820 39578
rect 2976 39420 3004 39782
rect 3054 39536 3110 39545
rect 3054 39471 3056 39480
rect 3108 39471 3110 39480
rect 3056 39442 3108 39448
rect 2884 39392 3004 39420
rect 2884 39284 2912 39392
rect 3056 39296 3108 39302
rect 2884 39256 3004 39284
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2608 37998 2728 38026
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2332 37726 2452 37754
rect 2504 37800 2556 37806
rect 2504 37742 2556 37748
rect 2228 37664 2280 37670
rect 2228 37606 2280 37612
rect 2134 37496 2190 37505
rect 2134 37431 2190 37440
rect 2042 35728 2098 35737
rect 1952 35692 2004 35698
rect 2042 35663 2098 35672
rect 1952 35634 2004 35640
rect 1952 35148 2004 35154
rect 1952 35090 2004 35096
rect 1860 34400 1912 34406
rect 1860 34342 1912 34348
rect 1964 34184 1992 35090
rect 2056 34746 2084 35663
rect 2148 35222 2176 37431
rect 2240 37330 2268 37606
rect 2228 37324 2280 37330
rect 2228 37266 2280 37272
rect 2332 36666 2360 37726
rect 2516 36689 2544 37742
rect 2240 36638 2360 36666
rect 2502 36680 2558 36689
rect 2136 35216 2188 35222
rect 2136 35158 2188 35164
rect 2044 34740 2096 34746
rect 2044 34682 2096 34688
rect 2240 34626 2268 36638
rect 2502 36615 2558 36624
rect 2412 35828 2464 35834
rect 2412 35770 2464 35776
rect 2424 34678 2452 35770
rect 2516 35698 2544 36615
rect 2504 35692 2556 35698
rect 2504 35634 2556 35640
rect 2608 35329 2636 37810
rect 2700 37194 2728 37998
rect 2688 37188 2740 37194
rect 2688 37130 2740 37136
rect 2700 35834 2728 37130
rect 2792 36786 2820 38830
rect 2872 37936 2924 37942
rect 2872 37878 2924 37884
rect 2884 37777 2912 37878
rect 2870 37768 2926 37777
rect 2870 37703 2926 37712
rect 2872 37664 2924 37670
rect 2872 37606 2924 37612
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2688 35828 2740 35834
rect 2688 35770 2740 35776
rect 2688 35692 2740 35698
rect 2688 35634 2740 35640
rect 2594 35320 2650 35329
rect 2594 35255 2650 35264
rect 2596 34740 2648 34746
rect 2596 34682 2648 34688
rect 1780 34156 1992 34184
rect 2148 34598 2268 34626
rect 2412 34672 2464 34678
rect 2412 34614 2464 34620
rect 1676 32020 1728 32026
rect 1676 31962 1728 31968
rect 1780 31872 1808 34156
rect 1952 34060 2004 34066
rect 1952 34002 2004 34008
rect 1858 33688 1914 33697
rect 1858 33623 1914 33632
rect 1872 32201 1900 33623
rect 1964 33386 1992 34002
rect 2044 33652 2096 33658
rect 2044 33594 2096 33600
rect 1952 33380 2004 33386
rect 1952 33322 2004 33328
rect 1964 33289 1992 33322
rect 1950 33280 2006 33289
rect 1950 33215 2006 33224
rect 1858 32192 1914 32201
rect 1858 32127 1914 32136
rect 2056 32026 2084 33594
rect 2148 32570 2176 34598
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2240 34066 2268 34478
rect 2502 34232 2558 34241
rect 2502 34167 2558 34176
rect 2228 34060 2280 34066
rect 2228 34002 2280 34008
rect 2240 33522 2268 34002
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2240 33046 2268 33458
rect 2320 33448 2372 33454
rect 2318 33416 2320 33425
rect 2372 33416 2374 33425
rect 2318 33351 2374 33360
rect 2228 33040 2280 33046
rect 2228 32982 2280 32988
rect 2136 32564 2188 32570
rect 2136 32506 2188 32512
rect 2424 32450 2452 33798
rect 2516 33522 2544 34167
rect 2504 33516 2556 33522
rect 2504 33458 2556 33464
rect 2608 33402 2636 34682
rect 2700 33504 2728 35634
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2792 35290 2820 35566
rect 2780 35284 2832 35290
rect 2780 35226 2832 35232
rect 2884 33658 2912 37606
rect 2872 33652 2924 33658
rect 2872 33594 2924 33600
rect 2700 33476 2820 33504
rect 2608 33374 2728 33402
rect 2596 33312 2648 33318
rect 2596 33254 2648 33260
rect 2608 33153 2636 33254
rect 2594 33144 2650 33153
rect 2594 33079 2650 33088
rect 2700 33017 2728 33374
rect 2686 33008 2742 33017
rect 2504 32972 2556 32978
rect 2686 32943 2742 32952
rect 2504 32914 2556 32920
rect 2516 32570 2544 32914
rect 2688 32904 2740 32910
rect 2688 32846 2740 32852
rect 2504 32564 2556 32570
rect 2504 32506 2556 32512
rect 2148 32422 2544 32450
rect 2044 32020 2096 32026
rect 2044 31962 2096 31968
rect 2148 31890 2176 32422
rect 2412 32292 2464 32298
rect 2412 32234 2464 32240
rect 2424 31958 2452 32234
rect 2320 31952 2372 31958
rect 2320 31894 2372 31900
rect 2412 31952 2464 31958
rect 2412 31894 2464 31900
rect 1688 31844 1808 31872
rect 1952 31884 2004 31890
rect 1688 31521 1716 31844
rect 1952 31826 2004 31832
rect 2136 31884 2188 31890
rect 2136 31826 2188 31832
rect 2228 31884 2280 31890
rect 2228 31826 2280 31832
rect 1674 31512 1730 31521
rect 1674 31447 1730 31456
rect 1964 31278 1992 31826
rect 2042 31784 2098 31793
rect 2042 31719 2098 31728
rect 1952 31272 2004 31278
rect 1952 31214 2004 31220
rect 1676 31204 1728 31210
rect 1676 31146 1728 31152
rect 1688 29782 1716 31146
rect 1860 30592 1912 30598
rect 1860 30534 1912 30540
rect 1766 29880 1822 29889
rect 1766 29815 1768 29824
rect 1820 29815 1822 29824
rect 1768 29786 1820 29792
rect 1676 29776 1728 29782
rect 1676 29718 1728 29724
rect 1584 29232 1636 29238
rect 1584 29174 1636 29180
rect 1596 29102 1624 29174
rect 1584 29096 1636 29102
rect 1688 29073 1716 29718
rect 1768 29640 1820 29646
rect 1768 29582 1820 29588
rect 1584 29038 1636 29044
rect 1674 29064 1730 29073
rect 1674 28999 1730 29008
rect 1320 28886 1624 28914
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1308 26784 1360 26790
rect 1308 26726 1360 26732
rect 1320 26586 1348 26726
rect 1308 26580 1360 26586
rect 1308 26522 1360 26528
rect 1412 26518 1440 27950
rect 1492 27328 1544 27334
rect 1492 27270 1544 27276
rect 1504 26926 1532 27270
rect 1492 26920 1544 26926
rect 1492 26862 1544 26868
rect 1400 26512 1452 26518
rect 1400 26454 1452 26460
rect 1412 25430 1440 26454
rect 1504 26450 1532 26862
rect 1492 26444 1544 26450
rect 1492 26386 1544 26392
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 25838 1532 26182
rect 1492 25832 1544 25838
rect 1492 25774 1544 25780
rect 1400 25424 1452 25430
rect 1400 25366 1452 25372
rect 1308 24744 1360 24750
rect 1308 24686 1360 24692
rect 1216 23792 1268 23798
rect 1216 23734 1268 23740
rect 1320 23662 1348 24686
rect 1412 24342 1440 25366
rect 1504 24750 1532 25774
rect 1492 24744 1544 24750
rect 1492 24686 1544 24692
rect 1492 24608 1544 24614
rect 1492 24550 1544 24556
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1504 24274 1532 24550
rect 1492 24268 1544 24274
rect 1492 24210 1544 24216
rect 1596 24154 1624 28886
rect 1780 27538 1808 29582
rect 1872 29578 1900 30534
rect 1964 30394 1992 31214
rect 1952 30388 2004 30394
rect 1952 30330 2004 30336
rect 2056 30274 2084 31719
rect 2240 31482 2268 31826
rect 2228 31476 2280 31482
rect 2228 31418 2280 31424
rect 2332 31362 2360 31894
rect 1964 30246 2084 30274
rect 2148 31334 2360 31362
rect 1860 29572 1912 29578
rect 1860 29514 1912 29520
rect 1964 29238 1992 30246
rect 2148 29850 2176 31334
rect 2228 31272 2280 31278
rect 2228 31214 2280 31220
rect 2240 30734 2268 31214
rect 2424 30802 2452 31894
rect 2516 31822 2544 32422
rect 2596 31884 2648 31890
rect 2596 31826 2648 31832
rect 2504 31816 2556 31822
rect 2504 31758 2556 31764
rect 2502 31240 2558 31249
rect 2502 31175 2504 31184
rect 2556 31175 2558 31184
rect 2504 31146 2556 31152
rect 2608 30954 2636 31826
rect 2700 31414 2728 32846
rect 2792 31770 2820 33476
rect 2870 33144 2926 33153
rect 2870 33079 2872 33088
rect 2924 33079 2926 33088
rect 2872 33050 2924 33056
rect 2870 33008 2926 33017
rect 2870 32943 2926 32952
rect 2884 31890 2912 32943
rect 2872 31884 2924 31890
rect 2872 31826 2924 31832
rect 2792 31742 2912 31770
rect 2780 31680 2832 31686
rect 2780 31622 2832 31628
rect 2688 31408 2740 31414
rect 2688 31350 2740 31356
rect 2688 31272 2740 31278
rect 2688 31214 2740 31220
rect 2516 30926 2636 30954
rect 2412 30796 2464 30802
rect 2332 30756 2412 30784
rect 2228 30728 2280 30734
rect 2228 30670 2280 30676
rect 2136 29844 2188 29850
rect 2136 29786 2188 29792
rect 2134 29608 2190 29617
rect 2134 29543 2190 29552
rect 1860 29232 1912 29238
rect 1860 29174 1912 29180
rect 1952 29232 2004 29238
rect 1952 29174 2004 29180
rect 2042 29200 2098 29209
rect 1872 28558 1900 29174
rect 2042 29135 2098 29144
rect 1952 29096 2004 29102
rect 1952 29038 2004 29044
rect 1860 28552 1912 28558
rect 1860 28494 1912 28500
rect 1768 27532 1820 27538
rect 1768 27474 1820 27480
rect 1768 27124 1820 27130
rect 1768 27066 1820 27072
rect 1676 27056 1728 27062
rect 1676 26998 1728 27004
rect 1688 25498 1716 26998
rect 1676 25492 1728 25498
rect 1676 25434 1728 25440
rect 1780 24857 1808 27066
rect 1872 26994 1900 28494
rect 1964 27946 1992 29038
rect 1952 27940 2004 27946
rect 1952 27882 2004 27888
rect 1964 27849 1992 27882
rect 1950 27840 2006 27849
rect 1950 27775 2006 27784
rect 2056 27690 2084 29135
rect 1964 27662 2084 27690
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 1872 26246 1900 26930
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1964 26194 1992 27662
rect 2044 27328 2096 27334
rect 2044 27270 2096 27276
rect 2056 26353 2084 27270
rect 2148 27130 2176 29543
rect 2240 28082 2268 30670
rect 2332 30190 2360 30756
rect 2412 30738 2464 30744
rect 2412 30320 2464 30326
rect 2410 30288 2412 30297
rect 2464 30288 2466 30297
rect 2410 30223 2466 30232
rect 2320 30184 2372 30190
rect 2320 30126 2372 30132
rect 2412 30184 2464 30190
rect 2412 30126 2464 30132
rect 2424 29850 2452 30126
rect 2320 29844 2372 29850
rect 2320 29786 2372 29792
rect 2412 29844 2464 29850
rect 2412 29786 2464 29792
rect 2332 29696 2360 29786
rect 2516 29714 2544 30926
rect 2596 30864 2648 30870
rect 2596 30806 2648 30812
rect 2608 30190 2636 30806
rect 2700 30258 2728 31214
rect 2792 30938 2820 31622
rect 2884 30977 2912 31742
rect 2870 30968 2926 30977
rect 2780 30932 2832 30938
rect 2870 30903 2926 30912
rect 2780 30874 2832 30880
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2596 30184 2648 30190
rect 2596 30126 2648 30132
rect 2778 30152 2834 30161
rect 2412 29708 2464 29714
rect 2332 29668 2412 29696
rect 2412 29650 2464 29656
rect 2504 29708 2556 29714
rect 2504 29650 2556 29656
rect 2320 29572 2372 29578
rect 2320 29514 2372 29520
rect 2332 29306 2360 29514
rect 2320 29300 2372 29306
rect 2320 29242 2372 29248
rect 2318 28928 2374 28937
rect 2318 28863 2374 28872
rect 2332 28694 2360 28863
rect 2320 28688 2372 28694
rect 2320 28630 2372 28636
rect 2228 28076 2280 28082
rect 2228 28018 2280 28024
rect 2136 27124 2188 27130
rect 2136 27066 2188 27072
rect 2134 26616 2190 26625
rect 2134 26551 2190 26560
rect 2148 26466 2176 26551
rect 2320 26512 2372 26518
rect 2148 26438 2268 26466
rect 2320 26454 2372 26460
rect 2136 26376 2188 26382
rect 2042 26344 2098 26353
rect 2136 26318 2188 26324
rect 2042 26279 2098 26288
rect 1964 26166 2084 26194
rect 1952 25900 2004 25906
rect 1952 25842 2004 25848
rect 1964 25362 1992 25842
rect 1952 25356 2004 25362
rect 1952 25298 2004 25304
rect 1766 24848 1822 24857
rect 1766 24783 1822 24792
rect 1768 24744 1820 24750
rect 1768 24686 1820 24692
rect 1412 24126 1624 24154
rect 1216 23656 1268 23662
rect 1216 23598 1268 23604
rect 1308 23656 1360 23662
rect 1308 23598 1360 23604
rect 1124 23180 1176 23186
rect 1124 23122 1176 23128
rect 1044 22766 1164 22794
rect 1032 22704 1084 22710
rect 1030 22672 1032 22681
rect 1084 22672 1086 22681
rect 1030 22607 1086 22616
rect 1032 22432 1084 22438
rect 1032 22374 1084 22380
rect 940 20052 992 20058
rect 940 19994 992 20000
rect 754 19272 810 19281
rect 860 19264 980 19292
rect 754 19207 810 19216
rect 662 17640 718 17649
rect 662 17575 718 17584
rect 676 12322 704 17575
rect 768 12442 796 19207
rect 952 18766 980 19264
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 952 17785 980 18702
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 846 17232 902 17241
rect 846 17167 902 17176
rect 860 14482 888 17167
rect 938 16960 994 16969
rect 938 16895 994 16904
rect 952 16726 980 16895
rect 940 16720 992 16726
rect 940 16662 992 16668
rect 938 16552 994 16561
rect 938 16487 994 16496
rect 848 14476 900 14482
rect 848 14418 900 14424
rect 848 12708 900 12714
rect 848 12650 900 12656
rect 860 12617 888 12650
rect 846 12608 902 12617
rect 846 12543 902 12552
rect 756 12436 808 12442
rect 952 12434 980 16487
rect 756 12378 808 12384
rect 860 12406 980 12434
rect 676 12294 796 12322
rect 584 12158 704 12186
rect 572 12096 624 12102
rect 572 12038 624 12044
rect 584 11257 612 12038
rect 570 11248 626 11257
rect 570 11183 626 11192
rect 676 10538 704 12158
rect 664 10532 716 10538
rect 664 10474 716 10480
rect 768 9654 796 12294
rect 756 9648 808 9654
rect 756 9590 808 9596
rect 860 9450 888 12406
rect 938 12064 994 12073
rect 938 11999 994 12008
rect 952 10674 980 11999
rect 1044 11898 1072 22374
rect 1136 21978 1164 22766
rect 1228 22094 1256 23598
rect 1306 23488 1362 23497
rect 1306 23423 1362 23432
rect 1320 22642 1348 23423
rect 1308 22636 1360 22642
rect 1308 22578 1360 22584
rect 1228 22066 1348 22094
rect 1136 21950 1256 21978
rect 1124 21888 1176 21894
rect 1124 21830 1176 21836
rect 1136 20913 1164 21830
rect 1228 21554 1256 21950
rect 1216 21548 1268 21554
rect 1216 21490 1268 21496
rect 1320 21486 1348 22066
rect 1412 21962 1440 24126
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1492 23656 1544 23662
rect 1492 23598 1544 23604
rect 1504 23474 1532 23598
rect 1504 23446 1624 23474
rect 1492 23316 1544 23322
rect 1492 23258 1544 23264
rect 1400 21956 1452 21962
rect 1400 21898 1452 21904
rect 1504 21690 1532 23258
rect 1596 22574 1624 23446
rect 1584 22568 1636 22574
rect 1584 22510 1636 22516
rect 1688 21894 1716 23666
rect 1780 23322 1808 24686
rect 1860 24676 1912 24682
rect 1860 24618 1912 24624
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1676 21888 1728 21894
rect 1676 21830 1728 21836
rect 1766 21856 1822 21865
rect 1766 21791 1822 21800
rect 1492 21684 1544 21690
rect 1492 21626 1544 21632
rect 1308 21480 1360 21486
rect 1308 21422 1360 21428
rect 1122 20904 1178 20913
rect 1122 20839 1178 20848
rect 1216 20800 1268 20806
rect 1216 20742 1268 20748
rect 1122 20632 1178 20641
rect 1122 20567 1178 20576
rect 1032 11892 1084 11898
rect 1032 11834 1084 11840
rect 1136 11694 1164 20567
rect 1228 20466 1256 20742
rect 1216 20460 1268 20466
rect 1216 20402 1268 20408
rect 1320 20346 1348 21422
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1674 21312 1730 21321
rect 1412 20398 1440 21286
rect 1674 21247 1730 21256
rect 1492 21004 1544 21010
rect 1492 20946 1544 20952
rect 1504 20398 1532 20946
rect 1688 20641 1716 21247
rect 1674 20632 1730 20641
rect 1674 20567 1730 20576
rect 1780 20482 1808 21791
rect 1688 20454 1808 20482
rect 1228 20318 1348 20346
rect 1400 20392 1452 20398
rect 1400 20334 1452 20340
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1228 16658 1256 20318
rect 1308 19712 1360 19718
rect 1308 19654 1360 19660
rect 1320 18154 1348 19654
rect 1412 18834 1440 20334
rect 1504 19514 1532 20334
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1492 19372 1544 19378
rect 1492 19314 1544 19320
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1308 18148 1360 18154
rect 1308 18090 1360 18096
rect 1308 17536 1360 17542
rect 1308 17478 1360 17484
rect 1320 17134 1348 17478
rect 1412 17134 1440 18770
rect 1308 17128 1360 17134
rect 1308 17070 1360 17076
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1306 16824 1362 16833
rect 1306 16759 1362 16768
rect 1216 16652 1268 16658
rect 1216 16594 1268 16600
rect 1214 11792 1270 11801
rect 1214 11727 1270 11736
rect 1124 11688 1176 11694
rect 1124 11630 1176 11636
rect 1032 11552 1084 11558
rect 1030 11520 1032 11529
rect 1084 11520 1086 11529
rect 1030 11455 1086 11464
rect 940 10668 992 10674
rect 940 10610 992 10616
rect 1228 9586 1256 11727
rect 1216 9580 1268 9586
rect 1216 9522 1268 9528
rect 848 9444 900 9450
rect 848 9386 900 9392
rect 1320 9178 1348 16759
rect 1412 14482 1440 17070
rect 1504 16674 1532 19314
rect 1596 19310 1624 20198
rect 1688 20058 1716 20454
rect 1768 20392 1820 20398
rect 1768 20334 1820 20340
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1688 19825 1716 19858
rect 1674 19816 1730 19825
rect 1674 19751 1730 19760
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1584 19304 1636 19310
rect 1584 19246 1636 19252
rect 1584 18828 1636 18834
rect 1584 18770 1636 18776
rect 1596 18426 1624 18770
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1596 17270 1624 18090
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1504 16646 1624 16674
rect 1490 16552 1546 16561
rect 1490 16487 1546 16496
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1412 12782 1440 14418
rect 1504 13938 1532 16487
rect 1596 16250 1624 16646
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1688 16130 1716 19654
rect 1780 18902 1808 20334
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1780 16794 1808 18838
rect 1768 16788 1820 16794
rect 1768 16730 1820 16736
rect 1768 16652 1820 16658
rect 1768 16594 1820 16600
rect 1596 16102 1716 16130
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12434 1440 12718
rect 1412 12406 1532 12434
rect 1400 12368 1452 12374
rect 1398 12336 1400 12345
rect 1452 12336 1454 12345
rect 1398 12271 1454 12280
rect 1400 12232 1452 12238
rect 1504 12220 1532 12406
rect 1596 12374 1624 16102
rect 1780 15978 1808 16594
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 1674 15736 1730 15745
rect 1780 15706 1808 15914
rect 1674 15671 1676 15680
rect 1728 15671 1730 15680
rect 1768 15700 1820 15706
rect 1676 15642 1728 15648
rect 1768 15642 1820 15648
rect 1674 15192 1730 15201
rect 1674 15127 1730 15136
rect 1688 14074 1716 15127
rect 1768 14272 1820 14278
rect 1768 14214 1820 14220
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1584 12368 1636 12374
rect 1584 12310 1636 12316
rect 1452 12192 1532 12220
rect 1400 12174 1452 12180
rect 1412 10606 1440 12174
rect 1596 11626 1624 12310
rect 1584 11620 1636 11626
rect 1584 11562 1636 11568
rect 1688 11286 1716 13874
rect 1676 11280 1728 11286
rect 1676 11222 1728 11228
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10674 1624 10950
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1400 10600 1452 10606
rect 1400 10542 1452 10548
rect 1412 9518 1440 10542
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1412 8430 1440 9454
rect 1780 8430 1808 14214
rect 1872 10198 1900 24618
rect 1964 24426 1992 25298
rect 2056 24596 2084 26166
rect 2148 24750 2176 26318
rect 2136 24744 2188 24750
rect 2240 24721 2268 26438
rect 2332 25158 2360 26454
rect 2424 26353 2452 29650
rect 2516 29617 2544 29650
rect 2502 29608 2558 29617
rect 2502 29543 2558 29552
rect 2608 29492 2636 30126
rect 2688 30116 2740 30122
rect 2778 30087 2780 30096
rect 2688 30058 2740 30064
rect 2832 30087 2834 30096
rect 2780 30058 2832 30064
rect 2700 29782 2728 30058
rect 2688 29776 2740 29782
rect 2688 29718 2740 29724
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2778 29608 2834 29617
rect 2516 29464 2636 29492
rect 2516 29102 2544 29464
rect 2700 29209 2728 29582
rect 2778 29543 2834 29552
rect 2686 29200 2742 29209
rect 2686 29135 2742 29144
rect 2504 29096 2556 29102
rect 2504 29038 2556 29044
rect 2596 29096 2648 29102
rect 2596 29038 2648 29044
rect 2516 27674 2544 29038
rect 2608 28218 2636 29038
rect 2688 29028 2740 29034
rect 2688 28970 2740 28976
rect 2700 28762 2728 28970
rect 2688 28756 2740 28762
rect 2688 28698 2740 28704
rect 2596 28212 2648 28218
rect 2596 28154 2648 28160
rect 2594 27704 2650 27713
rect 2504 27668 2556 27674
rect 2594 27639 2650 27648
rect 2504 27610 2556 27616
rect 2516 26450 2544 27610
rect 2608 27418 2636 27639
rect 2700 27538 2728 28698
rect 2792 28257 2820 29543
rect 2884 29510 2912 30534
rect 2976 30036 3004 39256
rect 3056 39238 3108 39244
rect 3068 37738 3096 39238
rect 3056 37732 3108 37738
rect 3056 37674 3108 37680
rect 3056 37120 3108 37126
rect 3056 37062 3108 37068
rect 3068 36854 3096 37062
rect 3160 36922 3188 39850
rect 3252 38978 3280 40598
rect 3332 40520 3384 40526
rect 3332 40462 3384 40468
rect 3344 39098 3372 40462
rect 3436 40089 3464 40870
rect 3528 40662 3556 41414
rect 3662 41372 3970 41381
rect 3662 41370 3668 41372
rect 3724 41370 3748 41372
rect 3804 41370 3828 41372
rect 3884 41370 3908 41372
rect 3964 41370 3970 41372
rect 3724 41318 3726 41370
rect 3906 41318 3908 41370
rect 3662 41316 3668 41318
rect 3724 41316 3748 41318
rect 3804 41316 3828 41318
rect 3884 41316 3908 41318
rect 3964 41316 3970 41318
rect 3662 41307 3970 41316
rect 4080 41002 4108 42502
rect 4158 42463 4214 42472
rect 4172 42362 4200 42463
rect 4160 42356 4212 42362
rect 4160 42298 4212 42304
rect 4172 42158 4200 42298
rect 4264 42226 4292 42599
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4160 42152 4212 42158
rect 4160 42094 4212 42100
rect 4160 42016 4212 42022
rect 4160 41958 4212 41964
rect 4172 41682 4200 41958
rect 4264 41698 4292 42162
rect 4344 42152 4396 42158
rect 4804 42152 4856 42158
rect 4396 42100 4752 42106
rect 4344 42094 4752 42100
rect 4804 42094 4856 42100
rect 4356 42078 4752 42094
rect 4322 41916 4630 41925
rect 4322 41914 4328 41916
rect 4384 41914 4408 41916
rect 4464 41914 4488 41916
rect 4544 41914 4568 41916
rect 4624 41914 4630 41916
rect 4384 41862 4386 41914
rect 4566 41862 4568 41914
rect 4322 41860 4328 41862
rect 4384 41860 4408 41862
rect 4464 41860 4488 41862
rect 4544 41860 4568 41862
rect 4624 41860 4630 41862
rect 4322 41851 4630 41860
rect 4160 41676 4212 41682
rect 4264 41670 4384 41698
rect 4160 41618 4212 41624
rect 4252 41608 4304 41614
rect 4252 41550 4304 41556
rect 4264 41070 4292 41550
rect 4252 41064 4304 41070
rect 4252 41006 4304 41012
rect 4068 40996 4120 41002
rect 4068 40938 4120 40944
rect 4356 40916 4384 41670
rect 4264 40888 4384 40916
rect 4160 40724 4212 40730
rect 4264 40712 4292 40888
rect 4322 40828 4630 40837
rect 4322 40826 4328 40828
rect 4384 40826 4408 40828
rect 4464 40826 4488 40828
rect 4544 40826 4568 40828
rect 4624 40826 4630 40828
rect 4384 40774 4386 40826
rect 4566 40774 4568 40826
rect 4322 40772 4328 40774
rect 4384 40772 4408 40774
rect 4464 40772 4488 40774
rect 4544 40772 4568 40774
rect 4624 40772 4630 40774
rect 4322 40763 4630 40772
rect 4264 40684 4568 40712
rect 4160 40666 4212 40672
rect 3516 40656 3568 40662
rect 3516 40598 3568 40604
rect 4172 40594 4200 40666
rect 4160 40588 4212 40594
rect 4160 40530 4212 40536
rect 4252 40588 4304 40594
rect 4252 40530 4304 40536
rect 3514 40352 3570 40361
rect 3514 40287 3570 40296
rect 3422 40080 3478 40089
rect 3422 40015 3478 40024
rect 3424 39432 3476 39438
rect 3424 39374 3476 39380
rect 3332 39092 3384 39098
rect 3332 39034 3384 39040
rect 3252 38950 3372 38978
rect 3240 38208 3292 38214
rect 3240 38150 3292 38156
rect 3252 36922 3280 38150
rect 3344 37874 3372 38950
rect 3436 38282 3464 39374
rect 3528 39098 3556 40287
rect 3662 40284 3970 40293
rect 3662 40282 3668 40284
rect 3724 40282 3748 40284
rect 3804 40282 3828 40284
rect 3884 40282 3908 40284
rect 3964 40282 3970 40284
rect 3724 40230 3726 40282
rect 3906 40230 3908 40282
rect 3662 40228 3668 40230
rect 3724 40228 3748 40230
rect 3804 40228 3828 40230
rect 3884 40228 3908 40230
rect 3964 40228 3970 40230
rect 3662 40219 3970 40228
rect 3700 40180 3752 40186
rect 3700 40122 3752 40128
rect 3712 39914 3740 40122
rect 4172 40118 4200 40530
rect 4264 40458 4292 40530
rect 4252 40452 4304 40458
rect 4252 40394 4304 40400
rect 4160 40112 4212 40118
rect 4160 40054 4212 40060
rect 4356 39982 4384 40684
rect 4540 40594 4568 40684
rect 4528 40588 4580 40594
rect 4528 40530 4580 40536
rect 4620 40520 4672 40526
rect 4620 40462 4672 40468
rect 4436 40384 4488 40390
rect 4436 40326 4488 40332
rect 4448 39982 4476 40326
rect 4528 40044 4580 40050
rect 4528 39986 4580 39992
rect 4160 39976 4212 39982
rect 4344 39976 4396 39982
rect 4160 39918 4212 39924
rect 4264 39936 4344 39964
rect 3700 39908 3752 39914
rect 3700 39850 3752 39856
rect 4068 39364 4120 39370
rect 4068 39306 4120 39312
rect 3662 39196 3970 39205
rect 3662 39194 3668 39196
rect 3724 39194 3748 39196
rect 3804 39194 3828 39196
rect 3884 39194 3908 39196
rect 3964 39194 3970 39196
rect 3724 39142 3726 39194
rect 3906 39142 3908 39194
rect 3662 39140 3668 39142
rect 3724 39140 3748 39142
rect 3804 39140 3828 39142
rect 3884 39140 3908 39142
rect 3964 39140 3970 39142
rect 3662 39131 3970 39140
rect 3516 39092 3568 39098
rect 3516 39034 3568 39040
rect 3884 39024 3936 39030
rect 3882 38992 3884 39001
rect 3936 38992 3938 39001
rect 3882 38927 3938 38936
rect 3516 38752 3568 38758
rect 4080 38706 4108 39306
rect 4172 38962 4200 39918
rect 4264 39506 4292 39936
rect 4344 39918 4396 39924
rect 4436 39976 4488 39982
rect 4436 39918 4488 39924
rect 4540 39846 4568 39986
rect 4632 39982 4660 40462
rect 4620 39976 4672 39982
rect 4620 39918 4672 39924
rect 4528 39840 4580 39846
rect 4528 39782 4580 39788
rect 4322 39740 4630 39749
rect 4322 39738 4328 39740
rect 4384 39738 4408 39740
rect 4464 39738 4488 39740
rect 4544 39738 4568 39740
rect 4624 39738 4630 39740
rect 4384 39686 4386 39738
rect 4566 39686 4568 39738
rect 4322 39684 4328 39686
rect 4384 39684 4408 39686
rect 4464 39684 4488 39686
rect 4544 39684 4568 39686
rect 4624 39684 4630 39686
rect 4322 39675 4630 39684
rect 4724 39642 4752 42078
rect 4816 41818 4844 42094
rect 4804 41812 4856 41818
rect 4804 41754 4856 41760
rect 4908 39982 4936 42638
rect 4986 42528 5042 42537
rect 4986 42463 5042 42472
rect 5000 40662 5028 42463
rect 5276 42362 5304 42638
rect 5368 42362 5396 42706
rect 5264 42356 5316 42362
rect 5264 42298 5316 42304
rect 5356 42356 5408 42362
rect 5356 42298 5408 42304
rect 5080 42152 5132 42158
rect 5080 42094 5132 42100
rect 5172 42152 5224 42158
rect 5172 42094 5224 42100
rect 5092 41274 5120 42094
rect 5080 41268 5132 41274
rect 5080 41210 5132 41216
rect 5080 41064 5132 41070
rect 5184 41052 5212 42094
rect 5264 42084 5316 42090
rect 5264 42026 5316 42032
rect 5276 41120 5304 42026
rect 5448 42016 5500 42022
rect 5448 41958 5500 41964
rect 5276 41092 5309 41120
rect 5132 41024 5212 41052
rect 5080 41006 5132 41012
rect 5281 41018 5309 41092
rect 4988 40656 5040 40662
rect 4988 40598 5040 40604
rect 4988 40384 5040 40390
rect 4988 40326 5040 40332
rect 5000 40118 5028 40326
rect 4988 40112 5040 40118
rect 4988 40054 5040 40060
rect 4896 39976 4948 39982
rect 4896 39918 4948 39924
rect 5000 39930 5028 40054
rect 5092 40050 5120 41006
rect 5281 40990 5396 41018
rect 5172 40928 5224 40934
rect 5172 40870 5224 40876
rect 5184 40769 5212 40870
rect 5170 40760 5226 40769
rect 5170 40695 5226 40704
rect 5262 40624 5318 40633
rect 5262 40559 5264 40568
rect 5316 40559 5318 40568
rect 5264 40530 5316 40536
rect 5080 40044 5132 40050
rect 5080 39986 5132 39992
rect 4804 39840 4856 39846
rect 4804 39782 4856 39788
rect 4712 39636 4764 39642
rect 4712 39578 4764 39584
rect 4252 39500 4304 39506
rect 4252 39442 4304 39448
rect 4712 39500 4764 39506
rect 4712 39442 4764 39448
rect 4252 39296 4304 39302
rect 4252 39238 4304 39244
rect 4160 38956 4212 38962
rect 4160 38898 4212 38904
rect 4160 38820 4212 38826
rect 4160 38762 4212 38768
rect 3516 38694 3568 38700
rect 3424 38276 3476 38282
rect 3424 38218 3476 38224
rect 3332 37868 3384 37874
rect 3332 37810 3384 37816
rect 3344 37126 3372 37810
rect 3422 37768 3478 37777
rect 3422 37703 3478 37712
rect 3332 37120 3384 37126
rect 3332 37062 3384 37068
rect 3436 36938 3464 37703
rect 3528 37670 3556 38694
rect 3988 38678 4108 38706
rect 3700 38412 3752 38418
rect 3700 38354 3752 38360
rect 3792 38412 3844 38418
rect 3988 38400 4016 38678
rect 4172 38554 4200 38762
rect 4160 38548 4212 38554
rect 4160 38490 4212 38496
rect 4068 38412 4120 38418
rect 3844 38372 3924 38400
rect 3988 38372 4068 38400
rect 3792 38354 3844 38360
rect 3712 38321 3740 38354
rect 3698 38312 3754 38321
rect 3896 38298 3924 38372
rect 4068 38354 4120 38360
rect 3896 38270 4108 38298
rect 3698 38247 3754 38256
rect 3662 38108 3970 38117
rect 3662 38106 3668 38108
rect 3724 38106 3748 38108
rect 3804 38106 3828 38108
rect 3884 38106 3908 38108
rect 3964 38106 3970 38108
rect 3724 38054 3726 38106
rect 3906 38054 3908 38106
rect 3662 38052 3668 38054
rect 3724 38052 3748 38054
rect 3804 38052 3828 38054
rect 3884 38052 3908 38054
rect 3964 38052 3970 38054
rect 3662 38043 3970 38052
rect 3976 38004 4028 38010
rect 3976 37946 4028 37952
rect 3988 37806 4016 37946
rect 3792 37800 3844 37806
rect 3976 37800 4028 37806
rect 3792 37742 3844 37748
rect 3974 37768 3976 37777
rect 4028 37768 4030 37777
rect 3516 37664 3568 37670
rect 3700 37664 3752 37670
rect 3516 37606 3568 37612
rect 3606 37632 3662 37641
rect 3528 37369 3556 37606
rect 3804 37641 3832 37742
rect 3974 37703 4030 37712
rect 3700 37606 3752 37612
rect 3790 37632 3846 37641
rect 3606 37567 3662 37576
rect 3514 37360 3570 37369
rect 3620 37330 3648 37567
rect 3514 37295 3570 37304
rect 3608 37324 3660 37330
rect 3608 37266 3660 37272
rect 3712 37108 3740 37606
rect 3790 37567 3846 37576
rect 3790 37496 3846 37505
rect 3790 37431 3846 37440
rect 3804 37330 3832 37431
rect 3792 37324 3844 37330
rect 3792 37266 3844 37272
rect 3148 36916 3200 36922
rect 3148 36858 3200 36864
rect 3240 36916 3292 36922
rect 3240 36858 3292 36864
rect 3344 36910 3464 36938
rect 3528 37080 3740 37108
rect 3056 36848 3108 36854
rect 3056 36790 3108 36796
rect 3148 36780 3200 36786
rect 3148 36722 3200 36728
rect 3056 36644 3108 36650
rect 3056 36586 3108 36592
rect 3068 35766 3096 36586
rect 3056 35760 3108 35766
rect 3056 35702 3108 35708
rect 3056 35556 3108 35562
rect 3056 35498 3108 35504
rect 3068 35193 3096 35498
rect 3054 35184 3110 35193
rect 3054 35119 3110 35128
rect 3054 34640 3110 34649
rect 3054 34575 3056 34584
rect 3108 34575 3110 34584
rect 3056 34546 3108 34552
rect 3068 33454 3096 34546
rect 3160 33946 3188 36722
rect 3240 35488 3292 35494
rect 3240 35430 3292 35436
rect 3252 35222 3280 35430
rect 3240 35216 3292 35222
rect 3240 35158 3292 35164
rect 3240 34400 3292 34406
rect 3240 34342 3292 34348
rect 3252 34134 3280 34342
rect 3344 34202 3372 36910
rect 3528 36854 3556 37080
rect 3662 37020 3970 37029
rect 3662 37018 3668 37020
rect 3724 37018 3748 37020
rect 3804 37018 3828 37020
rect 3884 37018 3908 37020
rect 3964 37018 3970 37020
rect 3724 36966 3726 37018
rect 3906 36966 3908 37018
rect 3662 36964 3668 36966
rect 3724 36964 3748 36966
rect 3804 36964 3828 36966
rect 3884 36964 3908 36966
rect 3964 36964 3970 36966
rect 3662 36955 3970 36964
rect 3884 36916 3936 36922
rect 3884 36858 3936 36864
rect 3516 36848 3568 36854
rect 3516 36790 3568 36796
rect 3528 36378 3556 36790
rect 3792 36576 3844 36582
rect 3792 36518 3844 36524
rect 3516 36372 3568 36378
rect 3516 36314 3568 36320
rect 3516 36236 3568 36242
rect 3516 36178 3568 36184
rect 3424 36032 3476 36038
rect 3424 35974 3476 35980
rect 3436 34746 3464 35974
rect 3424 34740 3476 34746
rect 3528 34728 3556 36178
rect 3804 36106 3832 36518
rect 3792 36100 3844 36106
rect 3792 36042 3844 36048
rect 3896 36038 3924 36858
rect 3974 36272 4030 36281
rect 3974 36207 4030 36216
rect 3988 36174 4016 36207
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3884 36032 3936 36038
rect 3884 35974 3936 35980
rect 3662 35932 3970 35941
rect 3662 35930 3668 35932
rect 3724 35930 3748 35932
rect 3804 35930 3828 35932
rect 3884 35930 3908 35932
rect 3964 35930 3970 35932
rect 3724 35878 3726 35930
rect 3906 35878 3908 35930
rect 3662 35876 3668 35878
rect 3724 35876 3748 35878
rect 3804 35876 3828 35878
rect 3884 35876 3908 35878
rect 3964 35876 3970 35878
rect 3662 35867 3970 35876
rect 4080 35766 4108 38270
rect 4264 37806 4292 39238
rect 4322 38652 4630 38661
rect 4322 38650 4328 38652
rect 4384 38650 4408 38652
rect 4464 38650 4488 38652
rect 4544 38650 4568 38652
rect 4624 38650 4630 38652
rect 4384 38598 4386 38650
rect 4566 38598 4568 38650
rect 4322 38596 4328 38598
rect 4384 38596 4408 38598
rect 4464 38596 4488 38598
rect 4544 38596 4568 38598
rect 4624 38596 4630 38598
rect 4322 38587 4630 38596
rect 4344 38548 4396 38554
rect 4344 38490 4396 38496
rect 4252 37800 4304 37806
rect 4252 37742 4304 37748
rect 4356 37652 4384 38490
rect 4436 38412 4488 38418
rect 4436 38354 4488 38360
rect 4448 37738 4476 38354
rect 4724 38010 4752 39442
rect 4816 38350 4844 39782
rect 4908 38554 4936 39918
rect 5000 39902 5212 39930
rect 4988 39840 5040 39846
rect 4988 39782 5040 39788
rect 5000 39642 5028 39782
rect 4988 39636 5040 39642
rect 4988 39578 5040 39584
rect 5080 39568 5132 39574
rect 5080 39510 5132 39516
rect 4986 39128 5042 39137
rect 4986 39063 5042 39072
rect 4896 38548 4948 38554
rect 4896 38490 4948 38496
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 4712 38004 4764 38010
rect 4712 37946 4764 37952
rect 4528 37936 4580 37942
rect 4528 37878 4580 37884
rect 4540 37738 4568 37878
rect 4804 37800 4856 37806
rect 4856 37760 4936 37788
rect 4804 37742 4856 37748
rect 4436 37732 4488 37738
rect 4436 37674 4488 37680
rect 4528 37732 4580 37738
rect 4528 37674 4580 37680
rect 4264 37624 4384 37652
rect 4620 37664 4672 37670
rect 4264 37448 4292 37624
rect 4672 37641 4844 37652
rect 4672 37632 4858 37641
rect 4672 37624 4802 37632
rect 4620 37606 4672 37612
rect 4322 37564 4630 37573
rect 4802 37567 4858 37576
rect 4322 37562 4328 37564
rect 4384 37562 4408 37564
rect 4464 37562 4488 37564
rect 4544 37562 4568 37564
rect 4624 37562 4630 37564
rect 4384 37510 4386 37562
rect 4566 37510 4568 37562
rect 4322 37508 4328 37510
rect 4384 37508 4408 37510
rect 4464 37508 4488 37510
rect 4544 37508 4568 37510
rect 4624 37508 4630 37510
rect 4322 37499 4630 37508
rect 4264 37420 4568 37448
rect 4434 37360 4490 37369
rect 4434 37295 4490 37304
rect 4160 37256 4212 37262
rect 4160 37198 4212 37204
rect 4342 37224 4398 37233
rect 4172 36242 4200 37198
rect 4448 37194 4476 37295
rect 4342 37159 4398 37168
rect 4436 37188 4488 37194
rect 4356 36650 4384 37159
rect 4436 37130 4488 37136
rect 4252 36644 4304 36650
rect 4252 36586 4304 36592
rect 4344 36644 4396 36650
rect 4344 36586 4396 36592
rect 4264 36242 4292 36586
rect 4540 36582 4568 37420
rect 4908 37274 4936 37760
rect 4816 37262 4936 37274
rect 4804 37256 4936 37262
rect 4856 37246 4936 37256
rect 4804 37198 4856 37204
rect 4896 36848 4948 36854
rect 5000 36825 5028 39063
rect 5092 38962 5120 39510
rect 5080 38956 5132 38962
rect 5080 38898 5132 38904
rect 5080 38752 5132 38758
rect 5080 38694 5132 38700
rect 5092 37330 5120 38694
rect 5184 37505 5212 39902
rect 5368 39846 5396 40990
rect 5460 40594 5488 41958
rect 5552 40934 5580 43500
rect 6656 42838 6684 43500
rect 7196 43376 7248 43382
rect 7196 43318 7248 43324
rect 6644 42832 6696 42838
rect 6644 42774 6696 42780
rect 6184 42764 6236 42770
rect 6184 42706 6236 42712
rect 6276 42764 6328 42770
rect 6276 42706 6328 42712
rect 5632 42560 5684 42566
rect 5632 42502 5684 42508
rect 5816 42560 5868 42566
rect 5816 42502 5868 42508
rect 5644 41750 5672 42502
rect 5724 42356 5776 42362
rect 5724 42298 5776 42304
rect 5632 41744 5684 41750
rect 5632 41686 5684 41692
rect 5736 41614 5764 42298
rect 5724 41608 5776 41614
rect 5724 41550 5776 41556
rect 5632 41472 5684 41478
rect 5632 41414 5684 41420
rect 5540 40928 5592 40934
rect 5644 40905 5672 41414
rect 5540 40870 5592 40876
rect 5630 40896 5686 40905
rect 5630 40831 5686 40840
rect 5540 40656 5592 40662
rect 5540 40598 5592 40604
rect 5448 40588 5500 40594
rect 5448 40530 5500 40536
rect 5356 39840 5408 39846
rect 5356 39782 5408 39788
rect 5368 38654 5396 39782
rect 5368 38626 5488 38654
rect 5262 38584 5318 38593
rect 5262 38519 5264 38528
rect 5316 38519 5318 38528
rect 5264 38490 5316 38496
rect 5356 38480 5408 38486
rect 5356 38422 5408 38428
rect 5368 38010 5396 38422
rect 5460 38049 5488 38626
rect 5552 38418 5580 40598
rect 5644 40089 5672 40831
rect 5630 40080 5686 40089
rect 5630 40015 5686 40024
rect 5540 38412 5592 38418
rect 5540 38354 5592 38360
rect 5446 38040 5502 38049
rect 5264 38004 5316 38010
rect 5264 37946 5316 37952
rect 5356 38004 5408 38010
rect 5446 37975 5502 37984
rect 5356 37946 5408 37952
rect 5170 37496 5226 37505
rect 5170 37431 5226 37440
rect 5170 37360 5226 37369
rect 5080 37324 5132 37330
rect 5170 37295 5226 37304
rect 5080 37266 5132 37272
rect 4896 36790 4948 36796
rect 4986 36816 5042 36825
rect 4528 36576 4580 36582
rect 4528 36518 4580 36524
rect 4712 36576 4764 36582
rect 4712 36518 4764 36524
rect 4322 36476 4630 36485
rect 4322 36474 4328 36476
rect 4384 36474 4408 36476
rect 4464 36474 4488 36476
rect 4544 36474 4568 36476
rect 4624 36474 4630 36476
rect 4384 36422 4386 36474
rect 4566 36422 4568 36474
rect 4322 36420 4328 36422
rect 4384 36420 4408 36422
rect 4464 36420 4488 36422
rect 4544 36420 4568 36422
rect 4624 36420 4630 36422
rect 4322 36411 4630 36420
rect 4160 36236 4212 36242
rect 4160 36178 4212 36184
rect 4252 36236 4304 36242
rect 4252 36178 4304 36184
rect 4344 36236 4396 36242
rect 4344 36178 4396 36184
rect 4160 36100 4212 36106
rect 4160 36042 4212 36048
rect 3792 35760 3844 35766
rect 3792 35702 3844 35708
rect 4068 35760 4120 35766
rect 4068 35702 4120 35708
rect 3608 35488 3660 35494
rect 3608 35430 3660 35436
rect 3620 35329 3648 35430
rect 3606 35320 3662 35329
rect 3606 35255 3662 35264
rect 3804 35086 3832 35702
rect 3884 35692 3936 35698
rect 3884 35634 3936 35640
rect 3976 35692 4028 35698
rect 3976 35634 4028 35640
rect 3896 35154 3924 35634
rect 3988 35170 4016 35634
rect 4066 35456 4122 35465
rect 4066 35391 4122 35400
rect 4080 35290 4108 35391
rect 4172 35290 4200 36042
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 4160 35284 4212 35290
rect 4160 35226 4212 35232
rect 4264 35222 4292 36178
rect 4356 35494 4384 36178
rect 4724 35873 4752 36518
rect 4804 36372 4856 36378
rect 4804 36314 4856 36320
rect 4710 35864 4766 35873
rect 4710 35799 4766 35808
rect 4712 35556 4764 35562
rect 4712 35498 4764 35504
rect 4344 35488 4396 35494
rect 4344 35430 4396 35436
rect 4322 35388 4630 35397
rect 4322 35386 4328 35388
rect 4384 35386 4408 35388
rect 4464 35386 4488 35388
rect 4544 35386 4568 35388
rect 4624 35386 4630 35388
rect 4384 35334 4386 35386
rect 4566 35334 4568 35386
rect 4322 35332 4328 35334
rect 4384 35332 4408 35334
rect 4464 35332 4488 35334
rect 4544 35332 4568 35334
rect 4624 35332 4630 35334
rect 4322 35323 4630 35332
rect 4724 35290 4752 35498
rect 4344 35284 4396 35290
rect 4344 35226 4396 35232
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 4252 35216 4304 35222
rect 3884 35148 3936 35154
rect 3988 35142 4200 35170
rect 4252 35158 4304 35164
rect 3884 35090 3936 35096
rect 3792 35080 3844 35086
rect 3792 35022 3844 35028
rect 3896 34932 3924 35090
rect 4172 35057 4200 35142
rect 4158 35048 4214 35057
rect 4158 34983 4214 34992
rect 3896 34904 4032 34932
rect 3662 34844 3970 34853
rect 3662 34842 3668 34844
rect 3724 34842 3748 34844
rect 3804 34842 3828 34844
rect 3884 34842 3908 34844
rect 3964 34842 3970 34844
rect 3724 34790 3726 34842
rect 3906 34790 3908 34842
rect 3662 34788 3668 34790
rect 3724 34788 3748 34790
rect 3804 34788 3828 34790
rect 3884 34788 3908 34790
rect 3964 34788 3970 34790
rect 3662 34779 3970 34788
rect 3700 34740 3752 34746
rect 3528 34700 3648 34728
rect 3424 34682 3476 34688
rect 3422 34504 3478 34513
rect 3422 34439 3478 34448
rect 3516 34468 3568 34474
rect 3436 34406 3464 34439
rect 3516 34410 3568 34416
rect 3424 34400 3476 34406
rect 3424 34342 3476 34348
rect 3332 34196 3384 34202
rect 3332 34138 3384 34144
rect 3240 34128 3292 34134
rect 3240 34070 3292 34076
rect 3424 34060 3476 34066
rect 3424 34002 3476 34008
rect 3330 33960 3386 33969
rect 3160 33918 3280 33946
rect 3056 33448 3108 33454
rect 3056 33390 3108 33396
rect 3148 33380 3200 33386
rect 3148 33322 3200 33328
rect 3056 33312 3108 33318
rect 3056 33254 3108 33260
rect 3068 33046 3096 33254
rect 3056 33040 3108 33046
rect 3056 32982 3108 32988
rect 3160 31346 3188 33322
rect 3252 32230 3280 33918
rect 3330 33895 3386 33904
rect 3344 32450 3372 33895
rect 3436 33046 3464 34002
rect 3528 33522 3556 34410
rect 3620 34202 3648 34700
rect 4004 34728 4032 34904
rect 3700 34682 3752 34688
rect 3804 34700 4032 34728
rect 4066 34776 4122 34785
rect 4066 34711 4122 34720
rect 3712 34406 3740 34682
rect 3804 34610 3832 34700
rect 4080 34660 4108 34711
rect 3988 34632 4108 34660
rect 3792 34604 3844 34610
rect 3792 34546 3844 34552
rect 3700 34400 3752 34406
rect 3804 34377 3832 34546
rect 3700 34342 3752 34348
rect 3790 34368 3846 34377
rect 3712 34241 3740 34342
rect 3790 34303 3846 34312
rect 3698 34232 3754 34241
rect 3608 34196 3660 34202
rect 3698 34167 3754 34176
rect 3608 34138 3660 34144
rect 3988 34066 4016 34632
rect 4264 34610 4292 35158
rect 4356 35086 4384 35226
rect 4344 35080 4396 35086
rect 4344 35022 4396 35028
rect 4252 34604 4304 34610
rect 4252 34546 4304 34552
rect 4356 34490 4384 35022
rect 4712 34944 4764 34950
rect 4712 34886 4764 34892
rect 4724 34678 4752 34886
rect 4712 34672 4764 34678
rect 4712 34614 4764 34620
rect 4068 34468 4120 34474
rect 4068 34410 4120 34416
rect 4264 34462 4384 34490
rect 3976 34060 4028 34066
rect 3976 34002 4028 34008
rect 3974 33960 4030 33969
rect 3974 33895 4030 33904
rect 3988 33862 4016 33895
rect 4080 33862 4108 34410
rect 4160 34400 4212 34406
rect 4160 34342 4212 34348
rect 3976 33856 4028 33862
rect 3976 33798 4028 33804
rect 4068 33856 4120 33862
rect 4068 33798 4120 33804
rect 3662 33756 3970 33765
rect 3662 33754 3668 33756
rect 3724 33754 3748 33756
rect 3804 33754 3828 33756
rect 3884 33754 3908 33756
rect 3964 33754 3970 33756
rect 3724 33702 3726 33754
rect 3906 33702 3908 33754
rect 3662 33700 3668 33702
rect 3724 33700 3748 33702
rect 3804 33700 3828 33702
rect 3884 33700 3908 33702
rect 3964 33700 3970 33702
rect 3662 33691 3970 33700
rect 4080 33658 4108 33798
rect 4068 33652 4120 33658
rect 4068 33594 4120 33600
rect 3516 33516 3568 33522
rect 3516 33458 3568 33464
rect 3700 33448 3752 33454
rect 3700 33390 3752 33396
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3436 32774 3464 32982
rect 3712 32842 3740 33390
rect 3700 32836 3752 32842
rect 3700 32778 3752 32784
rect 3424 32768 3476 32774
rect 3424 32710 3476 32716
rect 3662 32668 3970 32677
rect 3662 32666 3668 32668
rect 3724 32666 3748 32668
rect 3804 32666 3828 32668
rect 3884 32666 3908 32668
rect 3964 32666 3970 32668
rect 3724 32614 3726 32666
rect 3906 32614 3908 32666
rect 3662 32612 3668 32614
rect 3724 32612 3748 32614
rect 3804 32612 3828 32614
rect 3884 32612 3908 32614
rect 3964 32612 3970 32614
rect 3662 32603 3970 32612
rect 3344 32422 3648 32450
rect 3620 32366 3648 32422
rect 4080 32366 4108 33594
rect 4172 33386 4200 34342
rect 4264 33930 4292 34462
rect 4712 34400 4764 34406
rect 4712 34342 4764 34348
rect 4322 34300 4630 34309
rect 4322 34298 4328 34300
rect 4384 34298 4408 34300
rect 4464 34298 4488 34300
rect 4544 34298 4568 34300
rect 4624 34298 4630 34300
rect 4384 34246 4386 34298
rect 4566 34246 4568 34298
rect 4322 34244 4328 34246
rect 4384 34244 4408 34246
rect 4464 34244 4488 34246
rect 4544 34244 4568 34246
rect 4624 34244 4630 34246
rect 4322 34235 4630 34244
rect 4724 34082 4752 34342
rect 4540 34066 4752 34082
rect 4528 34060 4752 34066
rect 4580 34054 4752 34060
rect 4528 34002 4580 34008
rect 4816 33980 4844 36314
rect 4908 35465 4936 36790
rect 4986 36751 5042 36760
rect 4988 36712 5040 36718
rect 4988 36654 5040 36660
rect 5000 36009 5028 36654
rect 5080 36644 5132 36650
rect 5080 36586 5132 36592
rect 4986 36000 5042 36009
rect 4986 35935 5042 35944
rect 4988 35556 5040 35562
rect 4988 35498 5040 35504
rect 4894 35456 4950 35465
rect 4894 35391 4950 35400
rect 4908 35154 4936 35391
rect 4896 35148 4948 35154
rect 4896 35090 4948 35096
rect 5000 34950 5028 35498
rect 4988 34944 5040 34950
rect 4894 34912 4950 34921
rect 4988 34886 5040 34892
rect 4894 34847 4950 34856
rect 4724 33952 4844 33980
rect 4252 33924 4304 33930
rect 4252 33866 4304 33872
rect 4160 33380 4212 33386
rect 4160 33322 4212 33328
rect 4252 33312 4304 33318
rect 4252 33254 4304 33260
rect 4264 32434 4292 33254
rect 4322 33212 4630 33221
rect 4322 33210 4328 33212
rect 4384 33210 4408 33212
rect 4464 33210 4488 33212
rect 4544 33210 4568 33212
rect 4624 33210 4630 33212
rect 4384 33158 4386 33210
rect 4566 33158 4568 33210
rect 4322 33156 4328 33158
rect 4384 33156 4408 33158
rect 4464 33156 4488 33158
rect 4544 33156 4568 33158
rect 4624 33156 4630 33158
rect 4322 33147 4630 33156
rect 4436 32836 4488 32842
rect 4436 32778 4488 32784
rect 4448 32745 4476 32778
rect 4434 32736 4490 32745
rect 4434 32671 4490 32680
rect 4252 32428 4304 32434
rect 4252 32370 4304 32376
rect 4448 32366 4476 32671
rect 3332 32360 3384 32366
rect 3332 32302 3384 32308
rect 3608 32360 3660 32366
rect 3608 32302 3660 32308
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 4436 32360 4488 32366
rect 4436 32302 4488 32308
rect 3240 32224 3292 32230
rect 3240 32166 3292 32172
rect 3252 31822 3280 32166
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 3240 31476 3292 31482
rect 3240 31418 3292 31424
rect 3148 31340 3200 31346
rect 3148 31282 3200 31288
rect 3148 31204 3200 31210
rect 3148 31146 3200 31152
rect 3056 31136 3108 31142
rect 3160 31113 3188 31146
rect 3056 31078 3108 31084
rect 3146 31104 3202 31113
rect 3068 30954 3096 31078
rect 3146 31039 3202 31048
rect 3068 30926 3188 30954
rect 3160 30802 3188 30926
rect 3148 30796 3200 30802
rect 3148 30738 3200 30744
rect 3160 30138 3188 30738
rect 3252 30258 3280 31418
rect 3344 31362 3372 32302
rect 3792 32224 3844 32230
rect 3792 32166 3844 32172
rect 4160 32224 4212 32230
rect 4160 32166 4212 32172
rect 4252 32224 4304 32230
rect 4252 32166 4304 32172
rect 3804 31958 3832 32166
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 3424 31816 3476 31822
rect 3424 31758 3476 31764
rect 3436 31482 3464 31758
rect 4172 31754 4200 32166
rect 4264 32008 4292 32166
rect 4322 32124 4630 32133
rect 4322 32122 4328 32124
rect 4384 32122 4408 32124
rect 4464 32122 4488 32124
rect 4544 32122 4568 32124
rect 4624 32122 4630 32124
rect 4384 32070 4386 32122
rect 4566 32070 4568 32122
rect 4322 32068 4328 32070
rect 4384 32068 4408 32070
rect 4464 32068 4488 32070
rect 4544 32068 4568 32070
rect 4624 32068 4630 32070
rect 4322 32059 4630 32068
rect 4264 31980 4568 32008
rect 4160 31748 4212 31754
rect 4160 31690 4212 31696
rect 4068 31680 4120 31686
rect 3514 31648 3570 31657
rect 4436 31680 4488 31686
rect 4068 31622 4120 31628
rect 4158 31648 4214 31657
rect 3514 31583 3570 31592
rect 3424 31476 3476 31482
rect 3424 31418 3476 31424
rect 3344 31334 3464 31362
rect 3332 31272 3384 31278
rect 3332 31214 3384 31220
rect 3344 31113 3372 31214
rect 3330 31104 3386 31113
rect 3330 31039 3386 31048
rect 3436 30954 3464 31334
rect 3344 30926 3464 30954
rect 3528 30938 3556 31583
rect 3662 31580 3970 31589
rect 3662 31578 3668 31580
rect 3724 31578 3748 31580
rect 3804 31578 3828 31580
rect 3884 31578 3908 31580
rect 3964 31578 3970 31580
rect 3724 31526 3726 31578
rect 3906 31526 3908 31578
rect 3662 31524 3668 31526
rect 3724 31524 3748 31526
rect 3804 31524 3828 31526
rect 3884 31524 3908 31526
rect 3964 31524 3970 31526
rect 3662 31515 3970 31524
rect 3792 31272 3844 31278
rect 3792 31214 3844 31220
rect 3516 30932 3568 30938
rect 3344 30274 3372 30926
rect 3516 30874 3568 30880
rect 3804 30802 3832 31214
rect 4080 30870 4108 31622
rect 4436 31622 4488 31628
rect 4158 31583 4214 31592
rect 4068 30864 4120 30870
rect 4068 30806 4120 30812
rect 3516 30796 3568 30802
rect 3516 30738 3568 30744
rect 3792 30796 3844 30802
rect 3792 30738 3844 30744
rect 3528 30376 3556 30738
rect 4172 30682 4200 31583
rect 4250 31512 4306 31521
rect 4250 31447 4306 31456
rect 4264 30920 4292 31447
rect 4448 31210 4476 31622
rect 4540 31278 4568 31980
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 4528 31272 4580 31278
rect 4528 31214 4580 31220
rect 4436 31204 4488 31210
rect 4436 31146 4488 31152
rect 4632 31142 4660 31826
rect 4724 31754 4752 33952
rect 4908 33912 4936 34847
rect 4816 33884 4936 33912
rect 4712 31748 4764 31754
rect 4712 31690 4764 31696
rect 4620 31136 4672 31142
rect 4672 31096 4752 31124
rect 4620 31078 4672 31084
rect 4322 31036 4630 31045
rect 4322 31034 4328 31036
rect 4384 31034 4408 31036
rect 4464 31034 4488 31036
rect 4544 31034 4568 31036
rect 4624 31034 4630 31036
rect 4384 30982 4386 31034
rect 4566 30982 4568 31034
rect 4322 30980 4328 30982
rect 4384 30980 4408 30982
rect 4464 30980 4488 30982
rect 4544 30980 4568 30982
rect 4624 30980 4630 30982
rect 4322 30971 4630 30980
rect 4724 30938 4752 31096
rect 4436 30932 4488 30938
rect 4264 30892 4384 30920
rect 4250 30832 4306 30841
rect 4250 30767 4306 30776
rect 4080 30654 4200 30682
rect 3662 30492 3970 30501
rect 3662 30490 3668 30492
rect 3724 30490 3748 30492
rect 3804 30490 3828 30492
rect 3884 30490 3908 30492
rect 3964 30490 3970 30492
rect 3724 30438 3726 30490
rect 3906 30438 3908 30490
rect 3662 30436 3668 30438
rect 3724 30436 3748 30438
rect 3804 30436 3828 30438
rect 3884 30436 3908 30438
rect 3964 30436 3970 30438
rect 3662 30427 3970 30436
rect 3792 30388 3844 30394
rect 3528 30348 3740 30376
rect 3240 30252 3292 30258
rect 3344 30246 3556 30274
rect 3240 30194 3292 30200
rect 3332 30184 3384 30190
rect 3238 30152 3294 30161
rect 3160 30110 3238 30138
rect 3332 30126 3384 30132
rect 3238 30087 3294 30096
rect 2976 30008 3096 30036
rect 3068 29764 3096 30008
rect 2976 29736 3096 29764
rect 2872 29504 2924 29510
rect 2872 29446 2924 29452
rect 2870 29336 2926 29345
rect 2870 29271 2872 29280
rect 2924 29271 2926 29280
rect 2872 29242 2924 29248
rect 2976 29102 3004 29736
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 3054 29472 3110 29481
rect 3054 29407 3110 29416
rect 2964 29096 3016 29102
rect 2964 29038 3016 29044
rect 3068 28994 3096 29407
rect 3160 29073 3188 29650
rect 3146 29064 3202 29073
rect 3146 28999 3202 29008
rect 2976 28966 3096 28994
rect 2872 28416 2924 28422
rect 2872 28358 2924 28364
rect 2778 28248 2834 28257
rect 2778 28183 2834 28192
rect 2688 27532 2740 27538
rect 2688 27474 2740 27480
rect 2608 27390 2728 27418
rect 2700 27316 2728 27390
rect 2700 27288 2820 27316
rect 2504 26444 2556 26450
rect 2504 26386 2556 26392
rect 2596 26444 2648 26450
rect 2596 26386 2648 26392
rect 2410 26344 2466 26353
rect 2410 26279 2466 26288
rect 2412 26240 2464 26246
rect 2412 26182 2464 26188
rect 2424 26042 2452 26182
rect 2412 26036 2464 26042
rect 2412 25978 2464 25984
rect 2410 25936 2466 25945
rect 2410 25871 2466 25880
rect 2424 25294 2452 25871
rect 2516 25430 2544 26386
rect 2608 26042 2636 26386
rect 2792 26314 2820 27288
rect 2780 26308 2832 26314
rect 2780 26250 2832 26256
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2608 25906 2636 25978
rect 2596 25900 2648 25906
rect 2596 25842 2648 25848
rect 2608 25498 2636 25842
rect 2884 25838 2912 28358
rect 2976 26518 3004 28966
rect 3148 28688 3200 28694
rect 3148 28630 3200 28636
rect 3056 28008 3108 28014
rect 3054 27976 3056 27985
rect 3108 27976 3110 27985
rect 3160 27946 3188 28630
rect 3252 28626 3280 30087
rect 3240 28620 3292 28626
rect 3240 28562 3292 28568
rect 3240 28484 3292 28490
rect 3240 28426 3292 28432
rect 3054 27911 3110 27920
rect 3148 27940 3200 27946
rect 3148 27882 3200 27888
rect 3056 27872 3108 27878
rect 3056 27814 3108 27820
rect 3068 27538 3096 27814
rect 3160 27538 3188 27882
rect 3056 27532 3108 27538
rect 3056 27474 3108 27480
rect 3148 27532 3200 27538
rect 3148 27474 3200 27480
rect 2964 26512 3016 26518
rect 3016 26472 3096 26500
rect 2964 26454 3016 26460
rect 2872 25832 2924 25838
rect 2872 25774 2924 25780
rect 2964 25832 3016 25838
rect 2964 25774 3016 25780
rect 2884 25537 2912 25774
rect 2870 25528 2926 25537
rect 2596 25492 2648 25498
rect 2870 25463 2926 25472
rect 2596 25434 2648 25440
rect 2504 25424 2556 25430
rect 2504 25366 2556 25372
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2320 25152 2372 25158
rect 2320 25094 2372 25100
rect 2332 24750 2360 25094
rect 2320 24744 2372 24750
rect 2136 24686 2188 24692
rect 2226 24712 2282 24721
rect 2320 24686 2372 24692
rect 2226 24647 2282 24656
rect 2056 24568 2360 24596
rect 1964 24398 2176 24426
rect 2042 24304 2098 24313
rect 1952 24268 2004 24274
rect 2042 24239 2098 24248
rect 1952 24210 2004 24216
rect 1964 22574 1992 24210
rect 1952 22568 2004 22574
rect 1952 22510 2004 22516
rect 2056 21457 2084 24239
rect 2042 21448 2098 21457
rect 2042 21383 2098 21392
rect 2042 21040 2098 21049
rect 2042 20975 2098 20984
rect 1950 20904 2006 20913
rect 1950 20839 2006 20848
rect 1964 19446 1992 20839
rect 2056 19854 2084 20975
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2042 19680 2098 19689
rect 2042 19615 2098 19624
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 1952 19304 2004 19310
rect 1952 19246 2004 19252
rect 1964 18766 1992 19246
rect 1952 18760 2004 18766
rect 1952 18702 2004 18708
rect 1950 17640 2006 17649
rect 1950 17575 2006 17584
rect 1964 17066 1992 17575
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1964 16697 1992 17002
rect 1950 16688 2006 16697
rect 1950 16623 2006 16632
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1964 15042 1992 16186
rect 2056 15609 2084 19615
rect 2148 18970 2176 24398
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 2240 22642 2268 24006
rect 2332 23497 2360 24568
rect 2318 23488 2374 23497
rect 2318 23423 2374 23432
rect 2318 23352 2374 23361
rect 2318 23287 2374 23296
rect 2332 23186 2360 23287
rect 2320 23180 2372 23186
rect 2320 23122 2372 23128
rect 2228 22636 2280 22642
rect 2228 22578 2280 22584
rect 2332 22137 2360 23122
rect 2424 23066 2452 25230
rect 2516 23186 2544 25366
rect 2872 25220 2924 25226
rect 2872 25162 2924 25168
rect 2780 25152 2832 25158
rect 2780 25094 2832 25100
rect 2792 24750 2820 25094
rect 2780 24744 2832 24750
rect 2780 24686 2832 24692
rect 2780 24268 2832 24274
rect 2780 24210 2832 24216
rect 2792 23254 2820 24210
rect 2780 23248 2832 23254
rect 2686 23216 2742 23225
rect 2504 23180 2556 23186
rect 2780 23190 2832 23196
rect 2686 23151 2742 23160
rect 2504 23122 2556 23128
rect 2424 23038 2544 23066
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2318 22128 2374 22137
rect 2424 22098 2452 22918
rect 2318 22063 2374 22072
rect 2412 22092 2464 22098
rect 2412 22034 2464 22040
rect 2410 21992 2466 22001
rect 2410 21927 2466 21936
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2240 21486 2268 21830
rect 2228 21480 2280 21486
rect 2228 21422 2280 21428
rect 2240 20942 2268 21422
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2332 21010 2360 21286
rect 2424 21146 2452 21927
rect 2516 21486 2544 23038
rect 2596 22636 2648 22642
rect 2596 22578 2648 22584
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2412 21140 2464 21146
rect 2412 21082 2464 21088
rect 2320 21004 2372 21010
rect 2320 20946 2372 20952
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2148 18154 2176 18702
rect 2240 18222 2268 20878
rect 2332 19825 2360 20946
rect 2516 20890 2544 21422
rect 2608 21185 2636 22578
rect 2700 22030 2728 23151
rect 2780 22976 2832 22982
rect 2778 22944 2780 22953
rect 2832 22944 2834 22953
rect 2778 22879 2834 22888
rect 2884 22794 2912 25162
rect 2976 24018 3004 25774
rect 3068 25226 3096 26472
rect 3252 26432 3280 28426
rect 3160 26404 3280 26432
rect 3160 25974 3188 26404
rect 3240 26308 3292 26314
rect 3240 26250 3292 26256
rect 3148 25968 3200 25974
rect 3148 25910 3200 25916
rect 3148 25832 3200 25838
rect 3148 25774 3200 25780
rect 3160 25498 3188 25774
rect 3148 25492 3200 25498
rect 3148 25434 3200 25440
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3148 25220 3200 25226
rect 3148 25162 3200 25168
rect 2976 23990 3096 24018
rect 2962 23896 3018 23905
rect 2962 23831 3018 23840
rect 2792 22766 2912 22794
rect 2976 22778 3004 23831
rect 3068 23662 3096 23990
rect 3056 23656 3108 23662
rect 3160 23633 3188 25162
rect 3056 23598 3108 23604
rect 3146 23624 3202 23633
rect 3146 23559 3202 23568
rect 3054 23488 3110 23497
rect 3054 23423 3110 23432
rect 2964 22772 3016 22778
rect 2688 22024 2740 22030
rect 2688 21966 2740 21972
rect 2792 21622 2820 22766
rect 2964 22714 3016 22720
rect 2870 22672 2926 22681
rect 2870 22607 2926 22616
rect 2780 21616 2832 21622
rect 2780 21558 2832 21564
rect 2594 21176 2650 21185
rect 2594 21111 2650 21120
rect 2424 20862 2544 20890
rect 2424 20398 2452 20862
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2412 20392 2464 20398
rect 2412 20334 2464 20340
rect 2412 19984 2464 19990
rect 2410 19952 2412 19961
rect 2464 19952 2466 19961
rect 2410 19887 2466 19896
rect 2318 19816 2374 19825
rect 2318 19751 2374 19760
rect 2318 19272 2374 19281
rect 2318 19207 2374 19216
rect 2332 19174 2360 19207
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2332 18222 2360 18770
rect 2424 18714 2452 19887
rect 2516 19854 2544 20742
rect 2594 20632 2650 20641
rect 2594 20567 2650 20576
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2504 19712 2556 19718
rect 2608 19700 2636 20567
rect 2688 20528 2740 20534
rect 2792 20516 2820 21558
rect 2740 20488 2820 20516
rect 2688 20470 2740 20476
rect 2688 20052 2740 20058
rect 2688 19994 2740 20000
rect 2556 19672 2636 19700
rect 2504 19654 2556 19660
rect 2516 19242 2544 19654
rect 2700 19553 2728 19994
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2792 18970 2820 20488
rect 2884 19825 2912 22607
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2976 21962 3004 22510
rect 2964 21956 3016 21962
rect 2964 21898 3016 21904
rect 2962 21584 3018 21593
rect 2962 21519 2964 21528
rect 3016 21519 3018 21528
rect 2964 21490 3016 21496
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 19894 3004 21286
rect 3068 21146 3096 23423
rect 3252 23338 3280 26250
rect 3160 23310 3280 23338
rect 3160 22710 3188 23310
rect 3240 23248 3292 23254
rect 3240 23190 3292 23196
rect 3148 22704 3200 22710
rect 3148 22646 3200 22652
rect 3148 22568 3200 22574
rect 3148 22510 3200 22516
rect 3160 22234 3188 22510
rect 3148 22228 3200 22234
rect 3148 22170 3200 22176
rect 3160 21457 3188 22170
rect 3252 22166 3280 23190
rect 3240 22160 3292 22166
rect 3238 22128 3240 22137
rect 3292 22128 3294 22137
rect 3238 22063 3294 22072
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3344 21842 3372 30126
rect 3424 30048 3476 30054
rect 3424 29990 3476 29996
rect 3436 29730 3464 29990
rect 3528 29850 3556 30246
rect 3516 29844 3568 29850
rect 3516 29786 3568 29792
rect 3436 29702 3556 29730
rect 3620 29714 3648 30348
rect 3712 30190 3740 30348
rect 3792 30330 3844 30336
rect 3700 30184 3752 30190
rect 3700 30126 3752 30132
rect 3804 30036 3832 30330
rect 3974 30152 4030 30161
rect 3974 30087 3976 30096
rect 4028 30087 4030 30096
rect 3976 30058 4028 30064
rect 3712 30008 3832 30036
rect 3884 30048 3936 30054
rect 3424 29640 3476 29646
rect 3424 29582 3476 29588
rect 3436 29481 3464 29582
rect 3422 29472 3478 29481
rect 3422 29407 3478 29416
rect 3422 29200 3478 29209
rect 3422 29135 3478 29144
rect 3436 29102 3464 29135
rect 3424 29096 3476 29102
rect 3424 29038 3476 29044
rect 3424 28960 3476 28966
rect 3424 28902 3476 28908
rect 3436 28082 3464 28902
rect 3424 28076 3476 28082
rect 3424 28018 3476 28024
rect 3436 27674 3464 28018
rect 3424 27668 3476 27674
rect 3424 27610 3476 27616
rect 3424 27532 3476 27538
rect 3424 27474 3476 27480
rect 3436 25838 3464 27474
rect 3528 26314 3556 29702
rect 3608 29708 3660 29714
rect 3608 29650 3660 29656
rect 3712 29617 3740 30008
rect 3884 29990 3936 29996
rect 3974 30016 4030 30025
rect 3790 29880 3846 29889
rect 3790 29815 3792 29824
rect 3844 29815 3846 29824
rect 3792 29786 3844 29792
rect 3698 29608 3754 29617
rect 3698 29543 3754 29552
rect 3896 29492 3924 29990
rect 3974 29951 4030 29960
rect 3988 29646 4016 29951
rect 4080 29782 4108 30654
rect 4160 30320 4212 30326
rect 4160 30262 4212 30268
rect 4172 30190 4200 30262
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4172 29850 4200 30126
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 4068 29776 4120 29782
rect 4068 29718 4120 29724
rect 4264 29714 4292 30767
rect 4356 30161 4384 30892
rect 4436 30874 4488 30880
rect 4712 30932 4764 30938
rect 4712 30874 4764 30880
rect 4448 30376 4476 30874
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4712 30592 4764 30598
rect 4712 30534 4764 30540
rect 4448 30348 4568 30376
rect 4434 30288 4490 30297
rect 4434 30223 4490 30232
rect 4448 30190 4476 30223
rect 4436 30184 4488 30190
rect 4342 30152 4398 30161
rect 4436 30126 4488 30132
rect 4342 30087 4398 30096
rect 4540 30054 4568 30348
rect 4632 30161 4660 30534
rect 4724 30326 4752 30534
rect 4712 30320 4764 30326
rect 4816 30297 4844 33884
rect 4894 33688 4950 33697
rect 4894 33623 4950 33632
rect 4908 33114 4936 33623
rect 4896 33108 4948 33114
rect 4896 33050 4948 33056
rect 4894 33008 4950 33017
rect 4894 32943 4896 32952
rect 4948 32943 4950 32952
rect 4896 32914 4948 32920
rect 5000 32910 5028 34886
rect 4988 32904 5040 32910
rect 4988 32846 5040 32852
rect 5092 32609 5120 36586
rect 5078 32600 5134 32609
rect 4896 32564 4948 32570
rect 5078 32535 5134 32544
rect 4896 32506 4948 32512
rect 4712 30262 4764 30268
rect 4802 30288 4858 30297
rect 4802 30223 4858 30232
rect 4618 30152 4674 30161
rect 4618 30087 4674 30096
rect 4528 30048 4580 30054
rect 4528 29990 4580 29996
rect 4620 30048 4672 30054
rect 4804 30048 4856 30054
rect 4672 30008 4752 30036
rect 4620 29990 4672 29996
rect 4322 29948 4630 29957
rect 4322 29946 4328 29948
rect 4384 29946 4408 29948
rect 4464 29946 4488 29948
rect 4544 29946 4568 29948
rect 4624 29946 4630 29948
rect 4384 29894 4386 29946
rect 4566 29894 4568 29946
rect 4322 29892 4328 29894
rect 4384 29892 4408 29894
rect 4464 29892 4488 29894
rect 4544 29892 4568 29894
rect 4624 29892 4630 29894
rect 4322 29883 4630 29892
rect 4724 29832 4752 30008
rect 4804 29990 4856 29996
rect 4540 29804 4752 29832
rect 4252 29708 4304 29714
rect 4252 29650 4304 29656
rect 3976 29640 4028 29646
rect 4028 29600 4108 29628
rect 3976 29582 4028 29588
rect 3896 29464 4032 29492
rect 3662 29404 3970 29413
rect 3662 29402 3668 29404
rect 3724 29402 3748 29404
rect 3804 29402 3828 29404
rect 3884 29402 3908 29404
rect 3964 29402 3970 29404
rect 3724 29350 3726 29402
rect 3906 29350 3908 29402
rect 3662 29348 3668 29350
rect 3724 29348 3748 29350
rect 3804 29348 3828 29350
rect 3884 29348 3908 29350
rect 3964 29348 3970 29350
rect 3662 29339 3970 29348
rect 4004 29288 4032 29464
rect 3988 29260 4032 29288
rect 3988 29102 4016 29260
rect 3700 29096 3752 29102
rect 3700 29038 3752 29044
rect 3976 29096 4028 29102
rect 3976 29038 4028 29044
rect 3712 28404 3740 29038
rect 3884 28960 3936 28966
rect 3884 28902 3936 28908
rect 3976 28960 4028 28966
rect 3976 28902 4028 28908
rect 3790 28656 3846 28665
rect 3896 28626 3924 28902
rect 3988 28694 4016 28902
rect 3976 28688 4028 28694
rect 3976 28630 4028 28636
rect 3790 28591 3792 28600
rect 3844 28591 3846 28600
rect 3884 28620 3936 28626
rect 3792 28562 3844 28568
rect 3884 28562 3936 28568
rect 3976 28552 4028 28558
rect 3882 28520 3938 28529
rect 3938 28500 3976 28506
rect 4080 28529 4108 29600
rect 4160 29504 4212 29510
rect 4264 29481 4292 29650
rect 4160 29446 4212 29452
rect 4250 29472 4306 29481
rect 3938 28494 4028 28500
rect 4066 28520 4122 28529
rect 3938 28478 4016 28494
rect 3882 28455 3938 28464
rect 4066 28455 4122 28464
rect 3712 28376 4108 28404
rect 3662 28316 3970 28325
rect 3662 28314 3668 28316
rect 3724 28314 3748 28316
rect 3804 28314 3828 28316
rect 3884 28314 3908 28316
rect 3964 28314 3970 28316
rect 3724 28262 3726 28314
rect 3906 28262 3908 28314
rect 3662 28260 3668 28262
rect 3724 28260 3748 28262
rect 3804 28260 3828 28262
rect 3884 28260 3908 28262
rect 3964 28260 3970 28262
rect 3662 28251 3970 28260
rect 4080 27946 4108 28376
rect 4172 28150 4200 29446
rect 4250 29407 4306 29416
rect 4540 29073 4568 29804
rect 4816 29753 4844 29990
rect 4802 29744 4858 29753
rect 4802 29679 4858 29688
rect 4908 29639 4936 32506
rect 4988 32428 5040 32434
rect 4988 32370 5040 32376
rect 5000 31890 5028 32370
rect 5080 32224 5132 32230
rect 5080 32166 5132 32172
rect 5092 31890 5120 32166
rect 5184 32065 5212 37295
rect 5276 37274 5304 37946
rect 5448 37936 5500 37942
rect 5552 37924 5580 38354
rect 5632 38344 5684 38350
rect 5632 38286 5684 38292
rect 5500 37896 5580 37924
rect 5448 37878 5500 37884
rect 5356 37800 5408 37806
rect 5354 37768 5356 37777
rect 5408 37768 5410 37777
rect 5552 37738 5580 37896
rect 5354 37703 5410 37712
rect 5540 37732 5592 37738
rect 5540 37674 5592 37680
rect 5538 37632 5594 37641
rect 5538 37567 5594 37576
rect 5552 37330 5580 37567
rect 5540 37324 5592 37330
rect 5276 37246 5396 37274
rect 5540 37266 5592 37272
rect 5368 36417 5396 37246
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5448 36780 5500 36786
rect 5448 36722 5500 36728
rect 5354 36408 5410 36417
rect 5354 36343 5410 36352
rect 5460 36038 5488 36722
rect 5552 36145 5580 37130
rect 5644 36650 5672 38286
rect 5736 37670 5764 41550
rect 5828 41002 5856 42502
rect 5908 41676 5960 41682
rect 5908 41618 5960 41624
rect 6000 41676 6052 41682
rect 6000 41618 6052 41624
rect 5920 41070 5948 41618
rect 5908 41064 5960 41070
rect 5908 41006 5960 41012
rect 6012 41018 6040 41618
rect 6196 41614 6224 42706
rect 6184 41608 6236 41614
rect 6184 41550 6236 41556
rect 6012 41002 6132 41018
rect 5816 40996 5868 41002
rect 6012 40996 6144 41002
rect 6012 40990 6092 40996
rect 5816 40938 5868 40944
rect 6092 40938 6144 40944
rect 6196 40934 6224 41550
rect 6000 40928 6052 40934
rect 6000 40870 6052 40876
rect 6184 40928 6236 40934
rect 6184 40870 6236 40876
rect 5908 40384 5960 40390
rect 5908 40326 5960 40332
rect 5920 39982 5948 40326
rect 5908 39976 5960 39982
rect 5908 39918 5960 39924
rect 5908 39432 5960 39438
rect 5908 39374 5960 39380
rect 5816 38888 5868 38894
rect 5816 38830 5868 38836
rect 5828 38418 5856 38830
rect 5920 38457 5948 39374
rect 5906 38448 5962 38457
rect 5816 38412 5868 38418
rect 5906 38383 5962 38392
rect 5816 38354 5868 38360
rect 5816 38276 5868 38282
rect 5816 38218 5868 38224
rect 5724 37664 5776 37670
rect 5724 37606 5776 37612
rect 5632 36644 5684 36650
rect 5632 36586 5684 36592
rect 5630 36544 5686 36553
rect 5630 36479 5686 36488
rect 5644 36242 5672 36479
rect 5632 36236 5684 36242
rect 5632 36178 5684 36184
rect 5538 36136 5594 36145
rect 5828 36106 5856 38218
rect 5908 37664 5960 37670
rect 5908 37606 5960 37612
rect 5920 37466 5948 37606
rect 5908 37460 5960 37466
rect 5908 37402 5960 37408
rect 5908 36576 5960 36582
rect 5908 36518 5960 36524
rect 5920 36310 5948 36518
rect 5908 36304 5960 36310
rect 5908 36246 5960 36252
rect 5538 36071 5594 36080
rect 5816 36100 5868 36106
rect 5816 36042 5868 36048
rect 5448 36032 5500 36038
rect 5448 35974 5500 35980
rect 5354 35864 5410 35873
rect 5354 35799 5410 35808
rect 5264 34944 5316 34950
rect 5368 34921 5396 35799
rect 5460 35601 5488 35974
rect 5814 35864 5870 35873
rect 5814 35799 5870 35808
rect 5724 35624 5776 35630
rect 5446 35592 5502 35601
rect 5446 35527 5502 35536
rect 5630 35592 5686 35601
rect 5724 35566 5776 35572
rect 5630 35527 5632 35536
rect 5684 35527 5686 35536
rect 5632 35498 5684 35504
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 5264 34886 5316 34892
rect 5354 34912 5410 34921
rect 5276 33454 5304 34886
rect 5354 34847 5410 34856
rect 5356 34740 5408 34746
rect 5356 34682 5408 34688
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 5368 33318 5396 34682
rect 5460 34513 5488 34954
rect 5552 34649 5580 35090
rect 5632 35080 5684 35086
rect 5632 35022 5684 35028
rect 5538 34640 5594 34649
rect 5538 34575 5540 34584
rect 5592 34575 5594 34584
rect 5540 34546 5592 34552
rect 5446 34504 5502 34513
rect 5446 34439 5502 34448
rect 5540 34468 5592 34474
rect 5540 34410 5592 34416
rect 5446 34232 5502 34241
rect 5446 34167 5502 34176
rect 5460 33522 5488 34167
rect 5448 33516 5500 33522
rect 5448 33458 5500 33464
rect 5460 33425 5488 33458
rect 5446 33416 5502 33425
rect 5446 33351 5502 33360
rect 5264 33312 5316 33318
rect 5264 33254 5316 33260
rect 5356 33312 5408 33318
rect 5356 33254 5408 33260
rect 5170 32056 5226 32065
rect 5170 31991 5226 32000
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 5080 31884 5132 31890
rect 5080 31826 5132 31832
rect 4986 31784 5042 31793
rect 4986 31719 5042 31728
rect 5000 30190 5028 31719
rect 5276 31226 5304 33254
rect 5368 32978 5396 33254
rect 5552 32994 5580 34410
rect 5644 33998 5672 35022
rect 5632 33992 5684 33998
rect 5632 33934 5684 33940
rect 5630 33688 5686 33697
rect 5630 33623 5686 33632
rect 5356 32972 5408 32978
rect 5356 32914 5408 32920
rect 5460 32966 5580 32994
rect 5460 32910 5488 32966
rect 5448 32904 5500 32910
rect 5354 32872 5410 32881
rect 5448 32846 5500 32852
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5354 32807 5356 32816
rect 5408 32807 5410 32816
rect 5356 32778 5408 32784
rect 5356 32496 5408 32502
rect 5356 32438 5408 32444
rect 5368 31906 5396 32438
rect 5460 32026 5488 32846
rect 5552 32570 5580 32846
rect 5540 32564 5592 32570
rect 5540 32506 5592 32512
rect 5448 32020 5500 32026
rect 5448 31962 5500 31968
rect 5368 31890 5488 31906
rect 5552 31890 5580 32506
rect 5368 31884 5500 31890
rect 5368 31878 5448 31884
rect 5448 31826 5500 31832
rect 5540 31884 5592 31890
rect 5540 31826 5592 31832
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5368 31482 5396 31758
rect 5448 31748 5500 31754
rect 5448 31690 5500 31696
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 5276 31198 5396 31226
rect 5264 31136 5316 31142
rect 5264 31078 5316 31084
rect 5172 30932 5224 30938
rect 5172 30874 5224 30880
rect 5078 30424 5134 30433
rect 5078 30359 5134 30368
rect 4988 30184 5040 30190
rect 4988 30126 5040 30132
rect 5000 29850 5028 30126
rect 4988 29844 5040 29850
rect 4988 29786 5040 29792
rect 5092 29646 5120 30359
rect 4632 29611 4936 29639
rect 5080 29640 5132 29646
rect 4632 29510 4660 29611
rect 5000 29600 5080 29628
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4620 29504 4672 29510
rect 4620 29446 4672 29452
rect 4816 29170 4844 29514
rect 4894 29472 4950 29481
rect 4894 29407 4950 29416
rect 4804 29164 4856 29170
rect 4804 29106 4856 29112
rect 4712 29096 4764 29102
rect 4526 29064 4582 29073
rect 4712 29038 4764 29044
rect 4526 28999 4582 29008
rect 4252 28960 4304 28966
rect 4252 28902 4304 28908
rect 4264 28762 4292 28902
rect 4322 28860 4630 28869
rect 4322 28858 4328 28860
rect 4384 28858 4408 28860
rect 4464 28858 4488 28860
rect 4544 28858 4568 28860
rect 4624 28858 4630 28860
rect 4384 28806 4386 28858
rect 4566 28806 4568 28858
rect 4322 28804 4328 28806
rect 4384 28804 4408 28806
rect 4464 28804 4488 28806
rect 4544 28804 4568 28806
rect 4624 28804 4630 28806
rect 4322 28795 4630 28804
rect 4252 28756 4304 28762
rect 4304 28716 4384 28744
rect 4252 28698 4304 28704
rect 4250 28520 4306 28529
rect 4250 28455 4306 28464
rect 4160 28144 4212 28150
rect 4160 28086 4212 28092
rect 4160 28008 4212 28014
rect 4160 27950 4212 27956
rect 4068 27940 4120 27946
rect 4068 27882 4120 27888
rect 3662 27228 3970 27237
rect 3662 27226 3668 27228
rect 3724 27226 3748 27228
rect 3804 27226 3828 27228
rect 3884 27226 3908 27228
rect 3964 27226 3970 27228
rect 3724 27174 3726 27226
rect 3906 27174 3908 27226
rect 3662 27172 3668 27174
rect 3724 27172 3748 27174
rect 3804 27172 3828 27174
rect 3884 27172 3908 27174
rect 3964 27172 3970 27174
rect 3662 27163 3970 27172
rect 4080 26353 4108 27882
rect 4172 27606 4200 27950
rect 4160 27600 4212 27606
rect 4160 27542 4212 27548
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 26518 4200 26930
rect 4160 26512 4212 26518
rect 4160 26454 4212 26460
rect 4066 26344 4122 26353
rect 3516 26308 3568 26314
rect 4066 26279 4122 26288
rect 3516 26250 3568 26256
rect 3514 26208 3570 26217
rect 3514 26143 3570 26152
rect 3424 25832 3476 25838
rect 3424 25774 3476 25780
rect 3528 25770 3556 26143
rect 3662 26140 3970 26149
rect 3662 26138 3668 26140
rect 3724 26138 3748 26140
rect 3804 26138 3828 26140
rect 3884 26138 3908 26140
rect 3964 26138 3970 26140
rect 3724 26086 3726 26138
rect 3906 26086 3908 26138
rect 3662 26084 3668 26086
rect 3724 26084 3748 26086
rect 3804 26084 3828 26086
rect 3884 26084 3908 26086
rect 3964 26084 3970 26086
rect 3662 26075 3970 26084
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 3974 25936 4030 25945
rect 3974 25871 4030 25880
rect 3988 25838 4016 25871
rect 3700 25832 3752 25838
rect 3700 25774 3752 25780
rect 3976 25832 4028 25838
rect 3976 25774 4028 25780
rect 3516 25764 3568 25770
rect 3516 25706 3568 25712
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 3436 25362 3464 25638
rect 3528 25362 3556 25706
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3516 25356 3568 25362
rect 3516 25298 3568 25304
rect 3436 23662 3464 25298
rect 3712 25226 3740 25774
rect 4080 25498 4108 25978
rect 4172 25838 4200 26454
rect 4264 26246 4292 28455
rect 4356 27946 4384 28716
rect 4724 28694 4752 29038
rect 4712 28688 4764 28694
rect 4712 28630 4764 28636
rect 4528 28552 4580 28558
rect 4528 28494 4580 28500
rect 4434 28248 4490 28257
rect 4434 28183 4436 28192
rect 4488 28183 4490 28192
rect 4436 28154 4488 28160
rect 4434 28112 4490 28121
rect 4434 28047 4490 28056
rect 4540 28064 4568 28494
rect 4802 28112 4858 28121
rect 4620 28076 4672 28082
rect 4448 28014 4476 28047
rect 4540 28036 4620 28064
rect 4802 28047 4858 28056
rect 4620 28018 4672 28024
rect 4436 28008 4488 28014
rect 4436 27950 4488 27956
rect 4344 27940 4396 27946
rect 4344 27882 4396 27888
rect 4620 27872 4672 27878
rect 4672 27832 4752 27860
rect 4620 27814 4672 27820
rect 4322 27772 4630 27781
rect 4322 27770 4328 27772
rect 4384 27770 4408 27772
rect 4464 27770 4488 27772
rect 4544 27770 4568 27772
rect 4624 27770 4630 27772
rect 4384 27718 4386 27770
rect 4566 27718 4568 27770
rect 4322 27716 4328 27718
rect 4384 27716 4408 27718
rect 4464 27716 4488 27718
rect 4544 27716 4568 27718
rect 4624 27716 4630 27718
rect 4322 27707 4630 27716
rect 4344 27668 4396 27674
rect 4344 27610 4396 27616
rect 4356 27538 4384 27610
rect 4344 27532 4396 27538
rect 4344 27474 4396 27480
rect 4356 27334 4384 27474
rect 4620 27396 4672 27402
rect 4620 27338 4672 27344
rect 4344 27328 4396 27334
rect 4344 27270 4396 27276
rect 4632 26897 4660 27338
rect 4724 27062 4752 27832
rect 4816 27674 4844 28047
rect 4804 27668 4856 27674
rect 4804 27610 4856 27616
rect 4908 27538 4936 29407
rect 4896 27532 4948 27538
rect 4816 27492 4896 27520
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4618 26888 4674 26897
rect 4618 26823 4674 26832
rect 4322 26684 4630 26693
rect 4322 26682 4328 26684
rect 4384 26682 4408 26684
rect 4464 26682 4488 26684
rect 4544 26682 4568 26684
rect 4624 26682 4630 26684
rect 4384 26630 4386 26682
rect 4566 26630 4568 26682
rect 4322 26628 4328 26630
rect 4384 26628 4408 26630
rect 4464 26628 4488 26630
rect 4544 26628 4568 26630
rect 4624 26628 4630 26630
rect 4322 26619 4630 26628
rect 4724 26450 4752 26998
rect 4816 26926 4844 27492
rect 4896 27474 4948 27480
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4804 26784 4856 26790
rect 4804 26726 4856 26732
rect 4712 26444 4764 26450
rect 4712 26386 4764 26392
rect 4252 26240 4304 26246
rect 4252 26182 4304 26188
rect 4528 26240 4580 26246
rect 4528 26182 4580 26188
rect 4264 25838 4292 26182
rect 4540 25945 4568 26182
rect 4526 25936 4582 25945
rect 4526 25871 4582 25880
rect 4724 25838 4752 26386
rect 4160 25832 4212 25838
rect 4160 25774 4212 25780
rect 4252 25832 4304 25838
rect 4252 25774 4304 25780
rect 4712 25832 4764 25838
rect 4712 25774 4764 25780
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 3700 25220 3752 25226
rect 3700 25162 3752 25168
rect 3662 25052 3970 25061
rect 3662 25050 3668 25052
rect 3724 25050 3748 25052
rect 3804 25050 3828 25052
rect 3884 25050 3908 25052
rect 3964 25050 3970 25052
rect 3724 24998 3726 25050
rect 3906 24998 3908 25050
rect 3662 24996 3668 24998
rect 3724 24996 3748 24998
rect 3804 24996 3828 24998
rect 3884 24996 3908 24998
rect 3964 24996 3970 24998
rect 3662 24987 3970 24996
rect 3700 24948 3752 24954
rect 3700 24890 3752 24896
rect 3608 24744 3660 24750
rect 3608 24686 3660 24692
rect 3516 24336 3568 24342
rect 3516 24278 3568 24284
rect 3528 23730 3556 24278
rect 3620 24274 3648 24686
rect 3712 24313 3740 24890
rect 3884 24880 3936 24886
rect 3884 24822 3936 24828
rect 3792 24608 3844 24614
rect 3792 24550 3844 24556
rect 3698 24304 3754 24313
rect 3608 24268 3660 24274
rect 3804 24274 3832 24550
rect 3698 24239 3700 24248
rect 3608 24210 3660 24216
rect 3752 24239 3754 24248
rect 3792 24268 3844 24274
rect 3700 24210 3752 24216
rect 3792 24210 3844 24216
rect 3896 24138 3924 24822
rect 4172 24750 4200 25774
rect 4264 24818 4292 25774
rect 4322 25596 4630 25605
rect 4322 25594 4328 25596
rect 4384 25594 4408 25596
rect 4464 25594 4488 25596
rect 4544 25594 4568 25596
rect 4624 25594 4630 25596
rect 4384 25542 4386 25594
rect 4566 25542 4568 25594
rect 4322 25540 4328 25542
rect 4384 25540 4408 25542
rect 4464 25540 4488 25542
rect 4544 25540 4568 25542
rect 4624 25540 4630 25542
rect 4322 25531 4630 25540
rect 4724 25362 4752 25774
rect 4712 25356 4764 25362
rect 4712 25298 4764 25304
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4252 24812 4304 24818
rect 4252 24754 4304 24760
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4172 24410 4200 24686
rect 4160 24404 4212 24410
rect 4160 24346 4212 24352
rect 4264 24274 4292 24754
rect 4632 24664 4660 25162
rect 4724 24886 4752 25298
rect 4816 25226 4844 26726
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4802 24984 4858 24993
rect 4802 24919 4858 24928
rect 4712 24880 4764 24886
rect 4712 24822 4764 24828
rect 4712 24676 4764 24682
rect 4632 24636 4712 24664
rect 4712 24618 4764 24624
rect 4322 24508 4630 24517
rect 4322 24506 4328 24508
rect 4384 24506 4408 24508
rect 4464 24506 4488 24508
rect 4544 24506 4568 24508
rect 4624 24506 4630 24508
rect 4384 24454 4386 24506
rect 4566 24454 4568 24506
rect 4322 24452 4328 24454
rect 4384 24452 4408 24454
rect 4464 24452 4488 24454
rect 4544 24452 4568 24454
rect 4624 24452 4630 24454
rect 4322 24443 4630 24452
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4068 24268 4120 24274
rect 4068 24210 4120 24216
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4080 24177 4108 24210
rect 4066 24168 4122 24177
rect 3884 24132 3936 24138
rect 4632 24138 4660 24346
rect 4066 24103 4122 24112
rect 4160 24132 4212 24138
rect 3884 24074 3936 24080
rect 4160 24074 4212 24080
rect 4620 24132 4672 24138
rect 4620 24074 4672 24080
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 3662 23964 3970 23973
rect 3662 23962 3668 23964
rect 3724 23962 3748 23964
rect 3804 23962 3828 23964
rect 3884 23962 3908 23964
rect 3964 23962 3970 23964
rect 3724 23910 3726 23962
rect 3906 23910 3908 23962
rect 3662 23908 3668 23910
rect 3724 23908 3748 23910
rect 3804 23908 3828 23910
rect 3884 23908 3908 23910
rect 3964 23908 3970 23910
rect 3662 23899 3970 23908
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3424 23656 3476 23662
rect 3424 23598 3476 23604
rect 3424 23520 3476 23526
rect 3424 23462 3476 23468
rect 3436 22001 3464 23462
rect 3516 22976 3568 22982
rect 4080 22953 4108 24006
rect 3516 22918 3568 22924
rect 4066 22944 4122 22953
rect 3528 22642 3556 22918
rect 3662 22876 3970 22885
rect 4066 22879 4122 22888
rect 3662 22874 3668 22876
rect 3724 22874 3748 22876
rect 3804 22874 3828 22876
rect 3884 22874 3908 22876
rect 3964 22874 3970 22876
rect 3724 22822 3726 22874
rect 3906 22822 3908 22874
rect 3662 22820 3668 22822
rect 3724 22820 3748 22822
rect 3804 22820 3828 22822
rect 3884 22820 3908 22822
rect 3964 22820 3970 22822
rect 3662 22811 3970 22820
rect 4172 22778 4200 24074
rect 4528 24064 4580 24070
rect 4528 24006 4580 24012
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 4252 23792 4304 23798
rect 4252 23734 4304 23740
rect 4264 23186 4292 23734
rect 4356 23594 4384 23802
rect 4540 23662 4568 24006
rect 4620 23792 4672 23798
rect 4620 23734 4672 23740
rect 4632 23662 4660 23734
rect 4528 23656 4580 23662
rect 4528 23598 4580 23604
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4344 23588 4396 23594
rect 4344 23530 4396 23536
rect 4322 23420 4630 23429
rect 4322 23418 4328 23420
rect 4384 23418 4408 23420
rect 4464 23418 4488 23420
rect 4544 23418 4568 23420
rect 4624 23418 4630 23420
rect 4384 23366 4386 23418
rect 4566 23366 4568 23418
rect 4322 23364 4328 23366
rect 4384 23364 4408 23366
rect 4464 23364 4488 23366
rect 4544 23364 4568 23366
rect 4624 23364 4630 23366
rect 4322 23355 4630 23364
rect 4436 23248 4488 23254
rect 4434 23216 4436 23225
rect 4488 23216 4490 23225
rect 4252 23180 4304 23186
rect 4434 23151 4490 23160
rect 4252 23122 4304 23128
rect 4618 23080 4674 23089
rect 4618 23015 4674 23024
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 3516 22636 3568 22642
rect 3516 22578 3568 22584
rect 3422 21992 3478 22001
rect 3422 21927 3478 21936
rect 3252 21706 3280 21830
rect 3344 21814 3464 21842
rect 3252 21678 3372 21706
rect 3436 21690 3464 21814
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 3344 21049 3372 21678
rect 3424 21684 3476 21690
rect 3528 21672 3556 22578
rect 3712 22098 3740 22714
rect 4080 22438 4108 22714
rect 4172 22488 4200 22714
rect 4250 22672 4306 22681
rect 4250 22607 4252 22616
rect 4304 22607 4306 22616
rect 4252 22578 4304 22584
rect 4632 22506 4660 23015
rect 4620 22500 4672 22506
rect 4172 22460 4292 22488
rect 4068 22432 4120 22438
rect 4068 22374 4120 22380
rect 4080 22098 4108 22374
rect 4264 22098 4292 22460
rect 4620 22442 4672 22448
rect 4322 22332 4630 22341
rect 4322 22330 4328 22332
rect 4384 22330 4408 22332
rect 4464 22330 4488 22332
rect 4544 22330 4568 22332
rect 4624 22330 4630 22332
rect 4384 22278 4386 22330
rect 4566 22278 4568 22330
rect 4322 22276 4328 22278
rect 4384 22276 4408 22278
rect 4464 22276 4488 22278
rect 4544 22276 4568 22278
rect 4624 22276 4630 22278
rect 4322 22267 4630 22276
rect 4342 22128 4398 22137
rect 3700 22092 3752 22098
rect 3700 22034 3752 22040
rect 4068 22092 4120 22098
rect 4068 22034 4120 22040
rect 4252 22092 4304 22098
rect 4342 22063 4398 22072
rect 4252 22034 4304 22040
rect 4160 21888 4212 21894
rect 4080 21848 4160 21876
rect 3662 21788 3970 21797
rect 3662 21786 3668 21788
rect 3724 21786 3748 21788
rect 3804 21786 3828 21788
rect 3884 21786 3908 21788
rect 3964 21786 3970 21788
rect 3724 21734 3726 21786
rect 3906 21734 3908 21786
rect 3662 21732 3668 21734
rect 3724 21732 3748 21734
rect 3804 21732 3828 21734
rect 3884 21732 3908 21734
rect 3964 21732 3970 21734
rect 3662 21723 3970 21732
rect 3528 21644 3832 21672
rect 3424 21626 3476 21632
rect 3606 21584 3662 21593
rect 3516 21548 3568 21554
rect 3804 21570 3832 21644
rect 3804 21542 4016 21570
rect 3606 21519 3662 21528
rect 3516 21490 3568 21496
rect 3054 21040 3110 21049
rect 3330 21040 3386 21049
rect 3054 20975 3110 20984
rect 3148 21004 3200 21010
rect 3068 20942 3096 20975
rect 3528 21010 3556 21490
rect 3620 21486 3648 21519
rect 3988 21486 4016 21542
rect 3608 21480 3660 21486
rect 3792 21480 3844 21486
rect 3608 21422 3660 21428
rect 3790 21448 3792 21457
rect 3976 21480 4028 21486
rect 3844 21448 3846 21457
rect 3976 21422 4028 21428
rect 3790 21383 3846 21392
rect 3884 21412 3936 21418
rect 3884 21354 3936 21360
rect 3698 21312 3754 21321
rect 3698 21247 3754 21256
rect 3712 21146 3740 21247
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3792 21072 3844 21078
rect 3698 21040 3754 21049
rect 3330 20975 3386 20984
rect 3516 21004 3568 21010
rect 3148 20946 3200 20952
rect 3516 20946 3568 20952
rect 3608 21004 3660 21010
rect 3896 21060 3924 21354
rect 3844 21032 3924 21060
rect 3792 21014 3844 21020
rect 3698 20975 3754 20984
rect 3608 20946 3660 20952
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 3160 20398 3188 20946
rect 3330 20904 3386 20913
rect 3620 20890 3648 20946
rect 3712 20924 3740 20975
rect 3792 20936 3844 20942
rect 3712 20896 3792 20924
rect 3330 20839 3386 20848
rect 3436 20862 3648 20890
rect 3792 20878 3844 20884
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 2976 19866 3188 19894
rect 2870 19816 2926 19825
rect 2870 19751 2926 19760
rect 3054 19816 3110 19825
rect 3160 19786 3188 19866
rect 3054 19751 3056 19760
rect 3108 19751 3110 19760
rect 3148 19780 3200 19786
rect 3056 19722 3108 19728
rect 3148 19722 3200 19728
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 3146 19680 3202 19689
rect 2884 19530 2912 19654
rect 3146 19615 3202 19624
rect 3054 19544 3110 19553
rect 2884 19502 3004 19530
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 2424 18686 2544 18714
rect 2412 18624 2464 18630
rect 2412 18566 2464 18572
rect 2424 18426 2452 18566
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2136 18148 2188 18154
rect 2136 18090 2188 18096
rect 2134 18048 2190 18057
rect 2134 17983 2190 17992
rect 2148 17202 2176 17983
rect 2240 17678 2268 18158
rect 2332 17814 2360 18158
rect 2516 17954 2544 18686
rect 2596 18352 2648 18358
rect 2596 18294 2648 18300
rect 2424 17926 2544 17954
rect 2320 17808 2372 17814
rect 2320 17750 2372 17756
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2134 17096 2190 17105
rect 2134 17031 2136 17040
rect 2188 17031 2190 17040
rect 2136 17002 2188 17008
rect 2136 16584 2188 16590
rect 2136 16526 2188 16532
rect 2148 16250 2176 16526
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2240 16046 2268 17614
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2228 16040 2280 16046
rect 2228 15982 2280 15988
rect 2042 15600 2098 15609
rect 2042 15535 2098 15544
rect 2136 15564 2188 15570
rect 2136 15506 2188 15512
rect 2044 15360 2096 15366
rect 2044 15302 2096 15308
rect 2056 15162 2084 15302
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1964 15014 2084 15042
rect 1952 14884 2004 14890
rect 1952 14826 2004 14832
rect 1964 14414 1992 14826
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1952 13388 2004 13394
rect 2056 13376 2084 15014
rect 2148 14482 2176 15506
rect 2240 15026 2268 15982
rect 2332 15502 2360 17206
rect 2424 17066 2452 17926
rect 2608 17746 2636 18294
rect 2792 18170 2820 18906
rect 2884 18306 2912 19382
rect 2976 19310 3004 19502
rect 3054 19479 3110 19488
rect 2964 19304 3016 19310
rect 2964 19246 3016 19252
rect 3068 19242 3096 19479
rect 3160 19334 3188 19615
rect 3252 19514 3280 20402
rect 3344 20369 3372 20839
rect 3436 20534 3464 20862
rect 3516 20800 3568 20806
rect 3516 20742 3568 20748
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3330 20360 3386 20369
rect 3330 20295 3386 20304
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3344 19378 3372 20198
rect 3528 20058 3556 20742
rect 3662 20700 3970 20709
rect 3662 20698 3668 20700
rect 3724 20698 3748 20700
rect 3804 20698 3828 20700
rect 3884 20698 3908 20700
rect 3964 20698 3970 20700
rect 3724 20646 3726 20698
rect 3906 20646 3908 20698
rect 3662 20644 3668 20646
rect 3724 20644 3748 20646
rect 3804 20644 3828 20646
rect 3884 20644 3908 20646
rect 3964 20644 3970 20646
rect 3662 20635 3970 20644
rect 4080 20641 4108 21848
rect 4160 21830 4212 21836
rect 4160 21616 4212 21622
rect 4160 21558 4212 21564
rect 4066 20632 4122 20641
rect 3700 20596 3752 20602
rect 3700 20538 3752 20544
rect 3792 20596 3844 20602
rect 4066 20567 4122 20576
rect 3792 20538 3844 20544
rect 3712 20330 3740 20538
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3700 20324 3752 20330
rect 3700 20266 3752 20272
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3620 19922 3648 20266
rect 3516 19916 3568 19922
rect 3436 19876 3516 19904
rect 3332 19372 3384 19378
rect 3160 19306 3280 19334
rect 3332 19314 3384 19320
rect 3056 19236 3108 19242
rect 3056 19178 3108 19184
rect 2964 18964 3016 18970
rect 2964 18906 3016 18912
rect 2976 18714 3004 18906
rect 3054 18864 3110 18873
rect 3054 18799 3056 18808
rect 3108 18799 3110 18808
rect 3148 18828 3200 18834
rect 3056 18770 3108 18776
rect 3148 18770 3200 18776
rect 2976 18686 3096 18714
rect 2884 18278 3004 18306
rect 3068 18290 3096 18686
rect 2700 18142 2820 18170
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2596 17740 2648 17746
rect 2596 17682 2648 17688
rect 2700 17626 2728 18142
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2516 17598 2728 17626
rect 2792 17626 2820 18022
rect 2884 17746 2912 18158
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 2792 17598 2912 17626
rect 2412 17060 2464 17066
rect 2412 17002 2464 17008
rect 2516 16794 2544 17598
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2608 17270 2636 17478
rect 2700 17338 2728 17478
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 2596 17264 2648 17270
rect 2596 17206 2648 17212
rect 2594 17096 2650 17105
rect 2594 17031 2650 17040
rect 2412 16788 2464 16794
rect 2412 16730 2464 16736
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2424 16674 2452 16730
rect 2424 16646 2544 16674
rect 2516 16046 2544 16646
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2424 15570 2452 15846
rect 2516 15570 2544 15982
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2136 14476 2188 14482
rect 2136 14418 2188 14424
rect 2228 14408 2280 14414
rect 2332 14362 2360 15438
rect 2412 15428 2464 15434
rect 2412 15370 2464 15376
rect 2424 15162 2452 15370
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2608 14890 2636 17031
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2792 16250 2820 16730
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2686 16144 2742 16153
rect 2686 16079 2688 16088
rect 2740 16079 2742 16088
rect 2688 16050 2740 16056
rect 2688 15564 2740 15570
rect 2792 15552 2820 16186
rect 2740 15524 2820 15552
rect 2688 15506 2740 15512
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2780 15360 2832 15366
rect 2780 15302 2832 15308
rect 2596 14884 2648 14890
rect 2596 14826 2648 14832
rect 2700 14482 2728 15302
rect 2792 14822 2820 15302
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2792 14482 2820 14758
rect 2884 14618 2912 17598
rect 2976 16561 3004 18278
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3056 18148 3108 18154
rect 3056 18090 3108 18096
rect 2962 16552 3018 16561
rect 2962 16487 3018 16496
rect 2962 15328 3018 15337
rect 2962 15263 3018 15272
rect 2872 14612 2924 14618
rect 2872 14554 2924 14560
rect 2976 14498 3004 15263
rect 2688 14476 2740 14482
rect 2280 14356 2360 14362
rect 2228 14350 2360 14356
rect 2240 14334 2360 14350
rect 2332 14074 2360 14334
rect 2424 14436 2688 14464
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2228 13864 2280 13870
rect 2332 13852 2360 14010
rect 2424 13938 2452 14436
rect 2688 14418 2740 14424
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2884 14470 3004 14498
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2280 13824 2360 13852
rect 2504 13864 2556 13870
rect 2228 13806 2280 13812
rect 2504 13806 2556 13812
rect 2004 13348 2084 13376
rect 1952 13330 2004 13336
rect 2056 12782 2084 13348
rect 2044 12776 2096 12782
rect 2044 12718 2096 12724
rect 1950 11248 2006 11257
rect 1950 11183 1952 11192
rect 2004 11183 2006 11192
rect 1952 11154 2004 11160
rect 1964 10606 1992 11154
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1860 10192 1912 10198
rect 1860 10134 1912 10140
rect 1872 9518 1900 10134
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9586 1992 9862
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1124 8356 1176 8362
rect 1124 8298 1176 8304
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 480 6452 532 6458
rect 480 6394 532 6400
rect 952 5545 980 6734
rect 1032 6656 1084 6662
rect 1032 6598 1084 6604
rect 1044 6254 1072 6598
rect 1032 6248 1084 6254
rect 1032 6190 1084 6196
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 1136 5273 1164 8298
rect 1412 6866 1440 8366
rect 1780 8022 1808 8366
rect 1872 8090 1900 8366
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 1504 6186 1532 7278
rect 2148 7274 2176 13806
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2424 13530 2452 13670
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2240 11626 2268 13262
rect 2332 12986 2360 13330
rect 2516 13258 2544 13806
rect 2608 13802 2636 14214
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 2608 13462 2636 13738
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 2792 13394 2820 14418
rect 2884 13410 2912 14470
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13530 3004 13806
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2780 13388 2832 13394
rect 2884 13382 3004 13410
rect 2780 13330 2832 13336
rect 2504 13252 2556 13258
rect 2504 13194 2556 13200
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2792 12918 2820 13330
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12776 2740 12782
rect 2780 12776 2832 12782
rect 2688 12718 2740 12724
rect 2778 12744 2780 12753
rect 2832 12744 2834 12753
rect 2700 12442 2728 12718
rect 2778 12679 2834 12688
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2700 11898 2728 12174
rect 2884 11898 2912 12378
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 2228 11620 2280 11626
rect 2228 11562 2280 11568
rect 2240 11150 2268 11562
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10062 2268 11086
rect 2332 10810 2360 11154
rect 2504 11076 2556 11082
rect 2504 11018 2556 11024
rect 2516 10985 2544 11018
rect 2502 10976 2558 10985
rect 2502 10911 2558 10920
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2976 10606 3004 13382
rect 3068 12442 3096 18090
rect 3160 17882 3188 18770
rect 3252 17882 3280 19306
rect 3436 19145 3464 19876
rect 3516 19858 3568 19864
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3620 19802 3648 19858
rect 3528 19774 3648 19802
rect 3528 19496 3556 19774
rect 3804 19718 3832 20538
rect 3976 20528 4028 20534
rect 3976 20470 4028 20476
rect 3988 20346 4016 20470
rect 4080 20466 4108 20567
rect 4068 20460 4120 20466
rect 4068 20402 4120 20408
rect 3988 20318 4108 20346
rect 4172 20330 4200 21558
rect 4356 21486 4384 22063
rect 4724 21729 4752 24618
rect 4816 23730 4844 24919
rect 4908 24070 4936 27338
rect 5000 27062 5028 29600
rect 5080 29582 5132 29588
rect 5078 29472 5134 29481
rect 5078 29407 5134 29416
rect 5092 29306 5120 29407
rect 5080 29300 5132 29306
rect 5080 29242 5132 29248
rect 5092 27538 5120 29242
rect 5184 29102 5212 30874
rect 5276 30734 5304 31078
rect 5368 30938 5396 31198
rect 5356 30932 5408 30938
rect 5356 30874 5408 30880
rect 5356 30796 5408 30802
rect 5356 30738 5408 30744
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 5276 29578 5304 30670
rect 5368 30025 5396 30738
rect 5354 30016 5410 30025
rect 5354 29951 5410 29960
rect 5460 29850 5488 31690
rect 5552 31414 5580 31826
rect 5540 31408 5592 31414
rect 5540 31350 5592 31356
rect 5552 30598 5580 31350
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5644 30394 5672 33623
rect 5736 30705 5764 35566
rect 5828 35154 5856 35799
rect 6012 35494 6040 40870
rect 6288 40769 6316 42706
rect 6552 42560 6604 42566
rect 6552 42502 6604 42508
rect 6564 42158 6592 42502
rect 6920 42356 6972 42362
rect 6920 42298 6972 42304
rect 6552 42152 6604 42158
rect 6552 42094 6604 42100
rect 6828 42084 6880 42090
rect 6828 42026 6880 42032
rect 6460 42016 6512 42022
rect 6460 41958 6512 41964
rect 6366 41576 6422 41585
rect 6366 41511 6368 41520
rect 6420 41511 6422 41520
rect 6368 41482 6420 41488
rect 6366 41032 6422 41041
rect 6366 40967 6422 40976
rect 6274 40760 6330 40769
rect 6274 40695 6330 40704
rect 6184 40588 6236 40594
rect 6184 40530 6236 40536
rect 6196 39914 6224 40530
rect 6184 39908 6236 39914
rect 6184 39850 6236 39856
rect 6380 39846 6408 40967
rect 6368 39840 6420 39846
rect 6368 39782 6420 39788
rect 6274 39672 6330 39681
rect 6274 39607 6330 39616
rect 6184 39500 6236 39506
rect 6184 39442 6236 39448
rect 6092 38820 6144 38826
rect 6092 38762 6144 38768
rect 6104 37942 6132 38762
rect 6092 37936 6144 37942
rect 6092 37878 6144 37884
rect 6092 36780 6144 36786
rect 6092 36722 6144 36728
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 5998 35320 6054 35329
rect 6104 35306 6132 36722
rect 6196 35766 6224 39442
rect 6288 37754 6316 39607
rect 6472 39137 6500 41958
rect 6736 41744 6788 41750
rect 6642 41712 6698 41721
rect 6736 41686 6788 41692
rect 6642 41647 6698 41656
rect 6550 41440 6606 41449
rect 6550 41375 6606 41384
rect 6458 39128 6514 39137
rect 6458 39063 6514 39072
rect 6564 39001 6592 41375
rect 6656 41206 6684 41647
rect 6748 41206 6776 41686
rect 6644 41200 6696 41206
rect 6644 41142 6696 41148
rect 6736 41200 6788 41206
rect 6736 41142 6788 41148
rect 6644 41064 6696 41070
rect 6644 41006 6696 41012
rect 6840 41018 6868 42026
rect 6932 41274 6960 42298
rect 7208 42158 7236 43318
rect 7484 43110 7512 43574
rect 7746 43500 7802 43560
rect 8298 43500 8354 43900
rect 8850 43616 8906 43900
rect 8850 43500 8906 43560
rect 9402 43616 9458 43900
rect 9402 43500 9458 43560
rect 9954 43500 10010 43900
rect 7472 43104 7524 43110
rect 7472 43046 7524 43052
rect 8312 42906 8340 43500
rect 10048 43376 10100 43382
rect 10048 43318 10100 43324
rect 8668 43172 8720 43178
rect 8668 43114 8720 43120
rect 8300 42900 8352 42906
rect 7852 42860 8156 42888
rect 7748 42832 7800 42838
rect 7852 42820 7880 42860
rect 7800 42792 7880 42820
rect 7748 42774 7800 42780
rect 8128 42786 8156 42860
rect 8300 42842 8352 42848
rect 7472 42764 7524 42770
rect 7472 42706 7524 42712
rect 7288 42696 7340 42702
rect 7484 42673 7512 42706
rect 7288 42638 7340 42644
rect 7470 42664 7526 42673
rect 7196 42152 7248 42158
rect 7196 42094 7248 42100
rect 7012 42084 7064 42090
rect 7012 42026 7064 42032
rect 6920 41268 6972 41274
rect 6920 41210 6972 41216
rect 6656 40594 6684 41006
rect 6840 40990 6960 41018
rect 6828 40928 6880 40934
rect 6828 40870 6880 40876
rect 6840 40662 6868 40870
rect 6828 40656 6880 40662
rect 6828 40598 6880 40604
rect 6644 40588 6696 40594
rect 6644 40530 6696 40536
rect 6656 40186 6684 40530
rect 6932 40361 6960 40990
rect 6918 40352 6974 40361
rect 6918 40287 6974 40296
rect 6644 40180 6696 40186
rect 6644 40122 6696 40128
rect 6734 40080 6790 40089
rect 6734 40015 6790 40024
rect 6644 39296 6696 39302
rect 6644 39238 6696 39244
rect 6550 38992 6606 39001
rect 6550 38927 6606 38936
rect 6656 38876 6684 39238
rect 6564 38848 6684 38876
rect 6460 38480 6512 38486
rect 6460 38422 6512 38428
rect 6288 37726 6408 37754
rect 6276 36576 6328 36582
rect 6276 36518 6328 36524
rect 6288 36378 6316 36518
rect 6276 36372 6328 36378
rect 6276 36314 6328 36320
rect 6380 36258 6408 37726
rect 6472 37330 6500 38422
rect 6564 37330 6592 38848
rect 6644 37800 6696 37806
rect 6644 37742 6696 37748
rect 6460 37324 6512 37330
rect 6460 37266 6512 37272
rect 6552 37324 6604 37330
rect 6552 37266 6604 37272
rect 6288 36230 6408 36258
rect 6184 35760 6236 35766
rect 6184 35702 6236 35708
rect 6196 35630 6224 35702
rect 6184 35624 6236 35630
rect 6184 35566 6236 35572
rect 6184 35488 6236 35494
rect 6182 35456 6184 35465
rect 6236 35456 6238 35465
rect 6182 35391 6238 35400
rect 6104 35278 6224 35306
rect 5998 35255 6000 35264
rect 6052 35255 6054 35264
rect 6000 35226 6052 35232
rect 5816 35148 5868 35154
rect 5816 35090 5868 35096
rect 5998 34776 6054 34785
rect 5816 34740 5868 34746
rect 5998 34711 6054 34720
rect 5816 34682 5868 34688
rect 5828 33658 5856 34682
rect 6012 34678 6040 34711
rect 6000 34672 6052 34678
rect 6000 34614 6052 34620
rect 5908 34604 5960 34610
rect 5908 34546 5960 34552
rect 5816 33652 5868 33658
rect 5816 33594 5868 33600
rect 5816 32972 5868 32978
rect 5816 32914 5868 32920
rect 5828 32201 5856 32914
rect 5920 32230 5948 34546
rect 6012 33522 6040 34614
rect 6092 34400 6144 34406
rect 6092 34342 6144 34348
rect 6104 34066 6132 34342
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6090 33824 6146 33833
rect 6090 33759 6146 33768
rect 6000 33516 6052 33522
rect 6000 33458 6052 33464
rect 6104 33402 6132 33759
rect 6012 33374 6132 33402
rect 5908 32224 5960 32230
rect 5814 32192 5870 32201
rect 5908 32166 5960 32172
rect 5814 32127 5870 32136
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 5814 31784 5870 31793
rect 5920 31770 5948 31962
rect 6012 31890 6040 33374
rect 6196 32978 6224 35278
rect 6288 35222 6316 36230
rect 6472 36174 6500 37266
rect 6564 36786 6592 37266
rect 6552 36780 6604 36786
rect 6552 36722 6604 36728
rect 6656 36378 6684 37742
rect 6748 37210 6776 40015
rect 7024 39982 7052 42026
rect 7196 41608 7248 41614
rect 7196 41550 7248 41556
rect 7208 41478 7236 41550
rect 7104 41472 7156 41478
rect 7104 41414 7156 41420
rect 7196 41472 7248 41478
rect 7196 41414 7248 41420
rect 7116 40662 7144 41414
rect 7196 41064 7248 41070
rect 7196 41006 7248 41012
rect 7104 40656 7156 40662
rect 7104 40598 7156 40604
rect 7012 39976 7064 39982
rect 7012 39918 7064 39924
rect 7208 39846 7236 41006
rect 7300 40474 7328 42638
rect 7470 42599 7526 42608
rect 7760 42537 7788 42774
rect 8128 42770 8524 42786
rect 8680 42770 8708 43114
rect 9956 43104 10008 43110
rect 9956 43046 10008 43052
rect 9036 42832 9088 42838
rect 9036 42774 9088 42780
rect 7932 42764 7984 42770
rect 7932 42706 7984 42712
rect 8024 42764 8076 42770
rect 8128 42764 8536 42770
rect 8128 42758 8484 42764
rect 8024 42706 8076 42712
rect 8484 42706 8536 42712
rect 8668 42764 8720 42770
rect 8668 42706 8720 42712
rect 7746 42528 7802 42537
rect 7746 42463 7802 42472
rect 7944 42378 7972 42706
rect 7668 42350 7972 42378
rect 7472 42152 7524 42158
rect 7472 42094 7524 42100
rect 7380 41744 7432 41750
rect 7380 41686 7432 41692
rect 7392 41585 7420 41686
rect 7378 41576 7434 41585
rect 7378 41511 7434 41520
rect 7378 41304 7434 41313
rect 7378 41239 7434 41248
rect 7392 41070 7420 41239
rect 7484 41070 7512 42094
rect 7564 42016 7616 42022
rect 7564 41958 7616 41964
rect 7576 41154 7604 41958
rect 7668 41449 7696 42350
rect 7840 42288 7892 42294
rect 7840 42230 7892 42236
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 7654 41440 7710 41449
rect 7654 41375 7710 41384
rect 7760 41206 7788 42094
rect 7748 41200 7800 41206
rect 7576 41126 7696 41154
rect 7748 41142 7800 41148
rect 7852 41138 7880 42230
rect 7932 42152 7984 42158
rect 7932 42094 7984 42100
rect 7380 41064 7432 41070
rect 7380 41006 7432 41012
rect 7472 41064 7524 41070
rect 7668 41052 7696 41126
rect 7840 41132 7892 41138
rect 7840 41074 7892 41080
rect 7668 41024 7788 41052
rect 7472 41006 7524 41012
rect 7380 40928 7432 40934
rect 7380 40870 7432 40876
rect 7392 40594 7420 40870
rect 7656 40656 7708 40662
rect 7576 40616 7656 40644
rect 7380 40588 7432 40594
rect 7380 40530 7432 40536
rect 7472 40520 7524 40526
rect 7470 40488 7472 40497
rect 7524 40488 7526 40497
rect 7300 40446 7420 40474
rect 7288 40384 7340 40390
rect 7288 40326 7340 40332
rect 7300 40050 7328 40326
rect 7392 40118 7420 40446
rect 7470 40423 7526 40432
rect 7472 40384 7524 40390
rect 7472 40326 7524 40332
rect 7380 40112 7432 40118
rect 7380 40054 7432 40060
rect 7288 40044 7340 40050
rect 7288 39986 7340 39992
rect 7484 39982 7512 40326
rect 7576 39982 7604 40616
rect 7656 40598 7708 40604
rect 7656 40452 7708 40458
rect 7656 40394 7708 40400
rect 7668 40186 7696 40394
rect 7656 40180 7708 40186
rect 7656 40122 7708 40128
rect 7472 39976 7524 39982
rect 7472 39918 7524 39924
rect 7564 39976 7616 39982
rect 7564 39918 7616 39924
rect 7760 39846 7788 41024
rect 7852 40089 7880 41074
rect 7944 41070 7972 42094
rect 8036 42090 8064 42706
rect 8116 42696 8168 42702
rect 8300 42696 8352 42702
rect 8116 42638 8168 42644
rect 8298 42664 8300 42673
rect 8352 42664 8354 42673
rect 8128 42158 8156 42638
rect 8298 42599 8354 42608
rect 8208 42560 8260 42566
rect 8208 42502 8260 42508
rect 8392 42560 8444 42566
rect 8392 42502 8444 42508
rect 8116 42152 8168 42158
rect 8116 42094 8168 42100
rect 8024 42084 8076 42090
rect 8024 42026 8076 42032
rect 8116 42016 8168 42022
rect 8116 41958 8168 41964
rect 8128 41682 8156 41958
rect 8116 41676 8168 41682
rect 8116 41618 8168 41624
rect 8024 41200 8076 41206
rect 8024 41142 8076 41148
rect 7932 41064 7984 41070
rect 7932 41006 7984 41012
rect 8036 40662 8064 41142
rect 8116 41132 8168 41138
rect 8116 41074 8168 41080
rect 8024 40656 8076 40662
rect 8024 40598 8076 40604
rect 7932 40384 7984 40390
rect 7984 40332 8064 40338
rect 7932 40326 8064 40332
rect 7944 40310 8064 40326
rect 7838 40080 7894 40089
rect 7838 40015 7894 40024
rect 7196 39840 7248 39846
rect 7656 39840 7708 39846
rect 7196 39782 7248 39788
rect 7286 39808 7342 39817
rect 7656 39782 7708 39788
rect 7748 39840 7800 39846
rect 7748 39782 7800 39788
rect 7286 39743 7342 39752
rect 7196 39296 7248 39302
rect 7196 39238 7248 39244
rect 7208 39030 7236 39238
rect 7196 39024 7248 39030
rect 7196 38966 7248 38972
rect 7102 38856 7158 38865
rect 7300 38842 7328 39743
rect 7668 39545 7696 39782
rect 7378 39536 7434 39545
rect 7378 39471 7434 39480
rect 7654 39536 7710 39545
rect 7760 39506 7972 39522
rect 7654 39471 7710 39480
rect 7748 39500 7972 39506
rect 7392 39030 7420 39471
rect 7800 39494 7972 39500
rect 7748 39442 7800 39448
rect 7564 39432 7616 39438
rect 7564 39374 7616 39380
rect 7380 39024 7432 39030
rect 7380 38966 7432 38972
rect 7470 38992 7526 39001
rect 7470 38927 7526 38936
rect 7158 38814 7328 38842
rect 7102 38791 7158 38800
rect 7196 38752 7248 38758
rect 7196 38694 7248 38700
rect 6840 38406 7144 38434
rect 6840 38010 6868 38406
rect 7116 38350 7144 38406
rect 7104 38344 7156 38350
rect 7104 38286 7156 38292
rect 7104 38208 7156 38214
rect 7104 38150 7156 38156
rect 7116 38010 7144 38150
rect 7208 38049 7236 38694
rect 7194 38040 7250 38049
rect 6828 38004 6880 38010
rect 6828 37946 6880 37952
rect 7104 38004 7156 38010
rect 7194 37975 7250 37984
rect 7104 37946 7156 37952
rect 6840 37398 6868 37946
rect 6920 37800 6972 37806
rect 6920 37742 6972 37748
rect 7010 37768 7066 37777
rect 6828 37392 6880 37398
rect 6828 37334 6880 37340
rect 6932 37330 6960 37742
rect 7010 37703 7066 37712
rect 7104 37732 7156 37738
rect 6920 37324 6972 37330
rect 6920 37266 6972 37272
rect 6748 37182 6868 37210
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 6748 36582 6776 36790
rect 6736 36576 6788 36582
rect 6736 36518 6788 36524
rect 6644 36372 6696 36378
rect 6644 36314 6696 36320
rect 6736 36304 6788 36310
rect 6736 36246 6788 36252
rect 6552 36236 6604 36242
rect 6552 36178 6604 36184
rect 6644 36236 6696 36242
rect 6644 36178 6696 36184
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 6460 36168 6512 36174
rect 6460 36110 6512 36116
rect 6380 35834 6408 36110
rect 6460 36032 6512 36038
rect 6460 35974 6512 35980
rect 6472 35873 6500 35974
rect 6458 35864 6514 35873
rect 6368 35828 6420 35834
rect 6458 35799 6514 35808
rect 6368 35770 6420 35776
rect 6460 35624 6512 35630
rect 6460 35566 6512 35572
rect 6472 35290 6500 35566
rect 6460 35284 6512 35290
rect 6460 35226 6512 35232
rect 6564 35222 6592 36178
rect 6656 35714 6684 36178
rect 6748 35834 6776 36246
rect 6736 35828 6788 35834
rect 6736 35770 6788 35776
rect 6656 35686 6776 35714
rect 6644 35624 6696 35630
rect 6644 35566 6696 35572
rect 6276 35216 6328 35222
rect 6276 35158 6328 35164
rect 6552 35216 6604 35222
rect 6552 35158 6604 35164
rect 6656 35170 6684 35566
rect 6748 35290 6776 35686
rect 6736 35284 6788 35290
rect 6736 35226 6788 35232
rect 6656 35142 6776 35170
rect 6552 35080 6604 35086
rect 6552 35022 6604 35028
rect 6368 34944 6420 34950
rect 6368 34886 6420 34892
rect 6380 34649 6408 34886
rect 6366 34640 6422 34649
rect 6366 34575 6422 34584
rect 6380 34542 6408 34575
rect 6368 34536 6420 34542
rect 6288 34496 6368 34524
rect 6288 34202 6316 34496
rect 6368 34478 6420 34484
rect 6460 34536 6512 34542
rect 6460 34478 6512 34484
rect 6368 34400 6420 34406
rect 6368 34342 6420 34348
rect 6276 34196 6328 34202
rect 6276 34138 6328 34144
rect 6288 33522 6316 34138
rect 6380 33697 6408 34342
rect 6366 33688 6422 33697
rect 6366 33623 6422 33632
rect 6276 33516 6328 33522
rect 6276 33458 6328 33464
rect 6184 32972 6236 32978
rect 6184 32914 6236 32920
rect 6092 32768 6144 32774
rect 6092 32710 6144 32716
rect 6104 32570 6132 32710
rect 6092 32564 6144 32570
rect 6092 32506 6144 32512
rect 6104 31958 6132 32506
rect 6196 32434 6224 32914
rect 6288 32502 6316 33458
rect 6368 33448 6420 33454
rect 6366 33416 6368 33425
rect 6420 33416 6422 33425
rect 6366 33351 6422 33360
rect 6472 33114 6500 34478
rect 6460 33108 6512 33114
rect 6460 33050 6512 33056
rect 6460 32972 6512 32978
rect 6460 32914 6512 32920
rect 6276 32496 6328 32502
rect 6276 32438 6328 32444
rect 6472 32434 6500 32914
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 6276 32360 6328 32366
rect 6276 32302 6328 32308
rect 6366 32328 6422 32337
rect 6184 32292 6236 32298
rect 6184 32234 6236 32240
rect 6092 31952 6144 31958
rect 6092 31894 6144 31900
rect 6000 31884 6052 31890
rect 6000 31826 6052 31832
rect 5920 31742 6040 31770
rect 5814 31719 5870 31728
rect 5828 31482 5856 31719
rect 5908 31680 5960 31686
rect 5908 31622 5960 31628
rect 5816 31476 5868 31482
rect 5816 31418 5868 31424
rect 5814 31376 5870 31385
rect 5814 31311 5816 31320
rect 5868 31311 5870 31320
rect 5816 31282 5868 31288
rect 5814 31240 5870 31249
rect 5814 31175 5816 31184
rect 5868 31175 5870 31184
rect 5816 31146 5868 31152
rect 5814 30968 5870 30977
rect 5814 30903 5870 30912
rect 5722 30696 5778 30705
rect 5722 30631 5778 30640
rect 5724 30592 5776 30598
rect 5724 30534 5776 30540
rect 5736 30433 5764 30534
rect 5722 30424 5778 30433
rect 5632 30388 5684 30394
rect 5722 30359 5778 30368
rect 5632 30330 5684 30336
rect 5828 30326 5856 30903
rect 5816 30320 5868 30326
rect 5538 30288 5594 30297
rect 5920 30297 5948 31622
rect 6012 31346 6040 31742
rect 6000 31340 6052 31346
rect 6052 31300 6132 31328
rect 6000 31282 6052 31288
rect 6000 30660 6052 30666
rect 6000 30602 6052 30608
rect 6012 30394 6040 30602
rect 6000 30388 6052 30394
rect 6000 30330 6052 30336
rect 5816 30262 5868 30268
rect 5906 30288 5962 30297
rect 5538 30223 5594 30232
rect 5962 30246 6040 30274
rect 5906 30223 5962 30232
rect 5552 30190 5580 30223
rect 5540 30184 5592 30190
rect 5724 30184 5776 30190
rect 5540 30126 5592 30132
rect 5644 30144 5724 30172
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5448 29844 5500 29850
rect 5448 29786 5500 29792
rect 5356 29708 5408 29714
rect 5408 29668 5488 29696
rect 5356 29650 5408 29656
rect 5264 29572 5316 29578
rect 5264 29514 5316 29520
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5170 28792 5226 28801
rect 5170 28727 5226 28736
rect 5184 28694 5212 28727
rect 5172 28688 5224 28694
rect 5224 28648 5304 28676
rect 5172 28630 5224 28636
rect 5172 28008 5224 28014
rect 5172 27950 5224 27956
rect 5184 27538 5212 27950
rect 5276 27946 5304 28648
rect 5264 27940 5316 27946
rect 5264 27882 5316 27888
rect 5276 27674 5304 27882
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 5368 27538 5396 29446
rect 5460 29034 5488 29668
rect 5552 29238 5580 29990
rect 5644 29510 5672 30144
rect 5724 30126 5776 30132
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 5632 29504 5684 29510
rect 5632 29446 5684 29452
rect 5540 29232 5592 29238
rect 5540 29174 5592 29180
rect 5632 29164 5684 29170
rect 5632 29106 5684 29112
rect 5448 29028 5500 29034
rect 5448 28970 5500 28976
rect 5080 27532 5132 27538
rect 5080 27474 5132 27480
rect 5172 27532 5224 27538
rect 5172 27474 5224 27480
rect 5356 27532 5408 27538
rect 5356 27474 5408 27480
rect 5460 27402 5488 28970
rect 5644 28966 5672 29106
rect 5736 29102 5764 29786
rect 5814 29744 5870 29753
rect 5814 29679 5816 29688
rect 5868 29679 5870 29688
rect 5908 29708 5960 29714
rect 5816 29650 5868 29656
rect 5908 29650 5960 29656
rect 5724 29096 5776 29102
rect 5724 29038 5776 29044
rect 5632 28960 5684 28966
rect 5632 28902 5684 28908
rect 5724 28960 5776 28966
rect 5724 28902 5776 28908
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5552 28014 5580 28698
rect 5736 28694 5764 28902
rect 5724 28688 5776 28694
rect 5724 28630 5776 28636
rect 5828 28626 5856 29650
rect 5920 28762 5948 29650
rect 6012 29170 6040 30246
rect 6104 29850 6132 31300
rect 6092 29844 6144 29850
rect 6092 29786 6144 29792
rect 6196 29730 6224 32234
rect 6288 32201 6316 32302
rect 6564 32314 6592 35022
rect 6748 35018 6776 35142
rect 6644 35012 6696 35018
rect 6644 34954 6696 34960
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6656 34377 6684 34954
rect 6736 34468 6788 34474
rect 6736 34410 6788 34416
rect 6642 34368 6698 34377
rect 6642 34303 6698 34312
rect 6644 34196 6696 34202
rect 6644 34138 6696 34144
rect 6656 33590 6684 34138
rect 6644 33584 6696 33590
rect 6644 33526 6696 33532
rect 6644 33448 6696 33454
rect 6642 33416 6644 33425
rect 6696 33416 6698 33425
rect 6642 33351 6698 33360
rect 6748 33153 6776 34410
rect 6840 33289 6868 37182
rect 7024 36718 7052 37703
rect 7104 37674 7156 37680
rect 7196 37732 7248 37738
rect 7196 37674 7248 37680
rect 7116 36854 7144 37674
rect 7208 37466 7236 37674
rect 7196 37460 7248 37466
rect 7196 37402 7248 37408
rect 7300 37194 7328 38814
rect 7380 38752 7432 38758
rect 7380 38694 7432 38700
rect 7288 37188 7340 37194
rect 7288 37130 7340 37136
rect 7104 36848 7156 36854
rect 7156 36808 7236 36836
rect 7104 36790 7156 36796
rect 7012 36712 7064 36718
rect 7012 36654 7064 36660
rect 6918 36408 6974 36417
rect 6918 36343 6974 36352
rect 6932 36156 6960 36343
rect 7024 36310 7052 36654
rect 7104 36644 7156 36650
rect 7104 36586 7156 36592
rect 7012 36304 7064 36310
rect 7012 36246 7064 36252
rect 7012 36168 7064 36174
rect 6932 36128 7012 36156
rect 7012 36110 7064 36116
rect 7116 35834 7144 36586
rect 7104 35828 7156 35834
rect 7104 35770 7156 35776
rect 7208 35714 7236 36808
rect 7288 36712 7340 36718
rect 7286 36680 7288 36689
rect 7340 36680 7342 36689
rect 7286 36615 7342 36624
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7300 36417 7328 36518
rect 7286 36408 7342 36417
rect 7286 36343 7342 36352
rect 7392 36242 7420 38694
rect 7484 36961 7512 38927
rect 7576 38826 7604 39374
rect 7760 39302 7788 39442
rect 7840 39432 7892 39438
rect 7840 39374 7892 39380
rect 7748 39296 7800 39302
rect 7748 39238 7800 39244
rect 7656 38956 7708 38962
rect 7656 38898 7708 38904
rect 7564 38820 7616 38826
rect 7564 38762 7616 38768
rect 7470 36952 7526 36961
rect 7470 36887 7526 36896
rect 7472 36712 7524 36718
rect 7472 36654 7524 36660
rect 7380 36236 7432 36242
rect 7300 36196 7380 36224
rect 7300 35766 7328 36196
rect 7380 36178 7432 36184
rect 7380 36032 7432 36038
rect 7484 36009 7512 36654
rect 7576 36122 7604 38762
rect 7668 38758 7696 38898
rect 7748 38888 7800 38894
rect 7748 38830 7800 38836
rect 7760 38758 7788 38830
rect 7656 38752 7708 38758
rect 7656 38694 7708 38700
rect 7748 38752 7800 38758
rect 7748 38694 7800 38700
rect 7852 38350 7880 39374
rect 7944 38418 7972 39494
rect 8036 38894 8064 40310
rect 8128 39273 8156 41074
rect 8220 40662 8248 42502
rect 8404 42362 8432 42502
rect 8392 42356 8444 42362
rect 8392 42298 8444 42304
rect 8392 42152 8444 42158
rect 8392 42094 8444 42100
rect 8760 42152 8812 42158
rect 8760 42094 8812 42100
rect 8404 41002 8432 42094
rect 8484 42016 8536 42022
rect 8484 41958 8536 41964
rect 8496 41750 8524 41958
rect 8484 41744 8536 41750
rect 8484 41686 8536 41692
rect 8668 41676 8720 41682
rect 8668 41618 8720 41624
rect 8680 41478 8708 41618
rect 8668 41472 8720 41478
rect 8668 41414 8720 41420
rect 8772 41313 8800 42094
rect 8852 42084 8904 42090
rect 8852 42026 8904 42032
rect 8944 42084 8996 42090
rect 8944 42026 8996 42032
rect 8758 41304 8814 41313
rect 8758 41239 8814 41248
rect 8864 41002 8892 42026
rect 8956 41070 8984 42026
rect 9048 41546 9076 42774
rect 9680 42696 9732 42702
rect 9680 42638 9732 42644
rect 9772 42696 9824 42702
rect 9772 42638 9824 42644
rect 9404 42628 9456 42634
rect 9404 42570 9456 42576
rect 9128 42560 9180 42566
rect 9128 42502 9180 42508
rect 9140 42362 9168 42502
rect 9128 42356 9180 42362
rect 9128 42298 9180 42304
rect 9140 41993 9168 42298
rect 9220 42152 9272 42158
rect 9220 42094 9272 42100
rect 9126 41984 9182 41993
rect 9126 41919 9182 41928
rect 9232 41818 9260 42094
rect 9220 41812 9272 41818
rect 9220 41754 9272 41760
rect 9036 41540 9088 41546
rect 9036 41482 9088 41488
rect 9416 41478 9444 42570
rect 9404 41472 9456 41478
rect 9404 41414 9456 41420
rect 8944 41064 8996 41070
rect 8944 41006 8996 41012
rect 9312 41064 9364 41070
rect 9312 41006 9364 41012
rect 8392 40996 8444 41002
rect 8392 40938 8444 40944
rect 8852 40996 8904 41002
rect 8852 40938 8904 40944
rect 8300 40928 8352 40934
rect 8300 40870 8352 40876
rect 8208 40656 8260 40662
rect 8208 40598 8260 40604
rect 8206 40352 8262 40361
rect 8206 40287 8262 40296
rect 8220 40186 8248 40287
rect 8208 40180 8260 40186
rect 8208 40122 8260 40128
rect 8220 39302 8248 40122
rect 8208 39296 8260 39302
rect 8114 39264 8170 39273
rect 8208 39238 8260 39244
rect 8114 39199 8170 39208
rect 8220 39001 8248 39238
rect 8312 39030 8340 40870
rect 8404 40633 8432 40938
rect 8484 40928 8536 40934
rect 8484 40870 8536 40876
rect 8390 40624 8446 40633
rect 8390 40559 8446 40568
rect 8392 40452 8444 40458
rect 8392 40394 8444 40400
rect 8300 39024 8352 39030
rect 8206 38992 8262 39001
rect 8300 38966 8352 38972
rect 8206 38927 8262 38936
rect 8024 38888 8076 38894
rect 8024 38830 8076 38836
rect 8024 38752 8076 38758
rect 8024 38694 8076 38700
rect 7932 38412 7984 38418
rect 7932 38354 7984 38360
rect 7840 38344 7892 38350
rect 7840 38286 7892 38292
rect 7748 38276 7800 38282
rect 7748 38218 7800 38224
rect 7656 38208 7708 38214
rect 7656 38150 7708 38156
rect 7668 37398 7696 38150
rect 7656 37392 7708 37398
rect 7656 37334 7708 37340
rect 7656 37188 7708 37194
rect 7656 37130 7708 37136
rect 7668 36922 7696 37130
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 7760 36718 7788 38218
rect 7840 37664 7892 37670
rect 7840 37606 7892 37612
rect 7852 37466 7880 37606
rect 7840 37460 7892 37466
rect 7840 37402 7892 37408
rect 7748 36712 7800 36718
rect 7748 36654 7800 36660
rect 7840 36712 7892 36718
rect 7840 36654 7892 36660
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 7748 36576 7800 36582
rect 7852 36553 7880 36654
rect 7748 36518 7800 36524
rect 7838 36544 7894 36553
rect 7668 36281 7696 36518
rect 7654 36272 7710 36281
rect 7654 36207 7710 36216
rect 7760 36224 7788 36518
rect 7838 36479 7894 36488
rect 7840 36236 7892 36242
rect 7760 36196 7840 36224
rect 7840 36178 7892 36184
rect 7944 36174 7972 38354
rect 8036 37641 8064 38694
rect 8300 38344 8352 38350
rect 8300 38286 8352 38292
rect 8208 37800 8260 37806
rect 8208 37742 8260 37748
rect 8022 37632 8078 37641
rect 8022 37567 8078 37576
rect 8116 37256 8168 37262
rect 8116 37198 8168 37204
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 8036 36310 8064 37062
rect 8128 36961 8156 37198
rect 8114 36952 8170 36961
rect 8114 36887 8170 36896
rect 8114 36816 8170 36825
rect 8114 36751 8170 36760
rect 8024 36304 8076 36310
rect 8024 36246 8076 36252
rect 7932 36168 7984 36174
rect 7576 36094 7696 36122
rect 7932 36110 7984 36116
rect 7380 35974 7432 35980
rect 7470 36000 7526 36009
rect 7024 35686 7236 35714
rect 7288 35760 7340 35766
rect 7288 35702 7340 35708
rect 6920 35148 6972 35154
rect 6920 35090 6972 35096
rect 6932 34950 6960 35090
rect 6920 34944 6972 34950
rect 6920 34886 6972 34892
rect 6920 34468 6972 34474
rect 6920 34410 6972 34416
rect 6826 33280 6882 33289
rect 6826 33215 6882 33224
rect 6734 33144 6790 33153
rect 6734 33079 6790 33088
rect 6932 32978 6960 34410
rect 7024 34406 7052 35686
rect 7196 35624 7248 35630
rect 7196 35566 7248 35572
rect 7286 35592 7342 35601
rect 7104 35148 7156 35154
rect 7104 35090 7156 35096
rect 7116 34746 7144 35090
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 7012 34400 7064 34406
rect 7012 34342 7064 34348
rect 7104 33516 7156 33522
rect 7104 33458 7156 33464
rect 7116 33114 7144 33458
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 7104 33108 7156 33114
rect 7104 33050 7156 33056
rect 6644 32972 6696 32978
rect 6644 32914 6696 32920
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 6656 32570 6684 32914
rect 6736 32768 6788 32774
rect 6734 32736 6736 32745
rect 6788 32736 6790 32745
rect 6734 32671 6790 32680
rect 6734 32600 6790 32609
rect 6644 32564 6696 32570
rect 6840 32570 6868 32914
rect 6920 32836 6972 32842
rect 6920 32778 6972 32784
rect 6734 32535 6790 32544
rect 6828 32564 6880 32570
rect 6644 32506 6696 32512
rect 6366 32263 6422 32272
rect 6472 32286 6592 32314
rect 6274 32192 6330 32201
rect 6274 32127 6330 32136
rect 6288 31890 6316 32127
rect 6380 31958 6408 32263
rect 6368 31952 6420 31958
rect 6368 31894 6420 31900
rect 6276 31884 6328 31890
rect 6276 31826 6328 31832
rect 6288 30190 6316 31826
rect 6472 31822 6500 32286
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6368 31816 6420 31822
rect 6368 31758 6420 31764
rect 6460 31816 6512 31822
rect 6460 31758 6512 31764
rect 6380 31521 6408 31758
rect 6366 31512 6422 31521
rect 6366 31447 6422 31456
rect 6564 31396 6592 32166
rect 6748 32042 6776 32535
rect 6828 32506 6880 32512
rect 6828 32360 6880 32366
rect 6826 32328 6828 32337
rect 6880 32328 6882 32337
rect 6826 32263 6882 32272
rect 6656 32026 6776 32042
rect 6644 32020 6776 32026
rect 6696 32014 6776 32020
rect 6644 31962 6696 31968
rect 6736 31952 6788 31958
rect 6736 31894 6788 31900
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6656 31793 6684 31826
rect 6642 31784 6698 31793
rect 6642 31719 6698 31728
rect 6380 31368 6592 31396
rect 6380 30802 6408 31368
rect 6748 31278 6776 31894
rect 6826 31648 6882 31657
rect 6826 31583 6882 31592
rect 6460 31272 6512 31278
rect 6460 31214 6512 31220
rect 6552 31272 6604 31278
rect 6736 31272 6788 31278
rect 6552 31214 6604 31220
rect 6642 31240 6698 31249
rect 6472 30938 6500 31214
rect 6460 30932 6512 30938
rect 6460 30874 6512 30880
rect 6368 30796 6420 30802
rect 6368 30738 6420 30744
rect 6460 30796 6512 30802
rect 6460 30738 6512 30744
rect 6276 30184 6328 30190
rect 6276 30126 6328 30132
rect 6288 30025 6316 30126
rect 6274 30016 6330 30025
rect 6274 29951 6330 29960
rect 6380 29753 6408 30738
rect 6104 29714 6224 29730
rect 6092 29708 6224 29714
rect 6144 29702 6224 29708
rect 6366 29744 6422 29753
rect 6366 29679 6422 29688
rect 6092 29650 6144 29656
rect 6184 29651 6236 29657
rect 6184 29593 6236 29599
rect 6092 29504 6144 29510
rect 6092 29446 6144 29452
rect 6000 29164 6052 29170
rect 6000 29106 6052 29112
rect 5908 28756 5960 28762
rect 5908 28698 5960 28704
rect 6012 28626 6040 29106
rect 5816 28620 5868 28626
rect 5816 28562 5868 28568
rect 6000 28620 6052 28626
rect 6000 28562 6052 28568
rect 5828 28014 5856 28562
rect 5908 28416 5960 28422
rect 5908 28358 5960 28364
rect 5540 28008 5592 28014
rect 5540 27950 5592 27956
rect 5816 28008 5868 28014
rect 5816 27950 5868 27956
rect 5920 27962 5948 28358
rect 5920 27934 6040 27962
rect 5816 27872 5868 27878
rect 5816 27814 5868 27820
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5172 27328 5224 27334
rect 5172 27270 5224 27276
rect 4988 27056 5040 27062
rect 4988 26998 5040 27004
rect 5080 26240 5132 26246
rect 5184 26228 5212 27270
rect 5632 26988 5684 26994
rect 5632 26930 5684 26936
rect 5356 26784 5408 26790
rect 5356 26726 5408 26732
rect 5368 26450 5396 26726
rect 5356 26444 5408 26450
rect 5356 26386 5408 26392
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 5540 26376 5592 26382
rect 5540 26318 5592 26324
rect 5184 26200 5304 26228
rect 5080 26182 5132 26188
rect 4988 26036 5040 26042
rect 4988 25978 5040 25984
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4896 23792 4948 23798
rect 4896 23734 4948 23740
rect 4804 23724 4856 23730
rect 4804 23666 4856 23672
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4710 21720 4766 21729
rect 4710 21655 4766 21664
rect 4710 21584 4766 21593
rect 4710 21519 4766 21528
rect 4252 21480 4304 21486
rect 4250 21448 4252 21457
rect 4344 21480 4396 21486
rect 4304 21448 4306 21457
rect 4344 21422 4396 21428
rect 4250 21383 4306 21392
rect 4356 21332 4384 21422
rect 4264 21304 4384 21332
rect 4264 21128 4292 21304
rect 4322 21244 4630 21253
rect 4322 21242 4328 21244
rect 4384 21242 4408 21244
rect 4464 21242 4488 21244
rect 4544 21242 4568 21244
rect 4624 21242 4630 21244
rect 4384 21190 4386 21242
rect 4566 21190 4568 21242
rect 4322 21188 4328 21190
rect 4384 21188 4408 21190
rect 4464 21188 4488 21190
rect 4544 21188 4568 21190
rect 4624 21188 4630 21190
rect 4322 21179 4630 21188
rect 4264 21100 4568 21128
rect 4250 21040 4306 21049
rect 4250 20975 4252 20984
rect 4304 20975 4306 20984
rect 4434 21040 4490 21049
rect 4434 20975 4490 20984
rect 4252 20946 4304 20952
rect 4264 20806 4292 20946
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 4264 20398 4292 20742
rect 4252 20392 4304 20398
rect 4252 20334 4304 20340
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3988 20058 4016 20198
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4080 19922 4108 20318
rect 4160 20324 4212 20330
rect 4160 20266 4212 20272
rect 4448 20244 4476 20975
rect 4540 20942 4568 21100
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 4528 20936 4580 20942
rect 4528 20878 4580 20884
rect 4540 20398 4568 20878
rect 4632 20602 4660 20946
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4724 20448 4752 21519
rect 4632 20420 4752 20448
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4632 20262 4660 20420
rect 4710 20360 4766 20369
rect 4710 20295 4766 20304
rect 4816 20312 4844 23462
rect 4908 23118 4936 23734
rect 5000 23594 5028 25978
rect 5092 25430 5120 26182
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5080 25424 5132 25430
rect 5080 25366 5132 25372
rect 5080 25288 5132 25294
rect 5080 25230 5132 25236
rect 5092 24682 5120 25230
rect 5080 24676 5132 24682
rect 5080 24618 5132 24624
rect 5092 24410 5120 24618
rect 5080 24404 5132 24410
rect 5080 24346 5132 24352
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 4896 23112 4948 23118
rect 4896 23054 4948 23060
rect 4894 22944 4950 22953
rect 4894 22879 4950 22888
rect 4908 22098 4936 22879
rect 5000 22710 5028 23530
rect 5092 23322 5120 23802
rect 5080 23316 5132 23322
rect 5080 23258 5132 23264
rect 5080 23180 5132 23186
rect 5080 23122 5132 23128
rect 5092 22817 5120 23122
rect 5078 22808 5134 22817
rect 5078 22743 5134 22752
rect 4988 22704 5040 22710
rect 5184 22692 5212 25638
rect 5276 25129 5304 26200
rect 5460 25702 5488 26318
rect 5552 25906 5580 26318
rect 5644 26042 5672 26930
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5630 25800 5686 25809
rect 5540 25764 5592 25770
rect 5630 25735 5686 25744
rect 5540 25706 5592 25712
rect 5448 25696 5500 25702
rect 5448 25638 5500 25644
rect 5552 25294 5580 25706
rect 5540 25288 5592 25294
rect 5540 25230 5592 25236
rect 5262 25120 5318 25129
rect 5262 25055 5318 25064
rect 5264 24744 5316 24750
rect 5264 24686 5316 24692
rect 4988 22646 5040 22652
rect 5092 22664 5212 22692
rect 4988 22432 5040 22438
rect 4988 22374 5040 22380
rect 5000 22273 5028 22374
rect 4986 22264 5042 22273
rect 4986 22199 5042 22208
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4986 21992 5042 22001
rect 4986 21927 5042 21936
rect 4896 21888 4948 21894
rect 4894 21856 4896 21865
rect 4948 21856 4950 21865
rect 4894 21791 4950 21800
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4908 21146 4936 21422
rect 5000 21146 5028 21927
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4988 21140 5040 21146
rect 4988 21082 5040 21088
rect 4908 21010 4936 21082
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 4264 20216 4476 20244
rect 4620 20256 4672 20262
rect 4158 20088 4214 20097
rect 4158 20023 4160 20032
rect 4212 20023 4214 20032
rect 4160 19994 4212 20000
rect 4172 19922 4200 19994
rect 3884 19916 3936 19922
rect 4068 19916 4120 19922
rect 3936 19876 4016 19904
rect 3884 19858 3936 19864
rect 3988 19786 4016 19876
rect 4068 19858 4120 19864
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 3976 19780 4028 19786
rect 3976 19722 4028 19728
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 3662 19612 3970 19621
rect 3662 19610 3668 19612
rect 3724 19610 3748 19612
rect 3804 19610 3828 19612
rect 3884 19610 3908 19612
rect 3964 19610 3970 19612
rect 3724 19558 3726 19610
rect 3906 19558 3908 19610
rect 3662 19556 3668 19558
rect 3724 19556 3748 19558
rect 3804 19556 3828 19558
rect 3884 19556 3908 19558
rect 3964 19556 3970 19558
rect 3662 19547 3970 19556
rect 3528 19468 3648 19496
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 3422 19136 3478 19145
rect 3422 19071 3478 19080
rect 3528 18902 3556 19178
rect 3620 19009 3648 19468
rect 4172 19428 4200 19654
rect 4264 19530 4292 20216
rect 4620 20198 4672 20204
rect 4322 20156 4630 20165
rect 4322 20154 4328 20156
rect 4384 20154 4408 20156
rect 4464 20154 4488 20156
rect 4544 20154 4568 20156
rect 4624 20154 4630 20156
rect 4384 20102 4386 20154
rect 4566 20102 4568 20154
rect 4322 20100 4328 20102
rect 4384 20100 4408 20102
rect 4464 20100 4488 20102
rect 4544 20100 4568 20102
rect 4624 20100 4630 20102
rect 4322 20091 4630 20100
rect 4436 19916 4488 19922
rect 4436 19858 4488 19864
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4342 19544 4398 19553
rect 4264 19502 4342 19530
rect 4448 19514 4476 19858
rect 4540 19689 4568 19858
rect 4620 19712 4672 19718
rect 4526 19680 4582 19689
rect 4620 19654 4672 19660
rect 4526 19615 4582 19624
rect 4342 19479 4398 19488
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4080 19400 4200 19428
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3712 19281 3740 19314
rect 3698 19272 3754 19281
rect 3698 19207 3754 19216
rect 3606 19000 3662 19009
rect 3606 18935 3662 18944
rect 3516 18896 3568 18902
rect 3516 18838 3568 18844
rect 3528 18737 3556 18838
rect 3712 18766 3740 19207
rect 3790 19000 3846 19009
rect 3790 18935 3846 18944
rect 4080 18952 4108 19400
rect 4632 19156 4660 19654
rect 4724 19378 4752 20295
rect 4816 20284 4966 20312
rect 4938 19922 4966 20284
rect 4896 19916 4966 19922
rect 4948 19866 4966 19916
rect 4896 19858 4948 19864
rect 4894 19680 4950 19689
rect 4894 19615 4950 19624
rect 4804 19440 4856 19446
rect 4804 19382 4856 19388
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4632 19128 4752 19156
rect 4322 19068 4630 19077
rect 4322 19066 4328 19068
rect 4384 19066 4408 19068
rect 4464 19066 4488 19068
rect 4544 19066 4568 19068
rect 4624 19066 4630 19068
rect 4384 19014 4386 19066
rect 4566 19014 4568 19066
rect 4322 19012 4328 19014
rect 4384 19012 4408 19014
rect 4464 19012 4488 19014
rect 4544 19012 4568 19014
rect 4624 19012 4630 19014
rect 4322 19003 4630 19012
rect 3700 18760 3752 18766
rect 3514 18728 3570 18737
rect 3700 18702 3752 18708
rect 3804 18698 3832 18935
rect 4080 18924 4200 18952
rect 4066 18864 4122 18873
rect 4066 18799 4122 18808
rect 3514 18663 3570 18672
rect 3792 18692 3844 18698
rect 3792 18634 3844 18640
rect 3424 18624 3476 18630
rect 3608 18624 3660 18630
rect 3424 18566 3476 18572
rect 3528 18584 3608 18612
rect 3436 18136 3464 18566
rect 3528 18272 3556 18584
rect 3608 18566 3660 18572
rect 3662 18524 3970 18533
rect 3662 18522 3668 18524
rect 3724 18522 3748 18524
rect 3804 18522 3828 18524
rect 3884 18522 3908 18524
rect 3964 18522 3970 18524
rect 3724 18470 3726 18522
rect 3906 18470 3908 18522
rect 3662 18468 3668 18470
rect 3724 18468 3748 18470
rect 3804 18468 3828 18470
rect 3884 18468 3908 18470
rect 3964 18468 3970 18470
rect 3662 18459 3970 18468
rect 4080 18290 4108 18799
rect 3608 18284 3660 18290
rect 3528 18244 3608 18272
rect 3608 18226 3660 18232
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 4066 18184 4122 18193
rect 3516 18148 3568 18154
rect 3436 18108 3516 18136
rect 3332 18080 3384 18086
rect 3436 18057 3464 18108
rect 3516 18090 3568 18096
rect 3332 18022 3384 18028
rect 3422 18048 3478 18057
rect 3148 17876 3200 17882
rect 3148 17818 3200 17824
rect 3240 17876 3292 17882
rect 3240 17818 3292 17824
rect 3344 17814 3372 18022
rect 3422 17983 3478 17992
rect 3712 17882 3740 18158
rect 4066 18119 4122 18128
rect 4080 18086 4108 18119
rect 4068 18080 4120 18086
rect 4068 18022 4120 18028
rect 3424 17876 3476 17882
rect 3700 17876 3752 17882
rect 3476 17836 3556 17864
rect 3424 17818 3476 17824
rect 3332 17808 3384 17814
rect 3332 17750 3384 17756
rect 3422 17776 3478 17785
rect 3422 17711 3478 17720
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3240 17536 3292 17542
rect 3240 17478 3292 17484
rect 3160 17134 3188 17478
rect 3148 17128 3200 17134
rect 3252 17126 3280 17478
rect 3344 17338 3372 17614
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3252 17098 3372 17126
rect 3148 17070 3200 17076
rect 3240 17060 3292 17066
rect 3240 17002 3292 17008
rect 3148 14952 3200 14958
rect 3252 14940 3280 17002
rect 3344 16998 3372 17098
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3436 15178 3464 17711
rect 3528 15960 3556 17836
rect 3700 17818 3752 17824
rect 3884 17876 3936 17882
rect 3936 17836 4016 17864
rect 3884 17818 3936 17824
rect 3882 17776 3938 17785
rect 3882 17711 3938 17720
rect 3896 17678 3924 17711
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3988 17610 4016 17836
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 3976 17604 4028 17610
rect 3976 17546 4028 17552
rect 3662 17436 3970 17445
rect 3662 17434 3668 17436
rect 3724 17434 3748 17436
rect 3804 17434 3828 17436
rect 3884 17434 3908 17436
rect 3964 17434 3970 17436
rect 3724 17382 3726 17434
rect 3906 17382 3908 17434
rect 3662 17380 3668 17382
rect 3724 17380 3748 17382
rect 3804 17380 3828 17382
rect 3884 17380 3908 17382
rect 3964 17380 3970 17382
rect 3662 17371 3970 17380
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3896 16726 3924 17206
rect 4080 16794 4108 17750
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3662 16348 3970 16357
rect 3662 16346 3668 16348
rect 3724 16346 3748 16348
rect 3804 16346 3828 16348
rect 3884 16346 3908 16348
rect 3964 16346 3970 16348
rect 3724 16294 3726 16346
rect 3906 16294 3908 16346
rect 3662 16292 3668 16294
rect 3724 16292 3748 16294
rect 3804 16292 3828 16294
rect 3884 16292 3908 16294
rect 3964 16292 3970 16294
rect 3662 16283 3970 16292
rect 3528 15932 3648 15960
rect 3514 15872 3570 15881
rect 3514 15807 3570 15816
rect 3528 15706 3556 15807
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3620 15638 3648 15932
rect 4172 15706 4200 18924
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4252 18352 4304 18358
rect 4252 18294 4304 18300
rect 4264 18222 4292 18294
rect 4252 18216 4304 18222
rect 4356 18193 4384 18702
rect 4252 18158 4304 18164
rect 4342 18184 4398 18193
rect 4342 18119 4398 18128
rect 4540 18086 4568 18770
rect 4632 18154 4660 18770
rect 4724 18737 4752 19128
rect 4710 18728 4766 18737
rect 4710 18663 4766 18672
rect 4816 18358 4844 19382
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4620 18148 4672 18154
rect 4620 18090 4672 18096
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4528 18080 4580 18086
rect 4528 18022 4580 18028
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4264 17882 4292 18022
rect 4322 17980 4630 17989
rect 4322 17978 4328 17980
rect 4384 17978 4408 17980
rect 4464 17978 4488 17980
rect 4544 17978 4568 17980
rect 4624 17978 4630 17980
rect 4384 17926 4386 17978
rect 4566 17926 4568 17978
rect 4322 17924 4328 17926
rect 4384 17924 4408 17926
rect 4464 17924 4488 17926
rect 4544 17924 4568 17926
rect 4624 17924 4630 17926
rect 4322 17915 4630 17924
rect 4252 17876 4304 17882
rect 4252 17818 4304 17824
rect 4436 17876 4488 17882
rect 4436 17818 4488 17824
rect 4264 17746 4292 17818
rect 4252 17740 4304 17746
rect 4252 17682 4304 17688
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4160 15700 4212 15706
rect 4080 15660 4160 15688
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3516 15496 3568 15502
rect 3516 15438 3568 15444
rect 3200 14912 3280 14940
rect 3148 14894 3200 14900
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3160 12238 3188 14554
rect 3252 14482 3280 14912
rect 3344 15150 3464 15178
rect 3240 14476 3292 14482
rect 3240 14418 3292 14424
rect 3252 13802 3280 14418
rect 3240 13796 3292 13802
rect 3240 13738 3292 13744
rect 3240 13388 3292 13394
rect 3240 13330 3292 13336
rect 3252 12986 3280 13330
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10146 2820 10406
rect 2976 10282 3004 10542
rect 3148 10532 3200 10538
rect 3148 10474 3200 10480
rect 2700 10118 2820 10146
rect 2884 10254 3004 10282
rect 3056 10260 3108 10266
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9042 2268 9998
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2240 8838 2268 8978
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 7886 2268 8774
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7342 2268 7822
rect 2332 7342 2360 8366
rect 2424 8090 2452 9522
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2504 8424 2556 8430
rect 2504 8366 2556 8372
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2424 7546 2452 7822
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2136 7268 2188 7274
rect 2136 7210 2188 7216
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 6866 1716 7142
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1492 6180 1544 6186
rect 1492 6122 1544 6128
rect 1504 6066 1532 6122
rect 1412 6038 1532 6066
rect 1122 5264 1178 5273
rect 1122 5199 1178 5208
rect 386 4720 442 4729
rect 386 4655 442 4664
rect 1412 4078 1440 6038
rect 1872 5778 1900 6666
rect 1860 5772 1912 5778
rect 1860 5714 1912 5720
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 1358 1440 4014
rect 1676 4004 1728 4010
rect 1676 3946 1728 3952
rect 1688 3738 1716 3946
rect 1676 3732 1728 3738
rect 1676 3674 1728 3680
rect 1872 3534 1900 5714
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 3194 1532 3334
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1964 3058 1992 6938
rect 2148 6934 2176 7210
rect 2136 6928 2188 6934
rect 2136 6870 2188 6876
rect 2332 6866 2360 7278
rect 2424 7002 2452 7278
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2044 6792 2096 6798
rect 2044 6734 2096 6740
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2056 3398 2084 6734
rect 2148 5914 2176 6734
rect 2332 6458 2360 6802
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2332 5914 2360 6394
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2148 5624 2176 5850
rect 2412 5772 2464 5778
rect 2516 5760 2544 8366
rect 2608 7936 2636 8434
rect 2700 8242 2728 10118
rect 2884 9674 2912 10254
rect 3056 10202 3108 10208
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2792 9646 2912 9674
rect 2792 8344 2820 9646
rect 2872 9376 2924 9382
rect 2872 9318 2924 9324
rect 2884 9042 2912 9318
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2792 8316 2912 8344
rect 2700 8214 2820 8242
rect 2792 7954 2820 8214
rect 2688 7948 2740 7954
rect 2608 7908 2688 7936
rect 2688 7890 2740 7896
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2700 6914 2728 7890
rect 2884 7886 2912 8316
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2792 7546 2820 7686
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2884 7410 2912 7822
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2976 7342 3004 10066
rect 3068 8362 3096 10202
rect 3160 9722 3188 10474
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3160 8634 3188 8910
rect 3252 8634 3280 12038
rect 3344 10742 3372 15150
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3436 14482 3464 15030
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3424 13796 3476 13802
rect 3424 13738 3476 13744
rect 3436 12374 3464 13738
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3332 10736 3384 10742
rect 3528 10690 3556 15438
rect 3662 15260 3970 15269
rect 3662 15258 3668 15260
rect 3724 15258 3748 15260
rect 3804 15258 3828 15260
rect 3884 15258 3908 15260
rect 3964 15258 3970 15260
rect 3724 15206 3726 15258
rect 3906 15206 3908 15258
rect 3662 15204 3668 15206
rect 3724 15204 3748 15206
rect 3804 15204 3828 15206
rect 3884 15204 3908 15206
rect 3964 15204 3970 15206
rect 3662 15195 3970 15204
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 3698 14920 3754 14929
rect 3698 14855 3754 14864
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 3620 14278 3648 14418
rect 3712 14414 3740 14855
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3988 14278 4016 14991
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3662 14172 3970 14181
rect 3662 14170 3668 14172
rect 3724 14170 3748 14172
rect 3804 14170 3828 14172
rect 3884 14170 3908 14172
rect 3964 14170 3970 14172
rect 3724 14118 3726 14170
rect 3906 14118 3908 14170
rect 3662 14116 3668 14118
rect 3724 14116 3748 14118
rect 3804 14116 3828 14118
rect 3884 14116 3908 14118
rect 3964 14116 3970 14118
rect 3662 14107 3970 14116
rect 4080 13326 4108 15660
rect 4160 15642 4212 15648
rect 4264 15570 4292 17546
rect 4448 17270 4476 17818
rect 4816 17785 4844 18022
rect 4802 17776 4858 17785
rect 4802 17711 4804 17720
rect 4856 17711 4858 17720
rect 4804 17682 4856 17688
rect 4528 17536 4580 17542
rect 4528 17478 4580 17484
rect 4804 17536 4856 17542
rect 4804 17478 4856 17484
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4540 17202 4568 17478
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 4540 17105 4568 17138
rect 4816 17134 4844 17478
rect 4804 17128 4856 17134
rect 4526 17096 4582 17105
rect 4804 17070 4856 17076
rect 4526 17031 4582 17040
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4322 16892 4630 16901
rect 4322 16890 4328 16892
rect 4384 16890 4408 16892
rect 4464 16890 4488 16892
rect 4544 16890 4568 16892
rect 4624 16890 4630 16892
rect 4384 16838 4386 16890
rect 4566 16838 4568 16890
rect 4322 16836 4328 16838
rect 4384 16836 4408 16838
rect 4464 16836 4488 16838
rect 4544 16836 4568 16838
rect 4624 16836 4630 16838
rect 4322 16827 4630 16836
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4436 16584 4488 16590
rect 4434 16552 4436 16561
rect 4488 16552 4490 16561
rect 4434 16487 4490 16496
rect 4322 15804 4630 15813
rect 4322 15802 4328 15804
rect 4384 15802 4408 15804
rect 4464 15802 4488 15804
rect 4544 15802 4568 15804
rect 4624 15802 4630 15804
rect 4384 15750 4386 15802
rect 4566 15750 4568 15802
rect 4322 15748 4328 15750
rect 4384 15748 4408 15750
rect 4464 15748 4488 15750
rect 4544 15748 4568 15750
rect 4624 15748 4630 15750
rect 4322 15739 4630 15748
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4172 15065 4200 15438
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4158 15056 4214 15065
rect 4158 14991 4214 15000
rect 4540 14958 4568 15302
rect 4632 14958 4660 15506
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4528 14952 4580 14958
rect 4528 14894 4580 14900
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4172 14618 4200 14894
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4264 14550 4292 14894
rect 4322 14716 4630 14725
rect 4322 14714 4328 14716
rect 4384 14714 4408 14716
rect 4464 14714 4488 14716
rect 4544 14714 4568 14716
rect 4624 14714 4630 14716
rect 4384 14662 4386 14714
rect 4566 14662 4568 14714
rect 4322 14660 4328 14662
rect 4384 14660 4408 14662
rect 4464 14660 4488 14662
rect 4544 14660 4568 14662
rect 4624 14660 4630 14662
rect 4322 14651 4630 14660
rect 4252 14544 4304 14550
rect 4158 14512 4214 14521
rect 4252 14486 4304 14492
rect 4158 14447 4214 14456
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 4172 13138 4200 14447
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4356 13802 4384 14214
rect 4344 13796 4396 13802
rect 4344 13738 4396 13744
rect 4322 13628 4630 13637
rect 4322 13626 4328 13628
rect 4384 13626 4408 13628
rect 4464 13626 4488 13628
rect 4544 13626 4568 13628
rect 4624 13626 4630 13628
rect 4384 13574 4386 13626
rect 4566 13574 4568 13626
rect 4322 13572 4328 13574
rect 4384 13572 4408 13574
rect 4464 13572 4488 13574
rect 4544 13572 4568 13574
rect 4624 13572 4630 13574
rect 4322 13563 4630 13572
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4080 13110 4200 13138
rect 4436 13184 4488 13190
rect 4436 13126 4488 13132
rect 3662 13084 3970 13093
rect 3662 13082 3668 13084
rect 3724 13082 3748 13084
rect 3804 13082 3828 13084
rect 3884 13082 3908 13084
rect 3964 13082 3970 13084
rect 3724 13030 3726 13082
rect 3906 13030 3908 13082
rect 3662 13028 3668 13030
rect 3724 13028 3748 13030
rect 3804 13028 3828 13030
rect 3884 13028 3908 13030
rect 3964 13028 3970 13030
rect 3662 13019 3970 13028
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 3988 12306 4016 12650
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3662 11996 3970 12005
rect 3662 11994 3668 11996
rect 3724 11994 3748 11996
rect 3804 11994 3828 11996
rect 3884 11994 3908 11996
rect 3964 11994 3970 11996
rect 3724 11942 3726 11994
rect 3906 11942 3908 11994
rect 3662 11940 3668 11942
rect 3724 11940 3748 11942
rect 3804 11940 3828 11942
rect 3884 11940 3908 11942
rect 3964 11940 3970 11942
rect 3662 11931 3970 11940
rect 3662 10908 3970 10917
rect 3662 10906 3668 10908
rect 3724 10906 3748 10908
rect 3804 10906 3828 10908
rect 3884 10906 3908 10908
rect 3964 10906 3970 10908
rect 3724 10854 3726 10906
rect 3906 10854 3908 10906
rect 3662 10852 3668 10854
rect 3724 10852 3748 10854
rect 3804 10852 3828 10854
rect 3884 10852 3908 10854
rect 3964 10852 3970 10854
rect 3662 10843 3970 10852
rect 3976 10804 4028 10810
rect 3976 10746 4028 10752
rect 3332 10678 3384 10684
rect 3436 10662 3556 10690
rect 3332 9988 3384 9994
rect 3332 9930 3384 9936
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3344 8430 3372 9930
rect 3436 9654 3464 10662
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3424 9648 3476 9654
rect 3424 9590 3476 9596
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3436 9178 3464 9454
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 3422 8936 3478 8945
rect 3422 8871 3478 8880
rect 3436 8498 3464 8871
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 3056 7948 3108 7954
rect 3056 7890 3108 7896
rect 3068 7478 3096 7890
rect 3344 7886 3372 8366
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 3068 7154 3096 7414
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2976 7126 3096 7154
rect 2700 6886 2820 6914
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5846 2728 6054
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2464 5732 2544 5760
rect 2412 5714 2464 5720
rect 2228 5636 2280 5642
rect 2148 5596 2228 5624
rect 2228 5578 2280 5584
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2332 5166 2360 5510
rect 2320 5160 2372 5166
rect 2320 5102 2372 5108
rect 2424 5012 2452 5714
rect 2792 5370 2820 6886
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2884 5817 2912 6190
rect 2870 5808 2926 5817
rect 2870 5743 2872 5752
rect 2924 5743 2926 5752
rect 2872 5714 2924 5720
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2332 4984 2452 5012
rect 2044 3392 2096 3398
rect 2044 3334 2096 3340
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2056 1970 2084 3334
rect 2332 3058 2360 4984
rect 2884 4758 2912 5510
rect 2976 5302 3004 7126
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 6254 3096 6598
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5710 3096 6190
rect 3160 5846 3188 7346
rect 3528 6798 3556 10542
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3620 10033 3648 10066
rect 3988 10062 4016 10746
rect 4080 10674 4108 13110
rect 4158 13016 4214 13025
rect 4158 12951 4214 12960
rect 4172 12782 4200 12951
rect 4448 12782 4476 13126
rect 4632 12850 4660 13330
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4172 12345 4200 12718
rect 4264 12424 4292 12718
rect 4322 12540 4630 12549
rect 4322 12538 4328 12540
rect 4384 12538 4408 12540
rect 4464 12538 4488 12540
rect 4544 12538 4568 12540
rect 4624 12538 4630 12540
rect 4384 12486 4386 12538
rect 4566 12486 4568 12538
rect 4322 12484 4328 12486
rect 4384 12484 4408 12486
rect 4464 12484 4488 12486
rect 4544 12484 4568 12486
rect 4624 12484 4630 12486
rect 4322 12475 4630 12484
rect 4724 12442 4752 16730
rect 4816 16726 4844 16934
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14618 4844 14826
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4816 13394 4844 13942
rect 4908 13682 4936 19615
rect 5000 19174 5028 20878
rect 5092 20641 5120 22664
rect 5276 22642 5304 24686
rect 5354 24440 5410 24449
rect 5354 24375 5410 24384
rect 5644 24392 5672 25735
rect 5736 25514 5764 27610
rect 5828 27441 5856 27814
rect 5814 27432 5870 27441
rect 5814 27367 5870 27376
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5828 25702 5856 26522
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5736 25486 5856 25514
rect 5724 24880 5776 24886
rect 5828 24857 5856 25486
rect 5724 24822 5776 24828
rect 5814 24848 5870 24857
rect 5736 24585 5764 24822
rect 5814 24783 5870 24792
rect 5816 24744 5868 24750
rect 5814 24712 5816 24721
rect 5868 24712 5870 24721
rect 5814 24647 5870 24656
rect 5722 24576 5778 24585
rect 5722 24511 5778 24520
rect 5368 24274 5396 24375
rect 5644 24364 5856 24392
rect 5356 24268 5408 24274
rect 5356 24210 5408 24216
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5368 23798 5396 24210
rect 5448 24064 5500 24070
rect 5448 24006 5500 24012
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 5368 22778 5396 23598
rect 5460 23254 5488 24006
rect 5644 23866 5672 24210
rect 5724 24132 5776 24138
rect 5724 24074 5776 24080
rect 5632 23860 5684 23866
rect 5632 23802 5684 23808
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 5448 23248 5500 23254
rect 5448 23190 5500 23196
rect 5356 22772 5408 22778
rect 5356 22714 5408 22720
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5354 22264 5410 22273
rect 5354 22199 5410 22208
rect 5368 21842 5396 22199
rect 5184 21814 5396 21842
rect 5078 20632 5134 20641
rect 5078 20567 5134 20576
rect 5078 20496 5134 20505
rect 5078 20431 5134 20440
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5092 18766 5120 20431
rect 5184 19514 5212 21814
rect 5354 21720 5410 21729
rect 5264 21684 5316 21690
rect 5354 21655 5410 21664
rect 5264 21626 5316 21632
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 18760 5132 18766
rect 5080 18702 5132 18708
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 5000 18193 5028 18634
rect 4986 18184 5042 18193
rect 4986 18119 5042 18128
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 5000 17270 5028 18022
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 4988 17128 5040 17134
rect 4986 17096 4988 17105
rect 5040 17096 5042 17105
rect 4986 17031 5042 17040
rect 4988 16720 5040 16726
rect 4988 16662 5040 16668
rect 5000 13870 5028 16662
rect 5092 16658 5120 18702
rect 5184 18204 5212 19450
rect 5276 19417 5304 21626
rect 5368 21418 5396 21655
rect 5356 21412 5408 21418
rect 5356 21354 5408 21360
rect 5368 21049 5396 21354
rect 5354 21040 5410 21049
rect 5354 20975 5410 20984
rect 5356 20936 5408 20942
rect 5354 20904 5356 20913
rect 5408 20904 5410 20913
rect 5354 20839 5410 20848
rect 5356 20528 5408 20534
rect 5356 20470 5408 20476
rect 5262 19408 5318 19417
rect 5262 19343 5318 19352
rect 5368 18358 5396 20470
rect 5460 19922 5488 23190
rect 5552 21418 5580 23666
rect 5632 23520 5684 23526
rect 5632 23462 5684 23468
rect 5644 23186 5672 23462
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5736 23118 5764 24074
rect 5724 23112 5776 23118
rect 5644 23060 5724 23066
rect 5644 23054 5776 23060
rect 5644 23038 5764 23054
rect 5644 21865 5672 23038
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5736 22642 5764 22918
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5736 22166 5764 22578
rect 5724 22160 5776 22166
rect 5724 22102 5776 22108
rect 5828 22098 5856 24364
rect 5816 22092 5868 22098
rect 5816 22034 5868 22040
rect 5724 22024 5776 22030
rect 5722 21992 5724 22001
rect 5776 21992 5778 22001
rect 5722 21927 5778 21936
rect 5724 21888 5776 21894
rect 5630 21856 5686 21865
rect 5724 21830 5776 21836
rect 5814 21856 5870 21865
rect 5630 21791 5686 21800
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5540 21412 5592 21418
rect 5540 21354 5592 21360
rect 5538 21312 5594 21321
rect 5538 21247 5594 21256
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5446 19680 5502 19689
rect 5446 19615 5502 19624
rect 5460 19446 5488 19615
rect 5448 19440 5500 19446
rect 5448 19382 5500 19388
rect 5552 19310 5580 21247
rect 5644 20602 5672 21490
rect 5736 21486 5764 21830
rect 5814 21791 5870 21800
rect 5828 21690 5856 21791
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5632 20596 5684 20602
rect 5632 20538 5684 20544
rect 5724 20596 5776 20602
rect 5724 20538 5776 20544
rect 5630 20224 5686 20233
rect 5630 20159 5686 20168
rect 5644 20058 5672 20159
rect 5632 20052 5684 20058
rect 5632 19994 5684 20000
rect 5632 19916 5684 19922
rect 5632 19858 5684 19864
rect 5644 19310 5672 19858
rect 5736 19854 5764 20538
rect 5828 20505 5856 20946
rect 5814 20496 5870 20505
rect 5814 20431 5870 20440
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5540 19304 5592 19310
rect 5540 19246 5592 19252
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5446 19000 5502 19009
rect 5446 18935 5502 18944
rect 5460 18902 5488 18935
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5184 18176 5396 18204
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5080 16652 5132 16658
rect 5080 16594 5132 16600
rect 5080 16516 5132 16522
rect 5080 16458 5132 16464
rect 5092 16425 5120 16458
rect 5078 16416 5134 16425
rect 5078 16351 5134 16360
rect 5092 16114 5120 16351
rect 5080 16108 5132 16114
rect 5080 16050 5132 16056
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5092 15094 5120 15506
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5092 14958 5120 15030
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5080 14816 5132 14822
rect 5078 14784 5080 14793
rect 5132 14784 5134 14793
rect 5078 14719 5134 14728
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 5092 14074 5120 14350
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 4988 13864 5040 13870
rect 5040 13824 5120 13852
rect 4988 13806 5040 13812
rect 4908 13654 5028 13682
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4908 12782 4936 13126
rect 4896 12776 4948 12782
rect 4896 12718 4948 12724
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4528 12436 4580 12442
rect 4264 12396 4528 12424
rect 4158 12336 4214 12345
rect 4264 12306 4292 12396
rect 4528 12378 4580 12384
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4434 12336 4490 12345
rect 4158 12271 4214 12280
rect 4252 12300 4304 12306
rect 4252 12242 4304 12248
rect 4344 12300 4396 12306
rect 4434 12271 4436 12280
rect 4344 12242 4396 12248
rect 4488 12271 4490 12280
rect 4436 12242 4488 12248
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11762 4200 12106
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 4172 10810 4200 11698
rect 4356 11626 4384 12242
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11694 4660 12038
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4344 11620 4396 11626
rect 4344 11562 4396 11568
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4160 10600 4212 10606
rect 4160 10542 4212 10548
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10056 4028 10062
rect 3606 10024 3662 10033
rect 3976 9998 4028 10004
rect 3606 9959 3662 9968
rect 3662 9820 3970 9829
rect 3662 9818 3668 9820
rect 3724 9818 3748 9820
rect 3804 9818 3828 9820
rect 3884 9818 3908 9820
rect 3964 9818 3970 9820
rect 3724 9766 3726 9818
rect 3906 9766 3908 9818
rect 3662 9764 3668 9766
rect 3724 9764 3748 9766
rect 3804 9764 3828 9766
rect 3884 9764 3908 9766
rect 3964 9764 3970 9766
rect 3662 9755 3970 9764
rect 3608 9716 3660 9722
rect 3976 9716 4028 9722
rect 3608 9658 3660 9664
rect 3804 9664 3976 9674
rect 3804 9658 4028 9664
rect 3620 8945 3648 9658
rect 3804 9646 4016 9658
rect 4080 9654 4108 10406
rect 4172 10062 4200 10542
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9648 4120 9654
rect 3804 9382 3832 9646
rect 4068 9590 4120 9596
rect 4172 9518 4200 9862
rect 3976 9512 4028 9518
rect 4160 9512 4212 9518
rect 4028 9472 4108 9500
rect 3976 9454 4028 9460
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3792 9376 3844 9382
rect 3792 9318 3844 9324
rect 3896 9330 3924 9386
rect 4080 9382 4108 9472
rect 4160 9454 4212 9460
rect 4068 9376 4120 9382
rect 3896 9302 4016 9330
rect 4068 9318 4120 9324
rect 3988 9178 4016 9302
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3606 8936 3662 8945
rect 3606 8871 3662 8880
rect 3662 8732 3970 8741
rect 3662 8730 3668 8732
rect 3724 8730 3748 8732
rect 3804 8730 3828 8732
rect 3884 8730 3908 8732
rect 3964 8730 3970 8732
rect 3724 8678 3726 8730
rect 3906 8678 3908 8730
rect 3662 8676 3668 8678
rect 3724 8676 3748 8678
rect 3804 8676 3828 8678
rect 3884 8676 3908 8678
rect 3964 8676 3970 8678
rect 3662 8667 3970 8676
rect 4080 8430 4108 9318
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3620 8090 3648 8366
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3662 7644 3970 7653
rect 3662 7642 3668 7644
rect 3724 7642 3748 7644
rect 3804 7642 3828 7644
rect 3884 7642 3908 7644
rect 3964 7642 3970 7644
rect 3724 7590 3726 7642
rect 3906 7590 3908 7642
rect 3662 7588 3668 7590
rect 3724 7588 3748 7590
rect 3804 7588 3828 7590
rect 3884 7588 3908 7590
rect 3964 7588 3970 7590
rect 3662 7579 3970 7588
rect 4172 6848 4200 8774
rect 4264 6866 4292 11494
rect 4322 11452 4630 11461
rect 4322 11450 4328 11452
rect 4384 11450 4408 11452
rect 4464 11450 4488 11452
rect 4544 11450 4568 11452
rect 4624 11450 4630 11452
rect 4384 11398 4386 11450
rect 4566 11398 4568 11450
rect 4322 11396 4328 11398
rect 4384 11396 4408 11398
rect 4464 11396 4488 11398
rect 4544 11396 4568 11398
rect 4624 11396 4630 11398
rect 4322 11387 4630 11396
rect 4724 11354 4752 11562
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4322 10364 4630 10373
rect 4322 10362 4328 10364
rect 4384 10362 4408 10364
rect 4464 10362 4488 10364
rect 4544 10362 4568 10364
rect 4624 10362 4630 10364
rect 4384 10310 4386 10362
rect 4566 10310 4568 10362
rect 4322 10308 4328 10310
rect 4384 10308 4408 10310
rect 4464 10308 4488 10310
rect 4544 10308 4568 10310
rect 4624 10308 4630 10310
rect 4322 10299 4630 10308
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 4632 10130 4660 10202
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4356 9722 4384 9998
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4322 9276 4630 9285
rect 4322 9274 4328 9276
rect 4384 9274 4408 9276
rect 4464 9274 4488 9276
rect 4544 9274 4568 9276
rect 4624 9274 4630 9276
rect 4384 9222 4386 9274
rect 4566 9222 4568 9274
rect 4322 9220 4328 9222
rect 4384 9220 4408 9222
rect 4464 9220 4488 9222
rect 4544 9220 4568 9222
rect 4624 9220 4630 9222
rect 4322 9211 4630 9220
rect 4526 8936 4582 8945
rect 4526 8871 4582 8880
rect 4540 8430 4568 8871
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4632 8362 4660 8774
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4322 8188 4630 8197
rect 4322 8186 4328 8188
rect 4384 8186 4408 8188
rect 4464 8186 4488 8188
rect 4544 8186 4568 8188
rect 4624 8186 4630 8188
rect 4384 8134 4386 8186
rect 4566 8134 4568 8186
rect 4322 8132 4328 8134
rect 4384 8132 4408 8134
rect 4464 8132 4488 8134
rect 4544 8132 4568 8134
rect 4624 8132 4630 8134
rect 4322 8123 4630 8132
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4448 7818 4476 8026
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4540 7546 4568 7890
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4632 7274 4660 7686
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4322 7100 4630 7109
rect 4322 7098 4328 7100
rect 4384 7098 4408 7100
rect 4464 7098 4488 7100
rect 4544 7098 4568 7100
rect 4624 7098 4630 7100
rect 4384 7046 4386 7098
rect 4566 7046 4568 7098
rect 4322 7044 4328 7046
rect 4384 7044 4408 7046
rect 4464 7044 4488 7046
rect 4544 7044 4568 7046
rect 4624 7044 4630 7046
rect 4322 7035 4630 7044
rect 4724 6984 4752 11018
rect 4816 10130 4844 12582
rect 4908 12238 4936 12718
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 5000 12186 5028 13654
rect 5092 12288 5120 13824
rect 5184 12918 5212 17478
rect 5276 17338 5304 17750
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5262 16960 5318 16969
rect 5262 16895 5318 16904
rect 5276 16454 5304 16895
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5368 14906 5396 18176
rect 5460 17814 5488 18838
rect 5552 18766 5580 19246
rect 5632 18828 5684 18834
rect 5632 18770 5684 18776
rect 5540 18760 5592 18766
rect 5540 18702 5592 18708
rect 5644 18154 5672 18770
rect 5632 18148 5684 18154
rect 5632 18090 5684 18096
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5448 17604 5500 17610
rect 5448 17546 5500 17552
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5276 14878 5396 14906
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5276 12481 5304 14878
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5368 14414 5396 14758
rect 5356 14408 5408 14414
rect 5356 14350 5408 14356
rect 5460 14362 5488 17546
rect 5552 17134 5580 17546
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5644 16980 5672 18090
rect 5736 17814 5764 19654
rect 5828 18426 5856 20334
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5816 18216 5868 18222
rect 5816 18158 5868 18164
rect 5724 17808 5776 17814
rect 5724 17750 5776 17756
rect 5828 17660 5856 18158
rect 5736 17632 5856 17660
rect 5736 17134 5764 17632
rect 5920 17134 5948 27814
rect 6012 27010 6040 27934
rect 6104 27656 6132 29446
rect 6196 28218 6224 29593
rect 6368 29096 6420 29102
rect 6472 29073 6500 30738
rect 6564 30394 6592 31214
rect 6736 31214 6788 31220
rect 6642 31175 6698 31184
rect 6552 30388 6604 30394
rect 6552 30330 6604 30336
rect 6564 30297 6592 30330
rect 6550 30288 6606 30297
rect 6550 30223 6606 30232
rect 6656 30190 6684 31175
rect 6748 30394 6776 31214
rect 6736 30388 6788 30394
rect 6736 30330 6788 30336
rect 6736 30252 6788 30258
rect 6840 30240 6868 31583
rect 6932 31482 6960 32778
rect 7024 32502 7052 33050
rect 7104 32768 7156 32774
rect 7104 32710 7156 32716
rect 7116 32570 7144 32710
rect 7104 32564 7156 32570
rect 7104 32506 7156 32512
rect 7012 32496 7064 32502
rect 7012 32438 7064 32444
rect 7012 32292 7064 32298
rect 7012 32234 7064 32240
rect 7024 32026 7052 32234
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 7012 31748 7064 31754
rect 7012 31690 7064 31696
rect 7024 31521 7052 31690
rect 7116 31686 7144 32506
rect 7104 31680 7156 31686
rect 7104 31622 7156 31628
rect 7010 31512 7066 31521
rect 6920 31476 6972 31482
rect 7010 31447 7066 31456
rect 6920 31418 6972 31424
rect 7208 31414 7236 35566
rect 7286 35527 7288 35536
rect 7340 35527 7342 35536
rect 7288 35498 7340 35504
rect 7392 35086 7420 35974
rect 7470 35935 7526 35944
rect 7484 35766 7512 35935
rect 7472 35760 7524 35766
rect 7472 35702 7524 35708
rect 7472 35148 7524 35154
rect 7472 35090 7524 35096
rect 7564 35148 7616 35154
rect 7564 35090 7616 35096
rect 7380 35080 7432 35086
rect 7380 35022 7432 35028
rect 7288 34944 7340 34950
rect 7288 34886 7340 34892
rect 7300 33114 7328 34886
rect 7392 34542 7420 35022
rect 7484 35018 7512 35090
rect 7472 35012 7524 35018
rect 7472 34954 7524 34960
rect 7380 34536 7432 34542
rect 7380 34478 7432 34484
rect 7392 34066 7420 34478
rect 7380 34060 7432 34066
rect 7380 34002 7432 34008
rect 7380 33856 7432 33862
rect 7380 33798 7432 33804
rect 7392 33318 7420 33798
rect 7380 33312 7432 33318
rect 7380 33254 7432 33260
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7288 32972 7340 32978
rect 7288 32914 7340 32920
rect 7300 32745 7328 32914
rect 7286 32736 7342 32745
rect 7286 32671 7342 32680
rect 7286 32328 7342 32337
rect 7286 32263 7342 32272
rect 7300 32230 7328 32263
rect 7288 32224 7340 32230
rect 7288 32166 7340 32172
rect 7288 31680 7340 31686
rect 7288 31622 7340 31628
rect 7196 31408 7248 31414
rect 7196 31350 7248 31356
rect 7300 31278 7328 31622
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 7196 31272 7248 31278
rect 7196 31214 7248 31220
rect 7288 31272 7340 31278
rect 7288 31214 7340 31220
rect 6932 30326 6960 31214
rect 7012 31136 7064 31142
rect 7012 31078 7064 31084
rect 7024 30802 7052 31078
rect 7104 30932 7156 30938
rect 7104 30874 7156 30880
rect 7012 30796 7064 30802
rect 7012 30738 7064 30744
rect 7116 30705 7144 30874
rect 7102 30696 7158 30705
rect 7102 30631 7158 30640
rect 7208 30394 7236 31214
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 7012 30388 7064 30394
rect 7012 30330 7064 30336
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 6788 30212 6868 30240
rect 6736 30194 6788 30200
rect 6644 30184 6696 30190
rect 6644 30126 6696 30132
rect 6552 29708 6604 29714
rect 6552 29650 6604 29656
rect 6564 29510 6592 29650
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 6368 29038 6420 29044
rect 6458 29064 6514 29073
rect 6380 28937 6408 29038
rect 6458 28999 6514 29008
rect 6366 28928 6422 28937
rect 6366 28863 6422 28872
rect 6274 28792 6330 28801
rect 6274 28727 6330 28736
rect 6288 28694 6316 28727
rect 6276 28688 6328 28694
rect 6276 28630 6328 28636
rect 6564 28558 6592 29446
rect 6656 29102 6684 30126
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6368 28484 6420 28490
rect 6368 28426 6420 28432
rect 6276 28416 6328 28422
rect 6274 28384 6276 28393
rect 6328 28384 6330 28393
rect 6274 28319 6330 28328
rect 6184 28212 6236 28218
rect 6184 28154 6236 28160
rect 6104 27628 6316 27656
rect 6092 27532 6144 27538
rect 6092 27474 6144 27480
rect 6104 27130 6132 27474
rect 6184 27328 6236 27334
rect 6184 27270 6236 27276
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6196 27062 6224 27270
rect 6184 27056 6236 27062
rect 6012 26982 6132 27010
rect 6184 26998 6236 27004
rect 6000 26920 6052 26926
rect 6000 26862 6052 26868
rect 6012 26042 6040 26862
rect 6000 26036 6052 26042
rect 6000 25978 6052 25984
rect 6104 25242 6132 26982
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6196 26586 6224 26862
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6182 26480 6238 26489
rect 6182 26415 6238 26424
rect 6012 25214 6132 25242
rect 6012 21457 6040 25214
rect 6092 24676 6144 24682
rect 6092 24618 6144 24624
rect 6104 24206 6132 24618
rect 6092 24200 6144 24206
rect 6092 24142 6144 24148
rect 6092 24064 6144 24070
rect 6092 24006 6144 24012
rect 6104 23730 6132 24006
rect 6092 23724 6144 23730
rect 6092 23666 6144 23672
rect 6090 23352 6146 23361
rect 6090 23287 6092 23296
rect 6144 23287 6146 23296
rect 6092 23258 6144 23264
rect 6104 23118 6132 23258
rect 6092 23112 6144 23118
rect 6092 23054 6144 23060
rect 6104 22273 6132 23054
rect 6090 22264 6146 22273
rect 6090 22199 6146 22208
rect 6196 22094 6224 26415
rect 6288 24585 6316 27628
rect 6380 26994 6408 28426
rect 6460 27668 6512 27674
rect 6460 27610 6512 27616
rect 6368 26988 6420 26994
rect 6368 26930 6420 26936
rect 6368 26784 6420 26790
rect 6368 26726 6420 26732
rect 6380 26450 6408 26726
rect 6368 26444 6420 26450
rect 6368 26386 6420 26392
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6380 25362 6408 26250
rect 6368 25356 6420 25362
rect 6368 25298 6420 25304
rect 6274 24576 6330 24585
rect 6274 24511 6330 24520
rect 6274 24440 6330 24449
rect 6274 24375 6330 24384
rect 6288 24274 6316 24375
rect 6380 24313 6408 25298
rect 6472 24834 6500 27610
rect 6564 27577 6592 28494
rect 6656 28082 6684 28562
rect 6644 28076 6696 28082
rect 6644 28018 6696 28024
rect 6642 27840 6698 27849
rect 6642 27775 6698 27784
rect 6550 27568 6606 27577
rect 6550 27503 6606 27512
rect 6656 26874 6684 27775
rect 6748 27441 6776 30194
rect 7024 30122 7052 30330
rect 7300 30274 7328 30670
rect 7208 30246 7328 30274
rect 7104 30184 7156 30190
rect 7102 30152 7104 30161
rect 7156 30152 7158 30161
rect 6920 30116 6972 30122
rect 6920 30058 6972 30064
rect 7012 30116 7064 30122
rect 7102 30087 7158 30096
rect 7012 30058 7064 30064
rect 6932 29832 6960 30058
rect 7104 29844 7156 29850
rect 6932 29804 7104 29832
rect 7104 29786 7156 29792
rect 6920 29640 6972 29646
rect 6972 29600 7052 29628
rect 6920 29582 6972 29588
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 6828 29028 6880 29034
rect 6828 28970 6880 28976
rect 6840 28150 6868 28970
rect 6828 28144 6880 28150
rect 6828 28086 6880 28092
rect 6932 27826 6960 29038
rect 6840 27798 6960 27826
rect 6840 27538 6868 27798
rect 6918 27704 6974 27713
rect 7024 27674 7052 29600
rect 7116 29034 7144 29786
rect 7104 29028 7156 29034
rect 7104 28970 7156 28976
rect 7116 28121 7144 28970
rect 7208 28665 7236 30246
rect 7288 30184 7340 30190
rect 7288 30126 7340 30132
rect 7300 28966 7328 30126
rect 7392 29782 7420 33254
rect 7484 32842 7512 34954
rect 7576 34202 7604 35090
rect 7668 34542 7696 36094
rect 7840 36100 7892 36106
rect 7840 36042 7892 36048
rect 7852 35034 7880 36042
rect 8128 36038 8156 36751
rect 8220 36310 8248 37742
rect 8312 37330 8340 38286
rect 8404 37369 8432 40394
rect 8496 38321 8524 40870
rect 8668 40724 8720 40730
rect 8668 40666 8720 40672
rect 8680 39982 8708 40666
rect 8760 40520 8812 40526
rect 8760 40462 8812 40468
rect 8668 39976 8720 39982
rect 8668 39918 8720 39924
rect 8576 39364 8628 39370
rect 8576 39306 8628 39312
rect 8588 38654 8616 39306
rect 8666 39264 8722 39273
rect 8666 39199 8722 39208
rect 8680 38962 8708 39199
rect 8668 38956 8720 38962
rect 8668 38898 8720 38904
rect 8772 38894 8800 40462
rect 8956 39982 8984 41006
rect 9128 40928 9180 40934
rect 9180 40888 9260 40916
rect 9128 40870 9180 40876
rect 9232 40594 9260 40888
rect 9128 40588 9180 40594
rect 9128 40530 9180 40536
rect 9220 40588 9272 40594
rect 9220 40530 9272 40536
rect 9140 40186 9168 40530
rect 9220 40384 9272 40390
rect 9220 40326 9272 40332
rect 9128 40180 9180 40186
rect 9128 40122 9180 40128
rect 9232 40066 9260 40326
rect 9324 40225 9352 41006
rect 9310 40216 9366 40225
rect 9310 40151 9366 40160
rect 9140 40038 9260 40066
rect 8944 39976 8996 39982
rect 8944 39918 8996 39924
rect 8852 39500 8904 39506
rect 8852 39442 8904 39448
rect 8760 38888 8812 38894
rect 8760 38830 8812 38836
rect 8864 38654 8892 39442
rect 8944 39296 8996 39302
rect 8944 39238 8996 39244
rect 8956 38758 8984 39238
rect 9036 38820 9088 38826
rect 9036 38762 9088 38768
rect 8944 38752 8996 38758
rect 8944 38694 8996 38700
rect 8588 38626 8708 38654
rect 8864 38626 8984 38654
rect 8680 38350 8708 38626
rect 8668 38344 8720 38350
rect 8482 38312 8538 38321
rect 8666 38312 8668 38321
rect 8720 38312 8722 38321
rect 8482 38247 8538 38256
rect 8576 38276 8628 38282
rect 8666 38247 8722 38256
rect 8576 38218 8628 38224
rect 8588 37806 8616 38218
rect 8668 38208 8720 38214
rect 8666 38176 8668 38185
rect 8760 38208 8812 38214
rect 8720 38176 8722 38185
rect 8760 38150 8812 38156
rect 8666 38111 8722 38120
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 8576 37800 8628 37806
rect 8576 37742 8628 37748
rect 8668 37800 8720 37806
rect 8772 37788 8800 38150
rect 8956 37806 8984 38626
rect 9048 38554 9076 38762
rect 9036 38548 9088 38554
rect 9036 38490 9088 38496
rect 9034 38448 9090 38457
rect 9034 38383 9036 38392
rect 9088 38383 9090 38392
rect 9036 38354 9088 38360
rect 8720 37760 8800 37788
rect 8944 37800 8996 37806
rect 8850 37768 8906 37777
rect 8668 37742 8720 37748
rect 8390 37360 8446 37369
rect 8300 37324 8352 37330
rect 8390 37295 8446 37304
rect 8300 37266 8352 37272
rect 8496 37233 8524 37742
rect 8482 37224 8538 37233
rect 8392 37188 8444 37194
rect 8482 37159 8538 37168
rect 8392 37130 8444 37136
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8312 36700 8340 36858
rect 8404 36854 8432 37130
rect 8392 36848 8444 36854
rect 8392 36790 8444 36796
rect 8496 36802 8524 37159
rect 8576 37120 8628 37126
rect 8576 37062 8628 37068
rect 8588 36922 8616 37062
rect 8680 36922 8708 37742
rect 8944 37742 8996 37748
rect 8850 37703 8906 37712
rect 8864 37466 8892 37703
rect 8852 37460 8904 37466
rect 8852 37402 8904 37408
rect 8760 37324 8812 37330
rect 8760 37266 8812 37272
rect 8852 37324 8904 37330
rect 8852 37266 8904 37272
rect 8772 37097 8800 37266
rect 8758 37088 8814 37097
rect 8758 37023 8814 37032
rect 8758 36952 8814 36961
rect 8576 36916 8628 36922
rect 8576 36858 8628 36864
rect 8668 36916 8720 36922
rect 8758 36887 8760 36896
rect 8668 36858 8720 36864
rect 8812 36887 8814 36896
rect 8760 36858 8812 36864
rect 8496 36774 8635 36802
rect 8304 36672 8340 36700
rect 8607 36700 8635 36774
rect 8760 36780 8812 36786
rect 8760 36722 8812 36728
rect 8607 36684 8704 36700
rect 8607 36678 8716 36684
rect 8607 36672 8664 36678
rect 8304 36530 8332 36672
rect 8392 36644 8444 36650
rect 8444 36604 8609 36632
rect 8664 36620 8716 36626
rect 8392 36586 8444 36592
rect 8304 36502 8340 36530
rect 8208 36304 8260 36310
rect 8206 36272 8208 36281
rect 8260 36272 8262 36281
rect 8206 36207 8262 36216
rect 8312 36224 8340 36502
rect 8581 36394 8609 36604
rect 8581 36366 8616 36394
rect 8312 36196 8524 36224
rect 8206 36136 8262 36145
rect 8206 36071 8208 36080
rect 8260 36071 8262 36080
rect 8208 36042 8260 36048
rect 8496 36038 8524 36196
rect 8588 36174 8616 36366
rect 8772 36310 8800 36722
rect 8760 36304 8812 36310
rect 8760 36246 8812 36252
rect 8576 36168 8628 36174
rect 8864 36122 8892 37266
rect 8956 37097 8984 37742
rect 9036 37188 9088 37194
rect 9036 37130 9088 37136
rect 8942 37088 8998 37097
rect 8942 37023 8998 37032
rect 8944 36848 8996 36854
rect 8944 36790 8996 36796
rect 8956 36689 8984 36790
rect 9048 36786 9076 37130
rect 9140 37126 9168 40038
rect 9220 39976 9272 39982
rect 9220 39918 9272 39924
rect 9232 38729 9260 39918
rect 9312 39908 9364 39914
rect 9312 39850 9364 39856
rect 9324 39386 9352 39850
rect 9416 39817 9444 41414
rect 9692 41177 9720 42638
rect 9784 42294 9812 42638
rect 9772 42288 9824 42294
rect 9772 42230 9824 42236
rect 9678 41168 9734 41177
rect 9678 41103 9734 41112
rect 9784 40712 9812 42230
rect 9968 42158 9996 43046
rect 10060 42770 10088 43318
rect 10722 43004 11030 43013
rect 10722 43002 10728 43004
rect 10784 43002 10808 43004
rect 10864 43002 10888 43004
rect 10944 43002 10968 43004
rect 11024 43002 11030 43004
rect 10784 42950 10786 43002
rect 10966 42950 10968 43002
rect 10722 42948 10728 42950
rect 10784 42948 10808 42950
rect 10864 42948 10888 42950
rect 10944 42948 10968 42950
rect 11024 42948 11030 42950
rect 10722 42939 11030 42948
rect 11704 42832 11756 42838
rect 11704 42774 11756 42780
rect 10048 42764 10100 42770
rect 10048 42706 10100 42712
rect 10784 42764 10836 42770
rect 10784 42706 10836 42712
rect 11152 42764 11204 42770
rect 11152 42706 11204 42712
rect 10062 42460 10370 42469
rect 10062 42458 10068 42460
rect 10124 42458 10148 42460
rect 10204 42458 10228 42460
rect 10284 42458 10308 42460
rect 10364 42458 10370 42460
rect 10124 42406 10126 42458
rect 10306 42406 10308 42458
rect 10062 42404 10068 42406
rect 10124 42404 10148 42406
rect 10204 42404 10228 42406
rect 10284 42404 10308 42406
rect 10364 42404 10370 42406
rect 10062 42395 10370 42404
rect 9956 42152 10008 42158
rect 9956 42094 10008 42100
rect 10600 42152 10652 42158
rect 10600 42094 10652 42100
rect 10416 42084 10468 42090
rect 10416 42026 10468 42032
rect 9864 42016 9916 42022
rect 9864 41958 9916 41964
rect 10048 42016 10100 42022
rect 10048 41958 10100 41964
rect 9692 40684 9812 40712
rect 9588 40588 9640 40594
rect 9588 40530 9640 40536
rect 9402 39808 9458 39817
rect 9402 39743 9458 39752
rect 9404 39500 9456 39506
rect 9456 39460 9536 39488
rect 9404 39442 9456 39448
rect 9324 39358 9444 39386
rect 9416 38758 9444 39358
rect 9508 38962 9536 39460
rect 9600 39030 9628 40530
rect 9692 39982 9720 40684
rect 9876 40662 9904 41958
rect 10060 41478 10088 41958
rect 10428 41721 10456 42026
rect 10508 42016 10560 42022
rect 10508 41958 10560 41964
rect 10414 41712 10470 41721
rect 10414 41647 10470 41656
rect 10048 41472 10100 41478
rect 10048 41414 10100 41420
rect 10520 41414 10548 41958
rect 10612 41478 10640 42094
rect 10796 42090 10824 42706
rect 10876 42628 10928 42634
rect 10876 42570 10928 42576
rect 10888 42294 10916 42570
rect 10968 42560 11020 42566
rect 10968 42502 11020 42508
rect 10876 42288 10928 42294
rect 10876 42230 10928 42236
rect 10980 42106 11008 42502
rect 10784 42084 10836 42090
rect 10980 42078 11100 42106
rect 10784 42026 10836 42032
rect 10722 41916 11030 41925
rect 10722 41914 10728 41916
rect 10784 41914 10808 41916
rect 10864 41914 10888 41916
rect 10944 41914 10968 41916
rect 11024 41914 11030 41916
rect 10784 41862 10786 41914
rect 10966 41862 10968 41914
rect 10722 41860 10728 41862
rect 10784 41860 10808 41862
rect 10864 41860 10888 41862
rect 10944 41860 10968 41862
rect 11024 41860 11030 41862
rect 10722 41851 11030 41860
rect 10784 41812 10836 41818
rect 10784 41754 10836 41760
rect 10796 41585 10824 41754
rect 11072 41750 11100 42078
rect 10876 41744 10928 41750
rect 10876 41686 10928 41692
rect 11060 41744 11112 41750
rect 11060 41686 11112 41692
rect 10782 41576 10838 41585
rect 10782 41511 10838 41520
rect 10600 41472 10652 41478
rect 10600 41414 10652 41420
rect 10428 41386 10548 41414
rect 10062 41372 10370 41381
rect 10062 41370 10068 41372
rect 10124 41370 10148 41372
rect 10204 41370 10228 41372
rect 10284 41370 10308 41372
rect 10364 41370 10370 41372
rect 10124 41318 10126 41370
rect 10306 41318 10308 41370
rect 10062 41316 10068 41318
rect 10124 41316 10148 41318
rect 10204 41316 10228 41318
rect 10284 41316 10308 41318
rect 10364 41316 10370 41318
rect 10062 41307 10370 41316
rect 9956 40996 10008 41002
rect 9956 40938 10008 40944
rect 10048 40996 10100 41002
rect 10048 40938 10100 40944
rect 9968 40905 9996 40938
rect 9954 40896 10010 40905
rect 9954 40831 10010 40840
rect 10060 40746 10088 40938
rect 9968 40718 10088 40746
rect 9864 40656 9916 40662
rect 9864 40598 9916 40604
rect 9772 40588 9824 40594
rect 9772 40530 9824 40536
rect 9680 39976 9732 39982
rect 9680 39918 9732 39924
rect 9680 39840 9732 39846
rect 9680 39782 9732 39788
rect 9588 39024 9640 39030
rect 9588 38966 9640 38972
rect 9496 38956 9548 38962
rect 9496 38898 9548 38904
rect 9312 38752 9364 38758
rect 9218 38720 9274 38729
rect 9312 38694 9364 38700
rect 9404 38752 9456 38758
rect 9404 38694 9456 38700
rect 9218 38655 9274 38664
rect 9324 38554 9352 38694
rect 9312 38548 9364 38554
rect 9312 38490 9364 38496
rect 9416 38457 9444 38694
rect 9402 38448 9458 38457
rect 9402 38383 9458 38392
rect 9402 38312 9458 38321
rect 9402 38247 9458 38256
rect 9416 38214 9444 38247
rect 9404 38208 9456 38214
rect 9404 38150 9456 38156
rect 9402 38040 9458 38049
rect 9402 37975 9458 37984
rect 9220 37800 9272 37806
rect 9218 37768 9220 37777
rect 9272 37768 9274 37777
rect 9416 37754 9444 37975
rect 9508 37856 9536 38898
rect 9692 38457 9720 39782
rect 9784 38978 9812 40530
rect 9864 39840 9916 39846
rect 9864 39782 9916 39788
rect 9876 39574 9904 39782
rect 9968 39681 9996 40718
rect 10062 40284 10370 40293
rect 10062 40282 10068 40284
rect 10124 40282 10148 40284
rect 10204 40282 10228 40284
rect 10284 40282 10308 40284
rect 10364 40282 10370 40284
rect 10124 40230 10126 40282
rect 10306 40230 10308 40282
rect 10062 40228 10068 40230
rect 10124 40228 10148 40230
rect 10204 40228 10228 40230
rect 10284 40228 10308 40230
rect 10364 40228 10370 40230
rect 10062 40219 10370 40228
rect 10428 40168 10456 41386
rect 10508 41064 10560 41070
rect 10612 41052 10640 41414
rect 10560 41024 10640 41052
rect 10888 41041 10916 41686
rect 11060 41608 11112 41614
rect 11060 41550 11112 41556
rect 10968 41472 11020 41478
rect 10968 41414 11020 41420
rect 10980 41070 11008 41414
rect 10968 41064 11020 41070
rect 10508 41006 10560 41012
rect 10336 40140 10456 40168
rect 10508 40180 10560 40186
rect 10138 39944 10194 39953
rect 10138 39879 10140 39888
rect 10192 39879 10194 39888
rect 10232 39908 10284 39914
rect 10140 39850 10192 39856
rect 10232 39850 10284 39856
rect 10048 39840 10100 39846
rect 10048 39782 10100 39788
rect 9954 39672 10010 39681
rect 9954 39607 10010 39616
rect 9864 39568 9916 39574
rect 9864 39510 9916 39516
rect 9876 39098 9904 39510
rect 9956 39500 10008 39506
rect 9956 39442 10008 39448
rect 9968 39098 9996 39442
rect 10060 39409 10088 39782
rect 10244 39642 10272 39850
rect 10232 39636 10284 39642
rect 10232 39578 10284 39584
rect 10336 39506 10364 40140
rect 10508 40122 10560 40128
rect 10416 40044 10468 40050
rect 10416 39986 10468 39992
rect 10324 39500 10376 39506
rect 10324 39442 10376 39448
rect 10046 39400 10102 39409
rect 10046 39335 10102 39344
rect 10062 39196 10370 39205
rect 10062 39194 10068 39196
rect 10124 39194 10148 39196
rect 10204 39194 10228 39196
rect 10284 39194 10308 39196
rect 10364 39194 10370 39196
rect 10124 39142 10126 39194
rect 10306 39142 10308 39194
rect 10062 39140 10068 39142
rect 10124 39140 10148 39142
rect 10204 39140 10228 39142
rect 10284 39140 10308 39142
rect 10364 39140 10370 39142
rect 10062 39131 10370 39140
rect 9864 39092 9916 39098
rect 9864 39034 9916 39040
rect 9956 39092 10008 39098
rect 9956 39034 10008 39040
rect 10048 39024 10100 39030
rect 9784 38950 9996 38978
rect 10048 38966 10100 38972
rect 10230 38992 10286 39001
rect 9772 38888 9824 38894
rect 9772 38830 9824 38836
rect 9784 38729 9812 38830
rect 9770 38720 9826 38729
rect 9770 38655 9826 38664
rect 9678 38448 9734 38457
rect 9588 38412 9640 38418
rect 9678 38383 9734 38392
rect 9772 38412 9824 38418
rect 9588 38354 9640 38360
rect 9772 38354 9824 38360
rect 9864 38412 9916 38418
rect 9864 38354 9916 38360
rect 9600 38049 9628 38354
rect 9784 38321 9812 38354
rect 9770 38312 9826 38321
rect 9770 38247 9826 38256
rect 9586 38040 9642 38049
rect 9586 37975 9642 37984
rect 9508 37828 9608 37856
rect 9580 37806 9608 37828
rect 9580 37800 9640 37806
rect 9580 37760 9588 37800
rect 9218 37703 9274 37712
rect 9312 37732 9364 37738
rect 9416 37726 9536 37754
rect 9588 37742 9640 37748
rect 9312 37674 9364 37680
rect 9220 37664 9272 37670
rect 9220 37606 9272 37612
rect 9128 37120 9180 37126
rect 9128 37062 9180 37068
rect 9232 36922 9260 37606
rect 9220 36916 9272 36922
rect 9220 36858 9272 36864
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 9218 36816 9274 36825
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 8942 36680 8998 36689
rect 8942 36615 8998 36624
rect 9036 36644 9088 36650
rect 9036 36586 9088 36592
rect 8942 36544 8998 36553
rect 8942 36479 8998 36488
rect 8956 36310 8984 36479
rect 8944 36304 8996 36310
rect 9048 36281 9076 36586
rect 8944 36246 8996 36252
rect 9034 36272 9090 36281
rect 9034 36207 9090 36216
rect 9140 36122 9168 36790
rect 9218 36751 9274 36760
rect 8576 36110 8628 36116
rect 8772 36094 8892 36122
rect 9048 36094 9168 36122
rect 8116 36032 8168 36038
rect 8116 35974 8168 35980
rect 8392 36032 8444 36038
rect 8392 35974 8444 35980
rect 8484 36032 8536 36038
rect 8484 35974 8536 35980
rect 8404 35834 8432 35974
rect 8666 35864 8722 35873
rect 8392 35828 8444 35834
rect 8666 35799 8722 35808
rect 8392 35770 8444 35776
rect 8114 35592 8170 35601
rect 8298 35592 8354 35601
rect 8114 35527 8116 35536
rect 8168 35527 8170 35536
rect 8208 35556 8260 35562
rect 8116 35498 8168 35504
rect 8298 35527 8354 35536
rect 8208 35498 8260 35504
rect 7748 35012 7800 35018
rect 7852 35006 8156 35034
rect 7748 34954 7800 34960
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7760 34474 7788 34954
rect 7932 34944 7984 34950
rect 7932 34886 7984 34892
rect 7748 34468 7800 34474
rect 7748 34410 7800 34416
rect 7840 34400 7892 34406
rect 7840 34342 7892 34348
rect 7564 34196 7616 34202
rect 7564 34138 7616 34144
rect 7656 34196 7708 34202
rect 7656 34138 7708 34144
rect 7668 33454 7696 34138
rect 7748 33856 7800 33862
rect 7748 33798 7800 33804
rect 7656 33448 7708 33454
rect 7562 33416 7618 33425
rect 7656 33390 7708 33396
rect 7562 33351 7618 33360
rect 7576 33318 7604 33351
rect 7564 33312 7616 33318
rect 7564 33254 7616 33260
rect 7576 32892 7604 33254
rect 7656 32904 7708 32910
rect 7576 32864 7656 32892
rect 7472 32836 7524 32842
rect 7472 32778 7524 32784
rect 7576 32366 7604 32864
rect 7656 32846 7708 32852
rect 7564 32360 7616 32366
rect 7564 32302 7616 32308
rect 7472 32224 7524 32230
rect 7576 32201 7604 32302
rect 7472 32166 7524 32172
rect 7562 32192 7618 32201
rect 7484 30802 7512 32166
rect 7562 32127 7618 32136
rect 7564 31952 7616 31958
rect 7616 31912 7696 31940
rect 7564 31894 7616 31900
rect 7564 31680 7616 31686
rect 7668 31657 7696 31912
rect 7564 31622 7616 31628
rect 7654 31648 7710 31657
rect 7576 31210 7604 31622
rect 7654 31583 7710 31592
rect 7654 31376 7710 31385
rect 7654 31311 7710 31320
rect 7668 31278 7696 31311
rect 7656 31272 7708 31278
rect 7656 31214 7708 31220
rect 7564 31204 7616 31210
rect 7564 31146 7616 31152
rect 7656 31136 7708 31142
rect 7562 31104 7618 31113
rect 7656 31078 7708 31084
rect 7562 31039 7618 31048
rect 7472 30796 7524 30802
rect 7472 30738 7524 30744
rect 7576 30734 7604 31039
rect 7668 30802 7696 31078
rect 7656 30796 7708 30802
rect 7656 30738 7708 30744
rect 7564 30728 7616 30734
rect 7564 30670 7616 30676
rect 7472 30660 7524 30666
rect 7472 30602 7524 30608
rect 7656 30660 7708 30666
rect 7656 30602 7708 30608
rect 7484 30297 7512 30602
rect 7562 30424 7618 30433
rect 7562 30359 7618 30368
rect 7470 30288 7526 30297
rect 7470 30223 7526 30232
rect 7380 29776 7432 29782
rect 7380 29718 7432 29724
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7288 28960 7340 28966
rect 7288 28902 7340 28908
rect 7194 28656 7250 28665
rect 7194 28591 7250 28600
rect 7102 28112 7158 28121
rect 7300 28082 7328 28902
rect 7102 28047 7158 28056
rect 7288 28076 7340 28082
rect 7288 28018 7340 28024
rect 7104 28008 7156 28014
rect 7104 27950 7156 27956
rect 6918 27639 6974 27648
rect 7012 27668 7064 27674
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6734 27432 6790 27441
rect 6734 27367 6790 27376
rect 6734 27296 6790 27305
rect 6734 27231 6790 27240
rect 6564 26846 6684 26874
rect 6564 26489 6592 26846
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6656 26518 6684 26726
rect 6644 26512 6696 26518
rect 6550 26480 6606 26489
rect 6644 26454 6696 26460
rect 6550 26415 6606 26424
rect 6656 26246 6684 26454
rect 6644 26240 6696 26246
rect 6644 26182 6696 26188
rect 6656 25838 6684 26182
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6642 25392 6698 25401
rect 6642 25327 6698 25336
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 6564 24954 6592 25094
rect 6656 24954 6684 25327
rect 6552 24948 6604 24954
rect 6552 24890 6604 24896
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6472 24806 6684 24834
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 6366 24304 6422 24313
rect 6276 24268 6328 24274
rect 6472 24274 6500 24686
rect 6656 24449 6684 24806
rect 6642 24440 6698 24449
rect 6642 24375 6698 24384
rect 6656 24274 6684 24375
rect 6366 24239 6422 24248
rect 6460 24268 6512 24274
rect 6276 24210 6328 24216
rect 6274 24168 6330 24177
rect 6274 24103 6330 24112
rect 6288 23730 6316 24103
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6104 22066 6224 22094
rect 5998 21448 6054 21457
rect 5998 21383 6054 21392
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 6012 19417 6040 21286
rect 5998 19408 6054 19417
rect 5998 19343 6054 19352
rect 6104 18698 6132 22066
rect 6184 21956 6236 21962
rect 6288 21944 6316 23666
rect 6380 23089 6408 24239
rect 6460 24210 6512 24216
rect 6552 24268 6604 24274
rect 6552 24210 6604 24216
rect 6644 24268 6696 24274
rect 6644 24210 6696 24216
rect 6366 23080 6422 23089
rect 6366 23015 6422 23024
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6236 21916 6316 21944
rect 6184 21898 6236 21904
rect 6196 19378 6224 21898
rect 6276 21344 6328 21350
rect 6276 21286 6328 21292
rect 6288 21078 6316 21286
rect 6276 21072 6328 21078
rect 6276 21014 6328 21020
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6288 20398 6316 20878
rect 6380 20806 6408 22510
rect 6368 20800 6420 20806
rect 6368 20742 6420 20748
rect 6276 20392 6328 20398
rect 6276 20334 6328 20340
rect 6274 20088 6330 20097
rect 6274 20023 6330 20032
rect 6368 20052 6420 20058
rect 6288 19990 6316 20023
rect 6368 19994 6420 20000
rect 6276 19984 6328 19990
rect 6276 19926 6328 19932
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6196 18766 6224 19314
rect 6288 19009 6316 19790
rect 6274 19000 6330 19009
rect 6274 18935 6330 18944
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6092 18692 6144 18698
rect 6092 18634 6144 18640
rect 5998 18184 6054 18193
rect 5998 18119 6054 18128
rect 6012 17746 6040 18119
rect 6104 18057 6132 18634
rect 6184 18420 6236 18426
rect 6184 18362 6236 18368
rect 6090 18048 6146 18057
rect 6090 17983 6146 17992
rect 6090 17912 6146 17921
rect 6090 17847 6146 17856
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 6104 17678 6132 17847
rect 6092 17672 6144 17678
rect 5998 17640 6054 17649
rect 6092 17614 6144 17620
rect 5998 17575 6054 17584
rect 5724 17128 5776 17134
rect 5908 17128 5960 17134
rect 5724 17070 5776 17076
rect 5828 17088 5908 17116
rect 5644 16952 5764 16980
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 15162 5580 15370
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5552 14482 5580 14894
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5460 14334 5580 14362
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5262 12472 5318 12481
rect 5262 12407 5318 12416
rect 5460 12434 5488 14214
rect 5552 13512 5580 14334
rect 5644 13870 5672 16662
rect 5736 16522 5764 16952
rect 5828 16794 5856 17088
rect 5908 17070 5960 17076
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5736 15978 5764 16458
rect 5828 16046 5856 16730
rect 5920 16590 5948 16934
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 15162 5856 15846
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5920 15008 5948 16050
rect 6012 15638 6040 17575
rect 6104 16697 6132 17614
rect 6090 16688 6146 16697
rect 6090 16623 6146 16632
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6000 15632 6052 15638
rect 6000 15574 6052 15580
rect 6104 15570 6132 16390
rect 6196 15706 6224 18362
rect 6288 17882 6316 18935
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6288 17338 6316 17614
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6288 16046 6316 17274
rect 6380 17105 6408 19994
rect 6472 19786 6500 24210
rect 6564 23866 6592 24210
rect 6656 24070 6684 24210
rect 6748 24177 6776 27231
rect 6840 27062 6868 27474
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 26246 6868 26862
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6840 25430 6868 25978
rect 6828 25424 6880 25430
rect 6828 25366 6880 25372
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6734 24168 6790 24177
rect 6734 24103 6790 24112
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6564 23254 6592 23802
rect 6734 23760 6790 23769
rect 6644 23724 6696 23730
rect 6696 23704 6734 23712
rect 6696 23695 6790 23704
rect 6696 23684 6776 23695
rect 6644 23666 6696 23672
rect 6840 23338 6868 25230
rect 6748 23310 6868 23338
rect 6552 23248 6604 23254
rect 6552 23190 6604 23196
rect 6644 23044 6696 23050
rect 6644 22986 6696 22992
rect 6656 22710 6684 22986
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6748 22574 6776 23310
rect 6932 23225 6960 27639
rect 7012 27610 7064 27616
rect 7024 27538 7052 27610
rect 7012 27532 7064 27538
rect 7012 27474 7064 27480
rect 7116 27334 7144 27950
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 7012 27328 7064 27334
rect 7012 27270 7064 27276
rect 7104 27328 7156 27334
rect 7208 27305 7236 27814
rect 7300 27538 7328 27814
rect 7288 27532 7340 27538
rect 7288 27474 7340 27480
rect 7104 27270 7156 27276
rect 7194 27296 7250 27305
rect 7024 26994 7052 27270
rect 7012 26988 7064 26994
rect 7012 26930 7064 26936
rect 7116 26926 7144 27270
rect 7194 27231 7250 27240
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7196 27056 7248 27062
rect 7196 26998 7248 27004
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 7104 26376 7156 26382
rect 7104 26318 7156 26324
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 7024 25770 7052 26182
rect 7116 25838 7144 26318
rect 7104 25832 7156 25838
rect 7104 25774 7156 25780
rect 7012 25764 7064 25770
rect 7012 25706 7064 25712
rect 7024 25673 7052 25706
rect 7010 25664 7066 25673
rect 7010 25599 7066 25608
rect 7116 25498 7144 25774
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 7024 25226 7052 25298
rect 7012 25220 7064 25226
rect 7012 25162 7064 25168
rect 7208 25158 7236 26998
rect 7300 26382 7328 27066
rect 7392 26926 7420 29582
rect 7576 29578 7604 30359
rect 7668 29850 7696 30602
rect 7656 29844 7708 29850
rect 7656 29786 7708 29792
rect 7760 29714 7788 33798
rect 7852 32434 7880 34342
rect 7944 34241 7972 34886
rect 8024 34468 8076 34474
rect 8024 34410 8076 34416
rect 7930 34232 7986 34241
rect 7930 34167 7986 34176
rect 8036 33998 8064 34410
rect 8128 34066 8156 35006
rect 8220 34649 8248 35498
rect 8312 35193 8340 35527
rect 8298 35184 8354 35193
rect 8298 35119 8354 35128
rect 8206 34640 8262 34649
rect 8206 34575 8262 34584
rect 8208 34536 8260 34542
rect 8208 34478 8260 34484
rect 8116 34060 8168 34066
rect 8116 34002 8168 34008
rect 8024 33992 8076 33998
rect 8024 33934 8076 33940
rect 7932 33652 7984 33658
rect 7932 33594 7984 33600
rect 7944 33454 7972 33594
rect 7932 33448 7984 33454
rect 7932 33390 7984 33396
rect 7944 33114 7972 33390
rect 7932 33108 7984 33114
rect 7932 33050 7984 33056
rect 7944 32842 7972 33050
rect 7932 32836 7984 32842
rect 7932 32778 7984 32784
rect 7944 32570 7972 32778
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 7840 32428 7892 32434
rect 7840 32370 7892 32376
rect 7840 32292 7892 32298
rect 7840 32234 7892 32240
rect 7852 32201 7880 32234
rect 7932 32224 7984 32230
rect 7838 32192 7894 32201
rect 7932 32166 7984 32172
rect 7838 32127 7894 32136
rect 7944 32026 7972 32166
rect 7932 32020 7984 32026
rect 7852 31980 7932 32008
rect 7852 31249 7880 31980
rect 7932 31962 7984 31968
rect 7930 31920 7986 31929
rect 7930 31855 7986 31864
rect 7944 31822 7972 31855
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 7838 31240 7894 31249
rect 7838 31175 7894 31184
rect 7840 31136 7892 31142
rect 7840 31078 7892 31084
rect 7852 30938 7880 31078
rect 7840 30932 7892 30938
rect 7840 30874 7892 30880
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7852 30666 7880 30738
rect 7840 30660 7892 30666
rect 7840 30602 7892 30608
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7852 30190 7880 30330
rect 7944 30258 7972 31622
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7840 30184 7892 30190
rect 7840 30126 7892 30132
rect 7748 29708 7800 29714
rect 7748 29650 7800 29656
rect 7852 29578 7880 30126
rect 7932 29708 7984 29714
rect 7932 29650 7984 29656
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7840 29572 7892 29578
rect 7840 29514 7892 29520
rect 7472 28960 7524 28966
rect 7472 28902 7524 28908
rect 7564 28960 7616 28966
rect 7564 28902 7616 28908
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7484 28626 7512 28902
rect 7576 28762 7604 28902
rect 7564 28756 7616 28762
rect 7564 28698 7616 28704
rect 7748 28688 7800 28694
rect 7668 28648 7748 28676
rect 7472 28620 7524 28626
rect 7472 28562 7524 28568
rect 7564 27464 7616 27470
rect 7564 27406 7616 27412
rect 7576 27130 7604 27406
rect 7564 27124 7616 27130
rect 7564 27066 7616 27072
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7472 26920 7524 26926
rect 7472 26862 7524 26868
rect 7378 26616 7434 26625
rect 7378 26551 7380 26560
rect 7432 26551 7434 26560
rect 7380 26522 7432 26528
rect 7288 26376 7340 26382
rect 7288 26318 7340 26324
rect 7288 26240 7340 26246
rect 7288 26182 7340 26188
rect 7300 25974 7328 26182
rect 7288 25968 7340 25974
rect 7288 25910 7340 25916
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 7392 24954 7420 25230
rect 7380 24948 7432 24954
rect 7380 24890 7432 24896
rect 7102 24848 7158 24857
rect 7012 24812 7064 24818
rect 7484 24834 7512 26862
rect 7564 26852 7616 26858
rect 7564 26794 7616 26800
rect 7576 25158 7604 26794
rect 7668 26314 7696 28648
rect 7748 28630 7800 28636
rect 7852 28626 7880 28902
rect 7840 28620 7892 28626
rect 7840 28562 7892 28568
rect 7840 28484 7892 28490
rect 7840 28426 7892 28432
rect 7852 28218 7880 28426
rect 7944 28370 7972 29650
rect 8036 29034 8064 33934
rect 8116 32972 8168 32978
rect 8116 32914 8168 32920
rect 8128 32026 8156 32914
rect 8220 32026 8248 34478
rect 8312 32609 8340 35119
rect 8404 34105 8432 35770
rect 8576 35556 8628 35562
rect 8576 35498 8628 35504
rect 8484 35148 8536 35154
rect 8484 35090 8536 35096
rect 8390 34096 8446 34105
rect 8390 34031 8392 34040
rect 8444 34031 8446 34040
rect 8392 34002 8444 34008
rect 8496 33930 8524 35090
rect 8588 34785 8616 35498
rect 8680 35494 8708 35799
rect 8772 35630 8800 36094
rect 8852 36032 8904 36038
rect 9048 36020 9076 36094
rect 8852 35974 8904 35980
rect 8956 35992 9076 36020
rect 9128 36032 9180 36038
rect 8760 35624 8812 35630
rect 8760 35566 8812 35572
rect 8864 35562 8892 35974
rect 8852 35556 8904 35562
rect 8852 35498 8904 35504
rect 8668 35488 8720 35494
rect 8668 35430 8720 35436
rect 8852 35012 8904 35018
rect 8852 34954 8904 34960
rect 8574 34776 8630 34785
rect 8574 34711 8630 34720
rect 8758 34640 8814 34649
rect 8864 34610 8892 34954
rect 8758 34575 8814 34584
rect 8852 34604 8904 34610
rect 8772 34542 8800 34575
rect 8852 34546 8904 34552
rect 8956 34542 8984 35992
rect 9128 35974 9180 35980
rect 9034 35864 9090 35873
rect 9034 35799 9090 35808
rect 9048 34542 9076 35799
rect 9140 35737 9168 35974
rect 9126 35728 9182 35737
rect 9126 35663 9182 35672
rect 9128 35624 9180 35630
rect 9128 35566 9180 35572
rect 9140 35465 9168 35566
rect 9126 35456 9182 35465
rect 9126 35391 9182 35400
rect 8760 34536 8812 34542
rect 8760 34478 8812 34484
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 9036 34536 9088 34542
rect 9036 34478 9088 34484
rect 8484 33924 8536 33930
rect 8484 33866 8536 33872
rect 8392 33448 8444 33454
rect 8392 33390 8444 33396
rect 8404 32774 8432 33390
rect 8484 33380 8536 33386
rect 8484 33322 8536 33328
rect 8496 33114 8524 33322
rect 8668 33312 8720 33318
rect 8668 33254 8720 33260
rect 8484 33108 8536 33114
rect 8484 33050 8536 33056
rect 8680 32978 8708 33254
rect 8772 33130 8800 34478
rect 9048 34134 9076 34478
rect 9036 34128 9088 34134
rect 9036 34070 9088 34076
rect 9034 33552 9090 33561
rect 9034 33487 9090 33496
rect 8772 33102 8892 33130
rect 8668 32972 8720 32978
rect 8668 32914 8720 32920
rect 8760 32972 8812 32978
rect 8760 32914 8812 32920
rect 8392 32768 8444 32774
rect 8392 32710 8444 32716
rect 8298 32600 8354 32609
rect 8298 32535 8354 32544
rect 8300 32496 8352 32502
rect 8300 32438 8352 32444
rect 8576 32496 8628 32502
rect 8576 32438 8628 32444
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 8208 32020 8260 32026
rect 8208 31962 8260 31968
rect 8128 31278 8156 31962
rect 8312 31890 8340 32438
rect 8390 32056 8446 32065
rect 8588 32026 8616 32438
rect 8390 31991 8446 32000
rect 8484 32020 8536 32026
rect 8404 31958 8432 31991
rect 8484 31962 8536 31968
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8392 31952 8444 31958
rect 8392 31894 8444 31900
rect 8300 31884 8352 31890
rect 8300 31826 8352 31832
rect 8208 31680 8260 31686
rect 8208 31622 8260 31628
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8116 31272 8168 31278
rect 8116 31214 8168 31220
rect 8128 30802 8156 31214
rect 8220 30802 8248 31622
rect 8312 31210 8340 31622
rect 8300 31204 8352 31210
rect 8300 31146 8352 31152
rect 8116 30796 8168 30802
rect 8116 30738 8168 30744
rect 8208 30796 8260 30802
rect 8208 30738 8260 30744
rect 8312 30598 8340 31146
rect 8300 30592 8352 30598
rect 8300 30534 8352 30540
rect 8114 30288 8170 30297
rect 8114 30223 8170 30232
rect 8128 30190 8156 30223
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 8128 29850 8156 30126
rect 8312 30122 8340 30534
rect 8300 30116 8352 30122
rect 8300 30058 8352 30064
rect 8116 29844 8168 29850
rect 8116 29786 8168 29792
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8024 29028 8076 29034
rect 8024 28970 8076 28976
rect 8128 28506 8156 29650
rect 8208 29504 8260 29510
rect 8208 29446 8260 29452
rect 8220 28966 8248 29446
rect 8208 28960 8260 28966
rect 8208 28902 8260 28908
rect 8220 28626 8248 28902
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 8128 28478 8340 28506
rect 7944 28342 8156 28370
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7932 28212 7984 28218
rect 7932 28154 7984 28160
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7748 27464 7800 27470
rect 7748 27406 7800 27412
rect 7760 27130 7788 27406
rect 7748 27124 7800 27130
rect 7748 27066 7800 27072
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7760 26450 7788 26930
rect 7748 26444 7800 26450
rect 7748 26386 7800 26392
rect 7656 26308 7708 26314
rect 7656 26250 7708 26256
rect 7748 26308 7800 26314
rect 7852 26296 7880 28018
rect 7944 27946 7972 28154
rect 7932 27940 7984 27946
rect 7932 27882 7984 27888
rect 8024 27940 8076 27946
rect 8024 27882 8076 27888
rect 8036 27033 8064 27882
rect 8128 27538 8156 28342
rect 8312 28014 8340 28478
rect 8404 28121 8432 31894
rect 8496 30190 8524 31962
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8588 30938 8616 31826
rect 8576 30932 8628 30938
rect 8576 30874 8628 30880
rect 8680 30870 8708 32914
rect 8772 32609 8800 32914
rect 8758 32600 8814 32609
rect 8758 32535 8814 32544
rect 8772 32502 8800 32535
rect 8760 32496 8812 32502
rect 8760 32438 8812 32444
rect 8864 32065 8892 33102
rect 8944 32768 8996 32774
rect 8942 32736 8944 32745
rect 8996 32736 8998 32745
rect 8942 32671 8998 32680
rect 8944 32428 8996 32434
rect 8944 32370 8996 32376
rect 8850 32056 8906 32065
rect 8772 32014 8850 32042
rect 8772 31958 8800 32014
rect 8850 31991 8906 32000
rect 8956 31958 8984 32370
rect 8760 31952 8812 31958
rect 8944 31952 8996 31958
rect 8760 31894 8812 31900
rect 8864 31912 8944 31940
rect 8760 31748 8812 31754
rect 8760 31690 8812 31696
rect 8668 30864 8720 30870
rect 8668 30806 8720 30812
rect 8668 30728 8720 30734
rect 8668 30670 8720 30676
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 8496 29714 8524 30126
rect 8484 29708 8536 29714
rect 8484 29650 8536 29656
rect 8680 29560 8708 30670
rect 8772 30326 8800 31690
rect 8864 30870 8892 31912
rect 8944 31894 8996 31900
rect 8944 31816 8996 31822
rect 8944 31758 8996 31764
rect 8956 31482 8984 31758
rect 8944 31476 8996 31482
rect 8944 31418 8996 31424
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 8852 30864 8904 30870
rect 8852 30806 8904 30812
rect 8956 30666 8984 31146
rect 8944 30660 8996 30666
rect 8944 30602 8996 30608
rect 8850 30560 8906 30569
rect 8850 30495 8906 30504
rect 8760 30320 8812 30326
rect 8760 30262 8812 30268
rect 8864 30190 8892 30495
rect 8852 30184 8904 30190
rect 8944 30184 8996 30190
rect 8852 30126 8904 30132
rect 8942 30152 8944 30161
rect 8996 30152 8998 30161
rect 8942 30087 8998 30096
rect 8852 30048 8904 30054
rect 8850 30016 8852 30025
rect 8904 30016 8906 30025
rect 8850 29951 8906 29960
rect 8680 29532 8800 29560
rect 8772 29306 8800 29532
rect 8760 29300 8812 29306
rect 8760 29242 8812 29248
rect 8484 29232 8536 29238
rect 8484 29174 8536 29180
rect 8496 28966 8524 29174
rect 8772 29102 8800 29242
rect 8668 29096 8720 29102
rect 8668 29038 8720 29044
rect 8760 29096 8812 29102
rect 8864 29073 8892 29951
rect 8956 29782 8984 30087
rect 8944 29776 8996 29782
rect 8944 29718 8996 29724
rect 9048 29170 9076 33487
rect 9126 33008 9182 33017
rect 9126 32943 9182 32952
rect 9140 32842 9168 32943
rect 9128 32836 9180 32842
rect 9128 32778 9180 32784
rect 9140 32298 9168 32778
rect 9128 32292 9180 32298
rect 9128 32234 9180 32240
rect 9128 31884 9180 31890
rect 9128 31826 9180 31832
rect 9140 31278 9168 31826
rect 9128 31272 9180 31278
rect 9128 31214 9180 31220
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9140 30802 9168 31078
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 9232 30190 9260 36751
rect 9324 36174 9352 37674
rect 9508 37312 9536 37726
rect 9600 37466 9628 37742
rect 9588 37460 9640 37466
rect 9588 37402 9640 37408
rect 9680 37392 9732 37398
rect 9680 37334 9732 37340
rect 9588 37324 9640 37330
rect 9508 37284 9588 37312
rect 9588 37266 9640 37272
rect 9404 37120 9456 37126
rect 9404 37062 9456 37068
rect 9416 36718 9444 37062
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9600 36632 9628 37266
rect 9692 36854 9720 37334
rect 9772 37120 9824 37126
rect 9772 37062 9824 37068
rect 9680 36848 9732 36854
rect 9680 36790 9732 36796
rect 9784 36666 9812 37062
rect 9580 36604 9628 36632
rect 9692 36638 9812 36666
rect 9876 36666 9904 38354
rect 9968 36768 9996 38950
rect 10060 38418 10088 38966
rect 10230 38927 10286 38936
rect 10138 38856 10194 38865
rect 10138 38791 10194 38800
rect 10152 38758 10180 38791
rect 10140 38752 10192 38758
rect 10140 38694 10192 38700
rect 10244 38554 10272 38927
rect 10324 38888 10376 38894
rect 10428 38865 10456 39986
rect 10324 38830 10376 38836
rect 10414 38856 10470 38865
rect 10232 38548 10284 38554
rect 10232 38490 10284 38496
rect 10048 38412 10100 38418
rect 10048 38354 10100 38360
rect 10336 38196 10364 38830
rect 10414 38791 10470 38800
rect 10416 38752 10468 38758
rect 10416 38694 10468 38700
rect 10428 38486 10456 38694
rect 10520 38554 10548 40122
rect 10612 39030 10640 41024
rect 10874 41032 10930 41041
rect 10968 41006 11020 41012
rect 10874 40967 10930 40976
rect 10722 40828 11030 40837
rect 10722 40826 10728 40828
rect 10784 40826 10808 40828
rect 10864 40826 10888 40828
rect 10944 40826 10968 40828
rect 11024 40826 11030 40828
rect 10784 40774 10786 40826
rect 10966 40774 10968 40826
rect 10722 40772 10728 40774
rect 10784 40772 10808 40774
rect 10864 40772 10888 40774
rect 10944 40772 10968 40774
rect 11024 40772 11030 40774
rect 10722 40763 11030 40772
rect 10692 40452 10744 40458
rect 10692 40394 10744 40400
rect 10704 40225 10732 40394
rect 10690 40216 10746 40225
rect 10690 40151 10692 40160
rect 10744 40151 10746 40160
rect 10692 40122 10744 40128
rect 11072 40118 11100 41550
rect 11164 41070 11192 42706
rect 11244 42628 11296 42634
rect 11244 42570 11296 42576
rect 11152 41064 11204 41070
rect 11152 41006 11204 41012
rect 11152 40928 11204 40934
rect 11152 40870 11204 40876
rect 11060 40112 11112 40118
rect 11164 40089 11192 40870
rect 11256 40458 11284 42570
rect 11520 42084 11572 42090
rect 11520 42026 11572 42032
rect 11532 41614 11560 42026
rect 11520 41608 11572 41614
rect 11572 41556 11652 41562
rect 11520 41550 11652 41556
rect 11532 41534 11652 41550
rect 11520 41472 11572 41478
rect 11520 41414 11572 41420
rect 11532 41274 11560 41414
rect 11520 41268 11572 41274
rect 11520 41210 11572 41216
rect 11520 40724 11572 40730
rect 11520 40666 11572 40672
rect 11428 40588 11480 40594
rect 11428 40530 11480 40536
rect 11336 40520 11388 40526
rect 11336 40462 11388 40468
rect 11244 40452 11296 40458
rect 11244 40394 11296 40400
rect 11060 40054 11112 40060
rect 11150 40080 11206 40089
rect 11150 40015 11206 40024
rect 11244 40044 11296 40050
rect 11348 40032 11376 40462
rect 11440 40089 11468 40530
rect 11296 40004 11376 40032
rect 11426 40080 11482 40089
rect 11426 40015 11482 40024
rect 11244 39986 11296 39992
rect 10874 39944 10930 39953
rect 10874 39879 10930 39888
rect 11060 39908 11112 39914
rect 10888 39846 10916 39879
rect 11060 39850 11112 39856
rect 10876 39840 10928 39846
rect 10876 39782 10928 39788
rect 10722 39740 11030 39749
rect 10722 39738 10728 39740
rect 10784 39738 10808 39740
rect 10864 39738 10888 39740
rect 10944 39738 10968 39740
rect 11024 39738 11030 39740
rect 10784 39686 10786 39738
rect 10966 39686 10968 39738
rect 10722 39684 10728 39686
rect 10784 39684 10808 39686
rect 10864 39684 10888 39686
rect 10944 39684 10968 39686
rect 11024 39684 11030 39686
rect 10722 39675 11030 39684
rect 10690 39536 10746 39545
rect 10690 39471 10746 39480
rect 10704 39370 10732 39471
rect 10692 39364 10744 39370
rect 10692 39306 10744 39312
rect 10968 39296 11020 39302
rect 10968 39238 11020 39244
rect 10980 39098 11008 39238
rect 10968 39092 11020 39098
rect 10968 39034 11020 39040
rect 10600 39024 10652 39030
rect 10600 38966 10652 38972
rect 10722 38652 11030 38661
rect 10722 38650 10728 38652
rect 10784 38650 10808 38652
rect 10864 38650 10888 38652
rect 10944 38650 10968 38652
rect 11024 38650 11030 38652
rect 10784 38598 10786 38650
rect 10966 38598 10968 38650
rect 10722 38596 10728 38598
rect 10784 38596 10808 38598
rect 10864 38596 10888 38598
rect 10944 38596 10968 38598
rect 11024 38596 11030 38598
rect 10722 38587 11030 38596
rect 10508 38548 10560 38554
rect 10508 38490 10560 38496
rect 10416 38480 10468 38486
rect 10416 38422 10468 38428
rect 10600 38480 10652 38486
rect 10968 38480 11020 38486
rect 10600 38422 10652 38428
rect 10966 38448 10968 38457
rect 11020 38448 11022 38457
rect 10508 38208 10560 38214
rect 10336 38168 10456 38196
rect 10062 38108 10370 38117
rect 10062 38106 10068 38108
rect 10124 38106 10148 38108
rect 10204 38106 10228 38108
rect 10284 38106 10308 38108
rect 10364 38106 10370 38108
rect 10124 38054 10126 38106
rect 10306 38054 10308 38106
rect 10062 38052 10068 38054
rect 10124 38052 10148 38054
rect 10204 38052 10228 38054
rect 10284 38052 10308 38054
rect 10364 38052 10370 38054
rect 10062 38043 10370 38052
rect 10428 37992 10456 38168
rect 10508 38150 10560 38156
rect 10336 37964 10456 37992
rect 10336 37330 10364 37964
rect 10416 37664 10468 37670
rect 10416 37606 10468 37612
rect 10324 37324 10376 37330
rect 10324 37266 10376 37272
rect 10062 37020 10370 37029
rect 10062 37018 10068 37020
rect 10124 37018 10148 37020
rect 10204 37018 10228 37020
rect 10284 37018 10308 37020
rect 10364 37018 10370 37020
rect 10124 36966 10126 37018
rect 10306 36966 10308 37018
rect 10062 36964 10068 36966
rect 10124 36964 10148 36966
rect 10204 36964 10228 36966
rect 10284 36964 10308 36966
rect 10364 36964 10370 36966
rect 10062 36955 10370 36964
rect 10322 36816 10378 36825
rect 9968 36740 10272 36768
rect 10322 36751 10324 36760
rect 10138 36680 10194 36689
rect 9876 36638 10088 36666
rect 9404 36576 9456 36582
rect 9404 36518 9456 36524
rect 9496 36576 9548 36582
rect 9496 36518 9548 36524
rect 9416 36417 9444 36518
rect 9402 36408 9458 36417
rect 9402 36343 9458 36352
rect 9404 36236 9456 36242
rect 9404 36178 9456 36184
rect 9312 36168 9364 36174
rect 9312 36110 9364 36116
rect 9324 35766 9352 36110
rect 9312 35760 9364 35766
rect 9312 35702 9364 35708
rect 9312 35488 9364 35494
rect 9312 35430 9364 35436
rect 9324 35154 9352 35430
rect 9416 35154 9444 36178
rect 9508 35630 9536 36518
rect 9580 36394 9608 36604
rect 9580 36366 9628 36394
rect 9496 35624 9548 35630
rect 9600 35601 9628 36366
rect 9692 36174 9720 36638
rect 9772 36576 9824 36582
rect 9770 36544 9772 36553
rect 9864 36576 9916 36582
rect 9824 36544 9826 36553
rect 9864 36518 9916 36524
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 9770 36479 9826 36488
rect 9770 36272 9826 36281
rect 9770 36207 9826 36216
rect 9680 36168 9732 36174
rect 9680 36110 9732 36116
rect 9678 36000 9734 36009
rect 9678 35935 9734 35944
rect 9692 35834 9720 35935
rect 9680 35828 9732 35834
rect 9680 35770 9732 35776
rect 9680 35624 9732 35630
rect 9496 35566 9548 35572
rect 9586 35592 9642 35601
rect 9508 35290 9536 35566
rect 9784 35612 9812 36207
rect 9876 35630 9904 36518
rect 9968 35834 9996 36518
rect 10060 36174 10088 36638
rect 10138 36615 10194 36624
rect 10152 36242 10180 36615
rect 10244 36310 10272 36740
rect 10376 36751 10378 36760
rect 10324 36722 10376 36728
rect 10428 36718 10456 37606
rect 10416 36712 10468 36718
rect 10416 36654 10468 36660
rect 10416 36576 10468 36582
rect 10416 36518 10468 36524
rect 10428 36378 10456 36518
rect 10324 36372 10376 36378
rect 10324 36314 10376 36320
rect 10416 36372 10468 36378
rect 10416 36314 10468 36320
rect 10232 36304 10284 36310
rect 10232 36246 10284 36252
rect 10140 36236 10192 36242
rect 10140 36178 10192 36184
rect 10048 36168 10100 36174
rect 10048 36110 10100 36116
rect 10138 36136 10194 36145
rect 10138 36071 10140 36080
rect 10192 36071 10194 36080
rect 10140 36042 10192 36048
rect 10336 36038 10364 36314
rect 10416 36236 10468 36242
rect 10416 36178 10468 36184
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10062 35932 10370 35941
rect 10062 35930 10068 35932
rect 10124 35930 10148 35932
rect 10204 35930 10228 35932
rect 10284 35930 10308 35932
rect 10364 35930 10370 35932
rect 10124 35878 10126 35930
rect 10306 35878 10308 35930
rect 10062 35876 10068 35878
rect 10124 35876 10148 35878
rect 10204 35876 10228 35878
rect 10284 35876 10308 35878
rect 10364 35876 10370 35878
rect 10062 35867 10370 35876
rect 10428 35834 10456 36178
rect 10520 36038 10548 38150
rect 10612 37913 10640 38422
rect 10966 38383 11022 38392
rect 10692 38276 10744 38282
rect 10692 38218 10744 38224
rect 10598 37904 10654 37913
rect 10598 37839 10654 37848
rect 10704 37652 10732 38218
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 10796 37874 10824 38150
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 10612 37624 10732 37652
rect 10612 36904 10640 37624
rect 10722 37564 11030 37573
rect 10722 37562 10728 37564
rect 10784 37562 10808 37564
rect 10864 37562 10888 37564
rect 10944 37562 10968 37564
rect 11024 37562 11030 37564
rect 10784 37510 10786 37562
rect 10966 37510 10968 37562
rect 10722 37508 10728 37510
rect 10784 37508 10808 37510
rect 10864 37508 10888 37510
rect 10944 37508 10968 37510
rect 11024 37508 11030 37510
rect 10722 37499 11030 37508
rect 10876 37460 10928 37466
rect 10876 37402 10928 37408
rect 10612 36876 10732 36904
rect 10600 36780 10652 36786
rect 10600 36722 10652 36728
rect 10508 36032 10560 36038
rect 10508 35974 10560 35980
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 10416 35828 10468 35834
rect 10416 35770 10468 35776
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 10324 35692 10376 35698
rect 10324 35634 10376 35640
rect 9732 35584 9812 35612
rect 9864 35624 9916 35630
rect 9680 35566 9732 35572
rect 9864 35566 9916 35572
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 9586 35527 9642 35536
rect 9876 35476 9904 35566
rect 10048 35556 10100 35562
rect 10048 35498 10100 35504
rect 9600 35448 9904 35476
rect 9496 35284 9548 35290
rect 9496 35226 9548 35232
rect 9312 35148 9364 35154
rect 9312 35090 9364 35096
rect 9404 35148 9456 35154
rect 9404 35090 9456 35096
rect 9312 34944 9364 34950
rect 9312 34886 9364 34892
rect 9324 33114 9352 34886
rect 9416 34592 9444 35090
rect 9416 34564 9536 34592
rect 9508 34474 9536 34564
rect 9404 34468 9456 34474
rect 9404 34410 9456 34416
rect 9496 34468 9548 34474
rect 9496 34410 9548 34416
rect 9416 33930 9444 34410
rect 9600 34066 9628 35448
rect 9680 35284 9732 35290
rect 9680 35226 9732 35232
rect 9692 35086 9720 35226
rect 9956 35216 10008 35222
rect 10060 35193 10088 35498
rect 10152 35222 10180 35566
rect 10140 35216 10192 35222
rect 9956 35158 10008 35164
rect 10046 35184 10102 35193
rect 9680 35080 9732 35086
rect 9864 35080 9916 35086
rect 9680 35022 9732 35028
rect 9784 35040 9864 35068
rect 9784 34542 9812 35040
rect 9864 35022 9916 35028
rect 9864 34944 9916 34950
rect 9864 34886 9916 34892
rect 9772 34536 9824 34542
rect 9772 34478 9824 34484
rect 9680 34400 9732 34406
rect 9680 34342 9732 34348
rect 9692 34202 9720 34342
rect 9680 34196 9732 34202
rect 9680 34138 9732 34144
rect 9678 34096 9734 34105
rect 9496 34060 9548 34066
rect 9496 34002 9548 34008
rect 9588 34060 9640 34066
rect 9784 34066 9812 34478
rect 9876 34066 9904 34886
rect 9968 34474 9996 35158
rect 10140 35158 10192 35164
rect 10046 35119 10102 35128
rect 10244 34932 10272 35634
rect 10336 35601 10364 35634
rect 10322 35592 10378 35601
rect 10322 35527 10378 35536
rect 10428 35465 10456 35770
rect 10520 35562 10548 35974
rect 10612 35737 10640 36722
rect 10704 36689 10732 36876
rect 10888 36786 10916 37402
rect 10876 36780 10928 36786
rect 10876 36722 10928 36728
rect 10690 36680 10746 36689
rect 10690 36615 10746 36624
rect 10722 36476 11030 36485
rect 10722 36474 10728 36476
rect 10784 36474 10808 36476
rect 10864 36474 10888 36476
rect 10944 36474 10968 36476
rect 11024 36474 11030 36476
rect 10784 36422 10786 36474
rect 10966 36422 10968 36474
rect 10722 36420 10728 36422
rect 10784 36420 10808 36422
rect 10864 36420 10888 36422
rect 10944 36420 10968 36422
rect 11024 36420 11030 36422
rect 10722 36411 11030 36420
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10598 35728 10654 35737
rect 10598 35663 10654 35672
rect 10612 35630 10640 35663
rect 10600 35624 10652 35630
rect 10600 35566 10652 35572
rect 10508 35556 10560 35562
rect 10508 35498 10560 35504
rect 10704 35476 10732 36314
rect 10966 36272 11022 36281
rect 10966 36207 11022 36216
rect 10980 36174 11008 36207
rect 10968 36168 11020 36174
rect 10874 36136 10930 36145
rect 10968 36110 11020 36116
rect 10874 36071 10930 36080
rect 10888 35766 10916 36071
rect 10876 35760 10928 35766
rect 10876 35702 10928 35708
rect 10888 35494 10916 35702
rect 10414 35456 10470 35465
rect 10414 35391 10470 35400
rect 10612 35448 10732 35476
rect 10876 35488 10928 35494
rect 10428 35222 10456 35391
rect 10416 35216 10468 35222
rect 10416 35158 10468 35164
rect 10244 34904 10456 34932
rect 10062 34844 10370 34853
rect 10062 34842 10068 34844
rect 10124 34842 10148 34844
rect 10204 34842 10228 34844
rect 10284 34842 10308 34844
rect 10364 34842 10370 34844
rect 10124 34790 10126 34842
rect 10306 34790 10308 34842
rect 10062 34788 10068 34790
rect 10124 34788 10148 34790
rect 10204 34788 10228 34790
rect 10284 34788 10308 34790
rect 10364 34788 10370 34790
rect 10062 34779 10370 34788
rect 10140 34740 10192 34746
rect 10428 34728 10456 34904
rect 10140 34682 10192 34688
rect 10336 34700 10456 34728
rect 9956 34468 10008 34474
rect 9956 34410 10008 34416
rect 10048 34128 10100 34134
rect 10046 34096 10048 34105
rect 10100 34096 10102 34105
rect 9678 34031 9680 34040
rect 9588 34002 9640 34008
rect 9732 34031 9734 34040
rect 9772 34060 9824 34066
rect 9680 34002 9732 34008
rect 9772 34002 9824 34008
rect 9864 34060 9916 34066
rect 10046 34031 10102 34040
rect 9864 34002 9916 34008
rect 9404 33924 9456 33930
rect 9404 33866 9456 33872
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9508 32774 9536 34002
rect 9678 33960 9734 33969
rect 10152 33930 10180 34682
rect 10336 33946 10364 34700
rect 10508 34672 10560 34678
rect 10508 34614 10560 34620
rect 10520 34598 10557 34614
rect 10416 34468 10468 34474
rect 10416 34410 10468 34416
rect 10428 34066 10456 34410
rect 10416 34060 10468 34066
rect 10416 34002 10468 34008
rect 9678 33895 9734 33904
rect 10140 33924 10192 33930
rect 9692 33386 9720 33895
rect 10336 33918 10456 33946
rect 10140 33866 10192 33872
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9680 33380 9732 33386
rect 9680 33322 9732 33328
rect 9772 33108 9824 33114
rect 9772 33050 9824 33056
rect 9588 32972 9640 32978
rect 9588 32914 9640 32920
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 9496 32768 9548 32774
rect 9496 32710 9548 32716
rect 9324 31521 9352 32710
rect 9404 32496 9456 32502
rect 9404 32438 9456 32444
rect 9416 31890 9444 32438
rect 9508 32026 9536 32710
rect 9600 32570 9628 32914
rect 9588 32564 9640 32570
rect 9588 32506 9640 32512
rect 9680 32496 9732 32502
rect 9678 32464 9680 32473
rect 9732 32464 9734 32473
rect 9678 32399 9734 32408
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9692 32201 9720 32302
rect 9678 32192 9734 32201
rect 9784 32178 9812 33050
rect 9876 33046 9904 33798
rect 10062 33756 10370 33765
rect 10062 33754 10068 33756
rect 10124 33754 10148 33756
rect 10204 33754 10228 33756
rect 10284 33754 10308 33756
rect 10364 33754 10370 33756
rect 10124 33702 10126 33754
rect 10306 33702 10308 33754
rect 10062 33700 10068 33702
rect 10124 33700 10148 33702
rect 10204 33700 10228 33702
rect 10284 33700 10308 33702
rect 10364 33700 10370 33702
rect 10062 33691 10370 33700
rect 10140 33652 10192 33658
rect 10140 33594 10192 33600
rect 9956 33380 10008 33386
rect 9956 33322 10008 33328
rect 9864 33040 9916 33046
rect 9864 32982 9916 32988
rect 9862 32600 9918 32609
rect 9862 32535 9918 32544
rect 9876 32434 9904 32535
rect 9968 32484 9996 33322
rect 10152 32774 10180 33594
rect 10232 33380 10284 33386
rect 10232 33322 10284 33328
rect 10140 32768 10192 32774
rect 10244 32756 10272 33322
rect 10428 32994 10456 33918
rect 10520 33561 10548 34598
rect 10612 34406 10640 35448
rect 10876 35430 10928 35436
rect 10722 35388 11030 35397
rect 10722 35386 10728 35388
rect 10784 35386 10808 35388
rect 10864 35386 10888 35388
rect 10944 35386 10968 35388
rect 11024 35386 11030 35388
rect 10784 35334 10786 35386
rect 10966 35334 10968 35386
rect 10722 35332 10728 35334
rect 10784 35332 10808 35334
rect 10864 35332 10888 35334
rect 10944 35332 10968 35334
rect 11024 35332 11030 35334
rect 10722 35323 11030 35332
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10612 34082 10640 34342
rect 10722 34300 11030 34309
rect 10722 34298 10728 34300
rect 10784 34298 10808 34300
rect 10864 34298 10888 34300
rect 10944 34298 10968 34300
rect 11024 34298 11030 34300
rect 10784 34246 10786 34298
rect 10966 34246 10968 34298
rect 10722 34244 10728 34246
rect 10784 34244 10808 34246
rect 10864 34244 10888 34246
rect 10944 34244 10968 34246
rect 11024 34244 11030 34246
rect 10722 34235 11030 34244
rect 11072 34082 11100 39850
rect 11244 39840 11296 39846
rect 11244 39782 11296 39788
rect 11152 39636 11204 39642
rect 11152 39578 11204 39584
rect 11164 38554 11192 39578
rect 11256 39370 11284 39782
rect 11244 39364 11296 39370
rect 11244 39306 11296 39312
rect 11256 39001 11284 39306
rect 11242 38992 11298 39001
rect 11242 38927 11298 38936
rect 11152 38548 11204 38554
rect 11152 38490 11204 38496
rect 11244 38412 11296 38418
rect 11244 38354 11296 38360
rect 11152 38276 11204 38282
rect 11152 38218 11204 38224
rect 11164 37641 11192 38218
rect 11256 38185 11284 38354
rect 11242 38176 11298 38185
rect 11242 38111 11298 38120
rect 11244 38004 11296 38010
rect 11244 37946 11296 37952
rect 11150 37632 11206 37641
rect 11150 37567 11206 37576
rect 11152 37460 11204 37466
rect 11152 37402 11204 37408
rect 11164 37369 11192 37402
rect 11256 37398 11284 37946
rect 11244 37392 11296 37398
rect 11150 37360 11206 37369
rect 11244 37334 11296 37340
rect 11150 37295 11206 37304
rect 11244 37256 11296 37262
rect 11242 37224 11244 37233
rect 11296 37224 11298 37233
rect 11242 37159 11298 37168
rect 11152 37120 11204 37126
rect 11152 37062 11204 37068
rect 11164 36825 11192 37062
rect 11256 36922 11284 37159
rect 11244 36916 11296 36922
rect 11244 36858 11296 36864
rect 11150 36816 11206 36825
rect 11150 36751 11206 36760
rect 11152 36644 11204 36650
rect 11152 36586 11204 36592
rect 11164 36378 11192 36586
rect 11244 36576 11296 36582
rect 11244 36518 11296 36524
rect 11152 36372 11204 36378
rect 11152 36314 11204 36320
rect 11152 36100 11204 36106
rect 11152 36042 11204 36048
rect 11164 35154 11192 36042
rect 11152 35148 11204 35154
rect 11152 35090 11204 35096
rect 11150 34504 11206 34513
rect 11150 34439 11206 34448
rect 11164 34406 11192 34439
rect 11152 34400 11204 34406
rect 11152 34342 11204 34348
rect 10612 34054 10824 34082
rect 10796 33998 10824 34054
rect 10980 34054 11100 34082
rect 11164 34066 11192 34342
rect 11256 34202 11284 36518
rect 11348 34950 11376 40004
rect 11428 39364 11480 39370
rect 11428 39306 11480 39312
rect 11440 38350 11468 39306
rect 11428 38344 11480 38350
rect 11426 38312 11428 38321
rect 11480 38312 11482 38321
rect 11426 38247 11482 38256
rect 11426 38176 11482 38185
rect 11426 38111 11482 38120
rect 11440 37262 11468 38111
rect 11428 37256 11480 37262
rect 11428 37198 11480 37204
rect 11426 36952 11482 36961
rect 11426 36887 11482 36896
rect 11440 36145 11468 36887
rect 11426 36136 11482 36145
rect 11426 36071 11482 36080
rect 11532 35986 11560 40666
rect 11624 39914 11652 41534
rect 11716 40526 11744 42774
rect 12072 42764 12124 42770
rect 12072 42706 12124 42712
rect 11796 42560 11848 42566
rect 11796 42502 11848 42508
rect 11888 42560 11940 42566
rect 11888 42502 11940 42508
rect 11808 41818 11836 42502
rect 11900 41993 11928 42502
rect 11886 41984 11942 41993
rect 11886 41919 11942 41928
rect 11796 41812 11848 41818
rect 11796 41754 11848 41760
rect 12084 41414 12112 42706
rect 12164 42696 12216 42702
rect 12164 42638 12216 42644
rect 11992 41386 12112 41414
rect 11796 40996 11848 41002
rect 11796 40938 11848 40944
rect 11704 40520 11756 40526
rect 11704 40462 11756 40468
rect 11612 39908 11664 39914
rect 11612 39850 11664 39856
rect 11612 39432 11664 39438
rect 11612 39374 11664 39380
rect 11440 35958 11560 35986
rect 11440 35154 11468 35958
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11348 34082 11376 34886
rect 11440 34202 11468 35090
rect 11428 34196 11480 34202
rect 11428 34138 11480 34144
rect 11440 34105 11468 34138
rect 11152 34060 11204 34066
rect 10600 33992 10652 33998
rect 10600 33934 10652 33940
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10506 33552 10562 33561
rect 10506 33487 10562 33496
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10520 33114 10548 33390
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10428 32966 10548 32994
rect 10244 32728 10456 32756
rect 10140 32710 10192 32716
rect 10062 32668 10370 32677
rect 10062 32666 10068 32668
rect 10124 32666 10148 32668
rect 10204 32666 10228 32668
rect 10284 32666 10308 32668
rect 10364 32666 10370 32668
rect 10124 32614 10126 32666
rect 10306 32614 10308 32666
rect 10062 32612 10068 32614
rect 10124 32612 10148 32614
rect 10204 32612 10228 32614
rect 10284 32612 10308 32614
rect 10364 32612 10370 32614
rect 10062 32603 10370 32612
rect 10232 32496 10284 32502
rect 9968 32456 10180 32484
rect 9864 32428 9916 32434
rect 9864 32370 9916 32376
rect 10152 32230 10180 32456
rect 10232 32438 10284 32444
rect 10322 32464 10378 32473
rect 10244 32366 10272 32438
rect 10322 32399 10378 32408
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 10140 32224 10192 32230
rect 9784 32150 9904 32178
rect 10140 32166 10192 32172
rect 9678 32127 9734 32136
rect 9586 32056 9642 32065
rect 9496 32020 9548 32026
rect 9692 32042 9720 32127
rect 9692 32014 9812 32042
rect 9586 31991 9642 32000
rect 9496 31962 9548 31968
rect 9404 31884 9456 31890
rect 9404 31826 9456 31832
rect 9600 31754 9628 31991
rect 9508 31726 9628 31754
rect 9678 31784 9734 31793
rect 9402 31648 9458 31657
rect 9402 31583 9458 31592
rect 9310 31512 9366 31521
rect 9310 31447 9366 31456
rect 9324 30870 9352 31447
rect 9312 30864 9364 30870
rect 9312 30806 9364 30812
rect 9416 30734 9444 31583
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9416 30376 9444 30670
rect 9508 30394 9536 31726
rect 9678 31719 9734 31728
rect 9588 31204 9640 31210
rect 9588 31146 9640 31152
rect 9600 30938 9628 31146
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 9588 30660 9640 30666
rect 9588 30602 9640 30608
rect 9324 30348 9444 30376
rect 9496 30388 9548 30394
rect 9220 30184 9272 30190
rect 9220 30126 9272 30132
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9232 29714 9260 29990
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 8760 29038 8812 29044
rect 8850 29064 8906 29073
rect 8484 28960 8536 28966
rect 8484 28902 8536 28908
rect 8680 28762 8708 29038
rect 8668 28756 8720 28762
rect 8668 28698 8720 28704
rect 8772 28626 8800 29038
rect 8850 28999 8906 29008
rect 9324 28966 9352 30348
rect 9496 30330 9548 30336
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9416 29850 9444 30194
rect 9404 29844 9456 29850
rect 9404 29786 9456 29792
rect 8852 28960 8904 28966
rect 8852 28902 8904 28908
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 8864 28694 8892 28902
rect 8852 28688 8904 28694
rect 8852 28630 8904 28636
rect 8944 28688 8996 28694
rect 8944 28630 8996 28636
rect 8760 28620 8812 28626
rect 8760 28562 8812 28568
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8390 28112 8446 28121
rect 8390 28047 8446 28056
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 8588 27946 8616 28358
rect 8956 28257 8984 28630
rect 9128 28620 9180 28626
rect 9128 28562 9180 28568
rect 9312 28620 9364 28626
rect 9312 28562 9364 28568
rect 8942 28248 8998 28257
rect 8942 28183 8998 28192
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8576 27940 8628 27946
rect 8576 27882 8628 27888
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8208 27532 8260 27538
rect 8208 27474 8260 27480
rect 8022 27024 8078 27033
rect 8022 26959 8078 26968
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 7932 26784 7984 26790
rect 7932 26726 7984 26732
rect 7944 26450 7972 26726
rect 7932 26444 7984 26450
rect 7932 26386 7984 26392
rect 7800 26268 7880 26296
rect 7748 26250 7800 26256
rect 7760 25362 7788 26250
rect 7944 25498 7972 26386
rect 8036 25809 8064 26862
rect 8022 25800 8078 25809
rect 8022 25735 8078 25744
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 8128 25401 8156 27474
rect 8220 26450 8248 27474
rect 8404 26926 8432 27882
rect 8588 27577 8616 27882
rect 9048 27878 9076 28154
rect 8760 27872 8812 27878
rect 8760 27814 8812 27820
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 8772 27674 8800 27814
rect 8760 27668 8812 27674
rect 8760 27610 8812 27616
rect 8668 27600 8720 27606
rect 8574 27568 8630 27577
rect 8668 27542 8720 27548
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8574 27503 8630 27512
rect 8576 27328 8628 27334
rect 8576 27270 8628 27276
rect 8392 26920 8444 26926
rect 8312 26880 8392 26908
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 8312 26246 8340 26880
rect 8392 26862 8444 26868
rect 8484 26852 8536 26858
rect 8484 26794 8536 26800
rect 8300 26240 8352 26246
rect 8300 26182 8352 26188
rect 8390 26208 8446 26217
rect 8312 25786 8340 26182
rect 8390 26143 8446 26152
rect 8220 25758 8340 25786
rect 8114 25392 8170 25401
rect 7748 25356 7800 25362
rect 8220 25362 8248 25758
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 8114 25327 8170 25336
rect 8208 25356 8260 25362
rect 7748 25298 7800 25304
rect 7564 25152 7616 25158
rect 7564 25094 7616 25100
rect 7760 24954 7788 25298
rect 7840 25288 7892 25294
rect 8128 25242 8156 25327
rect 8208 25298 8260 25304
rect 7840 25230 7892 25236
rect 7852 24954 7880 25230
rect 8036 25214 8156 25242
rect 7748 24948 7800 24954
rect 7748 24890 7800 24896
rect 7840 24948 7892 24954
rect 7840 24890 7892 24896
rect 7484 24818 7788 24834
rect 7102 24783 7158 24792
rect 7472 24812 7788 24818
rect 7012 24754 7064 24760
rect 7024 24410 7052 24754
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 7012 24132 7064 24138
rect 7012 24074 7064 24080
rect 6918 23216 6974 23225
rect 6828 23180 6880 23186
rect 7024 23186 7052 24074
rect 7116 23730 7144 24783
rect 7524 24806 7788 24812
rect 7472 24754 7524 24760
rect 7760 24750 7788 24806
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7656 24744 7708 24750
rect 7656 24686 7708 24692
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7564 24676 7616 24682
rect 7564 24618 7616 24624
rect 7194 24576 7250 24585
rect 7194 24511 7250 24520
rect 7208 23798 7236 24511
rect 7576 24410 7604 24618
rect 7668 24410 7696 24686
rect 7564 24404 7616 24410
rect 7564 24346 7616 24352
rect 7656 24404 7708 24410
rect 7656 24346 7708 24352
rect 7288 24268 7340 24274
rect 7288 24210 7340 24216
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7300 24177 7328 24210
rect 7286 24168 7342 24177
rect 7484 24138 7512 24210
rect 7286 24103 7342 24112
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7564 23860 7616 23866
rect 7564 23802 7616 23808
rect 7196 23792 7248 23798
rect 7196 23734 7248 23740
rect 7472 23792 7524 23798
rect 7472 23734 7524 23740
rect 7104 23724 7156 23730
rect 7104 23666 7156 23672
rect 7116 23610 7144 23666
rect 7116 23582 7236 23610
rect 6918 23151 6974 23160
rect 7012 23180 7064 23186
rect 6828 23122 6880 23128
rect 6840 23089 6868 23122
rect 6826 23080 6882 23089
rect 6826 23015 6882 23024
rect 6932 22778 6960 23151
rect 7012 23122 7064 23128
rect 7104 23044 7156 23050
rect 7104 22986 7156 22992
rect 7012 22976 7064 22982
rect 7012 22918 7064 22924
rect 6920 22772 6972 22778
rect 6920 22714 6972 22720
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6828 22500 6880 22506
rect 6828 22442 6880 22448
rect 6734 22264 6790 22273
rect 6734 22199 6790 22208
rect 6748 22098 6776 22199
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6734 21992 6790 22001
rect 6734 21927 6790 21936
rect 6748 21894 6776 21927
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6552 21616 6604 21622
rect 6550 21584 6552 21593
rect 6604 21584 6606 21593
rect 6550 21519 6606 21528
rect 6656 21486 6684 21830
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6748 21332 6776 21830
rect 6840 21554 6868 22442
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6932 21486 6960 22374
rect 7024 21622 7052 22918
rect 7116 21622 7144 22986
rect 7208 22030 7236 23582
rect 7286 22128 7342 22137
rect 7286 22063 7342 22072
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7012 21616 7064 21622
rect 7012 21558 7064 21564
rect 7104 21616 7156 21622
rect 7104 21558 7156 21564
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6564 21304 6776 21332
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6564 19310 6592 21304
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6644 21004 6696 21010
rect 6644 20946 6696 20952
rect 6656 20602 6684 20946
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 6644 20392 6696 20398
rect 6644 20334 6696 20340
rect 6656 19514 6684 20334
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6748 19310 6776 21082
rect 6828 20936 6880 20942
rect 6932 20924 6960 21422
rect 7208 21146 7236 21966
rect 7196 21140 7248 21146
rect 7196 21082 7248 21088
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 6880 20896 6960 20924
rect 7104 20936 7156 20942
rect 6828 20878 6880 20884
rect 7104 20878 7156 20884
rect 6840 20398 6868 20878
rect 6920 20800 6972 20806
rect 6920 20742 6972 20748
rect 6932 20534 6960 20742
rect 6920 20528 6972 20534
rect 6920 20470 6972 20476
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 6828 20392 6880 20398
rect 6828 20334 6880 20340
rect 6920 20324 6972 20330
rect 6920 20266 6972 20272
rect 6932 19922 6960 20266
rect 6920 19916 6972 19922
rect 6920 19858 6972 19864
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19394 6868 19654
rect 6840 19366 6960 19394
rect 6460 19304 6512 19310
rect 6458 19272 6460 19281
rect 6552 19304 6604 19310
rect 6512 19272 6514 19281
rect 6552 19246 6604 19252
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6826 19272 6882 19281
rect 6458 19207 6514 19216
rect 6564 18970 6592 19246
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6656 18170 6684 19110
rect 6748 18873 6776 19246
rect 6826 19207 6882 19216
rect 6734 18864 6790 18873
rect 6840 18834 6868 19207
rect 6734 18799 6790 18808
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6932 18170 6960 19366
rect 7024 18970 7052 20402
rect 7116 20058 7144 20878
rect 7208 20777 7236 20946
rect 7194 20768 7250 20777
rect 7194 20703 7250 20712
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7208 20262 7236 20538
rect 7300 20398 7328 22063
rect 7484 21962 7512 23734
rect 7576 22710 7604 23802
rect 7654 23760 7710 23769
rect 7654 23695 7710 23704
rect 7668 23662 7696 23695
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7760 23322 7788 24686
rect 7852 24274 7880 24754
rect 8036 24698 8064 25214
rect 8116 25152 8168 25158
rect 8116 25094 8168 25100
rect 7944 24670 8064 24698
rect 7944 24410 7972 24670
rect 8024 24608 8076 24614
rect 8024 24550 8076 24556
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 8036 24342 8064 24550
rect 8024 24336 8076 24342
rect 8024 24278 8076 24284
rect 7840 24268 7892 24274
rect 7840 24210 7892 24216
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7656 23180 7708 23186
rect 7708 23140 7788 23168
rect 7656 23122 7708 23128
rect 7760 23066 7788 23140
rect 7852 23066 7880 24210
rect 7932 24200 7984 24206
rect 7930 24168 7932 24177
rect 8024 24200 8076 24206
rect 7984 24168 7986 24177
rect 8128 24188 8156 25094
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8220 24274 8248 24550
rect 8208 24268 8260 24274
rect 8208 24210 8260 24216
rect 8076 24160 8156 24188
rect 8024 24142 8076 24148
rect 7930 24103 7986 24112
rect 7944 23322 7972 24103
rect 8036 23866 8064 24142
rect 8024 23860 8076 23866
rect 8024 23802 8076 23808
rect 8220 23798 8248 24210
rect 8312 24177 8340 25638
rect 8298 24168 8354 24177
rect 8298 24103 8354 24112
rect 8300 24064 8352 24070
rect 8300 24006 8352 24012
rect 8208 23792 8260 23798
rect 8208 23734 8260 23740
rect 8220 23610 8248 23734
rect 8128 23582 8248 23610
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 8128 23202 8156 23582
rect 8206 23488 8262 23497
rect 8206 23423 8262 23432
rect 7944 23186 8156 23202
rect 7932 23180 8156 23186
rect 7984 23174 8156 23180
rect 7932 23122 7984 23128
rect 7656 23044 7708 23050
rect 7760 23038 8064 23066
rect 7656 22986 7708 22992
rect 7564 22704 7616 22710
rect 7564 22646 7616 22652
rect 7576 22030 7604 22646
rect 7564 22024 7616 22030
rect 7564 21966 7616 21972
rect 7472 21956 7524 21962
rect 7472 21898 7524 21904
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 21554 7420 21830
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7380 21412 7432 21418
rect 7380 21354 7432 21360
rect 7392 21010 7420 21354
rect 7484 21321 7512 21898
rect 7668 21876 7696 22986
rect 7932 22976 7984 22982
rect 7932 22918 7984 22924
rect 7748 22024 7800 22030
rect 7800 21984 7880 22012
rect 7748 21966 7800 21972
rect 7576 21848 7696 21876
rect 7470 21312 7526 21321
rect 7470 21247 7526 21256
rect 7380 21004 7432 21010
rect 7380 20946 7432 20952
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7392 20913 7420 20946
rect 7378 20904 7434 20913
rect 7378 20839 7434 20848
rect 7378 20632 7434 20641
rect 7378 20567 7434 20576
rect 7288 20392 7340 20398
rect 7288 20334 7340 20340
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7208 19334 7236 20198
rect 7300 19854 7328 20334
rect 7392 20233 7420 20567
rect 7378 20224 7434 20233
rect 7378 20159 7434 20168
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7116 19306 7236 19334
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7010 18864 7066 18873
rect 7010 18799 7012 18808
rect 7064 18799 7066 18808
rect 7012 18770 7064 18776
rect 6656 18142 6776 18170
rect 6460 18080 6512 18086
rect 6460 18022 6512 18028
rect 6472 17746 6500 18022
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6472 17649 6500 17682
rect 6458 17640 6514 17649
rect 6458 17575 6514 17584
rect 6460 17332 6512 17338
rect 6564 17320 6592 17750
rect 6512 17292 6592 17320
rect 6644 17332 6696 17338
rect 6460 17274 6512 17280
rect 6644 17274 6696 17280
rect 6366 17096 6422 17105
rect 6366 17031 6422 17040
rect 6380 16658 6408 17031
rect 6472 16726 6500 17274
rect 6656 17241 6684 17274
rect 6642 17232 6698 17241
rect 6642 17167 6698 17176
rect 6552 17128 6604 17134
rect 6550 17096 6552 17105
rect 6748 17105 6776 18142
rect 6840 18142 6960 18170
rect 7116 18154 7144 19306
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 7208 18154 7236 19110
rect 7392 18154 7420 20159
rect 7484 20058 7512 20946
rect 7576 20602 7604 21848
rect 7656 20936 7708 20942
rect 7656 20878 7708 20884
rect 7748 20936 7800 20942
rect 7748 20878 7800 20884
rect 7564 20596 7616 20602
rect 7564 20538 7616 20544
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7576 18630 7604 20334
rect 7668 19894 7696 20878
rect 7760 20602 7788 20878
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7852 20244 7880 21984
rect 7944 21554 7972 22918
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 7944 20466 7972 20538
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8036 20398 8064 23038
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 8128 22506 8156 22986
rect 8220 22574 8248 23423
rect 8312 23186 8340 24006
rect 8404 23610 8432 26143
rect 8496 25294 8524 26794
rect 8588 26450 8616 27270
rect 8680 26926 8708 27542
rect 8956 27062 8984 27542
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8668 26920 8720 26926
rect 8852 26920 8904 26926
rect 8720 26880 8800 26908
rect 8668 26862 8720 26868
rect 8772 26450 8800 26880
rect 8852 26862 8904 26868
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 8576 26444 8628 26450
rect 8760 26444 8812 26450
rect 8628 26404 8708 26432
rect 8576 26386 8628 26392
rect 8574 25936 8630 25945
rect 8574 25871 8630 25880
rect 8588 25838 8616 25871
rect 8576 25832 8628 25838
rect 8576 25774 8628 25780
rect 8680 25702 8708 26404
rect 8760 26386 8812 26392
rect 8668 25696 8720 25702
rect 8668 25638 8720 25644
rect 8668 25492 8720 25498
rect 8668 25434 8720 25440
rect 8680 25362 8708 25434
rect 8668 25356 8720 25362
rect 8668 25298 8720 25304
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8496 24410 8524 25230
rect 8574 25120 8630 25129
rect 8574 25055 8630 25064
rect 8588 24750 8616 25055
rect 8576 24744 8628 24750
rect 8576 24686 8628 24692
rect 8588 24585 8616 24686
rect 8574 24576 8630 24585
rect 8574 24511 8630 24520
rect 8484 24404 8536 24410
rect 8484 24346 8536 24352
rect 8576 24268 8628 24274
rect 8576 24210 8628 24216
rect 8404 23582 8524 23610
rect 8300 23180 8352 23186
rect 8300 23122 8352 23128
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8390 22944 8446 22953
rect 8208 22568 8260 22574
rect 8208 22510 8260 22516
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 8208 22432 8260 22438
rect 8208 22374 8260 22380
rect 8114 22128 8170 22137
rect 8114 22063 8116 22072
rect 8168 22063 8170 22072
rect 8116 22034 8168 22040
rect 8116 21888 8168 21894
rect 8116 21830 8168 21836
rect 8128 21593 8156 21830
rect 8220 21690 8248 22374
rect 8312 22098 8340 22918
rect 8390 22879 8446 22888
rect 8404 22574 8432 22879
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 8496 22273 8524 23582
rect 8588 23050 8616 24210
rect 8576 23044 8628 23050
rect 8576 22986 8628 22992
rect 8482 22264 8538 22273
rect 8482 22199 8538 22208
rect 8390 22128 8446 22137
rect 8300 22092 8352 22098
rect 8390 22063 8446 22072
rect 8484 22092 8536 22098
rect 8300 22034 8352 22040
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8114 21584 8170 21593
rect 8114 21519 8170 21528
rect 8220 20806 8248 21626
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 8116 20324 8168 20330
rect 8116 20266 8168 20272
rect 7852 20216 8064 20244
rect 7932 19916 7984 19922
rect 7668 19866 7880 19894
rect 7748 19780 7800 19786
rect 7748 19722 7800 19728
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7668 19009 7696 19246
rect 7654 19000 7710 19009
rect 7654 18935 7710 18944
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18222 7696 18566
rect 7760 18222 7788 19722
rect 7852 19446 7880 19866
rect 7932 19858 7984 19864
rect 7944 19514 7972 19858
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7840 19440 7892 19446
rect 7840 19382 7892 19388
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7104 18148 7156 18154
rect 6604 17096 6606 17105
rect 6550 17031 6606 17040
rect 6734 17096 6790 17105
rect 6734 17031 6790 17040
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6644 16992 6696 16998
rect 6840 16980 6868 18142
rect 7104 18090 7156 18096
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7380 18148 7432 18154
rect 7380 18090 7432 18096
rect 6920 18080 6972 18086
rect 6920 18022 6972 18028
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 7194 18048 7250 18057
rect 6644 16934 6696 16940
rect 6748 16952 6868 16980
rect 6460 16720 6512 16726
rect 6564 16697 6592 16934
rect 6460 16662 6512 16668
rect 6550 16688 6606 16697
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6472 16590 6500 16662
rect 6550 16623 6606 16632
rect 6564 16590 6592 16623
rect 6460 16584 6512 16590
rect 6458 16552 6460 16561
rect 6552 16584 6604 16590
rect 6512 16552 6514 16561
rect 6552 16526 6604 16532
rect 6656 16522 6684 16934
rect 6458 16487 6514 16496
rect 6644 16516 6696 16522
rect 6644 16458 6696 16464
rect 6550 16280 6606 16289
rect 6550 16215 6606 16224
rect 6564 16182 6592 16215
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6656 15910 6684 16458
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6368 15564 6420 15570
rect 6368 15506 6420 15512
rect 6104 15026 6132 15506
rect 6184 15088 6236 15094
rect 6184 15030 6236 15036
rect 5828 14980 5948 15008
rect 6092 15020 6144 15026
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5736 14006 5764 14214
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5552 13484 5764 13512
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5552 12918 5580 13330
rect 5540 12912 5592 12918
rect 5540 12854 5592 12860
rect 5632 12776 5684 12782
rect 5632 12718 5684 12724
rect 5460 12406 5580 12434
rect 5262 12336 5318 12345
rect 5172 12300 5224 12306
rect 5092 12260 5172 12288
rect 5262 12271 5318 12280
rect 5448 12300 5500 12306
rect 5172 12242 5224 12248
rect 4908 11608 4936 12174
rect 5000 12158 5120 12186
rect 5092 11914 5120 12158
rect 5092 11886 5212 11914
rect 5080 11688 5132 11694
rect 5080 11630 5132 11636
rect 4988 11620 5040 11626
rect 4908 11580 4988 11608
rect 4988 11562 5040 11568
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 10198 4936 10542
rect 5000 10470 5028 11562
rect 5092 11218 5120 11630
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4896 10056 4948 10062
rect 4802 10024 4858 10033
rect 4896 9998 4948 10004
rect 4802 9959 4804 9968
rect 4856 9959 4858 9968
rect 4804 9930 4856 9936
rect 4908 9382 4936 9998
rect 5000 9586 5028 10066
rect 5092 9926 5120 11154
rect 5184 10606 5212 11886
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10198 5212 10406
rect 5276 10266 5304 12271
rect 5448 12242 5500 12248
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11218 5396 12038
rect 5460 11830 5488 12242
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 5368 9654 5396 10542
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 4988 9580 5040 9586
rect 5040 9540 5120 9568
rect 4988 9522 5040 9528
rect 4988 9444 5040 9450
rect 4988 9386 5040 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8498 4844 8774
rect 4908 8566 4936 8978
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4896 8424 4948 8430
rect 4894 8392 4896 8401
rect 4948 8392 4950 8401
rect 4804 8356 4856 8362
rect 4894 8327 4950 8336
rect 4804 8298 4856 8304
rect 4632 6956 4752 6984
rect 4632 6866 4660 6956
rect 4080 6820 4200 6848
rect 4252 6860 4304 6866
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3662 6556 3970 6565
rect 3662 6554 3668 6556
rect 3724 6554 3748 6556
rect 3804 6554 3828 6556
rect 3884 6554 3908 6556
rect 3964 6554 3970 6556
rect 3724 6502 3726 6554
rect 3906 6502 3908 6554
rect 3662 6500 3668 6502
rect 3724 6500 3748 6502
rect 3804 6500 3828 6502
rect 3884 6500 3908 6502
rect 3964 6500 3970 6502
rect 3662 6491 3970 6500
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3528 5914 3556 6258
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3620 6118 3648 6190
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3620 5914 3648 6054
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 4080 5846 4108 6820
rect 4252 6802 4304 6808
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 3148 5840 3200 5846
rect 4068 5840 4120 5846
rect 3148 5782 3200 5788
rect 3422 5808 3478 5817
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2964 5296 3016 5302
rect 2964 5238 3016 5244
rect 2872 4752 2924 4758
rect 2872 4694 2924 4700
rect 2884 4282 2912 4694
rect 2976 4622 3004 5238
rect 3160 5114 3188 5782
rect 3240 5772 3292 5778
rect 4068 5782 4120 5788
rect 3700 5772 3752 5778
rect 3478 5752 3700 5760
rect 3422 5743 3424 5752
rect 3240 5714 3292 5720
rect 3476 5732 3700 5752
rect 3424 5714 3476 5720
rect 3700 5714 3752 5720
rect 3252 5574 3280 5714
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3662 5468 3970 5477
rect 3662 5466 3668 5468
rect 3724 5466 3748 5468
rect 3804 5466 3828 5468
rect 3884 5466 3908 5468
rect 3964 5466 3970 5468
rect 3724 5414 3726 5466
rect 3906 5414 3908 5466
rect 3662 5412 3668 5414
rect 3724 5412 3748 5414
rect 3804 5412 3828 5414
rect 3884 5412 3908 5414
rect 3964 5412 3970 5414
rect 3662 5403 3970 5412
rect 4172 5370 4200 6666
rect 4540 6458 4568 6666
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4436 6248 4488 6254
rect 4436 6190 4488 6196
rect 4448 6118 4476 6190
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4436 6112 4488 6118
rect 4632 6100 4660 6598
rect 4724 6458 4752 6802
rect 4816 6730 4844 8298
rect 4908 7002 4936 8327
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4908 6458 4936 6802
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4804 6112 4856 6118
rect 4632 6072 4752 6100
rect 4436 6054 4488 6060
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4264 5302 4292 6054
rect 4322 6012 4630 6021
rect 4322 6010 4328 6012
rect 4384 6010 4408 6012
rect 4464 6010 4488 6012
rect 4544 6010 4568 6012
rect 4624 6010 4630 6012
rect 4384 5958 4386 6010
rect 4566 5958 4568 6010
rect 4322 5956 4328 5958
rect 4384 5956 4408 5958
rect 4464 5956 4488 5958
rect 4544 5956 4568 5958
rect 4624 5956 4630 5958
rect 4322 5947 4630 5956
rect 4724 5370 4752 6072
rect 4804 6054 4856 6060
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4816 5302 4844 6054
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4804 5296 4856 5302
rect 5000 5250 5028 9386
rect 5092 8090 5120 9540
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5184 7818 5212 9454
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 8090 5396 8366
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7206 5212 7754
rect 5368 7478 5396 7890
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5460 6984 5488 11630
rect 5552 11014 5580 12406
rect 5644 12306 5672 12718
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5644 11694 5672 12038
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 9586 5580 10406
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 8974 5580 9522
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5538 8664 5594 8673
rect 5538 8599 5540 8608
rect 5592 8599 5594 8608
rect 5540 8570 5592 8576
rect 5644 7936 5672 11222
rect 5736 10810 5764 13484
rect 5828 11694 5856 14980
rect 6092 14962 6144 14968
rect 5908 14884 5960 14890
rect 5908 14826 5960 14832
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5920 10674 5948 14826
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6104 14074 6132 14554
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6196 13954 6224 15030
rect 6380 14618 6408 15506
rect 6656 14890 6684 15846
rect 6748 15026 6776 16952
rect 6828 16652 6880 16658
rect 6828 16594 6880 16600
rect 6840 16250 6868 16594
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6932 16046 6960 18022
rect 7024 17814 7052 18022
rect 7194 17983 7250 17992
rect 7012 17808 7064 17814
rect 7012 17750 7064 17756
rect 7024 17338 7052 17750
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7024 16046 7052 16526
rect 7116 16046 7144 17478
rect 7208 17202 7236 17983
rect 7392 17610 7420 18090
rect 7760 17882 7788 18158
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7564 17808 7616 17814
rect 7564 17750 7616 17756
rect 7576 17649 7604 17750
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7562 17640 7618 17649
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7484 17598 7562 17626
rect 7484 17252 7512 17598
rect 7562 17575 7618 17584
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7300 17224 7512 17252
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7208 17066 7236 17138
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7208 16522 7236 17002
rect 7300 16658 7328 17224
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7392 16697 7420 17070
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7378 16688 7434 16697
rect 7288 16652 7340 16658
rect 7378 16623 7434 16632
rect 7288 16594 7340 16600
rect 7286 16552 7342 16561
rect 7196 16516 7248 16522
rect 7392 16522 7420 16623
rect 7286 16487 7288 16496
rect 7196 16458 7248 16464
rect 7340 16487 7342 16496
rect 7380 16516 7432 16522
rect 7288 16458 7340 16464
rect 7380 16458 7432 16464
rect 7208 16046 7236 16458
rect 7300 16046 7328 16458
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7104 16040 7156 16046
rect 7104 15982 7156 15988
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6368 14612 6420 14618
rect 6368 14554 6420 14560
rect 6276 14544 6328 14550
rect 6276 14486 6328 14492
rect 6012 13926 6224 13954
rect 6012 12102 6040 13926
rect 6288 13852 6316 14486
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6104 13824 6316 13852
rect 6366 13832 6422 13841
rect 6104 12753 6132 13824
rect 6366 13767 6422 13776
rect 6380 13734 6408 13767
rect 6368 13728 6420 13734
rect 6182 13696 6238 13705
rect 6368 13670 6420 13676
rect 6182 13631 6238 13640
rect 6090 12744 6146 12753
rect 6090 12679 6146 12688
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6012 11694 6040 11766
rect 6000 11688 6052 11694
rect 6000 11630 6052 11636
rect 6012 11218 6040 11630
rect 6104 11218 6132 12679
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5368 6956 5488 6984
rect 5552 7908 5672 7936
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5184 6118 5212 6802
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 6390 5304 6598
rect 5264 6384 5316 6390
rect 5264 6326 5316 6332
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5184 5370 5212 5850
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4804 5238 4856 5244
rect 3700 5228 3752 5234
rect 3700 5170 3752 5176
rect 4908 5222 5028 5250
rect 5264 5296 5316 5302
rect 5264 5238 5316 5244
rect 3424 5160 3476 5166
rect 3160 5086 3280 5114
rect 3424 5102 3476 5108
rect 3148 5024 3200 5030
rect 3148 4966 3200 4972
rect 3160 4826 3188 4966
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2700 3738 2728 4082
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2688 3732 2740 3738
rect 2688 3674 2740 3680
rect 2424 3534 2452 3674
rect 2700 3584 2728 3674
rect 2884 3670 2912 4218
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2516 3556 2728 3584
rect 2412 3528 2464 3534
rect 2412 3470 2464 3476
rect 2516 3194 2544 3556
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2240 2446 2268 2994
rect 2516 2990 2544 3130
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2516 2106 2544 2450
rect 2700 2310 2728 3402
rect 2884 2922 2912 3606
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 2976 2774 3004 4558
rect 3252 3602 3280 5086
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3344 4690 3372 5034
rect 3436 4826 3464 5102
rect 3712 4826 3740 5170
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3662 4380 3970 4389
rect 3662 4378 3668 4380
rect 3724 4378 3748 4380
rect 3804 4378 3828 4380
rect 3884 4378 3908 4380
rect 3964 4378 3970 4380
rect 3724 4326 3726 4378
rect 3906 4326 3908 4378
rect 3662 4324 3668 4326
rect 3724 4324 3748 4326
rect 3804 4324 3828 4326
rect 3884 4324 3908 4326
rect 3964 4324 3970 4326
rect 3662 4315 3970 4324
rect 4264 4282 4292 4966
rect 4322 4924 4630 4933
rect 4322 4922 4328 4924
rect 4384 4922 4408 4924
rect 4464 4922 4488 4924
rect 4544 4922 4568 4924
rect 4624 4922 4630 4924
rect 4384 4870 4386 4922
rect 4566 4870 4568 4922
rect 4322 4868 4328 4870
rect 4384 4868 4408 4870
rect 4464 4868 4488 4870
rect 4544 4868 4568 4870
rect 4624 4868 4630 4870
rect 4322 4859 4630 4868
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 2792 2746 3004 2774
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 2504 2100 2556 2106
rect 2504 2042 2556 2048
rect 2596 2032 2648 2038
rect 2596 1974 2648 1980
rect 2044 1964 2096 1970
rect 2044 1906 2096 1912
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 2516 1465 2544 1906
rect 2608 1494 2636 1974
rect 2700 1902 2728 2246
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 2596 1488 2648 1494
rect 2502 1456 2558 1465
rect 2596 1430 2648 1436
rect 2502 1391 2558 1400
rect 1400 1352 1452 1358
rect 1400 1294 1452 1300
rect 2792 814 2820 2746
rect 3160 2514 3188 2994
rect 3252 2990 3280 3538
rect 4080 3534 4108 3878
rect 4172 3738 4200 4082
rect 4448 4010 4476 4422
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4322 3836 4630 3845
rect 4322 3834 4328 3836
rect 4384 3834 4408 3836
rect 4464 3834 4488 3836
rect 4544 3834 4568 3836
rect 4624 3834 4630 3836
rect 4384 3782 4386 3834
rect 4566 3782 4568 3834
rect 4322 3780 4328 3782
rect 4384 3780 4408 3782
rect 4464 3780 4488 3782
rect 4544 3780 4568 3782
rect 4624 3780 4630 3782
rect 4322 3771 4630 3780
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3436 2922 3464 3470
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3528 2650 3556 3470
rect 3662 3292 3970 3301
rect 3662 3290 3668 3292
rect 3724 3290 3748 3292
rect 3804 3290 3828 3292
rect 3884 3290 3908 3292
rect 3964 3290 3970 3292
rect 3724 3238 3726 3290
rect 3906 3238 3908 3290
rect 3662 3236 3668 3238
rect 3724 3236 3748 3238
rect 3804 3236 3828 3238
rect 3884 3236 3908 3238
rect 3964 3236 3970 3238
rect 3662 3227 3970 3236
rect 4724 3194 4752 3538
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3662 2204 3970 2213
rect 3662 2202 3668 2204
rect 3724 2202 3748 2204
rect 3804 2202 3828 2204
rect 3884 2202 3908 2204
rect 3964 2202 3970 2204
rect 3724 2150 3726 2202
rect 3906 2150 3908 2202
rect 3662 2148 3668 2150
rect 3724 2148 3748 2150
rect 3804 2148 3828 2150
rect 3884 2148 3908 2150
rect 3964 2148 3970 2150
rect 3662 2139 3970 2148
rect 3332 2100 3384 2106
rect 3332 2042 3384 2048
rect 3344 1766 3372 2042
rect 4172 1970 4200 2926
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4264 2582 4292 2858
rect 4322 2748 4630 2757
rect 4322 2746 4328 2748
rect 4384 2746 4408 2748
rect 4464 2746 4488 2748
rect 4544 2746 4568 2748
rect 4624 2746 4630 2748
rect 4384 2694 4386 2746
rect 4566 2694 4568 2746
rect 4322 2692 4328 2694
rect 4384 2692 4408 2694
rect 4464 2692 4488 2694
rect 4544 2692 4568 2694
rect 4624 2692 4630 2694
rect 4322 2683 4630 2692
rect 4252 2576 4304 2582
rect 4252 2518 4304 2524
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 3424 1896 3476 1902
rect 3424 1838 3476 1844
rect 3332 1760 3384 1766
rect 3332 1702 3384 1708
rect 2780 808 2832 814
rect 2780 750 2832 756
rect 3344 746 3372 1702
rect 3436 882 3464 1838
rect 3528 1426 3556 1906
rect 3608 1896 3660 1902
rect 3608 1838 3660 1844
rect 3792 1896 3844 1902
rect 3792 1838 3844 1844
rect 3516 1420 3568 1426
rect 3516 1362 3568 1368
rect 3528 1018 3556 1362
rect 3620 1290 3648 1838
rect 3804 1562 3832 1838
rect 3792 1556 3844 1562
rect 3792 1498 3844 1504
rect 4264 1426 4292 2518
rect 4322 1660 4630 1669
rect 4322 1658 4328 1660
rect 4384 1658 4408 1660
rect 4464 1658 4488 1660
rect 4544 1658 4568 1660
rect 4624 1658 4630 1660
rect 4384 1606 4386 1658
rect 4566 1606 4568 1658
rect 4322 1604 4328 1606
rect 4384 1604 4408 1606
rect 4464 1604 4488 1606
rect 4544 1604 4568 1606
rect 4624 1604 4630 1606
rect 4322 1595 4630 1604
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 3662 1116 3970 1125
rect 3662 1114 3668 1116
rect 3724 1114 3748 1116
rect 3804 1114 3828 1116
rect 3884 1114 3908 1116
rect 3964 1114 3970 1116
rect 3724 1062 3726 1114
rect 3906 1062 3908 1114
rect 3662 1060 3668 1062
rect 3724 1060 3748 1062
rect 3804 1060 3828 1062
rect 3884 1060 3908 1062
rect 3964 1060 3970 1062
rect 3662 1051 3970 1060
rect 3516 1012 3568 1018
rect 3516 954 3568 960
rect 3424 876 3476 882
rect 3424 818 3476 824
rect 3976 808 4028 814
rect 3976 750 4028 756
rect 3332 740 3384 746
rect 3332 682 3384 688
rect 3988 678 4016 750
rect 4080 746 4108 1294
rect 4816 1222 4844 5102
rect 4908 3398 4936 5222
rect 4988 5160 5040 5166
rect 4988 5102 5040 5108
rect 5000 4690 5028 5102
rect 5276 5098 5304 5238
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 5000 4282 5028 4626
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 4988 4276 5040 4282
rect 4988 4218 5040 4224
rect 5276 4146 5304 4490
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 4988 4072 5040 4078
rect 4988 4014 5040 4020
rect 5000 3670 5028 4014
rect 4988 3664 5040 3670
rect 4988 3606 5040 3612
rect 5184 3602 5212 4082
rect 5276 3738 5304 4082
rect 5264 3732 5316 3738
rect 5264 3674 5316 3680
rect 5368 3602 5396 6956
rect 5552 6914 5580 7908
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7342 5672 7686
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5736 7274 5764 8434
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 5460 6886 5580 6914
rect 5460 6798 5488 6886
rect 5632 6860 5684 6866
rect 5552 6820 5632 6848
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5552 6254 5580 6820
rect 5632 6802 5684 6808
rect 5828 6798 5856 9862
rect 5920 9602 5948 10610
rect 6104 10538 6132 11154
rect 6196 10674 6224 13631
rect 6380 13530 6408 13670
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6472 12782 6500 13874
rect 6564 13870 6592 14758
rect 6932 14482 6960 14758
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6736 14340 6788 14346
rect 6736 14282 6788 14288
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6644 13864 6696 13870
rect 6644 13806 6696 13812
rect 6656 13394 6684 13806
rect 6748 13530 6776 14282
rect 6840 14074 6868 14282
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6840 13410 6868 13670
rect 6644 13388 6696 13394
rect 6644 13330 6696 13336
rect 6748 13382 6868 13410
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6564 12782 6592 12922
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6368 12300 6420 12306
rect 6368 12242 6420 12248
rect 6276 12164 6328 12170
rect 6276 12106 6328 12112
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10532 6144 10538
rect 6092 10474 6144 10480
rect 6288 10130 6316 12106
rect 6380 11898 6408 12242
rect 6368 11892 6420 11898
rect 6368 11834 6420 11840
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 5920 9574 6040 9602
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5920 9042 5948 9454
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 5920 7410 5948 7890
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6012 7342 6040 9574
rect 6288 9518 6316 9862
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6380 8922 6408 11562
rect 6564 11218 6592 12718
rect 6656 12442 6684 13330
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6748 12306 6776 13382
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12306 6868 12854
rect 7024 12782 7052 15506
rect 7116 14278 7144 15982
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7208 15366 7236 15506
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7208 14958 7236 15302
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7288 14952 7340 14958
rect 7340 14912 7420 14940
rect 7288 14894 7340 14900
rect 7104 14272 7156 14278
rect 7104 14214 7156 14220
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6748 12209 6776 12242
rect 6734 12200 6790 12209
rect 6656 12158 6734 12186
rect 6656 11354 6684 12158
rect 6734 12135 6790 12144
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6748 11694 6776 12038
rect 6736 11688 6788 11694
rect 6736 11630 6788 11636
rect 6932 11354 6960 12650
rect 7024 12617 7052 12718
rect 7010 12608 7066 12617
rect 7010 12543 7066 12552
rect 7012 12368 7064 12374
rect 7010 12336 7012 12345
rect 7064 12336 7066 12345
rect 7116 12306 7144 13330
rect 7208 12782 7236 14894
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7300 13462 7328 14350
rect 7392 13802 7420 14912
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7300 12434 7328 13126
rect 7208 12406 7328 12434
rect 7010 12271 7066 12280
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7104 12096 7156 12102
rect 7102 12064 7104 12073
rect 7156 12064 7158 12073
rect 7102 11999 7158 12008
rect 7012 11688 7064 11694
rect 7064 11648 7144 11676
rect 7012 11630 7064 11636
rect 7012 11552 7064 11558
rect 7012 11494 7064 11500
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7024 11218 7052 11494
rect 7116 11354 7144 11648
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 6932 10742 6960 11154
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6460 10668 6512 10674
rect 6460 10610 6512 10616
rect 6472 9042 6500 10610
rect 6932 10606 6960 10678
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6564 9654 6592 10542
rect 7104 10532 7156 10538
rect 7104 10474 7156 10480
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6828 9988 6880 9994
rect 6828 9930 6880 9936
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 6380 8894 6500 8922
rect 6368 8832 6420 8838
rect 6368 8774 6420 8780
rect 6380 8430 6408 8774
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6104 7478 6132 8366
rect 6196 8090 6224 8366
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 6000 7336 6052 7342
rect 6000 7278 6052 7284
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5920 6254 5948 6734
rect 6012 6254 6040 7278
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 6104 6458 6132 6802
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5540 6248 5592 6254
rect 5540 6190 5592 6196
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5460 4690 5488 5102
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5460 3738 5488 4014
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 5184 2106 5212 3538
rect 5368 2774 5396 3538
rect 5368 2746 5488 2774
rect 5460 2514 5488 2746
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5552 2038 5580 6190
rect 6012 5166 6040 6190
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 5736 5030 5764 5102
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4758 5764 4966
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 4282 5856 4558
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5828 1902 5856 2450
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 5816 1896 5868 1902
rect 5816 1838 5868 1844
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 4908 1426 4936 1702
rect 5184 1562 5212 1838
rect 5172 1556 5224 1562
rect 5172 1498 5224 1504
rect 5828 1442 5856 1838
rect 5920 1834 5948 5034
rect 6472 4826 6500 8894
rect 6656 8634 6684 9454
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6748 8430 6776 9454
rect 6840 9178 6868 9930
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6840 9042 6868 9114
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6932 8974 6960 10406
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 7024 8498 7052 9590
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7342 6684 7754
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 6932 7342 6960 7686
rect 7024 7426 7052 7890
rect 7116 7546 7144 10474
rect 7208 7818 7236 12406
rect 7392 12345 7420 13738
rect 7484 12850 7512 16934
rect 7576 16046 7604 17274
rect 7668 17134 7696 17546
rect 7760 17202 7788 17682
rect 7852 17610 7880 19382
rect 7932 19304 7984 19310
rect 7930 19272 7932 19281
rect 7984 19272 7986 19281
rect 7930 19207 7986 19216
rect 7930 19000 7986 19009
rect 7930 18935 7986 18944
rect 7944 18290 7972 18935
rect 8036 18290 8064 20216
rect 8128 19310 8156 20266
rect 8220 20058 8248 20742
rect 8312 20641 8340 22034
rect 8404 21690 8432 22063
rect 8484 22034 8536 22040
rect 8392 21684 8444 21690
rect 8392 21626 8444 21632
rect 8496 21570 8524 22034
rect 8404 21542 8524 21570
rect 8404 21010 8432 21542
rect 8484 21412 8536 21418
rect 8484 21354 8536 21360
rect 8392 21004 8444 21010
rect 8392 20946 8444 20952
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8298 20632 8354 20641
rect 8298 20567 8354 20576
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8312 19922 8340 20402
rect 8404 20398 8432 20810
rect 8496 20398 8524 21354
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8484 20392 8536 20398
rect 8588 20380 8616 22986
rect 8680 22234 8708 25298
rect 8772 24954 8800 26386
rect 8864 26382 8892 26862
rect 8956 26586 8984 26862
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8852 26376 8904 26382
rect 8852 26318 8904 26324
rect 8944 26240 8996 26246
rect 8944 26182 8996 26188
rect 8852 25832 8904 25838
rect 8852 25774 8904 25780
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8758 24712 8814 24721
rect 8758 24647 8814 24656
rect 8772 22658 8800 24647
rect 8864 24426 8892 25774
rect 8956 24614 8984 26182
rect 9048 25838 9076 27814
rect 9140 27130 9168 28562
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 9232 28218 9260 28358
rect 9220 28212 9272 28218
rect 9220 28154 9272 28160
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 9232 27470 9260 27950
rect 9324 27674 9352 28562
rect 9312 27668 9364 27674
rect 9312 27610 9364 27616
rect 9220 27464 9272 27470
rect 9220 27406 9272 27412
rect 9324 27402 9352 27610
rect 9312 27396 9364 27402
rect 9312 27338 9364 27344
rect 9128 27124 9180 27130
rect 9128 27066 9180 27072
rect 9220 26920 9272 26926
rect 9416 26874 9444 29786
rect 9508 29170 9536 30194
rect 9496 29164 9548 29170
rect 9496 29106 9548 29112
rect 9600 28937 9628 30602
rect 9692 29714 9720 31719
rect 9784 31657 9812 32014
rect 9770 31648 9826 31657
rect 9770 31583 9826 31592
rect 9772 31272 9824 31278
rect 9876 31260 9904 32150
rect 10336 32042 10364 32399
rect 9824 31232 9904 31260
rect 9968 32014 10364 32042
rect 9772 31214 9824 31220
rect 9680 29708 9732 29714
rect 9680 29650 9732 29656
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 9586 28928 9642 28937
rect 9586 28863 9642 28872
rect 9588 28756 9640 28762
rect 9588 28698 9640 28704
rect 9600 27878 9628 28698
rect 9692 28626 9720 29106
rect 9680 28620 9732 28626
rect 9680 28562 9732 28568
rect 9784 28558 9812 31214
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9876 30569 9904 30670
rect 9862 30560 9918 30569
rect 9862 30495 9918 30504
rect 9862 30424 9918 30433
rect 9862 30359 9918 30368
rect 9876 29617 9904 30359
rect 9968 30190 9996 32014
rect 10062 31580 10370 31589
rect 10062 31578 10068 31580
rect 10124 31578 10148 31580
rect 10204 31578 10228 31580
rect 10284 31578 10308 31580
rect 10364 31578 10370 31580
rect 10124 31526 10126 31578
rect 10306 31526 10308 31578
rect 10062 31524 10068 31526
rect 10124 31524 10148 31526
rect 10204 31524 10228 31526
rect 10284 31524 10308 31526
rect 10364 31524 10370 31526
rect 10062 31515 10370 31524
rect 10428 31482 10456 32728
rect 10520 32473 10548 32966
rect 10612 32570 10640 33934
rect 10980 33300 11008 34054
rect 11152 34002 11204 34008
rect 11256 34054 11376 34082
rect 11426 34096 11482 34105
rect 11058 33960 11114 33969
rect 11058 33895 11060 33904
rect 11112 33895 11114 33904
rect 11152 33924 11204 33930
rect 11060 33866 11112 33872
rect 11152 33866 11204 33872
rect 10980 33272 11100 33300
rect 10722 33212 11030 33221
rect 10722 33210 10728 33212
rect 10784 33210 10808 33212
rect 10864 33210 10888 33212
rect 10944 33210 10968 33212
rect 11024 33210 11030 33212
rect 10784 33158 10786 33210
rect 10966 33158 10968 33210
rect 10722 33156 10728 33158
rect 10784 33156 10808 33158
rect 10864 33156 10888 33158
rect 10944 33156 10968 33158
rect 11024 33156 11030 33158
rect 10722 33147 11030 33156
rect 10876 33108 10928 33114
rect 10876 33050 10928 33056
rect 10692 33040 10744 33046
rect 10888 33017 10916 33050
rect 10692 32982 10744 32988
rect 10874 33008 10930 33017
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10506 32464 10562 32473
rect 10506 32399 10562 32408
rect 10600 32292 10652 32298
rect 10520 32252 10600 32280
rect 10140 31476 10192 31482
rect 10140 31418 10192 31424
rect 10416 31476 10468 31482
rect 10416 31418 10468 31424
rect 10152 30802 10180 31418
rect 10232 30864 10284 30870
rect 10230 30832 10232 30841
rect 10284 30832 10286 30841
rect 10048 30796 10100 30802
rect 10048 30738 10100 30744
rect 10140 30796 10192 30802
rect 10230 30767 10286 30776
rect 10140 30738 10192 30744
rect 10060 30705 10088 30738
rect 10046 30696 10102 30705
rect 10046 30631 10102 30640
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10062 30492 10370 30501
rect 10062 30490 10068 30492
rect 10124 30490 10148 30492
rect 10204 30490 10228 30492
rect 10284 30490 10308 30492
rect 10364 30490 10370 30492
rect 10124 30438 10126 30490
rect 10306 30438 10308 30490
rect 10062 30436 10068 30438
rect 10124 30436 10148 30438
rect 10204 30436 10228 30438
rect 10284 30436 10308 30438
rect 10364 30436 10370 30438
rect 10062 30427 10370 30436
rect 10232 30320 10284 30326
rect 10230 30288 10232 30297
rect 10284 30288 10286 30297
rect 10230 30223 10286 30232
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 10046 30152 10102 30161
rect 10046 30087 10102 30096
rect 10232 30116 10284 30122
rect 9956 30048 10008 30054
rect 10060 30036 10088 30087
rect 10232 30058 10284 30064
rect 10008 30008 10088 30036
rect 9956 29990 10008 29996
rect 9862 29608 9918 29617
rect 9862 29543 9918 29552
rect 9876 29209 9904 29543
rect 9862 29200 9918 29209
rect 9862 29135 9918 29144
rect 9968 29016 9996 29990
rect 10138 29880 10194 29889
rect 10138 29815 10140 29824
rect 10192 29815 10194 29824
rect 10140 29786 10192 29792
rect 10244 29753 10272 30058
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10336 29850 10364 29990
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10230 29744 10286 29753
rect 10230 29679 10286 29688
rect 10232 29640 10284 29646
rect 10230 29608 10232 29617
rect 10284 29608 10286 29617
rect 10230 29543 10286 29552
rect 10062 29404 10370 29413
rect 10062 29402 10068 29404
rect 10124 29402 10148 29404
rect 10204 29402 10228 29404
rect 10284 29402 10308 29404
rect 10364 29402 10370 29404
rect 10124 29350 10126 29402
rect 10306 29350 10308 29402
rect 10062 29348 10068 29350
rect 10124 29348 10148 29350
rect 10204 29348 10228 29350
rect 10284 29348 10308 29350
rect 10364 29348 10370 29350
rect 10062 29339 10370 29348
rect 10428 29102 10456 30534
rect 10520 30025 10548 32252
rect 10704 32280 10732 32982
rect 11072 32994 11100 33272
rect 10874 32943 10930 32952
rect 10980 32966 11100 32994
rect 10652 32252 10732 32280
rect 10980 32280 11008 32966
rect 11164 32910 11192 33866
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 10980 32252 11100 32280
rect 10600 32234 10652 32240
rect 10722 32124 11030 32133
rect 10722 32122 10728 32124
rect 10784 32122 10808 32124
rect 10864 32122 10888 32124
rect 10944 32122 10968 32124
rect 11024 32122 11030 32124
rect 10784 32070 10786 32122
rect 10966 32070 10968 32122
rect 10722 32068 10728 32070
rect 10784 32068 10808 32070
rect 10864 32068 10888 32070
rect 10944 32068 10968 32070
rect 11024 32068 11030 32070
rect 10722 32059 11030 32068
rect 10876 31952 10928 31958
rect 10876 31894 10928 31900
rect 10888 31754 10916 31894
rect 10968 31884 11020 31890
rect 10968 31826 11020 31832
rect 10876 31748 10928 31754
rect 10876 31690 10928 31696
rect 10692 31680 10744 31686
rect 10690 31648 10692 31657
rect 10744 31648 10746 31657
rect 10690 31583 10746 31592
rect 10888 31346 10916 31690
rect 10876 31340 10928 31346
rect 10876 31282 10928 31288
rect 10980 31226 11008 31826
rect 10612 31198 11008 31226
rect 10612 30938 10640 31198
rect 10722 31036 11030 31045
rect 10722 31034 10728 31036
rect 10784 31034 10808 31036
rect 10864 31034 10888 31036
rect 10944 31034 10968 31036
rect 11024 31034 11030 31036
rect 10784 30982 10786 31034
rect 10966 30982 10968 31034
rect 10722 30980 10728 30982
rect 10784 30980 10808 30982
rect 10864 30980 10888 30982
rect 10944 30980 10968 30982
rect 11024 30980 11030 30982
rect 10722 30971 11030 30980
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10612 30326 10640 30874
rect 10692 30864 10744 30870
rect 11072 30852 11100 32252
rect 11152 31680 11204 31686
rect 11152 31622 11204 31628
rect 11164 31278 11192 31622
rect 11152 31272 11204 31278
rect 11152 31214 11204 31220
rect 11152 31136 11204 31142
rect 11152 31078 11204 31084
rect 10692 30806 10744 30812
rect 10782 30832 10838 30841
rect 10600 30320 10652 30326
rect 10600 30262 10652 30268
rect 10704 30036 10732 30806
rect 10782 30767 10838 30776
rect 10980 30824 11100 30852
rect 10796 30394 10824 30767
rect 10980 30734 11008 30824
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10966 30424 11022 30433
rect 10784 30388 10836 30394
rect 10966 30359 11022 30368
rect 10784 30330 10836 30336
rect 10980 30138 11008 30359
rect 10980 30110 11100 30138
rect 10506 30016 10562 30025
rect 10506 29951 10562 29960
rect 10644 30008 10732 30036
rect 10508 29844 10560 29850
rect 10644 29832 10672 30008
rect 10722 29948 11030 29957
rect 10722 29946 10728 29948
rect 10784 29946 10808 29948
rect 10864 29946 10888 29948
rect 10944 29946 10968 29948
rect 11024 29946 11030 29948
rect 10784 29894 10786 29946
rect 10966 29894 10968 29946
rect 10722 29892 10728 29894
rect 10784 29892 10808 29894
rect 10864 29892 10888 29894
rect 10944 29892 10968 29894
rect 11024 29892 11030 29894
rect 10722 29883 11030 29892
rect 11072 29832 11100 30110
rect 10644 29804 10916 29832
rect 10508 29786 10560 29792
rect 10520 29238 10548 29786
rect 10690 29744 10746 29753
rect 10600 29708 10652 29714
rect 10690 29679 10746 29688
rect 10600 29650 10652 29656
rect 10612 29481 10640 29650
rect 10598 29472 10654 29481
rect 10598 29407 10654 29416
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10598 29200 10654 29209
rect 10598 29135 10654 29144
rect 10612 29102 10640 29135
rect 10416 29096 10468 29102
rect 10416 29038 10468 29044
rect 10600 29096 10652 29102
rect 10600 29038 10652 29044
rect 10048 29028 10100 29034
rect 9968 28988 10048 29016
rect 10048 28970 10100 28976
rect 10508 29028 10560 29034
rect 10704 28994 10732 29679
rect 10784 29504 10836 29510
rect 10784 29446 10836 29452
rect 10796 29170 10824 29446
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10508 28970 10560 28976
rect 9864 28960 9916 28966
rect 9864 28902 9916 28908
rect 9876 28626 9904 28902
rect 9864 28620 9916 28626
rect 9864 28562 9916 28568
rect 9772 28552 9824 28558
rect 9772 28494 9824 28500
rect 9680 28484 9732 28490
rect 9680 28426 9732 28432
rect 9588 27872 9640 27878
rect 9588 27814 9640 27820
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9588 27668 9640 27674
rect 9588 27610 9640 27616
rect 9220 26862 9272 26868
rect 9126 26616 9182 26625
rect 9232 26586 9260 26862
rect 9324 26846 9444 26874
rect 9126 26551 9182 26560
rect 9220 26580 9272 26586
rect 9140 26450 9168 26551
rect 9220 26522 9272 26528
rect 9128 26444 9180 26450
rect 9128 26386 9180 26392
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 9128 25764 9180 25770
rect 9128 25706 9180 25712
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 9048 24750 9076 25162
rect 9140 24750 9168 25706
rect 9232 24818 9260 26522
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9036 24744 9088 24750
rect 9128 24744 9180 24750
rect 9036 24686 9088 24692
rect 9126 24712 9128 24721
rect 9180 24712 9182 24721
rect 9126 24647 9182 24656
rect 9220 24676 9272 24682
rect 9220 24618 9272 24624
rect 8944 24608 8996 24614
rect 8944 24550 8996 24556
rect 8864 24398 8984 24426
rect 9232 24410 9260 24618
rect 8852 22976 8904 22982
rect 8852 22918 8904 22924
rect 8864 22778 8892 22918
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8956 22681 8984 24398
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9034 24168 9090 24177
rect 9034 24103 9090 24112
rect 9048 23254 9076 24103
rect 9036 23248 9088 23254
rect 9088 23208 9168 23236
rect 9036 23190 9088 23196
rect 8942 22672 8998 22681
rect 8772 22630 8892 22658
rect 8864 22574 8892 22630
rect 8942 22607 8998 22616
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8668 22228 8720 22234
rect 8668 22170 8720 22176
rect 8680 21486 8708 22170
rect 8760 21548 8812 21554
rect 8760 21490 8812 21496
rect 8668 21480 8720 21486
rect 8668 21422 8720 21428
rect 8680 20482 8708 21422
rect 8772 20602 8800 21490
rect 8864 20618 8892 22510
rect 8956 22098 8984 22607
rect 9036 22568 9088 22574
rect 9140 22556 9168 23208
rect 9232 23186 9260 24346
rect 9324 24274 9352 26846
rect 9404 26784 9456 26790
rect 9404 26726 9456 26732
rect 9416 26450 9444 26726
rect 9404 26444 9456 26450
rect 9404 26386 9456 26392
rect 9416 25838 9444 26386
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9508 25378 9536 27610
rect 9600 27577 9628 27610
rect 9586 27568 9642 27577
rect 9692 27538 9720 28426
rect 9586 27503 9642 27512
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9692 27441 9720 27474
rect 9678 27432 9734 27441
rect 9678 27367 9734 27376
rect 9678 27160 9734 27169
rect 9678 27095 9734 27104
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9600 25430 9628 25638
rect 9416 25350 9536 25378
rect 9588 25424 9640 25430
rect 9588 25366 9640 25372
rect 9416 24818 9444 25350
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9508 24954 9536 25230
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9404 24812 9456 24818
rect 9404 24754 9456 24760
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9312 24268 9364 24274
rect 9312 24210 9364 24216
rect 9220 23180 9272 23186
rect 9220 23122 9272 23128
rect 9324 23168 9352 24210
rect 9416 23322 9444 24346
rect 9600 24206 9628 24686
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9496 24132 9548 24138
rect 9496 24074 9548 24080
rect 9404 23316 9456 23322
rect 9404 23258 9456 23264
rect 9404 23180 9456 23186
rect 9324 23140 9404 23168
rect 9220 22568 9272 22574
rect 9140 22528 9220 22556
rect 9036 22510 9088 22516
rect 9220 22510 9272 22516
rect 8944 22092 8996 22098
rect 8944 22034 8996 22040
rect 8956 21146 8984 22034
rect 9048 21350 9076 22510
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 9140 22096 9168 22374
rect 9128 22090 9180 22096
rect 9128 22032 9180 22038
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9232 21865 9260 21966
rect 9218 21856 9274 21865
rect 9218 21791 9274 21800
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9034 21040 9090 21049
rect 9034 20975 9090 20984
rect 8760 20596 8812 20602
rect 8864 20590 8984 20618
rect 8760 20538 8812 20544
rect 8680 20454 8800 20482
rect 8772 20398 8800 20454
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8668 20392 8720 20398
rect 8588 20352 8668 20380
rect 8484 20334 8536 20340
rect 8668 20334 8720 20340
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8298 19816 8354 19825
rect 8298 19751 8300 19760
rect 8352 19751 8354 19760
rect 8300 19722 8352 19728
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8116 19304 8168 19310
rect 8116 19246 8168 19252
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8024 18080 8076 18086
rect 8024 18022 8076 18028
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7944 17785 7972 17818
rect 7930 17776 7986 17785
rect 7930 17711 7986 17720
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7852 17338 7880 17546
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7748 17196 7800 17202
rect 7748 17138 7800 17144
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7656 16992 7708 16998
rect 7656 16934 7708 16940
rect 7668 16561 7696 16934
rect 7760 16658 7788 17138
rect 7852 16794 7880 17274
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7944 16794 7972 17070
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7838 16688 7894 16697
rect 7748 16652 7800 16658
rect 8036 16658 8064 18022
rect 7838 16623 7894 16632
rect 8024 16652 8076 16658
rect 7748 16594 7800 16600
rect 7654 16552 7710 16561
rect 7654 16487 7710 16496
rect 7656 16448 7708 16454
rect 7656 16390 7708 16396
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7576 13938 7604 15846
rect 7668 15570 7696 16390
rect 7760 16114 7788 16594
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7852 15960 7880 16623
rect 8024 16594 8076 16600
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7932 15972 7984 15978
rect 7852 15932 7932 15960
rect 7852 15570 7880 15932
rect 7932 15914 7984 15920
rect 8036 15570 8064 15982
rect 7656 15564 7708 15570
rect 7840 15564 7892 15570
rect 7656 15506 7708 15512
rect 7760 15524 7840 15552
rect 7668 15094 7696 15506
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7472 12368 7524 12374
rect 7378 12336 7434 12345
rect 7472 12310 7524 12316
rect 7378 12271 7434 12280
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7300 11354 7328 12106
rect 7484 11778 7512 12310
rect 7392 11750 7512 11778
rect 7576 11778 7604 13466
rect 7668 12481 7696 14418
rect 7760 12986 7788 15524
rect 7840 15506 7892 15512
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 7838 15056 7894 15065
rect 7838 14991 7840 15000
rect 7892 14991 7894 15000
rect 7840 14962 7892 14968
rect 7840 14816 7892 14822
rect 7840 14758 7892 14764
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7746 12880 7802 12889
rect 7746 12815 7748 12824
rect 7800 12815 7802 12824
rect 7748 12786 7800 12792
rect 7852 12646 7880 14758
rect 7944 14346 7972 15506
rect 8128 14482 8156 18906
rect 8220 18834 8248 19654
rect 8404 19446 8432 20334
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19990 8524 20198
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8484 19984 8536 19990
rect 8484 19926 8536 19932
rect 8392 19440 8444 19446
rect 8392 19382 8444 19388
rect 8482 19408 8538 19417
rect 8482 19343 8538 19352
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8208 18828 8260 18834
rect 8208 18770 8260 18776
rect 8312 18426 8340 19246
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8404 18426 8432 18770
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8392 18420 8444 18426
rect 8392 18362 8444 18368
rect 8392 18080 8444 18086
rect 8392 18022 8444 18028
rect 8404 17814 8432 18022
rect 8392 17808 8444 17814
rect 8206 17776 8262 17785
rect 8392 17750 8444 17756
rect 8262 17720 8340 17728
rect 8206 17711 8208 17720
rect 8260 17700 8340 17720
rect 8208 17682 8260 17688
rect 8208 17128 8260 17134
rect 8208 17070 8260 17076
rect 8220 16250 8248 17070
rect 8312 16658 8340 17700
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8404 16590 8432 17614
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8496 16130 8524 19343
rect 8588 19310 8616 19994
rect 8680 19786 8708 20334
rect 8864 19990 8892 20402
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8668 19780 8720 19786
rect 8668 19722 8720 19728
rect 8772 19514 8800 19790
rect 8864 19514 8892 19926
rect 8760 19508 8812 19514
rect 8760 19450 8812 19456
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8666 19408 8722 19417
rect 8666 19343 8722 19352
rect 8576 19304 8628 19310
rect 8576 19246 8628 19252
rect 8588 18057 8616 19246
rect 8680 19174 8708 19343
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8956 18970 8984 20590
rect 9048 19854 9076 20975
rect 9324 20534 9352 23140
rect 9404 23122 9456 23128
rect 9404 22432 9456 22438
rect 9404 22374 9456 22380
rect 9416 22166 9444 22374
rect 9404 22160 9456 22166
rect 9404 22102 9456 22108
rect 9508 20777 9536 24074
rect 9692 23497 9720 27095
rect 9784 26994 9812 28494
rect 9876 28014 9904 28562
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9772 26852 9824 26858
rect 9772 26794 9824 26800
rect 9784 25770 9812 26794
rect 9864 25900 9916 25906
rect 9864 25842 9916 25848
rect 9772 25764 9824 25770
rect 9772 25706 9824 25712
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9784 24732 9812 25230
rect 9876 24886 9904 25842
rect 9968 25480 9996 28358
rect 10062 28316 10370 28325
rect 10062 28314 10068 28316
rect 10124 28314 10148 28316
rect 10204 28314 10228 28316
rect 10284 28314 10308 28316
rect 10364 28314 10370 28316
rect 10124 28262 10126 28314
rect 10306 28262 10308 28314
rect 10062 28260 10068 28262
rect 10124 28260 10148 28262
rect 10204 28260 10228 28262
rect 10284 28260 10308 28262
rect 10364 28260 10370 28262
rect 10062 28251 10370 28260
rect 10230 28112 10286 28121
rect 10230 28047 10286 28056
rect 10244 27674 10272 28047
rect 10428 28014 10456 28358
rect 10520 28121 10548 28970
rect 10612 28966 10732 28994
rect 10888 28994 10916 29804
rect 10980 29804 11100 29832
rect 10980 29306 11008 29804
rect 11058 29744 11114 29753
rect 11058 29679 11060 29688
rect 11112 29679 11114 29688
rect 11060 29650 11112 29656
rect 11058 29336 11114 29345
rect 10968 29300 11020 29306
rect 11058 29271 11060 29280
rect 10968 29242 11020 29248
rect 11112 29271 11114 29280
rect 11060 29242 11112 29248
rect 10888 28966 11100 28994
rect 10612 28218 10640 28966
rect 10722 28860 11030 28869
rect 10722 28858 10728 28860
rect 10784 28858 10808 28860
rect 10864 28858 10888 28860
rect 10944 28858 10968 28860
rect 11024 28858 11030 28860
rect 10784 28806 10786 28858
rect 10966 28806 10968 28858
rect 10722 28804 10728 28806
rect 10784 28804 10808 28806
rect 10864 28804 10888 28806
rect 10944 28804 10968 28806
rect 11024 28804 11030 28806
rect 10722 28795 11030 28804
rect 11072 28744 11100 28966
rect 10980 28716 11100 28744
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10506 28112 10562 28121
rect 10506 28047 10562 28056
rect 10416 28008 10468 28014
rect 10416 27950 10468 27956
rect 10508 28008 10560 28014
rect 10508 27950 10560 27956
rect 10980 27962 11008 28716
rect 11164 28642 11192 31078
rect 11256 29102 11284 34054
rect 11426 34031 11482 34040
rect 11336 33992 11388 33998
rect 11532 33969 11560 35770
rect 11624 34474 11652 39374
rect 11808 39370 11836 40938
rect 11888 40384 11940 40390
rect 11888 40326 11940 40332
rect 11900 39914 11928 40326
rect 11888 39908 11940 39914
rect 11888 39850 11940 39856
rect 11886 39536 11942 39545
rect 11886 39471 11942 39480
rect 11796 39364 11848 39370
rect 11796 39306 11848 39312
rect 11900 38944 11928 39471
rect 11808 38916 11928 38944
rect 11704 38548 11756 38554
rect 11704 38490 11756 38496
rect 11716 37330 11744 38490
rect 11808 38282 11836 38916
rect 11888 38820 11940 38826
rect 11888 38762 11940 38768
rect 11796 38276 11848 38282
rect 11796 38218 11848 38224
rect 11808 38010 11836 38218
rect 11796 38004 11848 38010
rect 11796 37946 11848 37952
rect 11796 37800 11848 37806
rect 11796 37742 11848 37748
rect 11808 37398 11836 37742
rect 11796 37392 11848 37398
rect 11796 37334 11848 37340
rect 11704 37324 11756 37330
rect 11704 37266 11756 37272
rect 11900 37233 11928 38762
rect 11992 38758 12020 41386
rect 12176 41290 12204 42638
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 12256 42152 12308 42158
rect 12256 42094 12308 42100
rect 12084 41262 12204 41290
rect 12084 40390 12112 41262
rect 12164 41064 12216 41070
rect 12164 41006 12216 41012
rect 12072 40384 12124 40390
rect 12072 40326 12124 40332
rect 12084 39846 12112 40326
rect 12072 39840 12124 39846
rect 12072 39782 12124 39788
rect 12072 39568 12124 39574
rect 12072 39510 12124 39516
rect 11980 38752 12032 38758
rect 11980 38694 12032 38700
rect 12084 38654 12112 39510
rect 11992 38626 12112 38654
rect 11992 37448 12020 38626
rect 12072 38412 12124 38418
rect 12072 38354 12124 38360
rect 12084 37806 12112 38354
rect 12072 37800 12124 37806
rect 12072 37742 12124 37748
rect 11992 37420 12112 37448
rect 11978 37360 12034 37369
rect 11978 37295 11980 37304
rect 12032 37295 12034 37304
rect 11980 37266 12032 37272
rect 11886 37224 11942 37233
rect 11704 37188 11756 37194
rect 11886 37159 11942 37168
rect 11704 37130 11756 37136
rect 11716 36106 11744 37130
rect 11796 36916 11848 36922
rect 11796 36858 11848 36864
rect 11704 36100 11756 36106
rect 11704 36042 11756 36048
rect 11808 35986 11836 36858
rect 11980 36712 12032 36718
rect 12084 36700 12112 37420
rect 12032 36672 12112 36700
rect 11980 36654 12032 36660
rect 11992 36242 12020 36654
rect 12072 36576 12124 36582
rect 12072 36518 12124 36524
rect 11888 36236 11940 36242
rect 11888 36178 11940 36184
rect 11980 36236 12032 36242
rect 11980 36178 12032 36184
rect 11716 35958 11836 35986
rect 11716 35193 11744 35958
rect 11900 35834 11928 36178
rect 11888 35828 11940 35834
rect 11888 35770 11940 35776
rect 11888 35488 11940 35494
rect 11888 35430 11940 35436
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 11702 35184 11758 35193
rect 11702 35119 11758 35128
rect 11612 34468 11664 34474
rect 11612 34410 11664 34416
rect 11716 34354 11744 35119
rect 11808 34406 11836 35226
rect 11900 35086 11928 35430
rect 11992 35222 12020 36178
rect 12084 36174 12112 36518
rect 12176 36378 12204 41006
rect 12268 40050 12296 42094
rect 12348 40588 12400 40594
rect 12348 40530 12400 40536
rect 12256 40044 12308 40050
rect 12256 39986 12308 39992
rect 12360 39302 12388 40530
rect 12452 39370 12480 42502
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12544 40662 12572 41414
rect 12624 41132 12676 41138
rect 12624 41074 12676 41080
rect 12532 40656 12584 40662
rect 12532 40598 12584 40604
rect 12440 39364 12492 39370
rect 12440 39306 12492 39312
rect 12348 39296 12400 39302
rect 12348 39238 12400 39244
rect 12256 38752 12308 38758
rect 12256 38694 12308 38700
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 12176 36281 12204 36314
rect 12162 36272 12218 36281
rect 12162 36207 12218 36216
rect 12072 36168 12124 36174
rect 12072 36110 12124 36116
rect 12164 36032 12216 36038
rect 12164 35974 12216 35980
rect 12072 35488 12124 35494
rect 12072 35430 12124 35436
rect 11980 35216 12032 35222
rect 11980 35158 12032 35164
rect 11888 35080 11940 35086
rect 11888 35022 11940 35028
rect 11980 35012 12032 35018
rect 11980 34954 12032 34960
rect 11886 34640 11942 34649
rect 11886 34575 11942 34584
rect 11624 34326 11744 34354
rect 11796 34400 11848 34406
rect 11796 34342 11848 34348
rect 11336 33934 11388 33940
rect 11518 33960 11574 33969
rect 11348 32978 11376 33934
rect 11518 33895 11574 33904
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11336 32972 11388 32978
rect 11336 32914 11388 32920
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11348 30802 11376 32710
rect 11440 31657 11468 33798
rect 11624 32881 11652 34326
rect 11808 33946 11836 34342
rect 11900 34134 11928 34575
rect 11992 34542 12020 34954
rect 11980 34536 12032 34542
rect 11980 34478 12032 34484
rect 11980 34400 12032 34406
rect 11980 34342 12032 34348
rect 11888 34128 11940 34134
rect 11888 34070 11940 34076
rect 11716 33918 11836 33946
rect 11716 33862 11744 33918
rect 11704 33856 11756 33862
rect 11704 33798 11756 33804
rect 11796 33856 11848 33862
rect 11796 33798 11848 33804
rect 11610 32872 11666 32881
rect 11716 32842 11744 33798
rect 11610 32807 11666 32816
rect 11704 32836 11756 32842
rect 11624 32722 11652 32807
rect 11704 32778 11756 32784
rect 11624 32694 11744 32722
rect 11520 32224 11572 32230
rect 11520 32166 11572 32172
rect 11532 31754 11560 32166
rect 11612 31884 11664 31890
rect 11612 31826 11664 31832
rect 11520 31748 11572 31754
rect 11520 31690 11572 31696
rect 11426 31648 11482 31657
rect 11426 31583 11482 31592
rect 11428 31136 11480 31142
rect 11428 31078 11480 31084
rect 11336 30796 11388 30802
rect 11336 30738 11388 30744
rect 11440 30734 11468 31078
rect 11624 30938 11652 31826
rect 11612 30932 11664 30938
rect 11612 30874 11664 30880
rect 11716 30870 11744 32694
rect 11808 32434 11836 33798
rect 11886 33688 11942 33697
rect 11886 33623 11888 33632
rect 11940 33623 11942 33632
rect 11888 33594 11940 33600
rect 11900 32978 11928 33594
rect 11992 33561 12020 34342
rect 11978 33552 12034 33561
rect 11978 33487 12034 33496
rect 11980 33380 12032 33386
rect 11980 33322 12032 33328
rect 11888 32972 11940 32978
rect 11888 32914 11940 32920
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11794 32328 11850 32337
rect 11794 32263 11850 32272
rect 11808 31890 11836 32263
rect 11900 32230 11928 32914
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11886 32056 11942 32065
rect 11886 31991 11942 32000
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11794 31784 11850 31793
rect 11794 31719 11850 31728
rect 11704 30864 11756 30870
rect 11704 30806 11756 30812
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11440 30376 11468 30670
rect 11624 30394 11652 30738
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11348 30348 11468 30376
rect 11612 30388 11664 30394
rect 11348 29578 11376 30348
rect 11612 30330 11664 30336
rect 11426 30288 11482 30297
rect 11426 30223 11482 30232
rect 11336 29572 11388 29578
rect 11336 29514 11388 29520
rect 11334 29472 11390 29481
rect 11334 29407 11390 29416
rect 11348 29306 11376 29407
rect 11336 29300 11388 29306
rect 11336 29242 11388 29248
rect 11440 29102 11468 30223
rect 11520 30116 11572 30122
rect 11520 30058 11572 30064
rect 11532 29306 11560 30058
rect 11624 29714 11652 30330
rect 11716 30190 11744 30534
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11716 29782 11744 30126
rect 11704 29776 11756 29782
rect 11704 29718 11756 29724
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 11520 29300 11572 29306
rect 11520 29242 11572 29248
rect 11624 29102 11652 29446
rect 11244 29096 11296 29102
rect 11244 29038 11296 29044
rect 11428 29096 11480 29102
rect 11428 29038 11480 29044
rect 11612 29096 11664 29102
rect 11612 29038 11664 29044
rect 11164 28626 11284 28642
rect 11164 28620 11296 28626
rect 11164 28614 11244 28620
rect 11164 28150 11192 28614
rect 11244 28562 11296 28568
rect 11336 28416 11388 28422
rect 11336 28358 11388 28364
rect 11428 28416 11480 28422
rect 11428 28358 11480 28364
rect 11152 28144 11204 28150
rect 11152 28086 11204 28092
rect 11348 28014 11376 28358
rect 11440 28082 11468 28358
rect 11428 28076 11480 28082
rect 11428 28018 11480 28024
rect 11244 28008 11296 28014
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10062 27228 10370 27237
rect 10062 27226 10068 27228
rect 10124 27226 10148 27228
rect 10204 27226 10228 27228
rect 10284 27226 10308 27228
rect 10364 27226 10370 27228
rect 10124 27174 10126 27226
rect 10306 27174 10308 27226
rect 10062 27172 10068 27174
rect 10124 27172 10148 27174
rect 10204 27172 10228 27174
rect 10284 27172 10308 27174
rect 10364 27172 10370 27174
rect 10062 27163 10370 27172
rect 10062 26140 10370 26149
rect 10062 26138 10068 26140
rect 10124 26138 10148 26140
rect 10204 26138 10228 26140
rect 10284 26138 10308 26140
rect 10364 26138 10370 26140
rect 10124 26086 10126 26138
rect 10306 26086 10308 26138
rect 10062 26084 10068 26086
rect 10124 26084 10148 26086
rect 10204 26084 10228 26086
rect 10284 26084 10308 26086
rect 10364 26084 10370 26086
rect 10062 26075 10370 26084
rect 10428 26042 10456 27338
rect 10520 27130 10548 27950
rect 10980 27934 11100 27962
rect 11244 27950 11296 27956
rect 11336 28008 11388 28014
rect 11624 27962 11652 29038
rect 11716 28762 11744 29718
rect 11808 29034 11836 31719
rect 11900 30841 11928 31991
rect 11886 30832 11942 30841
rect 11886 30767 11942 30776
rect 11900 30734 11928 30767
rect 11888 30728 11940 30734
rect 11888 30670 11940 30676
rect 11888 30592 11940 30598
rect 11888 30534 11940 30540
rect 11900 29850 11928 30534
rect 11888 29844 11940 29850
rect 11888 29786 11940 29792
rect 11992 29306 12020 33322
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 11796 29028 11848 29034
rect 11796 28970 11848 28976
rect 12084 28762 12112 35430
rect 12176 35290 12204 35974
rect 12164 35284 12216 35290
rect 12164 35226 12216 35232
rect 12268 35222 12296 38694
rect 12360 37777 12388 39238
rect 12346 37768 12402 37777
rect 12346 37703 12402 37712
rect 12256 35216 12308 35222
rect 12256 35158 12308 35164
rect 12256 34536 12308 34542
rect 12256 34478 12308 34484
rect 12164 33312 12216 33318
rect 12164 33254 12216 33260
rect 12176 32910 12204 33254
rect 12268 33046 12296 34478
rect 12256 33040 12308 33046
rect 12256 32982 12308 32988
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 12268 32366 12296 32982
rect 12256 32360 12308 32366
rect 12256 32302 12308 32308
rect 12164 32224 12216 32230
rect 12164 32166 12216 32172
rect 11704 28756 11756 28762
rect 11704 28698 11756 28704
rect 11980 28756 12032 28762
rect 11980 28698 12032 28704
rect 12072 28756 12124 28762
rect 12072 28698 12124 28704
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11704 28212 11756 28218
rect 11704 28154 11756 28160
rect 11336 27950 11388 27956
rect 10600 27872 10652 27878
rect 10600 27814 10652 27820
rect 10612 27606 10640 27814
rect 10722 27772 11030 27781
rect 10722 27770 10728 27772
rect 10784 27770 10808 27772
rect 10864 27770 10888 27772
rect 10944 27770 10968 27772
rect 11024 27770 11030 27772
rect 10784 27718 10786 27770
rect 10966 27718 10968 27770
rect 10722 27716 10728 27718
rect 10784 27716 10808 27718
rect 10864 27716 10888 27718
rect 10944 27716 10968 27718
rect 11024 27716 11030 27718
rect 10722 27707 11030 27716
rect 10600 27600 10652 27606
rect 11072 27554 11100 27934
rect 10600 27542 10652 27548
rect 10980 27526 11100 27554
rect 11256 27538 11284 27950
rect 11440 27934 11652 27962
rect 11152 27532 11204 27538
rect 10508 27124 10560 27130
rect 10508 27066 10560 27072
rect 10508 26852 10560 26858
rect 10508 26794 10560 26800
rect 10520 26586 10548 26794
rect 10980 26772 11008 27526
rect 11152 27474 11204 27480
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11072 26926 11100 27406
rect 11164 26926 11192 27474
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 11152 26920 11204 26926
rect 11152 26862 11204 26868
rect 11336 26784 11388 26790
rect 10980 26744 11100 26772
rect 10722 26684 11030 26693
rect 10722 26682 10728 26684
rect 10784 26682 10808 26684
rect 10864 26682 10888 26684
rect 10944 26682 10968 26684
rect 11024 26682 11030 26684
rect 10784 26630 10786 26682
rect 10966 26630 10968 26682
rect 10722 26628 10728 26630
rect 10784 26628 10808 26630
rect 10864 26628 10888 26630
rect 10944 26628 10968 26630
rect 11024 26628 11030 26630
rect 10722 26619 11030 26628
rect 10508 26580 10560 26586
rect 10508 26522 10560 26528
rect 11072 26228 11100 26744
rect 11336 26726 11388 26732
rect 11072 26200 11192 26228
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10508 25832 10560 25838
rect 10508 25774 10560 25780
rect 11060 25832 11112 25838
rect 11060 25774 11112 25780
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 9968 25452 10364 25480
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9968 24954 9996 25298
rect 10336 25208 10364 25452
rect 10428 25430 10456 25638
rect 10520 25498 10548 25774
rect 10600 25764 10652 25770
rect 10600 25706 10652 25712
rect 10508 25492 10560 25498
rect 10508 25434 10560 25440
rect 10416 25424 10468 25430
rect 10416 25366 10468 25372
rect 10612 25362 10640 25706
rect 10722 25596 11030 25605
rect 10722 25594 10728 25596
rect 10784 25594 10808 25596
rect 10864 25594 10888 25596
rect 10944 25594 10968 25596
rect 11024 25594 11030 25596
rect 10784 25542 10786 25594
rect 10966 25542 10968 25594
rect 10722 25540 10728 25542
rect 10784 25540 10808 25542
rect 10864 25540 10888 25542
rect 10944 25540 10968 25542
rect 11024 25540 11030 25542
rect 10722 25531 11030 25540
rect 10600 25356 10652 25362
rect 10600 25298 10652 25304
rect 10508 25288 10560 25294
rect 10508 25230 10560 25236
rect 10336 25180 10456 25208
rect 10062 25052 10370 25061
rect 10062 25050 10068 25052
rect 10124 25050 10148 25052
rect 10204 25050 10228 25052
rect 10284 25050 10308 25052
rect 10364 25050 10370 25052
rect 10124 24998 10126 25050
rect 10306 24998 10308 25050
rect 10062 24996 10068 24998
rect 10124 24996 10148 24998
rect 10204 24996 10228 24998
rect 10284 24996 10308 24998
rect 10364 24996 10370 24998
rect 10062 24987 10370 24996
rect 9956 24948 10008 24954
rect 9956 24890 10008 24896
rect 9864 24880 9916 24886
rect 9864 24822 9916 24828
rect 9864 24744 9916 24750
rect 9784 24704 9864 24732
rect 9864 24686 9916 24692
rect 9864 24608 9916 24614
rect 9770 24576 9826 24585
rect 9864 24550 9916 24556
rect 9770 24511 9826 24520
rect 9784 23633 9812 24511
rect 9876 24070 9904 24550
rect 9968 24274 9996 24890
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 9956 24268 10008 24274
rect 9956 24210 10008 24216
rect 10060 24154 10088 24822
rect 10324 24812 10376 24818
rect 10324 24754 10376 24760
rect 10336 24274 10364 24754
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 9968 24126 10088 24154
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9770 23624 9826 23633
rect 9770 23559 9826 23568
rect 9678 23488 9734 23497
rect 9678 23423 9734 23432
rect 9876 23202 9904 24006
rect 9784 23174 9904 23202
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9600 22778 9628 23054
rect 9680 22976 9732 22982
rect 9680 22918 9732 22924
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9600 22438 9628 22510
rect 9588 22432 9640 22438
rect 9588 22374 9640 22380
rect 9600 21622 9628 22374
rect 9588 21616 9640 21622
rect 9588 21558 9640 21564
rect 9692 21486 9720 22918
rect 9784 22624 9812 23174
rect 9968 22681 9996 24126
rect 10062 23964 10370 23973
rect 10062 23962 10068 23964
rect 10124 23962 10148 23964
rect 10204 23962 10228 23964
rect 10284 23962 10308 23964
rect 10364 23962 10370 23964
rect 10124 23910 10126 23962
rect 10306 23910 10308 23962
rect 10062 23908 10068 23910
rect 10124 23908 10148 23910
rect 10204 23908 10228 23910
rect 10284 23908 10308 23910
rect 10364 23908 10370 23910
rect 10062 23899 10370 23908
rect 10324 23656 10376 23662
rect 10324 23598 10376 23604
rect 10336 23186 10364 23598
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10428 23089 10456 25180
rect 10520 23866 10548 25230
rect 10692 24812 10744 24818
rect 10612 24772 10692 24800
rect 10612 24342 10640 24772
rect 10692 24754 10744 24760
rect 10722 24508 11030 24517
rect 10722 24506 10728 24508
rect 10784 24506 10808 24508
rect 10864 24506 10888 24508
rect 10944 24506 10968 24508
rect 11024 24506 11030 24508
rect 10784 24454 10786 24506
rect 10966 24454 10968 24506
rect 10722 24452 10728 24454
rect 10784 24452 10808 24454
rect 10864 24452 10888 24454
rect 10944 24452 10968 24454
rect 11024 24452 11030 24454
rect 10722 24443 11030 24452
rect 10600 24336 10652 24342
rect 10600 24278 10652 24284
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10612 23798 10640 24278
rect 11072 24274 11100 25774
rect 11060 24268 11112 24274
rect 11060 24210 11112 24216
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10600 23792 10652 23798
rect 10600 23734 10652 23740
rect 10612 23304 10640 23734
rect 10704 23662 10732 24074
rect 10692 23656 10744 23662
rect 10692 23598 10744 23604
rect 11072 23526 11100 24210
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10722 23420 11030 23429
rect 10722 23418 10728 23420
rect 10784 23418 10808 23420
rect 10864 23418 10888 23420
rect 10944 23418 10968 23420
rect 11024 23418 11030 23420
rect 10784 23366 10786 23418
rect 10966 23366 10968 23418
rect 10722 23364 10728 23366
rect 10784 23364 10808 23366
rect 10864 23364 10888 23366
rect 10944 23364 10968 23366
rect 11024 23364 11030 23366
rect 10722 23355 11030 23364
rect 10612 23276 10916 23304
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10414 23080 10470 23089
rect 10414 23015 10470 23024
rect 10508 23044 10560 23050
rect 10508 22986 10560 22992
rect 10416 22976 10468 22982
rect 10416 22918 10468 22924
rect 10062 22876 10370 22885
rect 10062 22874 10068 22876
rect 10124 22874 10148 22876
rect 10204 22874 10228 22876
rect 10284 22874 10308 22876
rect 10364 22874 10370 22876
rect 10124 22822 10126 22874
rect 10306 22822 10308 22874
rect 10062 22820 10068 22822
rect 10124 22820 10148 22822
rect 10204 22820 10228 22822
rect 10284 22820 10308 22822
rect 10364 22820 10370 22822
rect 10062 22811 10370 22820
rect 9954 22672 10010 22681
rect 9784 22596 9904 22624
rect 9954 22607 10010 22616
rect 10138 22672 10194 22681
rect 10138 22607 10140 22616
rect 9876 22386 9904 22596
rect 10192 22607 10194 22616
rect 10140 22578 10192 22584
rect 9956 22568 10008 22574
rect 10008 22528 10088 22556
rect 9956 22510 10008 22516
rect 9876 22358 9996 22386
rect 9968 22234 9996 22358
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9600 21298 9628 21422
rect 9876 21418 9904 22170
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9968 21622 9996 22034
rect 10060 21894 10088 22528
rect 10048 21888 10100 21894
rect 10152 21876 10180 22578
rect 10428 22166 10456 22918
rect 10416 22160 10468 22166
rect 10416 22102 10468 22108
rect 10520 22098 10548 22986
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10612 22710 10640 22918
rect 10600 22704 10652 22710
rect 10600 22646 10652 22652
rect 10704 22522 10732 23122
rect 10888 22642 10916 23276
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10980 22778 11008 23122
rect 10968 22772 11020 22778
rect 10968 22714 11020 22720
rect 10876 22636 10928 22642
rect 10928 22596 11100 22624
rect 10876 22578 10928 22584
rect 10784 22568 10836 22574
rect 10612 22494 10732 22522
rect 10782 22536 10784 22545
rect 10836 22536 10838 22545
rect 10612 22234 10640 22494
rect 10782 22471 10838 22480
rect 10722 22332 11030 22341
rect 10722 22330 10728 22332
rect 10784 22330 10808 22332
rect 10864 22330 10888 22332
rect 10944 22330 10968 22332
rect 11024 22330 11030 22332
rect 10784 22278 10786 22330
rect 10966 22278 10968 22330
rect 10722 22276 10728 22278
rect 10784 22276 10808 22278
rect 10864 22276 10888 22278
rect 10944 22276 10968 22278
rect 11024 22276 11030 22278
rect 10722 22267 11030 22276
rect 10600 22228 10652 22234
rect 11072 22216 11100 22596
rect 10600 22170 10652 22176
rect 10888 22188 11100 22216
rect 10508 22092 10560 22098
rect 10508 22034 10560 22040
rect 10692 22092 10744 22098
rect 10692 22034 10744 22040
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10508 21888 10560 21894
rect 10152 21848 10456 21876
rect 10048 21830 10100 21836
rect 10062 21788 10370 21797
rect 10062 21786 10068 21788
rect 10124 21786 10148 21788
rect 10204 21786 10228 21788
rect 10284 21786 10308 21788
rect 10364 21786 10370 21788
rect 10124 21734 10126 21786
rect 10306 21734 10308 21786
rect 10062 21732 10068 21734
rect 10124 21732 10148 21734
rect 10204 21732 10228 21734
rect 10284 21732 10308 21734
rect 10364 21732 10370 21734
rect 10062 21723 10370 21732
rect 9956 21616 10008 21622
rect 9956 21558 10008 21564
rect 10048 21616 10100 21622
rect 10048 21558 10100 21564
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9600 21270 9720 21298
rect 9494 20768 9550 20777
rect 9494 20703 9550 20712
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9312 20528 9364 20534
rect 9126 20496 9182 20505
rect 9312 20470 9364 20476
rect 9126 20431 9182 20440
rect 9140 20398 9168 20431
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9404 20324 9456 20330
rect 9404 20266 9456 20272
rect 9220 20256 9272 20262
rect 9272 20216 9352 20244
rect 9220 20198 9272 20204
rect 9218 20088 9274 20097
rect 9218 20023 9274 20032
rect 9128 19916 9180 19922
rect 9128 19858 9180 19864
rect 9036 19848 9088 19854
rect 9036 19790 9088 19796
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9048 19281 9076 19654
rect 9140 19378 9168 19858
rect 9128 19372 9180 19378
rect 9128 19314 9180 19320
rect 9034 19272 9090 19281
rect 9034 19207 9090 19216
rect 9128 19236 9180 19242
rect 9128 19178 9180 19184
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9140 18902 9168 19178
rect 8668 18896 8720 18902
rect 8668 18838 8720 18844
rect 9128 18896 9180 18902
rect 9128 18838 9180 18844
rect 8680 18222 8708 18838
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8944 18216 8996 18222
rect 8944 18158 8996 18164
rect 8574 18048 8630 18057
rect 8574 17983 8630 17992
rect 8574 17912 8630 17921
rect 8574 17847 8630 17856
rect 8758 17912 8814 17921
rect 8758 17847 8814 17856
rect 8588 17746 8616 17847
rect 8772 17814 8800 17847
rect 8760 17808 8812 17814
rect 8680 17768 8760 17796
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8588 16658 8616 17682
rect 8680 16658 8708 17768
rect 8760 17750 8812 17756
rect 8850 17640 8906 17649
rect 8850 17575 8906 17584
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8680 16182 8708 16594
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8404 16102 8524 16130
rect 8668 16176 8720 16182
rect 8668 16118 8720 16124
rect 8206 15600 8262 15609
rect 8206 15535 8208 15544
rect 8260 15535 8262 15544
rect 8208 15506 8260 15512
rect 8312 14890 8340 16050
rect 8404 15162 8432 16102
rect 8772 16046 8800 17478
rect 8864 17134 8892 17575
rect 8852 17128 8904 17134
rect 8852 17070 8904 17076
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8760 16040 8812 16046
rect 8760 15982 8812 15988
rect 8496 15706 8524 15982
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8588 15434 8616 15506
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8482 15328 8538 15337
rect 8482 15263 8538 15272
rect 8392 15156 8444 15162
rect 8392 15098 8444 15104
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8300 14884 8352 14890
rect 8300 14826 8352 14832
rect 8404 14550 8432 14962
rect 8496 14618 8524 15263
rect 8680 15162 8708 15642
rect 8772 15502 8800 15982
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8392 14544 8444 14550
rect 8392 14486 8444 14492
rect 8116 14476 8168 14482
rect 8484 14476 8536 14482
rect 8168 14436 8248 14464
rect 8116 14418 8168 14424
rect 7932 14340 7984 14346
rect 7932 14282 7984 14288
rect 7932 14000 7984 14006
rect 7932 13942 7984 13948
rect 7944 13818 7972 13942
rect 7944 13790 8064 13818
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7944 12782 7972 12922
rect 7932 12776 7984 12782
rect 7932 12718 7984 12724
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7654 12472 7710 12481
rect 7654 12407 7710 12416
rect 7654 12336 7710 12345
rect 7654 12271 7656 12280
rect 7708 12271 7710 12280
rect 7656 12242 7708 12248
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11898 7696 12038
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7576 11750 7788 11778
rect 7392 11354 7420 11750
rect 7472 11688 7524 11694
rect 7472 11630 7524 11636
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7300 9674 7328 11290
rect 7484 11286 7512 11630
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10606 7420 11086
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7300 9646 7420 9674
rect 7288 9512 7340 9518
rect 7288 9454 7340 9460
rect 7300 9382 7328 9454
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 9178 7328 9318
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7300 8430 7328 8842
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7392 8090 7420 9646
rect 7484 8956 7512 11222
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 10606 7696 11018
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7576 9110 7604 10066
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7668 9654 7696 9998
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7564 9104 7616 9110
rect 7564 9046 7616 9052
rect 7468 8928 7512 8956
rect 7468 8888 7496 8928
rect 7468 8860 7512 8888
rect 7484 8401 7512 8860
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7470 8392 7526 8401
rect 7470 8327 7526 8336
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7024 7398 7144 7426
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6564 6254 6592 7278
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 6798 6960 7142
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6840 6458 6868 6734
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6932 6338 6960 6734
rect 7024 6458 7052 6734
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6932 6310 7052 6338
rect 7024 6254 7052 6310
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6460 4820 6512 4826
rect 6460 4762 6512 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6104 4078 6132 4694
rect 6564 4214 6592 6190
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6840 4690 6868 5102
rect 7116 5030 7144 7398
rect 7196 7336 7248 7342
rect 7196 7278 7248 7284
rect 7208 6458 7236 7278
rect 7300 7002 7328 7890
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7300 6254 7328 6938
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 7288 6248 7340 6254
rect 7288 6190 7340 6196
rect 7208 6100 7236 6190
rect 7392 6100 7420 7890
rect 7484 7410 7512 8327
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7208 6072 7420 6100
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6828 4684 6880 4690
rect 6828 4626 6880 4632
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6748 3670 6776 4626
rect 6840 3738 6868 4626
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 3738 7052 4082
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 6736 3664 6788 3670
rect 6736 3606 6788 3612
rect 6840 3602 6868 3674
rect 6828 3596 6880 3602
rect 6828 3538 6880 3544
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6276 2304 6328 2310
rect 6276 2246 6328 2252
rect 5908 1828 5960 1834
rect 5908 1770 5960 1776
rect 5460 1426 5856 1442
rect 4896 1420 4948 1426
rect 4896 1362 4948 1368
rect 5448 1420 5856 1426
rect 5500 1414 5856 1420
rect 5448 1362 5500 1368
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 5552 882 5580 1414
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 5540 876 5592 882
rect 5540 818 5592 824
rect 6104 814 6132 1158
rect 6288 814 6316 2246
rect 6380 1902 6408 2926
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6368 1896 6420 1902
rect 6368 1838 6420 1844
rect 6472 1426 6500 2450
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6564 1494 6592 2382
rect 6656 1902 6684 2926
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6552 1488 6604 1494
rect 6552 1430 6604 1436
rect 6460 1420 6512 1426
rect 6460 1362 6512 1368
rect 6472 1018 6500 1362
rect 6656 1018 6684 1838
rect 6748 1426 6776 2790
rect 7208 2774 7236 6072
rect 7300 5222 7512 5250
rect 7300 5166 7328 5222
rect 7484 5166 7512 5222
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7024 2746 7236 2774
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6840 1358 6868 1702
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 7024 1222 7052 2746
rect 7300 2650 7328 5102
rect 7392 4282 7420 5102
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7484 4078 7512 4422
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7392 2774 7420 3538
rect 7484 3534 7512 4014
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7576 2774 7604 8434
rect 7760 5386 7788 11750
rect 7852 11558 7880 12582
rect 7932 12368 7984 12374
rect 7932 12310 7984 12316
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7944 11336 7972 12310
rect 8036 11694 8064 13790
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12782 8156 13126
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8220 12442 8248 14436
rect 8484 14418 8536 14424
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 8312 12322 8340 12718
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8220 12294 8340 12322
rect 8404 12306 8432 14350
rect 8392 12300 8444 12306
rect 8128 12073 8156 12242
rect 8114 12064 8170 12073
rect 8114 11999 8170 12008
rect 8220 11762 8248 12294
rect 8392 12242 8444 12248
rect 8496 12186 8524 14418
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8312 12158 8524 12186
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7852 11308 7972 11336
rect 7852 10674 7880 11308
rect 7932 11212 7984 11218
rect 8036 11200 8064 11630
rect 8208 11620 8260 11626
rect 8208 11562 8260 11568
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 11218 8156 11494
rect 8220 11354 8248 11562
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 7984 11172 8064 11200
rect 8116 11212 8168 11218
rect 7932 11154 7984 11160
rect 8116 11154 8168 11160
rect 8114 11112 8170 11121
rect 8114 11047 8170 11056
rect 8128 10810 8156 11047
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 7840 10668 7892 10674
rect 7840 10610 7892 10616
rect 7932 10192 7984 10198
rect 7932 10134 7984 10140
rect 7944 9382 7972 10134
rect 8220 9586 8248 11290
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8220 8906 8248 9522
rect 8312 8922 8340 12158
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8404 11762 8432 12038
rect 8496 11762 8524 12038
rect 8588 11898 8616 13398
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12481 8708 12786
rect 8666 12472 8722 12481
rect 8666 12407 8722 12416
rect 8680 11898 8708 12407
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8588 10266 8616 11630
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8404 9518 8432 9998
rect 8392 9512 8444 9518
rect 8392 9454 8444 9460
rect 8496 9110 8524 10066
rect 8772 9110 8800 14214
rect 8864 12306 8892 16934
rect 8956 16658 8984 18158
rect 9048 17882 9076 18566
rect 9232 18358 9260 20023
rect 9324 19922 9352 20216
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9312 19780 9364 19786
rect 9312 19722 9364 19728
rect 9324 19310 9352 19722
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9416 18902 9444 20266
rect 9508 18970 9536 20538
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9600 19378 9628 20402
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 18970 9628 19178
rect 9496 18964 9548 18970
rect 9496 18906 9548 18912
rect 9588 18964 9640 18970
rect 9588 18906 9640 18912
rect 9312 18896 9364 18902
rect 9312 18838 9364 18844
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9508 18850 9536 18906
rect 9220 18352 9272 18358
rect 9220 18294 9272 18300
rect 9232 18222 9260 18294
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 9140 17882 9168 18090
rect 9036 17876 9088 17882
rect 9036 17818 9088 17824
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9048 16658 9076 17818
rect 9126 17776 9182 17785
rect 9126 17711 9128 17720
rect 9180 17711 9182 17720
rect 9324 17728 9352 18838
rect 9508 18822 9628 18850
rect 9404 18760 9456 18766
rect 9456 18720 9536 18748
rect 9404 18702 9456 18708
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 17921 9444 18158
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9404 17740 9456 17746
rect 9324 17700 9404 17728
rect 9128 17682 9180 17688
rect 9404 17682 9456 17688
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9126 17368 9182 17377
rect 9126 17303 9128 17312
rect 9180 17303 9182 17312
rect 9128 17274 9180 17280
rect 8944 16652 8996 16658
rect 8944 16594 8996 16600
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 8956 15570 8984 16594
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8956 15065 8984 15506
rect 8942 15056 8998 15065
rect 8942 14991 8998 15000
rect 8956 14550 8984 14991
rect 8944 14544 8996 14550
rect 8944 14486 8996 14492
rect 9048 14498 9076 16594
rect 9232 15026 9260 17478
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9324 16697 9352 16934
rect 9310 16688 9366 16697
rect 9310 16623 9366 16632
rect 9416 16590 9444 17682
rect 9404 16584 9456 16590
rect 9404 16526 9456 16532
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9324 15178 9352 15982
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9416 15570 9444 15846
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9416 15366 9444 15506
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9324 15150 9444 15178
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9140 14618 9168 14758
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 9048 14470 9168 14498
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 8956 13802 8984 14350
rect 9048 14278 9076 14350
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 8942 12880 8998 12889
rect 8942 12815 8998 12824
rect 8956 12782 8984 12815
rect 9140 12782 9168 14470
rect 9232 13530 9260 14962
rect 9310 14512 9366 14521
rect 9310 14447 9366 14456
rect 9324 14414 9352 14447
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9324 13410 9352 14350
rect 9416 13802 9444 15150
rect 9508 14414 9536 18720
rect 9600 17898 9628 18822
rect 9692 18698 9720 21270
rect 9772 21072 9824 21078
rect 9772 21014 9824 21020
rect 9784 19514 9812 21014
rect 9876 20602 9904 21354
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 18970 9812 19246
rect 9876 18970 9904 20198
rect 9968 19378 9996 21082
rect 10060 21078 10088 21558
rect 10428 21486 10456 21848
rect 10508 21830 10560 21836
rect 10520 21554 10548 21830
rect 10612 21690 10640 21898
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10704 21570 10732 22034
rect 10888 21690 10916 22188
rect 11058 22128 11114 22137
rect 11058 22063 11114 22072
rect 10968 21888 11020 21894
rect 10968 21830 11020 21836
rect 10876 21684 10928 21690
rect 10876 21626 10928 21632
rect 10508 21548 10560 21554
rect 10508 21490 10560 21496
rect 10612 21542 10732 21570
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10508 21412 10560 21418
rect 10508 21354 10560 21360
rect 10414 21312 10470 21321
rect 10414 21247 10470 21256
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 10062 20700 10370 20709
rect 10062 20698 10068 20700
rect 10124 20698 10148 20700
rect 10204 20698 10228 20700
rect 10284 20698 10308 20700
rect 10364 20698 10370 20700
rect 10124 20646 10126 20698
rect 10306 20646 10308 20698
rect 10062 20644 10068 20646
rect 10124 20644 10148 20646
rect 10204 20644 10228 20646
rect 10284 20644 10308 20646
rect 10364 20644 10370 20646
rect 10062 20635 10370 20644
rect 10428 20330 10456 21247
rect 10520 21010 10548 21354
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10520 20398 10548 20946
rect 10508 20392 10560 20398
rect 10508 20334 10560 20340
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10612 20058 10640 21542
rect 10980 21350 11008 21830
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10722 21244 11030 21253
rect 10722 21242 10728 21244
rect 10784 21242 10808 21244
rect 10864 21242 10888 21244
rect 10944 21242 10968 21244
rect 11024 21242 11030 21244
rect 10784 21190 10786 21242
rect 10966 21190 10968 21242
rect 10722 21188 10728 21190
rect 10784 21188 10808 21190
rect 10864 21188 10888 21190
rect 10944 21188 10968 21190
rect 11024 21188 11030 21190
rect 10722 21179 11030 21188
rect 11072 21128 11100 22063
rect 11164 21962 11192 26200
rect 11244 25696 11296 25702
rect 11244 25638 11296 25644
rect 11256 25294 11284 25638
rect 11244 25288 11296 25294
rect 11244 25230 11296 25236
rect 11348 25106 11376 26726
rect 11440 26353 11468 27934
rect 11716 27538 11744 28154
rect 11900 28014 11928 28494
rect 11888 28008 11940 28014
rect 11888 27950 11940 27956
rect 11796 27872 11848 27878
rect 11796 27814 11848 27820
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 11426 26344 11482 26353
rect 11426 26279 11482 26288
rect 11428 25764 11480 25770
rect 11428 25706 11480 25712
rect 11256 25078 11376 25106
rect 11256 24342 11284 25078
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11244 24336 11296 24342
rect 11244 24278 11296 24284
rect 11348 24206 11376 24686
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11440 24154 11468 25706
rect 11532 25226 11560 27406
rect 11624 26994 11652 27406
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11716 26994 11744 27270
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11624 25480 11652 26930
rect 11808 26926 11836 27814
rect 11900 27674 11928 27950
rect 11888 27668 11940 27674
rect 11888 27610 11940 27616
rect 11888 27532 11940 27538
rect 11888 27474 11940 27480
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11900 26586 11928 27474
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11900 25888 11928 26522
rect 11808 25860 11928 25888
rect 11808 25702 11836 25860
rect 11992 25820 12020 28698
rect 12070 28656 12126 28665
rect 12070 28591 12072 28600
rect 12124 28591 12126 28600
rect 12072 28562 12124 28568
rect 12072 28484 12124 28490
rect 12072 28426 12124 28432
rect 12084 28014 12112 28426
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 12084 27130 12112 27950
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12176 26874 12204 32166
rect 12268 31686 12296 32302
rect 12360 32065 12388 37703
rect 12346 32056 12402 32065
rect 12346 31991 12402 32000
rect 12348 31748 12400 31754
rect 12348 31690 12400 31696
rect 12256 31680 12308 31686
rect 12256 31622 12308 31628
rect 12268 30258 12296 31622
rect 12360 30734 12388 31690
rect 12348 30728 12400 30734
rect 12348 30670 12400 30676
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12268 29646 12296 29990
rect 12256 29640 12308 29646
rect 12256 29582 12308 29588
rect 12452 28626 12480 39306
rect 12636 37942 12664 41074
rect 12716 38344 12768 38350
rect 12716 38286 12768 38292
rect 12624 37936 12676 37942
rect 12624 37878 12676 37884
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12544 34514 12572 37198
rect 12636 36038 12664 37878
rect 12728 37126 12756 38286
rect 12716 37120 12768 37126
rect 12716 37062 12768 37068
rect 12716 36100 12768 36106
rect 12716 36042 12768 36048
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12544 34486 12664 34514
rect 12532 33448 12584 33454
rect 12532 33390 12584 33396
rect 12544 31822 12572 33390
rect 12636 31929 12664 34486
rect 12728 33114 12756 36042
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12622 31920 12678 31929
rect 12622 31855 12678 31864
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12544 29170 12572 31758
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12636 29617 12664 30670
rect 12622 29608 12678 29617
rect 12622 29543 12678 29552
rect 12532 29164 12584 29170
rect 12532 29106 12584 29112
rect 12440 28620 12492 28626
rect 12440 28562 12492 28568
rect 12256 27872 12308 27878
rect 12256 27814 12308 27820
rect 12268 27713 12296 27814
rect 12254 27704 12310 27713
rect 12254 27639 12310 27648
rect 12176 26846 12296 26874
rect 11900 25792 12020 25820
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11624 25452 11836 25480
rect 11612 25356 11664 25362
rect 11612 25298 11664 25304
rect 11520 25220 11572 25226
rect 11520 25162 11572 25168
rect 11532 24750 11560 25162
rect 11624 24818 11652 25298
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11716 24886 11744 25230
rect 11704 24880 11756 24886
rect 11704 24822 11756 24828
rect 11612 24812 11664 24818
rect 11612 24754 11664 24760
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11624 24274 11652 24754
rect 11704 24608 11756 24614
rect 11704 24550 11756 24556
rect 11612 24268 11664 24274
rect 11612 24210 11664 24216
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11256 23322 11284 23666
rect 11348 23662 11376 24142
rect 11440 24126 11652 24154
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11336 23656 11388 23662
rect 11336 23598 11388 23604
rect 11440 23497 11468 24006
rect 11520 23860 11572 23866
rect 11520 23802 11572 23808
rect 11532 23594 11560 23802
rect 11520 23588 11572 23594
rect 11520 23530 11572 23536
rect 11426 23488 11482 23497
rect 11426 23423 11482 23432
rect 11244 23316 11296 23322
rect 11428 23316 11480 23322
rect 11296 23276 11376 23304
rect 11244 23258 11296 23264
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11256 22506 11284 23054
rect 11348 22574 11376 23276
rect 11428 23258 11480 23264
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11244 22500 11296 22506
rect 11244 22442 11296 22448
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11348 22030 11376 22374
rect 11440 22098 11468 23258
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11532 22234 11560 23122
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11624 22137 11652 24126
rect 11716 23497 11744 24550
rect 11808 23798 11836 25452
rect 11900 24410 11928 25792
rect 12072 25764 12124 25770
rect 12072 25706 12124 25712
rect 11980 25696 12032 25702
rect 11980 25638 12032 25644
rect 11992 24750 12020 25638
rect 12084 25362 12112 25706
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11992 24290 12020 24686
rect 11900 24262 12020 24290
rect 12084 24274 12112 25298
rect 12176 24818 12204 25638
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12072 24268 12124 24274
rect 11900 24070 11928 24262
rect 12072 24210 12124 24216
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 11888 24064 11940 24070
rect 11888 24006 11940 24012
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11702 23488 11758 23497
rect 11702 23423 11758 23432
rect 11808 23322 11836 23734
rect 11796 23316 11848 23322
rect 11796 23258 11848 23264
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11704 22976 11756 22982
rect 11704 22918 11756 22924
rect 11610 22128 11666 22137
rect 11428 22092 11480 22098
rect 11610 22063 11666 22072
rect 11428 22034 11480 22040
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11152 21956 11204 21962
rect 11152 21898 11204 21904
rect 11348 21298 11376 21966
rect 11716 21962 11744 22918
rect 11808 22778 11836 23122
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11704 21956 11756 21962
rect 11704 21898 11756 21904
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11348 21270 11468 21298
rect 11072 21100 11284 21128
rect 11152 21004 11204 21010
rect 11152 20946 11204 20952
rect 10690 20904 10746 20913
rect 10690 20839 10746 20848
rect 10704 20330 10732 20839
rect 11060 20800 11112 20806
rect 11060 20742 11112 20748
rect 10692 20324 10744 20330
rect 10692 20266 10744 20272
rect 10722 20156 11030 20165
rect 10722 20154 10728 20156
rect 10784 20154 10808 20156
rect 10864 20154 10888 20156
rect 10944 20154 10968 20156
rect 11024 20154 11030 20156
rect 10784 20102 10786 20154
rect 10966 20102 10968 20154
rect 10722 20100 10728 20102
rect 10784 20100 10808 20102
rect 10864 20100 10888 20102
rect 10944 20100 10968 20102
rect 11024 20100 11030 20102
rect 10722 20091 11030 20100
rect 10600 20052 10652 20058
rect 10600 19994 10652 20000
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 10876 19984 10928 19990
rect 10874 19952 10876 19961
rect 10928 19952 10930 19961
rect 10600 19916 10652 19922
rect 10652 19876 10732 19904
rect 10874 19887 10930 19896
rect 10600 19858 10652 19864
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10062 19612 10370 19621
rect 10062 19610 10068 19612
rect 10124 19610 10148 19612
rect 10204 19610 10228 19612
rect 10284 19610 10308 19612
rect 10364 19610 10370 19612
rect 10124 19558 10126 19610
rect 10306 19558 10308 19610
rect 10062 19556 10068 19558
rect 10124 19556 10148 19558
rect 10204 19556 10228 19558
rect 10284 19556 10308 19558
rect 10364 19556 10370 19558
rect 10062 19547 10370 19556
rect 10428 19514 10456 19654
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10060 18834 10088 19450
rect 10520 19310 10548 19654
rect 10612 19310 10640 19722
rect 10704 19689 10732 19876
rect 10980 19802 11008 19994
rect 11072 19922 11100 20742
rect 11164 20602 11192 20946
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11164 19922 11192 20538
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 10980 19774 11100 19802
rect 11072 19718 11100 19774
rect 10968 19712 11020 19718
rect 10690 19680 10746 19689
rect 10690 19615 10746 19624
rect 10966 19680 10968 19689
rect 11060 19712 11112 19718
rect 11020 19680 11022 19689
rect 11060 19654 11112 19660
rect 10966 19615 11022 19624
rect 11256 19310 11284 21100
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11348 20058 11376 20946
rect 11440 20874 11468 21270
rect 11532 21010 11560 21626
rect 11716 21350 11744 21898
rect 11704 21344 11756 21350
rect 11704 21286 11756 21292
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11612 21004 11664 21010
rect 11612 20946 11664 20952
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11440 19922 11468 20810
rect 11428 19916 11480 19922
rect 11428 19858 11480 19864
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 10722 19068 11030 19077
rect 10722 19066 10728 19068
rect 10784 19066 10808 19068
rect 10864 19066 10888 19068
rect 10944 19066 10968 19068
rect 11024 19066 11030 19068
rect 10784 19014 10786 19066
rect 10966 19014 10968 19066
rect 10722 19012 10728 19014
rect 10784 19012 10808 19014
rect 10864 19012 10888 19014
rect 10944 19012 10968 19014
rect 11024 19012 11030 19014
rect 10722 19003 11030 19012
rect 9864 18828 9916 18834
rect 10048 18828 10100 18834
rect 9916 18788 10048 18816
rect 9864 18770 9916 18776
rect 9680 18692 9732 18698
rect 9680 18634 9732 18640
rect 9772 18352 9824 18358
rect 9772 18294 9824 18300
rect 9600 17870 9720 17898
rect 9588 17740 9640 17746
rect 9588 17682 9640 17688
rect 9600 16794 9628 17682
rect 9692 17270 9720 17870
rect 9784 17814 9812 18294
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9784 17542 9812 17750
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9770 17232 9826 17241
rect 9770 17167 9826 17176
rect 9784 17134 9812 17167
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9692 16794 9720 17070
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9770 16688 9826 16697
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9680 16652 9732 16658
rect 9770 16623 9826 16632
rect 9680 16594 9732 16600
rect 9600 16454 9628 16594
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9692 16289 9720 16594
rect 9784 16590 9812 16623
rect 9772 16584 9824 16590
rect 9772 16526 9824 16532
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9678 16280 9734 16289
rect 9678 16215 9680 16224
rect 9732 16215 9734 16224
rect 9680 16186 9732 16192
rect 9586 16144 9642 16153
rect 9586 16079 9588 16088
rect 9640 16079 9642 16088
rect 9588 16050 9640 16056
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9600 15638 9628 15846
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 9692 15502 9720 15982
rect 9784 15638 9812 16390
rect 9772 15632 9824 15638
rect 9772 15574 9824 15580
rect 9680 15496 9732 15502
rect 9876 15484 9904 17818
rect 9968 17320 9996 18788
rect 10048 18770 10100 18776
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10062 18524 10370 18533
rect 10062 18522 10068 18524
rect 10124 18522 10148 18524
rect 10204 18522 10228 18524
rect 10284 18522 10308 18524
rect 10364 18522 10370 18524
rect 10124 18470 10126 18522
rect 10306 18470 10308 18522
rect 10062 18468 10068 18470
rect 10124 18468 10148 18470
rect 10204 18468 10228 18470
rect 10284 18468 10308 18470
rect 10364 18468 10370 18470
rect 10062 18459 10370 18468
rect 10428 18426 10456 18770
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10416 18216 10468 18222
rect 10416 18158 10468 18164
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 10152 17746 10180 17818
rect 10140 17740 10192 17746
rect 10140 17682 10192 17688
rect 10428 17678 10456 18158
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 10062 17436 10370 17445
rect 10062 17434 10068 17436
rect 10124 17434 10148 17436
rect 10204 17434 10228 17436
rect 10284 17434 10308 17436
rect 10364 17434 10370 17436
rect 10124 17382 10126 17434
rect 10306 17382 10308 17434
rect 10062 17380 10068 17382
rect 10124 17380 10148 17382
rect 10204 17380 10228 17382
rect 10284 17380 10308 17382
rect 10364 17380 10370 17382
rect 10062 17371 10370 17380
rect 9968 17292 10364 17320
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 9954 17096 10010 17105
rect 9954 17031 10010 17040
rect 9968 16232 9996 17031
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 10060 16522 10088 16934
rect 10152 16726 10180 17138
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10336 17082 10364 17292
rect 10428 17270 10456 17614
rect 10520 17542 10548 18158
rect 10612 17882 10640 18770
rect 11072 18766 11100 19178
rect 11624 19174 11652 20946
rect 11716 19310 11744 21286
rect 11808 19514 11836 22714
rect 11900 22438 11928 24006
rect 11992 23866 12020 24142
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 11980 23588 12032 23594
rect 11980 23530 12032 23536
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22234 11928 22374
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11992 20398 12020 23530
rect 12084 22545 12112 24210
rect 12164 23792 12216 23798
rect 12164 23734 12216 23740
rect 12176 23662 12204 23734
rect 12164 23656 12216 23662
rect 12164 23598 12216 23604
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12070 22536 12126 22545
rect 12176 22506 12204 23462
rect 12070 22471 12126 22480
rect 12164 22500 12216 22506
rect 12084 21010 12112 22471
rect 12164 22442 12216 22448
rect 12176 22166 12204 22442
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 11980 20392 12032 20398
rect 11980 20334 12032 20340
rect 11888 19984 11940 19990
rect 11886 19952 11888 19961
rect 11940 19952 11942 19961
rect 11886 19887 11942 19896
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 19718 11928 19790
rect 11888 19712 11940 19718
rect 11888 19654 11940 19660
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11704 19304 11756 19310
rect 11704 19246 11756 19252
rect 11612 19168 11664 19174
rect 11612 19110 11664 19116
rect 11624 18834 11652 19110
rect 11612 18828 11664 18834
rect 11532 18788 11612 18816
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 11072 18290 11100 18702
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 10722 17980 11030 17989
rect 10722 17978 10728 17980
rect 10784 17978 10808 17980
rect 10864 17978 10888 17980
rect 10944 17978 10968 17980
rect 11024 17978 11030 17980
rect 10784 17926 10786 17978
rect 10966 17926 10968 17978
rect 10722 17924 10728 17926
rect 10784 17924 10808 17926
rect 10864 17924 10888 17926
rect 10944 17924 10968 17926
rect 11024 17924 11030 17926
rect 10722 17915 11030 17924
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10612 17338 10640 17546
rect 11072 17338 11100 18226
rect 11532 18086 11560 18788
rect 11612 18770 11664 18776
rect 11612 18624 11664 18630
rect 11612 18566 11664 18572
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17882 11560 18022
rect 11520 17876 11572 17882
rect 11520 17818 11572 17824
rect 11426 17776 11482 17785
rect 11336 17740 11388 17746
rect 11426 17711 11482 17720
rect 11336 17682 11388 17688
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 11072 17202 11100 17274
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10244 16794 10272 17070
rect 10336 17054 10548 17082
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10140 16720 10192 16726
rect 10336 16674 10364 16934
rect 10140 16662 10192 16668
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10152 16454 10180 16662
rect 10244 16646 10364 16674
rect 10244 16454 10272 16646
rect 10140 16448 10192 16454
rect 10140 16390 10192 16396
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10062 16348 10370 16357
rect 10062 16346 10068 16348
rect 10124 16346 10148 16348
rect 10204 16346 10228 16348
rect 10284 16346 10308 16348
rect 10364 16346 10370 16348
rect 10124 16294 10126 16346
rect 10306 16294 10308 16346
rect 10062 16292 10068 16294
rect 10124 16292 10148 16294
rect 10204 16292 10228 16294
rect 10284 16292 10308 16294
rect 10364 16292 10370 16294
rect 10062 16283 10370 16292
rect 9968 16204 10180 16232
rect 10152 15910 10180 16204
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 9680 15438 9732 15444
rect 9784 15456 9904 15484
rect 9956 15496 10008 15502
rect 9588 15360 9640 15366
rect 9784 15348 9812 15456
rect 9956 15438 10008 15444
rect 9588 15302 9640 15308
rect 9692 15320 9812 15348
rect 9864 15360 9916 15366
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9232 13382 9352 13410
rect 9404 13388 9456 13394
rect 8944 12776 8996 12782
rect 9128 12776 9180 12782
rect 8944 12718 8996 12724
rect 9126 12744 9128 12753
rect 9180 12744 9182 12753
rect 9126 12679 9182 12688
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12374 8984 12582
rect 9232 12434 9260 13382
rect 9404 13330 9456 13336
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9048 12406 9260 12434
rect 8944 12368 8996 12374
rect 8944 12310 8996 12316
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8864 11354 8892 11630
rect 8956 11354 8984 12174
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8944 11348 8996 11354
rect 8944 11290 8996 11296
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 10130 8892 10474
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9722 8892 10066
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8208 8900 8260 8906
rect 8312 8894 8432 8922
rect 8208 8842 8260 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8312 8430 8340 8774
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8024 8016 8076 8022
rect 8024 7958 8076 7964
rect 8036 7274 8064 7958
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8036 7002 8064 7210
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7852 6458 7880 6802
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7668 5358 7788 5386
rect 7668 5302 7696 5358
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7852 4826 7880 5102
rect 7840 4820 7892 4826
rect 7840 4762 7892 4768
rect 7932 4616 7984 4622
rect 8036 4570 8064 5646
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 7984 4564 8064 4570
rect 7932 4558 8064 4564
rect 7944 4542 8064 4558
rect 8036 4078 8064 4542
rect 8128 4282 8156 5170
rect 8300 5092 8352 5098
rect 8300 5034 8352 5040
rect 8312 4622 8340 5034
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8404 4282 8432 8894
rect 8496 8634 8524 9046
rect 8772 8838 8800 9046
rect 9048 8906 9076 12406
rect 9126 12336 9182 12345
rect 9126 12271 9182 12280
rect 9140 12238 9168 12271
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9140 10062 9168 10678
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9178 9168 9998
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9232 9058 9260 12038
rect 9140 9030 9260 9058
rect 9036 8900 9088 8906
rect 9036 8842 9088 8848
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 7954 8708 8502
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8574 7440 8630 7449
rect 8574 7375 8630 7384
rect 8588 7342 8616 7375
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8496 6866 8524 7278
rect 8588 7002 8616 7278
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6730 8524 6802
rect 8772 6746 8800 8774
rect 9048 8514 9076 8842
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8956 8486 9076 8514
rect 8864 8022 8892 8434
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8864 6934 8892 7346
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8852 6792 8904 6798
rect 8772 6740 8852 6746
rect 8772 6734 8904 6740
rect 8484 6724 8536 6730
rect 8772 6718 8892 6734
rect 8484 6666 8536 6672
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8772 5234 8800 6598
rect 8864 5710 8892 6718
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8576 4752 8628 4758
rect 8576 4694 8628 4700
rect 8116 4276 8168 4282
rect 8116 4218 8168 4224
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7852 3670 7880 4014
rect 7840 3664 7892 3670
rect 7840 3606 7892 3612
rect 7392 2746 7512 2774
rect 7576 2746 7788 2774
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7288 2508 7340 2514
rect 7288 2450 7340 2456
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 1834 7236 2246
rect 7196 1828 7248 1834
rect 7196 1770 7248 1776
rect 7300 1562 7328 2450
rect 7484 2310 7512 2746
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 2106 7512 2246
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 7484 1834 7512 2042
rect 7472 1828 7524 1834
rect 7472 1770 7524 1776
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 7378 1456 7434 1465
rect 7378 1391 7434 1400
rect 7392 1358 7420 1391
rect 7484 1358 7512 1770
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 7576 1426 7604 1498
rect 7668 1426 7696 2518
rect 7760 2446 7788 2746
rect 8220 2514 8248 4014
rect 8496 3602 8524 4218
rect 8588 3738 8616 4694
rect 8680 4690 8708 4966
rect 8864 4826 8892 5238
rect 8852 4820 8904 4826
rect 8852 4762 8904 4768
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 4146 8800 4422
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8772 3602 8800 4082
rect 8956 4078 8984 8486
rect 9036 8424 9088 8430
rect 9036 8366 9088 8372
rect 9048 8090 9076 8366
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 9140 7886 9168 9030
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7954 9260 8230
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9140 7478 9168 7822
rect 9128 7472 9180 7478
rect 9128 7414 9180 7420
rect 9232 7410 9260 7890
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9324 7290 9352 13262
rect 9416 12986 9444 13330
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 11694 9536 12786
rect 9600 11830 9628 15302
rect 9692 14958 9720 15320
rect 9864 15302 9916 15308
rect 9876 15094 9904 15302
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9692 12918 9720 14894
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9784 14414 9812 14758
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9784 14074 9812 14350
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9876 13954 9904 15030
rect 9968 15026 9996 15438
rect 10152 15416 10180 15846
rect 10244 15706 10272 15846
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10336 15502 10364 16118
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10232 15428 10284 15434
rect 10152 15388 10232 15416
rect 10232 15370 10284 15376
rect 10062 15260 10370 15269
rect 10062 15258 10068 15260
rect 10124 15258 10148 15260
rect 10204 15258 10228 15260
rect 10284 15258 10308 15260
rect 10364 15258 10370 15260
rect 10124 15206 10126 15258
rect 10306 15206 10308 15258
rect 10062 15204 10068 15206
rect 10124 15204 10148 15206
rect 10204 15204 10228 15206
rect 10284 15204 10308 15206
rect 10364 15204 10370 15206
rect 10062 15195 10370 15204
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10060 14618 10088 14894
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9784 13926 9904 13954
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9784 12764 9812 13926
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9692 12736 9812 12764
rect 9692 12442 9720 12736
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9416 10130 9444 10406
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9508 9586 9536 11630
rect 9600 11286 9628 11766
rect 9692 11694 9720 12106
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9588 11280 9640 11286
rect 9588 11222 9640 11228
rect 9784 11218 9812 12582
rect 9876 12434 9904 13806
rect 9968 13802 9996 14418
rect 10062 14172 10370 14181
rect 10062 14170 10068 14172
rect 10124 14170 10148 14172
rect 10204 14170 10228 14172
rect 10284 14170 10308 14172
rect 10364 14170 10370 14172
rect 10124 14118 10126 14170
rect 10306 14118 10308 14170
rect 10062 14116 10068 14118
rect 10124 14116 10148 14118
rect 10204 14116 10228 14118
rect 10284 14116 10308 14118
rect 10364 14116 10370 14118
rect 10062 14107 10370 14116
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 12986 9996 13738
rect 10062 13084 10370 13093
rect 10062 13082 10068 13084
rect 10124 13082 10148 13084
rect 10204 13082 10228 13084
rect 10284 13082 10308 13084
rect 10364 13082 10370 13084
rect 10124 13030 10126 13082
rect 10306 13030 10308 13082
rect 10062 13028 10068 13030
rect 10124 13028 10148 13030
rect 10204 13028 10228 13030
rect 10284 13028 10308 13030
rect 10364 13028 10370 13030
rect 10062 13019 10370 13028
rect 9956 12980 10008 12986
rect 10428 12968 10456 16934
rect 10520 14414 10548 17054
rect 10722 16892 11030 16901
rect 10722 16890 10728 16892
rect 10784 16890 10808 16892
rect 10864 16890 10888 16892
rect 10944 16890 10968 16892
rect 11024 16890 11030 16892
rect 10784 16838 10786 16890
rect 10966 16838 10968 16890
rect 10722 16836 10728 16838
rect 10784 16836 10808 16838
rect 10864 16836 10888 16838
rect 10944 16836 10968 16838
rect 11024 16836 11030 16838
rect 10722 16827 11030 16836
rect 10966 16688 11022 16697
rect 11072 16674 11100 17138
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11072 16646 11192 16674
rect 11256 16658 11284 17002
rect 11348 16794 11376 17682
rect 11440 17678 11468 17711
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 17270 11468 17614
rect 11428 17264 11480 17270
rect 11428 17206 11480 17212
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11440 16658 11468 17070
rect 10966 16623 11022 16632
rect 10980 15892 11008 16623
rect 10980 15864 11100 15892
rect 10722 15804 11030 15813
rect 10722 15802 10728 15804
rect 10784 15802 10808 15804
rect 10864 15802 10888 15804
rect 10944 15802 10968 15804
rect 11024 15802 11030 15804
rect 10784 15750 10786 15802
rect 10966 15750 10968 15802
rect 10722 15748 10728 15750
rect 10784 15748 10808 15750
rect 10864 15748 10888 15750
rect 10944 15748 10968 15750
rect 11024 15748 11030 15750
rect 10722 15739 11030 15748
rect 11072 15706 11100 15864
rect 11164 15706 11192 16646
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11624 16250 11652 18566
rect 11716 18222 11744 19246
rect 11808 18358 11836 19450
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11900 16658 11928 19654
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11992 18766 12020 19246
rect 12176 18970 12204 19858
rect 12268 19310 12296 26846
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12360 24750 12388 26794
rect 12636 25838 12664 29543
rect 12728 29238 12756 33050
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12714 29064 12770 29073
rect 12714 28999 12770 29008
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12636 25294 12664 25774
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12360 23186 12388 24686
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12360 23089 12388 23122
rect 12346 23080 12402 23089
rect 12346 23015 12402 23024
rect 12348 22976 12400 22982
rect 12348 22918 12400 22924
rect 12360 22710 12388 22918
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 12360 21486 12388 22510
rect 12452 22438 12480 24346
rect 12636 23798 12664 25230
rect 12624 23792 12676 23798
rect 12624 23734 12676 23740
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 22234 12480 22374
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12348 20392 12400 20398
rect 12348 20334 12400 20340
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12268 18834 12296 19110
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 11992 18222 12020 18702
rect 12084 18426 12112 18770
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12268 18290 12296 18770
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 12254 18184 12310 18193
rect 12254 18119 12310 18128
rect 12164 17060 12216 17066
rect 12164 17002 12216 17008
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12072 16652 12124 16658
rect 12072 16594 12124 16600
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11808 16046 11836 16390
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11348 15706 11376 15982
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10704 15094 10732 15574
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10980 14804 11008 15370
rect 11072 15026 11100 15642
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11348 14958 11376 15642
rect 11532 15570 11560 15846
rect 11716 15706 11744 15982
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11336 14952 11388 14958
rect 11150 14920 11206 14929
rect 11336 14894 11388 14900
rect 11426 14920 11482 14929
rect 11150 14855 11206 14864
rect 11426 14855 11482 14864
rect 11164 14822 11192 14855
rect 11152 14816 11204 14822
rect 10980 14776 11100 14804
rect 10722 14716 11030 14725
rect 10722 14714 10728 14716
rect 10784 14714 10808 14716
rect 10864 14714 10888 14716
rect 10944 14714 10968 14716
rect 11024 14714 11030 14716
rect 10784 14662 10786 14714
rect 10966 14662 10968 14714
rect 10722 14660 10728 14662
rect 10784 14660 10808 14662
rect 10864 14660 10888 14662
rect 10944 14660 10968 14662
rect 11024 14660 11030 14662
rect 10722 14651 11030 14660
rect 11072 14600 11100 14776
rect 11152 14758 11204 14764
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11072 14572 11192 14600
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10600 14272 10652 14278
rect 10600 14214 10652 14220
rect 9956 12922 10008 12928
rect 10336 12940 10456 12968
rect 9876 12406 9996 12434
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9876 11898 9904 12310
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9968 11778 9996 12406
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10060 12209 10088 12242
rect 10046 12200 10102 12209
rect 10046 12135 10102 12144
rect 10336 12102 10364 12940
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10428 12374 10456 12786
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10062 11996 10370 12005
rect 10062 11994 10068 11996
rect 10124 11994 10148 11996
rect 10204 11994 10228 11996
rect 10284 11994 10308 11996
rect 10364 11994 10370 11996
rect 10124 11942 10126 11994
rect 10306 11942 10308 11994
rect 10062 11940 10068 11942
rect 10124 11940 10148 11942
rect 10204 11940 10228 11942
rect 10284 11940 10308 11942
rect 10364 11940 10370 11942
rect 10062 11931 10370 11940
rect 9876 11750 9996 11778
rect 10428 11762 10456 12038
rect 10416 11756 10468 11762
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9600 10810 9628 11086
rect 9692 10810 9720 11086
rect 9588 10804 9640 10810
rect 9588 10746 9640 10752
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9876 10690 9904 11750
rect 10416 11698 10468 11704
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9784 10662 9904 10690
rect 9496 9580 9548 9586
rect 9496 9522 9548 9528
rect 9508 9042 9536 9522
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9600 8922 9628 10610
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10266 9720 10474
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9110 9720 9862
rect 9680 9104 9732 9110
rect 9680 9046 9732 9052
rect 9496 8900 9548 8906
rect 9600 8894 9720 8922
rect 9496 8842 9548 8848
rect 9508 8566 9536 8842
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9508 8430 9536 8502
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9416 7410 9444 8298
rect 9494 8120 9550 8129
rect 9494 8055 9496 8064
rect 9548 8055 9550 8064
rect 9496 8026 9548 8032
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9324 7262 9444 7290
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9128 5772 9180 5778
rect 9128 5714 9180 5720
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4282 9076 5034
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8956 3602 8984 4014
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8772 2582 8800 3538
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8956 2514 8984 3538
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7760 2106 7788 2382
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 8128 1562 8156 2382
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8220 1426 8248 2450
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8496 1834 8524 2314
rect 8484 1828 8536 1834
rect 8484 1770 8536 1776
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 7564 1420 7616 1426
rect 7564 1362 7616 1368
rect 7656 1420 7708 1426
rect 7656 1362 7708 1368
rect 8208 1420 8260 1426
rect 8208 1362 8260 1368
rect 7380 1352 7432 1358
rect 7380 1294 7432 1300
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7012 1216 7064 1222
rect 7012 1158 7064 1164
rect 6460 1012 6512 1018
rect 6460 954 6512 960
rect 6644 1012 6696 1018
rect 6644 954 6696 960
rect 7484 814 7512 1294
rect 8312 1290 8340 1498
rect 8496 1426 8524 1770
rect 8588 1562 8616 2450
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 1834 8708 2246
rect 8668 1828 8720 1834
rect 8668 1770 8720 1776
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 8956 1494 8984 2450
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 8484 1420 8536 1426
rect 8484 1362 8536 1368
rect 9048 1358 9076 3538
rect 9140 2378 9168 5714
rect 9324 5166 9352 7142
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9232 4758 9260 4966
rect 9416 4826 9444 7262
rect 9508 5794 9536 7686
rect 9600 6866 9628 8774
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9692 6746 9720 8894
rect 9784 7313 9812 10662
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9876 10198 9904 10474
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 9864 10056 9916 10062
rect 9862 10024 9864 10033
rect 9916 10024 9918 10033
rect 9862 9959 9918 9968
rect 9968 9625 9996 11630
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10060 11218 10088 11494
rect 10244 11354 10272 11630
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10336 11082 10364 11494
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10062 10908 10370 10917
rect 10062 10906 10068 10908
rect 10124 10906 10148 10908
rect 10204 10906 10228 10908
rect 10284 10906 10308 10908
rect 10364 10906 10370 10908
rect 10124 10854 10126 10906
rect 10306 10854 10308 10906
rect 10062 10852 10068 10854
rect 10124 10852 10148 10854
rect 10204 10852 10228 10854
rect 10284 10852 10308 10854
rect 10364 10852 10370 10854
rect 10062 10843 10370 10852
rect 10428 9994 10456 11154
rect 10520 10606 10548 14214
rect 10612 14074 10640 14214
rect 10600 14068 10652 14074
rect 10600 14010 10652 14016
rect 11072 13938 11100 14418
rect 11060 13932 11112 13938
rect 11060 13874 11112 13880
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13530 10640 13806
rect 11164 13734 11192 14572
rect 11256 14414 11284 14758
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 13870 11284 14350
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 11152 13728 11204 13734
rect 11152 13670 11204 13676
rect 10722 13628 11030 13637
rect 10722 13626 10728 13628
rect 10784 13626 10808 13628
rect 10864 13626 10888 13628
rect 10944 13626 10968 13628
rect 11024 13626 11030 13628
rect 10784 13574 10786 13626
rect 10966 13574 10968 13626
rect 10722 13572 10728 13574
rect 10784 13572 10808 13574
rect 10864 13572 10888 13574
rect 10944 13572 10968 13574
rect 11024 13572 11030 13574
rect 10722 13563 11030 13572
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 11164 13394 11192 13670
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 11152 13388 11204 13394
rect 11152 13330 11204 13336
rect 10612 12434 10640 13330
rect 10722 12540 11030 12549
rect 10722 12538 10728 12540
rect 10784 12538 10808 12540
rect 10864 12538 10888 12540
rect 10944 12538 10968 12540
rect 11024 12538 11030 12540
rect 10784 12486 10786 12538
rect 10966 12486 10968 12538
rect 10722 12484 10728 12486
rect 10784 12484 10808 12486
rect 10864 12484 10888 12486
rect 10944 12484 10968 12486
rect 11024 12484 11030 12486
rect 10722 12475 11030 12484
rect 11164 12481 11192 13330
rect 11244 12776 11296 12782
rect 11244 12718 11296 12724
rect 11150 12472 11206 12481
rect 10612 12406 10732 12434
rect 11150 12407 11206 12416
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10612 10606 10640 12038
rect 10704 11694 10732 12406
rect 10966 12336 11022 12345
rect 10784 12300 10836 12306
rect 10966 12271 10968 12280
rect 10784 12242 10836 12248
rect 11020 12271 11022 12280
rect 11152 12300 11204 12306
rect 10968 12242 11020 12248
rect 11152 12242 11204 12248
rect 10796 11762 10824 12242
rect 10968 12164 11020 12170
rect 10968 12106 11020 12112
rect 10980 11830 11008 12106
rect 11164 11898 11192 12242
rect 11256 12170 11284 12718
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 11164 11694 11192 11834
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 10722 11452 11030 11461
rect 10722 11450 10728 11452
rect 10784 11450 10808 11452
rect 10864 11450 10888 11452
rect 10944 11450 10968 11452
rect 11024 11450 11030 11452
rect 10784 11398 10786 11450
rect 10966 11398 10968 11450
rect 10722 11396 10728 11398
rect 10784 11396 10808 11398
rect 10864 11396 10888 11398
rect 10944 11396 10968 11398
rect 11024 11396 11030 11398
rect 10722 11387 11030 11396
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10508 10464 10560 10470
rect 10704 10452 10732 11290
rect 10968 11280 11020 11286
rect 10968 11222 11020 11228
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10888 10470 10916 11086
rect 10980 10810 11008 11222
rect 11256 11014 11284 11494
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 11256 10674 11284 10950
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10508 10406 10560 10412
rect 10612 10424 10732 10452
rect 10876 10464 10928 10470
rect 10520 10062 10548 10406
rect 10612 10248 10640 10424
rect 10876 10406 10928 10412
rect 10722 10364 11030 10373
rect 10722 10362 10728 10364
rect 10784 10362 10808 10364
rect 10864 10362 10888 10364
rect 10944 10362 10968 10364
rect 11024 10362 11030 10364
rect 10784 10310 10786 10362
rect 10966 10310 10968 10362
rect 10722 10308 10728 10310
rect 10784 10308 10808 10310
rect 10864 10308 10888 10310
rect 10944 10308 10968 10310
rect 11024 10308 11030 10310
rect 10722 10299 11030 10308
rect 10612 10220 10732 10248
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10598 10024 10654 10033
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10062 9820 10370 9829
rect 10062 9818 10068 9820
rect 10124 9818 10148 9820
rect 10204 9818 10228 9820
rect 10284 9818 10308 9820
rect 10364 9818 10370 9820
rect 10124 9766 10126 9818
rect 10306 9766 10308 9818
rect 10062 9764 10068 9766
rect 10124 9764 10148 9766
rect 10204 9764 10228 9766
rect 10284 9764 10308 9766
rect 10364 9764 10370 9766
rect 10062 9755 10370 9764
rect 9954 9616 10010 9625
rect 10520 9586 10548 9998
rect 10598 9959 10654 9968
rect 9954 9551 10010 9560
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 9956 9512 10008 9518
rect 9956 9454 10008 9460
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9968 9042 9996 9454
rect 10060 9110 10088 9454
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 9956 9036 10008 9042
rect 9876 8996 9956 9024
rect 9876 8566 9904 8996
rect 9956 8978 10008 8984
rect 10152 8922 10180 9522
rect 10612 9518 10640 9959
rect 10600 9512 10652 9518
rect 10704 9489 10732 10220
rect 11072 10130 11100 10542
rect 11152 10464 11204 10470
rect 11152 10406 11204 10412
rect 11164 10130 11192 10406
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 10796 9722 10824 10066
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 9454 10652 9460
rect 10690 9480 10746 9489
rect 10690 9415 10746 9424
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10416 9036 10468 9042
rect 10416 8978 10468 8984
rect 10060 8906 10180 8922
rect 10048 8900 10180 8906
rect 10100 8894 10180 8900
rect 10048 8842 10100 8848
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9864 8560 9916 8566
rect 9864 8502 9916 8508
rect 9864 7948 9916 7954
rect 9864 7890 9916 7896
rect 9876 7546 9904 7890
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9770 7304 9826 7313
rect 9770 7239 9826 7248
rect 9770 6896 9826 6905
rect 9826 6840 9904 6848
rect 9770 6831 9772 6840
rect 9824 6820 9904 6840
rect 9772 6802 9824 6808
rect 9600 6718 9720 6746
rect 9600 6118 9628 6718
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9692 6254 9720 6598
rect 9680 6248 9732 6254
rect 9678 6216 9680 6225
rect 9732 6216 9734 6225
rect 9678 6151 9734 6160
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9508 5766 9628 5794
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9220 4752 9272 4758
rect 9220 4694 9272 4700
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9232 3738 9260 4014
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9324 3602 9352 4694
rect 9508 4690 9536 5646
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9508 3602 9536 4626
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9600 3398 9628 5766
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 4758 9720 5646
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4010 9720 4422
rect 9784 4214 9812 6598
rect 9876 5710 9904 6820
rect 9968 6338 9996 8774
rect 10062 8732 10370 8741
rect 10062 8730 10068 8732
rect 10124 8730 10148 8732
rect 10204 8730 10228 8732
rect 10284 8730 10308 8732
rect 10364 8730 10370 8732
rect 10124 8678 10126 8730
rect 10306 8678 10308 8730
rect 10062 8676 10068 8678
rect 10124 8676 10148 8678
rect 10204 8676 10228 8678
rect 10284 8676 10308 8678
rect 10364 8676 10370 8678
rect 10062 8667 10370 8676
rect 10428 8498 10456 8978
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10520 8430 10548 8842
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10322 8256 10378 8265
rect 10322 8191 10378 8200
rect 10336 8022 10364 8191
rect 10324 8016 10376 8022
rect 10324 7958 10376 7964
rect 10336 7750 10364 7958
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10062 7644 10370 7653
rect 10062 7642 10068 7644
rect 10124 7642 10148 7644
rect 10204 7642 10228 7644
rect 10284 7642 10308 7644
rect 10364 7642 10370 7644
rect 10124 7590 10126 7642
rect 10306 7590 10308 7642
rect 10062 7588 10068 7590
rect 10124 7588 10148 7590
rect 10204 7588 10228 7590
rect 10284 7588 10308 7590
rect 10364 7588 10370 7590
rect 10062 7579 10370 7588
rect 10612 7410 10640 9318
rect 10722 9276 11030 9285
rect 10722 9274 10728 9276
rect 10784 9274 10808 9276
rect 10864 9274 10888 9276
rect 10944 9274 10968 9276
rect 11024 9274 11030 9276
rect 10784 9222 10786 9274
rect 10966 9222 10968 9274
rect 10722 9220 10728 9222
rect 10784 9220 10808 9222
rect 10864 9220 10888 9222
rect 10944 9220 10968 9222
rect 11024 9220 11030 9222
rect 10722 9211 11030 9220
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8634 10732 8910
rect 11072 8906 11100 10066
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10980 8430 11008 8842
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10722 8188 11030 8197
rect 10722 8186 10728 8188
rect 10784 8186 10808 8188
rect 10864 8186 10888 8188
rect 10944 8186 10968 8188
rect 11024 8186 11030 8188
rect 10784 8134 10786 8186
rect 10966 8134 10968 8186
rect 10722 8132 10728 8134
rect 10784 8132 10808 8134
rect 10864 8132 10888 8134
rect 10944 8132 10968 8134
rect 11024 8132 11030 8134
rect 10722 8123 11030 8132
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 10600 7404 10652 7410
rect 10600 7346 10652 7352
rect 10062 6556 10370 6565
rect 10062 6554 10068 6556
rect 10124 6554 10148 6556
rect 10204 6554 10228 6556
rect 10284 6554 10308 6556
rect 10364 6554 10370 6556
rect 10124 6502 10126 6554
rect 10306 6502 10308 6554
rect 10062 6500 10068 6502
rect 10124 6500 10148 6502
rect 10204 6500 10228 6502
rect 10284 6500 10308 6502
rect 10364 6500 10370 6502
rect 10062 6491 10370 6500
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 9968 6310 10088 6338
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5914 9996 6190
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10060 5794 10088 6310
rect 10152 5846 10180 6394
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10336 6202 10364 6258
rect 10244 6174 10364 6202
rect 10416 6180 10468 6186
rect 9968 5766 10088 5794
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9772 4208 9824 4214
rect 9772 4150 9824 4156
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9692 3584 9720 3946
rect 9784 3738 9812 4014
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9772 3596 9824 3602
rect 9692 3556 9772 3584
rect 9772 3538 9824 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9692 2938 9720 3402
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9600 2910 9720 2938
rect 9600 2774 9628 2910
rect 9784 2774 9812 3334
rect 9508 2746 9628 2774
rect 9692 2746 9812 2774
rect 9508 2650 9536 2746
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 9508 2122 9536 2586
rect 9692 2514 9720 2746
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9324 2094 9536 2122
rect 8392 1352 8444 1358
rect 9036 1352 9088 1358
rect 8444 1300 8800 1306
rect 8392 1294 8800 1300
rect 9036 1294 9088 1300
rect 8404 1290 8800 1294
rect 9324 1290 9352 2094
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9416 1426 9444 1974
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 9508 1562 9536 1838
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9404 1420 9456 1426
rect 9404 1362 9456 1368
rect 8300 1284 8352 1290
rect 8404 1284 8812 1290
rect 8404 1278 8760 1284
rect 8300 1226 8352 1232
rect 8760 1226 8812 1232
rect 9312 1284 9364 1290
rect 9312 1226 9364 1232
rect 9508 814 9536 1498
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9600 1018 9628 1362
rect 9692 1358 9720 1770
rect 9784 1426 9812 2518
rect 9772 1420 9824 1426
rect 9772 1362 9824 1368
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 9876 1222 9904 5510
rect 9968 1834 9996 5766
rect 10244 5574 10272 6174
rect 10416 6122 10468 6128
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5846 10364 6054
rect 10428 5914 10456 6122
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10062 5468 10370 5477
rect 10062 5466 10068 5468
rect 10124 5466 10148 5468
rect 10204 5466 10228 5468
rect 10284 5466 10308 5468
rect 10364 5466 10370 5468
rect 10124 5414 10126 5466
rect 10306 5414 10308 5466
rect 10062 5412 10068 5414
rect 10124 5412 10148 5414
rect 10204 5412 10228 5414
rect 10284 5412 10308 5414
rect 10364 5412 10370 5414
rect 10062 5403 10370 5412
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10062 4380 10370 4389
rect 10062 4378 10068 4380
rect 10124 4378 10148 4380
rect 10204 4378 10228 4380
rect 10284 4378 10308 4380
rect 10364 4378 10370 4380
rect 10124 4326 10126 4378
rect 10306 4326 10308 4378
rect 10062 4324 10068 4326
rect 10124 4324 10148 4326
rect 10204 4324 10228 4326
rect 10284 4324 10308 4326
rect 10364 4324 10370 4326
rect 10062 4315 10370 4324
rect 10428 3602 10456 4422
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10612 4128 10640 7346
rect 10722 7100 11030 7109
rect 10722 7098 10728 7100
rect 10784 7098 10808 7100
rect 10864 7098 10888 7100
rect 10944 7098 10968 7100
rect 11024 7098 11030 7100
rect 10784 7046 10786 7098
rect 10966 7046 10968 7098
rect 10722 7044 10728 7046
rect 10784 7044 10808 7046
rect 10864 7044 10888 7046
rect 10944 7044 10968 7046
rect 11024 7044 11030 7046
rect 10722 7035 11030 7044
rect 11072 6798 11100 7822
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11164 6458 11192 9551
rect 11348 8786 11376 12038
rect 11440 10198 11468 14855
rect 11624 14822 11652 15370
rect 11716 15026 11744 15642
rect 11794 15600 11850 15609
rect 11794 15535 11850 15544
rect 11808 15502 11836 15535
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11808 15094 11836 15438
rect 11900 15162 11928 16594
rect 11992 16046 12020 16594
rect 12084 16250 12112 16594
rect 12176 16590 12204 17002
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11900 14906 11928 15098
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11808 14878 11928 14906
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11716 14074 11744 14826
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11440 9042 11468 10134
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11256 8758 11376 8786
rect 11256 7954 11284 8758
rect 11440 8650 11468 8978
rect 11348 8634 11468 8650
rect 11336 8628 11468 8634
rect 11388 8622 11468 8628
rect 11336 8570 11388 8576
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11256 7002 11284 7890
rect 11244 6996 11296 7002
rect 11244 6938 11296 6944
rect 11348 6866 11376 8434
rect 11532 7886 11560 13806
rect 11612 13796 11664 13802
rect 11612 13738 11664 13744
rect 11624 13462 11652 13738
rect 11702 13696 11758 13705
rect 11702 13631 11758 13640
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11716 12850 11744 13631
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11624 12442 11652 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11716 12306 11744 12786
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 11694 11652 12106
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11624 9178 11652 11630
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 11716 9518 11744 11562
rect 11808 10606 11836 14878
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11900 13870 11928 14418
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11992 12918 12020 15982
rect 12084 15434 12112 16186
rect 12072 15428 12124 15434
rect 12072 15370 12124 15376
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12084 13870 12112 14418
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11900 11898 11928 12174
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12176 11218 12204 16526
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11992 10130 12020 10678
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11808 9722 11836 10066
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11624 8634 11652 9114
rect 11992 9042 12020 10066
rect 12268 10062 12296 18119
rect 12360 16522 12388 20334
rect 12440 18148 12492 18154
rect 12440 18090 12492 18096
rect 12348 16516 12400 16522
rect 12348 16458 12400 16464
rect 12360 15502 12388 16458
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12256 10056 12308 10062
rect 12256 9998 12308 10004
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12084 9042 12112 9862
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12176 9178 12204 9386
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11624 8362 11652 8570
rect 11612 8356 11664 8362
rect 11612 8298 11664 8304
rect 11624 7954 11652 8298
rect 11716 7954 11744 8774
rect 11992 8430 12020 8978
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11900 7546 11928 8298
rect 12176 7954 12204 8502
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11992 7342 12020 7686
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11336 6860 11388 6866
rect 11388 6820 11468 6848
rect 11336 6802 11388 6808
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10874 6216 10930 6225
rect 10874 6151 10876 6160
rect 10928 6151 10930 6160
rect 10876 6122 10928 6128
rect 10722 6012 11030 6021
rect 10722 6010 10728 6012
rect 10784 6010 10808 6012
rect 10864 6010 10888 6012
rect 10944 6010 10968 6012
rect 11024 6010 11030 6012
rect 10784 5958 10786 6010
rect 10966 5958 10968 6010
rect 10722 5956 10728 5958
rect 10784 5956 10808 5958
rect 10864 5956 10888 5958
rect 10944 5956 10968 5958
rect 11024 5956 11030 5958
rect 10722 5947 11030 5956
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11060 5160 11112 5166
rect 11060 5102 11112 5108
rect 10722 4924 11030 4933
rect 10722 4922 10728 4924
rect 10784 4922 10808 4924
rect 10864 4922 10888 4924
rect 10944 4922 10968 4924
rect 11024 4922 11030 4924
rect 10784 4870 10786 4922
rect 10966 4870 10968 4922
rect 10722 4868 10728 4870
rect 10784 4868 10808 4870
rect 10864 4868 10888 4870
rect 10944 4868 10968 4870
rect 11024 4868 11030 4870
rect 10722 4859 11030 4868
rect 11072 4486 11100 5102
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11256 4690 11284 4966
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10692 4140 10744 4146
rect 10612 4100 10692 4128
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10062 3292 10370 3301
rect 10062 3290 10068 3292
rect 10124 3290 10148 3292
rect 10204 3290 10228 3292
rect 10284 3290 10308 3292
rect 10364 3290 10370 3292
rect 10124 3238 10126 3290
rect 10306 3238 10308 3290
rect 10062 3236 10068 3238
rect 10124 3236 10148 3238
rect 10204 3236 10228 3238
rect 10284 3236 10308 3238
rect 10364 3236 10370 3238
rect 10062 3227 10370 3236
rect 10520 2650 10548 4082
rect 10612 3058 10640 4100
rect 10692 4082 10744 4088
rect 11164 4078 11192 4558
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 10722 3836 11030 3845
rect 10722 3834 10728 3836
rect 10784 3834 10808 3836
rect 10864 3834 10888 3836
rect 10944 3834 10968 3836
rect 11024 3834 11030 3836
rect 10784 3782 10786 3834
rect 10966 3782 10968 3834
rect 10722 3780 10728 3782
rect 10784 3780 10808 3782
rect 10864 3780 10888 3782
rect 10944 3780 10968 3782
rect 11024 3780 11030 3782
rect 10722 3771 11030 3780
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10508 2644 10560 2650
rect 10508 2586 10560 2592
rect 10046 2544 10102 2553
rect 10046 2479 10102 2488
rect 10416 2508 10468 2514
rect 10060 2446 10088 2479
rect 10416 2450 10468 2456
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10062 2204 10370 2213
rect 10062 2202 10068 2204
rect 10124 2202 10148 2204
rect 10204 2202 10228 2204
rect 10284 2202 10308 2204
rect 10364 2202 10370 2204
rect 10124 2150 10126 2202
rect 10306 2150 10308 2202
rect 10062 2148 10068 2150
rect 10124 2148 10148 2150
rect 10204 2148 10228 2150
rect 10284 2148 10308 2150
rect 10364 2148 10370 2150
rect 10062 2139 10370 2148
rect 10428 2106 10456 2450
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 10416 1896 10468 1902
rect 10336 1856 10416 1884
rect 9956 1828 10008 1834
rect 9956 1770 10008 1776
rect 10336 1442 10364 1856
rect 10416 1838 10468 1844
rect 10416 1760 10468 1766
rect 10416 1702 10468 1708
rect 10428 1562 10456 1702
rect 10416 1556 10468 1562
rect 10416 1498 10468 1504
rect 10336 1414 10456 1442
rect 10520 1426 10548 2382
rect 10612 1970 10640 2994
rect 10722 2748 11030 2757
rect 10722 2746 10728 2748
rect 10784 2746 10808 2748
rect 10864 2746 10888 2748
rect 10944 2746 10968 2748
rect 11024 2746 11030 2748
rect 10784 2694 10786 2746
rect 10966 2694 10968 2746
rect 10722 2692 10728 2694
rect 10784 2692 10808 2694
rect 10864 2692 10888 2694
rect 10944 2692 10968 2694
rect 11024 2692 11030 2694
rect 10722 2683 11030 2692
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 10704 1850 10732 2518
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 1902 10824 2246
rect 11256 1902 11284 3538
rect 11348 3398 11376 5170
rect 11440 5166 11468 6820
rect 12176 5370 12204 7890
rect 12268 7886 12296 9998
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 11612 5364 11664 5370
rect 11612 5306 11664 5312
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11440 4622 11468 5102
rect 11520 5092 11572 5098
rect 11520 5034 11572 5040
rect 11532 4758 11560 5034
rect 11624 4826 11652 5306
rect 12268 5234 12296 7822
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12256 5092 12308 5098
rect 12256 5034 12308 5040
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11532 3602 11560 4694
rect 11624 4690 11652 4762
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 3670 11744 4422
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11336 3392 11388 3398
rect 11336 3334 11388 3340
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11348 2774 11376 3334
rect 11532 2990 11560 3334
rect 12268 3194 12296 5034
rect 12360 4690 12388 14894
rect 12452 9110 12480 18090
rect 12544 17746 12572 23530
rect 12636 22094 12664 23734
rect 12728 23497 12756 28999
rect 12714 23488 12770 23497
rect 12714 23423 12770 23432
rect 12636 22066 12756 22094
rect 12728 21554 12756 22066
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12544 12170 12572 17682
rect 12532 12164 12584 12170
rect 12532 12106 12584 12112
rect 12440 9104 12492 9110
rect 12440 9046 12492 9052
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12360 4282 12388 4626
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12256 3188 12308 3194
rect 12256 3130 12308 3136
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 11348 2746 11468 2774
rect 10612 1822 10732 1850
rect 10784 1896 10836 1902
rect 10784 1838 10836 1844
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 10612 1562 10640 1822
rect 10722 1660 11030 1669
rect 10722 1658 10728 1660
rect 10784 1658 10808 1660
rect 10864 1658 10888 1660
rect 10944 1658 10968 1660
rect 11024 1658 11030 1660
rect 10784 1606 10786 1658
rect 10966 1606 10968 1658
rect 10722 1604 10728 1606
rect 10784 1604 10808 1606
rect 10864 1604 10888 1606
rect 10944 1604 10968 1606
rect 11024 1604 11030 1606
rect 10722 1595 11030 1604
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 9864 1216 9916 1222
rect 9864 1158 9916 1164
rect 10062 1116 10370 1125
rect 10062 1114 10068 1116
rect 10124 1114 10148 1116
rect 10204 1114 10228 1116
rect 10284 1114 10308 1116
rect 10364 1114 10370 1116
rect 10124 1062 10126 1114
rect 10306 1062 10308 1114
rect 10062 1060 10068 1062
rect 10124 1060 10148 1062
rect 10204 1060 10228 1062
rect 10284 1060 10308 1062
rect 10364 1060 10370 1062
rect 10062 1051 10370 1060
rect 9588 1012 9640 1018
rect 9588 954 9640 960
rect 10428 814 10456 1414
rect 10508 1420 10560 1426
rect 10508 1362 10560 1368
rect 11440 1290 11468 2746
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 6092 808 6144 814
rect 6092 750 6144 756
rect 6276 808 6328 814
rect 6276 750 6328 756
rect 7472 808 7524 814
rect 7472 750 7524 756
rect 9496 808 9548 814
rect 9496 750 9548 756
rect 10416 808 10468 814
rect 10416 750 10468 756
rect 4068 740 4120 746
rect 4068 682 4120 688
rect 3976 672 4028 678
rect 3976 614 4028 620
rect 4322 572 4630 581
rect 4322 570 4328 572
rect 4384 570 4408 572
rect 4464 570 4488 572
rect 4544 570 4568 572
rect 4624 570 4630 572
rect 4384 518 4386 570
rect 4566 518 4568 570
rect 4322 516 4328 518
rect 4384 516 4408 518
rect 4464 516 4488 518
rect 4544 516 4568 518
rect 4624 516 4630 518
rect 4322 507 4630 516
rect 10722 572 11030 581
rect 10722 570 10728 572
rect 10784 570 10808 572
rect 10864 570 10888 572
rect 10944 570 10968 572
rect 11024 570 11030 572
rect 10784 518 10786 570
rect 10966 518 10968 570
rect 10722 516 10728 518
rect 10784 516 10808 518
rect 10864 516 10888 518
rect 10944 516 10968 518
rect 11024 516 11030 518
rect 10722 507 11030 516
<< via2 >>
rect 2226 43560 2282 43616
rect 4986 43560 5042 43616
rect 6090 43560 6146 43616
rect 846 42608 902 42664
rect 938 41384 994 41440
rect 386 41112 442 41168
rect 570 40840 626 40896
rect 478 39888 534 39944
rect 386 38528 442 38584
rect 478 34856 534 34912
rect 846 40432 902 40488
rect 754 39344 810 39400
rect 938 39480 994 39536
rect 938 39244 940 39264
rect 940 39244 992 39264
rect 992 39244 994 39264
rect 938 39208 994 39244
rect 938 39072 994 39128
rect 1214 40568 1270 40624
rect 1122 39616 1178 39672
rect 1214 38936 1270 38992
rect 1398 40024 1454 40080
rect 1398 38836 1400 38856
rect 1400 38836 1452 38856
rect 1452 38836 1454 38856
rect 1030 37848 1086 37904
rect 1398 38800 1454 38836
rect 1122 37576 1178 37632
rect 1122 36896 1178 36952
rect 938 36760 994 36816
rect 1214 36760 1270 36816
rect 1122 36488 1178 36544
rect 846 36216 902 36272
rect 386 34584 442 34640
rect 386 31048 442 31104
rect 1030 35536 1086 35592
rect 938 34312 994 34368
rect 754 32000 810 32056
rect 662 31728 718 31784
rect 202 27648 258 27704
rect 846 31320 902 31376
rect 1214 31728 1270 31784
rect 754 28328 810 28384
rect 570 25064 626 25120
rect 478 23704 534 23760
rect 386 21936 442 21992
rect 478 15272 534 15328
rect 386 7112 442 7168
rect 754 24248 810 24304
rect 1030 28600 1086 28656
rect 1030 28328 1086 28384
rect 1122 28056 1178 28112
rect 1030 23976 1086 24032
rect 2042 41656 2098 41712
rect 2594 41112 2650 41168
rect 2502 40568 2558 40624
rect 2042 39616 2098 39672
rect 1950 39344 2006 39400
rect 1858 38800 1914 38856
rect 1490 37440 1546 37496
rect 1766 37712 1822 37768
rect 1490 37032 1546 37088
rect 1766 37032 1822 37088
rect 1674 35808 1730 35864
rect 1398 30912 1454 30968
rect 1766 34992 1822 35048
rect 2502 40024 2558 40080
rect 2318 39208 2374 39264
rect 2042 38120 2098 38176
rect 1950 37168 2006 37224
rect 4328 43002 4384 43004
rect 4408 43002 4464 43004
rect 4488 43002 4544 43004
rect 4568 43002 4624 43004
rect 4328 42950 4374 43002
rect 4374 42950 4384 43002
rect 4408 42950 4438 43002
rect 4438 42950 4450 43002
rect 4450 42950 4464 43002
rect 4488 42950 4502 43002
rect 4502 42950 4514 43002
rect 4514 42950 4544 43002
rect 4568 42950 4578 43002
rect 4578 42950 4624 43002
rect 4328 42948 4384 42950
rect 4408 42948 4464 42950
rect 4488 42948 4544 42950
rect 4568 42948 4624 42950
rect 4250 42608 4306 42664
rect 3668 42458 3724 42460
rect 3748 42458 3804 42460
rect 3828 42458 3884 42460
rect 3908 42458 3964 42460
rect 3668 42406 3714 42458
rect 3714 42406 3724 42458
rect 3748 42406 3778 42458
rect 3778 42406 3790 42458
rect 3790 42406 3804 42458
rect 3828 42406 3842 42458
rect 3842 42406 3854 42458
rect 3854 42406 3884 42458
rect 3908 42406 3918 42458
rect 3918 42406 3964 42458
rect 3668 42404 3724 42406
rect 3748 42404 3804 42406
rect 3828 42404 3884 42406
rect 3908 42404 3964 42406
rect 2962 40568 3018 40624
rect 3054 40180 3110 40216
rect 3054 40160 3056 40180
rect 3056 40160 3108 40180
rect 3108 40160 3110 40180
rect 2870 40024 2926 40080
rect 2778 39888 2834 39944
rect 3330 40704 3386 40760
rect 3054 39500 3110 39536
rect 3054 39480 3056 39500
rect 3056 39480 3108 39500
rect 3108 39480 3110 39500
rect 2134 37440 2190 37496
rect 2042 35672 2098 35728
rect 2502 36624 2558 36680
rect 2870 37712 2926 37768
rect 2594 35264 2650 35320
rect 1858 33632 1914 33688
rect 1950 33224 2006 33280
rect 1858 32136 1914 32192
rect 2502 34176 2558 34232
rect 2318 33396 2320 33416
rect 2320 33396 2372 33416
rect 2372 33396 2374 33416
rect 2318 33360 2374 33396
rect 2594 33088 2650 33144
rect 2686 32952 2742 33008
rect 1674 31456 1730 31512
rect 2042 31728 2098 31784
rect 1766 29844 1822 29880
rect 1766 29824 1768 29844
rect 1768 29824 1820 29844
rect 1820 29824 1822 29844
rect 1674 29008 1730 29064
rect 2502 31204 2558 31240
rect 2502 31184 2504 31204
rect 2504 31184 2556 31204
rect 2556 31184 2558 31204
rect 2870 33108 2926 33144
rect 2870 33088 2872 33108
rect 2872 33088 2924 33108
rect 2924 33088 2926 33108
rect 2870 32952 2926 33008
rect 2134 29552 2190 29608
rect 2042 29144 2098 29200
rect 1950 27784 2006 27840
rect 2410 30268 2412 30288
rect 2412 30268 2464 30288
rect 2464 30268 2466 30288
rect 2410 30232 2466 30268
rect 2870 30912 2926 30968
rect 2318 28872 2374 28928
rect 2134 26560 2190 26616
rect 2042 26288 2098 26344
rect 1766 24792 1822 24848
rect 1030 22652 1032 22672
rect 1032 22652 1084 22672
rect 1084 22652 1086 22672
rect 1030 22616 1086 22652
rect 754 19216 810 19272
rect 662 17584 718 17640
rect 938 17720 994 17776
rect 846 17176 902 17232
rect 938 16904 994 16960
rect 938 16496 994 16552
rect 846 12552 902 12608
rect 570 11192 626 11248
rect 938 12008 994 12064
rect 1306 23432 1362 23488
rect 1766 21800 1822 21856
rect 1122 20848 1178 20904
rect 1122 20576 1178 20632
rect 1674 21256 1730 21312
rect 1674 20576 1730 20632
rect 1306 16768 1362 16824
rect 1214 11736 1270 11792
rect 1030 11500 1032 11520
rect 1032 11500 1084 11520
rect 1084 11500 1086 11520
rect 1030 11464 1086 11500
rect 1674 19760 1730 19816
rect 1490 16496 1546 16552
rect 1398 12316 1400 12336
rect 1400 12316 1452 12336
rect 1452 12316 1454 12336
rect 1398 12280 1454 12316
rect 1674 15700 1730 15736
rect 1674 15680 1676 15700
rect 1676 15680 1728 15700
rect 1728 15680 1730 15700
rect 1674 15136 1730 15192
rect 2502 29552 2558 29608
rect 2778 30116 2834 30152
rect 2778 30096 2780 30116
rect 2780 30096 2832 30116
rect 2832 30096 2834 30116
rect 2778 29552 2834 29608
rect 2686 29144 2742 29200
rect 2594 27648 2650 27704
rect 3668 41370 3724 41372
rect 3748 41370 3804 41372
rect 3828 41370 3884 41372
rect 3908 41370 3964 41372
rect 3668 41318 3714 41370
rect 3714 41318 3724 41370
rect 3748 41318 3778 41370
rect 3778 41318 3790 41370
rect 3790 41318 3804 41370
rect 3828 41318 3842 41370
rect 3842 41318 3854 41370
rect 3854 41318 3884 41370
rect 3908 41318 3918 41370
rect 3918 41318 3964 41370
rect 3668 41316 3724 41318
rect 3748 41316 3804 41318
rect 3828 41316 3884 41318
rect 3908 41316 3964 41318
rect 4158 42472 4214 42528
rect 4328 41914 4384 41916
rect 4408 41914 4464 41916
rect 4488 41914 4544 41916
rect 4568 41914 4624 41916
rect 4328 41862 4374 41914
rect 4374 41862 4384 41914
rect 4408 41862 4438 41914
rect 4438 41862 4450 41914
rect 4450 41862 4464 41914
rect 4488 41862 4502 41914
rect 4502 41862 4514 41914
rect 4514 41862 4544 41914
rect 4568 41862 4578 41914
rect 4578 41862 4624 41914
rect 4328 41860 4384 41862
rect 4408 41860 4464 41862
rect 4488 41860 4544 41862
rect 4568 41860 4624 41862
rect 4328 40826 4384 40828
rect 4408 40826 4464 40828
rect 4488 40826 4544 40828
rect 4568 40826 4624 40828
rect 4328 40774 4374 40826
rect 4374 40774 4384 40826
rect 4408 40774 4438 40826
rect 4438 40774 4450 40826
rect 4450 40774 4464 40826
rect 4488 40774 4502 40826
rect 4502 40774 4514 40826
rect 4514 40774 4544 40826
rect 4568 40774 4578 40826
rect 4578 40774 4624 40826
rect 4328 40772 4384 40774
rect 4408 40772 4464 40774
rect 4488 40772 4544 40774
rect 4568 40772 4624 40774
rect 3514 40296 3570 40352
rect 3422 40024 3478 40080
rect 3668 40282 3724 40284
rect 3748 40282 3804 40284
rect 3828 40282 3884 40284
rect 3908 40282 3964 40284
rect 3668 40230 3714 40282
rect 3714 40230 3724 40282
rect 3748 40230 3778 40282
rect 3778 40230 3790 40282
rect 3790 40230 3804 40282
rect 3828 40230 3842 40282
rect 3842 40230 3854 40282
rect 3854 40230 3884 40282
rect 3908 40230 3918 40282
rect 3918 40230 3964 40282
rect 3668 40228 3724 40230
rect 3748 40228 3804 40230
rect 3828 40228 3884 40230
rect 3908 40228 3964 40230
rect 3668 39194 3724 39196
rect 3748 39194 3804 39196
rect 3828 39194 3884 39196
rect 3908 39194 3964 39196
rect 3668 39142 3714 39194
rect 3714 39142 3724 39194
rect 3748 39142 3778 39194
rect 3778 39142 3790 39194
rect 3790 39142 3804 39194
rect 3828 39142 3842 39194
rect 3842 39142 3854 39194
rect 3854 39142 3884 39194
rect 3908 39142 3918 39194
rect 3918 39142 3964 39194
rect 3668 39140 3724 39142
rect 3748 39140 3804 39142
rect 3828 39140 3884 39142
rect 3908 39140 3964 39142
rect 3882 38972 3884 38992
rect 3884 38972 3936 38992
rect 3936 38972 3938 38992
rect 3882 38936 3938 38972
rect 4328 39738 4384 39740
rect 4408 39738 4464 39740
rect 4488 39738 4544 39740
rect 4568 39738 4624 39740
rect 4328 39686 4374 39738
rect 4374 39686 4384 39738
rect 4408 39686 4438 39738
rect 4438 39686 4450 39738
rect 4450 39686 4464 39738
rect 4488 39686 4502 39738
rect 4502 39686 4514 39738
rect 4514 39686 4544 39738
rect 4568 39686 4578 39738
rect 4578 39686 4624 39738
rect 4328 39684 4384 39686
rect 4408 39684 4464 39686
rect 4488 39684 4544 39686
rect 4568 39684 4624 39686
rect 4986 42472 5042 42528
rect 5170 40704 5226 40760
rect 5262 40588 5318 40624
rect 5262 40568 5264 40588
rect 5264 40568 5316 40588
rect 5316 40568 5318 40588
rect 3422 37712 3478 37768
rect 3698 38256 3754 38312
rect 3668 38106 3724 38108
rect 3748 38106 3804 38108
rect 3828 38106 3884 38108
rect 3908 38106 3964 38108
rect 3668 38054 3714 38106
rect 3714 38054 3724 38106
rect 3748 38054 3778 38106
rect 3778 38054 3790 38106
rect 3790 38054 3804 38106
rect 3828 38054 3842 38106
rect 3842 38054 3854 38106
rect 3854 38054 3884 38106
rect 3908 38054 3918 38106
rect 3918 38054 3964 38106
rect 3668 38052 3724 38054
rect 3748 38052 3804 38054
rect 3828 38052 3884 38054
rect 3908 38052 3964 38054
rect 3974 37748 3976 37768
rect 3976 37748 4028 37768
rect 4028 37748 4030 37768
rect 3606 37576 3662 37632
rect 3974 37712 4030 37748
rect 3514 37304 3570 37360
rect 3790 37576 3846 37632
rect 3790 37440 3846 37496
rect 3054 35128 3110 35184
rect 3054 34604 3110 34640
rect 3054 34584 3056 34604
rect 3056 34584 3108 34604
rect 3108 34584 3110 34604
rect 3668 37018 3724 37020
rect 3748 37018 3804 37020
rect 3828 37018 3884 37020
rect 3908 37018 3964 37020
rect 3668 36966 3714 37018
rect 3714 36966 3724 37018
rect 3748 36966 3778 37018
rect 3778 36966 3790 37018
rect 3790 36966 3804 37018
rect 3828 36966 3842 37018
rect 3842 36966 3854 37018
rect 3854 36966 3884 37018
rect 3908 36966 3918 37018
rect 3918 36966 3964 37018
rect 3668 36964 3724 36966
rect 3748 36964 3804 36966
rect 3828 36964 3884 36966
rect 3908 36964 3964 36966
rect 3974 36216 4030 36272
rect 3668 35930 3724 35932
rect 3748 35930 3804 35932
rect 3828 35930 3884 35932
rect 3908 35930 3964 35932
rect 3668 35878 3714 35930
rect 3714 35878 3724 35930
rect 3748 35878 3778 35930
rect 3778 35878 3790 35930
rect 3790 35878 3804 35930
rect 3828 35878 3842 35930
rect 3842 35878 3854 35930
rect 3854 35878 3884 35930
rect 3908 35878 3918 35930
rect 3918 35878 3964 35930
rect 3668 35876 3724 35878
rect 3748 35876 3804 35878
rect 3828 35876 3884 35878
rect 3908 35876 3964 35878
rect 4328 38650 4384 38652
rect 4408 38650 4464 38652
rect 4488 38650 4544 38652
rect 4568 38650 4624 38652
rect 4328 38598 4374 38650
rect 4374 38598 4384 38650
rect 4408 38598 4438 38650
rect 4438 38598 4450 38650
rect 4450 38598 4464 38650
rect 4488 38598 4502 38650
rect 4502 38598 4514 38650
rect 4514 38598 4544 38650
rect 4568 38598 4578 38650
rect 4578 38598 4624 38650
rect 4328 38596 4384 38598
rect 4408 38596 4464 38598
rect 4488 38596 4544 38598
rect 4568 38596 4624 38598
rect 4986 39072 5042 39128
rect 4802 37576 4858 37632
rect 4328 37562 4384 37564
rect 4408 37562 4464 37564
rect 4488 37562 4544 37564
rect 4568 37562 4624 37564
rect 4328 37510 4374 37562
rect 4374 37510 4384 37562
rect 4408 37510 4438 37562
rect 4438 37510 4450 37562
rect 4450 37510 4464 37562
rect 4488 37510 4502 37562
rect 4502 37510 4514 37562
rect 4514 37510 4544 37562
rect 4568 37510 4578 37562
rect 4578 37510 4624 37562
rect 4328 37508 4384 37510
rect 4408 37508 4464 37510
rect 4488 37508 4544 37510
rect 4568 37508 4624 37510
rect 4434 37304 4490 37360
rect 4342 37168 4398 37224
rect 5630 40840 5686 40896
rect 5262 38548 5318 38584
rect 5262 38528 5264 38548
rect 5264 38528 5316 38548
rect 5316 38528 5318 38548
rect 5630 40024 5686 40080
rect 5446 37984 5502 38040
rect 5170 37440 5226 37496
rect 5170 37304 5226 37360
rect 4328 36474 4384 36476
rect 4408 36474 4464 36476
rect 4488 36474 4544 36476
rect 4568 36474 4624 36476
rect 4328 36422 4374 36474
rect 4374 36422 4384 36474
rect 4408 36422 4438 36474
rect 4438 36422 4450 36474
rect 4450 36422 4464 36474
rect 4488 36422 4502 36474
rect 4502 36422 4514 36474
rect 4514 36422 4544 36474
rect 4568 36422 4578 36474
rect 4578 36422 4624 36474
rect 4328 36420 4384 36422
rect 4408 36420 4464 36422
rect 4488 36420 4544 36422
rect 4568 36420 4624 36422
rect 3606 35264 3662 35320
rect 4066 35400 4122 35456
rect 4710 35808 4766 35864
rect 4328 35386 4384 35388
rect 4408 35386 4464 35388
rect 4488 35386 4544 35388
rect 4568 35386 4624 35388
rect 4328 35334 4374 35386
rect 4374 35334 4384 35386
rect 4408 35334 4438 35386
rect 4438 35334 4450 35386
rect 4450 35334 4464 35386
rect 4488 35334 4502 35386
rect 4502 35334 4514 35386
rect 4514 35334 4544 35386
rect 4568 35334 4578 35386
rect 4578 35334 4624 35386
rect 4328 35332 4384 35334
rect 4408 35332 4464 35334
rect 4488 35332 4544 35334
rect 4568 35332 4624 35334
rect 4158 34992 4214 35048
rect 3668 34842 3724 34844
rect 3748 34842 3804 34844
rect 3828 34842 3884 34844
rect 3908 34842 3964 34844
rect 3668 34790 3714 34842
rect 3714 34790 3724 34842
rect 3748 34790 3778 34842
rect 3778 34790 3790 34842
rect 3790 34790 3804 34842
rect 3828 34790 3842 34842
rect 3842 34790 3854 34842
rect 3854 34790 3884 34842
rect 3908 34790 3918 34842
rect 3918 34790 3964 34842
rect 3668 34788 3724 34790
rect 3748 34788 3804 34790
rect 3828 34788 3884 34790
rect 3908 34788 3964 34790
rect 3422 34448 3478 34504
rect 3330 33904 3386 33960
rect 4066 34720 4122 34776
rect 3790 34312 3846 34368
rect 3698 34176 3754 34232
rect 3974 33904 4030 33960
rect 3668 33754 3724 33756
rect 3748 33754 3804 33756
rect 3828 33754 3884 33756
rect 3908 33754 3964 33756
rect 3668 33702 3714 33754
rect 3714 33702 3724 33754
rect 3748 33702 3778 33754
rect 3778 33702 3790 33754
rect 3790 33702 3804 33754
rect 3828 33702 3842 33754
rect 3842 33702 3854 33754
rect 3854 33702 3884 33754
rect 3908 33702 3918 33754
rect 3918 33702 3964 33754
rect 3668 33700 3724 33702
rect 3748 33700 3804 33702
rect 3828 33700 3884 33702
rect 3908 33700 3964 33702
rect 3668 32666 3724 32668
rect 3748 32666 3804 32668
rect 3828 32666 3884 32668
rect 3908 32666 3964 32668
rect 3668 32614 3714 32666
rect 3714 32614 3724 32666
rect 3748 32614 3778 32666
rect 3778 32614 3790 32666
rect 3790 32614 3804 32666
rect 3828 32614 3842 32666
rect 3842 32614 3854 32666
rect 3854 32614 3884 32666
rect 3908 32614 3918 32666
rect 3918 32614 3964 32666
rect 3668 32612 3724 32614
rect 3748 32612 3804 32614
rect 3828 32612 3884 32614
rect 3908 32612 3964 32614
rect 4328 34298 4384 34300
rect 4408 34298 4464 34300
rect 4488 34298 4544 34300
rect 4568 34298 4624 34300
rect 4328 34246 4374 34298
rect 4374 34246 4384 34298
rect 4408 34246 4438 34298
rect 4438 34246 4450 34298
rect 4450 34246 4464 34298
rect 4488 34246 4502 34298
rect 4502 34246 4514 34298
rect 4514 34246 4544 34298
rect 4568 34246 4578 34298
rect 4578 34246 4624 34298
rect 4328 34244 4384 34246
rect 4408 34244 4464 34246
rect 4488 34244 4544 34246
rect 4568 34244 4624 34246
rect 4986 36760 5042 36816
rect 4986 35944 5042 36000
rect 4894 35400 4950 35456
rect 4894 34856 4950 34912
rect 4328 33210 4384 33212
rect 4408 33210 4464 33212
rect 4488 33210 4544 33212
rect 4568 33210 4624 33212
rect 4328 33158 4374 33210
rect 4374 33158 4384 33210
rect 4408 33158 4438 33210
rect 4438 33158 4450 33210
rect 4450 33158 4464 33210
rect 4488 33158 4502 33210
rect 4502 33158 4514 33210
rect 4514 33158 4544 33210
rect 4568 33158 4578 33210
rect 4578 33158 4624 33210
rect 4328 33156 4384 33158
rect 4408 33156 4464 33158
rect 4488 33156 4544 33158
rect 4568 33156 4624 33158
rect 4434 32680 4490 32736
rect 3146 31048 3202 31104
rect 4328 32122 4384 32124
rect 4408 32122 4464 32124
rect 4488 32122 4544 32124
rect 4568 32122 4624 32124
rect 4328 32070 4374 32122
rect 4374 32070 4384 32122
rect 4408 32070 4438 32122
rect 4438 32070 4450 32122
rect 4450 32070 4464 32122
rect 4488 32070 4502 32122
rect 4502 32070 4514 32122
rect 4514 32070 4544 32122
rect 4568 32070 4578 32122
rect 4578 32070 4624 32122
rect 4328 32068 4384 32070
rect 4408 32068 4464 32070
rect 4488 32068 4544 32070
rect 4568 32068 4624 32070
rect 3514 31592 3570 31648
rect 3330 31048 3386 31104
rect 3668 31578 3724 31580
rect 3748 31578 3804 31580
rect 3828 31578 3884 31580
rect 3908 31578 3964 31580
rect 3668 31526 3714 31578
rect 3714 31526 3724 31578
rect 3748 31526 3778 31578
rect 3778 31526 3790 31578
rect 3790 31526 3804 31578
rect 3828 31526 3842 31578
rect 3842 31526 3854 31578
rect 3854 31526 3884 31578
rect 3908 31526 3918 31578
rect 3918 31526 3964 31578
rect 3668 31524 3724 31526
rect 3748 31524 3804 31526
rect 3828 31524 3884 31526
rect 3908 31524 3964 31526
rect 4158 31592 4214 31648
rect 4250 31456 4306 31512
rect 4328 31034 4384 31036
rect 4408 31034 4464 31036
rect 4488 31034 4544 31036
rect 4568 31034 4624 31036
rect 4328 30982 4374 31034
rect 4374 30982 4384 31034
rect 4408 30982 4438 31034
rect 4438 30982 4450 31034
rect 4450 30982 4464 31034
rect 4488 30982 4502 31034
rect 4502 30982 4514 31034
rect 4514 30982 4544 31034
rect 4568 30982 4578 31034
rect 4578 30982 4624 31034
rect 4328 30980 4384 30982
rect 4408 30980 4464 30982
rect 4488 30980 4544 30982
rect 4568 30980 4624 30982
rect 4250 30776 4306 30832
rect 3668 30490 3724 30492
rect 3748 30490 3804 30492
rect 3828 30490 3884 30492
rect 3908 30490 3964 30492
rect 3668 30438 3714 30490
rect 3714 30438 3724 30490
rect 3748 30438 3778 30490
rect 3778 30438 3790 30490
rect 3790 30438 3804 30490
rect 3828 30438 3842 30490
rect 3842 30438 3854 30490
rect 3854 30438 3884 30490
rect 3908 30438 3918 30490
rect 3918 30438 3964 30490
rect 3668 30436 3724 30438
rect 3748 30436 3804 30438
rect 3828 30436 3884 30438
rect 3908 30436 3964 30438
rect 3238 30096 3294 30152
rect 2870 29300 2926 29336
rect 2870 29280 2872 29300
rect 2872 29280 2924 29300
rect 2924 29280 2926 29300
rect 3054 29416 3110 29472
rect 3146 29008 3202 29064
rect 2778 28192 2834 28248
rect 2410 26288 2466 26344
rect 2410 25880 2466 25936
rect 3054 27956 3056 27976
rect 3056 27956 3108 27976
rect 3108 27956 3110 27976
rect 3054 27920 3110 27956
rect 2870 25472 2926 25528
rect 2226 24656 2282 24712
rect 2042 24248 2098 24304
rect 2042 21392 2098 21448
rect 2042 20984 2098 21040
rect 1950 20848 2006 20904
rect 2042 19624 2098 19680
rect 1950 17584 2006 17640
rect 1950 16632 2006 16688
rect 2318 23432 2374 23488
rect 2318 23296 2374 23352
rect 2686 23160 2742 23216
rect 2318 22072 2374 22128
rect 2410 21936 2466 21992
rect 2778 22924 2780 22944
rect 2780 22924 2832 22944
rect 2832 22924 2834 22944
rect 2778 22888 2834 22924
rect 2962 23840 3018 23896
rect 3146 23568 3202 23624
rect 3054 23432 3110 23488
rect 2870 22616 2926 22672
rect 2594 21120 2650 21176
rect 2410 19932 2412 19952
rect 2412 19932 2464 19952
rect 2464 19932 2466 19952
rect 2410 19896 2466 19932
rect 2318 19760 2374 19816
rect 2318 19216 2374 19272
rect 2594 20576 2650 20632
rect 2686 19488 2742 19544
rect 2962 21548 3018 21584
rect 2962 21528 2964 21548
rect 2964 21528 3016 21548
rect 3016 21528 3018 21548
rect 3238 22108 3240 22128
rect 3240 22108 3292 22128
rect 3292 22108 3294 22128
rect 3238 22072 3294 22108
rect 3974 30116 4030 30152
rect 3974 30096 3976 30116
rect 3976 30096 4028 30116
rect 4028 30096 4030 30116
rect 3422 29416 3478 29472
rect 3422 29144 3478 29200
rect 3790 29844 3846 29880
rect 3790 29824 3792 29844
rect 3792 29824 3844 29844
rect 3844 29824 3846 29844
rect 3698 29552 3754 29608
rect 3974 29960 4030 30016
rect 4434 30232 4490 30288
rect 4342 30096 4398 30152
rect 4894 33632 4950 33688
rect 4894 32972 4950 33008
rect 4894 32952 4896 32972
rect 4896 32952 4948 32972
rect 4948 32952 4950 32972
rect 5078 32544 5134 32600
rect 4802 30232 4858 30288
rect 4618 30096 4674 30152
rect 4328 29946 4384 29948
rect 4408 29946 4464 29948
rect 4488 29946 4544 29948
rect 4568 29946 4624 29948
rect 4328 29894 4374 29946
rect 4374 29894 4384 29946
rect 4408 29894 4438 29946
rect 4438 29894 4450 29946
rect 4450 29894 4464 29946
rect 4488 29894 4502 29946
rect 4502 29894 4514 29946
rect 4514 29894 4544 29946
rect 4568 29894 4578 29946
rect 4578 29894 4624 29946
rect 4328 29892 4384 29894
rect 4408 29892 4464 29894
rect 4488 29892 4544 29894
rect 4568 29892 4624 29894
rect 3668 29402 3724 29404
rect 3748 29402 3804 29404
rect 3828 29402 3884 29404
rect 3908 29402 3964 29404
rect 3668 29350 3714 29402
rect 3714 29350 3724 29402
rect 3748 29350 3778 29402
rect 3778 29350 3790 29402
rect 3790 29350 3804 29402
rect 3828 29350 3842 29402
rect 3842 29350 3854 29402
rect 3854 29350 3884 29402
rect 3908 29350 3918 29402
rect 3918 29350 3964 29402
rect 3668 29348 3724 29350
rect 3748 29348 3804 29350
rect 3828 29348 3884 29350
rect 3908 29348 3964 29350
rect 3790 28620 3846 28656
rect 3790 28600 3792 28620
rect 3792 28600 3844 28620
rect 3844 28600 3846 28620
rect 3882 28464 3938 28520
rect 4066 28464 4122 28520
rect 3668 28314 3724 28316
rect 3748 28314 3804 28316
rect 3828 28314 3884 28316
rect 3908 28314 3964 28316
rect 3668 28262 3714 28314
rect 3714 28262 3724 28314
rect 3748 28262 3778 28314
rect 3778 28262 3790 28314
rect 3790 28262 3804 28314
rect 3828 28262 3842 28314
rect 3842 28262 3854 28314
rect 3854 28262 3884 28314
rect 3908 28262 3918 28314
rect 3918 28262 3964 28314
rect 3668 28260 3724 28262
rect 3748 28260 3804 28262
rect 3828 28260 3884 28262
rect 3908 28260 3964 28262
rect 4250 29416 4306 29472
rect 4802 29688 4858 29744
rect 5354 37748 5356 37768
rect 5356 37748 5408 37768
rect 5408 37748 5410 37768
rect 5354 37712 5410 37748
rect 5538 37576 5594 37632
rect 5354 36352 5410 36408
rect 5906 38392 5962 38448
rect 5630 36488 5686 36544
rect 5538 36080 5594 36136
rect 5354 35808 5410 35864
rect 5814 35808 5870 35864
rect 5446 35536 5502 35592
rect 5630 35556 5686 35592
rect 5630 35536 5632 35556
rect 5632 35536 5684 35556
rect 5684 35536 5686 35556
rect 5354 34856 5410 34912
rect 5538 34604 5594 34640
rect 5538 34584 5540 34604
rect 5540 34584 5592 34604
rect 5592 34584 5594 34604
rect 5446 34448 5502 34504
rect 5446 34176 5502 34232
rect 5446 33360 5502 33416
rect 5170 32000 5226 32056
rect 4986 31728 5042 31784
rect 5630 33632 5686 33688
rect 5354 32836 5410 32872
rect 5354 32816 5356 32836
rect 5356 32816 5408 32836
rect 5408 32816 5410 32836
rect 5078 30368 5134 30424
rect 4894 29416 4950 29472
rect 4526 29008 4582 29064
rect 4328 28858 4384 28860
rect 4408 28858 4464 28860
rect 4488 28858 4544 28860
rect 4568 28858 4624 28860
rect 4328 28806 4374 28858
rect 4374 28806 4384 28858
rect 4408 28806 4438 28858
rect 4438 28806 4450 28858
rect 4450 28806 4464 28858
rect 4488 28806 4502 28858
rect 4502 28806 4514 28858
rect 4514 28806 4544 28858
rect 4568 28806 4578 28858
rect 4578 28806 4624 28858
rect 4328 28804 4384 28806
rect 4408 28804 4464 28806
rect 4488 28804 4544 28806
rect 4568 28804 4624 28806
rect 4250 28464 4306 28520
rect 3668 27226 3724 27228
rect 3748 27226 3804 27228
rect 3828 27226 3884 27228
rect 3908 27226 3964 27228
rect 3668 27174 3714 27226
rect 3714 27174 3724 27226
rect 3748 27174 3778 27226
rect 3778 27174 3790 27226
rect 3790 27174 3804 27226
rect 3828 27174 3842 27226
rect 3842 27174 3854 27226
rect 3854 27174 3884 27226
rect 3908 27174 3918 27226
rect 3918 27174 3964 27226
rect 3668 27172 3724 27174
rect 3748 27172 3804 27174
rect 3828 27172 3884 27174
rect 3908 27172 3964 27174
rect 4066 26288 4122 26344
rect 3514 26152 3570 26208
rect 3668 26138 3724 26140
rect 3748 26138 3804 26140
rect 3828 26138 3884 26140
rect 3908 26138 3964 26140
rect 3668 26086 3714 26138
rect 3714 26086 3724 26138
rect 3748 26086 3778 26138
rect 3778 26086 3790 26138
rect 3790 26086 3804 26138
rect 3828 26086 3842 26138
rect 3842 26086 3854 26138
rect 3854 26086 3884 26138
rect 3908 26086 3918 26138
rect 3918 26086 3964 26138
rect 3668 26084 3724 26086
rect 3748 26084 3804 26086
rect 3828 26084 3884 26086
rect 3908 26084 3964 26086
rect 3974 25880 4030 25936
rect 4434 28212 4490 28248
rect 4434 28192 4436 28212
rect 4436 28192 4488 28212
rect 4488 28192 4490 28212
rect 4434 28056 4490 28112
rect 4802 28056 4858 28112
rect 4328 27770 4384 27772
rect 4408 27770 4464 27772
rect 4488 27770 4544 27772
rect 4568 27770 4624 27772
rect 4328 27718 4374 27770
rect 4374 27718 4384 27770
rect 4408 27718 4438 27770
rect 4438 27718 4450 27770
rect 4450 27718 4464 27770
rect 4488 27718 4502 27770
rect 4502 27718 4514 27770
rect 4514 27718 4544 27770
rect 4568 27718 4578 27770
rect 4578 27718 4624 27770
rect 4328 27716 4384 27718
rect 4408 27716 4464 27718
rect 4488 27716 4544 27718
rect 4568 27716 4624 27718
rect 4618 26832 4674 26888
rect 4328 26682 4384 26684
rect 4408 26682 4464 26684
rect 4488 26682 4544 26684
rect 4568 26682 4624 26684
rect 4328 26630 4374 26682
rect 4374 26630 4384 26682
rect 4408 26630 4438 26682
rect 4438 26630 4450 26682
rect 4450 26630 4464 26682
rect 4488 26630 4502 26682
rect 4502 26630 4514 26682
rect 4514 26630 4544 26682
rect 4568 26630 4578 26682
rect 4578 26630 4624 26682
rect 4328 26628 4384 26630
rect 4408 26628 4464 26630
rect 4488 26628 4544 26630
rect 4568 26628 4624 26630
rect 4526 25880 4582 25936
rect 3668 25050 3724 25052
rect 3748 25050 3804 25052
rect 3828 25050 3884 25052
rect 3908 25050 3964 25052
rect 3668 24998 3714 25050
rect 3714 24998 3724 25050
rect 3748 24998 3778 25050
rect 3778 24998 3790 25050
rect 3790 24998 3804 25050
rect 3828 24998 3842 25050
rect 3842 24998 3854 25050
rect 3854 24998 3884 25050
rect 3908 24998 3918 25050
rect 3918 24998 3964 25050
rect 3668 24996 3724 24998
rect 3748 24996 3804 24998
rect 3828 24996 3884 24998
rect 3908 24996 3964 24998
rect 3698 24268 3754 24304
rect 3698 24248 3700 24268
rect 3700 24248 3752 24268
rect 3752 24248 3754 24268
rect 4328 25594 4384 25596
rect 4408 25594 4464 25596
rect 4488 25594 4544 25596
rect 4568 25594 4624 25596
rect 4328 25542 4374 25594
rect 4374 25542 4384 25594
rect 4408 25542 4438 25594
rect 4438 25542 4450 25594
rect 4450 25542 4464 25594
rect 4488 25542 4502 25594
rect 4502 25542 4514 25594
rect 4514 25542 4544 25594
rect 4568 25542 4578 25594
rect 4578 25542 4624 25594
rect 4328 25540 4384 25542
rect 4408 25540 4464 25542
rect 4488 25540 4544 25542
rect 4568 25540 4624 25542
rect 4802 24928 4858 24984
rect 4328 24506 4384 24508
rect 4408 24506 4464 24508
rect 4488 24506 4544 24508
rect 4568 24506 4624 24508
rect 4328 24454 4374 24506
rect 4374 24454 4384 24506
rect 4408 24454 4438 24506
rect 4438 24454 4450 24506
rect 4450 24454 4464 24506
rect 4488 24454 4502 24506
rect 4502 24454 4514 24506
rect 4514 24454 4544 24506
rect 4568 24454 4578 24506
rect 4578 24454 4624 24506
rect 4328 24452 4384 24454
rect 4408 24452 4464 24454
rect 4488 24452 4544 24454
rect 4568 24452 4624 24454
rect 4066 24112 4122 24168
rect 3668 23962 3724 23964
rect 3748 23962 3804 23964
rect 3828 23962 3884 23964
rect 3908 23962 3964 23964
rect 3668 23910 3714 23962
rect 3714 23910 3724 23962
rect 3748 23910 3778 23962
rect 3778 23910 3790 23962
rect 3790 23910 3804 23962
rect 3828 23910 3842 23962
rect 3842 23910 3854 23962
rect 3854 23910 3884 23962
rect 3908 23910 3918 23962
rect 3918 23910 3964 23962
rect 3668 23908 3724 23910
rect 3748 23908 3804 23910
rect 3828 23908 3884 23910
rect 3908 23908 3964 23910
rect 4066 22888 4122 22944
rect 3668 22874 3724 22876
rect 3748 22874 3804 22876
rect 3828 22874 3884 22876
rect 3908 22874 3964 22876
rect 3668 22822 3714 22874
rect 3714 22822 3724 22874
rect 3748 22822 3778 22874
rect 3778 22822 3790 22874
rect 3790 22822 3804 22874
rect 3828 22822 3842 22874
rect 3842 22822 3854 22874
rect 3854 22822 3884 22874
rect 3908 22822 3918 22874
rect 3918 22822 3964 22874
rect 3668 22820 3724 22822
rect 3748 22820 3804 22822
rect 3828 22820 3884 22822
rect 3908 22820 3964 22822
rect 4328 23418 4384 23420
rect 4408 23418 4464 23420
rect 4488 23418 4544 23420
rect 4568 23418 4624 23420
rect 4328 23366 4374 23418
rect 4374 23366 4384 23418
rect 4408 23366 4438 23418
rect 4438 23366 4450 23418
rect 4450 23366 4464 23418
rect 4488 23366 4502 23418
rect 4502 23366 4514 23418
rect 4514 23366 4544 23418
rect 4568 23366 4578 23418
rect 4578 23366 4624 23418
rect 4328 23364 4384 23366
rect 4408 23364 4464 23366
rect 4488 23364 4544 23366
rect 4568 23364 4624 23366
rect 4434 23196 4436 23216
rect 4436 23196 4488 23216
rect 4488 23196 4490 23216
rect 4434 23160 4490 23196
rect 4618 23024 4674 23080
rect 3422 21936 3478 21992
rect 3146 21392 3202 21448
rect 4250 22636 4306 22672
rect 4250 22616 4252 22636
rect 4252 22616 4304 22636
rect 4304 22616 4306 22636
rect 4328 22330 4384 22332
rect 4408 22330 4464 22332
rect 4488 22330 4544 22332
rect 4568 22330 4624 22332
rect 4328 22278 4374 22330
rect 4374 22278 4384 22330
rect 4408 22278 4438 22330
rect 4438 22278 4450 22330
rect 4450 22278 4464 22330
rect 4488 22278 4502 22330
rect 4502 22278 4514 22330
rect 4514 22278 4544 22330
rect 4568 22278 4578 22330
rect 4578 22278 4624 22330
rect 4328 22276 4384 22278
rect 4408 22276 4464 22278
rect 4488 22276 4544 22278
rect 4568 22276 4624 22278
rect 4342 22072 4398 22128
rect 3668 21786 3724 21788
rect 3748 21786 3804 21788
rect 3828 21786 3884 21788
rect 3908 21786 3964 21788
rect 3668 21734 3714 21786
rect 3714 21734 3724 21786
rect 3748 21734 3778 21786
rect 3778 21734 3790 21786
rect 3790 21734 3804 21786
rect 3828 21734 3842 21786
rect 3842 21734 3854 21786
rect 3854 21734 3884 21786
rect 3908 21734 3918 21786
rect 3918 21734 3964 21786
rect 3668 21732 3724 21734
rect 3748 21732 3804 21734
rect 3828 21732 3884 21734
rect 3908 21732 3964 21734
rect 3606 21528 3662 21584
rect 3054 20984 3110 21040
rect 3330 20984 3386 21040
rect 3790 21428 3792 21448
rect 3792 21428 3844 21448
rect 3844 21428 3846 21448
rect 3790 21392 3846 21428
rect 3698 21256 3754 21312
rect 3698 20984 3754 21040
rect 3330 20848 3386 20904
rect 2870 19760 2926 19816
rect 3054 19780 3110 19816
rect 3054 19760 3056 19780
rect 3056 19760 3108 19780
rect 3108 19760 3110 19780
rect 3146 19624 3202 19680
rect 2134 17992 2190 18048
rect 2134 17060 2190 17096
rect 2134 17040 2136 17060
rect 2136 17040 2188 17060
rect 2188 17040 2190 17060
rect 2042 15544 2098 15600
rect 3054 19488 3110 19544
rect 3330 20304 3386 20360
rect 3668 20698 3724 20700
rect 3748 20698 3804 20700
rect 3828 20698 3884 20700
rect 3908 20698 3964 20700
rect 3668 20646 3714 20698
rect 3714 20646 3724 20698
rect 3748 20646 3778 20698
rect 3778 20646 3790 20698
rect 3790 20646 3804 20698
rect 3828 20646 3842 20698
rect 3842 20646 3854 20698
rect 3854 20646 3884 20698
rect 3908 20646 3918 20698
rect 3918 20646 3964 20698
rect 3668 20644 3724 20646
rect 3748 20644 3804 20646
rect 3828 20644 3884 20646
rect 3908 20644 3964 20646
rect 4066 20576 4122 20632
rect 3054 18828 3110 18864
rect 3054 18808 3056 18828
rect 3056 18808 3108 18828
rect 3108 18808 3110 18828
rect 2594 17040 2650 17096
rect 2686 16108 2742 16144
rect 2686 16088 2688 16108
rect 2688 16088 2740 16108
rect 2740 16088 2742 16108
rect 2962 16496 3018 16552
rect 2962 15272 3018 15328
rect 1950 11212 2006 11248
rect 1950 11192 1952 11212
rect 1952 11192 2004 11212
rect 2004 11192 2006 11212
rect 938 5480 994 5536
rect 2778 12724 2780 12744
rect 2780 12724 2832 12744
rect 2832 12724 2834 12744
rect 2778 12688 2834 12724
rect 2502 10920 2558 10976
rect 5078 29416 5134 29472
rect 5354 29960 5410 30016
rect 6366 41540 6422 41576
rect 6366 41520 6368 41540
rect 6368 41520 6420 41540
rect 6420 41520 6422 41540
rect 6366 40976 6422 41032
rect 6274 40704 6330 40760
rect 6274 39616 6330 39672
rect 5998 35284 6054 35320
rect 5998 35264 6000 35284
rect 6000 35264 6052 35284
rect 6052 35264 6054 35284
rect 6642 41656 6698 41712
rect 6550 41384 6606 41440
rect 6458 39072 6514 39128
rect 7746 43560 7802 43616
rect 8850 43560 8906 43616
rect 9402 43560 9458 43616
rect 6918 40296 6974 40352
rect 6734 40024 6790 40080
rect 6550 38936 6606 38992
rect 6182 35436 6184 35456
rect 6184 35436 6236 35456
rect 6236 35436 6238 35456
rect 6182 35400 6238 35436
rect 5998 34720 6054 34776
rect 6090 33768 6146 33824
rect 5814 32136 5870 32192
rect 5814 31728 5870 31784
rect 7470 42608 7526 42664
rect 7746 42472 7802 42528
rect 7378 41520 7434 41576
rect 7378 41248 7434 41304
rect 7654 41384 7710 41440
rect 7470 40468 7472 40488
rect 7472 40468 7524 40488
rect 7524 40468 7526 40488
rect 7470 40432 7526 40468
rect 8298 42644 8300 42664
rect 8300 42644 8352 42664
rect 8352 42644 8354 42664
rect 8298 42608 8354 42644
rect 7838 40024 7894 40080
rect 7286 39752 7342 39808
rect 7102 38800 7158 38856
rect 7378 39480 7434 39536
rect 7654 39480 7710 39536
rect 7470 38936 7526 38992
rect 7194 37984 7250 38040
rect 7010 37712 7066 37768
rect 6458 35808 6514 35864
rect 6366 34584 6422 34640
rect 6366 33632 6422 33688
rect 6366 33396 6368 33416
rect 6368 33396 6420 33416
rect 6420 33396 6422 33416
rect 6366 33360 6422 33396
rect 5814 31340 5870 31376
rect 5814 31320 5816 31340
rect 5816 31320 5868 31340
rect 5868 31320 5870 31340
rect 5814 31204 5870 31240
rect 5814 31184 5816 31204
rect 5816 31184 5868 31204
rect 5868 31184 5870 31204
rect 5814 30912 5870 30968
rect 5722 30640 5778 30696
rect 5722 30368 5778 30424
rect 5538 30232 5594 30288
rect 5906 30232 5962 30288
rect 5170 28736 5226 28792
rect 5814 29708 5870 29744
rect 5814 29688 5816 29708
rect 5816 29688 5868 29708
rect 5868 29688 5870 29708
rect 6366 32272 6422 32328
rect 6642 34312 6698 34368
rect 6642 33396 6644 33416
rect 6644 33396 6696 33416
rect 6696 33396 6698 33416
rect 6642 33360 6698 33396
rect 6918 36352 6974 36408
rect 7286 36660 7288 36680
rect 7288 36660 7340 36680
rect 7340 36660 7342 36680
rect 7286 36624 7342 36660
rect 7286 36352 7342 36408
rect 7470 36896 7526 36952
rect 8758 41248 8814 41304
rect 9126 41928 9182 41984
rect 8206 40296 8262 40352
rect 8114 39208 8170 39264
rect 8390 40568 8446 40624
rect 8206 38936 8262 38992
rect 7654 36216 7710 36272
rect 7838 36488 7894 36544
rect 8022 37576 8078 37632
rect 8114 36896 8170 36952
rect 8114 36760 8170 36816
rect 6826 33224 6882 33280
rect 6734 33088 6790 33144
rect 6734 32716 6736 32736
rect 6736 32716 6788 32736
rect 6788 32716 6790 32736
rect 6734 32680 6790 32716
rect 6734 32544 6790 32600
rect 6274 32136 6330 32192
rect 6366 31456 6422 31512
rect 6826 32308 6828 32328
rect 6828 32308 6880 32328
rect 6880 32308 6882 32328
rect 6826 32272 6882 32308
rect 6642 31728 6698 31784
rect 6826 31592 6882 31648
rect 6274 29960 6330 30016
rect 6366 29688 6422 29744
rect 4710 21664 4766 21720
rect 4710 21528 4766 21584
rect 4250 21428 4252 21448
rect 4252 21428 4304 21448
rect 4304 21428 4306 21448
rect 4250 21392 4306 21428
rect 4328 21242 4384 21244
rect 4408 21242 4464 21244
rect 4488 21242 4544 21244
rect 4568 21242 4624 21244
rect 4328 21190 4374 21242
rect 4374 21190 4384 21242
rect 4408 21190 4438 21242
rect 4438 21190 4450 21242
rect 4450 21190 4464 21242
rect 4488 21190 4502 21242
rect 4502 21190 4514 21242
rect 4514 21190 4544 21242
rect 4568 21190 4578 21242
rect 4578 21190 4624 21242
rect 4328 21188 4384 21190
rect 4408 21188 4464 21190
rect 4488 21188 4544 21190
rect 4568 21188 4624 21190
rect 4250 21004 4306 21040
rect 4250 20984 4252 21004
rect 4252 20984 4304 21004
rect 4304 20984 4306 21004
rect 4434 20984 4490 21040
rect 4710 20304 4766 20360
rect 4894 22888 4950 22944
rect 5078 22752 5134 22808
rect 5630 25744 5686 25800
rect 5262 25064 5318 25120
rect 4986 22208 5042 22264
rect 4986 21936 5042 21992
rect 4894 21836 4896 21856
rect 4896 21836 4948 21856
rect 4948 21836 4950 21856
rect 4894 21800 4950 21836
rect 4158 20052 4214 20088
rect 4158 20032 4160 20052
rect 4160 20032 4212 20052
rect 4212 20032 4214 20052
rect 3668 19610 3724 19612
rect 3748 19610 3804 19612
rect 3828 19610 3884 19612
rect 3908 19610 3964 19612
rect 3668 19558 3714 19610
rect 3714 19558 3724 19610
rect 3748 19558 3778 19610
rect 3778 19558 3790 19610
rect 3790 19558 3804 19610
rect 3828 19558 3842 19610
rect 3842 19558 3854 19610
rect 3854 19558 3884 19610
rect 3908 19558 3918 19610
rect 3918 19558 3964 19610
rect 3668 19556 3724 19558
rect 3748 19556 3804 19558
rect 3828 19556 3884 19558
rect 3908 19556 3964 19558
rect 3422 19080 3478 19136
rect 4328 20154 4384 20156
rect 4408 20154 4464 20156
rect 4488 20154 4544 20156
rect 4568 20154 4624 20156
rect 4328 20102 4374 20154
rect 4374 20102 4384 20154
rect 4408 20102 4438 20154
rect 4438 20102 4450 20154
rect 4450 20102 4464 20154
rect 4488 20102 4502 20154
rect 4502 20102 4514 20154
rect 4514 20102 4544 20154
rect 4568 20102 4578 20154
rect 4578 20102 4624 20154
rect 4328 20100 4384 20102
rect 4408 20100 4464 20102
rect 4488 20100 4544 20102
rect 4568 20100 4624 20102
rect 4342 19488 4398 19544
rect 4526 19624 4582 19680
rect 3698 19216 3754 19272
rect 3606 18944 3662 19000
rect 3790 18944 3846 19000
rect 4894 19624 4950 19680
rect 4328 19066 4384 19068
rect 4408 19066 4464 19068
rect 4488 19066 4544 19068
rect 4568 19066 4624 19068
rect 4328 19014 4374 19066
rect 4374 19014 4384 19066
rect 4408 19014 4438 19066
rect 4438 19014 4450 19066
rect 4450 19014 4464 19066
rect 4488 19014 4502 19066
rect 4502 19014 4514 19066
rect 4514 19014 4544 19066
rect 4568 19014 4578 19066
rect 4578 19014 4624 19066
rect 4328 19012 4384 19014
rect 4408 19012 4464 19014
rect 4488 19012 4544 19014
rect 4568 19012 4624 19014
rect 3514 18672 3570 18728
rect 4066 18808 4122 18864
rect 3668 18522 3724 18524
rect 3748 18522 3804 18524
rect 3828 18522 3884 18524
rect 3908 18522 3964 18524
rect 3668 18470 3714 18522
rect 3714 18470 3724 18522
rect 3748 18470 3778 18522
rect 3778 18470 3790 18522
rect 3790 18470 3804 18522
rect 3828 18470 3842 18522
rect 3842 18470 3854 18522
rect 3854 18470 3884 18522
rect 3908 18470 3918 18522
rect 3918 18470 3964 18522
rect 3668 18468 3724 18470
rect 3748 18468 3804 18470
rect 3828 18468 3884 18470
rect 3908 18468 3964 18470
rect 3422 17992 3478 18048
rect 4066 18128 4122 18184
rect 3422 17720 3478 17776
rect 3882 17720 3938 17776
rect 3668 17434 3724 17436
rect 3748 17434 3804 17436
rect 3828 17434 3884 17436
rect 3908 17434 3964 17436
rect 3668 17382 3714 17434
rect 3714 17382 3724 17434
rect 3748 17382 3778 17434
rect 3778 17382 3790 17434
rect 3790 17382 3804 17434
rect 3828 17382 3842 17434
rect 3842 17382 3854 17434
rect 3854 17382 3884 17434
rect 3908 17382 3918 17434
rect 3918 17382 3964 17434
rect 3668 17380 3724 17382
rect 3748 17380 3804 17382
rect 3828 17380 3884 17382
rect 3908 17380 3964 17382
rect 3668 16346 3724 16348
rect 3748 16346 3804 16348
rect 3828 16346 3884 16348
rect 3908 16346 3964 16348
rect 3668 16294 3714 16346
rect 3714 16294 3724 16346
rect 3748 16294 3778 16346
rect 3778 16294 3790 16346
rect 3790 16294 3804 16346
rect 3828 16294 3842 16346
rect 3842 16294 3854 16346
rect 3854 16294 3884 16346
rect 3908 16294 3918 16346
rect 3918 16294 3964 16346
rect 3668 16292 3724 16294
rect 3748 16292 3804 16294
rect 3828 16292 3884 16294
rect 3908 16292 3964 16294
rect 3514 15816 3570 15872
rect 4342 18128 4398 18184
rect 4710 18672 4766 18728
rect 4328 17978 4384 17980
rect 4408 17978 4464 17980
rect 4488 17978 4544 17980
rect 4568 17978 4624 17980
rect 4328 17926 4374 17978
rect 4374 17926 4384 17978
rect 4408 17926 4438 17978
rect 4438 17926 4450 17978
rect 4450 17926 4464 17978
rect 4488 17926 4502 17978
rect 4502 17926 4514 17978
rect 4514 17926 4544 17978
rect 4568 17926 4578 17978
rect 4578 17926 4624 17978
rect 4328 17924 4384 17926
rect 4408 17924 4464 17926
rect 4488 17924 4544 17926
rect 4568 17924 4624 17926
rect 1122 5208 1178 5264
rect 386 4664 442 4720
rect 3668 15258 3724 15260
rect 3748 15258 3804 15260
rect 3828 15258 3884 15260
rect 3908 15258 3964 15260
rect 3668 15206 3714 15258
rect 3714 15206 3724 15258
rect 3748 15206 3778 15258
rect 3778 15206 3790 15258
rect 3790 15206 3804 15258
rect 3828 15206 3842 15258
rect 3842 15206 3854 15258
rect 3854 15206 3884 15258
rect 3908 15206 3918 15258
rect 3918 15206 3964 15258
rect 3668 15204 3724 15206
rect 3748 15204 3804 15206
rect 3828 15204 3884 15206
rect 3908 15204 3964 15206
rect 3974 15000 4030 15056
rect 3698 14864 3754 14920
rect 3668 14170 3724 14172
rect 3748 14170 3804 14172
rect 3828 14170 3884 14172
rect 3908 14170 3964 14172
rect 3668 14118 3714 14170
rect 3714 14118 3724 14170
rect 3748 14118 3778 14170
rect 3778 14118 3790 14170
rect 3790 14118 3804 14170
rect 3828 14118 3842 14170
rect 3842 14118 3854 14170
rect 3854 14118 3884 14170
rect 3908 14118 3918 14170
rect 3918 14118 3964 14170
rect 3668 14116 3724 14118
rect 3748 14116 3804 14118
rect 3828 14116 3884 14118
rect 3908 14116 3964 14118
rect 4802 17740 4858 17776
rect 4802 17720 4804 17740
rect 4804 17720 4856 17740
rect 4856 17720 4858 17740
rect 4526 17040 4582 17096
rect 4328 16890 4384 16892
rect 4408 16890 4464 16892
rect 4488 16890 4544 16892
rect 4568 16890 4624 16892
rect 4328 16838 4374 16890
rect 4374 16838 4384 16890
rect 4408 16838 4438 16890
rect 4438 16838 4450 16890
rect 4450 16838 4464 16890
rect 4488 16838 4502 16890
rect 4502 16838 4514 16890
rect 4514 16838 4544 16890
rect 4568 16838 4578 16890
rect 4578 16838 4624 16890
rect 4328 16836 4384 16838
rect 4408 16836 4464 16838
rect 4488 16836 4544 16838
rect 4568 16836 4624 16838
rect 4434 16532 4436 16552
rect 4436 16532 4488 16552
rect 4488 16532 4490 16552
rect 4434 16496 4490 16532
rect 4328 15802 4384 15804
rect 4408 15802 4464 15804
rect 4488 15802 4544 15804
rect 4568 15802 4624 15804
rect 4328 15750 4374 15802
rect 4374 15750 4384 15802
rect 4408 15750 4438 15802
rect 4438 15750 4450 15802
rect 4450 15750 4464 15802
rect 4488 15750 4502 15802
rect 4502 15750 4514 15802
rect 4514 15750 4544 15802
rect 4568 15750 4578 15802
rect 4578 15750 4624 15802
rect 4328 15748 4384 15750
rect 4408 15748 4464 15750
rect 4488 15748 4544 15750
rect 4568 15748 4624 15750
rect 4158 15000 4214 15056
rect 4328 14714 4384 14716
rect 4408 14714 4464 14716
rect 4488 14714 4544 14716
rect 4568 14714 4624 14716
rect 4328 14662 4374 14714
rect 4374 14662 4384 14714
rect 4408 14662 4438 14714
rect 4438 14662 4450 14714
rect 4450 14662 4464 14714
rect 4488 14662 4502 14714
rect 4502 14662 4514 14714
rect 4514 14662 4544 14714
rect 4568 14662 4578 14714
rect 4578 14662 4624 14714
rect 4328 14660 4384 14662
rect 4408 14660 4464 14662
rect 4488 14660 4544 14662
rect 4568 14660 4624 14662
rect 4158 14456 4214 14512
rect 4328 13626 4384 13628
rect 4408 13626 4464 13628
rect 4488 13626 4544 13628
rect 4568 13626 4624 13628
rect 4328 13574 4374 13626
rect 4374 13574 4384 13626
rect 4408 13574 4438 13626
rect 4438 13574 4450 13626
rect 4450 13574 4464 13626
rect 4488 13574 4502 13626
rect 4502 13574 4514 13626
rect 4514 13574 4544 13626
rect 4568 13574 4578 13626
rect 4578 13574 4624 13626
rect 4328 13572 4384 13574
rect 4408 13572 4464 13574
rect 4488 13572 4544 13574
rect 4568 13572 4624 13574
rect 3668 13082 3724 13084
rect 3748 13082 3804 13084
rect 3828 13082 3884 13084
rect 3908 13082 3964 13084
rect 3668 13030 3714 13082
rect 3714 13030 3724 13082
rect 3748 13030 3778 13082
rect 3778 13030 3790 13082
rect 3790 13030 3804 13082
rect 3828 13030 3842 13082
rect 3842 13030 3854 13082
rect 3854 13030 3884 13082
rect 3908 13030 3918 13082
rect 3918 13030 3964 13082
rect 3668 13028 3724 13030
rect 3748 13028 3804 13030
rect 3828 13028 3884 13030
rect 3908 13028 3964 13030
rect 3668 11994 3724 11996
rect 3748 11994 3804 11996
rect 3828 11994 3884 11996
rect 3908 11994 3964 11996
rect 3668 11942 3714 11994
rect 3714 11942 3724 11994
rect 3748 11942 3778 11994
rect 3778 11942 3790 11994
rect 3790 11942 3804 11994
rect 3828 11942 3842 11994
rect 3842 11942 3854 11994
rect 3854 11942 3884 11994
rect 3908 11942 3918 11994
rect 3918 11942 3964 11994
rect 3668 11940 3724 11942
rect 3748 11940 3804 11942
rect 3828 11940 3884 11942
rect 3908 11940 3964 11942
rect 3668 10906 3724 10908
rect 3748 10906 3804 10908
rect 3828 10906 3884 10908
rect 3908 10906 3964 10908
rect 3668 10854 3714 10906
rect 3714 10854 3724 10906
rect 3748 10854 3778 10906
rect 3778 10854 3790 10906
rect 3790 10854 3804 10906
rect 3828 10854 3842 10906
rect 3842 10854 3854 10906
rect 3854 10854 3884 10906
rect 3908 10854 3918 10906
rect 3918 10854 3964 10906
rect 3668 10852 3724 10854
rect 3748 10852 3804 10854
rect 3828 10852 3884 10854
rect 3908 10852 3964 10854
rect 3422 8880 3478 8936
rect 2870 5772 2926 5808
rect 2870 5752 2872 5772
rect 2872 5752 2924 5772
rect 2924 5752 2926 5772
rect 4158 12960 4214 13016
rect 4328 12538 4384 12540
rect 4408 12538 4464 12540
rect 4488 12538 4544 12540
rect 4568 12538 4624 12540
rect 4328 12486 4374 12538
rect 4374 12486 4384 12538
rect 4408 12486 4438 12538
rect 4438 12486 4450 12538
rect 4450 12486 4464 12538
rect 4488 12486 4502 12538
rect 4502 12486 4514 12538
rect 4514 12486 4544 12538
rect 4568 12486 4578 12538
rect 4578 12486 4624 12538
rect 4328 12484 4384 12486
rect 4408 12484 4464 12486
rect 4488 12484 4544 12486
rect 4568 12484 4624 12486
rect 5354 24384 5410 24440
rect 5814 27376 5870 27432
rect 5814 24792 5870 24848
rect 5814 24692 5816 24712
rect 5816 24692 5868 24712
rect 5868 24692 5870 24712
rect 5814 24656 5870 24692
rect 5722 24520 5778 24576
rect 5354 22208 5410 22264
rect 5078 20576 5134 20632
rect 5078 20440 5134 20496
rect 5354 21664 5410 21720
rect 4986 18128 5042 18184
rect 4986 17076 4988 17096
rect 4988 17076 5040 17096
rect 5040 17076 5042 17096
rect 4986 17040 5042 17076
rect 5354 20984 5410 21040
rect 5354 20884 5356 20904
rect 5356 20884 5408 20904
rect 5408 20884 5410 20904
rect 5354 20848 5410 20884
rect 5262 19352 5318 19408
rect 5722 21972 5724 21992
rect 5724 21972 5776 21992
rect 5776 21972 5778 21992
rect 5722 21936 5778 21972
rect 5630 21800 5686 21856
rect 5538 21256 5594 21312
rect 5446 19624 5502 19680
rect 5814 21800 5870 21856
rect 5630 20168 5686 20224
rect 5814 20440 5870 20496
rect 5446 18944 5502 19000
rect 5078 16360 5134 16416
rect 5078 14764 5080 14784
rect 5080 14764 5132 14784
rect 5132 14764 5134 14784
rect 5078 14728 5134 14764
rect 4158 12280 4214 12336
rect 4434 12300 4490 12336
rect 4434 12280 4436 12300
rect 4436 12280 4488 12300
rect 4488 12280 4490 12300
rect 3606 9968 3662 10024
rect 3668 9818 3724 9820
rect 3748 9818 3804 9820
rect 3828 9818 3884 9820
rect 3908 9818 3964 9820
rect 3668 9766 3714 9818
rect 3714 9766 3724 9818
rect 3748 9766 3778 9818
rect 3778 9766 3790 9818
rect 3790 9766 3804 9818
rect 3828 9766 3842 9818
rect 3842 9766 3854 9818
rect 3854 9766 3884 9818
rect 3908 9766 3918 9818
rect 3918 9766 3964 9818
rect 3668 9764 3724 9766
rect 3748 9764 3804 9766
rect 3828 9764 3884 9766
rect 3908 9764 3964 9766
rect 3606 8880 3662 8936
rect 3668 8730 3724 8732
rect 3748 8730 3804 8732
rect 3828 8730 3884 8732
rect 3908 8730 3964 8732
rect 3668 8678 3714 8730
rect 3714 8678 3724 8730
rect 3748 8678 3778 8730
rect 3778 8678 3790 8730
rect 3790 8678 3804 8730
rect 3828 8678 3842 8730
rect 3842 8678 3854 8730
rect 3854 8678 3884 8730
rect 3908 8678 3918 8730
rect 3918 8678 3964 8730
rect 3668 8676 3724 8678
rect 3748 8676 3804 8678
rect 3828 8676 3884 8678
rect 3908 8676 3964 8678
rect 3668 7642 3724 7644
rect 3748 7642 3804 7644
rect 3828 7642 3884 7644
rect 3908 7642 3964 7644
rect 3668 7590 3714 7642
rect 3714 7590 3724 7642
rect 3748 7590 3778 7642
rect 3778 7590 3790 7642
rect 3790 7590 3804 7642
rect 3828 7590 3842 7642
rect 3842 7590 3854 7642
rect 3854 7590 3884 7642
rect 3908 7590 3918 7642
rect 3918 7590 3964 7642
rect 3668 7588 3724 7590
rect 3748 7588 3804 7590
rect 3828 7588 3884 7590
rect 3908 7588 3964 7590
rect 4328 11450 4384 11452
rect 4408 11450 4464 11452
rect 4488 11450 4544 11452
rect 4568 11450 4624 11452
rect 4328 11398 4374 11450
rect 4374 11398 4384 11450
rect 4408 11398 4438 11450
rect 4438 11398 4450 11450
rect 4450 11398 4464 11450
rect 4488 11398 4502 11450
rect 4502 11398 4514 11450
rect 4514 11398 4544 11450
rect 4568 11398 4578 11450
rect 4578 11398 4624 11450
rect 4328 11396 4384 11398
rect 4408 11396 4464 11398
rect 4488 11396 4544 11398
rect 4568 11396 4624 11398
rect 4328 10362 4384 10364
rect 4408 10362 4464 10364
rect 4488 10362 4544 10364
rect 4568 10362 4624 10364
rect 4328 10310 4374 10362
rect 4374 10310 4384 10362
rect 4408 10310 4438 10362
rect 4438 10310 4450 10362
rect 4450 10310 4464 10362
rect 4488 10310 4502 10362
rect 4502 10310 4514 10362
rect 4514 10310 4544 10362
rect 4568 10310 4578 10362
rect 4578 10310 4624 10362
rect 4328 10308 4384 10310
rect 4408 10308 4464 10310
rect 4488 10308 4544 10310
rect 4568 10308 4624 10310
rect 4328 9274 4384 9276
rect 4408 9274 4464 9276
rect 4488 9274 4544 9276
rect 4568 9274 4624 9276
rect 4328 9222 4374 9274
rect 4374 9222 4384 9274
rect 4408 9222 4438 9274
rect 4438 9222 4450 9274
rect 4450 9222 4464 9274
rect 4488 9222 4502 9274
rect 4502 9222 4514 9274
rect 4514 9222 4544 9274
rect 4568 9222 4578 9274
rect 4578 9222 4624 9274
rect 4328 9220 4384 9222
rect 4408 9220 4464 9222
rect 4488 9220 4544 9222
rect 4568 9220 4624 9222
rect 4526 8880 4582 8936
rect 4328 8186 4384 8188
rect 4408 8186 4464 8188
rect 4488 8186 4544 8188
rect 4568 8186 4624 8188
rect 4328 8134 4374 8186
rect 4374 8134 4384 8186
rect 4408 8134 4438 8186
rect 4438 8134 4450 8186
rect 4450 8134 4464 8186
rect 4488 8134 4502 8186
rect 4502 8134 4514 8186
rect 4514 8134 4544 8186
rect 4568 8134 4578 8186
rect 4578 8134 4624 8186
rect 4328 8132 4384 8134
rect 4408 8132 4464 8134
rect 4488 8132 4544 8134
rect 4568 8132 4624 8134
rect 4328 7098 4384 7100
rect 4408 7098 4464 7100
rect 4488 7098 4544 7100
rect 4568 7098 4624 7100
rect 4328 7046 4374 7098
rect 4374 7046 4384 7098
rect 4408 7046 4438 7098
rect 4438 7046 4450 7098
rect 4450 7046 4464 7098
rect 4488 7046 4502 7098
rect 4502 7046 4514 7098
rect 4514 7046 4544 7098
rect 4568 7046 4578 7098
rect 4578 7046 4624 7098
rect 4328 7044 4384 7046
rect 4408 7044 4464 7046
rect 4488 7044 4544 7046
rect 4568 7044 4624 7046
rect 5262 16904 5318 16960
rect 6642 31184 6698 31240
rect 6550 30232 6606 30288
rect 7010 31456 7066 31512
rect 7286 35556 7342 35592
rect 7286 35536 7288 35556
rect 7288 35536 7340 35556
rect 7340 35536 7342 35556
rect 7470 35944 7526 36000
rect 7286 32680 7342 32736
rect 7286 32272 7342 32328
rect 7102 30640 7158 30696
rect 6458 29008 6514 29064
rect 6366 28872 6422 28928
rect 6274 28736 6330 28792
rect 6274 28364 6276 28384
rect 6276 28364 6328 28384
rect 6328 28364 6330 28384
rect 6274 28328 6330 28364
rect 6182 26424 6238 26480
rect 6090 23316 6146 23352
rect 6090 23296 6092 23316
rect 6092 23296 6144 23316
rect 6144 23296 6146 23316
rect 6090 22208 6146 22264
rect 6274 24520 6330 24576
rect 6274 24384 6330 24440
rect 6642 27784 6698 27840
rect 6550 27512 6606 27568
rect 7102 30132 7104 30152
rect 7104 30132 7156 30152
rect 7156 30132 7158 30152
rect 7102 30096 7158 30132
rect 6918 27648 6974 27704
rect 8666 39208 8722 39264
rect 9310 40160 9366 40216
rect 8482 38256 8538 38312
rect 8666 38292 8668 38312
rect 8668 38292 8720 38312
rect 8720 38292 8722 38312
rect 8666 38256 8722 38292
rect 8666 38156 8668 38176
rect 8668 38156 8720 38176
rect 8720 38156 8722 38176
rect 8666 38120 8722 38156
rect 9034 38412 9090 38448
rect 9034 38392 9036 38412
rect 9036 38392 9088 38412
rect 9088 38392 9090 38412
rect 8390 37304 8446 37360
rect 8482 37168 8538 37224
rect 8850 37712 8906 37768
rect 8758 37032 8814 37088
rect 8758 36916 8814 36952
rect 8758 36896 8760 36916
rect 8760 36896 8812 36916
rect 8812 36896 8814 36916
rect 8206 36252 8208 36272
rect 8208 36252 8260 36272
rect 8260 36252 8262 36272
rect 8206 36216 8262 36252
rect 8206 36100 8262 36136
rect 8206 36080 8208 36100
rect 8208 36080 8260 36100
rect 8260 36080 8262 36100
rect 8942 37032 8998 37088
rect 9678 41112 9734 41168
rect 10728 43002 10784 43004
rect 10808 43002 10864 43004
rect 10888 43002 10944 43004
rect 10968 43002 11024 43004
rect 10728 42950 10774 43002
rect 10774 42950 10784 43002
rect 10808 42950 10838 43002
rect 10838 42950 10850 43002
rect 10850 42950 10864 43002
rect 10888 42950 10902 43002
rect 10902 42950 10914 43002
rect 10914 42950 10944 43002
rect 10968 42950 10978 43002
rect 10978 42950 11024 43002
rect 10728 42948 10784 42950
rect 10808 42948 10864 42950
rect 10888 42948 10944 42950
rect 10968 42948 11024 42950
rect 10068 42458 10124 42460
rect 10148 42458 10204 42460
rect 10228 42458 10284 42460
rect 10308 42458 10364 42460
rect 10068 42406 10114 42458
rect 10114 42406 10124 42458
rect 10148 42406 10178 42458
rect 10178 42406 10190 42458
rect 10190 42406 10204 42458
rect 10228 42406 10242 42458
rect 10242 42406 10254 42458
rect 10254 42406 10284 42458
rect 10308 42406 10318 42458
rect 10318 42406 10364 42458
rect 10068 42404 10124 42406
rect 10148 42404 10204 42406
rect 10228 42404 10284 42406
rect 10308 42404 10364 42406
rect 9402 39752 9458 39808
rect 10414 41656 10470 41712
rect 10728 41914 10784 41916
rect 10808 41914 10864 41916
rect 10888 41914 10944 41916
rect 10968 41914 11024 41916
rect 10728 41862 10774 41914
rect 10774 41862 10784 41914
rect 10808 41862 10838 41914
rect 10838 41862 10850 41914
rect 10850 41862 10864 41914
rect 10888 41862 10902 41914
rect 10902 41862 10914 41914
rect 10914 41862 10944 41914
rect 10968 41862 10978 41914
rect 10978 41862 11024 41914
rect 10728 41860 10784 41862
rect 10808 41860 10864 41862
rect 10888 41860 10944 41862
rect 10968 41860 11024 41862
rect 10782 41520 10838 41576
rect 10068 41370 10124 41372
rect 10148 41370 10204 41372
rect 10228 41370 10284 41372
rect 10308 41370 10364 41372
rect 10068 41318 10114 41370
rect 10114 41318 10124 41370
rect 10148 41318 10178 41370
rect 10178 41318 10190 41370
rect 10190 41318 10204 41370
rect 10228 41318 10242 41370
rect 10242 41318 10254 41370
rect 10254 41318 10284 41370
rect 10308 41318 10318 41370
rect 10318 41318 10364 41370
rect 10068 41316 10124 41318
rect 10148 41316 10204 41318
rect 10228 41316 10284 41318
rect 10308 41316 10364 41318
rect 9954 40840 10010 40896
rect 9218 38664 9274 38720
rect 9402 38392 9458 38448
rect 9402 38256 9458 38312
rect 9402 37984 9458 38040
rect 9218 37748 9220 37768
rect 9220 37748 9272 37768
rect 9272 37748 9274 37768
rect 9218 37712 9274 37748
rect 10068 40282 10124 40284
rect 10148 40282 10204 40284
rect 10228 40282 10284 40284
rect 10308 40282 10364 40284
rect 10068 40230 10114 40282
rect 10114 40230 10124 40282
rect 10148 40230 10178 40282
rect 10178 40230 10190 40282
rect 10190 40230 10204 40282
rect 10228 40230 10242 40282
rect 10242 40230 10254 40282
rect 10254 40230 10284 40282
rect 10308 40230 10318 40282
rect 10318 40230 10364 40282
rect 10068 40228 10124 40230
rect 10148 40228 10204 40230
rect 10228 40228 10284 40230
rect 10308 40228 10364 40230
rect 10138 39908 10194 39944
rect 10138 39888 10140 39908
rect 10140 39888 10192 39908
rect 10192 39888 10194 39908
rect 9954 39616 10010 39672
rect 10046 39344 10102 39400
rect 10068 39194 10124 39196
rect 10148 39194 10204 39196
rect 10228 39194 10284 39196
rect 10308 39194 10364 39196
rect 10068 39142 10114 39194
rect 10114 39142 10124 39194
rect 10148 39142 10178 39194
rect 10178 39142 10190 39194
rect 10190 39142 10204 39194
rect 10228 39142 10242 39194
rect 10242 39142 10254 39194
rect 10254 39142 10284 39194
rect 10308 39142 10318 39194
rect 10318 39142 10364 39194
rect 10068 39140 10124 39142
rect 10148 39140 10204 39142
rect 10228 39140 10284 39142
rect 10308 39140 10364 39142
rect 9770 38664 9826 38720
rect 9678 38392 9734 38448
rect 9770 38256 9826 38312
rect 9586 37984 9642 38040
rect 8942 36624 8998 36680
rect 8942 36488 8998 36544
rect 9034 36216 9090 36272
rect 9218 36760 9274 36816
rect 8666 35808 8722 35864
rect 8114 35556 8170 35592
rect 8114 35536 8116 35556
rect 8116 35536 8168 35556
rect 8168 35536 8170 35556
rect 8298 35536 8354 35592
rect 7562 33360 7618 33416
rect 7562 32136 7618 32192
rect 7654 31592 7710 31648
rect 7654 31320 7710 31376
rect 7562 31048 7618 31104
rect 7562 30368 7618 30424
rect 7470 30232 7526 30288
rect 7194 28600 7250 28656
rect 7102 28056 7158 28112
rect 6734 27376 6790 27432
rect 6734 27240 6790 27296
rect 6550 26424 6606 26480
rect 6642 25336 6698 25392
rect 6366 24248 6422 24304
rect 6642 24384 6698 24440
rect 6274 24112 6330 24168
rect 5998 21392 6054 21448
rect 5998 19352 6054 19408
rect 6366 23024 6422 23080
rect 6274 20032 6330 20088
rect 6274 18944 6330 19000
rect 5998 18128 6054 18184
rect 6090 17992 6146 18048
rect 6090 17856 6146 17912
rect 5998 17584 6054 17640
rect 5262 12416 5318 12472
rect 6090 16632 6146 16688
rect 6734 24112 6790 24168
rect 6734 23704 6790 23760
rect 7194 27240 7250 27296
rect 7010 25608 7066 25664
rect 7930 34176 7986 34232
rect 8298 35128 8354 35184
rect 8206 34584 8262 34640
rect 7838 32136 7894 32192
rect 7930 31864 7986 31920
rect 7838 31184 7894 31240
rect 7378 26580 7434 26616
rect 7378 26560 7380 26580
rect 7380 26560 7432 26580
rect 7432 26560 7434 26580
rect 7102 24792 7158 24848
rect 8390 34060 8446 34096
rect 8390 34040 8392 34060
rect 8392 34040 8444 34060
rect 8444 34040 8446 34060
rect 8574 34720 8630 34776
rect 8758 34584 8814 34640
rect 9034 35808 9090 35864
rect 9126 35672 9182 35728
rect 9126 35400 9182 35456
rect 9034 33496 9090 33552
rect 8298 32544 8354 32600
rect 8390 32000 8446 32056
rect 8114 30232 8170 30288
rect 8758 32544 8814 32600
rect 8942 32716 8944 32736
rect 8944 32716 8996 32736
rect 8996 32716 8998 32736
rect 8942 32680 8998 32716
rect 8850 32000 8906 32056
rect 8850 30504 8906 30560
rect 8942 30132 8944 30152
rect 8944 30132 8996 30152
rect 8996 30132 8998 30152
rect 8942 30096 8998 30132
rect 8850 29996 8852 30016
rect 8852 29996 8904 30016
rect 8904 29996 8906 30016
rect 8850 29960 8906 29996
rect 9126 32952 9182 33008
rect 10230 38936 10286 38992
rect 10138 38800 10194 38856
rect 10414 38800 10470 38856
rect 10874 40976 10930 41032
rect 10728 40826 10784 40828
rect 10808 40826 10864 40828
rect 10888 40826 10944 40828
rect 10968 40826 11024 40828
rect 10728 40774 10774 40826
rect 10774 40774 10784 40826
rect 10808 40774 10838 40826
rect 10838 40774 10850 40826
rect 10850 40774 10864 40826
rect 10888 40774 10902 40826
rect 10902 40774 10914 40826
rect 10914 40774 10944 40826
rect 10968 40774 10978 40826
rect 10978 40774 11024 40826
rect 10728 40772 10784 40774
rect 10808 40772 10864 40774
rect 10888 40772 10944 40774
rect 10968 40772 11024 40774
rect 10690 40180 10746 40216
rect 10690 40160 10692 40180
rect 10692 40160 10744 40180
rect 10744 40160 10746 40180
rect 11150 40024 11206 40080
rect 11426 40024 11482 40080
rect 10874 39888 10930 39944
rect 10728 39738 10784 39740
rect 10808 39738 10864 39740
rect 10888 39738 10944 39740
rect 10968 39738 11024 39740
rect 10728 39686 10774 39738
rect 10774 39686 10784 39738
rect 10808 39686 10838 39738
rect 10838 39686 10850 39738
rect 10850 39686 10864 39738
rect 10888 39686 10902 39738
rect 10902 39686 10914 39738
rect 10914 39686 10944 39738
rect 10968 39686 10978 39738
rect 10978 39686 11024 39738
rect 10728 39684 10784 39686
rect 10808 39684 10864 39686
rect 10888 39684 10944 39686
rect 10968 39684 11024 39686
rect 10690 39480 10746 39536
rect 10728 38650 10784 38652
rect 10808 38650 10864 38652
rect 10888 38650 10944 38652
rect 10968 38650 11024 38652
rect 10728 38598 10774 38650
rect 10774 38598 10784 38650
rect 10808 38598 10838 38650
rect 10838 38598 10850 38650
rect 10850 38598 10864 38650
rect 10888 38598 10902 38650
rect 10902 38598 10914 38650
rect 10914 38598 10944 38650
rect 10968 38598 10978 38650
rect 10978 38598 11024 38650
rect 10728 38596 10784 38598
rect 10808 38596 10864 38598
rect 10888 38596 10944 38598
rect 10968 38596 11024 38598
rect 10966 38428 10968 38448
rect 10968 38428 11020 38448
rect 11020 38428 11022 38448
rect 10068 38106 10124 38108
rect 10148 38106 10204 38108
rect 10228 38106 10284 38108
rect 10308 38106 10364 38108
rect 10068 38054 10114 38106
rect 10114 38054 10124 38106
rect 10148 38054 10178 38106
rect 10178 38054 10190 38106
rect 10190 38054 10204 38106
rect 10228 38054 10242 38106
rect 10242 38054 10254 38106
rect 10254 38054 10284 38106
rect 10308 38054 10318 38106
rect 10318 38054 10364 38106
rect 10068 38052 10124 38054
rect 10148 38052 10204 38054
rect 10228 38052 10284 38054
rect 10308 38052 10364 38054
rect 10068 37018 10124 37020
rect 10148 37018 10204 37020
rect 10228 37018 10284 37020
rect 10308 37018 10364 37020
rect 10068 36966 10114 37018
rect 10114 36966 10124 37018
rect 10148 36966 10178 37018
rect 10178 36966 10190 37018
rect 10190 36966 10204 37018
rect 10228 36966 10242 37018
rect 10242 36966 10254 37018
rect 10254 36966 10284 37018
rect 10308 36966 10318 37018
rect 10318 36966 10364 37018
rect 10068 36964 10124 36966
rect 10148 36964 10204 36966
rect 10228 36964 10284 36966
rect 10308 36964 10364 36966
rect 10322 36780 10378 36816
rect 10322 36760 10324 36780
rect 10324 36760 10376 36780
rect 10376 36760 10378 36780
rect 9402 36352 9458 36408
rect 9770 36524 9772 36544
rect 9772 36524 9824 36544
rect 9824 36524 9826 36544
rect 9770 36488 9826 36524
rect 9770 36216 9826 36272
rect 9678 35944 9734 36000
rect 9586 35536 9642 35592
rect 10138 36624 10194 36680
rect 10138 36100 10194 36136
rect 10138 36080 10140 36100
rect 10140 36080 10192 36100
rect 10192 36080 10194 36100
rect 10068 35930 10124 35932
rect 10148 35930 10204 35932
rect 10228 35930 10284 35932
rect 10308 35930 10364 35932
rect 10068 35878 10114 35930
rect 10114 35878 10124 35930
rect 10148 35878 10178 35930
rect 10178 35878 10190 35930
rect 10190 35878 10204 35930
rect 10228 35878 10242 35930
rect 10242 35878 10254 35930
rect 10254 35878 10284 35930
rect 10308 35878 10318 35930
rect 10318 35878 10364 35930
rect 10068 35876 10124 35878
rect 10148 35876 10204 35878
rect 10228 35876 10284 35878
rect 10308 35876 10364 35878
rect 10966 38392 11022 38428
rect 10598 37848 10654 37904
rect 10728 37562 10784 37564
rect 10808 37562 10864 37564
rect 10888 37562 10944 37564
rect 10968 37562 11024 37564
rect 10728 37510 10774 37562
rect 10774 37510 10784 37562
rect 10808 37510 10838 37562
rect 10838 37510 10850 37562
rect 10850 37510 10864 37562
rect 10888 37510 10902 37562
rect 10902 37510 10914 37562
rect 10914 37510 10944 37562
rect 10968 37510 10978 37562
rect 10978 37510 11024 37562
rect 10728 37508 10784 37510
rect 10808 37508 10864 37510
rect 10888 37508 10944 37510
rect 10968 37508 11024 37510
rect 9678 34060 9734 34096
rect 10046 35128 10102 35184
rect 10322 35536 10378 35592
rect 10690 36624 10746 36680
rect 10728 36474 10784 36476
rect 10808 36474 10864 36476
rect 10888 36474 10944 36476
rect 10968 36474 11024 36476
rect 10728 36422 10774 36474
rect 10774 36422 10784 36474
rect 10808 36422 10838 36474
rect 10838 36422 10850 36474
rect 10850 36422 10864 36474
rect 10888 36422 10902 36474
rect 10902 36422 10914 36474
rect 10914 36422 10944 36474
rect 10968 36422 10978 36474
rect 10978 36422 11024 36474
rect 10728 36420 10784 36422
rect 10808 36420 10864 36422
rect 10888 36420 10944 36422
rect 10968 36420 11024 36422
rect 10598 35672 10654 35728
rect 10966 36216 11022 36272
rect 10874 36080 10930 36136
rect 10414 35400 10470 35456
rect 10068 34842 10124 34844
rect 10148 34842 10204 34844
rect 10228 34842 10284 34844
rect 10308 34842 10364 34844
rect 10068 34790 10114 34842
rect 10114 34790 10124 34842
rect 10148 34790 10178 34842
rect 10178 34790 10190 34842
rect 10190 34790 10204 34842
rect 10228 34790 10242 34842
rect 10242 34790 10254 34842
rect 10254 34790 10284 34842
rect 10308 34790 10318 34842
rect 10318 34790 10364 34842
rect 10068 34788 10124 34790
rect 10148 34788 10204 34790
rect 10228 34788 10284 34790
rect 10308 34788 10364 34790
rect 10046 34076 10048 34096
rect 10048 34076 10100 34096
rect 10100 34076 10102 34096
rect 9678 34040 9680 34060
rect 9680 34040 9732 34060
rect 9732 34040 9734 34060
rect 10046 34040 10102 34076
rect 9678 33904 9734 33960
rect 9678 32444 9680 32464
rect 9680 32444 9732 32464
rect 9732 32444 9734 32464
rect 9678 32408 9734 32444
rect 9678 32136 9734 32192
rect 10068 33754 10124 33756
rect 10148 33754 10204 33756
rect 10228 33754 10284 33756
rect 10308 33754 10364 33756
rect 10068 33702 10114 33754
rect 10114 33702 10124 33754
rect 10148 33702 10178 33754
rect 10178 33702 10190 33754
rect 10190 33702 10204 33754
rect 10228 33702 10242 33754
rect 10242 33702 10254 33754
rect 10254 33702 10284 33754
rect 10308 33702 10318 33754
rect 10318 33702 10364 33754
rect 10068 33700 10124 33702
rect 10148 33700 10204 33702
rect 10228 33700 10284 33702
rect 10308 33700 10364 33702
rect 9862 32544 9918 32600
rect 10728 35386 10784 35388
rect 10808 35386 10864 35388
rect 10888 35386 10944 35388
rect 10968 35386 11024 35388
rect 10728 35334 10774 35386
rect 10774 35334 10784 35386
rect 10808 35334 10838 35386
rect 10838 35334 10850 35386
rect 10850 35334 10864 35386
rect 10888 35334 10902 35386
rect 10902 35334 10914 35386
rect 10914 35334 10944 35386
rect 10968 35334 10978 35386
rect 10978 35334 11024 35386
rect 10728 35332 10784 35334
rect 10808 35332 10864 35334
rect 10888 35332 10944 35334
rect 10968 35332 11024 35334
rect 10728 34298 10784 34300
rect 10808 34298 10864 34300
rect 10888 34298 10944 34300
rect 10968 34298 11024 34300
rect 10728 34246 10774 34298
rect 10774 34246 10784 34298
rect 10808 34246 10838 34298
rect 10838 34246 10850 34298
rect 10850 34246 10864 34298
rect 10888 34246 10902 34298
rect 10902 34246 10914 34298
rect 10914 34246 10944 34298
rect 10968 34246 10978 34298
rect 10978 34246 11024 34298
rect 10728 34244 10784 34246
rect 10808 34244 10864 34246
rect 10888 34244 10944 34246
rect 10968 34244 11024 34246
rect 11242 38936 11298 38992
rect 11242 38120 11298 38176
rect 11150 37576 11206 37632
rect 11150 37304 11206 37360
rect 11242 37204 11244 37224
rect 11244 37204 11296 37224
rect 11296 37204 11298 37224
rect 11242 37168 11298 37204
rect 11150 36760 11206 36816
rect 11150 34448 11206 34504
rect 11426 38292 11428 38312
rect 11428 38292 11480 38312
rect 11480 38292 11482 38312
rect 11426 38256 11482 38292
rect 11426 38120 11482 38176
rect 11426 36896 11482 36952
rect 11426 36080 11482 36136
rect 11886 41928 11942 41984
rect 10506 33496 10562 33552
rect 10068 32666 10124 32668
rect 10148 32666 10204 32668
rect 10228 32666 10284 32668
rect 10308 32666 10364 32668
rect 10068 32614 10114 32666
rect 10114 32614 10124 32666
rect 10148 32614 10178 32666
rect 10178 32614 10190 32666
rect 10190 32614 10204 32666
rect 10228 32614 10242 32666
rect 10242 32614 10254 32666
rect 10254 32614 10284 32666
rect 10308 32614 10318 32666
rect 10318 32614 10364 32666
rect 10068 32612 10124 32614
rect 10148 32612 10204 32614
rect 10228 32612 10284 32614
rect 10308 32612 10364 32614
rect 10322 32408 10378 32464
rect 9586 32000 9642 32056
rect 9678 31728 9734 31784
rect 9402 31592 9458 31648
rect 9310 31456 9366 31512
rect 8850 29008 8906 29064
rect 8390 28056 8446 28112
rect 8942 28192 8998 28248
rect 8022 26968 8078 27024
rect 8022 25744 8078 25800
rect 8574 27512 8630 27568
rect 8390 26152 8446 26208
rect 8114 25336 8170 25392
rect 6918 23160 6974 23216
rect 7194 24520 7250 24576
rect 7286 24112 7342 24168
rect 6826 23024 6882 23080
rect 6734 22208 6790 22264
rect 6734 21936 6790 21992
rect 6550 21564 6552 21584
rect 6552 21564 6604 21584
rect 6604 21564 6606 21584
rect 6550 21528 6606 21564
rect 7286 22072 7342 22128
rect 6458 19252 6460 19272
rect 6460 19252 6512 19272
rect 6512 19252 6514 19272
rect 6458 19216 6514 19252
rect 6826 19216 6882 19272
rect 6734 18808 6790 18864
rect 7194 20712 7250 20768
rect 7654 23704 7710 23760
rect 7930 24148 7932 24168
rect 7932 24148 7984 24168
rect 7984 24148 7986 24168
rect 7930 24112 7986 24148
rect 8298 24112 8354 24168
rect 8206 23432 8262 23488
rect 7470 21256 7526 21312
rect 7378 20848 7434 20904
rect 7378 20576 7434 20632
rect 7378 20168 7434 20224
rect 7010 18828 7066 18864
rect 7010 18808 7012 18828
rect 7012 18808 7064 18828
rect 7064 18808 7066 18828
rect 6458 17584 6514 17640
rect 6366 17040 6422 17096
rect 6642 17176 6698 17232
rect 8574 25880 8630 25936
rect 8574 25064 8630 25120
rect 8574 24520 8630 24576
rect 8114 22092 8170 22128
rect 8114 22072 8116 22092
rect 8116 22072 8168 22092
rect 8168 22072 8170 22092
rect 8390 22888 8446 22944
rect 8482 22208 8538 22264
rect 8390 22072 8446 22128
rect 8114 21528 8170 21584
rect 7654 18944 7710 19000
rect 6550 17076 6552 17096
rect 6552 17076 6604 17096
rect 6604 17076 6606 17096
rect 6550 17040 6606 17076
rect 6734 17040 6790 17096
rect 6550 16632 6606 16688
rect 6458 16532 6460 16552
rect 6460 16532 6512 16552
rect 6512 16532 6514 16552
rect 6458 16496 6514 16532
rect 6550 16224 6606 16280
rect 5262 12280 5318 12336
rect 4802 9988 4858 10024
rect 4802 9968 4804 9988
rect 4804 9968 4856 9988
rect 4856 9968 4858 9988
rect 4894 8372 4896 8392
rect 4896 8372 4948 8392
rect 4948 8372 4950 8392
rect 4894 8336 4950 8372
rect 3668 6554 3724 6556
rect 3748 6554 3804 6556
rect 3828 6554 3884 6556
rect 3908 6554 3964 6556
rect 3668 6502 3714 6554
rect 3714 6502 3724 6554
rect 3748 6502 3778 6554
rect 3778 6502 3790 6554
rect 3790 6502 3804 6554
rect 3828 6502 3842 6554
rect 3842 6502 3854 6554
rect 3854 6502 3884 6554
rect 3908 6502 3918 6554
rect 3918 6502 3964 6554
rect 3668 6500 3724 6502
rect 3748 6500 3804 6502
rect 3828 6500 3884 6502
rect 3908 6500 3964 6502
rect 3422 5772 3478 5808
rect 3422 5752 3424 5772
rect 3424 5752 3476 5772
rect 3476 5752 3478 5772
rect 3668 5466 3724 5468
rect 3748 5466 3804 5468
rect 3828 5466 3884 5468
rect 3908 5466 3964 5468
rect 3668 5414 3714 5466
rect 3714 5414 3724 5466
rect 3748 5414 3778 5466
rect 3778 5414 3790 5466
rect 3790 5414 3804 5466
rect 3828 5414 3842 5466
rect 3842 5414 3854 5466
rect 3854 5414 3884 5466
rect 3908 5414 3918 5466
rect 3918 5414 3964 5466
rect 3668 5412 3724 5414
rect 3748 5412 3804 5414
rect 3828 5412 3884 5414
rect 3908 5412 3964 5414
rect 4328 6010 4384 6012
rect 4408 6010 4464 6012
rect 4488 6010 4544 6012
rect 4568 6010 4624 6012
rect 4328 5958 4374 6010
rect 4374 5958 4384 6010
rect 4408 5958 4438 6010
rect 4438 5958 4450 6010
rect 4450 5958 4464 6010
rect 4488 5958 4502 6010
rect 4502 5958 4514 6010
rect 4514 5958 4544 6010
rect 4568 5958 4578 6010
rect 4578 5958 4624 6010
rect 4328 5956 4384 5958
rect 4408 5956 4464 5958
rect 4488 5956 4544 5958
rect 4568 5956 4624 5958
rect 5538 8628 5594 8664
rect 5538 8608 5540 8628
rect 5540 8608 5592 8628
rect 5592 8608 5594 8628
rect 7194 17992 7250 18048
rect 7562 17584 7618 17640
rect 7378 16632 7434 16688
rect 7286 16516 7342 16552
rect 7286 16496 7288 16516
rect 7288 16496 7340 16516
rect 7340 16496 7342 16516
rect 6366 13776 6422 13832
rect 6182 13640 6238 13696
rect 6090 12688 6146 12744
rect 3668 4378 3724 4380
rect 3748 4378 3804 4380
rect 3828 4378 3884 4380
rect 3908 4378 3964 4380
rect 3668 4326 3714 4378
rect 3714 4326 3724 4378
rect 3748 4326 3778 4378
rect 3778 4326 3790 4378
rect 3790 4326 3804 4378
rect 3828 4326 3842 4378
rect 3842 4326 3854 4378
rect 3854 4326 3884 4378
rect 3908 4326 3918 4378
rect 3918 4326 3964 4378
rect 3668 4324 3724 4326
rect 3748 4324 3804 4326
rect 3828 4324 3884 4326
rect 3908 4324 3964 4326
rect 4328 4922 4384 4924
rect 4408 4922 4464 4924
rect 4488 4922 4544 4924
rect 4568 4922 4624 4924
rect 4328 4870 4374 4922
rect 4374 4870 4384 4922
rect 4408 4870 4438 4922
rect 4438 4870 4450 4922
rect 4450 4870 4464 4922
rect 4488 4870 4502 4922
rect 4502 4870 4514 4922
rect 4514 4870 4544 4922
rect 4568 4870 4578 4922
rect 4578 4870 4624 4922
rect 4328 4868 4384 4870
rect 4408 4868 4464 4870
rect 4488 4868 4544 4870
rect 4568 4868 4624 4870
rect 2502 1400 2558 1456
rect 4328 3834 4384 3836
rect 4408 3834 4464 3836
rect 4488 3834 4544 3836
rect 4568 3834 4624 3836
rect 4328 3782 4374 3834
rect 4374 3782 4384 3834
rect 4408 3782 4438 3834
rect 4438 3782 4450 3834
rect 4450 3782 4464 3834
rect 4488 3782 4502 3834
rect 4502 3782 4514 3834
rect 4514 3782 4544 3834
rect 4568 3782 4578 3834
rect 4578 3782 4624 3834
rect 4328 3780 4384 3782
rect 4408 3780 4464 3782
rect 4488 3780 4544 3782
rect 4568 3780 4624 3782
rect 3668 3290 3724 3292
rect 3748 3290 3804 3292
rect 3828 3290 3884 3292
rect 3908 3290 3964 3292
rect 3668 3238 3714 3290
rect 3714 3238 3724 3290
rect 3748 3238 3778 3290
rect 3778 3238 3790 3290
rect 3790 3238 3804 3290
rect 3828 3238 3842 3290
rect 3842 3238 3854 3290
rect 3854 3238 3884 3290
rect 3908 3238 3918 3290
rect 3918 3238 3964 3290
rect 3668 3236 3724 3238
rect 3748 3236 3804 3238
rect 3828 3236 3884 3238
rect 3908 3236 3964 3238
rect 3668 2202 3724 2204
rect 3748 2202 3804 2204
rect 3828 2202 3884 2204
rect 3908 2202 3964 2204
rect 3668 2150 3714 2202
rect 3714 2150 3724 2202
rect 3748 2150 3778 2202
rect 3778 2150 3790 2202
rect 3790 2150 3804 2202
rect 3828 2150 3842 2202
rect 3842 2150 3854 2202
rect 3854 2150 3884 2202
rect 3908 2150 3918 2202
rect 3918 2150 3964 2202
rect 3668 2148 3724 2150
rect 3748 2148 3804 2150
rect 3828 2148 3884 2150
rect 3908 2148 3964 2150
rect 4328 2746 4384 2748
rect 4408 2746 4464 2748
rect 4488 2746 4544 2748
rect 4568 2746 4624 2748
rect 4328 2694 4374 2746
rect 4374 2694 4384 2746
rect 4408 2694 4438 2746
rect 4438 2694 4450 2746
rect 4450 2694 4464 2746
rect 4488 2694 4502 2746
rect 4502 2694 4514 2746
rect 4514 2694 4544 2746
rect 4568 2694 4578 2746
rect 4578 2694 4624 2746
rect 4328 2692 4384 2694
rect 4408 2692 4464 2694
rect 4488 2692 4544 2694
rect 4568 2692 4624 2694
rect 4328 1658 4384 1660
rect 4408 1658 4464 1660
rect 4488 1658 4544 1660
rect 4568 1658 4624 1660
rect 4328 1606 4374 1658
rect 4374 1606 4384 1658
rect 4408 1606 4438 1658
rect 4438 1606 4450 1658
rect 4450 1606 4464 1658
rect 4488 1606 4502 1658
rect 4502 1606 4514 1658
rect 4514 1606 4544 1658
rect 4568 1606 4578 1658
rect 4578 1606 4624 1658
rect 4328 1604 4384 1606
rect 4408 1604 4464 1606
rect 4488 1604 4544 1606
rect 4568 1604 4624 1606
rect 3668 1114 3724 1116
rect 3748 1114 3804 1116
rect 3828 1114 3884 1116
rect 3908 1114 3964 1116
rect 3668 1062 3714 1114
rect 3714 1062 3724 1114
rect 3748 1062 3778 1114
rect 3778 1062 3790 1114
rect 3790 1062 3804 1114
rect 3828 1062 3842 1114
rect 3842 1062 3854 1114
rect 3854 1062 3884 1114
rect 3908 1062 3918 1114
rect 3918 1062 3964 1114
rect 3668 1060 3724 1062
rect 3748 1060 3804 1062
rect 3828 1060 3884 1062
rect 3908 1060 3964 1062
rect 6734 12144 6790 12200
rect 7010 12552 7066 12608
rect 7010 12316 7012 12336
rect 7012 12316 7064 12336
rect 7064 12316 7066 12336
rect 7010 12280 7066 12316
rect 7102 12044 7104 12064
rect 7104 12044 7156 12064
rect 7156 12044 7158 12064
rect 7102 12008 7158 12044
rect 7930 19252 7932 19272
rect 7932 19252 7984 19272
rect 7984 19252 7986 19272
rect 7930 19216 7986 19252
rect 7930 18944 7986 19000
rect 8298 20576 8354 20632
rect 8758 24656 8814 24712
rect 9770 31592 9826 31648
rect 9586 28872 9642 28928
rect 9862 30504 9918 30560
rect 9862 30368 9918 30424
rect 10068 31578 10124 31580
rect 10148 31578 10204 31580
rect 10228 31578 10284 31580
rect 10308 31578 10364 31580
rect 10068 31526 10114 31578
rect 10114 31526 10124 31578
rect 10148 31526 10178 31578
rect 10178 31526 10190 31578
rect 10190 31526 10204 31578
rect 10228 31526 10242 31578
rect 10242 31526 10254 31578
rect 10254 31526 10284 31578
rect 10308 31526 10318 31578
rect 10318 31526 10364 31578
rect 10068 31524 10124 31526
rect 10148 31524 10204 31526
rect 10228 31524 10284 31526
rect 10308 31524 10364 31526
rect 11058 33924 11114 33960
rect 11058 33904 11060 33924
rect 11060 33904 11112 33924
rect 11112 33904 11114 33924
rect 10728 33210 10784 33212
rect 10808 33210 10864 33212
rect 10888 33210 10944 33212
rect 10968 33210 11024 33212
rect 10728 33158 10774 33210
rect 10774 33158 10784 33210
rect 10808 33158 10838 33210
rect 10838 33158 10850 33210
rect 10850 33158 10864 33210
rect 10888 33158 10902 33210
rect 10902 33158 10914 33210
rect 10914 33158 10944 33210
rect 10968 33158 10978 33210
rect 10978 33158 11024 33210
rect 10728 33156 10784 33158
rect 10808 33156 10864 33158
rect 10888 33156 10944 33158
rect 10968 33156 11024 33158
rect 10506 32408 10562 32464
rect 10230 30812 10232 30832
rect 10232 30812 10284 30832
rect 10284 30812 10286 30832
rect 10230 30776 10286 30812
rect 10046 30640 10102 30696
rect 10068 30490 10124 30492
rect 10148 30490 10204 30492
rect 10228 30490 10284 30492
rect 10308 30490 10364 30492
rect 10068 30438 10114 30490
rect 10114 30438 10124 30490
rect 10148 30438 10178 30490
rect 10178 30438 10190 30490
rect 10190 30438 10204 30490
rect 10228 30438 10242 30490
rect 10242 30438 10254 30490
rect 10254 30438 10284 30490
rect 10308 30438 10318 30490
rect 10318 30438 10364 30490
rect 10068 30436 10124 30438
rect 10148 30436 10204 30438
rect 10228 30436 10284 30438
rect 10308 30436 10364 30438
rect 10230 30268 10232 30288
rect 10232 30268 10284 30288
rect 10284 30268 10286 30288
rect 10230 30232 10286 30268
rect 10046 30096 10102 30152
rect 9862 29552 9918 29608
rect 9862 29144 9918 29200
rect 10138 29844 10194 29880
rect 10138 29824 10140 29844
rect 10140 29824 10192 29844
rect 10192 29824 10194 29844
rect 10230 29688 10286 29744
rect 10230 29588 10232 29608
rect 10232 29588 10284 29608
rect 10284 29588 10286 29608
rect 10230 29552 10286 29588
rect 10068 29402 10124 29404
rect 10148 29402 10204 29404
rect 10228 29402 10284 29404
rect 10308 29402 10364 29404
rect 10068 29350 10114 29402
rect 10114 29350 10124 29402
rect 10148 29350 10178 29402
rect 10178 29350 10190 29402
rect 10190 29350 10204 29402
rect 10228 29350 10242 29402
rect 10242 29350 10254 29402
rect 10254 29350 10284 29402
rect 10308 29350 10318 29402
rect 10318 29350 10364 29402
rect 10068 29348 10124 29350
rect 10148 29348 10204 29350
rect 10228 29348 10284 29350
rect 10308 29348 10364 29350
rect 10874 32952 10930 33008
rect 10728 32122 10784 32124
rect 10808 32122 10864 32124
rect 10888 32122 10944 32124
rect 10968 32122 11024 32124
rect 10728 32070 10774 32122
rect 10774 32070 10784 32122
rect 10808 32070 10838 32122
rect 10838 32070 10850 32122
rect 10850 32070 10864 32122
rect 10888 32070 10902 32122
rect 10902 32070 10914 32122
rect 10914 32070 10944 32122
rect 10968 32070 10978 32122
rect 10978 32070 11024 32122
rect 10728 32068 10784 32070
rect 10808 32068 10864 32070
rect 10888 32068 10944 32070
rect 10968 32068 11024 32070
rect 10690 31628 10692 31648
rect 10692 31628 10744 31648
rect 10744 31628 10746 31648
rect 10690 31592 10746 31628
rect 10728 31034 10784 31036
rect 10808 31034 10864 31036
rect 10888 31034 10944 31036
rect 10968 31034 11024 31036
rect 10728 30982 10774 31034
rect 10774 30982 10784 31034
rect 10808 30982 10838 31034
rect 10838 30982 10850 31034
rect 10850 30982 10864 31034
rect 10888 30982 10902 31034
rect 10902 30982 10914 31034
rect 10914 30982 10944 31034
rect 10968 30982 10978 31034
rect 10978 30982 11024 31034
rect 10728 30980 10784 30982
rect 10808 30980 10864 30982
rect 10888 30980 10944 30982
rect 10968 30980 11024 30982
rect 10782 30776 10838 30832
rect 10966 30368 11022 30424
rect 10506 29960 10562 30016
rect 10728 29946 10784 29948
rect 10808 29946 10864 29948
rect 10888 29946 10944 29948
rect 10968 29946 11024 29948
rect 10728 29894 10774 29946
rect 10774 29894 10784 29946
rect 10808 29894 10838 29946
rect 10838 29894 10850 29946
rect 10850 29894 10864 29946
rect 10888 29894 10902 29946
rect 10902 29894 10914 29946
rect 10914 29894 10944 29946
rect 10968 29894 10978 29946
rect 10978 29894 11024 29946
rect 10728 29892 10784 29894
rect 10808 29892 10864 29894
rect 10888 29892 10944 29894
rect 10968 29892 11024 29894
rect 10690 29688 10746 29744
rect 10598 29416 10654 29472
rect 10598 29144 10654 29200
rect 9126 26560 9182 26616
rect 9126 24692 9128 24712
rect 9128 24692 9180 24712
rect 9180 24692 9182 24712
rect 9126 24656 9182 24692
rect 9034 24112 9090 24168
rect 8942 22616 8998 22672
rect 9586 27512 9642 27568
rect 9678 27376 9734 27432
rect 9678 27104 9734 27160
rect 9218 21800 9274 21856
rect 9034 20984 9090 21040
rect 8298 19780 8354 19816
rect 8298 19760 8300 19780
rect 8300 19760 8352 19780
rect 8352 19760 8354 19780
rect 7930 17720 7986 17776
rect 7838 16632 7894 16688
rect 7654 16496 7710 16552
rect 7378 12280 7434 12336
rect 7838 15020 7894 15056
rect 7838 15000 7840 15020
rect 7840 15000 7892 15020
rect 7892 15000 7894 15020
rect 7746 12844 7802 12880
rect 7746 12824 7748 12844
rect 7748 12824 7800 12844
rect 7800 12824 7802 12844
rect 8482 19352 8538 19408
rect 8206 17740 8262 17776
rect 8206 17720 8208 17740
rect 8208 17720 8260 17740
rect 8260 17720 8262 17740
rect 8666 19352 8722 19408
rect 10068 28314 10124 28316
rect 10148 28314 10204 28316
rect 10228 28314 10284 28316
rect 10308 28314 10364 28316
rect 10068 28262 10114 28314
rect 10114 28262 10124 28314
rect 10148 28262 10178 28314
rect 10178 28262 10190 28314
rect 10190 28262 10204 28314
rect 10228 28262 10242 28314
rect 10242 28262 10254 28314
rect 10254 28262 10284 28314
rect 10308 28262 10318 28314
rect 10318 28262 10364 28314
rect 10068 28260 10124 28262
rect 10148 28260 10204 28262
rect 10228 28260 10284 28262
rect 10308 28260 10364 28262
rect 10230 28056 10286 28112
rect 11058 29708 11114 29744
rect 11058 29688 11060 29708
rect 11060 29688 11112 29708
rect 11112 29688 11114 29708
rect 11058 29300 11114 29336
rect 11058 29280 11060 29300
rect 11060 29280 11112 29300
rect 11112 29280 11114 29300
rect 10728 28858 10784 28860
rect 10808 28858 10864 28860
rect 10888 28858 10944 28860
rect 10968 28858 11024 28860
rect 10728 28806 10774 28858
rect 10774 28806 10784 28858
rect 10808 28806 10838 28858
rect 10838 28806 10850 28858
rect 10850 28806 10864 28858
rect 10888 28806 10902 28858
rect 10902 28806 10914 28858
rect 10914 28806 10944 28858
rect 10968 28806 10978 28858
rect 10978 28806 11024 28858
rect 10728 28804 10784 28806
rect 10808 28804 10864 28806
rect 10888 28804 10944 28806
rect 10968 28804 11024 28806
rect 10506 28056 10562 28112
rect 11426 34040 11482 34096
rect 11886 39480 11942 39536
rect 11978 37324 12034 37360
rect 11978 37304 11980 37324
rect 11980 37304 12032 37324
rect 12032 37304 12034 37324
rect 11886 37168 11942 37224
rect 11702 35128 11758 35184
rect 12162 36216 12218 36272
rect 11886 34584 11942 34640
rect 11518 33904 11574 33960
rect 11610 32816 11666 32872
rect 11426 31592 11482 31648
rect 11886 33652 11942 33688
rect 11886 33632 11888 33652
rect 11888 33632 11940 33652
rect 11940 33632 11942 33652
rect 11978 33496 12034 33552
rect 11794 32272 11850 32328
rect 11886 32000 11942 32056
rect 11794 31728 11850 31784
rect 11426 30232 11482 30288
rect 11334 29416 11390 29472
rect 10068 27226 10124 27228
rect 10148 27226 10204 27228
rect 10228 27226 10284 27228
rect 10308 27226 10364 27228
rect 10068 27174 10114 27226
rect 10114 27174 10124 27226
rect 10148 27174 10178 27226
rect 10178 27174 10190 27226
rect 10190 27174 10204 27226
rect 10228 27174 10242 27226
rect 10242 27174 10254 27226
rect 10254 27174 10284 27226
rect 10308 27174 10318 27226
rect 10318 27174 10364 27226
rect 10068 27172 10124 27174
rect 10148 27172 10204 27174
rect 10228 27172 10284 27174
rect 10308 27172 10364 27174
rect 10068 26138 10124 26140
rect 10148 26138 10204 26140
rect 10228 26138 10284 26140
rect 10308 26138 10364 26140
rect 10068 26086 10114 26138
rect 10114 26086 10124 26138
rect 10148 26086 10178 26138
rect 10178 26086 10190 26138
rect 10190 26086 10204 26138
rect 10228 26086 10242 26138
rect 10242 26086 10254 26138
rect 10254 26086 10284 26138
rect 10308 26086 10318 26138
rect 10318 26086 10364 26138
rect 10068 26084 10124 26086
rect 10148 26084 10204 26086
rect 10228 26084 10284 26086
rect 10308 26084 10364 26086
rect 11886 30776 11942 30832
rect 12346 37712 12402 37768
rect 10728 27770 10784 27772
rect 10808 27770 10864 27772
rect 10888 27770 10944 27772
rect 10968 27770 11024 27772
rect 10728 27718 10774 27770
rect 10774 27718 10784 27770
rect 10808 27718 10838 27770
rect 10838 27718 10850 27770
rect 10850 27718 10864 27770
rect 10888 27718 10902 27770
rect 10902 27718 10914 27770
rect 10914 27718 10944 27770
rect 10968 27718 10978 27770
rect 10978 27718 11024 27770
rect 10728 27716 10784 27718
rect 10808 27716 10864 27718
rect 10888 27716 10944 27718
rect 10968 27716 11024 27718
rect 10728 26682 10784 26684
rect 10808 26682 10864 26684
rect 10888 26682 10944 26684
rect 10968 26682 11024 26684
rect 10728 26630 10774 26682
rect 10774 26630 10784 26682
rect 10808 26630 10838 26682
rect 10838 26630 10850 26682
rect 10850 26630 10864 26682
rect 10888 26630 10902 26682
rect 10902 26630 10914 26682
rect 10914 26630 10944 26682
rect 10968 26630 10978 26682
rect 10978 26630 11024 26682
rect 10728 26628 10784 26630
rect 10808 26628 10864 26630
rect 10888 26628 10944 26630
rect 10968 26628 11024 26630
rect 10728 25594 10784 25596
rect 10808 25594 10864 25596
rect 10888 25594 10944 25596
rect 10968 25594 11024 25596
rect 10728 25542 10774 25594
rect 10774 25542 10784 25594
rect 10808 25542 10838 25594
rect 10838 25542 10850 25594
rect 10850 25542 10864 25594
rect 10888 25542 10902 25594
rect 10902 25542 10914 25594
rect 10914 25542 10944 25594
rect 10968 25542 10978 25594
rect 10978 25542 11024 25594
rect 10728 25540 10784 25542
rect 10808 25540 10864 25542
rect 10888 25540 10944 25542
rect 10968 25540 11024 25542
rect 10068 25050 10124 25052
rect 10148 25050 10204 25052
rect 10228 25050 10284 25052
rect 10308 25050 10364 25052
rect 10068 24998 10114 25050
rect 10114 24998 10124 25050
rect 10148 24998 10178 25050
rect 10178 24998 10190 25050
rect 10190 24998 10204 25050
rect 10228 24998 10242 25050
rect 10242 24998 10254 25050
rect 10254 24998 10284 25050
rect 10308 24998 10318 25050
rect 10318 24998 10364 25050
rect 10068 24996 10124 24998
rect 10148 24996 10204 24998
rect 10228 24996 10284 24998
rect 10308 24996 10364 24998
rect 9770 24520 9826 24576
rect 9770 23568 9826 23624
rect 9678 23432 9734 23488
rect 10068 23962 10124 23964
rect 10148 23962 10204 23964
rect 10228 23962 10284 23964
rect 10308 23962 10364 23964
rect 10068 23910 10114 23962
rect 10114 23910 10124 23962
rect 10148 23910 10178 23962
rect 10178 23910 10190 23962
rect 10190 23910 10204 23962
rect 10228 23910 10242 23962
rect 10242 23910 10254 23962
rect 10254 23910 10284 23962
rect 10308 23910 10318 23962
rect 10318 23910 10364 23962
rect 10068 23908 10124 23910
rect 10148 23908 10204 23910
rect 10228 23908 10284 23910
rect 10308 23908 10364 23910
rect 10728 24506 10784 24508
rect 10808 24506 10864 24508
rect 10888 24506 10944 24508
rect 10968 24506 11024 24508
rect 10728 24454 10774 24506
rect 10774 24454 10784 24506
rect 10808 24454 10838 24506
rect 10838 24454 10850 24506
rect 10850 24454 10864 24506
rect 10888 24454 10902 24506
rect 10902 24454 10914 24506
rect 10914 24454 10944 24506
rect 10968 24454 10978 24506
rect 10978 24454 11024 24506
rect 10728 24452 10784 24454
rect 10808 24452 10864 24454
rect 10888 24452 10944 24454
rect 10968 24452 11024 24454
rect 10728 23418 10784 23420
rect 10808 23418 10864 23420
rect 10888 23418 10944 23420
rect 10968 23418 11024 23420
rect 10728 23366 10774 23418
rect 10774 23366 10784 23418
rect 10808 23366 10838 23418
rect 10838 23366 10850 23418
rect 10850 23366 10864 23418
rect 10888 23366 10902 23418
rect 10902 23366 10914 23418
rect 10914 23366 10944 23418
rect 10968 23366 10978 23418
rect 10978 23366 11024 23418
rect 10728 23364 10784 23366
rect 10808 23364 10864 23366
rect 10888 23364 10944 23366
rect 10968 23364 11024 23366
rect 10414 23024 10470 23080
rect 10068 22874 10124 22876
rect 10148 22874 10204 22876
rect 10228 22874 10284 22876
rect 10308 22874 10364 22876
rect 10068 22822 10114 22874
rect 10114 22822 10124 22874
rect 10148 22822 10178 22874
rect 10178 22822 10190 22874
rect 10190 22822 10204 22874
rect 10228 22822 10242 22874
rect 10242 22822 10254 22874
rect 10254 22822 10284 22874
rect 10308 22822 10318 22874
rect 10318 22822 10364 22874
rect 10068 22820 10124 22822
rect 10148 22820 10204 22822
rect 10228 22820 10284 22822
rect 10308 22820 10364 22822
rect 9954 22616 10010 22672
rect 10138 22636 10194 22672
rect 10138 22616 10140 22636
rect 10140 22616 10192 22636
rect 10192 22616 10194 22636
rect 10782 22516 10784 22536
rect 10784 22516 10836 22536
rect 10836 22516 10838 22536
rect 10782 22480 10838 22516
rect 10728 22330 10784 22332
rect 10808 22330 10864 22332
rect 10888 22330 10944 22332
rect 10968 22330 11024 22332
rect 10728 22278 10774 22330
rect 10774 22278 10784 22330
rect 10808 22278 10838 22330
rect 10838 22278 10850 22330
rect 10850 22278 10864 22330
rect 10888 22278 10902 22330
rect 10902 22278 10914 22330
rect 10914 22278 10944 22330
rect 10968 22278 10978 22330
rect 10978 22278 11024 22330
rect 10728 22276 10784 22278
rect 10808 22276 10864 22278
rect 10888 22276 10944 22278
rect 10968 22276 11024 22278
rect 10068 21786 10124 21788
rect 10148 21786 10204 21788
rect 10228 21786 10284 21788
rect 10308 21786 10364 21788
rect 10068 21734 10114 21786
rect 10114 21734 10124 21786
rect 10148 21734 10178 21786
rect 10178 21734 10190 21786
rect 10190 21734 10204 21786
rect 10228 21734 10242 21786
rect 10242 21734 10254 21786
rect 10254 21734 10284 21786
rect 10308 21734 10318 21786
rect 10318 21734 10364 21786
rect 10068 21732 10124 21734
rect 10148 21732 10204 21734
rect 10228 21732 10284 21734
rect 10308 21732 10364 21734
rect 9494 20712 9550 20768
rect 9126 20440 9182 20496
rect 9218 20032 9274 20088
rect 9034 19216 9090 19272
rect 8574 17992 8630 18048
rect 8574 17856 8630 17912
rect 8758 17856 8814 17912
rect 8850 17584 8906 17640
rect 8206 15564 8262 15600
rect 8206 15544 8208 15564
rect 8208 15544 8260 15564
rect 8260 15544 8262 15564
rect 8482 15272 8538 15328
rect 7654 12416 7710 12472
rect 7654 12300 7710 12336
rect 7654 12280 7656 12300
rect 7656 12280 7708 12300
rect 7708 12280 7710 12300
rect 7470 8336 7526 8392
rect 8114 12008 8170 12064
rect 8114 11056 8170 11112
rect 8666 12416 8722 12472
rect 9126 17740 9182 17776
rect 9126 17720 9128 17740
rect 9128 17720 9180 17740
rect 9180 17720 9182 17740
rect 9402 17856 9458 17912
rect 9126 17332 9182 17368
rect 9126 17312 9128 17332
rect 9128 17312 9180 17332
rect 9180 17312 9182 17332
rect 8942 15000 8998 15056
rect 9310 16632 9366 16688
rect 8942 12824 8998 12880
rect 9310 14456 9366 14512
rect 11058 22072 11114 22128
rect 10414 21256 10470 21312
rect 10068 20698 10124 20700
rect 10148 20698 10204 20700
rect 10228 20698 10284 20700
rect 10308 20698 10364 20700
rect 10068 20646 10114 20698
rect 10114 20646 10124 20698
rect 10148 20646 10178 20698
rect 10178 20646 10190 20698
rect 10190 20646 10204 20698
rect 10228 20646 10242 20698
rect 10242 20646 10254 20698
rect 10254 20646 10284 20698
rect 10308 20646 10318 20698
rect 10318 20646 10364 20698
rect 10068 20644 10124 20646
rect 10148 20644 10204 20646
rect 10228 20644 10284 20646
rect 10308 20644 10364 20646
rect 10728 21242 10784 21244
rect 10808 21242 10864 21244
rect 10888 21242 10944 21244
rect 10968 21242 11024 21244
rect 10728 21190 10774 21242
rect 10774 21190 10784 21242
rect 10808 21190 10838 21242
rect 10838 21190 10850 21242
rect 10850 21190 10864 21242
rect 10888 21190 10902 21242
rect 10902 21190 10914 21242
rect 10914 21190 10944 21242
rect 10968 21190 10978 21242
rect 10978 21190 11024 21242
rect 10728 21188 10784 21190
rect 10808 21188 10864 21190
rect 10888 21188 10944 21190
rect 10968 21188 11024 21190
rect 11426 26288 11482 26344
rect 12070 28620 12126 28656
rect 12070 28600 12072 28620
rect 12072 28600 12124 28620
rect 12124 28600 12126 28620
rect 12346 32000 12402 32056
rect 12622 31864 12678 31920
rect 12622 29552 12678 29608
rect 12254 27648 12310 27704
rect 11426 23432 11482 23488
rect 11702 23432 11758 23488
rect 11610 22072 11666 22128
rect 10690 20848 10746 20904
rect 10728 20154 10784 20156
rect 10808 20154 10864 20156
rect 10888 20154 10944 20156
rect 10968 20154 11024 20156
rect 10728 20102 10774 20154
rect 10774 20102 10784 20154
rect 10808 20102 10838 20154
rect 10838 20102 10850 20154
rect 10850 20102 10864 20154
rect 10888 20102 10902 20154
rect 10902 20102 10914 20154
rect 10914 20102 10944 20154
rect 10968 20102 10978 20154
rect 10978 20102 11024 20154
rect 10728 20100 10784 20102
rect 10808 20100 10864 20102
rect 10888 20100 10944 20102
rect 10968 20100 11024 20102
rect 10874 19932 10876 19952
rect 10876 19932 10928 19952
rect 10928 19932 10930 19952
rect 10874 19896 10930 19932
rect 10068 19610 10124 19612
rect 10148 19610 10204 19612
rect 10228 19610 10284 19612
rect 10308 19610 10364 19612
rect 10068 19558 10114 19610
rect 10114 19558 10124 19610
rect 10148 19558 10178 19610
rect 10178 19558 10190 19610
rect 10190 19558 10204 19610
rect 10228 19558 10242 19610
rect 10242 19558 10254 19610
rect 10254 19558 10284 19610
rect 10308 19558 10318 19610
rect 10318 19558 10364 19610
rect 10068 19556 10124 19558
rect 10148 19556 10204 19558
rect 10228 19556 10284 19558
rect 10308 19556 10364 19558
rect 10690 19624 10746 19680
rect 10966 19660 10968 19680
rect 10968 19660 11020 19680
rect 11020 19660 11022 19680
rect 10966 19624 11022 19660
rect 10728 19066 10784 19068
rect 10808 19066 10864 19068
rect 10888 19066 10944 19068
rect 10968 19066 11024 19068
rect 10728 19014 10774 19066
rect 10774 19014 10784 19066
rect 10808 19014 10838 19066
rect 10838 19014 10850 19066
rect 10850 19014 10864 19066
rect 10888 19014 10902 19066
rect 10902 19014 10914 19066
rect 10914 19014 10944 19066
rect 10968 19014 10978 19066
rect 10978 19014 11024 19066
rect 10728 19012 10784 19014
rect 10808 19012 10864 19014
rect 10888 19012 10944 19014
rect 10968 19012 11024 19014
rect 9770 17176 9826 17232
rect 9770 16632 9826 16688
rect 9678 16244 9734 16280
rect 9678 16224 9680 16244
rect 9680 16224 9732 16244
rect 9732 16224 9734 16244
rect 9586 16108 9642 16144
rect 9586 16088 9588 16108
rect 9588 16088 9640 16108
rect 9640 16088 9642 16108
rect 10068 18522 10124 18524
rect 10148 18522 10204 18524
rect 10228 18522 10284 18524
rect 10308 18522 10364 18524
rect 10068 18470 10114 18522
rect 10114 18470 10124 18522
rect 10148 18470 10178 18522
rect 10178 18470 10190 18522
rect 10190 18470 10204 18522
rect 10228 18470 10242 18522
rect 10242 18470 10254 18522
rect 10254 18470 10284 18522
rect 10308 18470 10318 18522
rect 10318 18470 10364 18522
rect 10068 18468 10124 18470
rect 10148 18468 10204 18470
rect 10228 18468 10284 18470
rect 10308 18468 10364 18470
rect 10068 17434 10124 17436
rect 10148 17434 10204 17436
rect 10228 17434 10284 17436
rect 10308 17434 10364 17436
rect 10068 17382 10114 17434
rect 10114 17382 10124 17434
rect 10148 17382 10178 17434
rect 10178 17382 10190 17434
rect 10190 17382 10204 17434
rect 10228 17382 10242 17434
rect 10242 17382 10254 17434
rect 10254 17382 10284 17434
rect 10308 17382 10318 17434
rect 10318 17382 10364 17434
rect 10068 17380 10124 17382
rect 10148 17380 10204 17382
rect 10228 17380 10284 17382
rect 10308 17380 10364 17382
rect 9954 17040 10010 17096
rect 12070 22480 12126 22536
rect 11886 19932 11888 19952
rect 11888 19932 11940 19952
rect 11940 19932 11942 19952
rect 11886 19896 11942 19932
rect 10728 17978 10784 17980
rect 10808 17978 10864 17980
rect 10888 17978 10944 17980
rect 10968 17978 11024 17980
rect 10728 17926 10774 17978
rect 10774 17926 10784 17978
rect 10808 17926 10838 17978
rect 10838 17926 10850 17978
rect 10850 17926 10864 17978
rect 10888 17926 10902 17978
rect 10902 17926 10914 17978
rect 10914 17926 10944 17978
rect 10968 17926 10978 17978
rect 10978 17926 11024 17978
rect 10728 17924 10784 17926
rect 10808 17924 10864 17926
rect 10888 17924 10944 17926
rect 10968 17924 11024 17926
rect 11426 17720 11482 17776
rect 10068 16346 10124 16348
rect 10148 16346 10204 16348
rect 10228 16346 10284 16348
rect 10308 16346 10364 16348
rect 10068 16294 10114 16346
rect 10114 16294 10124 16346
rect 10148 16294 10178 16346
rect 10178 16294 10190 16346
rect 10190 16294 10204 16346
rect 10228 16294 10242 16346
rect 10242 16294 10254 16346
rect 10254 16294 10284 16346
rect 10308 16294 10318 16346
rect 10318 16294 10364 16346
rect 10068 16292 10124 16294
rect 10148 16292 10204 16294
rect 10228 16292 10284 16294
rect 10308 16292 10364 16294
rect 9126 12724 9128 12744
rect 9128 12724 9180 12744
rect 9180 12724 9182 12744
rect 9126 12688 9182 12724
rect 9126 12280 9182 12336
rect 8574 7384 8630 7440
rect 7378 1400 7434 1456
rect 10068 15258 10124 15260
rect 10148 15258 10204 15260
rect 10228 15258 10284 15260
rect 10308 15258 10364 15260
rect 10068 15206 10114 15258
rect 10114 15206 10124 15258
rect 10148 15206 10178 15258
rect 10178 15206 10190 15258
rect 10190 15206 10204 15258
rect 10228 15206 10242 15258
rect 10242 15206 10254 15258
rect 10254 15206 10284 15258
rect 10308 15206 10318 15258
rect 10318 15206 10364 15258
rect 10068 15204 10124 15206
rect 10148 15204 10204 15206
rect 10228 15204 10284 15206
rect 10308 15204 10364 15206
rect 10068 14170 10124 14172
rect 10148 14170 10204 14172
rect 10228 14170 10284 14172
rect 10308 14170 10364 14172
rect 10068 14118 10114 14170
rect 10114 14118 10124 14170
rect 10148 14118 10178 14170
rect 10178 14118 10190 14170
rect 10190 14118 10204 14170
rect 10228 14118 10242 14170
rect 10242 14118 10254 14170
rect 10254 14118 10284 14170
rect 10308 14118 10318 14170
rect 10318 14118 10364 14170
rect 10068 14116 10124 14118
rect 10148 14116 10204 14118
rect 10228 14116 10284 14118
rect 10308 14116 10364 14118
rect 10068 13082 10124 13084
rect 10148 13082 10204 13084
rect 10228 13082 10284 13084
rect 10308 13082 10364 13084
rect 10068 13030 10114 13082
rect 10114 13030 10124 13082
rect 10148 13030 10178 13082
rect 10178 13030 10190 13082
rect 10190 13030 10204 13082
rect 10228 13030 10242 13082
rect 10242 13030 10254 13082
rect 10254 13030 10284 13082
rect 10308 13030 10318 13082
rect 10318 13030 10364 13082
rect 10068 13028 10124 13030
rect 10148 13028 10204 13030
rect 10228 13028 10284 13030
rect 10308 13028 10364 13030
rect 10728 16890 10784 16892
rect 10808 16890 10864 16892
rect 10888 16890 10944 16892
rect 10968 16890 11024 16892
rect 10728 16838 10774 16890
rect 10774 16838 10784 16890
rect 10808 16838 10838 16890
rect 10838 16838 10850 16890
rect 10850 16838 10864 16890
rect 10888 16838 10902 16890
rect 10902 16838 10914 16890
rect 10914 16838 10944 16890
rect 10968 16838 10978 16890
rect 10978 16838 11024 16890
rect 10728 16836 10784 16838
rect 10808 16836 10864 16838
rect 10888 16836 10944 16838
rect 10968 16836 11024 16838
rect 10966 16632 11022 16688
rect 10728 15802 10784 15804
rect 10808 15802 10864 15804
rect 10888 15802 10944 15804
rect 10968 15802 11024 15804
rect 10728 15750 10774 15802
rect 10774 15750 10784 15802
rect 10808 15750 10838 15802
rect 10838 15750 10850 15802
rect 10850 15750 10864 15802
rect 10888 15750 10902 15802
rect 10902 15750 10914 15802
rect 10914 15750 10944 15802
rect 10968 15750 10978 15802
rect 10978 15750 11024 15802
rect 10728 15748 10784 15750
rect 10808 15748 10864 15750
rect 10888 15748 10944 15750
rect 10968 15748 11024 15750
rect 12714 29008 12770 29064
rect 12346 23024 12402 23080
rect 12254 18128 12310 18184
rect 11150 14864 11206 14920
rect 11426 14864 11482 14920
rect 10728 14714 10784 14716
rect 10808 14714 10864 14716
rect 10888 14714 10944 14716
rect 10968 14714 11024 14716
rect 10728 14662 10774 14714
rect 10774 14662 10784 14714
rect 10808 14662 10838 14714
rect 10838 14662 10850 14714
rect 10850 14662 10864 14714
rect 10888 14662 10902 14714
rect 10902 14662 10914 14714
rect 10914 14662 10944 14714
rect 10968 14662 10978 14714
rect 10978 14662 11024 14714
rect 10728 14660 10784 14662
rect 10808 14660 10864 14662
rect 10888 14660 10944 14662
rect 10968 14660 11024 14662
rect 10046 12144 10102 12200
rect 10068 11994 10124 11996
rect 10148 11994 10204 11996
rect 10228 11994 10284 11996
rect 10308 11994 10364 11996
rect 10068 11942 10114 11994
rect 10114 11942 10124 11994
rect 10148 11942 10178 11994
rect 10178 11942 10190 11994
rect 10190 11942 10204 11994
rect 10228 11942 10242 11994
rect 10242 11942 10254 11994
rect 10254 11942 10284 11994
rect 10308 11942 10318 11994
rect 10318 11942 10364 11994
rect 10068 11940 10124 11942
rect 10148 11940 10204 11942
rect 10228 11940 10284 11942
rect 10308 11940 10364 11942
rect 9494 8084 9550 8120
rect 9494 8064 9496 8084
rect 9496 8064 9548 8084
rect 9548 8064 9550 8084
rect 9862 10004 9864 10024
rect 9864 10004 9916 10024
rect 9916 10004 9918 10024
rect 9862 9968 9918 10004
rect 10068 10906 10124 10908
rect 10148 10906 10204 10908
rect 10228 10906 10284 10908
rect 10308 10906 10364 10908
rect 10068 10854 10114 10906
rect 10114 10854 10124 10906
rect 10148 10854 10178 10906
rect 10178 10854 10190 10906
rect 10190 10854 10204 10906
rect 10228 10854 10242 10906
rect 10242 10854 10254 10906
rect 10254 10854 10284 10906
rect 10308 10854 10318 10906
rect 10318 10854 10364 10906
rect 10068 10852 10124 10854
rect 10148 10852 10204 10854
rect 10228 10852 10284 10854
rect 10308 10852 10364 10854
rect 10728 13626 10784 13628
rect 10808 13626 10864 13628
rect 10888 13626 10944 13628
rect 10968 13626 11024 13628
rect 10728 13574 10774 13626
rect 10774 13574 10784 13626
rect 10808 13574 10838 13626
rect 10838 13574 10850 13626
rect 10850 13574 10864 13626
rect 10888 13574 10902 13626
rect 10902 13574 10914 13626
rect 10914 13574 10944 13626
rect 10968 13574 10978 13626
rect 10978 13574 11024 13626
rect 10728 13572 10784 13574
rect 10808 13572 10864 13574
rect 10888 13572 10944 13574
rect 10968 13572 11024 13574
rect 10728 12538 10784 12540
rect 10808 12538 10864 12540
rect 10888 12538 10944 12540
rect 10968 12538 11024 12540
rect 10728 12486 10774 12538
rect 10774 12486 10784 12538
rect 10808 12486 10838 12538
rect 10838 12486 10850 12538
rect 10850 12486 10864 12538
rect 10888 12486 10902 12538
rect 10902 12486 10914 12538
rect 10914 12486 10944 12538
rect 10968 12486 10978 12538
rect 10978 12486 11024 12538
rect 10728 12484 10784 12486
rect 10808 12484 10864 12486
rect 10888 12484 10944 12486
rect 10968 12484 11024 12486
rect 11150 12416 11206 12472
rect 10966 12300 11022 12336
rect 10966 12280 10968 12300
rect 10968 12280 11020 12300
rect 11020 12280 11022 12300
rect 10728 11450 10784 11452
rect 10808 11450 10864 11452
rect 10888 11450 10944 11452
rect 10968 11450 11024 11452
rect 10728 11398 10774 11450
rect 10774 11398 10784 11450
rect 10808 11398 10838 11450
rect 10838 11398 10850 11450
rect 10850 11398 10864 11450
rect 10888 11398 10902 11450
rect 10902 11398 10914 11450
rect 10914 11398 10944 11450
rect 10968 11398 10978 11450
rect 10978 11398 11024 11450
rect 10728 11396 10784 11398
rect 10808 11396 10864 11398
rect 10888 11396 10944 11398
rect 10968 11396 11024 11398
rect 10728 10362 10784 10364
rect 10808 10362 10864 10364
rect 10888 10362 10944 10364
rect 10968 10362 11024 10364
rect 10728 10310 10774 10362
rect 10774 10310 10784 10362
rect 10808 10310 10838 10362
rect 10838 10310 10850 10362
rect 10850 10310 10864 10362
rect 10888 10310 10902 10362
rect 10902 10310 10914 10362
rect 10914 10310 10944 10362
rect 10968 10310 10978 10362
rect 10978 10310 11024 10362
rect 10728 10308 10784 10310
rect 10808 10308 10864 10310
rect 10888 10308 10944 10310
rect 10968 10308 11024 10310
rect 10068 9818 10124 9820
rect 10148 9818 10204 9820
rect 10228 9818 10284 9820
rect 10308 9818 10364 9820
rect 10068 9766 10114 9818
rect 10114 9766 10124 9818
rect 10148 9766 10178 9818
rect 10178 9766 10190 9818
rect 10190 9766 10204 9818
rect 10228 9766 10242 9818
rect 10242 9766 10254 9818
rect 10254 9766 10284 9818
rect 10308 9766 10318 9818
rect 10318 9766 10364 9818
rect 10068 9764 10124 9766
rect 10148 9764 10204 9766
rect 10228 9764 10284 9766
rect 10308 9764 10364 9766
rect 9954 9560 10010 9616
rect 10598 9968 10654 10024
rect 10690 9424 10746 9480
rect 9770 7248 9826 7304
rect 9770 6860 9826 6896
rect 9770 6840 9772 6860
rect 9772 6840 9824 6860
rect 9824 6840 9826 6860
rect 9678 6196 9680 6216
rect 9680 6196 9732 6216
rect 9732 6196 9734 6216
rect 9678 6160 9734 6196
rect 10068 8730 10124 8732
rect 10148 8730 10204 8732
rect 10228 8730 10284 8732
rect 10308 8730 10364 8732
rect 10068 8678 10114 8730
rect 10114 8678 10124 8730
rect 10148 8678 10178 8730
rect 10178 8678 10190 8730
rect 10190 8678 10204 8730
rect 10228 8678 10242 8730
rect 10242 8678 10254 8730
rect 10254 8678 10284 8730
rect 10308 8678 10318 8730
rect 10318 8678 10364 8730
rect 10068 8676 10124 8678
rect 10148 8676 10204 8678
rect 10228 8676 10284 8678
rect 10308 8676 10364 8678
rect 10322 8200 10378 8256
rect 10068 7642 10124 7644
rect 10148 7642 10204 7644
rect 10228 7642 10284 7644
rect 10308 7642 10364 7644
rect 10068 7590 10114 7642
rect 10114 7590 10124 7642
rect 10148 7590 10178 7642
rect 10178 7590 10190 7642
rect 10190 7590 10204 7642
rect 10228 7590 10242 7642
rect 10242 7590 10254 7642
rect 10254 7590 10284 7642
rect 10308 7590 10318 7642
rect 10318 7590 10364 7642
rect 10068 7588 10124 7590
rect 10148 7588 10204 7590
rect 10228 7588 10284 7590
rect 10308 7588 10364 7590
rect 10728 9274 10784 9276
rect 10808 9274 10864 9276
rect 10888 9274 10944 9276
rect 10968 9274 11024 9276
rect 10728 9222 10774 9274
rect 10774 9222 10784 9274
rect 10808 9222 10838 9274
rect 10838 9222 10850 9274
rect 10850 9222 10864 9274
rect 10888 9222 10902 9274
rect 10902 9222 10914 9274
rect 10914 9222 10944 9274
rect 10968 9222 10978 9274
rect 10978 9222 11024 9274
rect 10728 9220 10784 9222
rect 10808 9220 10864 9222
rect 10888 9220 10944 9222
rect 10968 9220 11024 9222
rect 11150 9560 11206 9616
rect 10728 8186 10784 8188
rect 10808 8186 10864 8188
rect 10888 8186 10944 8188
rect 10968 8186 11024 8188
rect 10728 8134 10774 8186
rect 10774 8134 10784 8186
rect 10808 8134 10838 8186
rect 10838 8134 10850 8186
rect 10850 8134 10864 8186
rect 10888 8134 10902 8186
rect 10902 8134 10914 8186
rect 10914 8134 10944 8186
rect 10968 8134 10978 8186
rect 10978 8134 11024 8186
rect 10728 8132 10784 8134
rect 10808 8132 10864 8134
rect 10888 8132 10944 8134
rect 10968 8132 11024 8134
rect 10068 6554 10124 6556
rect 10148 6554 10204 6556
rect 10228 6554 10284 6556
rect 10308 6554 10364 6556
rect 10068 6502 10114 6554
rect 10114 6502 10124 6554
rect 10148 6502 10178 6554
rect 10178 6502 10190 6554
rect 10190 6502 10204 6554
rect 10228 6502 10242 6554
rect 10242 6502 10254 6554
rect 10254 6502 10284 6554
rect 10308 6502 10318 6554
rect 10318 6502 10364 6554
rect 10068 6500 10124 6502
rect 10148 6500 10204 6502
rect 10228 6500 10284 6502
rect 10308 6500 10364 6502
rect 10068 5466 10124 5468
rect 10148 5466 10204 5468
rect 10228 5466 10284 5468
rect 10308 5466 10364 5468
rect 10068 5414 10114 5466
rect 10114 5414 10124 5466
rect 10148 5414 10178 5466
rect 10178 5414 10190 5466
rect 10190 5414 10204 5466
rect 10228 5414 10242 5466
rect 10242 5414 10254 5466
rect 10254 5414 10284 5466
rect 10308 5414 10318 5466
rect 10318 5414 10364 5466
rect 10068 5412 10124 5414
rect 10148 5412 10204 5414
rect 10228 5412 10284 5414
rect 10308 5412 10364 5414
rect 10068 4378 10124 4380
rect 10148 4378 10204 4380
rect 10228 4378 10284 4380
rect 10308 4378 10364 4380
rect 10068 4326 10114 4378
rect 10114 4326 10124 4378
rect 10148 4326 10178 4378
rect 10178 4326 10190 4378
rect 10190 4326 10204 4378
rect 10228 4326 10242 4378
rect 10242 4326 10254 4378
rect 10254 4326 10284 4378
rect 10308 4326 10318 4378
rect 10318 4326 10364 4378
rect 10068 4324 10124 4326
rect 10148 4324 10204 4326
rect 10228 4324 10284 4326
rect 10308 4324 10364 4326
rect 10728 7098 10784 7100
rect 10808 7098 10864 7100
rect 10888 7098 10944 7100
rect 10968 7098 11024 7100
rect 10728 7046 10774 7098
rect 10774 7046 10784 7098
rect 10808 7046 10838 7098
rect 10838 7046 10850 7098
rect 10850 7046 10864 7098
rect 10888 7046 10902 7098
rect 10902 7046 10914 7098
rect 10914 7046 10944 7098
rect 10968 7046 10978 7098
rect 10978 7046 11024 7098
rect 10728 7044 10784 7046
rect 10808 7044 10864 7046
rect 10888 7044 10944 7046
rect 10968 7044 11024 7046
rect 11794 15544 11850 15600
rect 11702 13640 11758 13696
rect 10874 6180 10930 6216
rect 10874 6160 10876 6180
rect 10876 6160 10928 6180
rect 10928 6160 10930 6180
rect 10728 6010 10784 6012
rect 10808 6010 10864 6012
rect 10888 6010 10944 6012
rect 10968 6010 11024 6012
rect 10728 5958 10774 6010
rect 10774 5958 10784 6010
rect 10808 5958 10838 6010
rect 10838 5958 10850 6010
rect 10850 5958 10864 6010
rect 10888 5958 10902 6010
rect 10902 5958 10914 6010
rect 10914 5958 10944 6010
rect 10968 5958 10978 6010
rect 10978 5958 11024 6010
rect 10728 5956 10784 5958
rect 10808 5956 10864 5958
rect 10888 5956 10944 5958
rect 10968 5956 11024 5958
rect 10728 4922 10784 4924
rect 10808 4922 10864 4924
rect 10888 4922 10944 4924
rect 10968 4922 11024 4924
rect 10728 4870 10774 4922
rect 10774 4870 10784 4922
rect 10808 4870 10838 4922
rect 10838 4870 10850 4922
rect 10850 4870 10864 4922
rect 10888 4870 10902 4922
rect 10902 4870 10914 4922
rect 10914 4870 10944 4922
rect 10968 4870 10978 4922
rect 10978 4870 11024 4922
rect 10728 4868 10784 4870
rect 10808 4868 10864 4870
rect 10888 4868 10944 4870
rect 10968 4868 11024 4870
rect 10068 3290 10124 3292
rect 10148 3290 10204 3292
rect 10228 3290 10284 3292
rect 10308 3290 10364 3292
rect 10068 3238 10114 3290
rect 10114 3238 10124 3290
rect 10148 3238 10178 3290
rect 10178 3238 10190 3290
rect 10190 3238 10204 3290
rect 10228 3238 10242 3290
rect 10242 3238 10254 3290
rect 10254 3238 10284 3290
rect 10308 3238 10318 3290
rect 10318 3238 10364 3290
rect 10068 3236 10124 3238
rect 10148 3236 10204 3238
rect 10228 3236 10284 3238
rect 10308 3236 10364 3238
rect 10728 3834 10784 3836
rect 10808 3834 10864 3836
rect 10888 3834 10944 3836
rect 10968 3834 11024 3836
rect 10728 3782 10774 3834
rect 10774 3782 10784 3834
rect 10808 3782 10838 3834
rect 10838 3782 10850 3834
rect 10850 3782 10864 3834
rect 10888 3782 10902 3834
rect 10902 3782 10914 3834
rect 10914 3782 10944 3834
rect 10968 3782 10978 3834
rect 10978 3782 11024 3834
rect 10728 3780 10784 3782
rect 10808 3780 10864 3782
rect 10888 3780 10944 3782
rect 10968 3780 11024 3782
rect 10046 2488 10102 2544
rect 10068 2202 10124 2204
rect 10148 2202 10204 2204
rect 10228 2202 10284 2204
rect 10308 2202 10364 2204
rect 10068 2150 10114 2202
rect 10114 2150 10124 2202
rect 10148 2150 10178 2202
rect 10178 2150 10190 2202
rect 10190 2150 10204 2202
rect 10228 2150 10242 2202
rect 10242 2150 10254 2202
rect 10254 2150 10284 2202
rect 10308 2150 10318 2202
rect 10318 2150 10364 2202
rect 10068 2148 10124 2150
rect 10148 2148 10204 2150
rect 10228 2148 10284 2150
rect 10308 2148 10364 2150
rect 10728 2746 10784 2748
rect 10808 2746 10864 2748
rect 10888 2746 10944 2748
rect 10968 2746 11024 2748
rect 10728 2694 10774 2746
rect 10774 2694 10784 2746
rect 10808 2694 10838 2746
rect 10838 2694 10850 2746
rect 10850 2694 10864 2746
rect 10888 2694 10902 2746
rect 10902 2694 10914 2746
rect 10914 2694 10944 2746
rect 10968 2694 10978 2746
rect 10978 2694 11024 2746
rect 10728 2692 10784 2694
rect 10808 2692 10864 2694
rect 10888 2692 10944 2694
rect 10968 2692 11024 2694
rect 12714 23432 12770 23488
rect 10728 1658 10784 1660
rect 10808 1658 10864 1660
rect 10888 1658 10944 1660
rect 10968 1658 11024 1660
rect 10728 1606 10774 1658
rect 10774 1606 10784 1658
rect 10808 1606 10838 1658
rect 10838 1606 10850 1658
rect 10850 1606 10864 1658
rect 10888 1606 10902 1658
rect 10902 1606 10914 1658
rect 10914 1606 10944 1658
rect 10968 1606 10978 1658
rect 10978 1606 11024 1658
rect 10728 1604 10784 1606
rect 10808 1604 10864 1606
rect 10888 1604 10944 1606
rect 10968 1604 11024 1606
rect 10068 1114 10124 1116
rect 10148 1114 10204 1116
rect 10228 1114 10284 1116
rect 10308 1114 10364 1116
rect 10068 1062 10114 1114
rect 10114 1062 10124 1114
rect 10148 1062 10178 1114
rect 10178 1062 10190 1114
rect 10190 1062 10204 1114
rect 10228 1062 10242 1114
rect 10242 1062 10254 1114
rect 10254 1062 10284 1114
rect 10308 1062 10318 1114
rect 10318 1062 10364 1114
rect 10068 1060 10124 1062
rect 10148 1060 10204 1062
rect 10228 1060 10284 1062
rect 10308 1060 10364 1062
rect 4328 570 4384 572
rect 4408 570 4464 572
rect 4488 570 4544 572
rect 4568 570 4624 572
rect 4328 518 4374 570
rect 4374 518 4384 570
rect 4408 518 4438 570
rect 4438 518 4450 570
rect 4450 518 4464 570
rect 4488 518 4502 570
rect 4502 518 4514 570
rect 4514 518 4544 570
rect 4568 518 4578 570
rect 4578 518 4624 570
rect 4328 516 4384 518
rect 4408 516 4464 518
rect 4488 516 4544 518
rect 4568 516 4624 518
rect 10728 570 10784 572
rect 10808 570 10864 572
rect 10888 570 10944 572
rect 10968 570 11024 572
rect 10728 518 10774 570
rect 10774 518 10784 570
rect 10808 518 10838 570
rect 10838 518 10850 570
rect 10850 518 10864 570
rect 10888 518 10902 570
rect 10902 518 10914 570
rect 10914 518 10944 570
rect 10968 518 10978 570
rect 10978 518 11024 570
rect 10728 516 10784 518
rect 10808 516 10864 518
rect 10888 516 10944 518
rect 10968 516 11024 518
<< metal3 >>
rect 1342 43556 1348 43620
rect 1412 43618 1418 43620
rect 2221 43618 2287 43621
rect 1412 43616 2287 43618
rect 1412 43560 2226 43616
rect 2282 43560 2287 43616
rect 1412 43558 2287 43560
rect 1412 43556 1418 43558
rect 2221 43555 2287 43558
rect 4981 43618 5047 43621
rect 5390 43618 5396 43620
rect 4981 43616 5396 43618
rect 4981 43560 4986 43616
rect 5042 43560 5396 43616
rect 4981 43558 5396 43560
rect 4981 43555 5047 43558
rect 5390 43556 5396 43558
rect 5460 43556 5466 43620
rect 5574 43556 5580 43620
rect 5644 43618 5650 43620
rect 6085 43618 6151 43621
rect 5644 43616 6151 43618
rect 5644 43560 6090 43616
rect 6146 43560 6151 43616
rect 5644 43558 6151 43560
rect 5644 43556 5650 43558
rect 6085 43555 6151 43558
rect 7741 43618 7807 43621
rect 8150 43618 8156 43620
rect 7741 43616 8156 43618
rect 7741 43560 7746 43616
rect 7802 43560 8156 43616
rect 7741 43558 8156 43560
rect 7741 43555 7807 43558
rect 8150 43556 8156 43558
rect 8220 43556 8226 43620
rect 8845 43618 8911 43621
rect 9254 43618 9260 43620
rect 8845 43616 9260 43618
rect 8845 43560 8850 43616
rect 8906 43560 9260 43616
rect 8845 43558 9260 43560
rect 8845 43555 8911 43558
rect 9254 43556 9260 43558
rect 9324 43556 9330 43620
rect 9397 43618 9463 43621
rect 9622 43618 9628 43620
rect 9397 43616 9628 43618
rect 9397 43560 9402 43616
rect 9458 43560 9628 43616
rect 9397 43558 9628 43560
rect 9397 43555 9463 43558
rect 9622 43556 9628 43558
rect 9692 43556 9698 43620
rect 4318 43008 4634 43009
rect 4318 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4634 43008
rect 4318 42943 4634 42944
rect 10718 43008 11034 43009
rect 10718 42944 10724 43008
rect 10788 42944 10804 43008
rect 10868 42944 10884 43008
rect 10948 42944 10964 43008
rect 11028 42944 11034 43008
rect 10718 42943 11034 42944
rect 841 42666 907 42669
rect 4245 42666 4311 42669
rect 7465 42666 7531 42669
rect 8293 42666 8359 42669
rect 841 42664 8359 42666
rect 841 42608 846 42664
rect 902 42608 4250 42664
rect 4306 42608 7470 42664
rect 7526 42608 8298 42664
rect 8354 42608 8359 42664
rect 841 42606 8359 42608
rect 841 42603 907 42606
rect 4245 42603 4311 42606
rect 7465 42603 7531 42606
rect 8293 42603 8359 42606
rect 4153 42530 4219 42533
rect 4981 42530 5047 42533
rect 7741 42530 7807 42533
rect 4153 42528 7807 42530
rect 4153 42472 4158 42528
rect 4214 42472 4986 42528
rect 5042 42472 7746 42528
rect 7802 42472 7807 42528
rect 4153 42470 7807 42472
rect 4153 42467 4219 42470
rect 4981 42467 5047 42470
rect 7741 42467 7807 42470
rect 3658 42464 3974 42465
rect 3658 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3974 42464
rect 3658 42399 3974 42400
rect 10058 42464 10374 42465
rect 10058 42400 10064 42464
rect 10128 42400 10144 42464
rect 10208 42400 10224 42464
rect 10288 42400 10304 42464
rect 10368 42400 10374 42464
rect 10058 42399 10374 42400
rect 8702 41924 8708 41988
rect 8772 41986 8778 41988
rect 9121 41986 9187 41989
rect 8772 41984 9187 41986
rect 8772 41928 9126 41984
rect 9182 41928 9187 41984
rect 8772 41926 9187 41928
rect 8772 41924 8778 41926
rect 9121 41923 9187 41926
rect 11462 41924 11468 41988
rect 11532 41986 11538 41988
rect 11881 41986 11947 41989
rect 11532 41984 11947 41986
rect 11532 41928 11886 41984
rect 11942 41928 11947 41984
rect 11532 41926 11947 41928
rect 11532 41924 11538 41926
rect 11881 41923 11947 41926
rect 4318 41920 4634 41921
rect 4318 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4634 41920
rect 4318 41855 4634 41856
rect 10718 41920 11034 41921
rect 10718 41856 10724 41920
rect 10788 41856 10804 41920
rect 10868 41856 10884 41920
rect 10948 41856 10964 41920
rect 11028 41856 11034 41920
rect 10718 41855 11034 41856
rect 0 41716 400 41744
rect 0 41652 382 41716
rect 446 41652 452 41716
rect 2037 41714 2103 41717
rect 6637 41714 6703 41717
rect 2037 41712 6703 41714
rect 2037 41656 2042 41712
rect 2098 41656 6642 41712
rect 6698 41656 6703 41712
rect 2037 41654 6703 41656
rect 0 41624 400 41652
rect 2037 41651 2103 41654
rect 6637 41651 6703 41654
rect 9806 41652 9812 41716
rect 9876 41714 9882 41716
rect 10409 41714 10475 41717
rect 9876 41712 10475 41714
rect 9876 41656 10414 41712
rect 10470 41656 10475 41712
rect 9876 41654 10475 41656
rect 9876 41652 9882 41654
rect 10409 41651 10475 41654
rect 3366 41516 3372 41580
rect 3436 41578 3442 41580
rect 6361 41578 6427 41581
rect 3436 41576 6427 41578
rect 3436 41520 6366 41576
rect 6422 41520 6427 41576
rect 3436 41518 6427 41520
rect 3436 41516 3442 41518
rect 6361 41515 6427 41518
rect 6494 41516 6500 41580
rect 6564 41578 6570 41580
rect 7373 41578 7439 41581
rect 6564 41576 7439 41578
rect 6564 41520 7378 41576
rect 7434 41520 7439 41576
rect 6564 41518 7439 41520
rect 6564 41516 6570 41518
rect 7373 41515 7439 41518
rect 10777 41578 10843 41581
rect 11646 41578 11652 41580
rect 10777 41576 11652 41578
rect 10777 41520 10782 41576
rect 10838 41520 11652 41576
rect 10777 41518 11652 41520
rect 10777 41515 10843 41518
rect 11646 41516 11652 41518
rect 11716 41516 11722 41580
rect 0 41442 400 41472
rect 933 41442 999 41445
rect 0 41440 999 41442
rect 0 41384 938 41440
rect 994 41384 999 41440
rect 0 41382 999 41384
rect 0 41352 400 41382
rect 933 41379 999 41382
rect 6545 41442 6611 41445
rect 7649 41442 7715 41445
rect 6545 41440 7715 41442
rect 6545 41384 6550 41440
rect 6606 41384 7654 41440
rect 7710 41384 7715 41440
rect 6545 41382 7715 41384
rect 6545 41379 6611 41382
rect 7649 41379 7715 41382
rect 3658 41376 3974 41377
rect 3658 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3974 41376
rect 3658 41311 3974 41312
rect 10058 41376 10374 41377
rect 10058 41312 10064 41376
rect 10128 41312 10144 41376
rect 10208 41312 10224 41376
rect 10288 41312 10304 41376
rect 10368 41312 10374 41376
rect 10058 41311 10374 41312
rect 7046 41244 7052 41308
rect 7116 41306 7122 41308
rect 7373 41306 7439 41309
rect 8753 41306 8819 41309
rect 7116 41304 8819 41306
rect 7116 41248 7378 41304
rect 7434 41248 8758 41304
rect 8814 41248 8819 41304
rect 7116 41246 8819 41248
rect 7116 41244 7122 41246
rect 7373 41243 7439 41246
rect 8753 41243 8819 41246
rect 0 41173 400 41200
rect 0 41168 447 41173
rect 0 41112 386 41168
rect 442 41112 447 41168
rect 0 41107 447 41112
rect 2589 41170 2655 41173
rect 9673 41170 9739 41173
rect 2589 41168 9739 41170
rect 2589 41112 2594 41168
rect 2650 41112 9678 41168
rect 9734 41112 9739 41168
rect 2589 41110 9739 41112
rect 2589 41107 2655 41110
rect 9673 41107 9739 41110
rect 0 41080 400 41107
rect 1158 40972 1164 41036
rect 1228 41034 1234 41036
rect 6361 41034 6427 41037
rect 1228 41032 6427 41034
rect 1228 40976 6366 41032
rect 6422 40976 6427 41032
rect 1228 40974 6427 40976
rect 1228 40972 1234 40974
rect 6361 40971 6427 40974
rect 8518 40972 8524 41036
rect 8588 41034 8594 41036
rect 10869 41034 10935 41037
rect 8588 41032 10935 41034
rect 8588 40976 10874 41032
rect 10930 40976 10935 41032
rect 8588 40974 10935 40976
rect 8588 40972 8594 40974
rect 10869 40971 10935 40974
rect 0 40898 400 40928
rect 565 40898 631 40901
rect 0 40896 631 40898
rect 0 40840 570 40896
rect 626 40840 631 40896
rect 0 40838 631 40840
rect 0 40808 400 40838
rect 565 40835 631 40838
rect 5625 40898 5691 40901
rect 9949 40898 10015 40901
rect 5625 40896 10015 40898
rect 5625 40840 5630 40896
rect 5686 40840 9954 40896
rect 10010 40840 10015 40896
rect 5625 40838 10015 40840
rect 5625 40835 5691 40838
rect 9949 40835 10015 40838
rect 4318 40832 4634 40833
rect 4318 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4634 40832
rect 4318 40767 4634 40768
rect 10718 40832 11034 40833
rect 10718 40768 10724 40832
rect 10788 40768 10804 40832
rect 10868 40768 10884 40832
rect 10948 40768 10964 40832
rect 11028 40768 11034 40832
rect 10718 40767 11034 40768
rect 3325 40762 3391 40765
rect 5165 40764 5231 40765
rect 5165 40762 5212 40764
rect 2500 40760 3391 40762
rect 2500 40704 3330 40760
rect 3386 40704 3391 40760
rect 2500 40702 3391 40704
rect 5124 40760 5212 40762
rect 5276 40762 5282 40764
rect 6269 40762 6335 40765
rect 5276 40760 6335 40762
rect 5124 40704 5170 40760
rect 5276 40704 6274 40760
rect 6330 40704 6335 40760
rect 5124 40702 5212 40704
rect 0 40626 400 40656
rect 2500 40629 2560 40702
rect 3325 40699 3391 40702
rect 5165 40700 5212 40702
rect 5276 40702 6335 40704
rect 5276 40700 5282 40702
rect 5165 40699 5231 40700
rect 6269 40699 6335 40702
rect 1209 40626 1275 40629
rect 0 40624 1275 40626
rect 0 40568 1214 40624
rect 1270 40568 1275 40624
rect 0 40566 1275 40568
rect 0 40536 400 40566
rect 1209 40563 1275 40566
rect 2497 40624 2563 40629
rect 2497 40568 2502 40624
rect 2558 40568 2563 40624
rect 2497 40563 2563 40568
rect 2957 40626 3023 40629
rect 5257 40626 5323 40629
rect 8385 40626 8451 40629
rect 2957 40624 5323 40626
rect 2957 40568 2962 40624
rect 3018 40568 5262 40624
rect 5318 40568 5323 40624
rect 2957 40566 5323 40568
rect 2957 40563 3023 40566
rect 5257 40563 5323 40566
rect 7238 40624 8451 40626
rect 7238 40568 8390 40624
rect 8446 40568 8451 40624
rect 7238 40566 8451 40568
rect 841 40490 907 40493
rect 7238 40490 7298 40566
rect 8385 40563 8451 40566
rect 7465 40492 7531 40493
rect 841 40488 7298 40490
rect 841 40432 846 40488
rect 902 40432 7298 40488
rect 841 40430 7298 40432
rect 841 40427 907 40430
rect 7414 40428 7420 40492
rect 7484 40490 7531 40492
rect 7484 40488 7576 40490
rect 7526 40432 7576 40488
rect 7484 40430 7576 40432
rect 7484 40428 7531 40430
rect 7465 40427 7531 40428
rect 0 40354 400 40384
rect 3509 40354 3575 40357
rect 0 40352 3575 40354
rect 0 40296 3514 40352
rect 3570 40296 3575 40352
rect 0 40294 3575 40296
rect 0 40264 400 40294
rect 3509 40291 3575 40294
rect 6913 40354 6979 40357
rect 8201 40354 8267 40357
rect 6913 40352 8267 40354
rect 6913 40296 6918 40352
rect 6974 40296 8206 40352
rect 8262 40296 8267 40352
rect 6913 40294 8267 40296
rect 6913 40291 6979 40294
rect 8201 40291 8267 40294
rect 3658 40288 3974 40289
rect 3658 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3974 40288
rect 3658 40223 3974 40224
rect 10058 40288 10374 40289
rect 10058 40224 10064 40288
rect 10128 40224 10144 40288
rect 10208 40224 10224 40288
rect 10288 40224 10304 40288
rect 10368 40224 10374 40288
rect 10058 40223 10374 40224
rect 3049 40218 3115 40221
rect 3182 40218 3188 40220
rect 3049 40216 3188 40218
rect 3049 40160 3054 40216
rect 3110 40160 3188 40216
rect 3049 40158 3188 40160
rect 3049 40155 3115 40158
rect 3182 40156 3188 40158
rect 3252 40156 3258 40220
rect 5942 40156 5948 40220
rect 6012 40218 6018 40220
rect 9305 40218 9371 40221
rect 6012 40216 9371 40218
rect 6012 40160 9310 40216
rect 9366 40160 9371 40216
rect 6012 40158 9371 40160
rect 6012 40156 6018 40158
rect 9305 40155 9371 40158
rect 10542 40156 10548 40220
rect 10612 40218 10618 40220
rect 10685 40218 10751 40221
rect 10612 40216 10751 40218
rect 10612 40160 10690 40216
rect 10746 40160 10751 40216
rect 10612 40158 10751 40160
rect 10612 40156 10618 40158
rect 10685 40155 10751 40158
rect 0 40082 400 40112
rect 1393 40082 1459 40085
rect 0 40080 1459 40082
rect 0 40024 1398 40080
rect 1454 40024 1459 40080
rect 0 40022 1459 40024
rect 0 39992 400 40022
rect 1393 40019 1459 40022
rect 2497 40082 2563 40085
rect 2865 40082 2931 40085
rect 2497 40080 2931 40082
rect 2497 40024 2502 40080
rect 2558 40024 2870 40080
rect 2926 40024 2931 40080
rect 2497 40022 2931 40024
rect 2497 40019 2563 40022
rect 2865 40019 2931 40022
rect 3417 40082 3483 40085
rect 4102 40082 4108 40084
rect 3417 40080 4108 40082
rect 3417 40024 3422 40080
rect 3478 40024 4108 40080
rect 3417 40022 4108 40024
rect 3417 40019 3483 40022
rect 4102 40020 4108 40022
rect 4172 40020 4178 40084
rect 5625 40082 5691 40085
rect 5758 40082 5764 40084
rect 5625 40080 5764 40082
rect 5625 40024 5630 40080
rect 5686 40024 5764 40080
rect 5625 40022 5764 40024
rect 5625 40019 5691 40022
rect 5758 40020 5764 40022
rect 5828 40020 5834 40084
rect 6729 40082 6795 40085
rect 7833 40082 7899 40085
rect 6729 40080 7899 40082
rect 6729 40024 6734 40080
rect 6790 40024 7838 40080
rect 7894 40024 7899 40080
rect 6729 40022 7899 40024
rect 6729 40019 6795 40022
rect 7833 40019 7899 40022
rect 8886 40020 8892 40084
rect 8956 40082 8962 40084
rect 11145 40082 11211 40085
rect 8956 40080 11211 40082
rect 8956 40024 11150 40080
rect 11206 40024 11211 40080
rect 8956 40022 11211 40024
rect 8956 40020 8962 40022
rect 11145 40019 11211 40022
rect 11278 40020 11284 40084
rect 11348 40082 11354 40084
rect 11421 40082 11487 40085
rect 11348 40080 11487 40082
rect 11348 40024 11426 40080
rect 11482 40024 11487 40080
rect 11348 40022 11487 40024
rect 11348 40020 11354 40022
rect 11421 40019 11487 40022
rect 473 39946 539 39949
rect 2078 39946 2084 39948
rect 473 39944 2084 39946
rect 473 39888 478 39944
rect 534 39888 2084 39944
rect 473 39886 2084 39888
rect 473 39883 539 39886
rect 2078 39884 2084 39886
rect 2148 39946 2154 39948
rect 2773 39946 2839 39949
rect 2148 39944 2839 39946
rect 2148 39888 2778 39944
rect 2834 39888 2839 39944
rect 2148 39886 2839 39888
rect 2148 39884 2154 39886
rect 2773 39883 2839 39886
rect 5390 39884 5396 39948
rect 5460 39946 5466 39948
rect 10133 39946 10199 39949
rect 10869 39946 10935 39949
rect 5460 39944 10199 39946
rect 5460 39888 10138 39944
rect 10194 39888 10199 39944
rect 5460 39886 10199 39888
rect 5460 39884 5466 39886
rect 10133 39883 10199 39886
rect 10366 39944 10935 39946
rect 10366 39888 10874 39944
rect 10930 39888 10935 39944
rect 10366 39886 10935 39888
rect 0 39810 400 39840
rect 7281 39810 7347 39813
rect 9397 39810 9463 39813
rect 0 39750 2790 39810
rect 0 39720 400 39750
rect 1117 39674 1183 39677
rect 2037 39674 2103 39677
rect 1117 39672 2103 39674
rect 1117 39616 1122 39672
rect 1178 39616 2042 39672
rect 2098 39616 2103 39672
rect 1117 39614 2103 39616
rect 2730 39674 2790 39750
rect 7281 39808 9463 39810
rect 7281 39752 7286 39808
rect 7342 39752 9402 39808
rect 9458 39752 9463 39808
rect 7281 39750 9463 39752
rect 7281 39747 7347 39750
rect 9397 39747 9463 39750
rect 4318 39744 4634 39745
rect 4318 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4634 39744
rect 4318 39679 4634 39680
rect 6269 39674 6335 39677
rect 9949 39674 10015 39677
rect 10366 39674 10426 39886
rect 10869 39883 10935 39886
rect 10718 39744 11034 39745
rect 10718 39680 10724 39744
rect 10788 39680 10804 39744
rect 10868 39680 10884 39744
rect 10948 39680 10964 39744
rect 11028 39680 11034 39744
rect 10718 39679 11034 39680
rect 2730 39614 4216 39674
rect 1117 39611 1183 39614
rect 2037 39611 2103 39614
rect 0 39538 400 39568
rect 933 39538 999 39541
rect 3049 39538 3115 39541
rect 0 39536 999 39538
rect 0 39480 938 39536
rect 994 39480 999 39536
rect 0 39478 999 39480
rect 0 39448 400 39478
rect 933 39475 999 39478
rect 1166 39536 3115 39538
rect 1166 39480 3054 39536
rect 3110 39480 3115 39536
rect 1166 39478 3115 39480
rect 4156 39538 4216 39614
rect 6269 39672 10426 39674
rect 6269 39616 6274 39672
rect 6330 39616 9954 39672
rect 10010 39616 10426 39672
rect 6269 39614 10426 39616
rect 6269 39611 6335 39614
rect 9949 39611 10015 39614
rect 7373 39538 7439 39541
rect 4156 39536 7439 39538
rect 4156 39480 7378 39536
rect 7434 39480 7439 39536
rect 4156 39478 7439 39480
rect 749 39402 815 39405
rect 1166 39402 1226 39478
rect 3049 39475 3115 39478
rect 7373 39475 7439 39478
rect 7649 39538 7715 39541
rect 7782 39538 7788 39540
rect 7649 39536 7788 39538
rect 7649 39480 7654 39536
rect 7710 39480 7788 39536
rect 7649 39478 7788 39480
rect 7649 39475 7715 39478
rect 7782 39476 7788 39478
rect 7852 39538 7858 39540
rect 10685 39538 10751 39541
rect 11881 39538 11947 39541
rect 7852 39536 11947 39538
rect 7852 39480 10690 39536
rect 10746 39480 11886 39536
rect 11942 39480 11947 39536
rect 7852 39478 11947 39480
rect 7852 39476 7858 39478
rect 10685 39475 10751 39478
rect 11881 39475 11947 39478
rect 749 39400 1226 39402
rect 749 39344 754 39400
rect 810 39344 1226 39400
rect 749 39342 1226 39344
rect 1945 39402 2011 39405
rect 1945 39400 4170 39402
rect 1945 39344 1950 39400
rect 2006 39344 4170 39400
rect 1945 39342 4170 39344
rect 749 39339 815 39342
rect 1945 39339 2011 39342
rect 0 39266 400 39296
rect 933 39266 999 39269
rect 2313 39266 2379 39269
rect 0 39264 999 39266
rect 0 39208 938 39264
rect 994 39208 999 39264
rect 0 39206 999 39208
rect 0 39176 400 39206
rect 933 39203 999 39206
rect 1212 39264 2379 39266
rect 1212 39208 2318 39264
rect 2374 39208 2379 39264
rect 1212 39206 2379 39208
rect 4110 39266 4170 39342
rect 4838 39340 4844 39404
rect 4908 39402 4914 39404
rect 10041 39402 10107 39405
rect 4908 39400 10107 39402
rect 4908 39344 10046 39400
rect 10102 39344 10107 39400
rect 4908 39342 10107 39344
rect 4908 39340 4914 39342
rect 10041 39339 10107 39342
rect 5206 39266 5212 39268
rect 4110 39206 5212 39266
rect 933 39130 999 39133
rect 1212 39130 1272 39206
rect 2313 39203 2379 39206
rect 5206 39204 5212 39206
rect 5276 39204 5282 39268
rect 8109 39266 8175 39269
rect 8661 39266 8727 39269
rect 8109 39264 8727 39266
rect 8109 39208 8114 39264
rect 8170 39208 8666 39264
rect 8722 39208 8727 39264
rect 8109 39206 8727 39208
rect 8109 39203 8175 39206
rect 8661 39203 8727 39206
rect 3658 39200 3974 39201
rect 3658 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3974 39200
rect 3658 39135 3974 39136
rect 10058 39200 10374 39201
rect 10058 39136 10064 39200
rect 10128 39136 10144 39200
rect 10208 39136 10224 39200
rect 10288 39136 10304 39200
rect 10368 39136 10374 39200
rect 10058 39135 10374 39136
rect 933 39128 1272 39130
rect 933 39072 938 39128
rect 994 39072 1272 39128
rect 933 39070 1272 39072
rect 4981 39130 5047 39133
rect 6453 39130 6519 39133
rect 4981 39128 6519 39130
rect 4981 39072 4986 39128
rect 5042 39072 6458 39128
rect 6514 39072 6519 39128
rect 4981 39070 6519 39072
rect 933 39067 999 39070
rect 4981 39067 5047 39070
rect 6453 39067 6519 39070
rect 1209 38994 1275 38997
rect 3877 38994 3943 38997
rect 6545 38994 6611 38997
rect 1209 38992 2790 38994
rect 1209 38936 1214 38992
rect 1270 38936 2790 38992
rect 1209 38934 2790 38936
rect 1209 38931 1275 38934
rect 1393 38858 1459 38861
rect 1526 38858 1532 38860
rect 1393 38856 1532 38858
rect 1393 38800 1398 38856
rect 1454 38800 1532 38856
rect 1393 38798 1532 38800
rect 1393 38795 1459 38798
rect 1526 38796 1532 38798
rect 1596 38858 1602 38860
rect 1853 38858 1919 38861
rect 1596 38856 1919 38858
rect 1596 38800 1858 38856
rect 1914 38800 1919 38856
rect 1596 38798 1919 38800
rect 2730 38858 2790 38934
rect 3877 38992 6611 38994
rect 3877 38936 3882 38992
rect 3938 38936 6550 38992
rect 6606 38936 6611 38992
rect 3877 38934 6611 38936
rect 3877 38931 3943 38934
rect 6545 38931 6611 38934
rect 7465 38994 7531 38997
rect 8201 38994 8267 38997
rect 7465 38992 8267 38994
rect 7465 38936 7470 38992
rect 7526 38936 8206 38992
rect 8262 38936 8267 38992
rect 7465 38934 8267 38936
rect 7465 38931 7531 38934
rect 8201 38931 8267 38934
rect 10225 38994 10291 38997
rect 11237 38994 11303 38997
rect 10225 38992 11303 38994
rect 10225 38936 10230 38992
rect 10286 38936 11242 38992
rect 11298 38936 11303 38992
rect 10225 38934 11303 38936
rect 10225 38931 10291 38934
rect 11237 38931 11303 38934
rect 7097 38858 7163 38861
rect 2730 38856 7163 38858
rect 2730 38800 7102 38856
rect 7158 38800 7163 38856
rect 2730 38798 7163 38800
rect 1596 38796 1602 38798
rect 1853 38795 1919 38798
rect 7097 38795 7163 38798
rect 7230 38796 7236 38860
rect 7300 38858 7306 38860
rect 9806 38858 9812 38860
rect 7300 38798 9812 38858
rect 7300 38796 7306 38798
rect 9806 38796 9812 38798
rect 9876 38796 9882 38860
rect 10133 38858 10199 38861
rect 10409 38858 10475 38861
rect 12014 38858 12020 38860
rect 10133 38856 12020 38858
rect 10133 38800 10138 38856
rect 10194 38800 10414 38856
rect 10470 38800 12020 38856
rect 10133 38798 12020 38800
rect 10133 38795 10199 38798
rect 10409 38795 10475 38798
rect 12014 38796 12020 38798
rect 12084 38796 12090 38860
rect 9213 38722 9279 38725
rect 6870 38720 9279 38722
rect 6870 38664 9218 38720
rect 9274 38664 9279 38720
rect 6870 38662 9279 38664
rect 4318 38656 4634 38657
rect 4318 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4634 38656
rect 4318 38591 4634 38592
rect 381 38586 447 38589
rect 1710 38586 1716 38588
rect 381 38584 1716 38586
rect 381 38528 386 38584
rect 442 38528 1716 38584
rect 381 38526 1716 38528
rect 381 38523 447 38526
rect 1710 38524 1716 38526
rect 1780 38524 1786 38588
rect 5257 38586 5323 38589
rect 6870 38588 6930 38662
rect 9213 38659 9279 38662
rect 9438 38660 9444 38724
rect 9508 38722 9514 38724
rect 9765 38722 9831 38725
rect 9508 38720 9831 38722
rect 9508 38664 9770 38720
rect 9826 38664 9831 38720
rect 9508 38662 9831 38664
rect 9508 38660 9514 38662
rect 9765 38659 9831 38662
rect 10718 38656 11034 38657
rect 10718 38592 10724 38656
rect 10788 38592 10804 38656
rect 10868 38592 10884 38656
rect 10948 38592 10964 38656
rect 11028 38592 11034 38656
rect 10718 38591 11034 38592
rect 5257 38584 5550 38586
rect 5257 38528 5262 38584
rect 5318 38528 5550 38584
rect 5257 38526 5550 38528
rect 5257 38523 5323 38526
rect 5490 38450 5550 38526
rect 6862 38524 6868 38588
rect 6932 38524 6938 38588
rect 5901 38450 5967 38453
rect 7598 38450 7604 38452
rect 5490 38448 7604 38450
rect 5490 38392 5906 38448
rect 5962 38392 7604 38448
rect 5490 38390 7604 38392
rect 5901 38387 5967 38390
rect 7598 38388 7604 38390
rect 7668 38388 7674 38452
rect 9029 38450 9095 38453
rect 9397 38450 9463 38453
rect 9029 38448 9463 38450
rect 9029 38392 9034 38448
rect 9090 38392 9402 38448
rect 9458 38392 9463 38448
rect 9029 38390 9463 38392
rect 9029 38387 9095 38390
rect 9397 38387 9463 38390
rect 9673 38450 9739 38453
rect 10961 38450 11027 38453
rect 9673 38448 11027 38450
rect 9673 38392 9678 38448
rect 9734 38392 10966 38448
rect 11022 38392 11027 38448
rect 9673 38390 11027 38392
rect 9673 38387 9739 38390
rect 10961 38387 11027 38390
rect 3693 38314 3759 38317
rect 3693 38312 5550 38314
rect 3693 38256 3698 38312
rect 3754 38256 5550 38312
rect 3693 38254 5550 38256
rect 3693 38251 3759 38254
rect 1894 38116 1900 38180
rect 1964 38178 1970 38180
rect 2037 38178 2103 38181
rect 1964 38176 2103 38178
rect 1964 38120 2042 38176
rect 2098 38120 2103 38176
rect 1964 38118 2103 38120
rect 5490 38178 5550 38254
rect 6310 38252 6316 38316
rect 6380 38314 6386 38316
rect 8477 38314 8543 38317
rect 6380 38312 8543 38314
rect 6380 38256 8482 38312
rect 8538 38256 8543 38312
rect 6380 38254 8543 38256
rect 6380 38252 6386 38254
rect 8477 38251 8543 38254
rect 8661 38314 8727 38317
rect 9397 38314 9463 38317
rect 8661 38312 9463 38314
rect 8661 38256 8666 38312
rect 8722 38256 9402 38312
rect 9458 38256 9463 38312
rect 8661 38254 9463 38256
rect 8661 38251 8727 38254
rect 9397 38251 9463 38254
rect 9765 38314 9831 38317
rect 10542 38314 10548 38316
rect 9765 38312 10548 38314
rect 9765 38256 9770 38312
rect 9826 38256 10548 38312
rect 9765 38254 10548 38256
rect 9765 38251 9831 38254
rect 10504 38252 10548 38254
rect 10612 38314 10618 38316
rect 10612 38254 10694 38314
rect 10612 38252 10618 38254
rect 11094 38252 11100 38316
rect 11164 38314 11170 38316
rect 11421 38314 11487 38317
rect 11164 38312 11487 38314
rect 11164 38256 11426 38312
rect 11482 38256 11487 38312
rect 11164 38254 11487 38256
rect 11164 38252 11170 38254
rect 8661 38178 8727 38181
rect 9768 38178 9828 38251
rect 5490 38176 9828 38178
rect 5490 38120 8666 38176
rect 8722 38120 9828 38176
rect 5490 38118 9828 38120
rect 10504 38178 10564 38252
rect 11421 38251 11487 38254
rect 11237 38178 11303 38181
rect 11421 38178 11487 38181
rect 10504 38176 11487 38178
rect 10504 38120 11242 38176
rect 11298 38120 11426 38176
rect 11482 38120 11487 38176
rect 10504 38118 11487 38120
rect 1964 38116 1970 38118
rect 2037 38115 2103 38118
rect 8661 38115 8727 38118
rect 11237 38115 11303 38118
rect 11421 38115 11487 38118
rect 3658 38112 3974 38113
rect 3658 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3974 38112
rect 3658 38047 3974 38048
rect 10058 38112 10374 38113
rect 10058 38048 10064 38112
rect 10128 38048 10144 38112
rect 10208 38048 10224 38112
rect 10288 38048 10304 38112
rect 10368 38048 10374 38112
rect 10058 38047 10374 38048
rect 5441 38042 5507 38045
rect 7189 38042 7255 38045
rect 9397 38042 9463 38045
rect 5441 38040 7114 38042
rect 5441 37984 5446 38040
rect 5502 37984 7114 38040
rect 5441 37982 7114 37984
rect 5441 37979 5507 37982
rect 1025 37906 1091 37909
rect 6862 37906 6868 37908
rect 1025 37904 6868 37906
rect 1025 37848 1030 37904
rect 1086 37848 6868 37904
rect 1025 37846 6868 37848
rect 1025 37843 1091 37846
rect 6862 37844 6868 37846
rect 6932 37844 6938 37908
rect 7054 37906 7114 37982
rect 7189 38040 9463 38042
rect 7189 37984 7194 38040
rect 7250 37984 9402 38040
rect 9458 37984 9463 38040
rect 7189 37982 9463 37984
rect 7189 37979 7255 37982
rect 9397 37979 9463 37982
rect 9581 38040 9647 38045
rect 9581 37984 9586 38040
rect 9642 37984 9647 38040
rect 9581 37979 9647 37984
rect 8334 37906 8340 37908
rect 7054 37846 8340 37906
rect 8334 37844 8340 37846
rect 8404 37906 8410 37908
rect 9584 37906 9644 37979
rect 8404 37846 9644 37906
rect 8404 37844 8410 37846
rect 9806 37844 9812 37908
rect 9876 37906 9882 37908
rect 10593 37906 10659 37909
rect 9876 37904 10659 37906
rect 9876 37848 10598 37904
rect 10654 37848 10659 37904
rect 9876 37846 10659 37848
rect 9876 37844 9882 37846
rect 10593 37843 10659 37846
rect 1761 37770 1827 37773
rect 2262 37770 2268 37772
rect 1761 37768 2268 37770
rect 1761 37712 1766 37768
rect 1822 37712 2268 37768
rect 1761 37710 2268 37712
rect 1761 37707 1827 37710
rect 2262 37708 2268 37710
rect 2332 37770 2338 37772
rect 2865 37770 2931 37773
rect 2332 37768 2931 37770
rect 2332 37712 2870 37768
rect 2926 37712 2931 37768
rect 2332 37710 2931 37712
rect 2332 37708 2338 37710
rect 2865 37707 2931 37710
rect 3417 37770 3483 37773
rect 3969 37770 4035 37773
rect 5349 37770 5415 37773
rect 3417 37768 4035 37770
rect 3417 37712 3422 37768
rect 3478 37712 3974 37768
rect 4030 37712 4035 37768
rect 3417 37710 4035 37712
rect 3417 37707 3483 37710
rect 3969 37707 4035 37710
rect 4110 37768 5415 37770
rect 4110 37712 5354 37768
rect 5410 37712 5415 37768
rect 4110 37710 5415 37712
rect 974 37572 980 37636
rect 1044 37634 1050 37636
rect 1117 37634 1183 37637
rect 3601 37634 3667 37637
rect 1044 37632 3667 37634
rect 1044 37576 1122 37632
rect 1178 37576 3606 37632
rect 3662 37576 3667 37632
rect 1044 37574 3667 37576
rect 1044 37572 1050 37574
rect 1117 37571 1183 37574
rect 3601 37571 3667 37574
rect 3785 37634 3851 37637
rect 4110 37634 4170 37710
rect 5349 37707 5415 37710
rect 7005 37770 7071 37773
rect 8845 37770 8911 37773
rect 7005 37768 8911 37770
rect 7005 37712 7010 37768
rect 7066 37712 8850 37768
rect 8906 37712 8911 37768
rect 7005 37710 8911 37712
rect 7005 37707 7071 37710
rect 8845 37707 8911 37710
rect 9213 37770 9279 37773
rect 12341 37770 12407 37773
rect 9213 37768 12407 37770
rect 9213 37712 9218 37768
rect 9274 37712 12346 37768
rect 12402 37712 12407 37768
rect 9213 37710 12407 37712
rect 9213 37707 9279 37710
rect 12341 37707 12407 37710
rect 3785 37632 4170 37634
rect 3785 37576 3790 37632
rect 3846 37576 4170 37632
rect 3785 37574 4170 37576
rect 4797 37634 4863 37637
rect 5533 37634 5599 37637
rect 4797 37632 5599 37634
rect 4797 37576 4802 37632
rect 4858 37576 5538 37632
rect 5594 37576 5599 37632
rect 4797 37574 5599 37576
rect 3785 37571 3851 37574
rect 4797 37571 4863 37574
rect 5533 37571 5599 37574
rect 8017 37634 8083 37637
rect 9070 37634 9076 37636
rect 8017 37632 9076 37634
rect 8017 37576 8022 37632
rect 8078 37576 9076 37632
rect 8017 37574 9076 37576
rect 8017 37571 8083 37574
rect 9070 37572 9076 37574
rect 9140 37572 9146 37636
rect 11145 37634 11211 37637
rect 11145 37632 11346 37634
rect 11145 37576 11150 37632
rect 11206 37576 11346 37632
rect 11145 37574 11346 37576
rect 11145 37571 11211 37574
rect 4318 37568 4634 37569
rect 4318 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4634 37568
rect 4318 37503 4634 37504
rect 10718 37568 11034 37569
rect 10718 37504 10724 37568
rect 10788 37504 10804 37568
rect 10868 37504 10884 37568
rect 10948 37504 10964 37568
rect 11028 37504 11034 37568
rect 10718 37503 11034 37504
rect 1485 37498 1551 37501
rect 2129 37498 2195 37501
rect 3785 37498 3851 37501
rect 5165 37500 5231 37501
rect 5165 37498 5212 37500
rect 1485 37496 3851 37498
rect 1485 37440 1490 37496
rect 1546 37440 2134 37496
rect 2190 37440 3790 37496
rect 3846 37440 3851 37496
rect 1485 37438 3851 37440
rect 5120 37496 5212 37498
rect 5120 37440 5170 37496
rect 5120 37438 5212 37440
rect 1485 37435 1551 37438
rect 2129 37435 2195 37438
rect 3785 37435 3851 37438
rect 5165 37436 5212 37438
rect 5276 37436 5282 37500
rect 5165 37435 5231 37436
rect 2630 37300 2636 37364
rect 2700 37362 2706 37364
rect 3509 37362 3575 37365
rect 2700 37360 3575 37362
rect 2700 37304 3514 37360
rect 3570 37304 3575 37360
rect 2700 37302 3575 37304
rect 2700 37300 2706 37302
rect 3509 37299 3575 37302
rect 4102 37300 4108 37364
rect 4172 37362 4178 37364
rect 4429 37362 4495 37365
rect 4172 37360 4495 37362
rect 4172 37304 4434 37360
rect 4490 37304 4495 37360
rect 4172 37302 4495 37304
rect 4172 37300 4178 37302
rect 4429 37299 4495 37302
rect 5165 37362 5231 37365
rect 5574 37362 5580 37364
rect 5165 37360 5580 37362
rect 5165 37304 5170 37360
rect 5226 37304 5580 37360
rect 5165 37302 5580 37304
rect 5165 37299 5231 37302
rect 5574 37300 5580 37302
rect 5644 37300 5650 37364
rect 7966 37300 7972 37364
rect 8036 37362 8042 37364
rect 8385 37362 8451 37365
rect 8036 37360 8451 37362
rect 8036 37304 8390 37360
rect 8446 37304 8451 37360
rect 8036 37302 8451 37304
rect 8036 37300 8042 37302
rect 8385 37299 8451 37302
rect 10542 37300 10548 37364
rect 10612 37362 10618 37364
rect 11145 37362 11211 37365
rect 10612 37360 11211 37362
rect 10612 37304 11150 37360
rect 11206 37304 11211 37360
rect 10612 37302 11211 37304
rect 10612 37300 10618 37302
rect 11145 37299 11211 37302
rect 11286 37229 11346 37574
rect 11830 37300 11836 37364
rect 11900 37362 11906 37364
rect 11973 37362 12039 37365
rect 11900 37360 12039 37362
rect 11900 37304 11978 37360
rect 12034 37304 12039 37360
rect 11900 37302 12039 37304
rect 11900 37300 11906 37302
rect 11973 37299 12039 37302
rect 1945 37226 2011 37229
rect 4337 37226 4403 37229
rect 1945 37224 4403 37226
rect 1945 37168 1950 37224
rect 2006 37168 4342 37224
rect 4398 37168 4403 37224
rect 1945 37166 4403 37168
rect 1945 37163 2011 37166
rect 4337 37163 4403 37166
rect 8477 37226 8543 37229
rect 9806 37226 9812 37228
rect 8477 37224 9812 37226
rect 8477 37168 8482 37224
rect 8538 37168 9812 37224
rect 8477 37166 9812 37168
rect 8477 37163 8543 37166
rect 9806 37164 9812 37166
rect 9876 37164 9882 37228
rect 11237 37224 11346 37229
rect 11237 37168 11242 37224
rect 11298 37168 11346 37224
rect 11237 37166 11346 37168
rect 11881 37226 11947 37229
rect 12198 37226 12204 37228
rect 11881 37224 12204 37226
rect 11881 37168 11886 37224
rect 11942 37168 12204 37224
rect 11881 37166 12204 37168
rect 11237 37163 11303 37166
rect 11881 37163 11947 37166
rect 12198 37164 12204 37166
rect 12268 37164 12274 37228
rect 0 37090 400 37120
rect 1485 37090 1551 37093
rect 0 37088 1551 37090
rect 0 37032 1490 37088
rect 1546 37032 1551 37088
rect 0 37030 1551 37032
rect 0 37000 400 37030
rect 1485 37027 1551 37030
rect 1761 37090 1827 37093
rect 1894 37090 1900 37092
rect 1761 37088 1900 37090
rect 1761 37032 1766 37088
rect 1822 37032 1900 37088
rect 1761 37030 1900 37032
rect 1761 37027 1827 37030
rect 1894 37028 1900 37030
rect 1964 37028 1970 37092
rect 7598 37028 7604 37092
rect 7668 37090 7674 37092
rect 8753 37090 8819 37093
rect 7668 37088 8819 37090
rect 7668 37032 8758 37088
rect 8814 37032 8819 37088
rect 7668 37030 8819 37032
rect 7668 37028 7674 37030
rect 8753 37027 8819 37030
rect 8937 37090 9003 37093
rect 8937 37088 9276 37090
rect 8937 37032 8942 37088
rect 8998 37032 9276 37088
rect 8937 37030 9276 37032
rect 8937 37027 9003 37030
rect 3658 37024 3974 37025
rect 3658 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3974 37024
rect 3658 36959 3974 36960
rect 1117 36954 1183 36957
rect 1342 36954 1348 36956
rect 1117 36952 1348 36954
rect 1117 36896 1122 36952
rect 1178 36896 1348 36952
rect 1117 36894 1348 36896
rect 1117 36891 1183 36894
rect 1342 36892 1348 36894
rect 1412 36892 1418 36956
rect 7465 36954 7531 36957
rect 8109 36954 8175 36957
rect 8753 36954 8819 36957
rect 4846 36952 8034 36954
rect 4846 36896 7470 36952
rect 7526 36896 8034 36952
rect 4846 36894 8034 36896
rect 0 36818 400 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 400 36758
rect 933 36755 999 36758
rect 1209 36818 1275 36821
rect 4846 36818 4906 36894
rect 7465 36891 7531 36894
rect 1209 36816 4906 36818
rect 1209 36760 1214 36816
rect 1270 36760 4906 36816
rect 1209 36758 4906 36760
rect 4981 36820 5047 36821
rect 4981 36816 5028 36820
rect 5092 36818 5098 36820
rect 7974 36818 8034 36894
rect 8109 36952 8819 36954
rect 8109 36896 8114 36952
rect 8170 36896 8758 36952
rect 8814 36896 8819 36952
rect 8109 36894 8819 36896
rect 8109 36891 8175 36894
rect 8753 36891 8819 36894
rect 9216 36821 9276 37030
rect 10058 37024 10374 37025
rect 10058 36960 10064 37024
rect 10128 36960 10144 37024
rect 10208 36960 10224 37024
rect 10288 36960 10304 37024
rect 10368 36960 10374 37024
rect 10058 36959 10374 36960
rect 11094 36892 11100 36956
rect 11164 36954 11170 36956
rect 11421 36954 11487 36957
rect 11164 36952 11487 36954
rect 11164 36896 11426 36952
rect 11482 36896 11487 36952
rect 11164 36894 11487 36896
rect 11164 36892 11170 36894
rect 11421 36891 11487 36894
rect 8109 36818 8175 36821
rect 4981 36760 4986 36816
rect 1209 36755 1275 36758
rect 4981 36756 5028 36760
rect 5092 36758 5138 36818
rect 7974 36816 8175 36818
rect 7974 36760 8114 36816
rect 8170 36760 8175 36816
rect 7974 36758 8175 36760
rect 5092 36756 5098 36758
rect 4981 36755 5047 36756
rect 8109 36755 8175 36758
rect 9213 36816 9279 36821
rect 9213 36760 9218 36816
rect 9274 36760 9279 36816
rect 9213 36755 9279 36760
rect 10317 36818 10383 36821
rect 11145 36820 11211 36821
rect 11094 36818 11100 36820
rect 10317 36816 11100 36818
rect 11164 36818 11211 36820
rect 11164 36816 11292 36818
rect 10317 36760 10322 36816
rect 10378 36760 11100 36816
rect 11206 36760 11292 36816
rect 10317 36758 11100 36760
rect 10317 36755 10383 36758
rect 11094 36756 11100 36758
rect 11164 36758 11292 36760
rect 11164 36756 11211 36758
rect 11145 36755 11211 36756
rect 2497 36682 2563 36685
rect 7281 36682 7347 36685
rect 2497 36680 7347 36682
rect 2497 36624 2502 36680
rect 2558 36624 7286 36680
rect 7342 36624 7347 36680
rect 2497 36622 7347 36624
rect 2497 36619 2563 36622
rect 7281 36619 7347 36622
rect 8937 36682 9003 36685
rect 10133 36682 10199 36685
rect 10685 36682 10751 36685
rect 8937 36680 10199 36682
rect 8937 36624 8942 36680
rect 8998 36624 10138 36680
rect 10194 36624 10199 36680
rect 8937 36622 10199 36624
rect 8937 36619 9003 36622
rect 10133 36619 10199 36622
rect 10320 36680 10751 36682
rect 10320 36624 10690 36680
rect 10746 36624 10751 36680
rect 10320 36622 10751 36624
rect 0 36546 400 36576
rect 1117 36546 1183 36549
rect 0 36544 1183 36546
rect 0 36488 1122 36544
rect 1178 36488 1183 36544
rect 0 36486 1183 36488
rect 0 36456 400 36486
rect 1117 36483 1183 36486
rect 5625 36546 5691 36549
rect 7046 36546 7052 36548
rect 5625 36544 7052 36546
rect 5625 36488 5630 36544
rect 5686 36488 7052 36544
rect 5625 36486 7052 36488
rect 5625 36483 5691 36486
rect 7046 36484 7052 36486
rect 7116 36484 7122 36548
rect 7833 36546 7899 36549
rect 8937 36546 9003 36549
rect 7833 36544 9003 36546
rect 7833 36488 7838 36544
rect 7894 36488 8942 36544
rect 8998 36488 9003 36544
rect 7833 36486 9003 36488
rect 7833 36483 7899 36486
rect 8937 36483 9003 36486
rect 9765 36544 9831 36549
rect 9765 36488 9770 36544
rect 9826 36488 9831 36544
rect 9765 36483 9831 36488
rect 4318 36480 4634 36481
rect 4318 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4634 36480
rect 4318 36415 4634 36416
rect 5349 36410 5415 36413
rect 6913 36410 6979 36413
rect 5349 36408 6979 36410
rect 5349 36352 5354 36408
rect 5410 36352 6918 36408
rect 6974 36352 6979 36408
rect 5349 36350 6979 36352
rect 5349 36347 5415 36350
rect 6913 36347 6979 36350
rect 7281 36410 7347 36413
rect 9397 36410 9463 36413
rect 7281 36408 9463 36410
rect 7281 36352 7286 36408
rect 7342 36352 9402 36408
rect 9458 36352 9463 36408
rect 7281 36350 9463 36352
rect 7281 36347 7347 36350
rect 9397 36347 9463 36350
rect 0 36274 400 36304
rect 9768 36277 9828 36483
rect 841 36274 907 36277
rect 0 36272 907 36274
rect 0 36216 846 36272
rect 902 36216 907 36272
rect 0 36214 907 36216
rect 0 36184 400 36214
rect 841 36211 907 36214
rect 3969 36274 4035 36277
rect 7649 36274 7715 36277
rect 3969 36272 7715 36274
rect 3969 36216 3974 36272
rect 4030 36216 7654 36272
rect 7710 36216 7715 36272
rect 3969 36214 7715 36216
rect 3969 36211 4035 36214
rect 7649 36211 7715 36214
rect 8201 36274 8267 36277
rect 9029 36274 9095 36277
rect 8201 36272 9095 36274
rect 8201 36216 8206 36272
rect 8262 36216 9034 36272
rect 9090 36216 9095 36272
rect 8201 36214 9095 36216
rect 8201 36211 8267 36214
rect 9029 36211 9095 36214
rect 9765 36272 9831 36277
rect 9765 36216 9770 36272
rect 9826 36216 9831 36272
rect 9765 36211 9831 36216
rect 5533 36138 5599 36141
rect 2730 36136 5599 36138
rect 2730 36080 5538 36136
rect 5594 36080 5599 36136
rect 2730 36078 5599 36080
rect 1669 35866 1735 35869
rect 2730 35866 2790 36078
rect 5533 36075 5599 36078
rect 7782 36076 7788 36140
rect 7852 36138 7858 36140
rect 8201 36138 8267 36141
rect 10133 36138 10199 36141
rect 10320 36138 10380 36622
rect 10685 36619 10751 36622
rect 10718 36480 11034 36481
rect 10718 36416 10724 36480
rect 10788 36416 10804 36480
rect 10868 36416 10884 36480
rect 10948 36416 10964 36480
rect 11028 36416 11034 36480
rect 10718 36415 11034 36416
rect 10961 36274 11027 36277
rect 12157 36274 12223 36277
rect 10961 36272 12223 36274
rect 10961 36216 10966 36272
rect 11022 36216 12162 36272
rect 12218 36216 12223 36272
rect 10961 36214 12223 36216
rect 10961 36211 11027 36214
rect 12157 36211 12223 36214
rect 7852 36136 9736 36138
rect 7852 36080 8206 36136
rect 8262 36080 9736 36136
rect 7852 36078 9736 36080
rect 7852 36076 7858 36078
rect 8201 36075 8267 36078
rect 9676 36005 9736 36078
rect 10133 36136 10380 36138
rect 10133 36080 10138 36136
rect 10194 36080 10380 36136
rect 10133 36078 10380 36080
rect 10869 36138 10935 36141
rect 11421 36138 11487 36141
rect 10869 36136 11487 36138
rect 10869 36080 10874 36136
rect 10930 36080 11426 36136
rect 11482 36080 11487 36136
rect 10869 36078 11487 36080
rect 10133 36075 10199 36078
rect 10869 36075 10935 36078
rect 11421 36075 11487 36078
rect 4981 36002 5047 36005
rect 5574 36002 5580 36004
rect 4981 36000 5580 36002
rect 4981 35944 4986 36000
rect 5042 35944 5580 36000
rect 4981 35942 5580 35944
rect 4981 35939 5047 35942
rect 5574 35940 5580 35942
rect 5644 36002 5650 36004
rect 7465 36002 7531 36005
rect 5644 36000 7531 36002
rect 5644 35944 7470 36000
rect 7526 35944 7531 36000
rect 5644 35942 7531 35944
rect 5644 35940 5650 35942
rect 7465 35939 7531 35942
rect 9673 36000 9739 36005
rect 9673 35944 9678 36000
rect 9734 35944 9739 36000
rect 9673 35939 9739 35944
rect 3658 35936 3974 35937
rect 3658 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3974 35936
rect 3658 35871 3974 35872
rect 10058 35936 10374 35937
rect 10058 35872 10064 35936
rect 10128 35872 10144 35936
rect 10208 35872 10224 35936
rect 10288 35872 10304 35936
rect 10368 35872 10374 35936
rect 10058 35871 10374 35872
rect 1669 35864 2790 35866
rect 1669 35808 1674 35864
rect 1730 35808 2790 35864
rect 1669 35806 2790 35808
rect 4705 35866 4771 35869
rect 5349 35866 5415 35869
rect 5809 35868 5875 35869
rect 5758 35866 5764 35868
rect 4705 35864 5415 35866
rect 4705 35808 4710 35864
rect 4766 35808 5354 35864
rect 5410 35808 5415 35864
rect 4705 35806 5415 35808
rect 5718 35806 5764 35866
rect 5828 35864 5875 35868
rect 5870 35808 5875 35864
rect 1669 35803 1735 35806
rect 4705 35803 4771 35806
rect 5349 35803 5415 35806
rect 5758 35804 5764 35806
rect 5828 35804 5875 35808
rect 5809 35803 5875 35804
rect 6453 35866 6519 35869
rect 8661 35866 8727 35869
rect 6453 35864 8727 35866
rect 6453 35808 6458 35864
rect 6514 35808 8666 35864
rect 8722 35808 8727 35864
rect 6453 35806 8727 35808
rect 6453 35803 6519 35806
rect 8661 35803 8727 35806
rect 9029 35866 9095 35869
rect 9029 35864 9322 35866
rect 9029 35808 9034 35864
rect 9090 35808 9322 35864
rect 9029 35806 9322 35808
rect 9029 35803 9095 35806
rect 2037 35730 2103 35733
rect 9121 35730 9187 35733
rect 2037 35728 9187 35730
rect 2037 35672 2042 35728
rect 2098 35672 9126 35728
rect 9182 35672 9187 35728
rect 2037 35670 9187 35672
rect 9262 35730 9322 35806
rect 10593 35730 10659 35733
rect 9262 35728 10659 35730
rect 9262 35672 10598 35728
rect 10654 35672 10659 35728
rect 9262 35670 10659 35672
rect 2037 35667 2103 35670
rect 9121 35667 9187 35670
rect 10593 35667 10659 35670
rect 1025 35594 1091 35597
rect 5441 35594 5507 35597
rect 1025 35592 5507 35594
rect 1025 35536 1030 35592
rect 1086 35536 5446 35592
rect 5502 35536 5507 35592
rect 1025 35534 5507 35536
rect 1025 35531 1091 35534
rect 5441 35531 5507 35534
rect 5625 35594 5691 35597
rect 7281 35594 7347 35597
rect 5625 35592 7347 35594
rect 5625 35536 5630 35592
rect 5686 35536 7286 35592
rect 7342 35536 7347 35592
rect 5625 35534 7347 35536
rect 5625 35531 5691 35534
rect 7281 35531 7347 35534
rect 7598 35532 7604 35596
rect 7668 35594 7674 35596
rect 8109 35594 8175 35597
rect 7668 35592 8175 35594
rect 7668 35536 8114 35592
rect 8170 35536 8175 35592
rect 7668 35534 8175 35536
rect 7668 35532 7674 35534
rect 8109 35531 8175 35534
rect 8293 35594 8359 35597
rect 9581 35594 9647 35597
rect 8293 35592 9647 35594
rect 8293 35536 8298 35592
rect 8354 35536 9586 35592
rect 9642 35536 9647 35592
rect 8293 35534 9647 35536
rect 8293 35531 8359 35534
rect 9581 35531 9647 35534
rect 9806 35532 9812 35596
rect 9876 35594 9882 35596
rect 10317 35594 10383 35597
rect 9876 35592 10383 35594
rect 9876 35536 10322 35592
rect 10378 35536 10383 35592
rect 9876 35534 10383 35536
rect 9876 35532 9882 35534
rect 10317 35531 10383 35534
rect 3366 35396 3372 35460
rect 3436 35458 3442 35460
rect 4061 35458 4127 35461
rect 3436 35456 4127 35458
rect 3436 35400 4066 35456
rect 4122 35400 4127 35456
rect 3436 35398 4127 35400
rect 3436 35396 3442 35398
rect 4061 35395 4127 35398
rect 4889 35458 4955 35461
rect 6177 35458 6243 35461
rect 4889 35456 6243 35458
rect 4889 35400 4894 35456
rect 4950 35400 6182 35456
rect 6238 35400 6243 35456
rect 4889 35398 6243 35400
rect 4889 35395 4955 35398
rect 6177 35395 6243 35398
rect 9121 35458 9187 35461
rect 10409 35458 10475 35461
rect 9121 35456 10475 35458
rect 9121 35400 9126 35456
rect 9182 35400 10414 35456
rect 10470 35400 10475 35456
rect 9121 35398 10475 35400
rect 9121 35395 9187 35398
rect 10409 35395 10475 35398
rect 4318 35392 4634 35393
rect 4318 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4634 35392
rect 4318 35327 4634 35328
rect 10718 35392 11034 35393
rect 10718 35328 10724 35392
rect 10788 35328 10804 35392
rect 10868 35328 10884 35392
rect 10948 35328 10964 35392
rect 11028 35328 11034 35392
rect 10718 35327 11034 35328
rect 2589 35322 2655 35325
rect 2998 35322 3004 35324
rect 2589 35320 3004 35322
rect 2589 35264 2594 35320
rect 2650 35264 3004 35320
rect 2589 35262 3004 35264
rect 2589 35259 2655 35262
rect 2998 35260 3004 35262
rect 3068 35322 3074 35324
rect 3601 35322 3667 35325
rect 3068 35320 3667 35322
rect 3068 35264 3606 35320
rect 3662 35264 3667 35320
rect 3068 35262 3667 35264
rect 3068 35260 3074 35262
rect 3601 35259 3667 35262
rect 5993 35322 6059 35325
rect 6862 35322 6868 35324
rect 5993 35320 6868 35322
rect 5993 35264 5998 35320
rect 6054 35264 6868 35320
rect 5993 35262 6868 35264
rect 5993 35259 6059 35262
rect 6862 35260 6868 35262
rect 6932 35260 6938 35324
rect 9438 35260 9444 35324
rect 9508 35322 9514 35324
rect 9806 35322 9812 35324
rect 9508 35262 9812 35322
rect 9508 35260 9514 35262
rect 9806 35260 9812 35262
rect 9876 35260 9882 35324
rect 3049 35186 3115 35189
rect 8293 35186 8359 35189
rect 3049 35184 8359 35186
rect 3049 35128 3054 35184
rect 3110 35128 8298 35184
rect 8354 35128 8359 35184
rect 3049 35126 8359 35128
rect 3049 35123 3115 35126
rect 8293 35123 8359 35126
rect 10041 35186 10107 35189
rect 11697 35186 11763 35189
rect 10041 35184 11763 35186
rect 10041 35128 10046 35184
rect 10102 35128 11702 35184
rect 11758 35128 11763 35184
rect 10041 35126 11763 35128
rect 10041 35123 10107 35126
rect 11697 35123 11763 35126
rect 1761 35050 1827 35053
rect 1894 35050 1900 35052
rect 1761 35048 1900 35050
rect 1761 34992 1766 35048
rect 1822 34992 1900 35048
rect 1761 34990 1900 34992
rect 1761 34987 1827 34990
rect 1894 34988 1900 34990
rect 1964 34988 1970 35052
rect 4153 35050 4219 35053
rect 11094 35050 11100 35052
rect 4153 35048 11100 35050
rect 4153 34992 4158 35048
rect 4214 34992 11100 35048
rect 4153 34990 11100 34992
rect 4153 34987 4219 34990
rect 11094 34988 11100 34990
rect 11164 34988 11170 35052
rect 0 34914 400 34944
rect 473 34914 539 34917
rect 0 34912 539 34914
rect 0 34856 478 34912
rect 534 34856 539 34912
rect 0 34854 539 34856
rect 0 34824 400 34854
rect 473 34851 539 34854
rect 4889 34914 4955 34917
rect 5349 34914 5415 34917
rect 4889 34912 5415 34914
rect 4889 34856 4894 34912
rect 4950 34856 5354 34912
rect 5410 34856 5415 34912
rect 4889 34854 5415 34856
rect 4889 34851 4955 34854
rect 5349 34851 5415 34854
rect 3658 34848 3974 34849
rect 3658 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3974 34848
rect 3658 34783 3974 34784
rect 10058 34848 10374 34849
rect 10058 34784 10064 34848
rect 10128 34784 10144 34848
rect 10208 34784 10224 34848
rect 10288 34784 10304 34848
rect 10368 34784 10374 34848
rect 10058 34783 10374 34784
rect 4061 34778 4127 34781
rect 5993 34778 6059 34781
rect 8569 34778 8635 34781
rect 4061 34776 5044 34778
rect 4061 34720 4066 34776
rect 4122 34720 5044 34776
rect 4061 34718 5044 34720
rect 4061 34715 4127 34718
rect 0 34645 400 34672
rect 0 34640 447 34645
rect 0 34584 386 34640
rect 442 34584 447 34640
rect 0 34579 447 34584
rect 3049 34642 3115 34645
rect 4838 34642 4844 34644
rect 3049 34640 4844 34642
rect 3049 34584 3054 34640
rect 3110 34584 4844 34640
rect 3049 34582 4844 34584
rect 3049 34579 3115 34582
rect 4838 34580 4844 34582
rect 4908 34580 4914 34644
rect 4984 34642 5044 34718
rect 5993 34776 8635 34778
rect 5993 34720 5998 34776
rect 6054 34720 8574 34776
rect 8630 34720 8635 34776
rect 5993 34718 8635 34720
rect 5993 34715 6059 34718
rect 8569 34715 8635 34718
rect 5533 34642 5599 34645
rect 4984 34640 5599 34642
rect 4984 34584 5538 34640
rect 5594 34584 5599 34640
rect 4984 34582 5599 34584
rect 5533 34579 5599 34582
rect 6361 34642 6427 34645
rect 8201 34642 8267 34645
rect 6361 34640 8267 34642
rect 6361 34584 6366 34640
rect 6422 34584 8206 34640
rect 8262 34584 8267 34640
rect 6361 34582 8267 34584
rect 6361 34579 6427 34582
rect 8201 34579 8267 34582
rect 8753 34642 8819 34645
rect 11881 34642 11947 34645
rect 8753 34640 11947 34642
rect 8753 34584 8758 34640
rect 8814 34584 11886 34640
rect 11942 34584 11947 34640
rect 8753 34582 11947 34584
rect 8753 34579 8819 34582
rect 11881 34579 11947 34582
rect 0 34552 400 34579
rect 3417 34506 3483 34509
rect 4102 34506 4108 34508
rect 3374 34504 4108 34506
rect 3374 34448 3422 34504
rect 3478 34448 4108 34504
rect 3374 34446 4108 34448
rect 3374 34443 3483 34446
rect 4102 34444 4108 34446
rect 4172 34444 4178 34508
rect 5441 34506 5507 34509
rect 11145 34506 11211 34509
rect 5441 34504 11211 34506
rect 5441 34448 5446 34504
rect 5502 34448 11150 34504
rect 11206 34448 11211 34504
rect 5441 34446 11211 34448
rect 5441 34443 5507 34446
rect 11145 34443 11211 34446
rect 0 34370 400 34400
rect 933 34370 999 34373
rect 0 34368 999 34370
rect 0 34312 938 34368
rect 994 34312 999 34368
rect 0 34310 999 34312
rect 0 34280 400 34310
rect 933 34307 999 34310
rect 1158 34308 1164 34372
rect 1228 34370 1234 34372
rect 3374 34370 3434 34443
rect 3785 34370 3851 34373
rect 1228 34310 3434 34370
rect 3558 34368 3851 34370
rect 3558 34312 3790 34368
rect 3846 34312 3851 34368
rect 3558 34310 3851 34312
rect 1228 34308 1234 34310
rect 2497 34234 2563 34237
rect 3558 34234 3618 34310
rect 3785 34307 3851 34310
rect 6637 34370 6703 34373
rect 6862 34370 6868 34372
rect 6637 34368 6868 34370
rect 6637 34312 6642 34368
rect 6698 34312 6868 34368
rect 6637 34310 6868 34312
rect 6637 34307 6703 34310
rect 6862 34308 6868 34310
rect 6932 34308 6938 34372
rect 4318 34304 4634 34305
rect 4318 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4634 34304
rect 4318 34239 4634 34240
rect 10718 34304 11034 34305
rect 10718 34240 10724 34304
rect 10788 34240 10804 34304
rect 10868 34240 10884 34304
rect 10948 34240 10964 34304
rect 11028 34240 11034 34304
rect 10718 34239 11034 34240
rect 2497 34232 3618 34234
rect 2497 34176 2502 34232
rect 2558 34176 3618 34232
rect 2497 34174 3618 34176
rect 3693 34234 3759 34237
rect 4102 34234 4108 34236
rect 3693 34232 4108 34234
rect 3693 34176 3698 34232
rect 3754 34176 4108 34232
rect 3693 34174 4108 34176
rect 2497 34171 2563 34174
rect 3693 34171 3759 34174
rect 4102 34172 4108 34174
rect 4172 34172 4178 34236
rect 5441 34234 5507 34237
rect 7925 34234 7991 34237
rect 5441 34232 7991 34234
rect 5441 34176 5446 34232
rect 5502 34176 7930 34232
rect 7986 34176 7991 34232
rect 5441 34174 7991 34176
rect 5441 34171 5507 34174
rect 7925 34171 7991 34174
rect 8385 34098 8451 34101
rect 9673 34098 9739 34101
rect 8385 34096 9739 34098
rect 8385 34040 8390 34096
rect 8446 34040 9678 34096
rect 9734 34040 9739 34096
rect 8385 34038 9739 34040
rect 8385 34035 8451 34038
rect 9673 34035 9739 34038
rect 10041 34098 10107 34101
rect 11421 34098 11487 34101
rect 10041 34096 11487 34098
rect 10041 34040 10046 34096
rect 10102 34040 11426 34096
rect 11482 34040 11487 34096
rect 10041 34038 11487 34040
rect 10041 34035 10107 34038
rect 11421 34035 11487 34038
rect 3325 33962 3391 33965
rect 3969 33962 4035 33965
rect 6862 33962 6868 33964
rect 3325 33960 6868 33962
rect 3325 33904 3330 33960
rect 3386 33904 3974 33960
rect 4030 33904 6868 33960
rect 3325 33902 6868 33904
rect 3325 33899 3391 33902
rect 3969 33899 4035 33902
rect 6862 33900 6868 33902
rect 6932 33900 6938 33964
rect 9673 33962 9739 33965
rect 11053 33962 11119 33965
rect 11513 33962 11579 33965
rect 9673 33960 11579 33962
rect 9673 33904 9678 33960
rect 9734 33904 11058 33960
rect 11114 33904 11518 33960
rect 11574 33904 11579 33960
rect 9673 33902 11579 33904
rect 9673 33899 9739 33902
rect 11053 33899 11119 33902
rect 11513 33899 11579 33902
rect 6085 33826 6151 33829
rect 9254 33826 9260 33828
rect 6085 33824 9260 33826
rect 6085 33768 6090 33824
rect 6146 33768 9260 33824
rect 6085 33766 9260 33768
rect 6085 33763 6151 33766
rect 9254 33764 9260 33766
rect 9324 33764 9330 33828
rect 3658 33760 3974 33761
rect 3658 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3974 33760
rect 3658 33695 3974 33696
rect 10058 33760 10374 33761
rect 10058 33696 10064 33760
rect 10128 33696 10144 33760
rect 10208 33696 10224 33760
rect 10288 33696 10304 33760
rect 10368 33696 10374 33760
rect 10058 33695 10374 33696
rect 1853 33690 1919 33693
rect 2078 33690 2084 33692
rect 1853 33688 2084 33690
rect 1853 33632 1858 33688
rect 1914 33632 2084 33688
rect 1853 33630 2084 33632
rect 1853 33627 1919 33630
rect 2078 33628 2084 33630
rect 2148 33628 2154 33692
rect 4889 33690 4955 33693
rect 5206 33690 5212 33692
rect 4889 33688 5212 33690
rect 4889 33632 4894 33688
rect 4950 33632 5212 33688
rect 4889 33630 5212 33632
rect 4889 33627 4955 33630
rect 5206 33628 5212 33630
rect 5276 33628 5282 33692
rect 5625 33690 5691 33693
rect 6361 33690 6427 33693
rect 11881 33692 11947 33693
rect 5625 33688 6427 33690
rect 5625 33632 5630 33688
rect 5686 33632 6366 33688
rect 6422 33632 6427 33688
rect 5625 33630 6427 33632
rect 5625 33627 5691 33630
rect 6361 33627 6427 33630
rect 8334 33628 8340 33692
rect 8404 33690 8410 33692
rect 9254 33690 9260 33692
rect 8404 33630 9260 33690
rect 8404 33628 8410 33630
rect 9254 33628 9260 33630
rect 9324 33628 9330 33692
rect 11830 33628 11836 33692
rect 11900 33690 11947 33692
rect 11900 33688 11992 33690
rect 11942 33632 11992 33688
rect 11900 33630 11992 33632
rect 11900 33628 11947 33630
rect 11881 33627 11947 33628
rect 1526 33492 1532 33556
rect 1596 33554 1602 33556
rect 1596 33494 2698 33554
rect 1596 33492 1602 33494
rect 2078 33356 2084 33420
rect 2148 33418 2154 33420
rect 2313 33418 2379 33421
rect 2148 33416 2379 33418
rect 2148 33360 2318 33416
rect 2374 33360 2379 33416
rect 2148 33358 2379 33360
rect 2638 33418 2698 33494
rect 5206 33492 5212 33556
rect 5276 33554 5282 33556
rect 5758 33554 5764 33556
rect 5276 33494 5764 33554
rect 5276 33492 5282 33494
rect 5758 33492 5764 33494
rect 5828 33492 5834 33556
rect 9029 33554 9095 33557
rect 10501 33554 10567 33557
rect 9029 33552 10567 33554
rect 9029 33496 9034 33552
rect 9090 33496 10506 33552
rect 10562 33496 10567 33552
rect 9029 33494 10567 33496
rect 9029 33491 9095 33494
rect 10501 33491 10567 33494
rect 11830 33492 11836 33556
rect 11900 33554 11906 33556
rect 11973 33554 12039 33557
rect 11900 33552 12039 33554
rect 11900 33496 11978 33552
rect 12034 33496 12039 33552
rect 11900 33494 12039 33496
rect 11900 33492 11906 33494
rect 11973 33491 12039 33494
rect 2814 33418 2820 33420
rect 2638 33358 2820 33418
rect 2148 33356 2154 33358
rect 2313 33355 2379 33358
rect 2814 33356 2820 33358
rect 2884 33356 2890 33420
rect 4838 33356 4844 33420
rect 4908 33418 4914 33420
rect 5441 33418 5507 33421
rect 4908 33416 5507 33418
rect 4908 33360 5446 33416
rect 5502 33360 5507 33416
rect 4908 33358 5507 33360
rect 4908 33356 4914 33358
rect 5441 33355 5507 33358
rect 5942 33356 5948 33420
rect 6012 33418 6018 33420
rect 6361 33418 6427 33421
rect 6012 33416 6427 33418
rect 6012 33360 6366 33416
rect 6422 33360 6427 33416
rect 6012 33358 6427 33360
rect 6012 33356 6018 33358
rect 6361 33355 6427 33358
rect 6637 33418 6703 33421
rect 7557 33418 7623 33421
rect 6637 33416 7623 33418
rect 6637 33360 6642 33416
rect 6698 33360 7562 33416
rect 7618 33360 7623 33416
rect 6637 33358 7623 33360
rect 6637 33355 6703 33358
rect 7557 33355 7623 33358
rect 1945 33282 2011 33285
rect 2446 33282 2452 33284
rect 1945 33280 2452 33282
rect 1945 33224 1950 33280
rect 2006 33224 2452 33280
rect 1945 33222 2452 33224
rect 1945 33219 2011 33222
rect 2446 33220 2452 33222
rect 2516 33220 2522 33284
rect 6821 33282 6887 33285
rect 7782 33282 7788 33284
rect 6821 33280 7788 33282
rect 6821 33224 6826 33280
rect 6882 33224 7788 33280
rect 6821 33222 7788 33224
rect 6821 33219 6887 33222
rect 7782 33220 7788 33222
rect 7852 33220 7858 33284
rect 4318 33216 4634 33217
rect 4318 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4634 33216
rect 4318 33151 4634 33152
rect 10718 33216 11034 33217
rect 10718 33152 10724 33216
rect 10788 33152 10804 33216
rect 10868 33152 10884 33216
rect 10948 33152 10964 33216
rect 11028 33152 11034 33216
rect 10718 33151 11034 33152
rect 2589 33146 2655 33149
rect 2865 33146 2931 33149
rect 2589 33144 2931 33146
rect 2589 33088 2594 33144
rect 2650 33088 2870 33144
rect 2926 33088 2931 33144
rect 2589 33086 2931 33088
rect 2589 33083 2655 33086
rect 2865 33083 2931 33086
rect 6729 33146 6795 33149
rect 6729 33144 9184 33146
rect 6729 33088 6734 33144
rect 6790 33088 9184 33144
rect 6729 33086 9184 33088
rect 6729 33083 6795 33086
rect 9124 33013 9184 33086
rect 2681 33010 2747 33013
rect 2865 33010 2931 33013
rect 2681 33008 2931 33010
rect 2681 32952 2686 33008
rect 2742 32952 2870 33008
rect 2926 32952 2931 33008
rect 2681 32950 2931 32952
rect 2681 32947 2747 32950
rect 2865 32947 2931 32950
rect 4889 33010 4955 33013
rect 9121 33010 9187 33013
rect 10869 33010 10935 33013
rect 4889 33008 6194 33010
rect 4889 32952 4894 33008
rect 4950 32952 6194 33008
rect 4889 32950 6194 32952
rect 4889 32947 4955 32950
rect 5349 32876 5415 32877
rect 5349 32872 5396 32876
rect 5460 32874 5466 32876
rect 6134 32874 6194 32950
rect 9121 33008 10935 33010
rect 9121 32952 9126 33008
rect 9182 32952 10874 33008
rect 10930 32952 10935 33008
rect 9121 32950 10935 32952
rect 9121 32947 9187 32950
rect 10869 32947 10935 32950
rect 11605 32874 11671 32877
rect 5349 32816 5354 32872
rect 5349 32812 5396 32816
rect 5460 32814 5506 32874
rect 6134 32872 11671 32874
rect 6134 32816 11610 32872
rect 11666 32816 11671 32872
rect 6134 32814 11671 32816
rect 5460 32812 5466 32814
rect 5349 32811 5415 32812
rect 11605 32811 11671 32814
rect 4429 32738 4495 32741
rect 6729 32738 6795 32741
rect 4429 32736 6795 32738
rect 4429 32680 4434 32736
rect 4490 32680 6734 32736
rect 6790 32680 6795 32736
rect 4429 32678 6795 32680
rect 4429 32675 4495 32678
rect 6729 32675 6795 32678
rect 6862 32676 6868 32740
rect 6932 32738 6938 32740
rect 7281 32738 7347 32741
rect 8334 32738 8340 32740
rect 6932 32736 8340 32738
rect 6932 32680 7286 32736
rect 7342 32680 8340 32736
rect 6932 32678 8340 32680
rect 6932 32676 6938 32678
rect 7281 32675 7347 32678
rect 8334 32676 8340 32678
rect 8404 32676 8410 32740
rect 8937 32738 9003 32741
rect 9438 32738 9444 32740
rect 8937 32736 9444 32738
rect 8937 32680 8942 32736
rect 8998 32680 9444 32736
rect 8937 32678 9444 32680
rect 8937 32675 9003 32678
rect 9438 32676 9444 32678
rect 9508 32676 9514 32740
rect 3658 32672 3974 32673
rect 3658 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3974 32672
rect 3658 32607 3974 32608
rect 10058 32672 10374 32673
rect 10058 32608 10064 32672
rect 10128 32608 10144 32672
rect 10208 32608 10224 32672
rect 10288 32608 10304 32672
rect 10368 32608 10374 32672
rect 10058 32607 10374 32608
rect 5073 32602 5139 32605
rect 6494 32602 6500 32604
rect 5073 32600 6500 32602
rect 5073 32544 5078 32600
rect 5134 32544 6500 32600
rect 5073 32542 6500 32544
rect 5073 32539 5139 32542
rect 6494 32540 6500 32542
rect 6564 32540 6570 32604
rect 6729 32602 6795 32605
rect 7230 32602 7236 32604
rect 6729 32600 7236 32602
rect 6729 32544 6734 32600
rect 6790 32544 7236 32600
rect 6729 32542 7236 32544
rect 6729 32539 6795 32542
rect 7230 32540 7236 32542
rect 7300 32540 7306 32604
rect 8293 32600 8359 32605
rect 8293 32544 8298 32600
rect 8354 32544 8359 32600
rect 8293 32539 8359 32544
rect 8753 32602 8819 32605
rect 9857 32602 9923 32605
rect 8753 32600 9923 32602
rect 8753 32544 8758 32600
rect 8814 32544 9862 32600
rect 9918 32544 9923 32600
rect 8753 32542 9923 32544
rect 8753 32539 8819 32542
rect 9857 32539 9923 32542
rect 3182 32404 3188 32468
rect 3252 32466 3258 32468
rect 5390 32466 5396 32468
rect 3252 32406 5396 32466
rect 3252 32404 3258 32406
rect 5390 32404 5396 32406
rect 5460 32404 5466 32468
rect 6126 32404 6132 32468
rect 6196 32466 6202 32468
rect 8296 32466 8356 32539
rect 9673 32466 9739 32469
rect 6196 32464 9739 32466
rect 6196 32408 9678 32464
rect 9734 32408 9739 32464
rect 6196 32406 9739 32408
rect 6196 32404 6202 32406
rect 9673 32403 9739 32406
rect 10317 32466 10383 32469
rect 10501 32466 10567 32469
rect 10317 32464 10567 32466
rect 10317 32408 10322 32464
rect 10378 32408 10506 32464
rect 10562 32408 10567 32464
rect 10317 32406 10567 32408
rect 10317 32403 10383 32406
rect 10501 32403 10567 32406
rect 790 32268 796 32332
rect 860 32330 866 32332
rect 1342 32330 1348 32332
rect 860 32270 1348 32330
rect 860 32268 866 32270
rect 1342 32268 1348 32270
rect 1412 32330 1418 32332
rect 6361 32330 6427 32333
rect 6821 32332 6887 32333
rect 6821 32330 6868 32332
rect 1412 32328 6427 32330
rect 1412 32272 6366 32328
rect 6422 32272 6427 32328
rect 1412 32270 6427 32272
rect 6776 32328 6868 32330
rect 6776 32272 6826 32328
rect 6776 32270 6868 32272
rect 1412 32268 1418 32270
rect 6361 32267 6427 32270
rect 6821 32268 6868 32270
rect 6932 32268 6938 32332
rect 7281 32330 7347 32333
rect 11789 32330 11855 32333
rect 7281 32328 11855 32330
rect 7281 32272 7286 32328
rect 7342 32272 11794 32328
rect 11850 32272 11855 32328
rect 7281 32270 11855 32272
rect 6821 32267 6887 32268
rect 7281 32267 7347 32270
rect 11789 32267 11855 32270
rect 1342 32132 1348 32196
rect 1412 32194 1418 32196
rect 1853 32194 1919 32197
rect 1412 32192 1919 32194
rect 1412 32136 1858 32192
rect 1914 32136 1919 32192
rect 1412 32134 1919 32136
rect 1412 32132 1418 32134
rect 1853 32131 1919 32134
rect 5809 32194 5875 32197
rect 6269 32194 6335 32197
rect 7557 32196 7623 32197
rect 7557 32194 7604 32196
rect 5809 32192 6335 32194
rect 5809 32136 5814 32192
rect 5870 32136 6274 32192
rect 6330 32136 6335 32192
rect 5809 32134 6335 32136
rect 7512 32192 7604 32194
rect 7512 32136 7562 32192
rect 7512 32134 7604 32136
rect 5809 32131 5875 32134
rect 6269 32131 6335 32134
rect 7557 32132 7604 32134
rect 7668 32132 7674 32196
rect 7833 32194 7899 32197
rect 9673 32194 9739 32197
rect 10542 32194 10548 32196
rect 7833 32192 10548 32194
rect 7833 32136 7838 32192
rect 7894 32136 9678 32192
rect 9734 32136 10548 32192
rect 7833 32134 10548 32136
rect 7557 32131 7623 32132
rect 7833 32131 7899 32134
rect 9673 32131 9739 32134
rect 10542 32132 10548 32134
rect 10612 32132 10618 32196
rect 4318 32128 4634 32129
rect 4318 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4634 32128
rect 4318 32063 4634 32064
rect 10718 32128 11034 32129
rect 10718 32064 10724 32128
rect 10788 32064 10804 32128
rect 10868 32064 10884 32128
rect 10948 32064 10964 32128
rect 11028 32064 11034 32128
rect 10718 32063 11034 32064
rect 749 32058 815 32061
rect 5165 32058 5231 32061
rect 749 32056 858 32058
rect 749 32000 754 32056
rect 810 32000 858 32056
rect 749 31995 858 32000
rect 798 31922 858 31995
rect 5030 32056 5231 32058
rect 5030 32000 5170 32056
rect 5226 32000 5231 32056
rect 5030 31998 5231 32000
rect 798 31862 4170 31922
rect 657 31786 723 31789
rect 1209 31786 1275 31789
rect 657 31784 1275 31786
rect 657 31728 662 31784
rect 718 31728 1214 31784
rect 1270 31728 1275 31784
rect 657 31726 1275 31728
rect 657 31723 723 31726
rect 1209 31723 1275 31726
rect 2037 31786 2103 31789
rect 2262 31786 2268 31788
rect 2037 31784 2268 31786
rect 2037 31728 2042 31784
rect 2098 31728 2268 31784
rect 2037 31726 2268 31728
rect 2037 31723 2103 31726
rect 2262 31724 2268 31726
rect 2332 31724 2338 31788
rect 4110 31653 4170 31862
rect 5030 31789 5090 31998
rect 5165 31995 5231 31998
rect 7966 31996 7972 32060
rect 8036 32058 8042 32060
rect 8385 32058 8451 32061
rect 8036 32056 8451 32058
rect 8036 32000 8390 32056
rect 8446 32000 8451 32056
rect 8036 31998 8451 32000
rect 8036 31996 8042 31998
rect 8385 31995 8451 31998
rect 8845 32058 8911 32061
rect 9581 32058 9647 32061
rect 8845 32056 9647 32058
rect 8845 32000 8850 32056
rect 8906 32000 9586 32056
rect 9642 32000 9647 32056
rect 8845 31998 9647 32000
rect 8845 31995 8911 31998
rect 9581 31995 9647 31998
rect 11881 32058 11947 32061
rect 12341 32058 12407 32061
rect 11881 32056 12407 32058
rect 11881 32000 11886 32056
rect 11942 32000 12346 32056
rect 12402 32000 12407 32056
rect 11881 31998 12407 32000
rect 11881 31995 11947 31998
rect 12341 31995 12407 31998
rect 7046 31860 7052 31924
rect 7116 31922 7122 31924
rect 7925 31922 7991 31925
rect 7116 31920 7991 31922
rect 7116 31864 7930 31920
rect 7986 31864 7991 31920
rect 7116 31862 7991 31864
rect 7116 31860 7122 31862
rect 7925 31859 7991 31862
rect 10542 31860 10548 31924
rect 10612 31922 10618 31924
rect 11094 31922 11100 31924
rect 10612 31862 11100 31922
rect 10612 31860 10618 31862
rect 11094 31860 11100 31862
rect 11164 31860 11170 31924
rect 12617 31922 12683 31925
rect 12574 31920 12683 31922
rect 12574 31864 12622 31920
rect 12678 31864 12683 31920
rect 12574 31859 12683 31864
rect 4981 31784 5090 31789
rect 5809 31788 5875 31789
rect 4981 31728 4986 31784
rect 5042 31728 5090 31784
rect 4981 31726 5090 31728
rect 4981 31723 5047 31726
rect 5758 31724 5764 31788
rect 5828 31786 5875 31788
rect 5828 31784 5920 31786
rect 5870 31728 5920 31784
rect 5828 31726 5920 31728
rect 5828 31724 5875 31726
rect 6310 31724 6316 31788
rect 6380 31786 6386 31788
rect 6637 31786 6703 31789
rect 6380 31784 6703 31786
rect 6380 31728 6642 31784
rect 6698 31728 6703 31784
rect 6380 31726 6703 31728
rect 6380 31724 6386 31726
rect 5809 31723 5875 31724
rect 6637 31723 6703 31726
rect 8702 31724 8708 31788
rect 8772 31786 8778 31788
rect 9673 31786 9739 31789
rect 8772 31784 9739 31786
rect 8772 31728 9678 31784
rect 9734 31728 9739 31784
rect 8772 31726 9739 31728
rect 8772 31724 8778 31726
rect 9673 31723 9739 31726
rect 11789 31786 11855 31789
rect 12574 31786 12634 31859
rect 11789 31784 12634 31786
rect 11789 31728 11794 31784
rect 11850 31728 12634 31784
rect 11789 31726 12634 31728
rect 11789 31723 11855 31726
rect 1710 31588 1716 31652
rect 1780 31650 1786 31652
rect 3509 31650 3575 31653
rect 1780 31648 3575 31650
rect 1780 31592 3514 31648
rect 3570 31592 3575 31648
rect 1780 31590 3575 31592
rect 4110 31648 4219 31653
rect 5942 31650 5948 31652
rect 4110 31592 4158 31648
rect 4214 31592 4219 31648
rect 4110 31590 4219 31592
rect 1780 31588 1786 31590
rect 3509 31587 3575 31590
rect 4153 31587 4219 31590
rect 5812 31590 5948 31650
rect 3658 31584 3974 31585
rect 3658 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3974 31584
rect 3658 31519 3974 31520
rect 1669 31516 1735 31517
rect 1669 31512 1716 31516
rect 1780 31514 1786 31516
rect 1669 31456 1674 31512
rect 1669 31452 1716 31456
rect 1780 31454 1826 31514
rect 1780 31452 1786 31454
rect 4102 31452 4108 31516
rect 4172 31514 4178 31516
rect 4245 31514 4311 31517
rect 4172 31512 4311 31514
rect 4172 31456 4250 31512
rect 4306 31456 4311 31512
rect 4172 31454 4311 31456
rect 4172 31452 4178 31454
rect 1669 31451 1735 31452
rect 4245 31451 4311 31454
rect 5812 31381 5872 31590
rect 5942 31588 5948 31590
rect 6012 31650 6018 31652
rect 6821 31650 6887 31653
rect 6012 31648 6887 31650
rect 6012 31592 6826 31648
rect 6882 31592 6887 31648
rect 6012 31590 6887 31592
rect 6012 31588 6018 31590
rect 6821 31587 6887 31590
rect 7414 31588 7420 31652
rect 7484 31650 7490 31652
rect 7649 31650 7715 31653
rect 7484 31648 7715 31650
rect 7484 31592 7654 31648
rect 7710 31592 7715 31648
rect 7484 31590 7715 31592
rect 7484 31588 7490 31590
rect 7649 31587 7715 31590
rect 9397 31650 9463 31653
rect 9765 31650 9831 31653
rect 9397 31648 9831 31650
rect 9397 31592 9402 31648
rect 9458 31592 9770 31648
rect 9826 31592 9831 31648
rect 9397 31590 9831 31592
rect 9397 31587 9463 31590
rect 9765 31587 9831 31590
rect 10685 31650 10751 31653
rect 11094 31650 11100 31652
rect 10685 31648 11100 31650
rect 10685 31592 10690 31648
rect 10746 31592 11100 31648
rect 10685 31590 11100 31592
rect 10685 31587 10751 31590
rect 11094 31588 11100 31590
rect 11164 31650 11170 31652
rect 11421 31650 11487 31653
rect 11164 31648 11487 31650
rect 11164 31592 11426 31648
rect 11482 31592 11487 31648
rect 11164 31590 11487 31592
rect 11164 31588 11170 31590
rect 11421 31587 11487 31590
rect 10058 31584 10374 31585
rect 10058 31520 10064 31584
rect 10128 31520 10144 31584
rect 10208 31520 10224 31584
rect 10288 31520 10304 31584
rect 10368 31520 10374 31584
rect 10058 31519 10374 31520
rect 6361 31514 6427 31517
rect 7005 31514 7071 31517
rect 9305 31514 9371 31517
rect 6361 31512 6700 31514
rect 6361 31456 6366 31512
rect 6422 31456 6700 31512
rect 6361 31454 6700 31456
rect 6361 31451 6427 31454
rect 841 31378 907 31381
rect 4102 31378 4108 31380
rect 841 31376 4108 31378
rect 841 31320 846 31376
rect 902 31320 4108 31376
rect 841 31318 4108 31320
rect 841 31315 907 31318
rect 4102 31316 4108 31318
rect 4172 31316 4178 31380
rect 5809 31376 5875 31381
rect 5809 31320 5814 31376
rect 5870 31320 5875 31376
rect 5809 31315 5875 31320
rect 6640 31378 6700 31454
rect 7005 31512 9371 31514
rect 7005 31456 7010 31512
rect 7066 31456 9310 31512
rect 9366 31456 9371 31512
rect 7005 31454 9371 31456
rect 7005 31451 7071 31454
rect 9305 31451 9371 31454
rect 7649 31378 7715 31381
rect 6640 31376 7715 31378
rect 6640 31320 7654 31376
rect 7710 31320 7715 31376
rect 6640 31318 7715 31320
rect 7649 31315 7715 31318
rect 2497 31242 2563 31245
rect 5809 31242 5875 31245
rect 6637 31242 6703 31245
rect 7833 31242 7899 31245
rect 2497 31240 5642 31242
rect 2497 31184 2502 31240
rect 2558 31184 5642 31240
rect 2497 31182 5642 31184
rect 2497 31179 2563 31182
rect 381 31106 447 31109
rect 3141 31106 3207 31109
rect 3325 31108 3391 31109
rect 3325 31106 3372 31108
rect 381 31104 3207 31106
rect 381 31048 386 31104
rect 442 31048 3146 31104
rect 3202 31048 3207 31104
rect 381 31046 3207 31048
rect 3280 31104 3372 31106
rect 3280 31048 3330 31104
rect 3280 31046 3372 31048
rect 381 31043 447 31046
rect 3141 31043 3207 31046
rect 3325 31044 3372 31046
rect 3436 31044 3442 31108
rect 5582 31106 5642 31182
rect 5809 31240 7899 31242
rect 5809 31184 5814 31240
rect 5870 31184 6642 31240
rect 6698 31184 7838 31240
rect 7894 31184 7899 31240
rect 5809 31182 7899 31184
rect 5809 31179 5875 31182
rect 6637 31179 6703 31182
rect 7833 31179 7899 31182
rect 7557 31106 7623 31109
rect 5582 31104 7623 31106
rect 5582 31048 7562 31104
rect 7618 31048 7623 31104
rect 5582 31046 7623 31048
rect 3325 31043 3391 31044
rect 7557 31043 7623 31046
rect 8702 31044 8708 31108
rect 8772 31106 8778 31108
rect 9070 31106 9076 31108
rect 8772 31046 9076 31106
rect 8772 31044 8778 31046
rect 9070 31044 9076 31046
rect 9140 31044 9146 31108
rect 4318 31040 4634 31041
rect 4318 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4634 31040
rect 4318 30975 4634 30976
rect 10718 31040 11034 31041
rect 10718 30976 10724 31040
rect 10788 30976 10804 31040
rect 10868 30976 10884 31040
rect 10948 30976 10964 31040
rect 11028 30976 11034 31040
rect 10718 30975 11034 30976
rect 1393 30970 1459 30973
rect 1393 30968 2330 30970
rect 1393 30912 1398 30968
rect 1454 30912 2330 30968
rect 1393 30910 2330 30912
rect 1393 30907 1459 30910
rect 2270 30428 2330 30910
rect 2865 30968 2931 30973
rect 2865 30912 2870 30968
rect 2926 30912 2931 30968
rect 2865 30907 2931 30912
rect 5809 30970 5875 30973
rect 9254 30970 9260 30972
rect 5809 30968 9260 30970
rect 5809 30912 5814 30968
rect 5870 30912 9260 30968
rect 5809 30910 9260 30912
rect 5809 30907 5875 30910
rect 9254 30908 9260 30910
rect 9324 30908 9330 30972
rect 2868 30834 2928 30907
rect 4245 30834 4311 30837
rect 2868 30832 4311 30834
rect 2868 30776 4250 30832
rect 4306 30776 4311 30832
rect 2868 30774 4311 30776
rect 4245 30771 4311 30774
rect 5758 30772 5764 30836
rect 5828 30834 5834 30836
rect 10225 30834 10291 30837
rect 10777 30834 10843 30837
rect 11881 30834 11947 30837
rect 5828 30832 11947 30834
rect 5828 30776 10230 30832
rect 10286 30776 10782 30832
rect 10838 30776 11886 30832
rect 11942 30776 11947 30832
rect 5828 30774 11947 30776
rect 5828 30772 5834 30774
rect 10225 30771 10291 30774
rect 10777 30771 10843 30774
rect 11881 30771 11947 30774
rect 5717 30698 5783 30701
rect 7097 30698 7163 30701
rect 5717 30696 7163 30698
rect 5717 30640 5722 30696
rect 5778 30640 7102 30696
rect 7158 30640 7163 30696
rect 5717 30638 7163 30640
rect 5717 30635 5783 30638
rect 7097 30635 7163 30638
rect 7414 30636 7420 30700
rect 7484 30698 7490 30700
rect 9070 30698 9076 30700
rect 7484 30638 9076 30698
rect 7484 30636 7490 30638
rect 9070 30636 9076 30638
rect 9140 30636 9146 30700
rect 10041 30698 10107 30701
rect 10041 30696 10564 30698
rect 10041 30640 10046 30696
rect 10102 30640 10564 30696
rect 10041 30638 10564 30640
rect 10041 30635 10107 30638
rect 5022 30500 5028 30564
rect 5092 30562 5098 30564
rect 8845 30562 8911 30565
rect 5092 30560 8911 30562
rect 5092 30504 8850 30560
rect 8906 30504 8911 30560
rect 5092 30502 8911 30504
rect 5092 30500 5098 30502
rect 8845 30499 8911 30502
rect 9254 30500 9260 30564
rect 9324 30562 9330 30564
rect 9857 30562 9923 30565
rect 9324 30560 9923 30562
rect 9324 30504 9862 30560
rect 9918 30504 9923 30560
rect 9324 30502 9923 30504
rect 9324 30500 9330 30502
rect 9857 30499 9923 30502
rect 3658 30496 3974 30497
rect 3658 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3974 30496
rect 3658 30431 3974 30432
rect 10058 30496 10374 30497
rect 10058 30432 10064 30496
rect 10128 30432 10144 30496
rect 10208 30432 10224 30496
rect 10288 30432 10304 30496
rect 10368 30432 10374 30496
rect 10058 30431 10374 30432
rect 2262 30364 2268 30428
rect 2332 30426 2338 30428
rect 5073 30426 5139 30429
rect 5574 30426 5580 30428
rect 2332 30366 2790 30426
rect 2332 30364 2338 30366
rect 2405 30288 2471 30293
rect 2405 30232 2410 30288
rect 2466 30232 2471 30288
rect 2405 30227 2471 30232
rect 2730 30290 2790 30366
rect 5073 30424 5580 30426
rect 5073 30368 5078 30424
rect 5134 30368 5580 30424
rect 5073 30366 5580 30368
rect 5073 30363 5139 30366
rect 5574 30364 5580 30366
rect 5644 30364 5650 30428
rect 5717 30426 5783 30429
rect 7557 30428 7623 30429
rect 6862 30426 6868 30428
rect 5717 30424 6868 30426
rect 5717 30368 5722 30424
rect 5778 30368 6868 30424
rect 5717 30366 6868 30368
rect 5717 30363 5783 30366
rect 6862 30364 6868 30366
rect 6932 30364 6938 30428
rect 7557 30424 7604 30428
rect 7668 30426 7674 30428
rect 7557 30368 7562 30424
rect 7557 30364 7604 30368
rect 7668 30366 7714 30426
rect 7668 30364 7674 30366
rect 8518 30364 8524 30428
rect 8588 30426 8594 30428
rect 9857 30426 9923 30429
rect 8588 30424 9923 30426
rect 8588 30368 9862 30424
rect 9918 30368 9923 30424
rect 8588 30366 9923 30368
rect 8588 30364 8594 30366
rect 7557 30363 7623 30364
rect 9857 30363 9923 30366
rect 4429 30290 4495 30293
rect 2730 30288 4495 30290
rect 2730 30232 4434 30288
rect 4490 30232 4495 30288
rect 2730 30230 4495 30232
rect 4429 30227 4495 30230
rect 4797 30290 4863 30293
rect 5022 30290 5028 30292
rect 4797 30288 5028 30290
rect 4797 30232 4802 30288
rect 4858 30232 5028 30288
rect 4797 30230 5028 30232
rect 4797 30227 4863 30230
rect 5022 30228 5028 30230
rect 5092 30228 5098 30292
rect 5533 30290 5599 30293
rect 5901 30290 5967 30293
rect 5533 30288 5967 30290
rect 5533 30232 5538 30288
rect 5594 30232 5906 30288
rect 5962 30232 5967 30288
rect 5533 30230 5967 30232
rect 5533 30227 5599 30230
rect 5901 30227 5967 30230
rect 6545 30290 6611 30293
rect 7465 30290 7531 30293
rect 8109 30292 8175 30293
rect 8109 30290 8156 30292
rect 6545 30288 7531 30290
rect 6545 30232 6550 30288
rect 6606 30232 7470 30288
rect 7526 30232 7531 30288
rect 6545 30230 7531 30232
rect 8064 30288 8156 30290
rect 8064 30232 8114 30288
rect 8064 30230 8156 30232
rect 6545 30227 6611 30230
rect 7465 30227 7531 30230
rect 8109 30228 8156 30230
rect 8220 30228 8226 30292
rect 9806 30228 9812 30292
rect 9876 30290 9882 30292
rect 10225 30290 10291 30293
rect 9876 30288 10291 30290
rect 9876 30232 10230 30288
rect 10286 30232 10291 30288
rect 9876 30230 10291 30232
rect 9876 30228 9882 30230
rect 8109 30227 8175 30228
rect 10225 30227 10291 30230
rect 2408 30154 2468 30227
rect 2408 30094 2698 30154
rect 1761 29882 1827 29885
rect 1894 29882 1900 29884
rect 1761 29880 1900 29882
rect 1761 29824 1766 29880
rect 1822 29824 1900 29880
rect 1761 29822 1900 29824
rect 1761 29819 1827 29822
rect 1894 29820 1900 29822
rect 1964 29820 1970 29884
rect 2638 29882 2698 30094
rect 2773 30152 2839 30157
rect 2773 30096 2778 30152
rect 2834 30096 2839 30152
rect 2773 30091 2839 30096
rect 3233 30154 3299 30157
rect 3969 30154 4035 30157
rect 4337 30154 4403 30157
rect 3233 30152 4035 30154
rect 3233 30096 3238 30152
rect 3294 30096 3974 30152
rect 4030 30096 4035 30152
rect 3233 30094 4035 30096
rect 3233 30091 3299 30094
rect 3969 30091 4035 30094
rect 4156 30152 4403 30154
rect 4156 30096 4342 30152
rect 4398 30096 4403 30152
rect 4156 30094 4403 30096
rect 2776 30018 2836 30091
rect 3366 30018 3372 30020
rect 2776 29958 3372 30018
rect 3366 29956 3372 29958
rect 3436 29956 3442 30020
rect 3969 30018 4035 30021
rect 4156 30018 4216 30094
rect 4337 30091 4403 30094
rect 4613 30154 4679 30157
rect 5942 30154 5948 30156
rect 4613 30152 5948 30154
rect 4613 30096 4618 30152
rect 4674 30096 5948 30152
rect 4613 30094 5948 30096
rect 4613 30091 4679 30094
rect 5942 30092 5948 30094
rect 6012 30092 6018 30156
rect 6310 30092 6316 30156
rect 6380 30154 6386 30156
rect 7097 30154 7163 30157
rect 6380 30152 7163 30154
rect 6380 30096 7102 30152
rect 7158 30096 7163 30152
rect 6380 30094 7163 30096
rect 6380 30092 6386 30094
rect 7097 30091 7163 30094
rect 7782 30092 7788 30156
rect 7852 30154 7858 30156
rect 8937 30154 9003 30157
rect 7852 30152 9003 30154
rect 7852 30096 8942 30152
rect 8998 30096 9003 30152
rect 7852 30094 9003 30096
rect 7852 30092 7858 30094
rect 8937 30091 9003 30094
rect 10041 30154 10107 30157
rect 10504 30154 10564 30638
rect 10961 30426 11027 30429
rect 11646 30426 11652 30428
rect 10961 30424 11652 30426
rect 10961 30368 10966 30424
rect 11022 30368 11652 30424
rect 10961 30366 11652 30368
rect 10961 30363 11027 30366
rect 11646 30364 11652 30366
rect 11716 30364 11722 30428
rect 11421 30292 11487 30293
rect 11421 30288 11468 30292
rect 11532 30290 11538 30292
rect 11421 30232 11426 30288
rect 11421 30228 11468 30232
rect 11532 30230 11578 30290
rect 11532 30228 11538 30230
rect 11421 30227 11487 30228
rect 10041 30152 10564 30154
rect 10041 30096 10046 30152
rect 10102 30096 10564 30152
rect 10041 30094 10564 30096
rect 10041 30091 10107 30094
rect 5349 30018 5415 30021
rect 6269 30018 6335 30021
rect 3969 30016 4216 30018
rect 3969 29960 3974 30016
rect 4030 29960 4216 30016
rect 3969 29958 4216 29960
rect 5076 30016 6335 30018
rect 5076 29960 5354 30016
rect 5410 29960 6274 30016
rect 6330 29960 6335 30016
rect 5076 29958 6335 29960
rect 3969 29955 4035 29958
rect 4318 29952 4634 29953
rect 4318 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4634 29952
rect 4318 29887 4634 29888
rect 3785 29882 3851 29885
rect 2638 29880 3851 29882
rect 2638 29824 3790 29880
rect 3846 29824 3851 29880
rect 2638 29822 3851 29824
rect 3785 29819 3851 29822
rect 54 29684 60 29748
rect 124 29746 130 29748
rect 4797 29746 4863 29749
rect 124 29744 4863 29746
rect 124 29688 4802 29744
rect 4858 29688 4863 29744
rect 124 29686 4863 29688
rect 124 29684 130 29686
rect 4797 29683 4863 29686
rect 2129 29610 2195 29613
rect 2262 29610 2268 29612
rect 2129 29608 2268 29610
rect 2129 29552 2134 29608
rect 2190 29552 2268 29608
rect 2129 29550 2268 29552
rect 2129 29547 2195 29550
rect 2262 29548 2268 29550
rect 2332 29548 2338 29612
rect 2497 29608 2563 29613
rect 2497 29552 2502 29608
rect 2558 29552 2563 29608
rect 2497 29547 2563 29552
rect 2773 29610 2839 29613
rect 3693 29610 3759 29613
rect 2773 29608 3759 29610
rect 2773 29552 2778 29608
rect 2834 29552 3698 29608
rect 3754 29552 3759 29608
rect 2773 29550 3759 29552
rect 2773 29547 2839 29550
rect 3693 29547 3759 29550
rect 2500 29474 2560 29547
rect 5076 29477 5136 29958
rect 5349 29955 5415 29958
rect 6269 29955 6335 29958
rect 6678 29956 6684 30020
rect 6748 30018 6754 30020
rect 8845 30018 8911 30021
rect 6748 30016 8911 30018
rect 6748 29960 8850 30016
rect 8906 29960 8911 30016
rect 6748 29958 8911 29960
rect 6748 29956 6754 29958
rect 8845 29955 8911 29958
rect 10501 30016 10567 30021
rect 10501 29960 10506 30016
rect 10562 29960 10567 30016
rect 10501 29955 10567 29960
rect 5206 29820 5212 29884
rect 5276 29882 5282 29884
rect 10133 29882 10199 29885
rect 5276 29880 10199 29882
rect 5276 29824 10138 29880
rect 10194 29824 10199 29880
rect 5276 29822 10199 29824
rect 5276 29820 5282 29822
rect 10133 29819 10199 29822
rect 5809 29746 5875 29749
rect 6361 29746 6427 29749
rect 5809 29744 6427 29746
rect 5809 29688 5814 29744
rect 5870 29688 6366 29744
rect 6422 29688 6427 29744
rect 5809 29686 6427 29688
rect 5809 29683 5875 29686
rect 6361 29683 6427 29686
rect 10225 29746 10291 29749
rect 10504 29746 10564 29955
rect 10718 29952 11034 29953
rect 10718 29888 10724 29952
rect 10788 29888 10804 29952
rect 10868 29888 10884 29952
rect 10948 29888 10964 29952
rect 11028 29888 11034 29952
rect 10718 29887 11034 29888
rect 10685 29746 10751 29749
rect 10225 29744 10426 29746
rect 10225 29688 10230 29744
rect 10286 29688 10426 29744
rect 10225 29686 10426 29688
rect 10504 29744 10751 29746
rect 10504 29688 10690 29744
rect 10746 29688 10751 29744
rect 10504 29686 10751 29688
rect 10225 29683 10291 29686
rect 9857 29610 9923 29613
rect 10225 29610 10291 29613
rect 9857 29608 10291 29610
rect 9857 29552 9862 29608
rect 9918 29552 10230 29608
rect 10286 29552 10291 29608
rect 9857 29550 10291 29552
rect 10366 29610 10426 29686
rect 10685 29683 10751 29686
rect 11053 29746 11119 29749
rect 12014 29746 12020 29748
rect 11053 29744 12020 29746
rect 11053 29688 11058 29744
rect 11114 29688 12020 29744
rect 11053 29686 12020 29688
rect 11053 29683 11119 29686
rect 12014 29684 12020 29686
rect 12084 29684 12090 29748
rect 12617 29610 12683 29613
rect 10366 29608 12683 29610
rect 10366 29552 12622 29608
rect 12678 29552 12683 29608
rect 10366 29550 12683 29552
rect 9857 29547 9923 29550
rect 10225 29547 10291 29550
rect 12617 29547 12683 29550
rect 3049 29474 3115 29477
rect 3417 29474 3483 29477
rect 2500 29472 3483 29474
rect 2500 29416 3054 29472
rect 3110 29416 3422 29472
rect 3478 29416 3483 29472
rect 2500 29414 3483 29416
rect 3049 29411 3115 29414
rect 3417 29411 3483 29414
rect 4245 29474 4311 29477
rect 4889 29474 4955 29477
rect 4245 29472 4955 29474
rect 4245 29416 4250 29472
rect 4306 29416 4894 29472
rect 4950 29416 4955 29472
rect 4245 29414 4955 29416
rect 4245 29411 4311 29414
rect 4889 29411 4955 29414
rect 5073 29472 5139 29477
rect 10593 29476 10659 29477
rect 10542 29474 10548 29476
rect 5073 29416 5078 29472
rect 5134 29416 5139 29472
rect 5073 29411 5139 29416
rect 10502 29414 10548 29474
rect 10612 29472 10659 29476
rect 10654 29416 10659 29472
rect 10542 29412 10548 29414
rect 10612 29412 10659 29416
rect 10593 29411 10659 29412
rect 11329 29474 11395 29477
rect 12198 29474 12204 29476
rect 11329 29472 12204 29474
rect 11329 29416 11334 29472
rect 11390 29416 12204 29472
rect 11329 29414 12204 29416
rect 11329 29411 11395 29414
rect 12198 29412 12204 29414
rect 12268 29412 12274 29476
rect 3658 29408 3974 29409
rect 3658 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3974 29408
rect 3658 29343 3974 29344
rect 10058 29408 10374 29409
rect 10058 29344 10064 29408
rect 10128 29344 10144 29408
rect 10208 29344 10224 29408
rect 10288 29344 10304 29408
rect 10368 29344 10374 29408
rect 10058 29343 10374 29344
rect 2865 29340 2931 29341
rect 2814 29276 2820 29340
rect 2884 29338 2931 29340
rect 11053 29338 11119 29341
rect 11278 29338 11284 29340
rect 2884 29336 2976 29338
rect 2926 29280 2976 29336
rect 2884 29278 2976 29280
rect 11053 29336 11284 29338
rect 11053 29280 11058 29336
rect 11114 29280 11284 29336
rect 11053 29278 11284 29280
rect 2884 29276 2931 29278
rect 2865 29275 2931 29276
rect 11053 29275 11119 29278
rect 11278 29276 11284 29278
rect 11348 29276 11354 29340
rect 974 29140 980 29204
rect 1044 29202 1050 29204
rect 2037 29202 2103 29205
rect 2681 29204 2747 29205
rect 2630 29202 2636 29204
rect 1044 29200 2103 29202
rect 1044 29144 2042 29200
rect 2098 29144 2103 29200
rect 1044 29142 2103 29144
rect 2590 29142 2636 29202
rect 2700 29202 2747 29204
rect 3417 29202 3483 29205
rect 7046 29202 7052 29204
rect 2700 29200 3483 29202
rect 2742 29144 3422 29200
rect 3478 29144 3483 29200
rect 1044 29140 1050 29142
rect 2037 29139 2103 29142
rect 2630 29140 2636 29142
rect 2700 29142 3483 29144
rect 2700 29140 2747 29142
rect 2681 29139 2747 29140
rect 3417 29139 3483 29142
rect 4846 29142 7052 29202
rect 1669 29066 1735 29069
rect 3141 29066 3207 29069
rect 4521 29066 4587 29069
rect 4846 29066 4906 29142
rect 7046 29140 7052 29142
rect 7116 29140 7122 29204
rect 9857 29202 9923 29205
rect 10593 29202 10659 29205
rect 9857 29200 10659 29202
rect 9857 29144 9862 29200
rect 9918 29144 10598 29200
rect 10654 29144 10659 29200
rect 9857 29142 10659 29144
rect 9857 29139 9923 29142
rect 10593 29139 10659 29142
rect 1669 29064 3207 29066
rect 1669 29008 1674 29064
rect 1730 29008 3146 29064
rect 3202 29008 3207 29064
rect 1669 29006 3207 29008
rect 1669 29003 1735 29006
rect 3141 29003 3207 29006
rect 4156 29064 4587 29066
rect 4156 29008 4526 29064
rect 4582 29008 4587 29064
rect 4156 29006 4587 29008
rect 0 28930 400 28960
rect 2313 28930 2379 28933
rect 0 28928 2379 28930
rect 0 28872 2318 28928
rect 2374 28872 2379 28928
rect 0 28870 2379 28872
rect 0 28840 400 28870
rect 2313 28867 2379 28870
rect 2998 28868 3004 28932
rect 3068 28930 3074 28932
rect 4156 28930 4216 29006
rect 4521 29003 4587 29006
rect 4800 29006 4906 29066
rect 6453 29068 6519 29069
rect 6453 29064 6500 29068
rect 6564 29066 6570 29068
rect 8845 29066 8911 29069
rect 12709 29066 12775 29069
rect 6453 29008 6458 29064
rect 3068 28870 4216 28930
rect 4800 28930 4860 29006
rect 6453 29004 6500 29008
rect 6564 29006 6610 29066
rect 8845 29064 12775 29066
rect 8845 29008 8850 29064
rect 8906 29008 12714 29064
rect 12770 29008 12775 29064
rect 8845 29006 12775 29008
rect 6564 29004 6570 29006
rect 6453 29003 6519 29004
rect 8845 29003 8911 29006
rect 12709 29003 12775 29006
rect 5206 28930 5212 28932
rect 4800 28870 5212 28930
rect 3068 28868 3074 28870
rect 5206 28868 5212 28870
rect 5276 28868 5282 28932
rect 6361 28930 6427 28933
rect 7414 28930 7420 28932
rect 6361 28928 7420 28930
rect 6361 28872 6366 28928
rect 6422 28872 7420 28928
rect 6361 28870 7420 28872
rect 6361 28867 6427 28870
rect 7414 28868 7420 28870
rect 7484 28868 7490 28932
rect 7966 28868 7972 28932
rect 8036 28930 8042 28932
rect 9581 28930 9647 28933
rect 8036 28928 9647 28930
rect 8036 28872 9586 28928
rect 9642 28872 9647 28928
rect 8036 28870 9647 28872
rect 8036 28868 8042 28870
rect 9581 28867 9647 28870
rect 4318 28864 4634 28865
rect 4318 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4634 28864
rect 4318 28799 4634 28800
rect 10718 28864 11034 28865
rect 10718 28800 10724 28864
rect 10788 28800 10804 28864
rect 10868 28800 10884 28864
rect 10948 28800 10964 28864
rect 11028 28800 11034 28864
rect 10718 28799 11034 28800
rect 5165 28794 5231 28797
rect 5390 28794 5396 28796
rect 5165 28792 5396 28794
rect 5165 28736 5170 28792
rect 5226 28736 5396 28792
rect 5165 28734 5396 28736
rect 5165 28731 5231 28734
rect 5390 28732 5396 28734
rect 5460 28732 5466 28796
rect 5574 28732 5580 28796
rect 5644 28794 5650 28796
rect 6269 28794 6335 28797
rect 5644 28792 6335 28794
rect 5644 28736 6274 28792
rect 6330 28736 6335 28792
rect 5644 28734 6335 28736
rect 5644 28732 5650 28734
rect 6269 28731 6335 28734
rect 0 28658 400 28688
rect 1025 28658 1091 28661
rect 0 28656 1091 28658
rect 0 28600 1030 28656
rect 1086 28600 1091 28656
rect 0 28598 1091 28600
rect 0 28568 400 28598
rect 1025 28595 1091 28598
rect 3785 28658 3851 28661
rect 7189 28658 7255 28661
rect 3785 28656 7255 28658
rect 3785 28600 3790 28656
rect 3846 28600 7194 28656
rect 7250 28600 7255 28656
rect 3785 28598 7255 28600
rect 3785 28595 3851 28598
rect 7189 28595 7255 28598
rect 8886 28596 8892 28660
rect 8956 28658 8962 28660
rect 12065 28658 12131 28661
rect 8956 28656 12131 28658
rect 8956 28600 12070 28656
rect 12126 28600 12131 28656
rect 8956 28598 12131 28600
rect 8956 28596 8962 28598
rect 12065 28595 12131 28598
rect 1710 28460 1716 28524
rect 1780 28522 1786 28524
rect 3877 28522 3943 28525
rect 1780 28520 3943 28522
rect 1780 28464 3882 28520
rect 3938 28464 3943 28520
rect 1780 28462 3943 28464
rect 1780 28460 1786 28462
rect 3877 28459 3943 28462
rect 4061 28522 4127 28525
rect 4245 28522 4311 28525
rect 4061 28520 4311 28522
rect 4061 28464 4066 28520
rect 4122 28464 4250 28520
rect 4306 28464 4311 28520
rect 4061 28462 4311 28464
rect 4061 28459 4127 28462
rect 4245 28459 4311 28462
rect 9070 28460 9076 28524
rect 9140 28522 9146 28524
rect 11278 28522 11284 28524
rect 9140 28462 11284 28522
rect 9140 28460 9146 28462
rect 11278 28460 11284 28462
rect 11348 28460 11354 28524
rect 0 28386 400 28416
rect 749 28386 815 28389
rect 1025 28386 1091 28389
rect 0 28384 1091 28386
rect 0 28328 754 28384
rect 810 28328 1030 28384
rect 1086 28328 1091 28384
rect 0 28326 1091 28328
rect 0 28296 400 28326
rect 749 28323 815 28326
rect 1025 28323 1091 28326
rect 6269 28386 6335 28389
rect 7046 28386 7052 28388
rect 6269 28384 7052 28386
rect 6269 28328 6274 28384
rect 6330 28328 7052 28384
rect 6269 28326 7052 28328
rect 6269 28323 6335 28326
rect 7046 28324 7052 28326
rect 7116 28324 7122 28388
rect 3658 28320 3974 28321
rect 3658 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3974 28320
rect 3658 28255 3974 28256
rect 10058 28320 10374 28321
rect 10058 28256 10064 28320
rect 10128 28256 10144 28320
rect 10208 28256 10224 28320
rect 10288 28256 10304 28320
rect 10368 28256 10374 28320
rect 10058 28255 10374 28256
rect 606 28188 612 28252
rect 676 28250 682 28252
rect 2773 28250 2839 28253
rect 676 28248 2839 28250
rect 676 28192 2778 28248
rect 2834 28192 2839 28248
rect 676 28190 2839 28192
rect 676 28188 682 28190
rect 2773 28187 2839 28190
rect 4429 28250 4495 28253
rect 8937 28250 9003 28253
rect 4429 28248 9003 28250
rect 4429 28192 4434 28248
rect 4490 28192 8942 28248
rect 8998 28192 9003 28248
rect 4429 28190 9003 28192
rect 4429 28187 4495 28190
rect 8937 28187 9003 28190
rect 0 28114 400 28144
rect 1117 28114 1183 28117
rect 0 28112 1183 28114
rect 0 28056 1122 28112
rect 1178 28056 1183 28112
rect 0 28054 1183 28056
rect 0 28024 400 28054
rect 1117 28051 1183 28054
rect 4429 28114 4495 28117
rect 4797 28114 4863 28117
rect 6678 28114 6684 28116
rect 4429 28112 6684 28114
rect 4429 28056 4434 28112
rect 4490 28056 4802 28112
rect 4858 28056 6684 28112
rect 4429 28054 6684 28056
rect 4429 28051 4495 28054
rect 4797 28051 4863 28054
rect 6678 28052 6684 28054
rect 6748 28052 6754 28116
rect 6862 28052 6868 28116
rect 6932 28114 6938 28116
rect 7097 28114 7163 28117
rect 6932 28112 7163 28114
rect 6932 28056 7102 28112
rect 7158 28056 7163 28112
rect 6932 28054 7163 28056
rect 6932 28052 6938 28054
rect 7097 28051 7163 28054
rect 7782 28052 7788 28116
rect 7852 28114 7858 28116
rect 8385 28114 8451 28117
rect 7852 28112 8451 28114
rect 7852 28056 8390 28112
rect 8446 28056 8451 28112
rect 7852 28054 8451 28056
rect 7852 28052 7858 28054
rect 8385 28051 8451 28054
rect 10225 28114 10291 28117
rect 10501 28114 10567 28117
rect 10225 28112 10567 28114
rect 10225 28056 10230 28112
rect 10286 28056 10506 28112
rect 10562 28056 10567 28112
rect 10225 28054 10567 28056
rect 10225 28051 10291 28054
rect 10501 28051 10567 28054
rect 3049 27978 3115 27981
rect 8150 27978 8156 27980
rect 3049 27976 8156 27978
rect 3049 27920 3054 27976
rect 3110 27920 8156 27976
rect 3049 27918 8156 27920
rect 3049 27915 3115 27918
rect 8150 27916 8156 27918
rect 8220 27916 8226 27980
rect 8518 27916 8524 27980
rect 8588 27978 8594 27980
rect 11094 27978 11100 27980
rect 8588 27918 11100 27978
rect 8588 27916 8594 27918
rect 11094 27916 11100 27918
rect 11164 27916 11170 27980
rect 1710 27780 1716 27844
rect 1780 27842 1786 27844
rect 1945 27842 2011 27845
rect 1780 27840 2011 27842
rect 1780 27784 1950 27840
rect 2006 27784 2011 27840
rect 1780 27782 2011 27784
rect 1780 27780 1786 27782
rect 1945 27779 2011 27782
rect 6637 27842 6703 27845
rect 8334 27842 8340 27844
rect 6637 27840 8340 27842
rect 6637 27784 6642 27840
rect 6698 27784 8340 27840
rect 6637 27782 8340 27784
rect 6637 27779 6703 27782
rect 8334 27780 8340 27782
rect 8404 27780 8410 27844
rect 4318 27776 4634 27777
rect 4318 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4634 27776
rect 4318 27711 4634 27712
rect 10718 27776 11034 27777
rect 10718 27712 10724 27776
rect 10788 27712 10804 27776
rect 10868 27712 10884 27776
rect 10948 27712 10964 27776
rect 11028 27712 11034 27776
rect 10718 27711 11034 27712
rect 197 27706 263 27709
rect 2262 27706 2268 27708
rect 197 27704 2268 27706
rect 197 27648 202 27704
rect 258 27648 2268 27704
rect 197 27646 2268 27648
rect 197 27643 263 27646
rect 2262 27644 2268 27646
rect 2332 27644 2338 27708
rect 2446 27644 2452 27708
rect 2516 27706 2522 27708
rect 2589 27706 2655 27709
rect 2516 27704 2655 27706
rect 2516 27648 2594 27704
rect 2650 27648 2655 27704
rect 2516 27646 2655 27648
rect 2516 27644 2522 27646
rect 2589 27643 2655 27646
rect 6126 27644 6132 27708
rect 6196 27706 6202 27708
rect 6913 27706 6979 27709
rect 6196 27704 6979 27706
rect 6196 27648 6918 27704
rect 6974 27648 6979 27704
rect 6196 27646 6979 27648
rect 6196 27644 6202 27646
rect 6913 27643 6979 27646
rect 11646 27644 11652 27708
rect 11716 27706 11722 27708
rect 12249 27706 12315 27709
rect 11716 27704 12315 27706
rect 11716 27648 12254 27704
rect 12310 27648 12315 27704
rect 11716 27646 12315 27648
rect 11716 27644 11722 27646
rect 12249 27643 12315 27646
rect 6545 27570 6611 27573
rect 7598 27570 7604 27572
rect 6545 27568 7604 27570
rect 6545 27512 6550 27568
rect 6606 27512 7604 27568
rect 6545 27510 7604 27512
rect 6545 27507 6611 27510
rect 7598 27508 7604 27510
rect 7668 27508 7674 27572
rect 8569 27570 8635 27573
rect 8886 27570 8892 27572
rect 8569 27568 8892 27570
rect 8569 27512 8574 27568
rect 8630 27512 8892 27568
rect 8569 27510 8892 27512
rect 8569 27507 8635 27510
rect 8886 27508 8892 27510
rect 8956 27570 8962 27572
rect 9581 27570 9647 27573
rect 8956 27568 9647 27570
rect 8956 27512 9586 27568
rect 9642 27512 9647 27568
rect 8956 27510 9647 27512
rect 8956 27508 8962 27510
rect 9581 27507 9647 27510
rect 5809 27434 5875 27437
rect 6729 27436 6795 27437
rect 6678 27434 6684 27436
rect 5809 27432 6684 27434
rect 6748 27434 6795 27436
rect 9673 27434 9739 27437
rect 10542 27434 10548 27436
rect 6748 27432 6876 27434
rect 5809 27376 5814 27432
rect 5870 27376 6684 27432
rect 6790 27376 6876 27432
rect 5809 27374 6684 27376
rect 5809 27371 5875 27374
rect 6678 27372 6684 27374
rect 6748 27374 6876 27376
rect 9673 27432 10548 27434
rect 9673 27376 9678 27432
rect 9734 27376 10548 27432
rect 9673 27374 10548 27376
rect 6748 27372 6795 27374
rect 6729 27371 6795 27372
rect 9673 27371 9739 27374
rect 10542 27372 10548 27374
rect 10612 27372 10618 27436
rect 6729 27298 6795 27301
rect 7189 27298 7255 27301
rect 6729 27296 7255 27298
rect 6729 27240 6734 27296
rect 6790 27240 7194 27296
rect 7250 27240 7255 27296
rect 6729 27238 7255 27240
rect 6729 27235 6795 27238
rect 7189 27235 7255 27238
rect 3658 27232 3974 27233
rect 3658 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3974 27232
rect 3658 27167 3974 27168
rect 10058 27232 10374 27233
rect 10058 27168 10064 27232
rect 10128 27168 10144 27232
rect 10208 27168 10224 27232
rect 10288 27168 10304 27232
rect 10368 27168 10374 27232
rect 10058 27167 10374 27168
rect 9673 27164 9739 27165
rect 9622 27162 9628 27164
rect 9582 27102 9628 27162
rect 9692 27160 9739 27164
rect 9734 27104 9739 27160
rect 9622 27100 9628 27102
rect 9692 27100 9739 27104
rect 9673 27099 9739 27100
rect 8017 27026 8083 27029
rect 7974 27024 8083 27026
rect 7974 26968 8022 27024
rect 8078 26968 8083 27024
rect 7974 26963 8083 26968
rect 4613 26890 4679 26893
rect 5390 26890 5396 26892
rect 4613 26888 5396 26890
rect 4613 26832 4618 26888
rect 4674 26832 5396 26888
rect 4613 26830 5396 26832
rect 4613 26827 4679 26830
rect 5390 26828 5396 26830
rect 5460 26890 5466 26892
rect 7974 26890 8034 26963
rect 5460 26830 8034 26890
rect 5460 26828 5466 26830
rect 4318 26688 4634 26689
rect 4318 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4634 26688
rect 4318 26623 4634 26624
rect 10718 26688 11034 26689
rect 10718 26624 10724 26688
rect 10788 26624 10804 26688
rect 10868 26624 10884 26688
rect 10948 26624 10964 26688
rect 11028 26624 11034 26688
rect 10718 26623 11034 26624
rect 2129 26620 2195 26621
rect 2078 26618 2084 26620
rect 2038 26558 2084 26618
rect 2148 26616 2195 26620
rect 2190 26560 2195 26616
rect 2078 26556 2084 26558
rect 2148 26556 2195 26560
rect 2129 26555 2195 26556
rect 7373 26618 7439 26621
rect 9121 26618 9187 26621
rect 7373 26616 9187 26618
rect 7373 26560 7378 26616
rect 7434 26560 9126 26616
rect 9182 26560 9187 26616
rect 7373 26558 9187 26560
rect 7373 26555 7439 26558
rect 9121 26555 9187 26558
rect 6177 26482 6243 26485
rect 6545 26482 6611 26485
rect 6177 26480 6611 26482
rect 6177 26424 6182 26480
rect 6238 26424 6550 26480
rect 6606 26424 6611 26480
rect 6177 26422 6611 26424
rect 6177 26419 6243 26422
rect 6545 26419 6611 26422
rect 7046 26420 7052 26484
rect 7116 26482 7122 26484
rect 9622 26482 9628 26484
rect 7116 26422 9628 26482
rect 7116 26420 7122 26422
rect 9622 26420 9628 26422
rect 9692 26420 9698 26484
rect 2037 26348 2103 26349
rect 2037 26344 2084 26348
rect 2148 26346 2154 26348
rect 2037 26288 2042 26344
rect 2037 26284 2084 26288
rect 2148 26286 2194 26346
rect 2405 26344 2471 26349
rect 4061 26346 4127 26349
rect 2405 26288 2410 26344
rect 2466 26288 2471 26344
rect 2148 26284 2154 26286
rect 2037 26283 2103 26284
rect 2405 26283 2471 26288
rect 3512 26344 4127 26346
rect 3512 26288 4066 26344
rect 4122 26288 4127 26344
rect 3512 26286 4127 26288
rect 2408 25941 2468 26283
rect 3512 26213 3572 26286
rect 4061 26283 4127 26286
rect 8150 26284 8156 26348
rect 8220 26346 8226 26348
rect 8220 26286 8448 26346
rect 8220 26284 8226 26286
rect 8388 26213 8448 26286
rect 9806 26284 9812 26348
rect 9876 26346 9882 26348
rect 11421 26346 11487 26349
rect 9876 26344 11487 26346
rect 9876 26288 11426 26344
rect 11482 26288 11487 26344
rect 9876 26286 11487 26288
rect 9876 26284 9882 26286
rect 11421 26283 11487 26286
rect 3509 26208 3575 26213
rect 3509 26152 3514 26208
rect 3570 26152 3575 26208
rect 3509 26147 3575 26152
rect 8385 26208 8451 26213
rect 8385 26152 8390 26208
rect 8446 26152 8451 26208
rect 8385 26147 8451 26152
rect 3658 26144 3974 26145
rect 3658 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3974 26144
rect 3658 26079 3974 26080
rect 10058 26144 10374 26145
rect 10058 26080 10064 26144
rect 10128 26080 10144 26144
rect 10208 26080 10224 26144
rect 10288 26080 10304 26144
rect 10368 26080 10374 26144
rect 10058 26079 10374 26080
rect 6310 26012 6316 26076
rect 6380 26074 6386 26076
rect 9438 26074 9444 26076
rect 6380 26014 9444 26074
rect 6380 26012 6386 26014
rect 9438 26012 9444 26014
rect 9508 26012 9514 26076
rect 2405 25936 2471 25941
rect 2405 25880 2410 25936
rect 2466 25880 2471 25936
rect 2405 25875 2471 25880
rect 3366 25876 3372 25940
rect 3436 25938 3442 25940
rect 3969 25938 4035 25941
rect 3436 25936 4035 25938
rect 3436 25880 3974 25936
rect 4030 25880 4035 25936
rect 3436 25878 4035 25880
rect 3436 25876 3442 25878
rect 3969 25875 4035 25878
rect 4521 25938 4587 25941
rect 8569 25938 8635 25941
rect 4521 25936 8635 25938
rect 4521 25880 4526 25936
rect 4582 25880 8574 25936
rect 8630 25880 8635 25936
rect 4521 25878 8635 25880
rect 4521 25875 4587 25878
rect 8569 25875 8635 25878
rect 3972 25802 4032 25875
rect 5625 25802 5691 25805
rect 8017 25802 8083 25805
rect 3972 25800 8083 25802
rect 3972 25744 5630 25800
rect 5686 25744 8022 25800
rect 8078 25744 8083 25800
rect 3972 25742 8083 25744
rect 5625 25739 5691 25742
rect 8017 25739 8083 25742
rect 7005 25668 7071 25669
rect 7005 25666 7052 25668
rect 6960 25664 7052 25666
rect 6960 25608 7010 25664
rect 6960 25606 7052 25608
rect 7005 25604 7052 25606
rect 7116 25604 7122 25668
rect 7005 25603 7071 25604
rect 4318 25600 4634 25601
rect 4318 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4634 25600
rect 4318 25535 4634 25536
rect 10718 25600 11034 25601
rect 10718 25536 10724 25600
rect 10788 25536 10804 25600
rect 10868 25536 10884 25600
rect 10948 25536 10964 25600
rect 11028 25536 11034 25600
rect 10718 25535 11034 25536
rect 2446 25468 2452 25532
rect 2516 25530 2522 25532
rect 2865 25530 2931 25533
rect 2516 25528 2931 25530
rect 2516 25472 2870 25528
rect 2926 25472 2931 25528
rect 2516 25470 2931 25472
rect 2516 25468 2522 25470
rect 2865 25467 2931 25470
rect 1158 25332 1164 25396
rect 1228 25394 1234 25396
rect 5574 25394 5580 25396
rect 1228 25334 5580 25394
rect 1228 25332 1234 25334
rect 5574 25332 5580 25334
rect 5644 25332 5650 25396
rect 6637 25394 6703 25397
rect 8109 25394 8175 25397
rect 6637 25392 8175 25394
rect 6637 25336 6642 25392
rect 6698 25336 8114 25392
rect 8170 25336 8175 25392
rect 6637 25334 8175 25336
rect 6637 25331 6703 25334
rect 8109 25331 8175 25334
rect 4838 25258 4844 25260
rect 3006 25198 4844 25258
rect 565 25122 631 25125
rect 3006 25122 3066 25198
rect 4838 25196 4844 25198
rect 4908 25196 4914 25260
rect 565 25120 3066 25122
rect 565 25064 570 25120
rect 626 25064 3066 25120
rect 565 25062 3066 25064
rect 5257 25122 5323 25125
rect 8569 25122 8635 25125
rect 5257 25120 8635 25122
rect 5257 25064 5262 25120
rect 5318 25064 8574 25120
rect 8630 25064 8635 25120
rect 5257 25062 8635 25064
rect 565 25059 631 25062
rect 5257 25059 5323 25062
rect 8569 25059 8635 25062
rect 3658 25056 3974 25057
rect 3658 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3974 25056
rect 3658 24991 3974 24992
rect 10058 25056 10374 25057
rect 10058 24992 10064 25056
rect 10128 24992 10144 25056
rect 10208 24992 10224 25056
rect 10288 24992 10304 25056
rect 10368 24992 10374 25056
rect 10058 24991 10374 24992
rect 4797 24986 4863 24989
rect 5758 24986 5764 24988
rect 4797 24984 5764 24986
rect 4797 24928 4802 24984
rect 4858 24928 5764 24984
rect 4797 24926 5764 24928
rect 4797 24923 4863 24926
rect 5758 24924 5764 24926
rect 5828 24924 5834 24988
rect 11830 24986 11836 24988
rect 10550 24926 11836 24986
rect 1761 24848 1827 24853
rect 1761 24792 1766 24848
rect 1822 24792 1827 24848
rect 1761 24787 1827 24792
rect 5809 24850 5875 24853
rect 7097 24850 7163 24853
rect 5809 24848 7163 24850
rect 5809 24792 5814 24848
rect 5870 24792 7102 24848
rect 7158 24792 7163 24848
rect 5809 24790 7163 24792
rect 5809 24787 5875 24790
rect 7097 24787 7163 24790
rect 0 24306 400 24336
rect 749 24306 815 24309
rect 0 24304 815 24306
rect 0 24248 754 24304
rect 810 24248 815 24304
rect 0 24246 815 24248
rect 1764 24306 1824 24787
rect 2221 24714 2287 24717
rect 5809 24714 5875 24717
rect 8753 24714 8819 24717
rect 2221 24712 2330 24714
rect 2221 24656 2226 24712
rect 2282 24656 2330 24712
rect 2221 24651 2330 24656
rect 5809 24712 8819 24714
rect 5809 24656 5814 24712
rect 5870 24656 8758 24712
rect 8814 24656 8819 24712
rect 5809 24654 8819 24656
rect 5809 24651 5875 24654
rect 8753 24651 8819 24654
rect 9121 24714 9187 24717
rect 9254 24714 9260 24716
rect 9121 24712 9260 24714
rect 9121 24656 9126 24712
rect 9182 24656 9260 24712
rect 9121 24654 9260 24656
rect 9121 24651 9187 24654
rect 9254 24652 9260 24654
rect 9324 24652 9330 24716
rect 2270 24578 2330 24651
rect 5717 24580 5783 24581
rect 3366 24578 3372 24580
rect 2270 24518 3372 24578
rect 3366 24516 3372 24518
rect 3436 24516 3442 24580
rect 5717 24576 5764 24580
rect 5828 24578 5834 24580
rect 6269 24578 6335 24581
rect 7189 24578 7255 24581
rect 5717 24520 5722 24576
rect 5717 24516 5764 24520
rect 5828 24518 5874 24578
rect 6269 24576 7255 24578
rect 6269 24520 6274 24576
rect 6330 24520 7194 24576
rect 7250 24520 7255 24576
rect 6269 24518 7255 24520
rect 5828 24516 5834 24518
rect 5717 24515 5783 24516
rect 6269 24515 6335 24518
rect 7189 24515 7255 24518
rect 8569 24578 8635 24581
rect 9070 24578 9076 24580
rect 8569 24576 9076 24578
rect 8569 24520 8574 24576
rect 8630 24520 9076 24576
rect 8569 24518 9076 24520
rect 8569 24515 8635 24518
rect 9070 24516 9076 24518
rect 9140 24516 9146 24580
rect 9765 24578 9831 24581
rect 10550 24578 10610 24926
rect 11830 24924 11836 24926
rect 11900 24924 11906 24988
rect 9765 24576 10610 24578
rect 9765 24520 9770 24576
rect 9826 24520 10610 24576
rect 9765 24518 10610 24520
rect 9765 24515 9831 24518
rect 4318 24512 4634 24513
rect 4318 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4634 24512
rect 4318 24447 4634 24448
rect 10718 24512 11034 24513
rect 10718 24448 10724 24512
rect 10788 24448 10804 24512
rect 10868 24448 10884 24512
rect 10948 24448 10964 24512
rect 11028 24448 11034 24512
rect 10718 24447 11034 24448
rect 5349 24442 5415 24445
rect 6269 24442 6335 24445
rect 6637 24442 6703 24445
rect 5349 24440 6703 24442
rect 5349 24384 5354 24440
rect 5410 24384 6274 24440
rect 6330 24384 6642 24440
rect 6698 24384 6703 24440
rect 5349 24382 6703 24384
rect 5349 24379 5415 24382
rect 6269 24379 6335 24382
rect 6637 24379 6703 24382
rect 2037 24306 2103 24309
rect 1764 24304 2103 24306
rect 1764 24248 2042 24304
rect 2098 24248 2103 24304
rect 1764 24246 2103 24248
rect 0 24216 400 24246
rect 749 24243 815 24246
rect 2037 24243 2103 24246
rect 3693 24306 3759 24309
rect 6361 24306 6427 24309
rect 3693 24304 6427 24306
rect 3693 24248 3698 24304
rect 3754 24248 6366 24304
rect 6422 24248 6427 24304
rect 3693 24246 6427 24248
rect 3693 24243 3759 24246
rect 6361 24243 6427 24246
rect 1894 24108 1900 24172
rect 1964 24170 1970 24172
rect 4061 24170 4127 24173
rect 1964 24168 4127 24170
rect 1964 24112 4066 24168
rect 4122 24112 4127 24168
rect 1964 24110 4127 24112
rect 1964 24108 1970 24110
rect 4061 24107 4127 24110
rect 6269 24170 6335 24173
rect 6729 24170 6795 24173
rect 6269 24168 6795 24170
rect 6269 24112 6274 24168
rect 6330 24112 6734 24168
rect 6790 24112 6795 24168
rect 6269 24110 6795 24112
rect 6269 24107 6335 24110
rect 6729 24107 6795 24110
rect 7281 24170 7347 24173
rect 7925 24170 7991 24173
rect 7281 24168 7991 24170
rect 7281 24112 7286 24168
rect 7342 24112 7930 24168
rect 7986 24112 7991 24168
rect 7281 24110 7991 24112
rect 7281 24107 7347 24110
rect 7925 24107 7991 24110
rect 8293 24170 8359 24173
rect 9029 24170 9095 24173
rect 8293 24168 9095 24170
rect 8293 24112 8298 24168
rect 8354 24112 9034 24168
rect 9090 24112 9095 24168
rect 8293 24110 9095 24112
rect 8293 24107 8359 24110
rect 9029 24107 9095 24110
rect 0 24034 400 24064
rect 1025 24034 1091 24037
rect 0 24032 1091 24034
rect 0 23976 1030 24032
rect 1086 23976 1091 24032
rect 0 23974 1091 23976
rect 0 23944 400 23974
rect 1025 23971 1091 23974
rect 3658 23968 3974 23969
rect 3658 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3974 23968
rect 3658 23903 3974 23904
rect 10058 23968 10374 23969
rect 10058 23904 10064 23968
rect 10128 23904 10144 23968
rect 10208 23904 10224 23968
rect 10288 23904 10304 23968
rect 10368 23904 10374 23968
rect 10058 23903 10374 23904
rect 1342 23836 1348 23900
rect 1412 23898 1418 23900
rect 2957 23898 3023 23901
rect 1412 23896 3023 23898
rect 1412 23840 2962 23896
rect 3018 23840 3023 23896
rect 1412 23838 3023 23840
rect 1412 23836 1418 23838
rect 2957 23835 3023 23838
rect 0 23762 400 23792
rect 473 23762 539 23765
rect 0 23760 539 23762
rect 0 23704 478 23760
rect 534 23704 539 23760
rect 0 23702 539 23704
rect 0 23672 400 23702
rect 473 23699 539 23702
rect 2630 23700 2636 23764
rect 2700 23762 2706 23764
rect 4102 23762 4108 23764
rect 2700 23702 4108 23762
rect 2700 23700 2706 23702
rect 4102 23700 4108 23702
rect 4172 23700 4178 23764
rect 6729 23762 6795 23765
rect 6862 23762 6868 23764
rect 6729 23760 6868 23762
rect 6729 23704 6734 23760
rect 6790 23704 6868 23760
rect 6729 23702 6868 23704
rect 6729 23699 6795 23702
rect 6862 23700 6868 23702
rect 6932 23700 6938 23764
rect 7414 23700 7420 23764
rect 7484 23762 7490 23764
rect 7649 23762 7715 23765
rect 7484 23760 7715 23762
rect 7484 23704 7654 23760
rect 7710 23704 7715 23760
rect 7484 23702 7715 23704
rect 7484 23700 7490 23702
rect 7649 23699 7715 23702
rect 3141 23626 3207 23629
rect 4102 23626 4108 23628
rect 3141 23624 4108 23626
rect 3141 23568 3146 23624
rect 3202 23568 4108 23624
rect 3141 23566 4108 23568
rect 3141 23563 3207 23566
rect 4102 23564 4108 23566
rect 4172 23564 4178 23628
rect 9765 23626 9831 23629
rect 7790 23624 9831 23626
rect 7790 23568 9770 23624
rect 9826 23568 9831 23624
rect 7790 23566 9831 23568
rect 0 23490 400 23520
rect 1301 23490 1367 23493
rect 0 23488 1367 23490
rect 0 23432 1306 23488
rect 1362 23432 1367 23488
rect 0 23430 1367 23432
rect 0 23400 400 23430
rect 1301 23427 1367 23430
rect 2313 23490 2379 23493
rect 3049 23490 3115 23493
rect 2313 23488 3115 23490
rect 2313 23432 2318 23488
rect 2374 23432 3054 23488
rect 3110 23432 3115 23488
rect 2313 23430 3115 23432
rect 2313 23427 2379 23430
rect 3049 23427 3115 23430
rect 6678 23428 6684 23492
rect 6748 23490 6754 23492
rect 7790 23490 7850 23566
rect 9765 23563 9831 23566
rect 6748 23430 7850 23490
rect 8201 23490 8267 23493
rect 9673 23490 9739 23493
rect 8201 23488 9739 23490
rect 8201 23432 8206 23488
rect 8262 23432 9678 23488
rect 9734 23432 9739 23488
rect 8201 23430 9739 23432
rect 6748 23428 6754 23430
rect 8201 23427 8267 23430
rect 9673 23427 9739 23430
rect 11421 23492 11487 23493
rect 11421 23488 11468 23492
rect 11532 23490 11538 23492
rect 11697 23490 11763 23493
rect 11830 23490 11836 23492
rect 11421 23432 11426 23488
rect 11421 23428 11468 23432
rect 11532 23430 11578 23490
rect 11697 23488 11836 23490
rect 11697 23432 11702 23488
rect 11758 23432 11836 23488
rect 11697 23430 11836 23432
rect 11532 23428 11538 23430
rect 11421 23427 11487 23428
rect 11697 23427 11763 23430
rect 11830 23428 11836 23430
rect 11900 23428 11906 23492
rect 12014 23428 12020 23492
rect 12084 23490 12090 23492
rect 12709 23490 12775 23493
rect 12084 23488 12775 23490
rect 12084 23432 12714 23488
rect 12770 23432 12775 23488
rect 12084 23430 12775 23432
rect 12084 23428 12090 23430
rect 12709 23427 12775 23430
rect 4318 23424 4634 23425
rect 4318 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4634 23424
rect 4318 23359 4634 23360
rect 10718 23424 11034 23425
rect 10718 23360 10724 23424
rect 10788 23360 10804 23424
rect 10868 23360 10884 23424
rect 10948 23360 10964 23424
rect 11028 23360 11034 23424
rect 10718 23359 11034 23360
rect 2313 23356 2379 23357
rect 2262 23292 2268 23356
rect 2332 23354 2379 23356
rect 6085 23354 6151 23357
rect 7966 23354 7972 23356
rect 2332 23352 2424 23354
rect 2374 23296 2424 23352
rect 2332 23294 2424 23296
rect 6085 23352 7972 23354
rect 6085 23296 6090 23352
rect 6146 23296 7972 23352
rect 6085 23294 7972 23296
rect 2332 23292 2379 23294
rect 2313 23291 2379 23292
rect 6085 23291 6151 23294
rect 7966 23292 7972 23294
rect 8036 23292 8042 23356
rect 0 23218 400 23248
rect 2681 23218 2747 23221
rect 0 23216 2747 23218
rect 0 23160 2686 23216
rect 2742 23160 2747 23216
rect 0 23158 2747 23160
rect 0 23128 400 23158
rect 2681 23155 2747 23158
rect 4429 23218 4495 23221
rect 6913 23218 6979 23221
rect 4429 23216 6979 23218
rect 4429 23160 4434 23216
rect 4490 23160 6918 23216
rect 6974 23160 6979 23216
rect 4429 23158 6979 23160
rect 4429 23155 4495 23158
rect 6913 23155 6979 23158
rect 3182 23020 3188 23084
rect 3252 23082 3258 23084
rect 4613 23082 4679 23085
rect 3252 23080 4679 23082
rect 3252 23024 4618 23080
rect 4674 23024 4679 23080
rect 3252 23022 4679 23024
rect 3252 23020 3258 23022
rect 4613 23019 4679 23022
rect 6361 23082 6427 23085
rect 6821 23082 6887 23085
rect 7966 23082 7972 23084
rect 6361 23080 7972 23082
rect 6361 23024 6366 23080
rect 6422 23024 6826 23080
rect 6882 23024 7972 23080
rect 6361 23022 7972 23024
rect 6361 23019 6427 23022
rect 6821 23019 6887 23022
rect 7966 23020 7972 23022
rect 8036 23020 8042 23084
rect 10409 23082 10475 23085
rect 12341 23082 12407 23085
rect 12566 23082 12572 23084
rect 10409 23080 10610 23082
rect 10409 23024 10414 23080
rect 10470 23024 10610 23080
rect 10409 23022 10610 23024
rect 10409 23019 10475 23022
rect 0 22946 400 22976
rect 2773 22946 2839 22949
rect 0 22944 2839 22946
rect 0 22888 2778 22944
rect 2834 22888 2839 22944
rect 0 22886 2839 22888
rect 0 22856 400 22886
rect 2773 22883 2839 22886
rect 4061 22946 4127 22949
rect 4889 22946 4955 22949
rect 8385 22946 8451 22949
rect 4061 22944 8451 22946
rect 4061 22888 4066 22944
rect 4122 22888 4894 22944
rect 4950 22888 8390 22944
rect 8446 22888 8451 22944
rect 4061 22886 8451 22888
rect 4061 22883 4127 22886
rect 4889 22883 4955 22886
rect 8385 22883 8451 22886
rect 3658 22880 3974 22881
rect 3658 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3974 22880
rect 3658 22815 3974 22816
rect 10058 22880 10374 22881
rect 10058 22816 10064 22880
rect 10128 22816 10144 22880
rect 10208 22816 10224 22880
rect 10288 22816 10304 22880
rect 10368 22816 10374 22880
rect 10058 22815 10374 22816
rect 4838 22748 4844 22812
rect 4908 22810 4914 22812
rect 5073 22810 5139 22813
rect 4908 22808 5139 22810
rect 4908 22752 5078 22808
rect 5134 22752 5139 22808
rect 4908 22750 5139 22752
rect 4908 22748 4914 22750
rect 5073 22747 5139 22750
rect 0 22674 400 22704
rect 1025 22674 1091 22677
rect 0 22672 1091 22674
rect 0 22616 1030 22672
rect 1086 22616 1091 22672
rect 0 22614 1091 22616
rect 0 22584 400 22614
rect 1025 22611 1091 22614
rect 2865 22674 2931 22677
rect 2998 22674 3004 22676
rect 2865 22672 3004 22674
rect 2865 22616 2870 22672
rect 2926 22616 3004 22672
rect 2865 22614 3004 22616
rect 2865 22611 2931 22614
rect 2998 22612 3004 22614
rect 3068 22612 3074 22676
rect 4245 22674 4311 22677
rect 8937 22674 9003 22677
rect 4245 22672 9003 22674
rect 4245 22616 4250 22672
rect 4306 22616 8942 22672
rect 8998 22616 9003 22672
rect 4245 22614 9003 22616
rect 4245 22611 4311 22614
rect 8937 22611 9003 22614
rect 9438 22612 9444 22676
rect 9508 22674 9514 22676
rect 9949 22674 10015 22677
rect 9508 22672 10015 22674
rect 9508 22616 9954 22672
rect 10010 22616 10015 22672
rect 9508 22614 10015 22616
rect 9508 22612 9514 22614
rect 9949 22611 10015 22614
rect 10133 22674 10199 22677
rect 10550 22674 10610 23022
rect 12341 23080 12572 23082
rect 12341 23024 12346 23080
rect 12402 23024 12572 23080
rect 12341 23022 12572 23024
rect 12341 23019 12407 23022
rect 12566 23020 12572 23022
rect 12636 23020 12642 23084
rect 10133 22672 10610 22674
rect 10133 22616 10138 22672
rect 10194 22616 10610 22672
rect 10133 22614 10610 22616
rect 10133 22611 10199 22614
rect 5022 22538 5028 22540
rect 2638 22478 5028 22538
rect 2313 22130 2379 22133
rect 2270 22128 2379 22130
rect 2270 22072 2318 22128
rect 2374 22072 2379 22128
rect 2270 22067 2379 22072
rect 381 21994 447 21997
rect 2270 21994 2330 22067
rect 381 21992 2330 21994
rect 381 21936 386 21992
rect 442 21936 2330 21992
rect 381 21934 2330 21936
rect 2405 21994 2471 21997
rect 2638 21994 2698 22478
rect 5022 22476 5028 22478
rect 5092 22476 5098 22540
rect 10777 22538 10843 22541
rect 12065 22538 12131 22541
rect 10777 22536 12131 22538
rect 10777 22480 10782 22536
rect 10838 22480 12070 22536
rect 12126 22480 12131 22536
rect 10777 22478 12131 22480
rect 10777 22475 10843 22478
rect 12065 22475 12131 22478
rect 4318 22336 4634 22337
rect 4318 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4634 22336
rect 4318 22271 4634 22272
rect 10718 22336 11034 22337
rect 10718 22272 10724 22336
rect 10788 22272 10804 22336
rect 10868 22272 10884 22336
rect 10948 22272 10964 22336
rect 11028 22272 11034 22336
rect 10718 22271 11034 22272
rect 4981 22268 5047 22269
rect 4981 22264 5028 22268
rect 5092 22266 5098 22268
rect 5349 22266 5415 22269
rect 6085 22266 6151 22269
rect 4981 22208 4986 22264
rect 4981 22204 5028 22208
rect 5092 22206 5138 22266
rect 5349 22264 6151 22266
rect 5349 22208 5354 22264
rect 5410 22208 6090 22264
rect 6146 22208 6151 22264
rect 5349 22206 6151 22208
rect 5092 22204 5098 22206
rect 4981 22203 5047 22204
rect 5349 22203 5415 22206
rect 6085 22203 6151 22206
rect 6729 22266 6795 22269
rect 7414 22266 7420 22268
rect 6729 22264 7420 22266
rect 6729 22208 6734 22264
rect 6790 22208 7420 22264
rect 6729 22206 7420 22208
rect 6729 22203 6795 22206
rect 7414 22204 7420 22206
rect 7484 22204 7490 22268
rect 8477 22266 8543 22269
rect 8342 22264 8543 22266
rect 8342 22208 8482 22264
rect 8538 22208 8543 22264
rect 8342 22206 8543 22208
rect 8342 22133 8402 22206
rect 8477 22203 8543 22206
rect 2814 22068 2820 22132
rect 2884 22130 2890 22132
rect 3233 22130 3299 22133
rect 2884 22128 3299 22130
rect 2884 22072 3238 22128
rect 3294 22072 3299 22128
rect 2884 22070 3299 22072
rect 2884 22068 2890 22070
rect 3233 22067 3299 22070
rect 4102 22068 4108 22132
rect 4172 22130 4178 22132
rect 4337 22130 4403 22133
rect 7281 22130 7347 22133
rect 8109 22130 8175 22133
rect 4172 22128 4403 22130
rect 4172 22072 4342 22128
rect 4398 22072 4403 22128
rect 4172 22070 4403 22072
rect 4172 22068 4178 22070
rect 4337 22067 4403 22070
rect 5720 22128 8175 22130
rect 5720 22072 7286 22128
rect 7342 22072 8114 22128
rect 8170 22072 8175 22128
rect 5720 22070 8175 22072
rect 8342 22128 8451 22133
rect 8342 22072 8390 22128
rect 8446 22072 8451 22128
rect 8342 22070 8451 22072
rect 5720 21997 5780 22070
rect 7281 22067 7347 22070
rect 8109 22067 8175 22070
rect 8385 22067 8451 22070
rect 11053 22130 11119 22133
rect 11605 22130 11671 22133
rect 11053 22128 11671 22130
rect 11053 22072 11058 22128
rect 11114 22072 11610 22128
rect 11666 22072 11671 22128
rect 11053 22070 11671 22072
rect 11053 22067 11119 22070
rect 11605 22067 11671 22070
rect 3417 21994 3483 21997
rect 4981 21994 5047 21997
rect 2405 21992 2698 21994
rect 2405 21936 2410 21992
rect 2466 21936 2698 21992
rect 2405 21934 2698 21936
rect 2776 21992 5047 21994
rect 2776 21936 3422 21992
rect 3478 21936 4986 21992
rect 5042 21936 5047 21992
rect 2776 21934 5047 21936
rect 381 21931 447 21934
rect 2405 21931 2471 21934
rect 1761 21858 1827 21861
rect 2776 21858 2836 21934
rect 3417 21931 3483 21934
rect 4981 21931 5047 21934
rect 5717 21992 5783 21997
rect 5717 21936 5722 21992
rect 5778 21936 5783 21992
rect 5717 21931 5783 21936
rect 6729 21994 6795 21997
rect 6862 21994 6868 21996
rect 6729 21992 6868 21994
rect 6729 21936 6734 21992
rect 6790 21936 6868 21992
rect 6729 21934 6868 21936
rect 6729 21931 6795 21934
rect 6862 21932 6868 21934
rect 6932 21932 6938 21996
rect 8334 21932 8340 21996
rect 8404 21994 8410 21996
rect 9806 21994 9812 21996
rect 8404 21934 9812 21994
rect 8404 21932 8410 21934
rect 9806 21932 9812 21934
rect 9876 21932 9882 21996
rect 1761 21856 2836 21858
rect 1761 21800 1766 21856
rect 1822 21800 2836 21856
rect 1761 21798 2836 21800
rect 4889 21858 4955 21861
rect 5625 21858 5691 21861
rect 4889 21856 5691 21858
rect 4889 21800 4894 21856
rect 4950 21800 5630 21856
rect 5686 21800 5691 21856
rect 4889 21798 5691 21800
rect 1761 21795 1827 21798
rect 4889 21795 4955 21798
rect 5625 21795 5691 21798
rect 5809 21858 5875 21861
rect 5942 21858 5948 21860
rect 5809 21856 5948 21858
rect 5809 21800 5814 21856
rect 5870 21800 5948 21856
rect 5809 21798 5948 21800
rect 5809 21795 5875 21798
rect 5942 21796 5948 21798
rect 6012 21796 6018 21860
rect 7966 21796 7972 21860
rect 8036 21858 8042 21860
rect 9213 21858 9279 21861
rect 8036 21856 9279 21858
rect 8036 21800 9218 21856
rect 9274 21800 9279 21856
rect 8036 21798 9279 21800
rect 8036 21796 8042 21798
rect 9213 21795 9279 21798
rect 3658 21792 3974 21793
rect 3658 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3974 21792
rect 3658 21727 3974 21728
rect 10058 21792 10374 21793
rect 10058 21728 10064 21792
rect 10128 21728 10144 21792
rect 10208 21728 10224 21792
rect 10288 21728 10304 21792
rect 10368 21728 10374 21792
rect 10058 21727 10374 21728
rect 4705 21722 4771 21725
rect 5349 21722 5415 21725
rect 4705 21720 5415 21722
rect 4705 21664 4710 21720
rect 4766 21664 5354 21720
rect 5410 21664 5415 21720
rect 4705 21662 5415 21664
rect 4705 21659 4771 21662
rect 5349 21659 5415 21662
rect 2957 21586 3023 21589
rect 3182 21586 3188 21588
rect 2957 21584 3188 21586
rect 2957 21528 2962 21584
rect 3018 21528 3188 21584
rect 2957 21526 3188 21528
rect 2957 21523 3023 21526
rect 3182 21524 3188 21526
rect 3252 21524 3258 21588
rect 3601 21586 3667 21589
rect 4705 21586 4771 21589
rect 3601 21584 4771 21586
rect 3601 21528 3606 21584
rect 3662 21528 4710 21584
rect 4766 21528 4771 21584
rect 3601 21526 4771 21528
rect 3601 21523 3667 21526
rect 4705 21523 4771 21526
rect 6545 21586 6611 21589
rect 8109 21586 8175 21589
rect 6545 21584 8175 21586
rect 6545 21528 6550 21584
rect 6606 21528 8114 21584
rect 8170 21528 8175 21584
rect 6545 21526 8175 21528
rect 6545 21523 6611 21526
rect 8109 21523 8175 21526
rect 2037 21450 2103 21453
rect 2998 21450 3004 21452
rect 2037 21448 3004 21450
rect 2037 21392 2042 21448
rect 2098 21392 3004 21448
rect 2037 21390 3004 21392
rect 2037 21387 2103 21390
rect 2998 21388 3004 21390
rect 3068 21388 3074 21452
rect 3141 21450 3207 21453
rect 3785 21450 3851 21453
rect 4245 21450 4311 21453
rect 3141 21448 3851 21450
rect 3141 21392 3146 21448
rect 3202 21392 3790 21448
rect 3846 21392 3851 21448
rect 3141 21390 3851 21392
rect 3141 21387 3207 21390
rect 3785 21387 3851 21390
rect 4110 21448 4311 21450
rect 4110 21392 4250 21448
rect 4306 21392 4311 21448
rect 4110 21390 4311 21392
rect 1669 21314 1735 21317
rect 3693 21314 3759 21317
rect 1669 21312 3759 21314
rect 1669 21256 1674 21312
rect 1730 21256 3698 21312
rect 3754 21256 3759 21312
rect 1669 21254 3759 21256
rect 1669 21251 1735 21254
rect 3693 21251 3759 21254
rect 2589 21178 2655 21181
rect 3182 21178 3188 21180
rect 2589 21176 3188 21178
rect 2589 21120 2594 21176
rect 2650 21120 3188 21176
rect 2589 21118 3188 21120
rect 2589 21115 2655 21118
rect 3182 21116 3188 21118
rect 3252 21116 3258 21180
rect 2037 21042 2103 21045
rect 3049 21042 3115 21045
rect 3325 21042 3391 21045
rect 3693 21042 3759 21045
rect 2037 21040 3759 21042
rect 2037 20984 2042 21040
rect 2098 20984 3054 21040
rect 3110 20984 3330 21040
rect 3386 20984 3698 21040
rect 3754 20984 3759 21040
rect 2037 20982 3759 20984
rect 4110 21042 4170 21390
rect 4245 21387 4311 21390
rect 5390 21388 5396 21452
rect 5460 21450 5466 21452
rect 5993 21450 6059 21453
rect 5460 21448 6059 21450
rect 5460 21392 5998 21448
rect 6054 21392 6059 21448
rect 5460 21390 6059 21392
rect 5460 21388 5466 21390
rect 5993 21387 6059 21390
rect 5533 21314 5599 21317
rect 7465 21314 7531 21317
rect 5533 21312 7531 21314
rect 5533 21256 5538 21312
rect 5594 21256 7470 21312
rect 7526 21256 7531 21312
rect 5533 21254 7531 21256
rect 5533 21251 5599 21254
rect 7465 21251 7531 21254
rect 10409 21314 10475 21317
rect 10542 21314 10548 21316
rect 10409 21312 10548 21314
rect 10409 21256 10414 21312
rect 10470 21256 10548 21312
rect 10409 21254 10548 21256
rect 10409 21251 10475 21254
rect 10542 21252 10548 21254
rect 10612 21252 10618 21316
rect 4318 21248 4634 21249
rect 4318 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4634 21248
rect 4318 21183 4634 21184
rect 10718 21248 11034 21249
rect 10718 21184 10724 21248
rect 10788 21184 10804 21248
rect 10868 21184 10884 21248
rect 10948 21184 10964 21248
rect 11028 21184 11034 21248
rect 10718 21183 11034 21184
rect 4245 21042 4311 21045
rect 4110 21040 4311 21042
rect 4110 20984 4250 21040
rect 4306 20984 4311 21040
rect 4110 20982 4311 20984
rect 2037 20979 2103 20982
rect 3049 20979 3115 20982
rect 3325 20979 3391 20982
rect 3693 20979 3759 20982
rect 4245 20979 4311 20982
rect 4429 21042 4495 21045
rect 5206 21042 5212 21044
rect 4429 21040 5212 21042
rect 4429 20984 4434 21040
rect 4490 20984 5212 21040
rect 4429 20982 5212 20984
rect 4429 20979 4495 20982
rect 5206 20980 5212 20982
rect 5276 20980 5282 21044
rect 5349 21042 5415 21045
rect 9029 21042 9095 21045
rect 5349 21040 9095 21042
rect 5349 20984 5354 21040
rect 5410 20984 9034 21040
rect 9090 20984 9095 21040
rect 5349 20982 9095 20984
rect 5349 20979 5415 20982
rect 9029 20979 9095 20982
rect 1117 20906 1183 20909
rect 1945 20906 2011 20909
rect 1117 20904 2011 20906
rect 1117 20848 1122 20904
rect 1178 20848 1950 20904
rect 2006 20848 2011 20904
rect 1117 20846 2011 20848
rect 1117 20843 1183 20846
rect 1945 20843 2011 20846
rect 3325 20906 3391 20909
rect 5349 20906 5415 20909
rect 3325 20904 5415 20906
rect 3325 20848 3330 20904
rect 3386 20848 5354 20904
rect 5410 20848 5415 20904
rect 3325 20846 5415 20848
rect 3325 20843 3391 20846
rect 5349 20843 5415 20846
rect 7373 20906 7439 20909
rect 7782 20906 7788 20908
rect 7373 20904 7788 20906
rect 7373 20848 7378 20904
rect 7434 20848 7788 20904
rect 7373 20846 7788 20848
rect 7373 20843 7439 20846
rect 7782 20844 7788 20846
rect 7852 20906 7858 20908
rect 10685 20906 10751 20909
rect 7852 20904 10751 20906
rect 7852 20848 10690 20904
rect 10746 20848 10751 20904
rect 7852 20846 10751 20848
rect 7852 20844 7858 20846
rect 10685 20843 10751 20846
rect 790 20708 796 20772
rect 860 20770 866 20772
rect 860 20710 2790 20770
rect 860 20708 866 20710
rect 1117 20634 1183 20637
rect 1342 20634 1348 20636
rect 1117 20632 1348 20634
rect 1117 20576 1122 20632
rect 1178 20576 1348 20632
rect 1117 20574 1348 20576
rect 1117 20571 1183 20574
rect 1342 20572 1348 20574
rect 1412 20572 1418 20636
rect 1669 20634 1735 20637
rect 2589 20634 2655 20637
rect 1669 20632 2655 20634
rect 1669 20576 1674 20632
rect 1730 20576 2594 20632
rect 2650 20576 2655 20632
rect 1669 20574 2655 20576
rect 1669 20571 1735 20574
rect 2589 20571 2655 20574
rect 2730 20498 2790 20710
rect 5206 20708 5212 20772
rect 5276 20770 5282 20772
rect 5574 20770 5580 20772
rect 5276 20710 5580 20770
rect 5276 20708 5282 20710
rect 5574 20708 5580 20710
rect 5644 20708 5650 20772
rect 7189 20770 7255 20773
rect 7782 20770 7788 20772
rect 7189 20768 7788 20770
rect 7189 20712 7194 20768
rect 7250 20712 7788 20768
rect 7189 20710 7788 20712
rect 7189 20707 7255 20710
rect 7782 20708 7788 20710
rect 7852 20708 7858 20772
rect 9489 20770 9555 20773
rect 9622 20770 9628 20772
rect 9489 20768 9628 20770
rect 9489 20712 9494 20768
rect 9550 20712 9628 20768
rect 9489 20710 9628 20712
rect 9489 20707 9555 20710
rect 9622 20708 9628 20710
rect 9692 20708 9698 20772
rect 3658 20704 3974 20705
rect 3658 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3974 20704
rect 3658 20639 3974 20640
rect 10058 20704 10374 20705
rect 10058 20640 10064 20704
rect 10128 20640 10144 20704
rect 10208 20640 10224 20704
rect 10288 20640 10304 20704
rect 10368 20640 10374 20704
rect 10058 20639 10374 20640
rect 4061 20636 4127 20637
rect 4061 20632 4108 20636
rect 4172 20634 4178 20636
rect 5073 20634 5139 20637
rect 5574 20634 5580 20636
rect 4061 20576 4066 20632
rect 4061 20572 4108 20576
rect 4172 20574 4218 20634
rect 5073 20632 5580 20634
rect 5073 20576 5078 20632
rect 5134 20576 5580 20632
rect 5073 20574 5580 20576
rect 4172 20572 4178 20574
rect 4061 20571 4127 20572
rect 5073 20571 5139 20574
rect 5574 20572 5580 20574
rect 5644 20572 5650 20636
rect 7373 20634 7439 20637
rect 8293 20634 8359 20637
rect 7373 20632 8359 20634
rect 7373 20576 7378 20632
rect 7434 20576 8298 20632
rect 8354 20576 8359 20632
rect 7373 20574 8359 20576
rect 7373 20571 7439 20574
rect 8293 20571 8359 20574
rect 5073 20498 5139 20501
rect 2730 20496 5139 20498
rect 2730 20440 5078 20496
rect 5134 20440 5139 20496
rect 2730 20438 5139 20440
rect 5073 20435 5139 20438
rect 5809 20496 5875 20501
rect 9121 20500 9187 20501
rect 5809 20440 5814 20496
rect 5870 20440 5875 20496
rect 5809 20435 5875 20440
rect 9070 20436 9076 20500
rect 9140 20498 9187 20500
rect 9140 20496 9232 20498
rect 9182 20440 9232 20496
rect 9140 20438 9232 20440
rect 9140 20436 9187 20438
rect 9121 20435 9187 20436
rect 2446 20300 2452 20364
rect 2516 20362 2522 20364
rect 3325 20362 3391 20365
rect 2516 20360 3391 20362
rect 2516 20304 3330 20360
rect 3386 20304 3391 20360
rect 2516 20302 3391 20304
rect 2516 20300 2522 20302
rect 3325 20299 3391 20302
rect 4705 20362 4771 20365
rect 5812 20362 5872 20435
rect 4705 20360 5872 20362
rect 4705 20304 4710 20360
rect 4766 20304 5872 20360
rect 4705 20302 5872 20304
rect 4705 20299 4771 20302
rect 1342 20164 1348 20228
rect 1412 20226 1418 20228
rect 2630 20226 2636 20228
rect 1412 20166 2636 20226
rect 1412 20164 1418 20166
rect 2630 20164 2636 20166
rect 2700 20164 2706 20228
rect 5625 20226 5691 20229
rect 7373 20226 7439 20229
rect 5625 20224 7439 20226
rect 5625 20168 5630 20224
rect 5686 20168 7378 20224
rect 7434 20168 7439 20224
rect 5625 20166 7439 20168
rect 5625 20163 5691 20166
rect 7373 20163 7439 20166
rect 4318 20160 4634 20161
rect 4318 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4634 20160
rect 4318 20095 4634 20096
rect 10718 20160 11034 20161
rect 10718 20096 10724 20160
rect 10788 20096 10804 20160
rect 10868 20096 10884 20160
rect 10948 20096 10964 20160
rect 11028 20096 11034 20160
rect 10718 20095 11034 20096
rect 1894 20028 1900 20092
rect 1964 20090 1970 20092
rect 4153 20090 4219 20093
rect 1964 20088 4219 20090
rect 1964 20032 4158 20088
rect 4214 20032 4219 20088
rect 1964 20030 4219 20032
rect 1964 20028 1970 20030
rect 4153 20027 4219 20030
rect 6269 20090 6335 20093
rect 8150 20090 8156 20092
rect 6269 20088 8156 20090
rect 6269 20032 6274 20088
rect 6330 20032 8156 20088
rect 6269 20030 8156 20032
rect 6269 20027 6335 20030
rect 8150 20028 8156 20030
rect 8220 20028 8226 20092
rect 9213 20090 9279 20093
rect 9438 20090 9444 20092
rect 9213 20088 9444 20090
rect 9213 20032 9218 20088
rect 9274 20032 9444 20088
rect 9213 20030 9444 20032
rect 9213 20027 9279 20030
rect 9438 20028 9444 20030
rect 9508 20028 9514 20092
rect 2405 19956 2471 19957
rect 2405 19952 2452 19956
rect 2516 19954 2522 19956
rect 5206 19954 5212 19956
rect 2405 19896 2410 19952
rect 2405 19892 2452 19896
rect 2516 19894 2562 19954
rect 2730 19894 5212 19954
rect 2516 19892 2522 19894
rect 2405 19891 2471 19892
rect 1669 19818 1735 19821
rect 2313 19818 2379 19821
rect 1669 19816 2379 19818
rect 1669 19760 1674 19816
rect 1730 19760 2318 19816
rect 2374 19760 2379 19816
rect 1669 19758 2379 19760
rect 1669 19755 1735 19758
rect 2313 19755 2379 19758
rect 2037 19682 2103 19685
rect 2730 19682 2790 19894
rect 5206 19892 5212 19894
rect 5276 19892 5282 19956
rect 10869 19954 10935 19957
rect 11881 19954 11947 19957
rect 10869 19952 11947 19954
rect 10869 19896 10874 19952
rect 10930 19896 11886 19952
rect 11942 19896 11947 19952
rect 10869 19894 11947 19896
rect 10869 19891 10935 19894
rect 11881 19891 11947 19894
rect 2865 19816 2931 19821
rect 2865 19760 2870 19816
rect 2926 19760 2931 19816
rect 2865 19755 2931 19760
rect 3049 19818 3115 19821
rect 8293 19818 8359 19821
rect 3049 19816 8359 19818
rect 3049 19760 3054 19816
rect 3110 19760 8298 19816
rect 8354 19760 8359 19816
rect 3049 19758 8359 19760
rect 3049 19755 3115 19758
rect 8293 19755 8359 19758
rect 2037 19680 2790 19682
rect 2037 19624 2042 19680
rect 2098 19624 2790 19680
rect 2037 19622 2790 19624
rect 2868 19682 2928 19755
rect 3141 19682 3207 19685
rect 2868 19680 3207 19682
rect 2868 19624 3146 19680
rect 3202 19624 3207 19680
rect 2868 19622 3207 19624
rect 2037 19619 2103 19622
rect 3141 19619 3207 19622
rect 4521 19682 4587 19685
rect 4889 19684 4955 19685
rect 4838 19682 4844 19684
rect 4521 19680 4844 19682
rect 4908 19682 4955 19684
rect 5441 19682 5507 19685
rect 5574 19682 5580 19684
rect 4908 19680 5036 19682
rect 4521 19624 4526 19680
rect 4582 19624 4844 19680
rect 4950 19624 5036 19680
rect 4521 19622 4844 19624
rect 4521 19619 4587 19622
rect 4838 19620 4844 19622
rect 4908 19622 5036 19624
rect 5441 19680 5580 19682
rect 5441 19624 5446 19680
rect 5502 19624 5580 19680
rect 5441 19622 5580 19624
rect 4908 19620 4955 19622
rect 4889 19619 4955 19620
rect 5441 19619 5507 19622
rect 5574 19620 5580 19622
rect 5644 19620 5650 19684
rect 10542 19620 10548 19684
rect 10612 19682 10618 19684
rect 10685 19682 10751 19685
rect 10961 19682 11027 19685
rect 10612 19680 11027 19682
rect 10612 19624 10690 19680
rect 10746 19624 10966 19680
rect 11022 19624 11027 19680
rect 10612 19622 11027 19624
rect 10612 19620 10618 19622
rect 10685 19619 10751 19622
rect 10961 19619 11027 19622
rect 3658 19616 3974 19617
rect 3658 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3974 19616
rect 3658 19551 3974 19552
rect 10058 19616 10374 19617
rect 10058 19552 10064 19616
rect 10128 19552 10144 19616
rect 10208 19552 10224 19616
rect 10288 19552 10304 19616
rect 10368 19552 10374 19616
rect 10058 19551 10374 19552
rect 2681 19546 2747 19549
rect 3049 19546 3115 19549
rect 2681 19544 3115 19546
rect 2681 19488 2686 19544
rect 2742 19488 3054 19544
rect 3110 19488 3115 19544
rect 2681 19486 3115 19488
rect 2681 19483 2747 19486
rect 3049 19483 3115 19486
rect 4337 19546 4403 19549
rect 4838 19546 4844 19548
rect 4337 19544 4844 19546
rect 4337 19488 4342 19544
rect 4398 19488 4844 19544
rect 4337 19486 4844 19488
rect 4337 19483 4403 19486
rect 4838 19484 4844 19486
rect 4908 19484 4914 19548
rect 5257 19410 5323 19413
rect 1350 19408 5323 19410
rect 1350 19352 5262 19408
rect 5318 19352 5323 19408
rect 1350 19350 5323 19352
rect 749 19274 815 19277
rect 1350 19274 1410 19350
rect 5257 19347 5323 19350
rect 5574 19348 5580 19412
rect 5644 19410 5650 19412
rect 5993 19410 6059 19413
rect 5644 19408 6059 19410
rect 5644 19352 5998 19408
rect 6054 19352 6059 19408
rect 5644 19350 6059 19352
rect 5644 19348 5650 19350
rect 5993 19347 6059 19350
rect 7598 19348 7604 19412
rect 7668 19410 7674 19412
rect 8477 19410 8543 19413
rect 7668 19408 8543 19410
rect 7668 19352 8482 19408
rect 8538 19352 8543 19408
rect 7668 19350 8543 19352
rect 7668 19348 7674 19350
rect 8477 19347 8543 19350
rect 8661 19412 8727 19413
rect 8661 19408 8708 19412
rect 8772 19410 8778 19412
rect 12014 19410 12020 19412
rect 8661 19352 8666 19408
rect 8661 19348 8708 19352
rect 8772 19350 12020 19410
rect 8772 19348 8778 19350
rect 12014 19348 12020 19350
rect 12084 19348 12090 19412
rect 8661 19347 8727 19348
rect 2313 19276 2379 19277
rect 749 19272 1410 19274
rect 749 19216 754 19272
rect 810 19216 1410 19272
rect 749 19214 1410 19216
rect 749 19211 815 19214
rect 2262 19212 2268 19276
rect 2332 19274 2379 19276
rect 3693 19274 3759 19277
rect 6453 19276 6519 19277
rect 5942 19274 5948 19276
rect 2332 19272 3759 19274
rect 2374 19216 3698 19272
rect 3754 19216 3759 19272
rect 2332 19214 3759 19216
rect 2332 19212 2379 19214
rect 2313 19211 2379 19212
rect 3693 19211 3759 19214
rect 4156 19214 5948 19274
rect 3417 19138 3483 19141
rect 4156 19138 4216 19214
rect 5942 19212 5948 19214
rect 6012 19212 6018 19276
rect 6453 19274 6500 19276
rect 6408 19272 6500 19274
rect 6564 19274 6570 19276
rect 6821 19274 6887 19277
rect 6564 19272 6887 19274
rect 6408 19216 6458 19272
rect 6564 19216 6826 19272
rect 6882 19216 6887 19272
rect 6408 19214 6500 19216
rect 6453 19212 6500 19214
rect 6564 19214 6887 19216
rect 6564 19212 6570 19214
rect 6453 19211 6519 19212
rect 6821 19211 6887 19214
rect 7925 19274 7991 19277
rect 9029 19274 9095 19277
rect 7925 19272 9095 19274
rect 7925 19216 7930 19272
rect 7986 19216 9034 19272
rect 9090 19216 9095 19272
rect 7925 19214 9095 19216
rect 7925 19211 7991 19214
rect 9029 19211 9095 19214
rect 3417 19136 4216 19138
rect 3417 19080 3422 19136
rect 3478 19080 4216 19136
rect 3417 19078 4216 19080
rect 3417 19075 3483 19078
rect 4318 19072 4634 19073
rect 4318 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4634 19072
rect 4318 19007 4634 19008
rect 10718 19072 11034 19073
rect 10718 19008 10724 19072
rect 10788 19008 10804 19072
rect 10868 19008 10884 19072
rect 10948 19008 10964 19072
rect 11028 19008 11034 19072
rect 10718 19007 11034 19008
rect 2814 18940 2820 19004
rect 2884 19002 2890 19004
rect 3601 19002 3667 19005
rect 2884 19000 3667 19002
rect 2884 18944 3606 19000
rect 3662 18944 3667 19000
rect 2884 18942 3667 18944
rect 2884 18940 2890 18942
rect 3601 18939 3667 18942
rect 3785 19002 3851 19005
rect 5441 19004 5507 19005
rect 4102 19002 4108 19004
rect 3785 19000 4108 19002
rect 3785 18944 3790 19000
rect 3846 18944 4108 19000
rect 3785 18942 4108 18944
rect 3785 18939 3851 18942
rect 4102 18940 4108 18942
rect 4172 18940 4178 19004
rect 5390 18940 5396 19004
rect 5460 19002 5507 19004
rect 6269 19002 6335 19005
rect 7649 19002 7715 19005
rect 7925 19004 7991 19005
rect 7925 19002 7972 19004
rect 5460 19000 5552 19002
rect 5502 18944 5552 19000
rect 5460 18942 5552 18944
rect 6269 19000 7972 19002
rect 8036 19002 8042 19004
rect 6269 18944 6274 19000
rect 6330 18944 7654 19000
rect 7710 18944 7930 19000
rect 6269 18942 7972 18944
rect 5460 18940 5507 18942
rect 5441 18939 5507 18940
rect 6269 18939 6335 18942
rect 7649 18939 7715 18942
rect 7925 18940 7972 18942
rect 8036 18942 8118 19002
rect 8036 18940 8042 18942
rect 7925 18939 7991 18940
rect 3049 18866 3115 18869
rect 3366 18866 3372 18868
rect 3049 18864 3372 18866
rect 3049 18808 3054 18864
rect 3110 18808 3372 18864
rect 3049 18806 3372 18808
rect 3049 18803 3115 18806
rect 3366 18804 3372 18806
rect 3436 18866 3442 18868
rect 4061 18866 4127 18869
rect 3436 18864 4127 18866
rect 3436 18808 4066 18864
rect 4122 18808 4127 18864
rect 3436 18806 4127 18808
rect 3436 18804 3442 18806
rect 4061 18803 4127 18806
rect 6729 18866 6795 18869
rect 7005 18866 7071 18869
rect 6729 18864 7071 18866
rect 6729 18808 6734 18864
rect 6790 18808 7010 18864
rect 7066 18808 7071 18864
rect 6729 18806 7071 18808
rect 6729 18803 6795 18806
rect 7005 18803 7071 18806
rect 3366 18668 3372 18732
rect 3436 18730 3442 18732
rect 3509 18730 3575 18733
rect 3436 18728 3575 18730
rect 3436 18672 3514 18728
rect 3570 18672 3575 18728
rect 3436 18670 3575 18672
rect 3436 18668 3442 18670
rect 3509 18667 3575 18670
rect 4102 18668 4108 18732
rect 4172 18730 4178 18732
rect 4705 18730 4771 18733
rect 4172 18728 4771 18730
rect 4172 18672 4710 18728
rect 4766 18672 4771 18728
rect 4172 18670 4771 18672
rect 4172 18668 4178 18670
rect 4705 18667 4771 18670
rect 3658 18528 3974 18529
rect 3658 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3974 18528
rect 3658 18463 3974 18464
rect 10058 18528 10374 18529
rect 10058 18464 10064 18528
rect 10128 18464 10144 18528
rect 10208 18464 10224 18528
rect 10288 18464 10304 18528
rect 10368 18464 10374 18528
rect 10058 18463 10374 18464
rect 4061 18186 4127 18189
rect 4337 18186 4403 18189
rect 4061 18184 4403 18186
rect 4061 18128 4066 18184
rect 4122 18128 4342 18184
rect 4398 18128 4403 18184
rect 4061 18126 4403 18128
rect 4061 18123 4127 18126
rect 4337 18123 4403 18126
rect 4981 18186 5047 18189
rect 5993 18186 6059 18189
rect 4981 18184 6332 18186
rect 4981 18128 4986 18184
rect 5042 18128 5998 18184
rect 6054 18128 6332 18184
rect 4981 18126 6332 18128
rect 4981 18123 5047 18126
rect 5993 18123 6059 18126
rect 2129 18050 2195 18053
rect 3417 18050 3483 18053
rect 2129 18048 3483 18050
rect 2129 17992 2134 18048
rect 2190 17992 3422 18048
rect 3478 17992 3483 18048
rect 2129 17990 3483 17992
rect 2129 17987 2195 17990
rect 3417 17987 3483 17990
rect 5390 17988 5396 18052
rect 5460 18050 5466 18052
rect 6085 18050 6151 18053
rect 5460 18048 6151 18050
rect 5460 17992 6090 18048
rect 6146 17992 6151 18048
rect 5460 17990 6151 17992
rect 6272 18050 6332 18126
rect 6678 18124 6684 18188
rect 6748 18186 6754 18188
rect 12249 18186 12315 18189
rect 6748 18184 12315 18186
rect 6748 18128 12254 18184
rect 12310 18128 12315 18184
rect 6748 18126 12315 18128
rect 6748 18124 6754 18126
rect 12249 18123 12315 18126
rect 7189 18050 7255 18053
rect 8569 18050 8635 18053
rect 6272 18048 8635 18050
rect 6272 17992 7194 18048
rect 7250 17992 8574 18048
rect 8630 17992 8635 18048
rect 6272 17990 8635 17992
rect 5460 17988 5466 17990
rect 6085 17987 6151 17990
rect 7189 17987 7255 17990
rect 8569 17987 8635 17990
rect 4318 17984 4634 17985
rect 4318 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4634 17984
rect 4318 17919 4634 17920
rect 10718 17984 11034 17985
rect 10718 17920 10724 17984
rect 10788 17920 10804 17984
rect 10868 17920 10884 17984
rect 10948 17920 10964 17984
rect 11028 17920 11034 17984
rect 10718 17919 11034 17920
rect 6085 17916 6151 17917
rect 6085 17912 6132 17916
rect 6196 17914 6202 17916
rect 6085 17856 6090 17912
rect 6085 17852 6132 17856
rect 6196 17854 6242 17914
rect 6196 17852 6202 17854
rect 7782 17852 7788 17916
rect 7852 17914 7858 17916
rect 8569 17914 8635 17917
rect 7852 17912 8635 17914
rect 7852 17856 8574 17912
rect 8630 17856 8635 17912
rect 7852 17854 8635 17856
rect 7852 17852 7858 17854
rect 6085 17851 6151 17852
rect 8569 17851 8635 17854
rect 8753 17914 8819 17917
rect 9397 17916 9463 17917
rect 8886 17914 8892 17916
rect 8753 17912 8892 17914
rect 8753 17856 8758 17912
rect 8814 17856 8892 17912
rect 8753 17854 8892 17856
rect 8753 17851 8819 17854
rect 8886 17852 8892 17854
rect 8956 17852 8962 17916
rect 9397 17912 9444 17916
rect 9508 17914 9514 17916
rect 9397 17856 9402 17912
rect 9397 17852 9444 17856
rect 9508 17854 9554 17914
rect 9508 17852 9514 17854
rect 9397 17851 9463 17852
rect 422 17716 428 17780
rect 492 17778 498 17780
rect 933 17778 999 17781
rect 3182 17778 3188 17780
rect 492 17776 999 17778
rect 492 17720 938 17776
rect 994 17720 999 17776
rect 492 17718 999 17720
rect 492 17716 498 17718
rect 933 17715 999 17718
rect 1166 17718 3188 17778
rect 657 17642 723 17645
rect 1166 17642 1226 17718
rect 3182 17716 3188 17718
rect 3252 17716 3258 17780
rect 3417 17778 3483 17781
rect 3877 17778 3943 17781
rect 3417 17776 3943 17778
rect 3417 17720 3422 17776
rect 3478 17720 3882 17776
rect 3938 17720 3943 17776
rect 3417 17718 3943 17720
rect 3417 17715 3483 17718
rect 3877 17715 3943 17718
rect 4797 17778 4863 17781
rect 7046 17778 7052 17780
rect 4797 17776 7052 17778
rect 4797 17720 4802 17776
rect 4858 17720 7052 17776
rect 4797 17718 7052 17720
rect 4797 17715 4863 17718
rect 5996 17645 6056 17718
rect 7046 17716 7052 17718
rect 7116 17778 7122 17780
rect 7925 17778 7991 17781
rect 7116 17776 7991 17778
rect 7116 17720 7930 17776
rect 7986 17720 7991 17776
rect 7116 17718 7991 17720
rect 7116 17716 7122 17718
rect 7925 17715 7991 17718
rect 8201 17778 8267 17781
rect 9121 17780 9187 17781
rect 8702 17778 8708 17780
rect 8201 17776 8708 17778
rect 8201 17720 8206 17776
rect 8262 17720 8708 17776
rect 8201 17718 8708 17720
rect 8201 17715 8267 17718
rect 8702 17716 8708 17718
rect 8772 17716 8778 17780
rect 9070 17716 9076 17780
rect 9140 17778 9187 17780
rect 11421 17780 11487 17781
rect 11421 17778 11468 17780
rect 9140 17776 9232 17778
rect 9182 17720 9232 17776
rect 9140 17718 9232 17720
rect 11376 17776 11468 17778
rect 11376 17720 11426 17776
rect 11376 17718 11468 17720
rect 9140 17716 9187 17718
rect 9121 17715 9187 17716
rect 11421 17716 11468 17718
rect 11532 17716 11538 17780
rect 11421 17715 11487 17716
rect 657 17640 1226 17642
rect 657 17584 662 17640
rect 718 17584 1226 17640
rect 657 17582 1226 17584
rect 1945 17642 2011 17645
rect 1945 17640 5642 17642
rect 1945 17584 1950 17640
rect 2006 17584 5642 17640
rect 1945 17582 5642 17584
rect 657 17579 723 17582
rect 1945 17579 2011 17582
rect 5582 17506 5642 17582
rect 5993 17640 6059 17645
rect 5993 17584 5998 17640
rect 6054 17584 6059 17640
rect 5993 17579 6059 17584
rect 6453 17642 6519 17645
rect 7414 17642 7420 17644
rect 6453 17640 7420 17642
rect 6453 17584 6458 17640
rect 6514 17584 7420 17640
rect 6453 17582 7420 17584
rect 6453 17579 6519 17582
rect 7414 17580 7420 17582
rect 7484 17580 7490 17644
rect 7557 17642 7623 17645
rect 8845 17642 8911 17645
rect 11278 17642 11284 17644
rect 7557 17640 11284 17642
rect 7557 17584 7562 17640
rect 7618 17584 8850 17640
rect 8906 17584 11284 17640
rect 7557 17582 11284 17584
rect 7557 17579 7623 17582
rect 8845 17579 8911 17582
rect 11278 17580 11284 17582
rect 11348 17580 11354 17644
rect 8518 17506 8524 17508
rect 5582 17446 8524 17506
rect 8518 17444 8524 17446
rect 8588 17444 8594 17508
rect 3658 17440 3974 17441
rect 3658 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3974 17440
rect 3658 17375 3974 17376
rect 10058 17440 10374 17441
rect 10058 17376 10064 17440
rect 10128 17376 10144 17440
rect 10208 17376 10224 17440
rect 10288 17376 10304 17440
rect 10368 17376 10374 17440
rect 10058 17375 10374 17376
rect 5758 17308 5764 17372
rect 5828 17370 5834 17372
rect 9121 17370 9187 17373
rect 5828 17368 9187 17370
rect 5828 17312 9126 17368
rect 9182 17312 9187 17368
rect 5828 17310 9187 17312
rect 5828 17308 5834 17310
rect 9121 17307 9187 17310
rect 0 17234 400 17264
rect 841 17234 907 17237
rect 0 17232 907 17234
rect 0 17176 846 17232
rect 902 17176 907 17232
rect 0 17174 907 17176
rect 0 17144 400 17174
rect 841 17171 907 17174
rect 6637 17236 6703 17237
rect 6637 17232 6684 17236
rect 6748 17234 6754 17236
rect 6637 17176 6642 17232
rect 6637 17172 6684 17176
rect 6748 17174 6794 17234
rect 6748 17172 6754 17174
rect 9622 17172 9628 17236
rect 9692 17234 9698 17236
rect 9765 17234 9831 17237
rect 9692 17232 9831 17234
rect 9692 17176 9770 17232
rect 9826 17176 9831 17232
rect 9692 17174 9831 17176
rect 9692 17172 9698 17174
rect 6637 17171 6703 17172
rect 9765 17171 9831 17174
rect 2129 17098 2195 17101
rect 2262 17098 2268 17100
rect 2129 17096 2268 17098
rect 2129 17040 2134 17096
rect 2190 17040 2268 17096
rect 2129 17038 2268 17040
rect 2129 17035 2195 17038
rect 2262 17036 2268 17038
rect 2332 17036 2338 17100
rect 2589 17098 2655 17101
rect 2814 17098 2820 17100
rect 2589 17096 2820 17098
rect 2589 17040 2594 17096
rect 2650 17040 2820 17096
rect 2589 17038 2820 17040
rect 2589 17035 2655 17038
rect 2814 17036 2820 17038
rect 2884 17036 2890 17100
rect 4521 17098 4587 17101
rect 4981 17098 5047 17101
rect 6361 17098 6427 17101
rect 6545 17098 6611 17101
rect 4521 17096 4906 17098
rect 4521 17040 4526 17096
rect 4582 17040 4906 17096
rect 4521 17038 4906 17040
rect 4521 17035 4587 17038
rect 0 16962 400 16992
rect 933 16962 999 16965
rect 0 16960 999 16962
rect 0 16904 938 16960
rect 994 16904 999 16960
rect 0 16902 999 16904
rect 0 16872 400 16902
rect 933 16899 999 16902
rect 4318 16896 4634 16897
rect 4318 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4634 16896
rect 4318 16831 4634 16832
rect 1301 16826 1367 16829
rect 2630 16826 2636 16828
rect 1301 16824 2636 16826
rect 1301 16768 1306 16824
rect 1362 16768 2636 16824
rect 1301 16766 2636 16768
rect 1301 16763 1367 16766
rect 2630 16764 2636 16766
rect 2700 16764 2706 16828
rect 4846 16826 4906 17038
rect 4981 17096 6611 17098
rect 4981 17040 4986 17096
rect 5042 17040 6366 17096
rect 6422 17040 6550 17096
rect 6606 17040 6611 17096
rect 4981 17038 6611 17040
rect 4981 17035 5047 17038
rect 6361 17035 6427 17038
rect 6545 17035 6611 17038
rect 6729 17098 6795 17101
rect 9949 17098 10015 17101
rect 6729 17096 10015 17098
rect 6729 17040 6734 17096
rect 6790 17040 9954 17096
rect 10010 17040 10015 17096
rect 6729 17038 10015 17040
rect 6729 17035 6795 17038
rect 9949 17035 10015 17038
rect 5257 16962 5323 16965
rect 6678 16962 6684 16964
rect 5257 16960 6684 16962
rect 5257 16904 5262 16960
rect 5318 16904 6684 16960
rect 5257 16902 6684 16904
rect 5257 16899 5323 16902
rect 6678 16900 6684 16902
rect 6748 16900 6754 16964
rect 10718 16896 11034 16897
rect 10718 16832 10724 16896
rect 10788 16832 10804 16896
rect 10868 16832 10884 16896
rect 10948 16832 10964 16896
rect 11028 16832 11034 16896
rect 10718 16831 11034 16832
rect 4846 16766 7712 16826
rect 0 16690 400 16720
rect 1945 16690 2011 16693
rect 0 16688 2011 16690
rect 0 16632 1950 16688
rect 2006 16632 2011 16688
rect 0 16630 2011 16632
rect 0 16600 400 16630
rect 1945 16627 2011 16630
rect 3182 16628 3188 16692
rect 3252 16690 3258 16692
rect 6085 16690 6151 16693
rect 3252 16688 6151 16690
rect 3252 16632 6090 16688
rect 6146 16632 6151 16688
rect 3252 16630 6151 16632
rect 3252 16628 3258 16630
rect 6085 16627 6151 16630
rect 6545 16690 6611 16693
rect 7373 16690 7439 16693
rect 6545 16688 7439 16690
rect 6545 16632 6550 16688
rect 6606 16632 7378 16688
rect 7434 16632 7439 16688
rect 6545 16630 7439 16632
rect 7652 16690 7712 16766
rect 7833 16690 7899 16693
rect 7652 16688 7899 16690
rect 7652 16632 7838 16688
rect 7894 16632 7899 16688
rect 7652 16630 7899 16632
rect 6545 16627 6611 16630
rect 7373 16627 7439 16630
rect 7833 16627 7899 16630
rect 9070 16628 9076 16692
rect 9140 16690 9146 16692
rect 9305 16690 9371 16693
rect 9140 16688 9371 16690
rect 9140 16632 9310 16688
rect 9366 16632 9371 16688
rect 9140 16630 9371 16632
rect 9140 16628 9146 16630
rect 9305 16627 9371 16630
rect 9765 16690 9831 16693
rect 10961 16690 11027 16693
rect 9765 16688 11027 16690
rect 9765 16632 9770 16688
rect 9826 16632 10966 16688
rect 11022 16632 11027 16688
rect 9765 16630 11027 16632
rect 9765 16627 9831 16630
rect 10961 16627 11027 16630
rect 933 16554 999 16557
rect 1158 16554 1164 16556
rect 933 16552 1164 16554
rect 933 16496 938 16552
rect 994 16496 1164 16552
rect 933 16494 1164 16496
rect 933 16491 999 16494
rect 1158 16492 1164 16494
rect 1228 16492 1234 16556
rect 1485 16554 1551 16557
rect 2957 16554 3023 16557
rect 1485 16552 3023 16554
rect 1485 16496 1490 16552
rect 1546 16496 2962 16552
rect 3018 16496 3023 16552
rect 1485 16494 3023 16496
rect 1485 16491 1551 16494
rect 2957 16491 3023 16494
rect 4429 16554 4495 16557
rect 6453 16554 6519 16557
rect 4429 16552 6519 16554
rect 4429 16496 4434 16552
rect 4490 16496 6458 16552
rect 6514 16496 6519 16552
rect 4429 16494 6519 16496
rect 4429 16491 4495 16494
rect 6453 16491 6519 16494
rect 7281 16554 7347 16557
rect 7649 16554 7715 16557
rect 7281 16552 7715 16554
rect 7281 16496 7286 16552
rect 7342 16496 7654 16552
rect 7710 16496 7715 16552
rect 7281 16494 7715 16496
rect 7281 16491 7347 16494
rect 7649 16491 7715 16494
rect 7782 16492 7788 16556
rect 7852 16554 7858 16556
rect 9806 16554 9812 16556
rect 7852 16494 9812 16554
rect 7852 16492 7858 16494
rect 9806 16492 9812 16494
rect 9876 16492 9882 16556
rect 0 16418 400 16448
rect 1342 16418 1348 16420
rect 0 16358 1348 16418
rect 0 16328 400 16358
rect 1342 16356 1348 16358
rect 1412 16356 1418 16420
rect 4838 16356 4844 16420
rect 4908 16418 4914 16420
rect 5073 16418 5139 16421
rect 4908 16416 5139 16418
rect 4908 16360 5078 16416
rect 5134 16360 5139 16416
rect 4908 16358 5139 16360
rect 4908 16356 4914 16358
rect 5073 16355 5139 16358
rect 3658 16352 3974 16353
rect 3658 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3974 16352
rect 3658 16287 3974 16288
rect 10058 16352 10374 16353
rect 10058 16288 10064 16352
rect 10128 16288 10144 16352
rect 10208 16288 10224 16352
rect 10288 16288 10304 16352
rect 10368 16288 10374 16352
rect 10058 16287 10374 16288
rect 4102 16220 4108 16284
rect 4172 16282 4178 16284
rect 6545 16282 6611 16285
rect 4172 16280 6611 16282
rect 4172 16224 6550 16280
rect 6606 16224 6611 16280
rect 4172 16222 6611 16224
rect 4172 16220 4178 16222
rect 6545 16219 6611 16222
rect 9673 16282 9739 16285
rect 9806 16282 9812 16284
rect 9673 16280 9812 16282
rect 9673 16224 9678 16280
rect 9734 16224 9812 16280
rect 9673 16222 9812 16224
rect 9673 16219 9739 16222
rect 9806 16220 9812 16222
rect 9876 16220 9882 16284
rect 974 16084 980 16148
rect 1044 16146 1050 16148
rect 2681 16146 2747 16149
rect 1044 16144 2747 16146
rect 1044 16088 2686 16144
rect 2742 16088 2747 16144
rect 1044 16086 2747 16088
rect 1044 16084 1050 16086
rect 2681 16083 2747 16086
rect 9254 16084 9260 16148
rect 9324 16146 9330 16148
rect 9581 16146 9647 16149
rect 9324 16144 9647 16146
rect 9324 16088 9586 16144
rect 9642 16088 9647 16144
rect 9324 16086 9647 16088
rect 9324 16084 9330 16086
rect 9581 16083 9647 16086
rect 606 15812 612 15876
rect 676 15874 682 15876
rect 3509 15874 3575 15877
rect 676 15872 3575 15874
rect 676 15816 3514 15872
rect 3570 15816 3575 15872
rect 676 15814 3575 15816
rect 676 15812 682 15814
rect 3509 15811 3575 15814
rect 4318 15808 4634 15809
rect 4318 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4634 15808
rect 4318 15743 4634 15744
rect 10718 15808 11034 15809
rect 10718 15744 10724 15808
rect 10788 15744 10804 15808
rect 10868 15744 10884 15808
rect 10948 15744 10964 15808
rect 11028 15744 11034 15808
rect 10718 15743 11034 15744
rect 1669 15740 1735 15741
rect 1669 15738 1716 15740
rect 1624 15736 1716 15738
rect 1624 15680 1674 15736
rect 1624 15678 1716 15680
rect 1669 15676 1716 15678
rect 1780 15676 1786 15740
rect 1669 15675 1735 15676
rect 2037 15602 2103 15605
rect 8201 15602 8267 15605
rect 11789 15604 11855 15605
rect 11789 15602 11836 15604
rect 2037 15600 8267 15602
rect 2037 15544 2042 15600
rect 2098 15544 8206 15600
rect 8262 15544 8267 15600
rect 2037 15542 8267 15544
rect 11744 15600 11836 15602
rect 11744 15544 11794 15600
rect 11744 15542 11836 15544
rect 2037 15539 2103 15542
rect 8201 15539 8267 15542
rect 11789 15540 11836 15542
rect 11900 15540 11906 15604
rect 11789 15539 11855 15540
rect 54 15404 60 15468
rect 124 15466 130 15468
rect 2630 15466 2636 15468
rect 124 15406 2636 15466
rect 124 15404 130 15406
rect 2630 15404 2636 15406
rect 2700 15404 2706 15468
rect 473 15330 539 15333
rect 2957 15330 3023 15333
rect 3182 15330 3188 15332
rect 473 15328 1594 15330
rect 473 15272 478 15328
rect 534 15272 1594 15328
rect 473 15270 1594 15272
rect 473 15267 539 15270
rect 1534 15194 1594 15270
rect 2957 15328 3188 15330
rect 2957 15272 2962 15328
rect 3018 15272 3188 15328
rect 2957 15270 3188 15272
rect 2957 15267 3023 15270
rect 3182 15268 3188 15270
rect 3252 15268 3258 15332
rect 8477 15330 8543 15333
rect 9254 15330 9260 15332
rect 8477 15328 9260 15330
rect 8477 15272 8482 15328
rect 8538 15272 9260 15328
rect 8477 15270 9260 15272
rect 8477 15267 8543 15270
rect 9254 15268 9260 15270
rect 9324 15268 9330 15332
rect 3658 15264 3974 15265
rect 3658 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3974 15264
rect 3658 15199 3974 15200
rect 10058 15264 10374 15265
rect 10058 15200 10064 15264
rect 10128 15200 10144 15264
rect 10208 15200 10224 15264
rect 10288 15200 10304 15264
rect 10368 15200 10374 15264
rect 10058 15199 10374 15200
rect 1669 15194 1735 15197
rect 1534 15192 1735 15194
rect 1534 15136 1674 15192
rect 1730 15136 1735 15192
rect 1534 15134 1735 15136
rect 1669 15131 1735 15134
rect 3969 15058 4035 15061
rect 4153 15058 4219 15061
rect 3969 15056 4219 15058
rect 3969 15000 3974 15056
rect 4030 15000 4158 15056
rect 4214 15000 4219 15056
rect 3969 14998 4219 15000
rect 3969 14995 4035 14998
rect 4153 14995 4219 14998
rect 7833 15058 7899 15061
rect 8937 15058 9003 15061
rect 7833 15056 9003 15058
rect 7833 15000 7838 15056
rect 7894 15000 8942 15056
rect 8998 15000 9003 15056
rect 7833 14998 9003 15000
rect 7833 14995 7899 14998
rect 8937 14995 9003 14998
rect 3366 14860 3372 14924
rect 3436 14922 3442 14924
rect 3693 14922 3759 14925
rect 11145 14922 11211 14925
rect 11421 14922 11487 14925
rect 12566 14922 12572 14924
rect 3436 14920 5136 14922
rect 3436 14864 3698 14920
rect 3754 14864 5136 14920
rect 3436 14862 5136 14864
rect 3436 14860 3442 14862
rect 3693 14859 3759 14862
rect 5076 14789 5136 14862
rect 11145 14920 12572 14922
rect 11145 14864 11150 14920
rect 11206 14864 11426 14920
rect 11482 14864 12572 14920
rect 11145 14862 12572 14864
rect 11145 14859 11211 14862
rect 11421 14859 11487 14862
rect 12566 14860 12572 14862
rect 12636 14860 12642 14924
rect 5073 14784 5139 14789
rect 5073 14728 5078 14784
rect 5134 14728 5139 14784
rect 5073 14723 5139 14728
rect 4318 14720 4634 14721
rect 4318 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4634 14720
rect 4318 14655 4634 14656
rect 10718 14720 11034 14721
rect 10718 14656 10724 14720
rect 10788 14656 10804 14720
rect 10868 14656 10884 14720
rect 10948 14656 10964 14720
rect 11028 14656 11034 14720
rect 10718 14655 11034 14656
rect 4153 14514 4219 14517
rect 5022 14514 5028 14516
rect 4153 14512 5028 14514
rect 4153 14456 4158 14512
rect 4214 14456 5028 14512
rect 4153 14454 5028 14456
rect 4153 14451 4219 14454
rect 5022 14452 5028 14454
rect 5092 14452 5098 14516
rect 6310 14452 6316 14516
rect 6380 14514 6386 14516
rect 9305 14514 9371 14517
rect 6380 14512 9371 14514
rect 6380 14456 9310 14512
rect 9366 14456 9371 14512
rect 6380 14454 9371 14456
rect 6380 14452 6386 14454
rect 9305 14451 9371 14454
rect 3658 14176 3974 14177
rect 3658 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3974 14176
rect 3658 14111 3974 14112
rect 10058 14176 10374 14177
rect 10058 14112 10064 14176
rect 10128 14112 10144 14176
rect 10208 14112 10224 14176
rect 10288 14112 10304 14176
rect 10368 14112 10374 14176
rect 10058 14111 10374 14112
rect 5758 13772 5764 13836
rect 5828 13834 5834 13836
rect 6361 13834 6427 13837
rect 5828 13832 6427 13834
rect 5828 13776 6366 13832
rect 6422 13776 6427 13832
rect 5828 13774 6427 13776
rect 5828 13772 5834 13774
rect 6361 13771 6427 13774
rect 6177 13698 6243 13701
rect 11697 13700 11763 13701
rect 7782 13698 7788 13700
rect 6177 13696 7788 13698
rect 6177 13640 6182 13696
rect 6238 13640 7788 13696
rect 6177 13638 7788 13640
rect 6177 13635 6243 13638
rect 7782 13636 7788 13638
rect 7852 13636 7858 13700
rect 11646 13636 11652 13700
rect 11716 13698 11763 13700
rect 11716 13696 11808 13698
rect 11758 13640 11808 13696
rect 11716 13638 11808 13640
rect 11716 13636 11763 13638
rect 11697 13635 11763 13636
rect 4318 13632 4634 13633
rect 4318 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4634 13632
rect 4318 13567 4634 13568
rect 10718 13632 11034 13633
rect 10718 13568 10724 13632
rect 10788 13568 10804 13632
rect 10868 13568 10884 13632
rect 10948 13568 10964 13632
rect 11028 13568 11034 13632
rect 10718 13567 11034 13568
rect 3658 13088 3974 13089
rect 3658 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3974 13088
rect 3658 13023 3974 13024
rect 10058 13088 10374 13089
rect 10058 13024 10064 13088
rect 10128 13024 10144 13088
rect 10208 13024 10224 13088
rect 10288 13024 10304 13088
rect 10368 13024 10374 13088
rect 10058 13023 10374 13024
rect 4153 13018 4219 13021
rect 4153 13016 8954 13018
rect 4153 12960 4158 13016
rect 4214 12960 8954 13016
rect 4153 12958 8954 12960
rect 4153 12955 4219 12958
rect 8894 12885 8954 12958
rect 5942 12820 5948 12884
rect 6012 12882 6018 12884
rect 7741 12882 7807 12885
rect 8894 12884 9003 12885
rect 6012 12880 7807 12882
rect 6012 12824 7746 12880
rect 7802 12824 7807 12880
rect 6012 12822 7807 12824
rect 6012 12820 6018 12822
rect 7741 12819 7807 12822
rect 8886 12820 8892 12884
rect 8956 12882 9003 12884
rect 8956 12880 9048 12882
rect 8998 12824 9048 12880
rect 8956 12822 9048 12824
rect 8956 12820 9003 12822
rect 8937 12819 9003 12820
rect 2773 12746 2839 12749
rect 6085 12746 6151 12749
rect 9121 12746 9187 12749
rect 2773 12744 6010 12746
rect 2773 12688 2778 12744
rect 2834 12688 6010 12744
rect 2773 12686 6010 12688
rect 2773 12683 2839 12686
rect 0 12610 400 12640
rect 841 12610 907 12613
rect 0 12608 907 12610
rect 0 12552 846 12608
rect 902 12552 907 12608
rect 0 12550 907 12552
rect 5950 12610 6010 12686
rect 6085 12744 9187 12746
rect 6085 12688 6090 12744
rect 6146 12688 9126 12744
rect 9182 12688 9187 12744
rect 6085 12686 9187 12688
rect 6085 12683 6151 12686
rect 9121 12683 9187 12686
rect 7005 12610 7071 12613
rect 5950 12608 7071 12610
rect 5950 12552 7010 12608
rect 7066 12552 7071 12608
rect 5950 12550 7071 12552
rect 0 12520 400 12550
rect 841 12547 907 12550
rect 7005 12547 7071 12550
rect 4318 12544 4634 12545
rect 4318 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4634 12544
rect 4318 12479 4634 12480
rect 10718 12544 11034 12545
rect 10718 12480 10724 12544
rect 10788 12480 10804 12544
rect 10868 12480 10884 12544
rect 10948 12480 10964 12544
rect 11028 12480 11034 12544
rect 10718 12479 11034 12480
rect 5257 12476 5323 12477
rect 5206 12412 5212 12476
rect 5276 12474 5323 12476
rect 7649 12474 7715 12477
rect 8661 12474 8727 12477
rect 11145 12476 11211 12477
rect 5276 12472 5368 12474
rect 5318 12416 5368 12472
rect 5276 12414 5368 12416
rect 7054 12472 8727 12474
rect 7054 12416 7654 12472
rect 7710 12416 8666 12472
rect 8722 12416 8727 12472
rect 7054 12414 8727 12416
rect 5276 12412 5323 12414
rect 5257 12411 5323 12412
rect 0 12338 400 12368
rect 7054 12341 7114 12414
rect 7649 12411 7715 12414
rect 8661 12411 8727 12414
rect 11094 12412 11100 12476
rect 11164 12474 11211 12476
rect 11164 12472 11256 12474
rect 11206 12416 11256 12472
rect 11164 12414 11256 12416
rect 11164 12412 11211 12414
rect 11145 12411 11211 12412
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 400 12278
rect 1393 12275 1459 12278
rect 4153 12338 4219 12341
rect 4429 12338 4495 12341
rect 5257 12340 5323 12341
rect 4153 12336 4495 12338
rect 4153 12280 4158 12336
rect 4214 12280 4434 12336
rect 4490 12280 4495 12336
rect 4153 12278 4495 12280
rect 4153 12275 4219 12278
rect 4429 12275 4495 12278
rect 5206 12276 5212 12340
rect 5276 12338 5323 12340
rect 5276 12336 5368 12338
rect 5318 12280 5368 12336
rect 5276 12278 5368 12280
rect 7005 12336 7114 12341
rect 7005 12280 7010 12336
rect 7066 12280 7114 12336
rect 7005 12278 7114 12280
rect 7373 12338 7439 12341
rect 7649 12338 7715 12341
rect 9121 12338 9187 12341
rect 7373 12336 9187 12338
rect 7373 12280 7378 12336
rect 7434 12280 7654 12336
rect 7710 12280 9126 12336
rect 9182 12280 9187 12336
rect 7373 12278 9187 12280
rect 5276 12276 5323 12278
rect 5257 12275 5323 12276
rect 7005 12275 7071 12278
rect 7373 12275 7439 12278
rect 7649 12275 7715 12278
rect 9121 12275 9187 12278
rect 10542 12276 10548 12340
rect 10612 12338 10618 12340
rect 10961 12338 11027 12341
rect 10612 12336 11027 12338
rect 10612 12280 10966 12336
rect 11022 12280 11027 12336
rect 10612 12278 11027 12280
rect 10612 12276 10618 12278
rect 10961 12275 11027 12278
rect 6729 12202 6795 12205
rect 10041 12202 10107 12205
rect 6729 12200 10107 12202
rect 6729 12144 6734 12200
rect 6790 12144 10046 12200
rect 10102 12144 10107 12200
rect 6729 12142 10107 12144
rect 6729 12139 6795 12142
rect 10041 12139 10107 12142
rect 0 12066 400 12096
rect 933 12066 999 12069
rect 0 12064 999 12066
rect 0 12008 938 12064
rect 994 12008 999 12064
rect 0 12006 999 12008
rect 0 11976 400 12006
rect 933 12003 999 12006
rect 7097 12066 7163 12069
rect 8109 12066 8175 12069
rect 7097 12064 8175 12066
rect 7097 12008 7102 12064
rect 7158 12008 8114 12064
rect 8170 12008 8175 12064
rect 7097 12006 8175 12008
rect 7097 12003 7163 12006
rect 8109 12003 8175 12006
rect 3658 12000 3974 12001
rect 3658 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3974 12000
rect 3658 11935 3974 11936
rect 10058 12000 10374 12001
rect 10058 11936 10064 12000
rect 10128 11936 10144 12000
rect 10208 11936 10224 12000
rect 10288 11936 10304 12000
rect 10368 11936 10374 12000
rect 10058 11935 10374 11936
rect 0 11794 400 11824
rect 1209 11794 1275 11797
rect 0 11792 1275 11794
rect 0 11736 1214 11792
rect 1270 11736 1275 11792
rect 0 11734 1275 11736
rect 0 11704 400 11734
rect 1209 11731 1275 11734
rect 0 11522 400 11552
rect 1025 11522 1091 11525
rect 0 11520 1091 11522
rect 0 11464 1030 11520
rect 1086 11464 1091 11520
rect 0 11462 1091 11464
rect 0 11432 400 11462
rect 1025 11459 1091 11462
rect 4318 11456 4634 11457
rect 4318 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4634 11456
rect 4318 11391 4634 11392
rect 10718 11456 11034 11457
rect 10718 11392 10724 11456
rect 10788 11392 10804 11456
rect 10868 11392 10884 11456
rect 10948 11392 10964 11456
rect 11028 11392 11034 11456
rect 10718 11391 11034 11392
rect 0 11250 400 11280
rect 565 11250 631 11253
rect 0 11248 631 11250
rect 0 11192 570 11248
rect 626 11192 631 11248
rect 0 11190 631 11192
rect 0 11160 400 11190
rect 565 11187 631 11190
rect 1945 11250 2011 11253
rect 2078 11250 2084 11252
rect 1945 11248 2084 11250
rect 1945 11192 1950 11248
rect 2006 11192 2084 11248
rect 1945 11190 2084 11192
rect 1945 11187 2011 11190
rect 2078 11188 2084 11190
rect 2148 11188 2154 11252
rect 8109 11116 8175 11117
rect 8109 11114 8156 11116
rect 8064 11112 8156 11114
rect 8064 11056 8114 11112
rect 8064 11054 8156 11056
rect 8109 11052 8156 11054
rect 8220 11052 8226 11116
rect 8109 11051 8175 11052
rect 0 10978 400 11008
rect 2497 10978 2563 10981
rect 0 10976 2563 10978
rect 0 10920 2502 10976
rect 2558 10920 2563 10976
rect 0 10918 2563 10920
rect 0 10888 400 10918
rect 2497 10915 2563 10918
rect 3658 10912 3974 10913
rect 3658 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3974 10912
rect 3658 10847 3974 10848
rect 10058 10912 10374 10913
rect 10058 10848 10064 10912
rect 10128 10848 10144 10912
rect 10208 10848 10224 10912
rect 10288 10848 10304 10912
rect 10368 10848 10374 10912
rect 10058 10847 10374 10848
rect 4318 10368 4634 10369
rect 4318 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4634 10368
rect 4318 10303 4634 10304
rect 10718 10368 11034 10369
rect 10718 10304 10724 10368
rect 10788 10304 10804 10368
rect 10868 10304 10884 10368
rect 10948 10304 10964 10368
rect 11028 10304 11034 10368
rect 10718 10303 11034 10304
rect 3601 10026 3667 10029
rect 4797 10026 4863 10029
rect 9857 10028 9923 10029
rect 5390 10026 5396 10028
rect 3601 10024 5396 10026
rect 3601 9968 3606 10024
rect 3662 9968 4802 10024
rect 4858 9968 5396 10024
rect 3601 9966 5396 9968
rect 3601 9963 3667 9966
rect 4797 9963 4863 9966
rect 5390 9964 5396 9966
rect 5460 9964 5466 10028
rect 9806 9964 9812 10028
rect 9876 10026 9923 10028
rect 10593 10026 10659 10029
rect 11094 10026 11100 10028
rect 9876 10024 9968 10026
rect 9918 9968 9968 10024
rect 9876 9966 9968 9968
rect 10593 10024 11100 10026
rect 10593 9968 10598 10024
rect 10654 9968 11100 10024
rect 10593 9966 11100 9968
rect 9876 9964 9923 9966
rect 9857 9963 9923 9964
rect 10593 9963 10659 9966
rect 11094 9964 11100 9966
rect 11164 9964 11170 10028
rect 3658 9824 3974 9825
rect 3658 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3974 9824
rect 3658 9759 3974 9760
rect 10058 9824 10374 9825
rect 10058 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10374 9824
rect 10058 9759 10374 9760
rect 9949 9618 10015 9621
rect 11145 9618 11211 9621
rect 9949 9616 11211 9618
rect 9949 9560 9954 9616
rect 10010 9560 11150 9616
rect 11206 9560 11211 9616
rect 9949 9558 11211 9560
rect 9949 9555 10015 9558
rect 11145 9555 11211 9558
rect 10542 9420 10548 9484
rect 10612 9482 10618 9484
rect 10685 9482 10751 9485
rect 10612 9480 10751 9482
rect 10612 9424 10690 9480
rect 10746 9424 10751 9480
rect 10612 9422 10751 9424
rect 10612 9420 10618 9422
rect 10685 9419 10751 9422
rect 4318 9280 4634 9281
rect 4318 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4634 9280
rect 4318 9215 4634 9216
rect 10718 9280 11034 9281
rect 10718 9216 10724 9280
rect 10788 9216 10804 9280
rect 10868 9216 10884 9280
rect 10948 9216 10964 9280
rect 11028 9216 11034 9280
rect 10718 9215 11034 9216
rect 3417 8938 3483 8941
rect 3601 8938 3667 8941
rect 4521 8938 4587 8941
rect 3417 8936 4587 8938
rect 3417 8880 3422 8936
rect 3478 8880 3606 8936
rect 3662 8880 4526 8936
rect 4582 8880 4587 8936
rect 3417 8878 4587 8880
rect 3417 8875 3483 8878
rect 3601 8875 3667 8878
rect 4521 8875 4587 8878
rect 3658 8736 3974 8737
rect 3658 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3974 8736
rect 3658 8671 3974 8672
rect 10058 8736 10374 8737
rect 10058 8672 10064 8736
rect 10128 8672 10144 8736
rect 10208 8672 10224 8736
rect 10288 8672 10304 8736
rect 10368 8672 10374 8736
rect 10058 8671 10374 8672
rect 5533 8668 5599 8669
rect 5533 8666 5580 8668
rect 5488 8664 5580 8666
rect 5488 8608 5538 8664
rect 5488 8606 5580 8608
rect 5533 8604 5580 8606
rect 5644 8604 5650 8668
rect 5533 8603 5599 8604
rect 4889 8394 4955 8397
rect 7465 8394 7531 8397
rect 4889 8392 7531 8394
rect 4889 8336 4894 8392
rect 4950 8336 7470 8392
rect 7526 8336 7531 8392
rect 4889 8334 7531 8336
rect 4889 8331 4955 8334
rect 7465 8331 7531 8334
rect 7414 8196 7420 8260
rect 7484 8258 7490 8260
rect 10317 8258 10383 8261
rect 7484 8256 10383 8258
rect 7484 8200 10322 8256
rect 10378 8200 10383 8256
rect 7484 8198 10383 8200
rect 7484 8196 7490 8198
rect 10317 8195 10383 8198
rect 4318 8192 4634 8193
rect 4318 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4634 8192
rect 4318 8127 4634 8128
rect 10718 8192 11034 8193
rect 10718 8128 10724 8192
rect 10788 8128 10804 8192
rect 10868 8128 10884 8192
rect 10948 8128 10964 8192
rect 11028 8128 11034 8192
rect 10718 8127 11034 8128
rect 9489 8124 9555 8125
rect 9438 8060 9444 8124
rect 9508 8122 9555 8124
rect 9508 8120 9600 8122
rect 9550 8064 9600 8120
rect 9508 8062 9600 8064
rect 9508 8060 9555 8062
rect 9489 8059 9555 8060
rect 3658 7648 3974 7649
rect 3658 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3974 7648
rect 3658 7583 3974 7584
rect 10058 7648 10374 7649
rect 10058 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10374 7648
rect 10058 7583 10374 7584
rect 8569 7442 8635 7445
rect 9070 7442 9076 7444
rect 8569 7440 9076 7442
rect 8569 7384 8574 7440
rect 8630 7384 9076 7440
rect 8569 7382 9076 7384
rect 8569 7379 8635 7382
rect 9070 7380 9076 7382
rect 9140 7380 9146 7444
rect 9765 7308 9831 7309
rect 9765 7304 9812 7308
rect 9876 7306 9882 7308
rect 9765 7248 9770 7304
rect 9765 7244 9812 7248
rect 9876 7246 9922 7306
rect 9876 7244 9882 7246
rect 9765 7243 9831 7244
rect 54 7108 60 7172
rect 124 7170 130 7172
rect 381 7170 447 7173
rect 124 7168 447 7170
rect 124 7112 386 7168
rect 442 7112 447 7168
rect 124 7110 447 7112
rect 124 7108 130 7110
rect 381 7107 447 7110
rect 4318 7104 4634 7105
rect 4318 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4634 7104
rect 4318 7039 4634 7040
rect 10718 7104 11034 7105
rect 10718 7040 10724 7104
rect 10788 7040 10804 7104
rect 10868 7040 10884 7104
rect 10948 7040 10964 7104
rect 11028 7040 11034 7104
rect 10718 7039 11034 7040
rect 9765 6898 9831 6901
rect 10542 6898 10548 6900
rect 9765 6896 10548 6898
rect 9765 6840 9770 6896
rect 9826 6840 10548 6896
rect 9765 6838 10548 6840
rect 9765 6835 9831 6838
rect 10542 6836 10548 6838
rect 10612 6836 10618 6900
rect 3658 6560 3974 6561
rect 3658 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3974 6560
rect 3658 6495 3974 6496
rect 10058 6560 10374 6561
rect 10058 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10374 6560
rect 10058 6495 10374 6496
rect 9673 6218 9739 6221
rect 10869 6218 10935 6221
rect 9673 6216 10935 6218
rect 9673 6160 9678 6216
rect 9734 6160 10874 6216
rect 10930 6160 10935 6216
rect 9673 6158 10935 6160
rect 9673 6155 9739 6158
rect 10869 6155 10935 6158
rect 4318 6016 4634 6017
rect 4318 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4634 6016
rect 4318 5951 4634 5952
rect 10718 6016 11034 6017
rect 10718 5952 10724 6016
rect 10788 5952 10804 6016
rect 10868 5952 10884 6016
rect 10948 5952 10964 6016
rect 11028 5952 11034 6016
rect 10718 5951 11034 5952
rect 2865 5810 2931 5813
rect 3417 5810 3483 5813
rect 2865 5808 3483 5810
rect 2865 5752 2870 5808
rect 2926 5752 3422 5808
rect 3478 5752 3483 5808
rect 2865 5750 3483 5752
rect 2865 5747 2931 5750
rect 3417 5747 3483 5750
rect 0 5538 400 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 400 5478
rect 933 5475 999 5478
rect 3658 5472 3974 5473
rect 3658 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3974 5472
rect 3658 5407 3974 5408
rect 10058 5472 10374 5473
rect 10058 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10374 5472
rect 10058 5407 10374 5408
rect 0 5266 400 5296
rect 1117 5266 1183 5269
rect 0 5264 1183 5266
rect 0 5208 1122 5264
rect 1178 5208 1183 5264
rect 0 5206 1183 5208
rect 0 5176 400 5206
rect 1117 5203 1183 5206
rect 0 4994 400 5024
rect 606 4994 612 4996
rect 0 4934 612 4994
rect 0 4904 400 4934
rect 606 4932 612 4934
rect 676 4932 682 4996
rect 4318 4928 4634 4929
rect 4318 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4634 4928
rect 4318 4863 4634 4864
rect 10718 4928 11034 4929
rect 10718 4864 10724 4928
rect 10788 4864 10804 4928
rect 10868 4864 10884 4928
rect 10948 4864 10964 4928
rect 11028 4864 11034 4928
rect 10718 4863 11034 4864
rect 0 4725 400 4752
rect 0 4720 447 4725
rect 0 4664 386 4720
rect 442 4664 447 4720
rect 0 4659 447 4664
rect 0 4632 400 4659
rect 3658 4384 3974 4385
rect 3658 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3974 4384
rect 3658 4319 3974 4320
rect 10058 4384 10374 4385
rect 10058 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10374 4384
rect 10058 4319 10374 4320
rect 4318 3840 4634 3841
rect 4318 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4634 3840
rect 4318 3775 4634 3776
rect 10718 3840 11034 3841
rect 10718 3776 10724 3840
rect 10788 3776 10804 3840
rect 10868 3776 10884 3840
rect 10948 3776 10964 3840
rect 11028 3776 11034 3840
rect 10718 3775 11034 3776
rect 3658 3296 3974 3297
rect 3658 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3974 3296
rect 3658 3231 3974 3232
rect 10058 3296 10374 3297
rect 10058 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10374 3296
rect 10058 3231 10374 3232
rect 4318 2752 4634 2753
rect 4318 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4634 2752
rect 4318 2687 4634 2688
rect 10718 2752 11034 2753
rect 10718 2688 10724 2752
rect 10788 2688 10804 2752
rect 10868 2688 10884 2752
rect 10948 2688 10964 2752
rect 11028 2688 11034 2752
rect 10718 2687 11034 2688
rect 9806 2484 9812 2548
rect 9876 2546 9882 2548
rect 10041 2546 10107 2549
rect 9876 2544 10107 2546
rect 9876 2488 10046 2544
rect 10102 2488 10107 2544
rect 9876 2486 10107 2488
rect 9876 2484 9882 2486
rect 10041 2483 10107 2486
rect 3658 2208 3974 2209
rect 3658 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3974 2208
rect 3658 2143 3974 2144
rect 10058 2208 10374 2209
rect 10058 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10374 2208
rect 10058 2143 10374 2144
rect 4318 1664 4634 1665
rect 4318 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4634 1664
rect 4318 1599 4634 1600
rect 10718 1664 11034 1665
rect 10718 1600 10724 1664
rect 10788 1600 10804 1664
rect 10868 1600 10884 1664
rect 10948 1600 10964 1664
rect 11028 1600 11034 1664
rect 10718 1599 11034 1600
rect 2497 1458 2563 1461
rect 7373 1458 7439 1461
rect 2497 1456 7439 1458
rect 2497 1400 2502 1456
rect 2558 1400 7378 1456
rect 7434 1400 7439 1456
rect 2497 1398 7439 1400
rect 2497 1395 2563 1398
rect 7373 1395 7439 1398
rect 3658 1120 3974 1121
rect 3658 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3974 1120
rect 3658 1055 3974 1056
rect 10058 1120 10374 1121
rect 10058 1056 10064 1120
rect 10128 1056 10144 1120
rect 10208 1056 10224 1120
rect 10288 1056 10304 1120
rect 10368 1056 10374 1120
rect 10058 1055 10374 1056
rect 4318 576 4634 577
rect 4318 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4634 576
rect 4318 511 4634 512
rect 10718 576 11034 577
rect 10718 512 10724 576
rect 10788 512 10804 576
rect 10868 512 10884 576
rect 10948 512 10964 576
rect 11028 512 11034 576
rect 10718 511 11034 512
<< via3 >>
rect 1348 43556 1412 43620
rect 5396 43556 5460 43620
rect 5580 43556 5644 43620
rect 8156 43556 8220 43620
rect 9260 43556 9324 43620
rect 9628 43556 9692 43620
rect 4324 43004 4388 43008
rect 4324 42948 4328 43004
rect 4328 42948 4384 43004
rect 4384 42948 4388 43004
rect 4324 42944 4388 42948
rect 4404 43004 4468 43008
rect 4404 42948 4408 43004
rect 4408 42948 4464 43004
rect 4464 42948 4468 43004
rect 4404 42944 4468 42948
rect 4484 43004 4548 43008
rect 4484 42948 4488 43004
rect 4488 42948 4544 43004
rect 4544 42948 4548 43004
rect 4484 42944 4548 42948
rect 4564 43004 4628 43008
rect 4564 42948 4568 43004
rect 4568 42948 4624 43004
rect 4624 42948 4628 43004
rect 4564 42944 4628 42948
rect 10724 43004 10788 43008
rect 10724 42948 10728 43004
rect 10728 42948 10784 43004
rect 10784 42948 10788 43004
rect 10724 42944 10788 42948
rect 10804 43004 10868 43008
rect 10804 42948 10808 43004
rect 10808 42948 10864 43004
rect 10864 42948 10868 43004
rect 10804 42944 10868 42948
rect 10884 43004 10948 43008
rect 10884 42948 10888 43004
rect 10888 42948 10944 43004
rect 10944 42948 10948 43004
rect 10884 42944 10948 42948
rect 10964 43004 11028 43008
rect 10964 42948 10968 43004
rect 10968 42948 11024 43004
rect 11024 42948 11028 43004
rect 10964 42944 11028 42948
rect 3664 42460 3728 42464
rect 3664 42404 3668 42460
rect 3668 42404 3724 42460
rect 3724 42404 3728 42460
rect 3664 42400 3728 42404
rect 3744 42460 3808 42464
rect 3744 42404 3748 42460
rect 3748 42404 3804 42460
rect 3804 42404 3808 42460
rect 3744 42400 3808 42404
rect 3824 42460 3888 42464
rect 3824 42404 3828 42460
rect 3828 42404 3884 42460
rect 3884 42404 3888 42460
rect 3824 42400 3888 42404
rect 3904 42460 3968 42464
rect 3904 42404 3908 42460
rect 3908 42404 3964 42460
rect 3964 42404 3968 42460
rect 3904 42400 3968 42404
rect 10064 42460 10128 42464
rect 10064 42404 10068 42460
rect 10068 42404 10124 42460
rect 10124 42404 10128 42460
rect 10064 42400 10128 42404
rect 10144 42460 10208 42464
rect 10144 42404 10148 42460
rect 10148 42404 10204 42460
rect 10204 42404 10208 42460
rect 10144 42400 10208 42404
rect 10224 42460 10288 42464
rect 10224 42404 10228 42460
rect 10228 42404 10284 42460
rect 10284 42404 10288 42460
rect 10224 42400 10288 42404
rect 10304 42460 10368 42464
rect 10304 42404 10308 42460
rect 10308 42404 10364 42460
rect 10364 42404 10368 42460
rect 10304 42400 10368 42404
rect 8708 41924 8772 41988
rect 11468 41924 11532 41988
rect 4324 41916 4388 41920
rect 4324 41860 4328 41916
rect 4328 41860 4384 41916
rect 4384 41860 4388 41916
rect 4324 41856 4388 41860
rect 4404 41916 4468 41920
rect 4404 41860 4408 41916
rect 4408 41860 4464 41916
rect 4464 41860 4468 41916
rect 4404 41856 4468 41860
rect 4484 41916 4548 41920
rect 4484 41860 4488 41916
rect 4488 41860 4544 41916
rect 4544 41860 4548 41916
rect 4484 41856 4548 41860
rect 4564 41916 4628 41920
rect 4564 41860 4568 41916
rect 4568 41860 4624 41916
rect 4624 41860 4628 41916
rect 4564 41856 4628 41860
rect 10724 41916 10788 41920
rect 10724 41860 10728 41916
rect 10728 41860 10784 41916
rect 10784 41860 10788 41916
rect 10724 41856 10788 41860
rect 10804 41916 10868 41920
rect 10804 41860 10808 41916
rect 10808 41860 10864 41916
rect 10864 41860 10868 41916
rect 10804 41856 10868 41860
rect 10884 41916 10948 41920
rect 10884 41860 10888 41916
rect 10888 41860 10944 41916
rect 10944 41860 10948 41916
rect 10884 41856 10948 41860
rect 10964 41916 11028 41920
rect 10964 41860 10968 41916
rect 10968 41860 11024 41916
rect 11024 41860 11028 41916
rect 10964 41856 11028 41860
rect 382 41652 446 41716
rect 9812 41652 9876 41716
rect 3372 41516 3436 41580
rect 6500 41516 6564 41580
rect 11652 41516 11716 41580
rect 3664 41372 3728 41376
rect 3664 41316 3668 41372
rect 3668 41316 3724 41372
rect 3724 41316 3728 41372
rect 3664 41312 3728 41316
rect 3744 41372 3808 41376
rect 3744 41316 3748 41372
rect 3748 41316 3804 41372
rect 3804 41316 3808 41372
rect 3744 41312 3808 41316
rect 3824 41372 3888 41376
rect 3824 41316 3828 41372
rect 3828 41316 3884 41372
rect 3884 41316 3888 41372
rect 3824 41312 3888 41316
rect 3904 41372 3968 41376
rect 3904 41316 3908 41372
rect 3908 41316 3964 41372
rect 3964 41316 3968 41372
rect 3904 41312 3968 41316
rect 10064 41372 10128 41376
rect 10064 41316 10068 41372
rect 10068 41316 10124 41372
rect 10124 41316 10128 41372
rect 10064 41312 10128 41316
rect 10144 41372 10208 41376
rect 10144 41316 10148 41372
rect 10148 41316 10204 41372
rect 10204 41316 10208 41372
rect 10144 41312 10208 41316
rect 10224 41372 10288 41376
rect 10224 41316 10228 41372
rect 10228 41316 10284 41372
rect 10284 41316 10288 41372
rect 10224 41312 10288 41316
rect 10304 41372 10368 41376
rect 10304 41316 10308 41372
rect 10308 41316 10364 41372
rect 10364 41316 10368 41372
rect 10304 41312 10368 41316
rect 7052 41244 7116 41308
rect 1164 40972 1228 41036
rect 8524 40972 8588 41036
rect 4324 40828 4388 40832
rect 4324 40772 4328 40828
rect 4328 40772 4384 40828
rect 4384 40772 4388 40828
rect 4324 40768 4388 40772
rect 4404 40828 4468 40832
rect 4404 40772 4408 40828
rect 4408 40772 4464 40828
rect 4464 40772 4468 40828
rect 4404 40768 4468 40772
rect 4484 40828 4548 40832
rect 4484 40772 4488 40828
rect 4488 40772 4544 40828
rect 4544 40772 4548 40828
rect 4484 40768 4548 40772
rect 4564 40828 4628 40832
rect 4564 40772 4568 40828
rect 4568 40772 4624 40828
rect 4624 40772 4628 40828
rect 4564 40768 4628 40772
rect 10724 40828 10788 40832
rect 10724 40772 10728 40828
rect 10728 40772 10784 40828
rect 10784 40772 10788 40828
rect 10724 40768 10788 40772
rect 10804 40828 10868 40832
rect 10804 40772 10808 40828
rect 10808 40772 10864 40828
rect 10864 40772 10868 40828
rect 10804 40768 10868 40772
rect 10884 40828 10948 40832
rect 10884 40772 10888 40828
rect 10888 40772 10944 40828
rect 10944 40772 10948 40828
rect 10884 40768 10948 40772
rect 10964 40828 11028 40832
rect 10964 40772 10968 40828
rect 10968 40772 11024 40828
rect 11024 40772 11028 40828
rect 10964 40768 11028 40772
rect 5212 40760 5276 40764
rect 5212 40704 5226 40760
rect 5226 40704 5276 40760
rect 5212 40700 5276 40704
rect 7420 40488 7484 40492
rect 7420 40432 7470 40488
rect 7470 40432 7484 40488
rect 7420 40428 7484 40432
rect 3664 40284 3728 40288
rect 3664 40228 3668 40284
rect 3668 40228 3724 40284
rect 3724 40228 3728 40284
rect 3664 40224 3728 40228
rect 3744 40284 3808 40288
rect 3744 40228 3748 40284
rect 3748 40228 3804 40284
rect 3804 40228 3808 40284
rect 3744 40224 3808 40228
rect 3824 40284 3888 40288
rect 3824 40228 3828 40284
rect 3828 40228 3884 40284
rect 3884 40228 3888 40284
rect 3824 40224 3888 40228
rect 3904 40284 3968 40288
rect 3904 40228 3908 40284
rect 3908 40228 3964 40284
rect 3964 40228 3968 40284
rect 3904 40224 3968 40228
rect 10064 40284 10128 40288
rect 10064 40228 10068 40284
rect 10068 40228 10124 40284
rect 10124 40228 10128 40284
rect 10064 40224 10128 40228
rect 10144 40284 10208 40288
rect 10144 40228 10148 40284
rect 10148 40228 10204 40284
rect 10204 40228 10208 40284
rect 10144 40224 10208 40228
rect 10224 40284 10288 40288
rect 10224 40228 10228 40284
rect 10228 40228 10284 40284
rect 10284 40228 10288 40284
rect 10224 40224 10288 40228
rect 10304 40284 10368 40288
rect 10304 40228 10308 40284
rect 10308 40228 10364 40284
rect 10364 40228 10368 40284
rect 10304 40224 10368 40228
rect 3188 40156 3252 40220
rect 5948 40156 6012 40220
rect 10548 40156 10612 40220
rect 4108 40020 4172 40084
rect 5764 40020 5828 40084
rect 8892 40020 8956 40084
rect 11284 40020 11348 40084
rect 2084 39884 2148 39948
rect 5396 39884 5460 39948
rect 4324 39740 4388 39744
rect 4324 39684 4328 39740
rect 4328 39684 4384 39740
rect 4384 39684 4388 39740
rect 4324 39680 4388 39684
rect 4404 39740 4468 39744
rect 4404 39684 4408 39740
rect 4408 39684 4464 39740
rect 4464 39684 4468 39740
rect 4404 39680 4468 39684
rect 4484 39740 4548 39744
rect 4484 39684 4488 39740
rect 4488 39684 4544 39740
rect 4544 39684 4548 39740
rect 4484 39680 4548 39684
rect 4564 39740 4628 39744
rect 4564 39684 4568 39740
rect 4568 39684 4624 39740
rect 4624 39684 4628 39740
rect 4564 39680 4628 39684
rect 10724 39740 10788 39744
rect 10724 39684 10728 39740
rect 10728 39684 10784 39740
rect 10784 39684 10788 39740
rect 10724 39680 10788 39684
rect 10804 39740 10868 39744
rect 10804 39684 10808 39740
rect 10808 39684 10864 39740
rect 10864 39684 10868 39740
rect 10804 39680 10868 39684
rect 10884 39740 10948 39744
rect 10884 39684 10888 39740
rect 10888 39684 10944 39740
rect 10944 39684 10948 39740
rect 10884 39680 10948 39684
rect 10964 39740 11028 39744
rect 10964 39684 10968 39740
rect 10968 39684 11024 39740
rect 11024 39684 11028 39740
rect 10964 39680 11028 39684
rect 7788 39476 7852 39540
rect 4844 39340 4908 39404
rect 5212 39204 5276 39268
rect 3664 39196 3728 39200
rect 3664 39140 3668 39196
rect 3668 39140 3724 39196
rect 3724 39140 3728 39196
rect 3664 39136 3728 39140
rect 3744 39196 3808 39200
rect 3744 39140 3748 39196
rect 3748 39140 3804 39196
rect 3804 39140 3808 39196
rect 3744 39136 3808 39140
rect 3824 39196 3888 39200
rect 3824 39140 3828 39196
rect 3828 39140 3884 39196
rect 3884 39140 3888 39196
rect 3824 39136 3888 39140
rect 3904 39196 3968 39200
rect 3904 39140 3908 39196
rect 3908 39140 3964 39196
rect 3964 39140 3968 39196
rect 3904 39136 3968 39140
rect 10064 39196 10128 39200
rect 10064 39140 10068 39196
rect 10068 39140 10124 39196
rect 10124 39140 10128 39196
rect 10064 39136 10128 39140
rect 10144 39196 10208 39200
rect 10144 39140 10148 39196
rect 10148 39140 10204 39196
rect 10204 39140 10208 39196
rect 10144 39136 10208 39140
rect 10224 39196 10288 39200
rect 10224 39140 10228 39196
rect 10228 39140 10284 39196
rect 10284 39140 10288 39196
rect 10224 39136 10288 39140
rect 10304 39196 10368 39200
rect 10304 39140 10308 39196
rect 10308 39140 10364 39196
rect 10364 39140 10368 39196
rect 10304 39136 10368 39140
rect 1532 38796 1596 38860
rect 7236 38796 7300 38860
rect 9812 38796 9876 38860
rect 12020 38796 12084 38860
rect 4324 38652 4388 38656
rect 4324 38596 4328 38652
rect 4328 38596 4384 38652
rect 4384 38596 4388 38652
rect 4324 38592 4388 38596
rect 4404 38652 4468 38656
rect 4404 38596 4408 38652
rect 4408 38596 4464 38652
rect 4464 38596 4468 38652
rect 4404 38592 4468 38596
rect 4484 38652 4548 38656
rect 4484 38596 4488 38652
rect 4488 38596 4544 38652
rect 4544 38596 4548 38652
rect 4484 38592 4548 38596
rect 4564 38652 4628 38656
rect 4564 38596 4568 38652
rect 4568 38596 4624 38652
rect 4624 38596 4628 38652
rect 4564 38592 4628 38596
rect 1716 38524 1780 38588
rect 9444 38660 9508 38724
rect 10724 38652 10788 38656
rect 10724 38596 10728 38652
rect 10728 38596 10784 38652
rect 10784 38596 10788 38652
rect 10724 38592 10788 38596
rect 10804 38652 10868 38656
rect 10804 38596 10808 38652
rect 10808 38596 10864 38652
rect 10864 38596 10868 38652
rect 10804 38592 10868 38596
rect 10884 38652 10948 38656
rect 10884 38596 10888 38652
rect 10888 38596 10944 38652
rect 10944 38596 10948 38652
rect 10884 38592 10948 38596
rect 10964 38652 11028 38656
rect 10964 38596 10968 38652
rect 10968 38596 11024 38652
rect 11024 38596 11028 38652
rect 10964 38592 11028 38596
rect 6868 38524 6932 38588
rect 7604 38388 7668 38452
rect 1900 38116 1964 38180
rect 6316 38252 6380 38316
rect 10548 38252 10612 38316
rect 11100 38252 11164 38316
rect 3664 38108 3728 38112
rect 3664 38052 3668 38108
rect 3668 38052 3724 38108
rect 3724 38052 3728 38108
rect 3664 38048 3728 38052
rect 3744 38108 3808 38112
rect 3744 38052 3748 38108
rect 3748 38052 3804 38108
rect 3804 38052 3808 38108
rect 3744 38048 3808 38052
rect 3824 38108 3888 38112
rect 3824 38052 3828 38108
rect 3828 38052 3884 38108
rect 3884 38052 3888 38108
rect 3824 38048 3888 38052
rect 3904 38108 3968 38112
rect 3904 38052 3908 38108
rect 3908 38052 3964 38108
rect 3964 38052 3968 38108
rect 3904 38048 3968 38052
rect 10064 38108 10128 38112
rect 10064 38052 10068 38108
rect 10068 38052 10124 38108
rect 10124 38052 10128 38108
rect 10064 38048 10128 38052
rect 10144 38108 10208 38112
rect 10144 38052 10148 38108
rect 10148 38052 10204 38108
rect 10204 38052 10208 38108
rect 10144 38048 10208 38052
rect 10224 38108 10288 38112
rect 10224 38052 10228 38108
rect 10228 38052 10284 38108
rect 10284 38052 10288 38108
rect 10224 38048 10288 38052
rect 10304 38108 10368 38112
rect 10304 38052 10308 38108
rect 10308 38052 10364 38108
rect 10364 38052 10368 38108
rect 10304 38048 10368 38052
rect 6868 37844 6932 37908
rect 8340 37844 8404 37908
rect 9812 37844 9876 37908
rect 2268 37708 2332 37772
rect 980 37572 1044 37636
rect 9076 37572 9140 37636
rect 4324 37564 4388 37568
rect 4324 37508 4328 37564
rect 4328 37508 4384 37564
rect 4384 37508 4388 37564
rect 4324 37504 4388 37508
rect 4404 37564 4468 37568
rect 4404 37508 4408 37564
rect 4408 37508 4464 37564
rect 4464 37508 4468 37564
rect 4404 37504 4468 37508
rect 4484 37564 4548 37568
rect 4484 37508 4488 37564
rect 4488 37508 4544 37564
rect 4544 37508 4548 37564
rect 4484 37504 4548 37508
rect 4564 37564 4628 37568
rect 4564 37508 4568 37564
rect 4568 37508 4624 37564
rect 4624 37508 4628 37564
rect 4564 37504 4628 37508
rect 10724 37564 10788 37568
rect 10724 37508 10728 37564
rect 10728 37508 10784 37564
rect 10784 37508 10788 37564
rect 10724 37504 10788 37508
rect 10804 37564 10868 37568
rect 10804 37508 10808 37564
rect 10808 37508 10864 37564
rect 10864 37508 10868 37564
rect 10804 37504 10868 37508
rect 10884 37564 10948 37568
rect 10884 37508 10888 37564
rect 10888 37508 10944 37564
rect 10944 37508 10948 37564
rect 10884 37504 10948 37508
rect 10964 37564 11028 37568
rect 10964 37508 10968 37564
rect 10968 37508 11024 37564
rect 11024 37508 11028 37564
rect 10964 37504 11028 37508
rect 5212 37496 5276 37500
rect 5212 37440 5226 37496
rect 5226 37440 5276 37496
rect 5212 37436 5276 37440
rect 2636 37300 2700 37364
rect 4108 37300 4172 37364
rect 5580 37300 5644 37364
rect 7972 37300 8036 37364
rect 10548 37300 10612 37364
rect 11836 37300 11900 37364
rect 9812 37164 9876 37228
rect 12204 37164 12268 37228
rect 1900 37028 1964 37092
rect 7604 37028 7668 37092
rect 3664 37020 3728 37024
rect 3664 36964 3668 37020
rect 3668 36964 3724 37020
rect 3724 36964 3728 37020
rect 3664 36960 3728 36964
rect 3744 37020 3808 37024
rect 3744 36964 3748 37020
rect 3748 36964 3804 37020
rect 3804 36964 3808 37020
rect 3744 36960 3808 36964
rect 3824 37020 3888 37024
rect 3824 36964 3828 37020
rect 3828 36964 3884 37020
rect 3884 36964 3888 37020
rect 3824 36960 3888 36964
rect 3904 37020 3968 37024
rect 3904 36964 3908 37020
rect 3908 36964 3964 37020
rect 3964 36964 3968 37020
rect 3904 36960 3968 36964
rect 1348 36892 1412 36956
rect 5028 36816 5092 36820
rect 10064 37020 10128 37024
rect 10064 36964 10068 37020
rect 10068 36964 10124 37020
rect 10124 36964 10128 37020
rect 10064 36960 10128 36964
rect 10144 37020 10208 37024
rect 10144 36964 10148 37020
rect 10148 36964 10204 37020
rect 10204 36964 10208 37020
rect 10144 36960 10208 36964
rect 10224 37020 10288 37024
rect 10224 36964 10228 37020
rect 10228 36964 10284 37020
rect 10284 36964 10288 37020
rect 10224 36960 10288 36964
rect 10304 37020 10368 37024
rect 10304 36964 10308 37020
rect 10308 36964 10364 37020
rect 10364 36964 10368 37020
rect 10304 36960 10368 36964
rect 11100 36892 11164 36956
rect 5028 36760 5042 36816
rect 5042 36760 5092 36816
rect 5028 36756 5092 36760
rect 11100 36816 11164 36820
rect 11100 36760 11150 36816
rect 11150 36760 11164 36816
rect 11100 36756 11164 36760
rect 7052 36484 7116 36548
rect 4324 36476 4388 36480
rect 4324 36420 4328 36476
rect 4328 36420 4384 36476
rect 4384 36420 4388 36476
rect 4324 36416 4388 36420
rect 4404 36476 4468 36480
rect 4404 36420 4408 36476
rect 4408 36420 4464 36476
rect 4464 36420 4468 36476
rect 4404 36416 4468 36420
rect 4484 36476 4548 36480
rect 4484 36420 4488 36476
rect 4488 36420 4544 36476
rect 4544 36420 4548 36476
rect 4484 36416 4548 36420
rect 4564 36476 4628 36480
rect 4564 36420 4568 36476
rect 4568 36420 4624 36476
rect 4624 36420 4628 36476
rect 4564 36416 4628 36420
rect 7788 36076 7852 36140
rect 10724 36476 10788 36480
rect 10724 36420 10728 36476
rect 10728 36420 10784 36476
rect 10784 36420 10788 36476
rect 10724 36416 10788 36420
rect 10804 36476 10868 36480
rect 10804 36420 10808 36476
rect 10808 36420 10864 36476
rect 10864 36420 10868 36476
rect 10804 36416 10868 36420
rect 10884 36476 10948 36480
rect 10884 36420 10888 36476
rect 10888 36420 10944 36476
rect 10944 36420 10948 36476
rect 10884 36416 10948 36420
rect 10964 36476 11028 36480
rect 10964 36420 10968 36476
rect 10968 36420 11024 36476
rect 11024 36420 11028 36476
rect 10964 36416 11028 36420
rect 5580 35940 5644 36004
rect 3664 35932 3728 35936
rect 3664 35876 3668 35932
rect 3668 35876 3724 35932
rect 3724 35876 3728 35932
rect 3664 35872 3728 35876
rect 3744 35932 3808 35936
rect 3744 35876 3748 35932
rect 3748 35876 3804 35932
rect 3804 35876 3808 35932
rect 3744 35872 3808 35876
rect 3824 35932 3888 35936
rect 3824 35876 3828 35932
rect 3828 35876 3884 35932
rect 3884 35876 3888 35932
rect 3824 35872 3888 35876
rect 3904 35932 3968 35936
rect 3904 35876 3908 35932
rect 3908 35876 3964 35932
rect 3964 35876 3968 35932
rect 3904 35872 3968 35876
rect 10064 35932 10128 35936
rect 10064 35876 10068 35932
rect 10068 35876 10124 35932
rect 10124 35876 10128 35932
rect 10064 35872 10128 35876
rect 10144 35932 10208 35936
rect 10144 35876 10148 35932
rect 10148 35876 10204 35932
rect 10204 35876 10208 35932
rect 10144 35872 10208 35876
rect 10224 35932 10288 35936
rect 10224 35876 10228 35932
rect 10228 35876 10284 35932
rect 10284 35876 10288 35932
rect 10224 35872 10288 35876
rect 10304 35932 10368 35936
rect 10304 35876 10308 35932
rect 10308 35876 10364 35932
rect 10364 35876 10368 35932
rect 10304 35872 10368 35876
rect 5764 35864 5828 35868
rect 5764 35808 5814 35864
rect 5814 35808 5828 35864
rect 5764 35804 5828 35808
rect 7604 35532 7668 35596
rect 9812 35532 9876 35596
rect 3372 35396 3436 35460
rect 4324 35388 4388 35392
rect 4324 35332 4328 35388
rect 4328 35332 4384 35388
rect 4384 35332 4388 35388
rect 4324 35328 4388 35332
rect 4404 35388 4468 35392
rect 4404 35332 4408 35388
rect 4408 35332 4464 35388
rect 4464 35332 4468 35388
rect 4404 35328 4468 35332
rect 4484 35388 4548 35392
rect 4484 35332 4488 35388
rect 4488 35332 4544 35388
rect 4544 35332 4548 35388
rect 4484 35328 4548 35332
rect 4564 35388 4628 35392
rect 4564 35332 4568 35388
rect 4568 35332 4624 35388
rect 4624 35332 4628 35388
rect 4564 35328 4628 35332
rect 10724 35388 10788 35392
rect 10724 35332 10728 35388
rect 10728 35332 10784 35388
rect 10784 35332 10788 35388
rect 10724 35328 10788 35332
rect 10804 35388 10868 35392
rect 10804 35332 10808 35388
rect 10808 35332 10864 35388
rect 10864 35332 10868 35388
rect 10804 35328 10868 35332
rect 10884 35388 10948 35392
rect 10884 35332 10888 35388
rect 10888 35332 10944 35388
rect 10944 35332 10948 35388
rect 10884 35328 10948 35332
rect 10964 35388 11028 35392
rect 10964 35332 10968 35388
rect 10968 35332 11024 35388
rect 11024 35332 11028 35388
rect 10964 35328 11028 35332
rect 3004 35260 3068 35324
rect 6868 35260 6932 35324
rect 9444 35260 9508 35324
rect 9812 35260 9876 35324
rect 1900 34988 1964 35052
rect 11100 34988 11164 35052
rect 3664 34844 3728 34848
rect 3664 34788 3668 34844
rect 3668 34788 3724 34844
rect 3724 34788 3728 34844
rect 3664 34784 3728 34788
rect 3744 34844 3808 34848
rect 3744 34788 3748 34844
rect 3748 34788 3804 34844
rect 3804 34788 3808 34844
rect 3744 34784 3808 34788
rect 3824 34844 3888 34848
rect 3824 34788 3828 34844
rect 3828 34788 3884 34844
rect 3884 34788 3888 34844
rect 3824 34784 3888 34788
rect 3904 34844 3968 34848
rect 3904 34788 3908 34844
rect 3908 34788 3964 34844
rect 3964 34788 3968 34844
rect 3904 34784 3968 34788
rect 10064 34844 10128 34848
rect 10064 34788 10068 34844
rect 10068 34788 10124 34844
rect 10124 34788 10128 34844
rect 10064 34784 10128 34788
rect 10144 34844 10208 34848
rect 10144 34788 10148 34844
rect 10148 34788 10204 34844
rect 10204 34788 10208 34844
rect 10144 34784 10208 34788
rect 10224 34844 10288 34848
rect 10224 34788 10228 34844
rect 10228 34788 10284 34844
rect 10284 34788 10288 34844
rect 10224 34784 10288 34788
rect 10304 34844 10368 34848
rect 10304 34788 10308 34844
rect 10308 34788 10364 34844
rect 10364 34788 10368 34844
rect 10304 34784 10368 34788
rect 4844 34580 4908 34644
rect 4108 34444 4172 34508
rect 1164 34308 1228 34372
rect 6868 34308 6932 34372
rect 4324 34300 4388 34304
rect 4324 34244 4328 34300
rect 4328 34244 4384 34300
rect 4384 34244 4388 34300
rect 4324 34240 4388 34244
rect 4404 34300 4468 34304
rect 4404 34244 4408 34300
rect 4408 34244 4464 34300
rect 4464 34244 4468 34300
rect 4404 34240 4468 34244
rect 4484 34300 4548 34304
rect 4484 34244 4488 34300
rect 4488 34244 4544 34300
rect 4544 34244 4548 34300
rect 4484 34240 4548 34244
rect 4564 34300 4628 34304
rect 4564 34244 4568 34300
rect 4568 34244 4624 34300
rect 4624 34244 4628 34300
rect 4564 34240 4628 34244
rect 10724 34300 10788 34304
rect 10724 34244 10728 34300
rect 10728 34244 10784 34300
rect 10784 34244 10788 34300
rect 10724 34240 10788 34244
rect 10804 34300 10868 34304
rect 10804 34244 10808 34300
rect 10808 34244 10864 34300
rect 10864 34244 10868 34300
rect 10804 34240 10868 34244
rect 10884 34300 10948 34304
rect 10884 34244 10888 34300
rect 10888 34244 10944 34300
rect 10944 34244 10948 34300
rect 10884 34240 10948 34244
rect 10964 34300 11028 34304
rect 10964 34244 10968 34300
rect 10968 34244 11024 34300
rect 11024 34244 11028 34300
rect 10964 34240 11028 34244
rect 4108 34172 4172 34236
rect 6868 33900 6932 33964
rect 9260 33764 9324 33828
rect 3664 33756 3728 33760
rect 3664 33700 3668 33756
rect 3668 33700 3724 33756
rect 3724 33700 3728 33756
rect 3664 33696 3728 33700
rect 3744 33756 3808 33760
rect 3744 33700 3748 33756
rect 3748 33700 3804 33756
rect 3804 33700 3808 33756
rect 3744 33696 3808 33700
rect 3824 33756 3888 33760
rect 3824 33700 3828 33756
rect 3828 33700 3884 33756
rect 3884 33700 3888 33756
rect 3824 33696 3888 33700
rect 3904 33756 3968 33760
rect 3904 33700 3908 33756
rect 3908 33700 3964 33756
rect 3964 33700 3968 33756
rect 3904 33696 3968 33700
rect 10064 33756 10128 33760
rect 10064 33700 10068 33756
rect 10068 33700 10124 33756
rect 10124 33700 10128 33756
rect 10064 33696 10128 33700
rect 10144 33756 10208 33760
rect 10144 33700 10148 33756
rect 10148 33700 10204 33756
rect 10204 33700 10208 33756
rect 10144 33696 10208 33700
rect 10224 33756 10288 33760
rect 10224 33700 10228 33756
rect 10228 33700 10284 33756
rect 10284 33700 10288 33756
rect 10224 33696 10288 33700
rect 10304 33756 10368 33760
rect 10304 33700 10308 33756
rect 10308 33700 10364 33756
rect 10364 33700 10368 33756
rect 10304 33696 10368 33700
rect 2084 33628 2148 33692
rect 5212 33628 5276 33692
rect 8340 33628 8404 33692
rect 9260 33628 9324 33692
rect 11836 33688 11900 33692
rect 11836 33632 11886 33688
rect 11886 33632 11900 33688
rect 11836 33628 11900 33632
rect 1532 33492 1596 33556
rect 2084 33356 2148 33420
rect 5212 33492 5276 33556
rect 5764 33492 5828 33556
rect 11836 33492 11900 33556
rect 2820 33356 2884 33420
rect 4844 33356 4908 33420
rect 5948 33356 6012 33420
rect 2452 33220 2516 33284
rect 7788 33220 7852 33284
rect 4324 33212 4388 33216
rect 4324 33156 4328 33212
rect 4328 33156 4384 33212
rect 4384 33156 4388 33212
rect 4324 33152 4388 33156
rect 4404 33212 4468 33216
rect 4404 33156 4408 33212
rect 4408 33156 4464 33212
rect 4464 33156 4468 33212
rect 4404 33152 4468 33156
rect 4484 33212 4548 33216
rect 4484 33156 4488 33212
rect 4488 33156 4544 33212
rect 4544 33156 4548 33212
rect 4484 33152 4548 33156
rect 4564 33212 4628 33216
rect 4564 33156 4568 33212
rect 4568 33156 4624 33212
rect 4624 33156 4628 33212
rect 4564 33152 4628 33156
rect 10724 33212 10788 33216
rect 10724 33156 10728 33212
rect 10728 33156 10784 33212
rect 10784 33156 10788 33212
rect 10724 33152 10788 33156
rect 10804 33212 10868 33216
rect 10804 33156 10808 33212
rect 10808 33156 10864 33212
rect 10864 33156 10868 33212
rect 10804 33152 10868 33156
rect 10884 33212 10948 33216
rect 10884 33156 10888 33212
rect 10888 33156 10944 33212
rect 10944 33156 10948 33212
rect 10884 33152 10948 33156
rect 10964 33212 11028 33216
rect 10964 33156 10968 33212
rect 10968 33156 11024 33212
rect 11024 33156 11028 33212
rect 10964 33152 11028 33156
rect 5396 32872 5460 32876
rect 5396 32816 5410 32872
rect 5410 32816 5460 32872
rect 5396 32812 5460 32816
rect 6868 32676 6932 32740
rect 8340 32676 8404 32740
rect 9444 32676 9508 32740
rect 3664 32668 3728 32672
rect 3664 32612 3668 32668
rect 3668 32612 3724 32668
rect 3724 32612 3728 32668
rect 3664 32608 3728 32612
rect 3744 32668 3808 32672
rect 3744 32612 3748 32668
rect 3748 32612 3804 32668
rect 3804 32612 3808 32668
rect 3744 32608 3808 32612
rect 3824 32668 3888 32672
rect 3824 32612 3828 32668
rect 3828 32612 3884 32668
rect 3884 32612 3888 32668
rect 3824 32608 3888 32612
rect 3904 32668 3968 32672
rect 3904 32612 3908 32668
rect 3908 32612 3964 32668
rect 3964 32612 3968 32668
rect 3904 32608 3968 32612
rect 10064 32668 10128 32672
rect 10064 32612 10068 32668
rect 10068 32612 10124 32668
rect 10124 32612 10128 32668
rect 10064 32608 10128 32612
rect 10144 32668 10208 32672
rect 10144 32612 10148 32668
rect 10148 32612 10204 32668
rect 10204 32612 10208 32668
rect 10144 32608 10208 32612
rect 10224 32668 10288 32672
rect 10224 32612 10228 32668
rect 10228 32612 10284 32668
rect 10284 32612 10288 32668
rect 10224 32608 10288 32612
rect 10304 32668 10368 32672
rect 10304 32612 10308 32668
rect 10308 32612 10364 32668
rect 10364 32612 10368 32668
rect 10304 32608 10368 32612
rect 6500 32540 6564 32604
rect 7236 32540 7300 32604
rect 3188 32404 3252 32468
rect 5396 32404 5460 32468
rect 6132 32404 6196 32468
rect 796 32268 860 32332
rect 1348 32268 1412 32332
rect 6868 32328 6932 32332
rect 6868 32272 6882 32328
rect 6882 32272 6932 32328
rect 6868 32268 6932 32272
rect 1348 32132 1412 32196
rect 7604 32192 7668 32196
rect 7604 32136 7618 32192
rect 7618 32136 7668 32192
rect 7604 32132 7668 32136
rect 10548 32132 10612 32196
rect 4324 32124 4388 32128
rect 4324 32068 4328 32124
rect 4328 32068 4384 32124
rect 4384 32068 4388 32124
rect 4324 32064 4388 32068
rect 4404 32124 4468 32128
rect 4404 32068 4408 32124
rect 4408 32068 4464 32124
rect 4464 32068 4468 32124
rect 4404 32064 4468 32068
rect 4484 32124 4548 32128
rect 4484 32068 4488 32124
rect 4488 32068 4544 32124
rect 4544 32068 4548 32124
rect 4484 32064 4548 32068
rect 4564 32124 4628 32128
rect 4564 32068 4568 32124
rect 4568 32068 4624 32124
rect 4624 32068 4628 32124
rect 4564 32064 4628 32068
rect 10724 32124 10788 32128
rect 10724 32068 10728 32124
rect 10728 32068 10784 32124
rect 10784 32068 10788 32124
rect 10724 32064 10788 32068
rect 10804 32124 10868 32128
rect 10804 32068 10808 32124
rect 10808 32068 10864 32124
rect 10864 32068 10868 32124
rect 10804 32064 10868 32068
rect 10884 32124 10948 32128
rect 10884 32068 10888 32124
rect 10888 32068 10944 32124
rect 10944 32068 10948 32124
rect 10884 32064 10948 32068
rect 10964 32124 11028 32128
rect 10964 32068 10968 32124
rect 10968 32068 11024 32124
rect 11024 32068 11028 32124
rect 10964 32064 11028 32068
rect 2268 31724 2332 31788
rect 7972 31996 8036 32060
rect 7052 31860 7116 31924
rect 10548 31860 10612 31924
rect 11100 31860 11164 31924
rect 5764 31784 5828 31788
rect 5764 31728 5814 31784
rect 5814 31728 5828 31784
rect 5764 31724 5828 31728
rect 6316 31724 6380 31788
rect 8708 31724 8772 31788
rect 1716 31588 1780 31652
rect 3664 31580 3728 31584
rect 3664 31524 3668 31580
rect 3668 31524 3724 31580
rect 3724 31524 3728 31580
rect 3664 31520 3728 31524
rect 3744 31580 3808 31584
rect 3744 31524 3748 31580
rect 3748 31524 3804 31580
rect 3804 31524 3808 31580
rect 3744 31520 3808 31524
rect 3824 31580 3888 31584
rect 3824 31524 3828 31580
rect 3828 31524 3884 31580
rect 3884 31524 3888 31580
rect 3824 31520 3888 31524
rect 3904 31580 3968 31584
rect 3904 31524 3908 31580
rect 3908 31524 3964 31580
rect 3964 31524 3968 31580
rect 3904 31520 3968 31524
rect 1716 31512 1780 31516
rect 1716 31456 1730 31512
rect 1730 31456 1780 31512
rect 1716 31452 1780 31456
rect 4108 31452 4172 31516
rect 5948 31588 6012 31652
rect 7420 31588 7484 31652
rect 11100 31588 11164 31652
rect 10064 31580 10128 31584
rect 10064 31524 10068 31580
rect 10068 31524 10124 31580
rect 10124 31524 10128 31580
rect 10064 31520 10128 31524
rect 10144 31580 10208 31584
rect 10144 31524 10148 31580
rect 10148 31524 10204 31580
rect 10204 31524 10208 31580
rect 10144 31520 10208 31524
rect 10224 31580 10288 31584
rect 10224 31524 10228 31580
rect 10228 31524 10284 31580
rect 10284 31524 10288 31580
rect 10224 31520 10288 31524
rect 10304 31580 10368 31584
rect 10304 31524 10308 31580
rect 10308 31524 10364 31580
rect 10364 31524 10368 31580
rect 10304 31520 10368 31524
rect 4108 31316 4172 31380
rect 3372 31104 3436 31108
rect 3372 31048 3386 31104
rect 3386 31048 3436 31104
rect 3372 31044 3436 31048
rect 8708 31044 8772 31108
rect 9076 31044 9140 31108
rect 4324 31036 4388 31040
rect 4324 30980 4328 31036
rect 4328 30980 4384 31036
rect 4384 30980 4388 31036
rect 4324 30976 4388 30980
rect 4404 31036 4468 31040
rect 4404 30980 4408 31036
rect 4408 30980 4464 31036
rect 4464 30980 4468 31036
rect 4404 30976 4468 30980
rect 4484 31036 4548 31040
rect 4484 30980 4488 31036
rect 4488 30980 4544 31036
rect 4544 30980 4548 31036
rect 4484 30976 4548 30980
rect 4564 31036 4628 31040
rect 4564 30980 4568 31036
rect 4568 30980 4624 31036
rect 4624 30980 4628 31036
rect 4564 30976 4628 30980
rect 10724 31036 10788 31040
rect 10724 30980 10728 31036
rect 10728 30980 10784 31036
rect 10784 30980 10788 31036
rect 10724 30976 10788 30980
rect 10804 31036 10868 31040
rect 10804 30980 10808 31036
rect 10808 30980 10864 31036
rect 10864 30980 10868 31036
rect 10804 30976 10868 30980
rect 10884 31036 10948 31040
rect 10884 30980 10888 31036
rect 10888 30980 10944 31036
rect 10944 30980 10948 31036
rect 10884 30976 10948 30980
rect 10964 31036 11028 31040
rect 10964 30980 10968 31036
rect 10968 30980 11024 31036
rect 11024 30980 11028 31036
rect 10964 30976 11028 30980
rect 9260 30908 9324 30972
rect 5764 30772 5828 30836
rect 7420 30636 7484 30700
rect 9076 30636 9140 30700
rect 5028 30500 5092 30564
rect 9260 30500 9324 30564
rect 3664 30492 3728 30496
rect 3664 30436 3668 30492
rect 3668 30436 3724 30492
rect 3724 30436 3728 30492
rect 3664 30432 3728 30436
rect 3744 30492 3808 30496
rect 3744 30436 3748 30492
rect 3748 30436 3804 30492
rect 3804 30436 3808 30492
rect 3744 30432 3808 30436
rect 3824 30492 3888 30496
rect 3824 30436 3828 30492
rect 3828 30436 3884 30492
rect 3884 30436 3888 30492
rect 3824 30432 3888 30436
rect 3904 30492 3968 30496
rect 3904 30436 3908 30492
rect 3908 30436 3964 30492
rect 3964 30436 3968 30492
rect 3904 30432 3968 30436
rect 10064 30492 10128 30496
rect 10064 30436 10068 30492
rect 10068 30436 10124 30492
rect 10124 30436 10128 30492
rect 10064 30432 10128 30436
rect 10144 30492 10208 30496
rect 10144 30436 10148 30492
rect 10148 30436 10204 30492
rect 10204 30436 10208 30492
rect 10144 30432 10208 30436
rect 10224 30492 10288 30496
rect 10224 30436 10228 30492
rect 10228 30436 10284 30492
rect 10284 30436 10288 30492
rect 10224 30432 10288 30436
rect 10304 30492 10368 30496
rect 10304 30436 10308 30492
rect 10308 30436 10364 30492
rect 10364 30436 10368 30492
rect 10304 30432 10368 30436
rect 2268 30364 2332 30428
rect 5580 30364 5644 30428
rect 6868 30364 6932 30428
rect 7604 30424 7668 30428
rect 7604 30368 7618 30424
rect 7618 30368 7668 30424
rect 7604 30364 7668 30368
rect 8524 30364 8588 30428
rect 5028 30228 5092 30292
rect 8156 30288 8220 30292
rect 8156 30232 8170 30288
rect 8170 30232 8220 30288
rect 8156 30228 8220 30232
rect 9812 30228 9876 30292
rect 1900 29820 1964 29884
rect 3372 29956 3436 30020
rect 5948 30092 6012 30156
rect 6316 30092 6380 30156
rect 7788 30092 7852 30156
rect 11652 30364 11716 30428
rect 11468 30288 11532 30292
rect 11468 30232 11482 30288
rect 11482 30232 11532 30288
rect 11468 30228 11532 30232
rect 4324 29948 4388 29952
rect 4324 29892 4328 29948
rect 4328 29892 4384 29948
rect 4384 29892 4388 29948
rect 4324 29888 4388 29892
rect 4404 29948 4468 29952
rect 4404 29892 4408 29948
rect 4408 29892 4464 29948
rect 4464 29892 4468 29948
rect 4404 29888 4468 29892
rect 4484 29948 4548 29952
rect 4484 29892 4488 29948
rect 4488 29892 4544 29948
rect 4544 29892 4548 29948
rect 4484 29888 4548 29892
rect 4564 29948 4628 29952
rect 4564 29892 4568 29948
rect 4568 29892 4624 29948
rect 4624 29892 4628 29948
rect 4564 29888 4628 29892
rect 60 29684 124 29748
rect 2268 29548 2332 29612
rect 6684 29956 6748 30020
rect 5212 29820 5276 29884
rect 10724 29948 10788 29952
rect 10724 29892 10728 29948
rect 10728 29892 10784 29948
rect 10784 29892 10788 29948
rect 10724 29888 10788 29892
rect 10804 29948 10868 29952
rect 10804 29892 10808 29948
rect 10808 29892 10864 29948
rect 10864 29892 10868 29948
rect 10804 29888 10868 29892
rect 10884 29948 10948 29952
rect 10884 29892 10888 29948
rect 10888 29892 10944 29948
rect 10944 29892 10948 29948
rect 10884 29888 10948 29892
rect 10964 29948 11028 29952
rect 10964 29892 10968 29948
rect 10968 29892 11024 29948
rect 11024 29892 11028 29948
rect 10964 29888 11028 29892
rect 12020 29684 12084 29748
rect 10548 29472 10612 29476
rect 10548 29416 10598 29472
rect 10598 29416 10612 29472
rect 10548 29412 10612 29416
rect 12204 29412 12268 29476
rect 3664 29404 3728 29408
rect 3664 29348 3668 29404
rect 3668 29348 3724 29404
rect 3724 29348 3728 29404
rect 3664 29344 3728 29348
rect 3744 29404 3808 29408
rect 3744 29348 3748 29404
rect 3748 29348 3804 29404
rect 3804 29348 3808 29404
rect 3744 29344 3808 29348
rect 3824 29404 3888 29408
rect 3824 29348 3828 29404
rect 3828 29348 3884 29404
rect 3884 29348 3888 29404
rect 3824 29344 3888 29348
rect 3904 29404 3968 29408
rect 3904 29348 3908 29404
rect 3908 29348 3964 29404
rect 3964 29348 3968 29404
rect 3904 29344 3968 29348
rect 10064 29404 10128 29408
rect 10064 29348 10068 29404
rect 10068 29348 10124 29404
rect 10124 29348 10128 29404
rect 10064 29344 10128 29348
rect 10144 29404 10208 29408
rect 10144 29348 10148 29404
rect 10148 29348 10204 29404
rect 10204 29348 10208 29404
rect 10144 29344 10208 29348
rect 10224 29404 10288 29408
rect 10224 29348 10228 29404
rect 10228 29348 10284 29404
rect 10284 29348 10288 29404
rect 10224 29344 10288 29348
rect 10304 29404 10368 29408
rect 10304 29348 10308 29404
rect 10308 29348 10364 29404
rect 10364 29348 10368 29404
rect 10304 29344 10368 29348
rect 2820 29336 2884 29340
rect 2820 29280 2870 29336
rect 2870 29280 2884 29336
rect 2820 29276 2884 29280
rect 11284 29276 11348 29340
rect 980 29140 1044 29204
rect 2636 29200 2700 29204
rect 2636 29144 2686 29200
rect 2686 29144 2700 29200
rect 2636 29140 2700 29144
rect 7052 29140 7116 29204
rect 3004 28868 3068 28932
rect 6500 29064 6564 29068
rect 6500 29008 6514 29064
rect 6514 29008 6564 29064
rect 6500 29004 6564 29008
rect 5212 28868 5276 28932
rect 7420 28868 7484 28932
rect 7972 28868 8036 28932
rect 4324 28860 4388 28864
rect 4324 28804 4328 28860
rect 4328 28804 4384 28860
rect 4384 28804 4388 28860
rect 4324 28800 4388 28804
rect 4404 28860 4468 28864
rect 4404 28804 4408 28860
rect 4408 28804 4464 28860
rect 4464 28804 4468 28860
rect 4404 28800 4468 28804
rect 4484 28860 4548 28864
rect 4484 28804 4488 28860
rect 4488 28804 4544 28860
rect 4544 28804 4548 28860
rect 4484 28800 4548 28804
rect 4564 28860 4628 28864
rect 4564 28804 4568 28860
rect 4568 28804 4624 28860
rect 4624 28804 4628 28860
rect 4564 28800 4628 28804
rect 10724 28860 10788 28864
rect 10724 28804 10728 28860
rect 10728 28804 10784 28860
rect 10784 28804 10788 28860
rect 10724 28800 10788 28804
rect 10804 28860 10868 28864
rect 10804 28804 10808 28860
rect 10808 28804 10864 28860
rect 10864 28804 10868 28860
rect 10804 28800 10868 28804
rect 10884 28860 10948 28864
rect 10884 28804 10888 28860
rect 10888 28804 10944 28860
rect 10944 28804 10948 28860
rect 10884 28800 10948 28804
rect 10964 28860 11028 28864
rect 10964 28804 10968 28860
rect 10968 28804 11024 28860
rect 11024 28804 11028 28860
rect 10964 28800 11028 28804
rect 5396 28732 5460 28796
rect 5580 28732 5644 28796
rect 8892 28596 8956 28660
rect 1716 28460 1780 28524
rect 9076 28460 9140 28524
rect 11284 28460 11348 28524
rect 7052 28324 7116 28388
rect 3664 28316 3728 28320
rect 3664 28260 3668 28316
rect 3668 28260 3724 28316
rect 3724 28260 3728 28316
rect 3664 28256 3728 28260
rect 3744 28316 3808 28320
rect 3744 28260 3748 28316
rect 3748 28260 3804 28316
rect 3804 28260 3808 28316
rect 3744 28256 3808 28260
rect 3824 28316 3888 28320
rect 3824 28260 3828 28316
rect 3828 28260 3884 28316
rect 3884 28260 3888 28316
rect 3824 28256 3888 28260
rect 3904 28316 3968 28320
rect 3904 28260 3908 28316
rect 3908 28260 3964 28316
rect 3964 28260 3968 28316
rect 3904 28256 3968 28260
rect 10064 28316 10128 28320
rect 10064 28260 10068 28316
rect 10068 28260 10124 28316
rect 10124 28260 10128 28316
rect 10064 28256 10128 28260
rect 10144 28316 10208 28320
rect 10144 28260 10148 28316
rect 10148 28260 10204 28316
rect 10204 28260 10208 28316
rect 10144 28256 10208 28260
rect 10224 28316 10288 28320
rect 10224 28260 10228 28316
rect 10228 28260 10284 28316
rect 10284 28260 10288 28316
rect 10224 28256 10288 28260
rect 10304 28316 10368 28320
rect 10304 28260 10308 28316
rect 10308 28260 10364 28316
rect 10364 28260 10368 28316
rect 10304 28256 10368 28260
rect 612 28188 676 28252
rect 6684 28052 6748 28116
rect 6868 28052 6932 28116
rect 7788 28052 7852 28116
rect 8156 27916 8220 27980
rect 8524 27916 8588 27980
rect 11100 27916 11164 27980
rect 1716 27780 1780 27844
rect 8340 27780 8404 27844
rect 4324 27772 4388 27776
rect 4324 27716 4328 27772
rect 4328 27716 4384 27772
rect 4384 27716 4388 27772
rect 4324 27712 4388 27716
rect 4404 27772 4468 27776
rect 4404 27716 4408 27772
rect 4408 27716 4464 27772
rect 4464 27716 4468 27772
rect 4404 27712 4468 27716
rect 4484 27772 4548 27776
rect 4484 27716 4488 27772
rect 4488 27716 4544 27772
rect 4544 27716 4548 27772
rect 4484 27712 4548 27716
rect 4564 27772 4628 27776
rect 4564 27716 4568 27772
rect 4568 27716 4624 27772
rect 4624 27716 4628 27772
rect 4564 27712 4628 27716
rect 10724 27772 10788 27776
rect 10724 27716 10728 27772
rect 10728 27716 10784 27772
rect 10784 27716 10788 27772
rect 10724 27712 10788 27716
rect 10804 27772 10868 27776
rect 10804 27716 10808 27772
rect 10808 27716 10864 27772
rect 10864 27716 10868 27772
rect 10804 27712 10868 27716
rect 10884 27772 10948 27776
rect 10884 27716 10888 27772
rect 10888 27716 10944 27772
rect 10944 27716 10948 27772
rect 10884 27712 10948 27716
rect 10964 27772 11028 27776
rect 10964 27716 10968 27772
rect 10968 27716 11024 27772
rect 11024 27716 11028 27772
rect 10964 27712 11028 27716
rect 2268 27644 2332 27708
rect 2452 27644 2516 27708
rect 6132 27644 6196 27708
rect 11652 27644 11716 27708
rect 7604 27508 7668 27572
rect 8892 27508 8956 27572
rect 6684 27432 6748 27436
rect 6684 27376 6734 27432
rect 6734 27376 6748 27432
rect 6684 27372 6748 27376
rect 10548 27372 10612 27436
rect 3664 27228 3728 27232
rect 3664 27172 3668 27228
rect 3668 27172 3724 27228
rect 3724 27172 3728 27228
rect 3664 27168 3728 27172
rect 3744 27228 3808 27232
rect 3744 27172 3748 27228
rect 3748 27172 3804 27228
rect 3804 27172 3808 27228
rect 3744 27168 3808 27172
rect 3824 27228 3888 27232
rect 3824 27172 3828 27228
rect 3828 27172 3884 27228
rect 3884 27172 3888 27228
rect 3824 27168 3888 27172
rect 3904 27228 3968 27232
rect 3904 27172 3908 27228
rect 3908 27172 3964 27228
rect 3964 27172 3968 27228
rect 3904 27168 3968 27172
rect 10064 27228 10128 27232
rect 10064 27172 10068 27228
rect 10068 27172 10124 27228
rect 10124 27172 10128 27228
rect 10064 27168 10128 27172
rect 10144 27228 10208 27232
rect 10144 27172 10148 27228
rect 10148 27172 10204 27228
rect 10204 27172 10208 27228
rect 10144 27168 10208 27172
rect 10224 27228 10288 27232
rect 10224 27172 10228 27228
rect 10228 27172 10284 27228
rect 10284 27172 10288 27228
rect 10224 27168 10288 27172
rect 10304 27228 10368 27232
rect 10304 27172 10308 27228
rect 10308 27172 10364 27228
rect 10364 27172 10368 27228
rect 10304 27168 10368 27172
rect 9628 27160 9692 27164
rect 9628 27104 9678 27160
rect 9678 27104 9692 27160
rect 9628 27100 9692 27104
rect 5396 26828 5460 26892
rect 4324 26684 4388 26688
rect 4324 26628 4328 26684
rect 4328 26628 4384 26684
rect 4384 26628 4388 26684
rect 4324 26624 4388 26628
rect 4404 26684 4468 26688
rect 4404 26628 4408 26684
rect 4408 26628 4464 26684
rect 4464 26628 4468 26684
rect 4404 26624 4468 26628
rect 4484 26684 4548 26688
rect 4484 26628 4488 26684
rect 4488 26628 4544 26684
rect 4544 26628 4548 26684
rect 4484 26624 4548 26628
rect 4564 26684 4628 26688
rect 4564 26628 4568 26684
rect 4568 26628 4624 26684
rect 4624 26628 4628 26684
rect 4564 26624 4628 26628
rect 10724 26684 10788 26688
rect 10724 26628 10728 26684
rect 10728 26628 10784 26684
rect 10784 26628 10788 26684
rect 10724 26624 10788 26628
rect 10804 26684 10868 26688
rect 10804 26628 10808 26684
rect 10808 26628 10864 26684
rect 10864 26628 10868 26684
rect 10804 26624 10868 26628
rect 10884 26684 10948 26688
rect 10884 26628 10888 26684
rect 10888 26628 10944 26684
rect 10944 26628 10948 26684
rect 10884 26624 10948 26628
rect 10964 26684 11028 26688
rect 10964 26628 10968 26684
rect 10968 26628 11024 26684
rect 11024 26628 11028 26684
rect 10964 26624 11028 26628
rect 2084 26616 2148 26620
rect 2084 26560 2134 26616
rect 2134 26560 2148 26616
rect 2084 26556 2148 26560
rect 7052 26420 7116 26484
rect 9628 26420 9692 26484
rect 2084 26344 2148 26348
rect 2084 26288 2098 26344
rect 2098 26288 2148 26344
rect 2084 26284 2148 26288
rect 8156 26284 8220 26348
rect 9812 26284 9876 26348
rect 3664 26140 3728 26144
rect 3664 26084 3668 26140
rect 3668 26084 3724 26140
rect 3724 26084 3728 26140
rect 3664 26080 3728 26084
rect 3744 26140 3808 26144
rect 3744 26084 3748 26140
rect 3748 26084 3804 26140
rect 3804 26084 3808 26140
rect 3744 26080 3808 26084
rect 3824 26140 3888 26144
rect 3824 26084 3828 26140
rect 3828 26084 3884 26140
rect 3884 26084 3888 26140
rect 3824 26080 3888 26084
rect 3904 26140 3968 26144
rect 3904 26084 3908 26140
rect 3908 26084 3964 26140
rect 3964 26084 3968 26140
rect 3904 26080 3968 26084
rect 10064 26140 10128 26144
rect 10064 26084 10068 26140
rect 10068 26084 10124 26140
rect 10124 26084 10128 26140
rect 10064 26080 10128 26084
rect 10144 26140 10208 26144
rect 10144 26084 10148 26140
rect 10148 26084 10204 26140
rect 10204 26084 10208 26140
rect 10144 26080 10208 26084
rect 10224 26140 10288 26144
rect 10224 26084 10228 26140
rect 10228 26084 10284 26140
rect 10284 26084 10288 26140
rect 10224 26080 10288 26084
rect 10304 26140 10368 26144
rect 10304 26084 10308 26140
rect 10308 26084 10364 26140
rect 10364 26084 10368 26140
rect 10304 26080 10368 26084
rect 6316 26012 6380 26076
rect 9444 26012 9508 26076
rect 3372 25876 3436 25940
rect 7052 25664 7116 25668
rect 7052 25608 7066 25664
rect 7066 25608 7116 25664
rect 7052 25604 7116 25608
rect 4324 25596 4388 25600
rect 4324 25540 4328 25596
rect 4328 25540 4384 25596
rect 4384 25540 4388 25596
rect 4324 25536 4388 25540
rect 4404 25596 4468 25600
rect 4404 25540 4408 25596
rect 4408 25540 4464 25596
rect 4464 25540 4468 25596
rect 4404 25536 4468 25540
rect 4484 25596 4548 25600
rect 4484 25540 4488 25596
rect 4488 25540 4544 25596
rect 4544 25540 4548 25596
rect 4484 25536 4548 25540
rect 4564 25596 4628 25600
rect 4564 25540 4568 25596
rect 4568 25540 4624 25596
rect 4624 25540 4628 25596
rect 4564 25536 4628 25540
rect 10724 25596 10788 25600
rect 10724 25540 10728 25596
rect 10728 25540 10784 25596
rect 10784 25540 10788 25596
rect 10724 25536 10788 25540
rect 10804 25596 10868 25600
rect 10804 25540 10808 25596
rect 10808 25540 10864 25596
rect 10864 25540 10868 25596
rect 10804 25536 10868 25540
rect 10884 25596 10948 25600
rect 10884 25540 10888 25596
rect 10888 25540 10944 25596
rect 10944 25540 10948 25596
rect 10884 25536 10948 25540
rect 10964 25596 11028 25600
rect 10964 25540 10968 25596
rect 10968 25540 11024 25596
rect 11024 25540 11028 25596
rect 10964 25536 11028 25540
rect 2452 25468 2516 25532
rect 1164 25332 1228 25396
rect 5580 25332 5644 25396
rect 4844 25196 4908 25260
rect 3664 25052 3728 25056
rect 3664 24996 3668 25052
rect 3668 24996 3724 25052
rect 3724 24996 3728 25052
rect 3664 24992 3728 24996
rect 3744 25052 3808 25056
rect 3744 24996 3748 25052
rect 3748 24996 3804 25052
rect 3804 24996 3808 25052
rect 3744 24992 3808 24996
rect 3824 25052 3888 25056
rect 3824 24996 3828 25052
rect 3828 24996 3884 25052
rect 3884 24996 3888 25052
rect 3824 24992 3888 24996
rect 3904 25052 3968 25056
rect 3904 24996 3908 25052
rect 3908 24996 3964 25052
rect 3964 24996 3968 25052
rect 3904 24992 3968 24996
rect 10064 25052 10128 25056
rect 10064 24996 10068 25052
rect 10068 24996 10124 25052
rect 10124 24996 10128 25052
rect 10064 24992 10128 24996
rect 10144 25052 10208 25056
rect 10144 24996 10148 25052
rect 10148 24996 10204 25052
rect 10204 24996 10208 25052
rect 10144 24992 10208 24996
rect 10224 25052 10288 25056
rect 10224 24996 10228 25052
rect 10228 24996 10284 25052
rect 10284 24996 10288 25052
rect 10224 24992 10288 24996
rect 10304 25052 10368 25056
rect 10304 24996 10308 25052
rect 10308 24996 10364 25052
rect 10364 24996 10368 25052
rect 10304 24992 10368 24996
rect 5764 24924 5828 24988
rect 9260 24652 9324 24716
rect 3372 24516 3436 24580
rect 5764 24576 5828 24580
rect 5764 24520 5778 24576
rect 5778 24520 5828 24576
rect 5764 24516 5828 24520
rect 9076 24516 9140 24580
rect 11836 24924 11900 24988
rect 4324 24508 4388 24512
rect 4324 24452 4328 24508
rect 4328 24452 4384 24508
rect 4384 24452 4388 24508
rect 4324 24448 4388 24452
rect 4404 24508 4468 24512
rect 4404 24452 4408 24508
rect 4408 24452 4464 24508
rect 4464 24452 4468 24508
rect 4404 24448 4468 24452
rect 4484 24508 4548 24512
rect 4484 24452 4488 24508
rect 4488 24452 4544 24508
rect 4544 24452 4548 24508
rect 4484 24448 4548 24452
rect 4564 24508 4628 24512
rect 4564 24452 4568 24508
rect 4568 24452 4624 24508
rect 4624 24452 4628 24508
rect 4564 24448 4628 24452
rect 10724 24508 10788 24512
rect 10724 24452 10728 24508
rect 10728 24452 10784 24508
rect 10784 24452 10788 24508
rect 10724 24448 10788 24452
rect 10804 24508 10868 24512
rect 10804 24452 10808 24508
rect 10808 24452 10864 24508
rect 10864 24452 10868 24508
rect 10804 24448 10868 24452
rect 10884 24508 10948 24512
rect 10884 24452 10888 24508
rect 10888 24452 10944 24508
rect 10944 24452 10948 24508
rect 10884 24448 10948 24452
rect 10964 24508 11028 24512
rect 10964 24452 10968 24508
rect 10968 24452 11024 24508
rect 11024 24452 11028 24508
rect 10964 24448 11028 24452
rect 1900 24108 1964 24172
rect 3664 23964 3728 23968
rect 3664 23908 3668 23964
rect 3668 23908 3724 23964
rect 3724 23908 3728 23964
rect 3664 23904 3728 23908
rect 3744 23964 3808 23968
rect 3744 23908 3748 23964
rect 3748 23908 3804 23964
rect 3804 23908 3808 23964
rect 3744 23904 3808 23908
rect 3824 23964 3888 23968
rect 3824 23908 3828 23964
rect 3828 23908 3884 23964
rect 3884 23908 3888 23964
rect 3824 23904 3888 23908
rect 3904 23964 3968 23968
rect 3904 23908 3908 23964
rect 3908 23908 3964 23964
rect 3964 23908 3968 23964
rect 3904 23904 3968 23908
rect 10064 23964 10128 23968
rect 10064 23908 10068 23964
rect 10068 23908 10124 23964
rect 10124 23908 10128 23964
rect 10064 23904 10128 23908
rect 10144 23964 10208 23968
rect 10144 23908 10148 23964
rect 10148 23908 10204 23964
rect 10204 23908 10208 23964
rect 10144 23904 10208 23908
rect 10224 23964 10288 23968
rect 10224 23908 10228 23964
rect 10228 23908 10284 23964
rect 10284 23908 10288 23964
rect 10224 23904 10288 23908
rect 10304 23964 10368 23968
rect 10304 23908 10308 23964
rect 10308 23908 10364 23964
rect 10364 23908 10368 23964
rect 10304 23904 10368 23908
rect 1348 23836 1412 23900
rect 2636 23700 2700 23764
rect 4108 23700 4172 23764
rect 6868 23700 6932 23764
rect 7420 23700 7484 23764
rect 4108 23564 4172 23628
rect 6684 23428 6748 23492
rect 11468 23488 11532 23492
rect 11468 23432 11482 23488
rect 11482 23432 11532 23488
rect 11468 23428 11532 23432
rect 11836 23428 11900 23492
rect 12020 23428 12084 23492
rect 4324 23420 4388 23424
rect 4324 23364 4328 23420
rect 4328 23364 4384 23420
rect 4384 23364 4388 23420
rect 4324 23360 4388 23364
rect 4404 23420 4468 23424
rect 4404 23364 4408 23420
rect 4408 23364 4464 23420
rect 4464 23364 4468 23420
rect 4404 23360 4468 23364
rect 4484 23420 4548 23424
rect 4484 23364 4488 23420
rect 4488 23364 4544 23420
rect 4544 23364 4548 23420
rect 4484 23360 4548 23364
rect 4564 23420 4628 23424
rect 4564 23364 4568 23420
rect 4568 23364 4624 23420
rect 4624 23364 4628 23420
rect 4564 23360 4628 23364
rect 10724 23420 10788 23424
rect 10724 23364 10728 23420
rect 10728 23364 10784 23420
rect 10784 23364 10788 23420
rect 10724 23360 10788 23364
rect 10804 23420 10868 23424
rect 10804 23364 10808 23420
rect 10808 23364 10864 23420
rect 10864 23364 10868 23420
rect 10804 23360 10868 23364
rect 10884 23420 10948 23424
rect 10884 23364 10888 23420
rect 10888 23364 10944 23420
rect 10944 23364 10948 23420
rect 10884 23360 10948 23364
rect 10964 23420 11028 23424
rect 10964 23364 10968 23420
rect 10968 23364 11024 23420
rect 11024 23364 11028 23420
rect 10964 23360 11028 23364
rect 2268 23352 2332 23356
rect 2268 23296 2318 23352
rect 2318 23296 2332 23352
rect 2268 23292 2332 23296
rect 7972 23292 8036 23356
rect 3188 23020 3252 23084
rect 7972 23020 8036 23084
rect 3664 22876 3728 22880
rect 3664 22820 3668 22876
rect 3668 22820 3724 22876
rect 3724 22820 3728 22876
rect 3664 22816 3728 22820
rect 3744 22876 3808 22880
rect 3744 22820 3748 22876
rect 3748 22820 3804 22876
rect 3804 22820 3808 22876
rect 3744 22816 3808 22820
rect 3824 22876 3888 22880
rect 3824 22820 3828 22876
rect 3828 22820 3884 22876
rect 3884 22820 3888 22876
rect 3824 22816 3888 22820
rect 3904 22876 3968 22880
rect 3904 22820 3908 22876
rect 3908 22820 3964 22876
rect 3964 22820 3968 22876
rect 3904 22816 3968 22820
rect 10064 22876 10128 22880
rect 10064 22820 10068 22876
rect 10068 22820 10124 22876
rect 10124 22820 10128 22876
rect 10064 22816 10128 22820
rect 10144 22876 10208 22880
rect 10144 22820 10148 22876
rect 10148 22820 10204 22876
rect 10204 22820 10208 22876
rect 10144 22816 10208 22820
rect 10224 22876 10288 22880
rect 10224 22820 10228 22876
rect 10228 22820 10284 22876
rect 10284 22820 10288 22876
rect 10224 22816 10288 22820
rect 10304 22876 10368 22880
rect 10304 22820 10308 22876
rect 10308 22820 10364 22876
rect 10364 22820 10368 22876
rect 10304 22816 10368 22820
rect 4844 22748 4908 22812
rect 3004 22612 3068 22676
rect 9444 22612 9508 22676
rect 12572 23020 12636 23084
rect 5028 22476 5092 22540
rect 4324 22332 4388 22336
rect 4324 22276 4328 22332
rect 4328 22276 4384 22332
rect 4384 22276 4388 22332
rect 4324 22272 4388 22276
rect 4404 22332 4468 22336
rect 4404 22276 4408 22332
rect 4408 22276 4464 22332
rect 4464 22276 4468 22332
rect 4404 22272 4468 22276
rect 4484 22332 4548 22336
rect 4484 22276 4488 22332
rect 4488 22276 4544 22332
rect 4544 22276 4548 22332
rect 4484 22272 4548 22276
rect 4564 22332 4628 22336
rect 4564 22276 4568 22332
rect 4568 22276 4624 22332
rect 4624 22276 4628 22332
rect 4564 22272 4628 22276
rect 10724 22332 10788 22336
rect 10724 22276 10728 22332
rect 10728 22276 10784 22332
rect 10784 22276 10788 22332
rect 10724 22272 10788 22276
rect 10804 22332 10868 22336
rect 10804 22276 10808 22332
rect 10808 22276 10864 22332
rect 10864 22276 10868 22332
rect 10804 22272 10868 22276
rect 10884 22332 10948 22336
rect 10884 22276 10888 22332
rect 10888 22276 10944 22332
rect 10944 22276 10948 22332
rect 10884 22272 10948 22276
rect 10964 22332 11028 22336
rect 10964 22276 10968 22332
rect 10968 22276 11024 22332
rect 11024 22276 11028 22332
rect 10964 22272 11028 22276
rect 5028 22264 5092 22268
rect 5028 22208 5042 22264
rect 5042 22208 5092 22264
rect 5028 22204 5092 22208
rect 7420 22204 7484 22268
rect 2820 22068 2884 22132
rect 4108 22068 4172 22132
rect 6868 21932 6932 21996
rect 8340 21932 8404 21996
rect 9812 21932 9876 21996
rect 5948 21796 6012 21860
rect 7972 21796 8036 21860
rect 3664 21788 3728 21792
rect 3664 21732 3668 21788
rect 3668 21732 3724 21788
rect 3724 21732 3728 21788
rect 3664 21728 3728 21732
rect 3744 21788 3808 21792
rect 3744 21732 3748 21788
rect 3748 21732 3804 21788
rect 3804 21732 3808 21788
rect 3744 21728 3808 21732
rect 3824 21788 3888 21792
rect 3824 21732 3828 21788
rect 3828 21732 3884 21788
rect 3884 21732 3888 21788
rect 3824 21728 3888 21732
rect 3904 21788 3968 21792
rect 3904 21732 3908 21788
rect 3908 21732 3964 21788
rect 3964 21732 3968 21788
rect 3904 21728 3968 21732
rect 10064 21788 10128 21792
rect 10064 21732 10068 21788
rect 10068 21732 10124 21788
rect 10124 21732 10128 21788
rect 10064 21728 10128 21732
rect 10144 21788 10208 21792
rect 10144 21732 10148 21788
rect 10148 21732 10204 21788
rect 10204 21732 10208 21788
rect 10144 21728 10208 21732
rect 10224 21788 10288 21792
rect 10224 21732 10228 21788
rect 10228 21732 10284 21788
rect 10284 21732 10288 21788
rect 10224 21728 10288 21732
rect 10304 21788 10368 21792
rect 10304 21732 10308 21788
rect 10308 21732 10364 21788
rect 10364 21732 10368 21788
rect 10304 21728 10368 21732
rect 3188 21524 3252 21588
rect 3004 21388 3068 21452
rect 3188 21116 3252 21180
rect 5396 21388 5460 21452
rect 10548 21252 10612 21316
rect 4324 21244 4388 21248
rect 4324 21188 4328 21244
rect 4328 21188 4384 21244
rect 4384 21188 4388 21244
rect 4324 21184 4388 21188
rect 4404 21244 4468 21248
rect 4404 21188 4408 21244
rect 4408 21188 4464 21244
rect 4464 21188 4468 21244
rect 4404 21184 4468 21188
rect 4484 21244 4548 21248
rect 4484 21188 4488 21244
rect 4488 21188 4544 21244
rect 4544 21188 4548 21244
rect 4484 21184 4548 21188
rect 4564 21244 4628 21248
rect 4564 21188 4568 21244
rect 4568 21188 4624 21244
rect 4624 21188 4628 21244
rect 4564 21184 4628 21188
rect 10724 21244 10788 21248
rect 10724 21188 10728 21244
rect 10728 21188 10784 21244
rect 10784 21188 10788 21244
rect 10724 21184 10788 21188
rect 10804 21244 10868 21248
rect 10804 21188 10808 21244
rect 10808 21188 10864 21244
rect 10864 21188 10868 21244
rect 10804 21184 10868 21188
rect 10884 21244 10948 21248
rect 10884 21188 10888 21244
rect 10888 21188 10944 21244
rect 10944 21188 10948 21244
rect 10884 21184 10948 21188
rect 10964 21244 11028 21248
rect 10964 21188 10968 21244
rect 10968 21188 11024 21244
rect 11024 21188 11028 21244
rect 10964 21184 11028 21188
rect 5212 20980 5276 21044
rect 7788 20844 7852 20908
rect 796 20708 860 20772
rect 1348 20572 1412 20636
rect 5212 20708 5276 20772
rect 5580 20708 5644 20772
rect 7788 20708 7852 20772
rect 9628 20708 9692 20772
rect 3664 20700 3728 20704
rect 3664 20644 3668 20700
rect 3668 20644 3724 20700
rect 3724 20644 3728 20700
rect 3664 20640 3728 20644
rect 3744 20700 3808 20704
rect 3744 20644 3748 20700
rect 3748 20644 3804 20700
rect 3804 20644 3808 20700
rect 3744 20640 3808 20644
rect 3824 20700 3888 20704
rect 3824 20644 3828 20700
rect 3828 20644 3884 20700
rect 3884 20644 3888 20700
rect 3824 20640 3888 20644
rect 3904 20700 3968 20704
rect 3904 20644 3908 20700
rect 3908 20644 3964 20700
rect 3964 20644 3968 20700
rect 3904 20640 3968 20644
rect 10064 20700 10128 20704
rect 10064 20644 10068 20700
rect 10068 20644 10124 20700
rect 10124 20644 10128 20700
rect 10064 20640 10128 20644
rect 10144 20700 10208 20704
rect 10144 20644 10148 20700
rect 10148 20644 10204 20700
rect 10204 20644 10208 20700
rect 10144 20640 10208 20644
rect 10224 20700 10288 20704
rect 10224 20644 10228 20700
rect 10228 20644 10284 20700
rect 10284 20644 10288 20700
rect 10224 20640 10288 20644
rect 10304 20700 10368 20704
rect 10304 20644 10308 20700
rect 10308 20644 10364 20700
rect 10364 20644 10368 20700
rect 10304 20640 10368 20644
rect 4108 20632 4172 20636
rect 4108 20576 4122 20632
rect 4122 20576 4172 20632
rect 4108 20572 4172 20576
rect 5580 20572 5644 20636
rect 9076 20496 9140 20500
rect 9076 20440 9126 20496
rect 9126 20440 9140 20496
rect 9076 20436 9140 20440
rect 2452 20300 2516 20364
rect 1348 20164 1412 20228
rect 2636 20164 2700 20228
rect 4324 20156 4388 20160
rect 4324 20100 4328 20156
rect 4328 20100 4384 20156
rect 4384 20100 4388 20156
rect 4324 20096 4388 20100
rect 4404 20156 4468 20160
rect 4404 20100 4408 20156
rect 4408 20100 4464 20156
rect 4464 20100 4468 20156
rect 4404 20096 4468 20100
rect 4484 20156 4548 20160
rect 4484 20100 4488 20156
rect 4488 20100 4544 20156
rect 4544 20100 4548 20156
rect 4484 20096 4548 20100
rect 4564 20156 4628 20160
rect 4564 20100 4568 20156
rect 4568 20100 4624 20156
rect 4624 20100 4628 20156
rect 4564 20096 4628 20100
rect 10724 20156 10788 20160
rect 10724 20100 10728 20156
rect 10728 20100 10784 20156
rect 10784 20100 10788 20156
rect 10724 20096 10788 20100
rect 10804 20156 10868 20160
rect 10804 20100 10808 20156
rect 10808 20100 10864 20156
rect 10864 20100 10868 20156
rect 10804 20096 10868 20100
rect 10884 20156 10948 20160
rect 10884 20100 10888 20156
rect 10888 20100 10944 20156
rect 10944 20100 10948 20156
rect 10884 20096 10948 20100
rect 10964 20156 11028 20160
rect 10964 20100 10968 20156
rect 10968 20100 11024 20156
rect 11024 20100 11028 20156
rect 10964 20096 11028 20100
rect 1900 20028 1964 20092
rect 8156 20028 8220 20092
rect 9444 20028 9508 20092
rect 2452 19952 2516 19956
rect 2452 19896 2466 19952
rect 2466 19896 2516 19952
rect 2452 19892 2516 19896
rect 5212 19892 5276 19956
rect 4844 19680 4908 19684
rect 4844 19624 4894 19680
rect 4894 19624 4908 19680
rect 4844 19620 4908 19624
rect 5580 19620 5644 19684
rect 10548 19620 10612 19684
rect 3664 19612 3728 19616
rect 3664 19556 3668 19612
rect 3668 19556 3724 19612
rect 3724 19556 3728 19612
rect 3664 19552 3728 19556
rect 3744 19612 3808 19616
rect 3744 19556 3748 19612
rect 3748 19556 3804 19612
rect 3804 19556 3808 19612
rect 3744 19552 3808 19556
rect 3824 19612 3888 19616
rect 3824 19556 3828 19612
rect 3828 19556 3884 19612
rect 3884 19556 3888 19612
rect 3824 19552 3888 19556
rect 3904 19612 3968 19616
rect 3904 19556 3908 19612
rect 3908 19556 3964 19612
rect 3964 19556 3968 19612
rect 3904 19552 3968 19556
rect 10064 19612 10128 19616
rect 10064 19556 10068 19612
rect 10068 19556 10124 19612
rect 10124 19556 10128 19612
rect 10064 19552 10128 19556
rect 10144 19612 10208 19616
rect 10144 19556 10148 19612
rect 10148 19556 10204 19612
rect 10204 19556 10208 19612
rect 10144 19552 10208 19556
rect 10224 19612 10288 19616
rect 10224 19556 10228 19612
rect 10228 19556 10284 19612
rect 10284 19556 10288 19612
rect 10224 19552 10288 19556
rect 10304 19612 10368 19616
rect 10304 19556 10308 19612
rect 10308 19556 10364 19612
rect 10364 19556 10368 19612
rect 10304 19552 10368 19556
rect 4844 19484 4908 19548
rect 5580 19348 5644 19412
rect 7604 19348 7668 19412
rect 8708 19408 8772 19412
rect 8708 19352 8722 19408
rect 8722 19352 8772 19408
rect 8708 19348 8772 19352
rect 12020 19348 12084 19412
rect 2268 19272 2332 19276
rect 2268 19216 2318 19272
rect 2318 19216 2332 19272
rect 2268 19212 2332 19216
rect 5948 19212 6012 19276
rect 6500 19272 6564 19276
rect 6500 19216 6514 19272
rect 6514 19216 6564 19272
rect 6500 19212 6564 19216
rect 4324 19068 4388 19072
rect 4324 19012 4328 19068
rect 4328 19012 4384 19068
rect 4384 19012 4388 19068
rect 4324 19008 4388 19012
rect 4404 19068 4468 19072
rect 4404 19012 4408 19068
rect 4408 19012 4464 19068
rect 4464 19012 4468 19068
rect 4404 19008 4468 19012
rect 4484 19068 4548 19072
rect 4484 19012 4488 19068
rect 4488 19012 4544 19068
rect 4544 19012 4548 19068
rect 4484 19008 4548 19012
rect 4564 19068 4628 19072
rect 4564 19012 4568 19068
rect 4568 19012 4624 19068
rect 4624 19012 4628 19068
rect 4564 19008 4628 19012
rect 10724 19068 10788 19072
rect 10724 19012 10728 19068
rect 10728 19012 10784 19068
rect 10784 19012 10788 19068
rect 10724 19008 10788 19012
rect 10804 19068 10868 19072
rect 10804 19012 10808 19068
rect 10808 19012 10864 19068
rect 10864 19012 10868 19068
rect 10804 19008 10868 19012
rect 10884 19068 10948 19072
rect 10884 19012 10888 19068
rect 10888 19012 10944 19068
rect 10944 19012 10948 19068
rect 10884 19008 10948 19012
rect 10964 19068 11028 19072
rect 10964 19012 10968 19068
rect 10968 19012 11024 19068
rect 11024 19012 11028 19068
rect 10964 19008 11028 19012
rect 2820 18940 2884 19004
rect 4108 18940 4172 19004
rect 5396 19000 5460 19004
rect 5396 18944 5446 19000
rect 5446 18944 5460 19000
rect 5396 18940 5460 18944
rect 7972 19000 8036 19004
rect 7972 18944 7986 19000
rect 7986 18944 8036 19000
rect 7972 18940 8036 18944
rect 3372 18804 3436 18868
rect 3372 18668 3436 18732
rect 4108 18668 4172 18732
rect 3664 18524 3728 18528
rect 3664 18468 3668 18524
rect 3668 18468 3724 18524
rect 3724 18468 3728 18524
rect 3664 18464 3728 18468
rect 3744 18524 3808 18528
rect 3744 18468 3748 18524
rect 3748 18468 3804 18524
rect 3804 18468 3808 18524
rect 3744 18464 3808 18468
rect 3824 18524 3888 18528
rect 3824 18468 3828 18524
rect 3828 18468 3884 18524
rect 3884 18468 3888 18524
rect 3824 18464 3888 18468
rect 3904 18524 3968 18528
rect 3904 18468 3908 18524
rect 3908 18468 3964 18524
rect 3964 18468 3968 18524
rect 3904 18464 3968 18468
rect 10064 18524 10128 18528
rect 10064 18468 10068 18524
rect 10068 18468 10124 18524
rect 10124 18468 10128 18524
rect 10064 18464 10128 18468
rect 10144 18524 10208 18528
rect 10144 18468 10148 18524
rect 10148 18468 10204 18524
rect 10204 18468 10208 18524
rect 10144 18464 10208 18468
rect 10224 18524 10288 18528
rect 10224 18468 10228 18524
rect 10228 18468 10284 18524
rect 10284 18468 10288 18524
rect 10224 18464 10288 18468
rect 10304 18524 10368 18528
rect 10304 18468 10308 18524
rect 10308 18468 10364 18524
rect 10364 18468 10368 18524
rect 10304 18464 10368 18468
rect 5396 17988 5460 18052
rect 6684 18124 6748 18188
rect 4324 17980 4388 17984
rect 4324 17924 4328 17980
rect 4328 17924 4384 17980
rect 4384 17924 4388 17980
rect 4324 17920 4388 17924
rect 4404 17980 4468 17984
rect 4404 17924 4408 17980
rect 4408 17924 4464 17980
rect 4464 17924 4468 17980
rect 4404 17920 4468 17924
rect 4484 17980 4548 17984
rect 4484 17924 4488 17980
rect 4488 17924 4544 17980
rect 4544 17924 4548 17980
rect 4484 17920 4548 17924
rect 4564 17980 4628 17984
rect 4564 17924 4568 17980
rect 4568 17924 4624 17980
rect 4624 17924 4628 17980
rect 4564 17920 4628 17924
rect 10724 17980 10788 17984
rect 10724 17924 10728 17980
rect 10728 17924 10784 17980
rect 10784 17924 10788 17980
rect 10724 17920 10788 17924
rect 10804 17980 10868 17984
rect 10804 17924 10808 17980
rect 10808 17924 10864 17980
rect 10864 17924 10868 17980
rect 10804 17920 10868 17924
rect 10884 17980 10948 17984
rect 10884 17924 10888 17980
rect 10888 17924 10944 17980
rect 10944 17924 10948 17980
rect 10884 17920 10948 17924
rect 10964 17980 11028 17984
rect 10964 17924 10968 17980
rect 10968 17924 11024 17980
rect 11024 17924 11028 17980
rect 10964 17920 11028 17924
rect 6132 17912 6196 17916
rect 6132 17856 6146 17912
rect 6146 17856 6196 17912
rect 6132 17852 6196 17856
rect 7788 17852 7852 17916
rect 8892 17852 8956 17916
rect 9444 17912 9508 17916
rect 9444 17856 9458 17912
rect 9458 17856 9508 17912
rect 9444 17852 9508 17856
rect 428 17716 492 17780
rect 3188 17716 3252 17780
rect 7052 17716 7116 17780
rect 8708 17716 8772 17780
rect 9076 17776 9140 17780
rect 9076 17720 9126 17776
rect 9126 17720 9140 17776
rect 9076 17716 9140 17720
rect 11468 17776 11532 17780
rect 11468 17720 11482 17776
rect 11482 17720 11532 17776
rect 11468 17716 11532 17720
rect 7420 17580 7484 17644
rect 11284 17580 11348 17644
rect 8524 17444 8588 17508
rect 3664 17436 3728 17440
rect 3664 17380 3668 17436
rect 3668 17380 3724 17436
rect 3724 17380 3728 17436
rect 3664 17376 3728 17380
rect 3744 17436 3808 17440
rect 3744 17380 3748 17436
rect 3748 17380 3804 17436
rect 3804 17380 3808 17436
rect 3744 17376 3808 17380
rect 3824 17436 3888 17440
rect 3824 17380 3828 17436
rect 3828 17380 3884 17436
rect 3884 17380 3888 17436
rect 3824 17376 3888 17380
rect 3904 17436 3968 17440
rect 3904 17380 3908 17436
rect 3908 17380 3964 17436
rect 3964 17380 3968 17436
rect 3904 17376 3968 17380
rect 10064 17436 10128 17440
rect 10064 17380 10068 17436
rect 10068 17380 10124 17436
rect 10124 17380 10128 17436
rect 10064 17376 10128 17380
rect 10144 17436 10208 17440
rect 10144 17380 10148 17436
rect 10148 17380 10204 17436
rect 10204 17380 10208 17436
rect 10144 17376 10208 17380
rect 10224 17436 10288 17440
rect 10224 17380 10228 17436
rect 10228 17380 10284 17436
rect 10284 17380 10288 17436
rect 10224 17376 10288 17380
rect 10304 17436 10368 17440
rect 10304 17380 10308 17436
rect 10308 17380 10364 17436
rect 10364 17380 10368 17436
rect 10304 17376 10368 17380
rect 5764 17308 5828 17372
rect 6684 17232 6748 17236
rect 6684 17176 6698 17232
rect 6698 17176 6748 17232
rect 6684 17172 6748 17176
rect 9628 17172 9692 17236
rect 2268 17036 2332 17100
rect 2820 17036 2884 17100
rect 4324 16892 4388 16896
rect 4324 16836 4328 16892
rect 4328 16836 4384 16892
rect 4384 16836 4388 16892
rect 4324 16832 4388 16836
rect 4404 16892 4468 16896
rect 4404 16836 4408 16892
rect 4408 16836 4464 16892
rect 4464 16836 4468 16892
rect 4404 16832 4468 16836
rect 4484 16892 4548 16896
rect 4484 16836 4488 16892
rect 4488 16836 4544 16892
rect 4544 16836 4548 16892
rect 4484 16832 4548 16836
rect 4564 16892 4628 16896
rect 4564 16836 4568 16892
rect 4568 16836 4624 16892
rect 4624 16836 4628 16892
rect 4564 16832 4628 16836
rect 2636 16764 2700 16828
rect 6684 16900 6748 16964
rect 10724 16892 10788 16896
rect 10724 16836 10728 16892
rect 10728 16836 10784 16892
rect 10784 16836 10788 16892
rect 10724 16832 10788 16836
rect 10804 16892 10868 16896
rect 10804 16836 10808 16892
rect 10808 16836 10864 16892
rect 10864 16836 10868 16892
rect 10804 16832 10868 16836
rect 10884 16892 10948 16896
rect 10884 16836 10888 16892
rect 10888 16836 10944 16892
rect 10944 16836 10948 16892
rect 10884 16832 10948 16836
rect 10964 16892 11028 16896
rect 10964 16836 10968 16892
rect 10968 16836 11024 16892
rect 11024 16836 11028 16892
rect 10964 16832 11028 16836
rect 3188 16628 3252 16692
rect 9076 16628 9140 16692
rect 1164 16492 1228 16556
rect 7788 16492 7852 16556
rect 9812 16492 9876 16556
rect 1348 16356 1412 16420
rect 4844 16356 4908 16420
rect 3664 16348 3728 16352
rect 3664 16292 3668 16348
rect 3668 16292 3724 16348
rect 3724 16292 3728 16348
rect 3664 16288 3728 16292
rect 3744 16348 3808 16352
rect 3744 16292 3748 16348
rect 3748 16292 3804 16348
rect 3804 16292 3808 16348
rect 3744 16288 3808 16292
rect 3824 16348 3888 16352
rect 3824 16292 3828 16348
rect 3828 16292 3884 16348
rect 3884 16292 3888 16348
rect 3824 16288 3888 16292
rect 3904 16348 3968 16352
rect 3904 16292 3908 16348
rect 3908 16292 3964 16348
rect 3964 16292 3968 16348
rect 3904 16288 3968 16292
rect 10064 16348 10128 16352
rect 10064 16292 10068 16348
rect 10068 16292 10124 16348
rect 10124 16292 10128 16348
rect 10064 16288 10128 16292
rect 10144 16348 10208 16352
rect 10144 16292 10148 16348
rect 10148 16292 10204 16348
rect 10204 16292 10208 16348
rect 10144 16288 10208 16292
rect 10224 16348 10288 16352
rect 10224 16292 10228 16348
rect 10228 16292 10284 16348
rect 10284 16292 10288 16348
rect 10224 16288 10288 16292
rect 10304 16348 10368 16352
rect 10304 16292 10308 16348
rect 10308 16292 10364 16348
rect 10364 16292 10368 16348
rect 10304 16288 10368 16292
rect 4108 16220 4172 16284
rect 9812 16220 9876 16284
rect 980 16084 1044 16148
rect 9260 16084 9324 16148
rect 612 15812 676 15876
rect 4324 15804 4388 15808
rect 4324 15748 4328 15804
rect 4328 15748 4384 15804
rect 4384 15748 4388 15804
rect 4324 15744 4388 15748
rect 4404 15804 4468 15808
rect 4404 15748 4408 15804
rect 4408 15748 4464 15804
rect 4464 15748 4468 15804
rect 4404 15744 4468 15748
rect 4484 15804 4548 15808
rect 4484 15748 4488 15804
rect 4488 15748 4544 15804
rect 4544 15748 4548 15804
rect 4484 15744 4548 15748
rect 4564 15804 4628 15808
rect 4564 15748 4568 15804
rect 4568 15748 4624 15804
rect 4624 15748 4628 15804
rect 4564 15744 4628 15748
rect 10724 15804 10788 15808
rect 10724 15748 10728 15804
rect 10728 15748 10784 15804
rect 10784 15748 10788 15804
rect 10724 15744 10788 15748
rect 10804 15804 10868 15808
rect 10804 15748 10808 15804
rect 10808 15748 10864 15804
rect 10864 15748 10868 15804
rect 10804 15744 10868 15748
rect 10884 15804 10948 15808
rect 10884 15748 10888 15804
rect 10888 15748 10944 15804
rect 10944 15748 10948 15804
rect 10884 15744 10948 15748
rect 10964 15804 11028 15808
rect 10964 15748 10968 15804
rect 10968 15748 11024 15804
rect 11024 15748 11028 15804
rect 10964 15744 11028 15748
rect 1716 15736 1780 15740
rect 1716 15680 1730 15736
rect 1730 15680 1780 15736
rect 1716 15676 1780 15680
rect 11836 15600 11900 15604
rect 11836 15544 11850 15600
rect 11850 15544 11900 15600
rect 11836 15540 11900 15544
rect 60 15404 124 15468
rect 2636 15404 2700 15468
rect 3188 15268 3252 15332
rect 9260 15268 9324 15332
rect 3664 15260 3728 15264
rect 3664 15204 3668 15260
rect 3668 15204 3724 15260
rect 3724 15204 3728 15260
rect 3664 15200 3728 15204
rect 3744 15260 3808 15264
rect 3744 15204 3748 15260
rect 3748 15204 3804 15260
rect 3804 15204 3808 15260
rect 3744 15200 3808 15204
rect 3824 15260 3888 15264
rect 3824 15204 3828 15260
rect 3828 15204 3884 15260
rect 3884 15204 3888 15260
rect 3824 15200 3888 15204
rect 3904 15260 3968 15264
rect 3904 15204 3908 15260
rect 3908 15204 3964 15260
rect 3964 15204 3968 15260
rect 3904 15200 3968 15204
rect 10064 15260 10128 15264
rect 10064 15204 10068 15260
rect 10068 15204 10124 15260
rect 10124 15204 10128 15260
rect 10064 15200 10128 15204
rect 10144 15260 10208 15264
rect 10144 15204 10148 15260
rect 10148 15204 10204 15260
rect 10204 15204 10208 15260
rect 10144 15200 10208 15204
rect 10224 15260 10288 15264
rect 10224 15204 10228 15260
rect 10228 15204 10284 15260
rect 10284 15204 10288 15260
rect 10224 15200 10288 15204
rect 10304 15260 10368 15264
rect 10304 15204 10308 15260
rect 10308 15204 10364 15260
rect 10364 15204 10368 15260
rect 10304 15200 10368 15204
rect 3372 14860 3436 14924
rect 12572 14860 12636 14924
rect 4324 14716 4388 14720
rect 4324 14660 4328 14716
rect 4328 14660 4384 14716
rect 4384 14660 4388 14716
rect 4324 14656 4388 14660
rect 4404 14716 4468 14720
rect 4404 14660 4408 14716
rect 4408 14660 4464 14716
rect 4464 14660 4468 14716
rect 4404 14656 4468 14660
rect 4484 14716 4548 14720
rect 4484 14660 4488 14716
rect 4488 14660 4544 14716
rect 4544 14660 4548 14716
rect 4484 14656 4548 14660
rect 4564 14716 4628 14720
rect 4564 14660 4568 14716
rect 4568 14660 4624 14716
rect 4624 14660 4628 14716
rect 4564 14656 4628 14660
rect 10724 14716 10788 14720
rect 10724 14660 10728 14716
rect 10728 14660 10784 14716
rect 10784 14660 10788 14716
rect 10724 14656 10788 14660
rect 10804 14716 10868 14720
rect 10804 14660 10808 14716
rect 10808 14660 10864 14716
rect 10864 14660 10868 14716
rect 10804 14656 10868 14660
rect 10884 14716 10948 14720
rect 10884 14660 10888 14716
rect 10888 14660 10944 14716
rect 10944 14660 10948 14716
rect 10884 14656 10948 14660
rect 10964 14716 11028 14720
rect 10964 14660 10968 14716
rect 10968 14660 11024 14716
rect 11024 14660 11028 14716
rect 10964 14656 11028 14660
rect 5028 14452 5092 14516
rect 6316 14452 6380 14516
rect 3664 14172 3728 14176
rect 3664 14116 3668 14172
rect 3668 14116 3724 14172
rect 3724 14116 3728 14172
rect 3664 14112 3728 14116
rect 3744 14172 3808 14176
rect 3744 14116 3748 14172
rect 3748 14116 3804 14172
rect 3804 14116 3808 14172
rect 3744 14112 3808 14116
rect 3824 14172 3888 14176
rect 3824 14116 3828 14172
rect 3828 14116 3884 14172
rect 3884 14116 3888 14172
rect 3824 14112 3888 14116
rect 3904 14172 3968 14176
rect 3904 14116 3908 14172
rect 3908 14116 3964 14172
rect 3964 14116 3968 14172
rect 3904 14112 3968 14116
rect 10064 14172 10128 14176
rect 10064 14116 10068 14172
rect 10068 14116 10124 14172
rect 10124 14116 10128 14172
rect 10064 14112 10128 14116
rect 10144 14172 10208 14176
rect 10144 14116 10148 14172
rect 10148 14116 10204 14172
rect 10204 14116 10208 14172
rect 10144 14112 10208 14116
rect 10224 14172 10288 14176
rect 10224 14116 10228 14172
rect 10228 14116 10284 14172
rect 10284 14116 10288 14172
rect 10224 14112 10288 14116
rect 10304 14172 10368 14176
rect 10304 14116 10308 14172
rect 10308 14116 10364 14172
rect 10364 14116 10368 14172
rect 10304 14112 10368 14116
rect 5764 13772 5828 13836
rect 7788 13636 7852 13700
rect 11652 13696 11716 13700
rect 11652 13640 11702 13696
rect 11702 13640 11716 13696
rect 11652 13636 11716 13640
rect 4324 13628 4388 13632
rect 4324 13572 4328 13628
rect 4328 13572 4384 13628
rect 4384 13572 4388 13628
rect 4324 13568 4388 13572
rect 4404 13628 4468 13632
rect 4404 13572 4408 13628
rect 4408 13572 4464 13628
rect 4464 13572 4468 13628
rect 4404 13568 4468 13572
rect 4484 13628 4548 13632
rect 4484 13572 4488 13628
rect 4488 13572 4544 13628
rect 4544 13572 4548 13628
rect 4484 13568 4548 13572
rect 4564 13628 4628 13632
rect 4564 13572 4568 13628
rect 4568 13572 4624 13628
rect 4624 13572 4628 13628
rect 4564 13568 4628 13572
rect 10724 13628 10788 13632
rect 10724 13572 10728 13628
rect 10728 13572 10784 13628
rect 10784 13572 10788 13628
rect 10724 13568 10788 13572
rect 10804 13628 10868 13632
rect 10804 13572 10808 13628
rect 10808 13572 10864 13628
rect 10864 13572 10868 13628
rect 10804 13568 10868 13572
rect 10884 13628 10948 13632
rect 10884 13572 10888 13628
rect 10888 13572 10944 13628
rect 10944 13572 10948 13628
rect 10884 13568 10948 13572
rect 10964 13628 11028 13632
rect 10964 13572 10968 13628
rect 10968 13572 11024 13628
rect 11024 13572 11028 13628
rect 10964 13568 11028 13572
rect 3664 13084 3728 13088
rect 3664 13028 3668 13084
rect 3668 13028 3724 13084
rect 3724 13028 3728 13084
rect 3664 13024 3728 13028
rect 3744 13084 3808 13088
rect 3744 13028 3748 13084
rect 3748 13028 3804 13084
rect 3804 13028 3808 13084
rect 3744 13024 3808 13028
rect 3824 13084 3888 13088
rect 3824 13028 3828 13084
rect 3828 13028 3884 13084
rect 3884 13028 3888 13084
rect 3824 13024 3888 13028
rect 3904 13084 3968 13088
rect 3904 13028 3908 13084
rect 3908 13028 3964 13084
rect 3964 13028 3968 13084
rect 3904 13024 3968 13028
rect 10064 13084 10128 13088
rect 10064 13028 10068 13084
rect 10068 13028 10124 13084
rect 10124 13028 10128 13084
rect 10064 13024 10128 13028
rect 10144 13084 10208 13088
rect 10144 13028 10148 13084
rect 10148 13028 10204 13084
rect 10204 13028 10208 13084
rect 10144 13024 10208 13028
rect 10224 13084 10288 13088
rect 10224 13028 10228 13084
rect 10228 13028 10284 13084
rect 10284 13028 10288 13084
rect 10224 13024 10288 13028
rect 10304 13084 10368 13088
rect 10304 13028 10308 13084
rect 10308 13028 10364 13084
rect 10364 13028 10368 13084
rect 10304 13024 10368 13028
rect 5948 12820 6012 12884
rect 8892 12880 8956 12884
rect 8892 12824 8942 12880
rect 8942 12824 8956 12880
rect 8892 12820 8956 12824
rect 4324 12540 4388 12544
rect 4324 12484 4328 12540
rect 4328 12484 4384 12540
rect 4384 12484 4388 12540
rect 4324 12480 4388 12484
rect 4404 12540 4468 12544
rect 4404 12484 4408 12540
rect 4408 12484 4464 12540
rect 4464 12484 4468 12540
rect 4404 12480 4468 12484
rect 4484 12540 4548 12544
rect 4484 12484 4488 12540
rect 4488 12484 4544 12540
rect 4544 12484 4548 12540
rect 4484 12480 4548 12484
rect 4564 12540 4628 12544
rect 4564 12484 4568 12540
rect 4568 12484 4624 12540
rect 4624 12484 4628 12540
rect 4564 12480 4628 12484
rect 10724 12540 10788 12544
rect 10724 12484 10728 12540
rect 10728 12484 10784 12540
rect 10784 12484 10788 12540
rect 10724 12480 10788 12484
rect 10804 12540 10868 12544
rect 10804 12484 10808 12540
rect 10808 12484 10864 12540
rect 10864 12484 10868 12540
rect 10804 12480 10868 12484
rect 10884 12540 10948 12544
rect 10884 12484 10888 12540
rect 10888 12484 10944 12540
rect 10944 12484 10948 12540
rect 10884 12480 10948 12484
rect 10964 12540 11028 12544
rect 10964 12484 10968 12540
rect 10968 12484 11024 12540
rect 11024 12484 11028 12540
rect 10964 12480 11028 12484
rect 5212 12472 5276 12476
rect 5212 12416 5262 12472
rect 5262 12416 5276 12472
rect 5212 12412 5276 12416
rect 11100 12472 11164 12476
rect 11100 12416 11150 12472
rect 11150 12416 11164 12472
rect 11100 12412 11164 12416
rect 5212 12336 5276 12340
rect 5212 12280 5262 12336
rect 5262 12280 5276 12336
rect 5212 12276 5276 12280
rect 10548 12276 10612 12340
rect 3664 11996 3728 12000
rect 3664 11940 3668 11996
rect 3668 11940 3724 11996
rect 3724 11940 3728 11996
rect 3664 11936 3728 11940
rect 3744 11996 3808 12000
rect 3744 11940 3748 11996
rect 3748 11940 3804 11996
rect 3804 11940 3808 11996
rect 3744 11936 3808 11940
rect 3824 11996 3888 12000
rect 3824 11940 3828 11996
rect 3828 11940 3884 11996
rect 3884 11940 3888 11996
rect 3824 11936 3888 11940
rect 3904 11996 3968 12000
rect 3904 11940 3908 11996
rect 3908 11940 3964 11996
rect 3964 11940 3968 11996
rect 3904 11936 3968 11940
rect 10064 11996 10128 12000
rect 10064 11940 10068 11996
rect 10068 11940 10124 11996
rect 10124 11940 10128 11996
rect 10064 11936 10128 11940
rect 10144 11996 10208 12000
rect 10144 11940 10148 11996
rect 10148 11940 10204 11996
rect 10204 11940 10208 11996
rect 10144 11936 10208 11940
rect 10224 11996 10288 12000
rect 10224 11940 10228 11996
rect 10228 11940 10284 11996
rect 10284 11940 10288 11996
rect 10224 11936 10288 11940
rect 10304 11996 10368 12000
rect 10304 11940 10308 11996
rect 10308 11940 10364 11996
rect 10364 11940 10368 11996
rect 10304 11936 10368 11940
rect 4324 11452 4388 11456
rect 4324 11396 4328 11452
rect 4328 11396 4384 11452
rect 4384 11396 4388 11452
rect 4324 11392 4388 11396
rect 4404 11452 4468 11456
rect 4404 11396 4408 11452
rect 4408 11396 4464 11452
rect 4464 11396 4468 11452
rect 4404 11392 4468 11396
rect 4484 11452 4548 11456
rect 4484 11396 4488 11452
rect 4488 11396 4544 11452
rect 4544 11396 4548 11452
rect 4484 11392 4548 11396
rect 4564 11452 4628 11456
rect 4564 11396 4568 11452
rect 4568 11396 4624 11452
rect 4624 11396 4628 11452
rect 4564 11392 4628 11396
rect 10724 11452 10788 11456
rect 10724 11396 10728 11452
rect 10728 11396 10784 11452
rect 10784 11396 10788 11452
rect 10724 11392 10788 11396
rect 10804 11452 10868 11456
rect 10804 11396 10808 11452
rect 10808 11396 10864 11452
rect 10864 11396 10868 11452
rect 10804 11392 10868 11396
rect 10884 11452 10948 11456
rect 10884 11396 10888 11452
rect 10888 11396 10944 11452
rect 10944 11396 10948 11452
rect 10884 11392 10948 11396
rect 10964 11452 11028 11456
rect 10964 11396 10968 11452
rect 10968 11396 11024 11452
rect 11024 11396 11028 11452
rect 10964 11392 11028 11396
rect 2084 11188 2148 11252
rect 8156 11112 8220 11116
rect 8156 11056 8170 11112
rect 8170 11056 8220 11112
rect 8156 11052 8220 11056
rect 3664 10908 3728 10912
rect 3664 10852 3668 10908
rect 3668 10852 3724 10908
rect 3724 10852 3728 10908
rect 3664 10848 3728 10852
rect 3744 10908 3808 10912
rect 3744 10852 3748 10908
rect 3748 10852 3804 10908
rect 3804 10852 3808 10908
rect 3744 10848 3808 10852
rect 3824 10908 3888 10912
rect 3824 10852 3828 10908
rect 3828 10852 3884 10908
rect 3884 10852 3888 10908
rect 3824 10848 3888 10852
rect 3904 10908 3968 10912
rect 3904 10852 3908 10908
rect 3908 10852 3964 10908
rect 3964 10852 3968 10908
rect 3904 10848 3968 10852
rect 10064 10908 10128 10912
rect 10064 10852 10068 10908
rect 10068 10852 10124 10908
rect 10124 10852 10128 10908
rect 10064 10848 10128 10852
rect 10144 10908 10208 10912
rect 10144 10852 10148 10908
rect 10148 10852 10204 10908
rect 10204 10852 10208 10908
rect 10144 10848 10208 10852
rect 10224 10908 10288 10912
rect 10224 10852 10228 10908
rect 10228 10852 10284 10908
rect 10284 10852 10288 10908
rect 10224 10848 10288 10852
rect 10304 10908 10368 10912
rect 10304 10852 10308 10908
rect 10308 10852 10364 10908
rect 10364 10852 10368 10908
rect 10304 10848 10368 10852
rect 4324 10364 4388 10368
rect 4324 10308 4328 10364
rect 4328 10308 4384 10364
rect 4384 10308 4388 10364
rect 4324 10304 4388 10308
rect 4404 10364 4468 10368
rect 4404 10308 4408 10364
rect 4408 10308 4464 10364
rect 4464 10308 4468 10364
rect 4404 10304 4468 10308
rect 4484 10364 4548 10368
rect 4484 10308 4488 10364
rect 4488 10308 4544 10364
rect 4544 10308 4548 10364
rect 4484 10304 4548 10308
rect 4564 10364 4628 10368
rect 4564 10308 4568 10364
rect 4568 10308 4624 10364
rect 4624 10308 4628 10364
rect 4564 10304 4628 10308
rect 10724 10364 10788 10368
rect 10724 10308 10728 10364
rect 10728 10308 10784 10364
rect 10784 10308 10788 10364
rect 10724 10304 10788 10308
rect 10804 10364 10868 10368
rect 10804 10308 10808 10364
rect 10808 10308 10864 10364
rect 10864 10308 10868 10364
rect 10804 10304 10868 10308
rect 10884 10364 10948 10368
rect 10884 10308 10888 10364
rect 10888 10308 10944 10364
rect 10944 10308 10948 10364
rect 10884 10304 10948 10308
rect 10964 10364 11028 10368
rect 10964 10308 10968 10364
rect 10968 10308 11024 10364
rect 11024 10308 11028 10364
rect 10964 10304 11028 10308
rect 5396 9964 5460 10028
rect 9812 10024 9876 10028
rect 9812 9968 9862 10024
rect 9862 9968 9876 10024
rect 9812 9964 9876 9968
rect 11100 9964 11164 10028
rect 3664 9820 3728 9824
rect 3664 9764 3668 9820
rect 3668 9764 3724 9820
rect 3724 9764 3728 9820
rect 3664 9760 3728 9764
rect 3744 9820 3808 9824
rect 3744 9764 3748 9820
rect 3748 9764 3804 9820
rect 3804 9764 3808 9820
rect 3744 9760 3808 9764
rect 3824 9820 3888 9824
rect 3824 9764 3828 9820
rect 3828 9764 3884 9820
rect 3884 9764 3888 9820
rect 3824 9760 3888 9764
rect 3904 9820 3968 9824
rect 3904 9764 3908 9820
rect 3908 9764 3964 9820
rect 3964 9764 3968 9820
rect 3904 9760 3968 9764
rect 10064 9820 10128 9824
rect 10064 9764 10068 9820
rect 10068 9764 10124 9820
rect 10124 9764 10128 9820
rect 10064 9760 10128 9764
rect 10144 9820 10208 9824
rect 10144 9764 10148 9820
rect 10148 9764 10204 9820
rect 10204 9764 10208 9820
rect 10144 9760 10208 9764
rect 10224 9820 10288 9824
rect 10224 9764 10228 9820
rect 10228 9764 10284 9820
rect 10284 9764 10288 9820
rect 10224 9760 10288 9764
rect 10304 9820 10368 9824
rect 10304 9764 10308 9820
rect 10308 9764 10364 9820
rect 10364 9764 10368 9820
rect 10304 9760 10368 9764
rect 10548 9420 10612 9484
rect 4324 9276 4388 9280
rect 4324 9220 4328 9276
rect 4328 9220 4384 9276
rect 4384 9220 4388 9276
rect 4324 9216 4388 9220
rect 4404 9276 4468 9280
rect 4404 9220 4408 9276
rect 4408 9220 4464 9276
rect 4464 9220 4468 9276
rect 4404 9216 4468 9220
rect 4484 9276 4548 9280
rect 4484 9220 4488 9276
rect 4488 9220 4544 9276
rect 4544 9220 4548 9276
rect 4484 9216 4548 9220
rect 4564 9276 4628 9280
rect 4564 9220 4568 9276
rect 4568 9220 4624 9276
rect 4624 9220 4628 9276
rect 4564 9216 4628 9220
rect 10724 9276 10788 9280
rect 10724 9220 10728 9276
rect 10728 9220 10784 9276
rect 10784 9220 10788 9276
rect 10724 9216 10788 9220
rect 10804 9276 10868 9280
rect 10804 9220 10808 9276
rect 10808 9220 10864 9276
rect 10864 9220 10868 9276
rect 10804 9216 10868 9220
rect 10884 9276 10948 9280
rect 10884 9220 10888 9276
rect 10888 9220 10944 9276
rect 10944 9220 10948 9276
rect 10884 9216 10948 9220
rect 10964 9276 11028 9280
rect 10964 9220 10968 9276
rect 10968 9220 11024 9276
rect 11024 9220 11028 9276
rect 10964 9216 11028 9220
rect 3664 8732 3728 8736
rect 3664 8676 3668 8732
rect 3668 8676 3724 8732
rect 3724 8676 3728 8732
rect 3664 8672 3728 8676
rect 3744 8732 3808 8736
rect 3744 8676 3748 8732
rect 3748 8676 3804 8732
rect 3804 8676 3808 8732
rect 3744 8672 3808 8676
rect 3824 8732 3888 8736
rect 3824 8676 3828 8732
rect 3828 8676 3884 8732
rect 3884 8676 3888 8732
rect 3824 8672 3888 8676
rect 3904 8732 3968 8736
rect 3904 8676 3908 8732
rect 3908 8676 3964 8732
rect 3964 8676 3968 8732
rect 3904 8672 3968 8676
rect 10064 8732 10128 8736
rect 10064 8676 10068 8732
rect 10068 8676 10124 8732
rect 10124 8676 10128 8732
rect 10064 8672 10128 8676
rect 10144 8732 10208 8736
rect 10144 8676 10148 8732
rect 10148 8676 10204 8732
rect 10204 8676 10208 8732
rect 10144 8672 10208 8676
rect 10224 8732 10288 8736
rect 10224 8676 10228 8732
rect 10228 8676 10284 8732
rect 10284 8676 10288 8732
rect 10224 8672 10288 8676
rect 10304 8732 10368 8736
rect 10304 8676 10308 8732
rect 10308 8676 10364 8732
rect 10364 8676 10368 8732
rect 10304 8672 10368 8676
rect 5580 8664 5644 8668
rect 5580 8608 5594 8664
rect 5594 8608 5644 8664
rect 5580 8604 5644 8608
rect 7420 8196 7484 8260
rect 4324 8188 4388 8192
rect 4324 8132 4328 8188
rect 4328 8132 4384 8188
rect 4384 8132 4388 8188
rect 4324 8128 4388 8132
rect 4404 8188 4468 8192
rect 4404 8132 4408 8188
rect 4408 8132 4464 8188
rect 4464 8132 4468 8188
rect 4404 8128 4468 8132
rect 4484 8188 4548 8192
rect 4484 8132 4488 8188
rect 4488 8132 4544 8188
rect 4544 8132 4548 8188
rect 4484 8128 4548 8132
rect 4564 8188 4628 8192
rect 4564 8132 4568 8188
rect 4568 8132 4624 8188
rect 4624 8132 4628 8188
rect 4564 8128 4628 8132
rect 10724 8188 10788 8192
rect 10724 8132 10728 8188
rect 10728 8132 10784 8188
rect 10784 8132 10788 8188
rect 10724 8128 10788 8132
rect 10804 8188 10868 8192
rect 10804 8132 10808 8188
rect 10808 8132 10864 8188
rect 10864 8132 10868 8188
rect 10804 8128 10868 8132
rect 10884 8188 10948 8192
rect 10884 8132 10888 8188
rect 10888 8132 10944 8188
rect 10944 8132 10948 8188
rect 10884 8128 10948 8132
rect 10964 8188 11028 8192
rect 10964 8132 10968 8188
rect 10968 8132 11024 8188
rect 11024 8132 11028 8188
rect 10964 8128 11028 8132
rect 9444 8120 9508 8124
rect 9444 8064 9494 8120
rect 9494 8064 9508 8120
rect 9444 8060 9508 8064
rect 3664 7644 3728 7648
rect 3664 7588 3668 7644
rect 3668 7588 3724 7644
rect 3724 7588 3728 7644
rect 3664 7584 3728 7588
rect 3744 7644 3808 7648
rect 3744 7588 3748 7644
rect 3748 7588 3804 7644
rect 3804 7588 3808 7644
rect 3744 7584 3808 7588
rect 3824 7644 3888 7648
rect 3824 7588 3828 7644
rect 3828 7588 3884 7644
rect 3884 7588 3888 7644
rect 3824 7584 3888 7588
rect 3904 7644 3968 7648
rect 3904 7588 3908 7644
rect 3908 7588 3964 7644
rect 3964 7588 3968 7644
rect 3904 7584 3968 7588
rect 10064 7644 10128 7648
rect 10064 7588 10068 7644
rect 10068 7588 10124 7644
rect 10124 7588 10128 7644
rect 10064 7584 10128 7588
rect 10144 7644 10208 7648
rect 10144 7588 10148 7644
rect 10148 7588 10204 7644
rect 10204 7588 10208 7644
rect 10144 7584 10208 7588
rect 10224 7644 10288 7648
rect 10224 7588 10228 7644
rect 10228 7588 10284 7644
rect 10284 7588 10288 7644
rect 10224 7584 10288 7588
rect 10304 7644 10368 7648
rect 10304 7588 10308 7644
rect 10308 7588 10364 7644
rect 10364 7588 10368 7644
rect 10304 7584 10368 7588
rect 9076 7380 9140 7444
rect 9812 7304 9876 7308
rect 9812 7248 9826 7304
rect 9826 7248 9876 7304
rect 9812 7244 9876 7248
rect 60 7108 124 7172
rect 4324 7100 4388 7104
rect 4324 7044 4328 7100
rect 4328 7044 4384 7100
rect 4384 7044 4388 7100
rect 4324 7040 4388 7044
rect 4404 7100 4468 7104
rect 4404 7044 4408 7100
rect 4408 7044 4464 7100
rect 4464 7044 4468 7100
rect 4404 7040 4468 7044
rect 4484 7100 4548 7104
rect 4484 7044 4488 7100
rect 4488 7044 4544 7100
rect 4544 7044 4548 7100
rect 4484 7040 4548 7044
rect 4564 7100 4628 7104
rect 4564 7044 4568 7100
rect 4568 7044 4624 7100
rect 4624 7044 4628 7100
rect 4564 7040 4628 7044
rect 10724 7100 10788 7104
rect 10724 7044 10728 7100
rect 10728 7044 10784 7100
rect 10784 7044 10788 7100
rect 10724 7040 10788 7044
rect 10804 7100 10868 7104
rect 10804 7044 10808 7100
rect 10808 7044 10864 7100
rect 10864 7044 10868 7100
rect 10804 7040 10868 7044
rect 10884 7100 10948 7104
rect 10884 7044 10888 7100
rect 10888 7044 10944 7100
rect 10944 7044 10948 7100
rect 10884 7040 10948 7044
rect 10964 7100 11028 7104
rect 10964 7044 10968 7100
rect 10968 7044 11024 7100
rect 11024 7044 11028 7100
rect 10964 7040 11028 7044
rect 10548 6836 10612 6900
rect 3664 6556 3728 6560
rect 3664 6500 3668 6556
rect 3668 6500 3724 6556
rect 3724 6500 3728 6556
rect 3664 6496 3728 6500
rect 3744 6556 3808 6560
rect 3744 6500 3748 6556
rect 3748 6500 3804 6556
rect 3804 6500 3808 6556
rect 3744 6496 3808 6500
rect 3824 6556 3888 6560
rect 3824 6500 3828 6556
rect 3828 6500 3884 6556
rect 3884 6500 3888 6556
rect 3824 6496 3888 6500
rect 3904 6556 3968 6560
rect 3904 6500 3908 6556
rect 3908 6500 3964 6556
rect 3964 6500 3968 6556
rect 3904 6496 3968 6500
rect 10064 6556 10128 6560
rect 10064 6500 10068 6556
rect 10068 6500 10124 6556
rect 10124 6500 10128 6556
rect 10064 6496 10128 6500
rect 10144 6556 10208 6560
rect 10144 6500 10148 6556
rect 10148 6500 10204 6556
rect 10204 6500 10208 6556
rect 10144 6496 10208 6500
rect 10224 6556 10288 6560
rect 10224 6500 10228 6556
rect 10228 6500 10284 6556
rect 10284 6500 10288 6556
rect 10224 6496 10288 6500
rect 10304 6556 10368 6560
rect 10304 6500 10308 6556
rect 10308 6500 10364 6556
rect 10364 6500 10368 6556
rect 10304 6496 10368 6500
rect 4324 6012 4388 6016
rect 4324 5956 4328 6012
rect 4328 5956 4384 6012
rect 4384 5956 4388 6012
rect 4324 5952 4388 5956
rect 4404 6012 4468 6016
rect 4404 5956 4408 6012
rect 4408 5956 4464 6012
rect 4464 5956 4468 6012
rect 4404 5952 4468 5956
rect 4484 6012 4548 6016
rect 4484 5956 4488 6012
rect 4488 5956 4544 6012
rect 4544 5956 4548 6012
rect 4484 5952 4548 5956
rect 4564 6012 4628 6016
rect 4564 5956 4568 6012
rect 4568 5956 4624 6012
rect 4624 5956 4628 6012
rect 4564 5952 4628 5956
rect 10724 6012 10788 6016
rect 10724 5956 10728 6012
rect 10728 5956 10784 6012
rect 10784 5956 10788 6012
rect 10724 5952 10788 5956
rect 10804 6012 10868 6016
rect 10804 5956 10808 6012
rect 10808 5956 10864 6012
rect 10864 5956 10868 6012
rect 10804 5952 10868 5956
rect 10884 6012 10948 6016
rect 10884 5956 10888 6012
rect 10888 5956 10944 6012
rect 10944 5956 10948 6012
rect 10884 5952 10948 5956
rect 10964 6012 11028 6016
rect 10964 5956 10968 6012
rect 10968 5956 11024 6012
rect 11024 5956 11028 6012
rect 10964 5952 11028 5956
rect 3664 5468 3728 5472
rect 3664 5412 3668 5468
rect 3668 5412 3724 5468
rect 3724 5412 3728 5468
rect 3664 5408 3728 5412
rect 3744 5468 3808 5472
rect 3744 5412 3748 5468
rect 3748 5412 3804 5468
rect 3804 5412 3808 5468
rect 3744 5408 3808 5412
rect 3824 5468 3888 5472
rect 3824 5412 3828 5468
rect 3828 5412 3884 5468
rect 3884 5412 3888 5468
rect 3824 5408 3888 5412
rect 3904 5468 3968 5472
rect 3904 5412 3908 5468
rect 3908 5412 3964 5468
rect 3964 5412 3968 5468
rect 3904 5408 3968 5412
rect 10064 5468 10128 5472
rect 10064 5412 10068 5468
rect 10068 5412 10124 5468
rect 10124 5412 10128 5468
rect 10064 5408 10128 5412
rect 10144 5468 10208 5472
rect 10144 5412 10148 5468
rect 10148 5412 10204 5468
rect 10204 5412 10208 5468
rect 10144 5408 10208 5412
rect 10224 5468 10288 5472
rect 10224 5412 10228 5468
rect 10228 5412 10284 5468
rect 10284 5412 10288 5468
rect 10224 5408 10288 5412
rect 10304 5468 10368 5472
rect 10304 5412 10308 5468
rect 10308 5412 10364 5468
rect 10364 5412 10368 5468
rect 10304 5408 10368 5412
rect 612 4932 676 4996
rect 4324 4924 4388 4928
rect 4324 4868 4328 4924
rect 4328 4868 4384 4924
rect 4384 4868 4388 4924
rect 4324 4864 4388 4868
rect 4404 4924 4468 4928
rect 4404 4868 4408 4924
rect 4408 4868 4464 4924
rect 4464 4868 4468 4924
rect 4404 4864 4468 4868
rect 4484 4924 4548 4928
rect 4484 4868 4488 4924
rect 4488 4868 4544 4924
rect 4544 4868 4548 4924
rect 4484 4864 4548 4868
rect 4564 4924 4628 4928
rect 4564 4868 4568 4924
rect 4568 4868 4624 4924
rect 4624 4868 4628 4924
rect 4564 4864 4628 4868
rect 10724 4924 10788 4928
rect 10724 4868 10728 4924
rect 10728 4868 10784 4924
rect 10784 4868 10788 4924
rect 10724 4864 10788 4868
rect 10804 4924 10868 4928
rect 10804 4868 10808 4924
rect 10808 4868 10864 4924
rect 10864 4868 10868 4924
rect 10804 4864 10868 4868
rect 10884 4924 10948 4928
rect 10884 4868 10888 4924
rect 10888 4868 10944 4924
rect 10944 4868 10948 4924
rect 10884 4864 10948 4868
rect 10964 4924 11028 4928
rect 10964 4868 10968 4924
rect 10968 4868 11024 4924
rect 11024 4868 11028 4924
rect 10964 4864 11028 4868
rect 3664 4380 3728 4384
rect 3664 4324 3668 4380
rect 3668 4324 3724 4380
rect 3724 4324 3728 4380
rect 3664 4320 3728 4324
rect 3744 4380 3808 4384
rect 3744 4324 3748 4380
rect 3748 4324 3804 4380
rect 3804 4324 3808 4380
rect 3744 4320 3808 4324
rect 3824 4380 3888 4384
rect 3824 4324 3828 4380
rect 3828 4324 3884 4380
rect 3884 4324 3888 4380
rect 3824 4320 3888 4324
rect 3904 4380 3968 4384
rect 3904 4324 3908 4380
rect 3908 4324 3964 4380
rect 3964 4324 3968 4380
rect 3904 4320 3968 4324
rect 10064 4380 10128 4384
rect 10064 4324 10068 4380
rect 10068 4324 10124 4380
rect 10124 4324 10128 4380
rect 10064 4320 10128 4324
rect 10144 4380 10208 4384
rect 10144 4324 10148 4380
rect 10148 4324 10204 4380
rect 10204 4324 10208 4380
rect 10144 4320 10208 4324
rect 10224 4380 10288 4384
rect 10224 4324 10228 4380
rect 10228 4324 10284 4380
rect 10284 4324 10288 4380
rect 10224 4320 10288 4324
rect 10304 4380 10368 4384
rect 10304 4324 10308 4380
rect 10308 4324 10364 4380
rect 10364 4324 10368 4380
rect 10304 4320 10368 4324
rect 4324 3836 4388 3840
rect 4324 3780 4328 3836
rect 4328 3780 4384 3836
rect 4384 3780 4388 3836
rect 4324 3776 4388 3780
rect 4404 3836 4468 3840
rect 4404 3780 4408 3836
rect 4408 3780 4464 3836
rect 4464 3780 4468 3836
rect 4404 3776 4468 3780
rect 4484 3836 4548 3840
rect 4484 3780 4488 3836
rect 4488 3780 4544 3836
rect 4544 3780 4548 3836
rect 4484 3776 4548 3780
rect 4564 3836 4628 3840
rect 4564 3780 4568 3836
rect 4568 3780 4624 3836
rect 4624 3780 4628 3836
rect 4564 3776 4628 3780
rect 10724 3836 10788 3840
rect 10724 3780 10728 3836
rect 10728 3780 10784 3836
rect 10784 3780 10788 3836
rect 10724 3776 10788 3780
rect 10804 3836 10868 3840
rect 10804 3780 10808 3836
rect 10808 3780 10864 3836
rect 10864 3780 10868 3836
rect 10804 3776 10868 3780
rect 10884 3836 10948 3840
rect 10884 3780 10888 3836
rect 10888 3780 10944 3836
rect 10944 3780 10948 3836
rect 10884 3776 10948 3780
rect 10964 3836 11028 3840
rect 10964 3780 10968 3836
rect 10968 3780 11024 3836
rect 11024 3780 11028 3836
rect 10964 3776 11028 3780
rect 3664 3292 3728 3296
rect 3664 3236 3668 3292
rect 3668 3236 3724 3292
rect 3724 3236 3728 3292
rect 3664 3232 3728 3236
rect 3744 3292 3808 3296
rect 3744 3236 3748 3292
rect 3748 3236 3804 3292
rect 3804 3236 3808 3292
rect 3744 3232 3808 3236
rect 3824 3292 3888 3296
rect 3824 3236 3828 3292
rect 3828 3236 3884 3292
rect 3884 3236 3888 3292
rect 3824 3232 3888 3236
rect 3904 3292 3968 3296
rect 3904 3236 3908 3292
rect 3908 3236 3964 3292
rect 3964 3236 3968 3292
rect 3904 3232 3968 3236
rect 10064 3292 10128 3296
rect 10064 3236 10068 3292
rect 10068 3236 10124 3292
rect 10124 3236 10128 3292
rect 10064 3232 10128 3236
rect 10144 3292 10208 3296
rect 10144 3236 10148 3292
rect 10148 3236 10204 3292
rect 10204 3236 10208 3292
rect 10144 3232 10208 3236
rect 10224 3292 10288 3296
rect 10224 3236 10228 3292
rect 10228 3236 10284 3292
rect 10284 3236 10288 3292
rect 10224 3232 10288 3236
rect 10304 3292 10368 3296
rect 10304 3236 10308 3292
rect 10308 3236 10364 3292
rect 10364 3236 10368 3292
rect 10304 3232 10368 3236
rect 4324 2748 4388 2752
rect 4324 2692 4328 2748
rect 4328 2692 4384 2748
rect 4384 2692 4388 2748
rect 4324 2688 4388 2692
rect 4404 2748 4468 2752
rect 4404 2692 4408 2748
rect 4408 2692 4464 2748
rect 4464 2692 4468 2748
rect 4404 2688 4468 2692
rect 4484 2748 4548 2752
rect 4484 2692 4488 2748
rect 4488 2692 4544 2748
rect 4544 2692 4548 2748
rect 4484 2688 4548 2692
rect 4564 2748 4628 2752
rect 4564 2692 4568 2748
rect 4568 2692 4624 2748
rect 4624 2692 4628 2748
rect 4564 2688 4628 2692
rect 10724 2748 10788 2752
rect 10724 2692 10728 2748
rect 10728 2692 10784 2748
rect 10784 2692 10788 2748
rect 10724 2688 10788 2692
rect 10804 2748 10868 2752
rect 10804 2692 10808 2748
rect 10808 2692 10864 2748
rect 10864 2692 10868 2748
rect 10804 2688 10868 2692
rect 10884 2748 10948 2752
rect 10884 2692 10888 2748
rect 10888 2692 10944 2748
rect 10944 2692 10948 2748
rect 10884 2688 10948 2692
rect 10964 2748 11028 2752
rect 10964 2692 10968 2748
rect 10968 2692 11024 2748
rect 11024 2692 11028 2748
rect 10964 2688 11028 2692
rect 9812 2484 9876 2548
rect 3664 2204 3728 2208
rect 3664 2148 3668 2204
rect 3668 2148 3724 2204
rect 3724 2148 3728 2204
rect 3664 2144 3728 2148
rect 3744 2204 3808 2208
rect 3744 2148 3748 2204
rect 3748 2148 3804 2204
rect 3804 2148 3808 2204
rect 3744 2144 3808 2148
rect 3824 2204 3888 2208
rect 3824 2148 3828 2204
rect 3828 2148 3884 2204
rect 3884 2148 3888 2204
rect 3824 2144 3888 2148
rect 3904 2204 3968 2208
rect 3904 2148 3908 2204
rect 3908 2148 3964 2204
rect 3964 2148 3968 2204
rect 3904 2144 3968 2148
rect 10064 2204 10128 2208
rect 10064 2148 10068 2204
rect 10068 2148 10124 2204
rect 10124 2148 10128 2204
rect 10064 2144 10128 2148
rect 10144 2204 10208 2208
rect 10144 2148 10148 2204
rect 10148 2148 10204 2204
rect 10204 2148 10208 2204
rect 10144 2144 10208 2148
rect 10224 2204 10288 2208
rect 10224 2148 10228 2204
rect 10228 2148 10284 2204
rect 10284 2148 10288 2204
rect 10224 2144 10288 2148
rect 10304 2204 10368 2208
rect 10304 2148 10308 2204
rect 10308 2148 10364 2204
rect 10364 2148 10368 2204
rect 10304 2144 10368 2148
rect 4324 1660 4388 1664
rect 4324 1604 4328 1660
rect 4328 1604 4384 1660
rect 4384 1604 4388 1660
rect 4324 1600 4388 1604
rect 4404 1660 4468 1664
rect 4404 1604 4408 1660
rect 4408 1604 4464 1660
rect 4464 1604 4468 1660
rect 4404 1600 4468 1604
rect 4484 1660 4548 1664
rect 4484 1604 4488 1660
rect 4488 1604 4544 1660
rect 4544 1604 4548 1660
rect 4484 1600 4548 1604
rect 4564 1660 4628 1664
rect 4564 1604 4568 1660
rect 4568 1604 4624 1660
rect 4624 1604 4628 1660
rect 4564 1600 4628 1604
rect 10724 1660 10788 1664
rect 10724 1604 10728 1660
rect 10728 1604 10784 1660
rect 10784 1604 10788 1660
rect 10724 1600 10788 1604
rect 10804 1660 10868 1664
rect 10804 1604 10808 1660
rect 10808 1604 10864 1660
rect 10864 1604 10868 1660
rect 10804 1600 10868 1604
rect 10884 1660 10948 1664
rect 10884 1604 10888 1660
rect 10888 1604 10944 1660
rect 10944 1604 10948 1660
rect 10884 1600 10948 1604
rect 10964 1660 11028 1664
rect 10964 1604 10968 1660
rect 10968 1604 11024 1660
rect 11024 1604 11028 1660
rect 10964 1600 11028 1604
rect 3664 1116 3728 1120
rect 3664 1060 3668 1116
rect 3668 1060 3724 1116
rect 3724 1060 3728 1116
rect 3664 1056 3728 1060
rect 3744 1116 3808 1120
rect 3744 1060 3748 1116
rect 3748 1060 3804 1116
rect 3804 1060 3808 1116
rect 3744 1056 3808 1060
rect 3824 1116 3888 1120
rect 3824 1060 3828 1116
rect 3828 1060 3884 1116
rect 3884 1060 3888 1116
rect 3824 1056 3888 1060
rect 3904 1116 3968 1120
rect 3904 1060 3908 1116
rect 3908 1060 3964 1116
rect 3964 1060 3968 1116
rect 3904 1056 3968 1060
rect 10064 1116 10128 1120
rect 10064 1060 10068 1116
rect 10068 1060 10124 1116
rect 10124 1060 10128 1116
rect 10064 1056 10128 1060
rect 10144 1116 10208 1120
rect 10144 1060 10148 1116
rect 10148 1060 10204 1116
rect 10204 1060 10208 1116
rect 10144 1056 10208 1060
rect 10224 1116 10288 1120
rect 10224 1060 10228 1116
rect 10228 1060 10284 1116
rect 10284 1060 10288 1116
rect 10224 1056 10288 1060
rect 10304 1116 10368 1120
rect 10304 1060 10308 1116
rect 10308 1060 10364 1116
rect 10364 1060 10368 1116
rect 10304 1056 10368 1060
rect 4324 572 4388 576
rect 4324 516 4328 572
rect 4328 516 4384 572
rect 4384 516 4388 572
rect 4324 512 4388 516
rect 4404 572 4468 576
rect 4404 516 4408 572
rect 4408 516 4464 572
rect 4464 516 4468 572
rect 4404 512 4468 516
rect 4484 572 4548 576
rect 4484 516 4488 572
rect 4488 516 4544 572
rect 4544 516 4548 572
rect 4484 512 4548 516
rect 4564 572 4628 576
rect 4564 516 4568 572
rect 4568 516 4624 572
rect 4624 516 4628 572
rect 4564 512 4628 516
rect 10724 572 10788 576
rect 10724 516 10728 572
rect 10728 516 10784 572
rect 10784 516 10788 572
rect 10724 512 10788 516
rect 10804 572 10868 576
rect 10804 516 10808 572
rect 10808 516 10864 572
rect 10864 516 10868 572
rect 10804 512 10868 516
rect 10884 572 10948 576
rect 10884 516 10888 572
rect 10888 516 10944 572
rect 10944 516 10948 572
rect 10884 512 10948 516
rect 10964 572 11028 576
rect 10964 516 10968 572
rect 10968 516 11024 572
rect 11024 516 11028 572
rect 10964 512 11028 516
<< metal4 >>
rect 1347 43620 1413 43621
rect 1347 43556 1348 43620
rect 1412 43556 1413 43620
rect 1347 43555 1413 43556
rect 5395 43620 5461 43621
rect 5395 43556 5396 43620
rect 5460 43556 5461 43620
rect 5395 43555 5461 43556
rect 5579 43620 5645 43621
rect 5579 43556 5580 43620
rect 5644 43556 5645 43620
rect 5579 43555 5645 43556
rect 8155 43620 8221 43621
rect 8155 43556 8156 43620
rect 8220 43556 8221 43620
rect 8155 43555 8221 43556
rect 9259 43620 9325 43621
rect 9259 43556 9260 43620
rect 9324 43556 9325 43620
rect 9259 43555 9325 43556
rect 9627 43620 9693 43621
rect 9627 43556 9628 43620
rect 9692 43556 9693 43620
rect 9627 43555 9693 43556
rect 381 41716 447 41717
rect 381 41714 382 41716
rect 62 41654 382 41714
rect 62 29749 122 41654
rect 381 41652 382 41654
rect 446 41652 447 41716
rect 381 41651 447 41652
rect 1163 41036 1229 41037
rect 1163 40972 1164 41036
rect 1228 40972 1229 41036
rect 1163 40971 1229 40972
rect 979 37636 1045 37637
rect 979 37572 980 37636
rect 1044 37572 1045 37636
rect 979 37571 1045 37572
rect 795 32332 861 32333
rect 795 32268 796 32332
rect 860 32268 861 32332
rect 795 32267 861 32268
rect 59 29748 125 29749
rect 59 29684 60 29748
rect 124 29684 125 29748
rect 59 29683 125 29684
rect 611 28252 677 28253
rect 611 28188 612 28252
rect 676 28188 677 28252
rect 611 28187 677 28188
rect 427 17780 493 17781
rect 427 17716 428 17780
rect 492 17716 493 17780
rect 427 17715 493 17716
rect 59 15468 125 15469
rect 59 15404 60 15468
rect 124 15404 125 15468
rect 59 15403 125 15404
rect 62 7173 122 15403
rect 430 12450 490 17715
rect 614 15877 674 28187
rect 798 20773 858 32267
rect 982 29205 1042 37571
rect 1166 35050 1226 40971
rect 1350 36957 1410 43555
rect 3656 42464 3976 43024
rect 3656 42400 3664 42464
rect 3728 42400 3744 42464
rect 3808 42400 3824 42464
rect 3888 42400 3904 42464
rect 3968 42400 3976 42464
rect 3371 41580 3437 41581
rect 3371 41516 3372 41580
rect 3436 41516 3437 41580
rect 3371 41515 3437 41516
rect 3187 40220 3253 40221
rect 3187 40156 3188 40220
rect 3252 40156 3253 40220
rect 3187 40155 3253 40156
rect 2083 39948 2149 39949
rect 2083 39884 2084 39948
rect 2148 39884 2149 39948
rect 2083 39883 2149 39884
rect 1531 38860 1597 38861
rect 1531 38796 1532 38860
rect 1596 38796 1597 38860
rect 1531 38795 1597 38796
rect 1347 36956 1413 36957
rect 1347 36892 1348 36956
rect 1412 36892 1413 36956
rect 1347 36891 1413 36892
rect 1166 34990 1410 35050
rect 1163 34372 1229 34373
rect 1163 34308 1164 34372
rect 1228 34308 1229 34372
rect 1163 34307 1229 34308
rect 979 29204 1045 29205
rect 979 29140 980 29204
rect 1044 29140 1045 29204
rect 979 29139 1045 29140
rect 1166 26890 1226 34307
rect 1350 32333 1410 34990
rect 1534 33557 1594 38795
rect 1715 38588 1781 38589
rect 1715 38524 1716 38588
rect 1780 38524 1781 38588
rect 1715 38523 1781 38524
rect 1531 33556 1597 33557
rect 1531 33492 1532 33556
rect 1596 33492 1597 33556
rect 1531 33491 1597 33492
rect 1347 32332 1413 32333
rect 1347 32268 1348 32332
rect 1412 32268 1413 32332
rect 1347 32267 1413 32268
rect 1347 32196 1413 32197
rect 1347 32132 1348 32196
rect 1412 32132 1413 32196
rect 1347 32131 1413 32132
rect 982 26830 1226 26890
rect 795 20772 861 20773
rect 795 20708 796 20772
rect 860 20708 861 20772
rect 795 20707 861 20708
rect 982 16149 1042 26830
rect 1163 25396 1229 25397
rect 1163 25332 1164 25396
rect 1228 25332 1229 25396
rect 1163 25331 1229 25332
rect 1166 16557 1226 25331
rect 1350 23901 1410 32131
rect 1718 31653 1778 38523
rect 1899 38180 1965 38181
rect 1899 38116 1900 38180
rect 1964 38116 1965 38180
rect 1899 38115 1965 38116
rect 1902 37093 1962 38115
rect 1899 37092 1965 37093
rect 1899 37028 1900 37092
rect 1964 37028 1965 37092
rect 1899 37027 1965 37028
rect 1899 35052 1965 35053
rect 1899 34988 1900 35052
rect 1964 34988 1965 35052
rect 1899 34987 1965 34988
rect 1715 31652 1781 31653
rect 1715 31588 1716 31652
rect 1780 31588 1781 31652
rect 1715 31587 1781 31588
rect 1715 31516 1781 31517
rect 1715 31452 1716 31516
rect 1780 31452 1781 31516
rect 1715 31451 1781 31452
rect 1718 28525 1778 31451
rect 1902 29885 1962 34987
rect 2086 33693 2146 39883
rect 2267 37772 2333 37773
rect 2267 37708 2268 37772
rect 2332 37708 2333 37772
rect 2267 37707 2333 37708
rect 2083 33692 2149 33693
rect 2083 33628 2084 33692
rect 2148 33628 2149 33692
rect 2083 33627 2149 33628
rect 2083 33420 2149 33421
rect 2083 33356 2084 33420
rect 2148 33356 2149 33420
rect 2083 33355 2149 33356
rect 1899 29884 1965 29885
rect 1899 29820 1900 29884
rect 1964 29820 1965 29884
rect 1899 29819 1965 29820
rect 1715 28524 1781 28525
rect 1715 28460 1716 28524
rect 1780 28460 1781 28524
rect 1715 28459 1781 28460
rect 1715 27844 1781 27845
rect 1715 27780 1716 27844
rect 1780 27780 1781 27844
rect 1715 27779 1781 27780
rect 1347 23900 1413 23901
rect 1347 23836 1348 23900
rect 1412 23836 1413 23900
rect 1347 23835 1413 23836
rect 1350 20637 1410 23835
rect 1347 20636 1413 20637
rect 1347 20572 1348 20636
rect 1412 20572 1413 20636
rect 1347 20571 1413 20572
rect 1347 20228 1413 20229
rect 1347 20164 1348 20228
rect 1412 20164 1413 20228
rect 1347 20163 1413 20164
rect 1163 16556 1229 16557
rect 1163 16492 1164 16556
rect 1228 16492 1229 16556
rect 1163 16491 1229 16492
rect 1350 16421 1410 20163
rect 1347 16420 1413 16421
rect 1347 16356 1348 16420
rect 1412 16356 1413 16420
rect 1347 16355 1413 16356
rect 979 16148 1045 16149
rect 979 16084 980 16148
rect 1044 16084 1045 16148
rect 979 16083 1045 16084
rect 611 15876 677 15877
rect 611 15812 612 15876
rect 676 15812 677 15876
rect 611 15811 677 15812
rect 1718 15741 1778 27779
rect 2086 26621 2146 33355
rect 2270 31789 2330 37707
rect 2635 37364 2701 37365
rect 2635 37300 2636 37364
rect 2700 37300 2701 37364
rect 2635 37299 2701 37300
rect 2451 33284 2517 33285
rect 2451 33220 2452 33284
rect 2516 33220 2517 33284
rect 2451 33219 2517 33220
rect 2267 31788 2333 31789
rect 2267 31724 2268 31788
rect 2332 31724 2333 31788
rect 2267 31723 2333 31724
rect 2267 30428 2333 30429
rect 2267 30364 2268 30428
rect 2332 30364 2333 30428
rect 2267 30363 2333 30364
rect 2270 29613 2330 30363
rect 2267 29612 2333 29613
rect 2267 29548 2268 29612
rect 2332 29548 2333 29612
rect 2267 29547 2333 29548
rect 2454 27709 2514 33219
rect 2638 29205 2698 37299
rect 3003 35324 3069 35325
rect 3003 35260 3004 35324
rect 3068 35260 3069 35324
rect 3003 35259 3069 35260
rect 2819 33420 2885 33421
rect 2819 33356 2820 33420
rect 2884 33356 2885 33420
rect 2819 33355 2885 33356
rect 2822 29341 2882 33355
rect 2819 29340 2885 29341
rect 2819 29276 2820 29340
rect 2884 29276 2885 29340
rect 2819 29275 2885 29276
rect 2635 29204 2701 29205
rect 2635 29140 2636 29204
rect 2700 29140 2701 29204
rect 2635 29139 2701 29140
rect 3006 28933 3066 35259
rect 3190 32469 3250 40155
rect 3374 35461 3434 41515
rect 3656 41376 3976 42400
rect 3656 41312 3664 41376
rect 3728 41312 3744 41376
rect 3808 41312 3824 41376
rect 3888 41312 3904 41376
rect 3968 41312 3976 41376
rect 3656 40288 3976 41312
rect 3656 40224 3664 40288
rect 3728 40224 3744 40288
rect 3808 40224 3824 40288
rect 3888 40224 3904 40288
rect 3968 40224 3976 40288
rect 3656 39200 3976 40224
rect 4316 43008 4636 43024
rect 4316 42944 4324 43008
rect 4388 42944 4404 43008
rect 4468 42944 4484 43008
rect 4548 42944 4564 43008
rect 4628 42944 4636 43008
rect 4316 41920 4636 42944
rect 4316 41856 4324 41920
rect 4388 41856 4404 41920
rect 4468 41856 4484 41920
rect 4548 41856 4564 41920
rect 4628 41856 4636 41920
rect 4316 40832 4636 41856
rect 4316 40768 4324 40832
rect 4388 40768 4404 40832
rect 4468 40768 4484 40832
rect 4548 40768 4564 40832
rect 4628 40768 4636 40832
rect 4107 40084 4173 40085
rect 4107 40020 4108 40084
rect 4172 40020 4173 40084
rect 4107 40019 4173 40020
rect 3656 39136 3664 39200
rect 3728 39136 3744 39200
rect 3808 39136 3824 39200
rect 3888 39136 3904 39200
rect 3968 39136 3976 39200
rect 3656 38112 3976 39136
rect 3656 38048 3664 38112
rect 3728 38048 3744 38112
rect 3808 38048 3824 38112
rect 3888 38048 3904 38112
rect 3968 38048 3976 38112
rect 3656 37024 3976 38048
rect 4110 37365 4170 40019
rect 4316 39744 4636 40768
rect 5211 40764 5277 40765
rect 5211 40700 5212 40764
rect 5276 40700 5277 40764
rect 5211 40699 5277 40700
rect 4316 39680 4324 39744
rect 4388 39680 4404 39744
rect 4468 39680 4484 39744
rect 4548 39680 4564 39744
rect 4628 39680 4636 39744
rect 4316 38656 4636 39680
rect 4843 39404 4909 39405
rect 4843 39340 4844 39404
rect 4908 39340 4909 39404
rect 4843 39339 4909 39340
rect 4316 38592 4324 38656
rect 4388 38592 4404 38656
rect 4468 38592 4484 38656
rect 4548 38592 4564 38656
rect 4628 38592 4636 38656
rect 4316 37568 4636 38592
rect 4316 37504 4324 37568
rect 4388 37504 4404 37568
rect 4468 37504 4484 37568
rect 4548 37504 4564 37568
rect 4628 37504 4636 37568
rect 4107 37364 4173 37365
rect 4107 37300 4108 37364
rect 4172 37300 4173 37364
rect 4107 37299 4173 37300
rect 3656 36960 3664 37024
rect 3728 36960 3744 37024
rect 3808 36960 3824 37024
rect 3888 36960 3904 37024
rect 3968 36960 3976 37024
rect 3656 35936 3976 36960
rect 3656 35872 3664 35936
rect 3728 35872 3744 35936
rect 3808 35872 3824 35936
rect 3888 35872 3904 35936
rect 3968 35872 3976 35936
rect 3371 35460 3437 35461
rect 3371 35396 3372 35460
rect 3436 35396 3437 35460
rect 3371 35395 3437 35396
rect 3187 32468 3253 32469
rect 3187 32404 3188 32468
rect 3252 32404 3253 32468
rect 3187 32403 3253 32404
rect 3374 31770 3434 35395
rect 3190 31710 3434 31770
rect 3656 34848 3976 35872
rect 3656 34784 3664 34848
rect 3728 34784 3744 34848
rect 3808 34784 3824 34848
rect 3888 34784 3904 34848
rect 3968 34784 3976 34848
rect 3656 33760 3976 34784
rect 4110 34509 4170 37299
rect 4316 36480 4636 37504
rect 4316 36416 4324 36480
rect 4388 36416 4404 36480
rect 4468 36416 4484 36480
rect 4548 36416 4564 36480
rect 4628 36416 4636 36480
rect 4316 35392 4636 36416
rect 4316 35328 4324 35392
rect 4388 35328 4404 35392
rect 4468 35328 4484 35392
rect 4548 35328 4564 35392
rect 4628 35328 4636 35392
rect 4107 34508 4173 34509
rect 4107 34444 4108 34508
rect 4172 34444 4173 34508
rect 4107 34443 4173 34444
rect 4316 34304 4636 35328
rect 4846 34645 4906 39339
rect 5214 39269 5274 40699
rect 5398 39949 5458 43555
rect 5395 39948 5461 39949
rect 5395 39884 5396 39948
rect 5460 39884 5461 39948
rect 5395 39883 5461 39884
rect 5211 39268 5277 39269
rect 5211 39204 5212 39268
rect 5276 39204 5277 39268
rect 5211 39203 5277 39204
rect 5214 38670 5274 39203
rect 5214 38610 5458 38670
rect 5211 37500 5277 37501
rect 5211 37436 5212 37500
rect 5276 37436 5277 37500
rect 5211 37435 5277 37436
rect 5027 36820 5093 36821
rect 5027 36756 5028 36820
rect 5092 36756 5093 36820
rect 5027 36755 5093 36756
rect 4843 34644 4909 34645
rect 4843 34580 4844 34644
rect 4908 34580 4909 34644
rect 4843 34579 4909 34580
rect 4316 34240 4324 34304
rect 4388 34240 4404 34304
rect 4468 34240 4484 34304
rect 4548 34240 4564 34304
rect 4628 34240 4636 34304
rect 4107 34236 4173 34237
rect 4107 34172 4108 34236
rect 4172 34172 4173 34236
rect 4107 34171 4173 34172
rect 3656 33696 3664 33760
rect 3728 33696 3744 33760
rect 3808 33696 3824 33760
rect 3888 33696 3904 33760
rect 3968 33696 3976 33760
rect 3656 32672 3976 33696
rect 3656 32608 3664 32672
rect 3728 32608 3744 32672
rect 3808 32608 3824 32672
rect 3888 32608 3904 32672
rect 3968 32608 3976 32672
rect 3003 28932 3069 28933
rect 3003 28868 3004 28932
rect 3068 28868 3069 28932
rect 3003 28867 3069 28868
rect 2267 27708 2333 27709
rect 2267 27644 2268 27708
rect 2332 27644 2333 27708
rect 2267 27643 2333 27644
rect 2451 27708 2517 27709
rect 2451 27644 2452 27708
rect 2516 27644 2517 27708
rect 2451 27643 2517 27644
rect 2083 26620 2149 26621
rect 2083 26556 2084 26620
rect 2148 26556 2149 26620
rect 2083 26555 2149 26556
rect 2083 26348 2149 26349
rect 2083 26284 2084 26348
rect 2148 26284 2149 26348
rect 2083 26283 2149 26284
rect 1899 24172 1965 24173
rect 1899 24108 1900 24172
rect 1964 24108 1965 24172
rect 1899 24107 1965 24108
rect 1902 20093 1962 24107
rect 1899 20092 1965 20093
rect 1899 20028 1900 20092
rect 1964 20028 1965 20092
rect 1899 20027 1965 20028
rect 1715 15740 1781 15741
rect 1715 15676 1716 15740
rect 1780 15676 1781 15740
rect 1715 15675 1781 15676
rect 430 12390 674 12450
rect 59 7172 125 7173
rect 59 7108 60 7172
rect 124 7108 125 7172
rect 59 7107 125 7108
rect 614 4997 674 12390
rect 2086 11253 2146 26283
rect 2270 23357 2330 27643
rect 2451 25532 2517 25533
rect 2451 25468 2452 25532
rect 2516 25468 2517 25532
rect 2451 25467 2517 25468
rect 2267 23356 2333 23357
rect 2267 23292 2268 23356
rect 2332 23292 2333 23356
rect 2267 23291 2333 23292
rect 2454 20634 2514 25467
rect 2635 23764 2701 23765
rect 2635 23700 2636 23764
rect 2700 23700 2701 23764
rect 2635 23699 2701 23700
rect 2270 20574 2514 20634
rect 2270 19277 2330 20574
rect 2451 20364 2517 20365
rect 2451 20300 2452 20364
rect 2516 20300 2517 20364
rect 2451 20299 2517 20300
rect 2454 19957 2514 20299
rect 2638 20229 2698 23699
rect 3006 22677 3066 28867
rect 3190 23085 3250 31710
rect 3656 31584 3976 32608
rect 3656 31520 3664 31584
rect 3728 31520 3744 31584
rect 3808 31520 3824 31584
rect 3888 31520 3904 31584
rect 3968 31520 3976 31584
rect 3371 31108 3437 31109
rect 3371 31044 3372 31108
rect 3436 31044 3437 31108
rect 3371 31043 3437 31044
rect 3374 30021 3434 31043
rect 3656 30496 3976 31520
rect 4110 31517 4170 34171
rect 4316 33216 4636 34240
rect 4843 33420 4909 33421
rect 4843 33356 4844 33420
rect 4908 33356 4909 33420
rect 4843 33355 4909 33356
rect 4316 33152 4324 33216
rect 4388 33152 4404 33216
rect 4468 33152 4484 33216
rect 4548 33152 4564 33216
rect 4628 33152 4636 33216
rect 4316 32128 4636 33152
rect 4316 32064 4324 32128
rect 4388 32064 4404 32128
rect 4468 32064 4484 32128
rect 4548 32064 4564 32128
rect 4628 32064 4636 32128
rect 4107 31516 4173 31517
rect 4107 31452 4108 31516
rect 4172 31452 4173 31516
rect 4107 31451 4173 31452
rect 4107 31380 4173 31381
rect 4107 31316 4108 31380
rect 4172 31316 4173 31380
rect 4107 31315 4173 31316
rect 3656 30432 3664 30496
rect 3728 30432 3744 30496
rect 3808 30432 3824 30496
rect 3888 30432 3904 30496
rect 3968 30432 3976 30496
rect 3371 30020 3437 30021
rect 3371 29956 3372 30020
rect 3436 29956 3437 30020
rect 3371 29955 3437 29956
rect 3374 25941 3434 29955
rect 3656 29408 3976 30432
rect 3656 29344 3664 29408
rect 3728 29344 3744 29408
rect 3808 29344 3824 29408
rect 3888 29344 3904 29408
rect 3968 29344 3976 29408
rect 3656 28320 3976 29344
rect 3656 28256 3664 28320
rect 3728 28256 3744 28320
rect 3808 28256 3824 28320
rect 3888 28256 3904 28320
rect 3968 28256 3976 28320
rect 3656 27232 3976 28256
rect 3656 27168 3664 27232
rect 3728 27168 3744 27232
rect 3808 27168 3824 27232
rect 3888 27168 3904 27232
rect 3968 27168 3976 27232
rect 3656 26144 3976 27168
rect 3656 26080 3664 26144
rect 3728 26080 3744 26144
rect 3808 26080 3824 26144
rect 3888 26080 3904 26144
rect 3968 26080 3976 26144
rect 3371 25940 3437 25941
rect 3371 25876 3372 25940
rect 3436 25876 3437 25940
rect 3371 25875 3437 25876
rect 3656 25056 3976 26080
rect 3656 24992 3664 25056
rect 3728 24992 3744 25056
rect 3808 24992 3824 25056
rect 3888 24992 3904 25056
rect 3968 24992 3976 25056
rect 3371 24580 3437 24581
rect 3371 24516 3372 24580
rect 3436 24516 3437 24580
rect 3371 24515 3437 24516
rect 3187 23084 3253 23085
rect 3187 23020 3188 23084
rect 3252 23020 3253 23084
rect 3187 23019 3253 23020
rect 3003 22676 3069 22677
rect 3003 22612 3004 22676
rect 3068 22612 3069 22676
rect 3003 22611 3069 22612
rect 2819 22132 2885 22133
rect 2819 22068 2820 22132
rect 2884 22068 2885 22132
rect 2819 22067 2885 22068
rect 2635 20228 2701 20229
rect 2635 20164 2636 20228
rect 2700 20164 2701 20228
rect 2635 20163 2701 20164
rect 2822 20090 2882 22067
rect 3190 21589 3250 23019
rect 3187 21588 3253 21589
rect 3187 21524 3188 21588
rect 3252 21524 3253 21588
rect 3187 21523 3253 21524
rect 3003 21452 3069 21453
rect 3003 21388 3004 21452
rect 3068 21388 3069 21452
rect 3003 21387 3069 21388
rect 2638 20030 2882 20090
rect 2451 19956 2517 19957
rect 2451 19892 2452 19956
rect 2516 19892 2517 19956
rect 2451 19891 2517 19892
rect 2267 19276 2333 19277
rect 2267 19212 2268 19276
rect 2332 19212 2333 19276
rect 2267 19211 2333 19212
rect 2270 17101 2330 19211
rect 2267 17100 2333 17101
rect 2267 17036 2268 17100
rect 2332 17036 2333 17100
rect 2267 17035 2333 17036
rect 2638 16829 2698 20030
rect 2819 19004 2885 19005
rect 2819 18940 2820 19004
rect 2884 18940 2885 19004
rect 2819 18939 2885 18940
rect 2822 17101 2882 18939
rect 2819 17100 2885 17101
rect 2819 17036 2820 17100
rect 2884 17036 2885 17100
rect 2819 17035 2885 17036
rect 2635 16828 2701 16829
rect 2635 16764 2636 16828
rect 2700 16764 2701 16828
rect 2635 16763 2701 16764
rect 3006 16590 3066 21387
rect 3187 21180 3253 21181
rect 3187 21116 3188 21180
rect 3252 21116 3253 21180
rect 3187 21115 3253 21116
rect 3190 17781 3250 21115
rect 3374 18869 3434 24515
rect 3656 23968 3976 24992
rect 3656 23904 3664 23968
rect 3728 23904 3744 23968
rect 3808 23904 3824 23968
rect 3888 23904 3904 23968
rect 3968 23904 3976 23968
rect 3656 22880 3976 23904
rect 4110 23765 4170 31315
rect 4316 31040 4636 32064
rect 4316 30976 4324 31040
rect 4388 30976 4404 31040
rect 4468 30976 4484 31040
rect 4548 30976 4564 31040
rect 4628 30976 4636 31040
rect 4316 29952 4636 30976
rect 4316 29888 4324 29952
rect 4388 29888 4404 29952
rect 4468 29888 4484 29952
rect 4548 29888 4564 29952
rect 4628 29888 4636 29952
rect 4316 28864 4636 29888
rect 4316 28800 4324 28864
rect 4388 28800 4404 28864
rect 4468 28800 4484 28864
rect 4548 28800 4564 28864
rect 4628 28800 4636 28864
rect 4316 27776 4636 28800
rect 4316 27712 4324 27776
rect 4388 27712 4404 27776
rect 4468 27712 4484 27776
rect 4548 27712 4564 27776
rect 4628 27712 4636 27776
rect 4316 26688 4636 27712
rect 4316 26624 4324 26688
rect 4388 26624 4404 26688
rect 4468 26624 4484 26688
rect 4548 26624 4564 26688
rect 4628 26624 4636 26688
rect 4316 25600 4636 26624
rect 4316 25536 4324 25600
rect 4388 25536 4404 25600
rect 4468 25536 4484 25600
rect 4548 25536 4564 25600
rect 4628 25536 4636 25600
rect 4316 24512 4636 25536
rect 4846 25261 4906 33355
rect 5030 30565 5090 36755
rect 5214 33693 5274 37435
rect 5211 33692 5277 33693
rect 5211 33628 5212 33692
rect 5276 33628 5277 33692
rect 5211 33627 5277 33628
rect 5211 33556 5277 33557
rect 5211 33492 5212 33556
rect 5276 33492 5277 33556
rect 5211 33491 5277 33492
rect 5027 30564 5093 30565
rect 5027 30500 5028 30564
rect 5092 30500 5093 30564
rect 5027 30499 5093 30500
rect 5027 30292 5093 30293
rect 5027 30228 5028 30292
rect 5092 30228 5093 30292
rect 5027 30227 5093 30228
rect 4843 25260 4909 25261
rect 4843 25196 4844 25260
rect 4908 25196 4909 25260
rect 4843 25195 4909 25196
rect 4316 24448 4324 24512
rect 4388 24448 4404 24512
rect 4468 24448 4484 24512
rect 4548 24448 4564 24512
rect 4628 24448 4636 24512
rect 4107 23764 4173 23765
rect 4107 23700 4108 23764
rect 4172 23700 4173 23764
rect 4107 23699 4173 23700
rect 4107 23628 4173 23629
rect 4107 23564 4108 23628
rect 4172 23564 4173 23628
rect 4107 23563 4173 23564
rect 3656 22816 3664 22880
rect 3728 22816 3744 22880
rect 3808 22816 3824 22880
rect 3888 22816 3904 22880
rect 3968 22816 3976 22880
rect 3656 21792 3976 22816
rect 4110 22133 4170 23563
rect 4316 23424 4636 24448
rect 4316 23360 4324 23424
rect 4388 23360 4404 23424
rect 4468 23360 4484 23424
rect 4548 23360 4564 23424
rect 4628 23360 4636 23424
rect 4316 22336 4636 23360
rect 4843 22812 4909 22813
rect 4843 22748 4844 22812
rect 4908 22748 4909 22812
rect 4843 22747 4909 22748
rect 4316 22272 4324 22336
rect 4388 22272 4404 22336
rect 4468 22272 4484 22336
rect 4548 22272 4564 22336
rect 4628 22272 4636 22336
rect 4107 22132 4173 22133
rect 4107 22068 4108 22132
rect 4172 22068 4173 22132
rect 4107 22067 4173 22068
rect 3656 21728 3664 21792
rect 3728 21728 3744 21792
rect 3808 21728 3824 21792
rect 3888 21728 3904 21792
rect 3968 21728 3976 21792
rect 3656 20704 3976 21728
rect 3656 20640 3664 20704
rect 3728 20640 3744 20704
rect 3808 20640 3824 20704
rect 3888 20640 3904 20704
rect 3968 20640 3976 20704
rect 3656 19616 3976 20640
rect 4316 21248 4636 22272
rect 4316 21184 4324 21248
rect 4388 21184 4404 21248
rect 4468 21184 4484 21248
rect 4548 21184 4564 21248
rect 4628 21184 4636 21248
rect 4107 20636 4173 20637
rect 4107 20572 4108 20636
rect 4172 20572 4173 20636
rect 4107 20571 4173 20572
rect 3656 19552 3664 19616
rect 3728 19552 3744 19616
rect 3808 19552 3824 19616
rect 3888 19552 3904 19616
rect 3968 19552 3976 19616
rect 3371 18868 3437 18869
rect 3371 18804 3372 18868
rect 3436 18804 3437 18868
rect 3371 18803 3437 18804
rect 3371 18732 3437 18733
rect 3371 18668 3372 18732
rect 3436 18668 3437 18732
rect 3371 18667 3437 18668
rect 3187 17780 3253 17781
rect 3187 17716 3188 17780
rect 3252 17716 3253 17780
rect 3187 17715 3253 17716
rect 3187 16692 3253 16693
rect 3187 16628 3188 16692
rect 3252 16628 3253 16692
rect 3187 16627 3253 16628
rect 2638 16530 3066 16590
rect 2638 15469 2698 16530
rect 2635 15468 2701 15469
rect 2635 15404 2636 15468
rect 2700 15404 2701 15468
rect 2635 15403 2701 15404
rect 3190 15333 3250 16627
rect 3187 15332 3253 15333
rect 3187 15268 3188 15332
rect 3252 15268 3253 15332
rect 3187 15267 3253 15268
rect 3374 14925 3434 18667
rect 3656 18528 3976 19552
rect 4110 19005 4170 20571
rect 4316 20160 4636 21184
rect 4316 20096 4324 20160
rect 4388 20096 4404 20160
rect 4468 20096 4484 20160
rect 4548 20096 4564 20160
rect 4628 20096 4636 20160
rect 4316 19072 4636 20096
rect 4846 19685 4906 22747
rect 5030 22541 5090 30227
rect 5214 29885 5274 33491
rect 5398 32877 5458 38610
rect 5582 37365 5642 43555
rect 6499 41580 6565 41581
rect 6499 41516 6500 41580
rect 6564 41516 6565 41580
rect 6499 41515 6565 41516
rect 5947 40220 6013 40221
rect 5947 40156 5948 40220
rect 6012 40156 6013 40220
rect 5947 40155 6013 40156
rect 5763 40084 5829 40085
rect 5763 40020 5764 40084
rect 5828 40020 5829 40084
rect 5763 40019 5829 40020
rect 5579 37364 5645 37365
rect 5579 37300 5580 37364
rect 5644 37300 5645 37364
rect 5579 37299 5645 37300
rect 5579 36004 5645 36005
rect 5579 35940 5580 36004
rect 5644 35940 5645 36004
rect 5579 35939 5645 35940
rect 5395 32876 5461 32877
rect 5395 32812 5396 32876
rect 5460 32812 5461 32876
rect 5395 32811 5461 32812
rect 5395 32468 5461 32469
rect 5395 32404 5396 32468
rect 5460 32404 5461 32468
rect 5395 32403 5461 32404
rect 5211 29884 5277 29885
rect 5211 29820 5212 29884
rect 5276 29820 5277 29884
rect 5211 29819 5277 29820
rect 5211 28932 5277 28933
rect 5211 28868 5212 28932
rect 5276 28868 5277 28932
rect 5211 28867 5277 28868
rect 5027 22540 5093 22541
rect 5027 22476 5028 22540
rect 5092 22476 5093 22540
rect 5027 22475 5093 22476
rect 5027 22268 5093 22269
rect 5027 22204 5028 22268
rect 5092 22204 5093 22268
rect 5027 22203 5093 22204
rect 4843 19684 4909 19685
rect 4843 19620 4844 19684
rect 4908 19620 4909 19684
rect 4843 19619 4909 19620
rect 4843 19548 4909 19549
rect 4843 19484 4844 19548
rect 4908 19484 4909 19548
rect 4843 19483 4909 19484
rect 4316 19008 4324 19072
rect 4388 19008 4404 19072
rect 4468 19008 4484 19072
rect 4548 19008 4564 19072
rect 4628 19008 4636 19072
rect 4107 19004 4173 19005
rect 4107 18940 4108 19004
rect 4172 18940 4173 19004
rect 4107 18939 4173 18940
rect 4107 18732 4173 18733
rect 4107 18668 4108 18732
rect 4172 18668 4173 18732
rect 4107 18667 4173 18668
rect 3656 18464 3664 18528
rect 3728 18464 3744 18528
rect 3808 18464 3824 18528
rect 3888 18464 3904 18528
rect 3968 18464 3976 18528
rect 3656 17440 3976 18464
rect 3656 17376 3664 17440
rect 3728 17376 3744 17440
rect 3808 17376 3824 17440
rect 3888 17376 3904 17440
rect 3968 17376 3976 17440
rect 3656 16352 3976 17376
rect 3656 16288 3664 16352
rect 3728 16288 3744 16352
rect 3808 16288 3824 16352
rect 3888 16288 3904 16352
rect 3968 16288 3976 16352
rect 3656 15264 3976 16288
rect 4110 16285 4170 18667
rect 4316 17984 4636 19008
rect 4316 17920 4324 17984
rect 4388 17920 4404 17984
rect 4468 17920 4484 17984
rect 4548 17920 4564 17984
rect 4628 17920 4636 17984
rect 4316 16896 4636 17920
rect 4316 16832 4324 16896
rect 4388 16832 4404 16896
rect 4468 16832 4484 16896
rect 4548 16832 4564 16896
rect 4628 16832 4636 16896
rect 4107 16284 4173 16285
rect 4107 16220 4108 16284
rect 4172 16220 4173 16284
rect 4107 16219 4173 16220
rect 3656 15200 3664 15264
rect 3728 15200 3744 15264
rect 3808 15200 3824 15264
rect 3888 15200 3904 15264
rect 3968 15200 3976 15264
rect 3371 14924 3437 14925
rect 3371 14860 3372 14924
rect 3436 14860 3437 14924
rect 3371 14859 3437 14860
rect 3656 14176 3976 15200
rect 3656 14112 3664 14176
rect 3728 14112 3744 14176
rect 3808 14112 3824 14176
rect 3888 14112 3904 14176
rect 3968 14112 3976 14176
rect 3656 13088 3976 14112
rect 3656 13024 3664 13088
rect 3728 13024 3744 13088
rect 3808 13024 3824 13088
rect 3888 13024 3904 13088
rect 3968 13024 3976 13088
rect 3656 12000 3976 13024
rect 3656 11936 3664 12000
rect 3728 11936 3744 12000
rect 3808 11936 3824 12000
rect 3888 11936 3904 12000
rect 3968 11936 3976 12000
rect 2083 11252 2149 11253
rect 2083 11188 2084 11252
rect 2148 11188 2149 11252
rect 2083 11187 2149 11188
rect 3656 10912 3976 11936
rect 3656 10848 3664 10912
rect 3728 10848 3744 10912
rect 3808 10848 3824 10912
rect 3888 10848 3904 10912
rect 3968 10848 3976 10912
rect 3656 9824 3976 10848
rect 3656 9760 3664 9824
rect 3728 9760 3744 9824
rect 3808 9760 3824 9824
rect 3888 9760 3904 9824
rect 3968 9760 3976 9824
rect 3656 8736 3976 9760
rect 3656 8672 3664 8736
rect 3728 8672 3744 8736
rect 3808 8672 3824 8736
rect 3888 8672 3904 8736
rect 3968 8672 3976 8736
rect 3656 7648 3976 8672
rect 3656 7584 3664 7648
rect 3728 7584 3744 7648
rect 3808 7584 3824 7648
rect 3888 7584 3904 7648
rect 3968 7584 3976 7648
rect 3656 6560 3976 7584
rect 3656 6496 3664 6560
rect 3728 6496 3744 6560
rect 3808 6496 3824 6560
rect 3888 6496 3904 6560
rect 3968 6496 3976 6560
rect 3656 5472 3976 6496
rect 3656 5408 3664 5472
rect 3728 5408 3744 5472
rect 3808 5408 3824 5472
rect 3888 5408 3904 5472
rect 3968 5408 3976 5472
rect 611 4996 677 4997
rect 611 4932 612 4996
rect 676 4932 677 4996
rect 611 4931 677 4932
rect 3656 4384 3976 5408
rect 3656 4320 3664 4384
rect 3728 4320 3744 4384
rect 3808 4320 3824 4384
rect 3888 4320 3904 4384
rect 3968 4320 3976 4384
rect 3656 3296 3976 4320
rect 3656 3232 3664 3296
rect 3728 3232 3744 3296
rect 3808 3232 3824 3296
rect 3888 3232 3904 3296
rect 3968 3232 3976 3296
rect 3656 2208 3976 3232
rect 3656 2144 3664 2208
rect 3728 2144 3744 2208
rect 3808 2144 3824 2208
rect 3888 2144 3904 2208
rect 3968 2144 3976 2208
rect 3656 1120 3976 2144
rect 3656 1056 3664 1120
rect 3728 1056 3744 1120
rect 3808 1056 3824 1120
rect 3888 1056 3904 1120
rect 3968 1056 3976 1120
rect 3656 496 3976 1056
rect 4316 15808 4636 16832
rect 4846 16421 4906 19483
rect 4843 16420 4909 16421
rect 4843 16356 4844 16420
rect 4908 16356 4909 16420
rect 4843 16355 4909 16356
rect 4316 15744 4324 15808
rect 4388 15744 4404 15808
rect 4468 15744 4484 15808
rect 4548 15744 4564 15808
rect 4628 15744 4636 15808
rect 4316 14720 4636 15744
rect 4316 14656 4324 14720
rect 4388 14656 4404 14720
rect 4468 14656 4484 14720
rect 4548 14656 4564 14720
rect 4628 14656 4636 14720
rect 4316 13632 4636 14656
rect 5030 14517 5090 22203
rect 5214 21045 5274 28867
rect 5398 28797 5458 32403
rect 5582 30429 5642 35939
rect 5766 35869 5826 40019
rect 5763 35868 5829 35869
rect 5763 35804 5764 35868
rect 5828 35804 5829 35868
rect 5763 35803 5829 35804
rect 5950 34370 6010 40155
rect 6315 38316 6381 38317
rect 6315 38252 6316 38316
rect 6380 38252 6381 38316
rect 6315 38251 6381 38252
rect 5766 34310 6010 34370
rect 6318 34370 6378 38251
rect 6502 34506 6562 41515
rect 7051 41308 7117 41309
rect 7051 41244 7052 41308
rect 7116 41244 7117 41308
rect 7051 41243 7117 41244
rect 6867 38588 6933 38589
rect 6867 38524 6868 38588
rect 6932 38524 6933 38588
rect 6867 38523 6933 38524
rect 6870 37909 6930 38523
rect 6867 37908 6933 37909
rect 6867 37844 6868 37908
rect 6932 37844 6933 37908
rect 6867 37843 6933 37844
rect 6870 35325 6930 37843
rect 7054 36549 7114 41243
rect 7419 40492 7485 40493
rect 7419 40428 7420 40492
rect 7484 40428 7485 40492
rect 7419 40427 7485 40428
rect 7235 38860 7301 38861
rect 7235 38796 7236 38860
rect 7300 38796 7301 38860
rect 7235 38795 7301 38796
rect 7051 36548 7117 36549
rect 7051 36484 7052 36548
rect 7116 36484 7117 36548
rect 7051 36483 7117 36484
rect 6867 35324 6933 35325
rect 6867 35260 6868 35324
rect 6932 35260 6933 35324
rect 6867 35259 6933 35260
rect 6502 34446 7114 34506
rect 6867 34372 6933 34373
rect 6318 34310 6746 34370
rect 5766 33557 5826 34310
rect 5763 33556 5829 33557
rect 5763 33492 5764 33556
rect 5828 33492 5829 33556
rect 5763 33491 5829 33492
rect 5947 33420 6013 33421
rect 5947 33356 5948 33420
rect 6012 33356 6013 33420
rect 5947 33355 6013 33356
rect 5763 31788 5829 31789
rect 5763 31724 5764 31788
rect 5828 31724 5829 31788
rect 5763 31723 5829 31724
rect 5766 30837 5826 31723
rect 5950 31653 6010 33355
rect 6499 32604 6565 32605
rect 6499 32540 6500 32604
rect 6564 32540 6565 32604
rect 6499 32539 6565 32540
rect 6131 32468 6197 32469
rect 6131 32404 6132 32468
rect 6196 32404 6197 32468
rect 6131 32403 6197 32404
rect 5947 31652 6013 31653
rect 5947 31588 5948 31652
rect 6012 31588 6013 31652
rect 5947 31587 6013 31588
rect 5763 30836 5829 30837
rect 5763 30772 5764 30836
rect 5828 30772 5829 30836
rect 5763 30771 5829 30772
rect 5579 30428 5645 30429
rect 5579 30364 5580 30428
rect 5644 30364 5645 30428
rect 5579 30363 5645 30364
rect 5395 28796 5461 28797
rect 5395 28732 5396 28796
rect 5460 28732 5461 28796
rect 5395 28731 5461 28732
rect 5579 28796 5645 28797
rect 5579 28732 5580 28796
rect 5644 28732 5645 28796
rect 5579 28731 5645 28732
rect 5395 26892 5461 26893
rect 5395 26828 5396 26892
rect 5460 26828 5461 26892
rect 5395 26827 5461 26828
rect 5398 23490 5458 26827
rect 5582 25397 5642 28731
rect 5579 25396 5645 25397
rect 5579 25332 5580 25396
rect 5644 25332 5645 25396
rect 5579 25331 5645 25332
rect 5766 24989 5826 30771
rect 5947 30156 6013 30157
rect 5947 30092 5948 30156
rect 6012 30092 6013 30156
rect 5947 30091 6013 30092
rect 5763 24988 5829 24989
rect 5763 24924 5764 24988
rect 5828 24924 5829 24988
rect 5763 24923 5829 24924
rect 5763 24580 5829 24581
rect 5763 24516 5764 24580
rect 5828 24516 5829 24580
rect 5763 24515 5829 24516
rect 5398 23430 5642 23490
rect 5395 21452 5461 21453
rect 5395 21388 5396 21452
rect 5460 21388 5461 21452
rect 5395 21387 5461 21388
rect 5211 21044 5277 21045
rect 5211 20980 5212 21044
rect 5276 20980 5277 21044
rect 5211 20979 5277 20980
rect 5211 20772 5277 20773
rect 5211 20708 5212 20772
rect 5276 20708 5277 20772
rect 5211 20707 5277 20708
rect 5214 19957 5274 20707
rect 5211 19956 5277 19957
rect 5211 19892 5212 19956
rect 5276 19892 5277 19956
rect 5211 19891 5277 19892
rect 5398 19005 5458 21387
rect 5582 20773 5642 23430
rect 5579 20772 5645 20773
rect 5579 20708 5580 20772
rect 5644 20708 5645 20772
rect 5579 20707 5645 20708
rect 5579 20636 5645 20637
rect 5579 20572 5580 20636
rect 5644 20572 5645 20636
rect 5579 20571 5645 20572
rect 5582 19685 5642 20571
rect 5579 19684 5645 19685
rect 5579 19620 5580 19684
rect 5644 19620 5645 19684
rect 5579 19619 5645 19620
rect 5579 19412 5645 19413
rect 5579 19348 5580 19412
rect 5644 19348 5645 19412
rect 5579 19347 5645 19348
rect 5395 19004 5461 19005
rect 5395 18940 5396 19004
rect 5460 18940 5461 19004
rect 5395 18939 5461 18940
rect 5395 18052 5461 18053
rect 5395 17988 5396 18052
rect 5460 17988 5461 18052
rect 5395 17987 5461 17988
rect 5027 14516 5093 14517
rect 5027 14452 5028 14516
rect 5092 14452 5093 14516
rect 5027 14451 5093 14452
rect 4316 13568 4324 13632
rect 4388 13568 4404 13632
rect 4468 13568 4484 13632
rect 4548 13568 4564 13632
rect 4628 13568 4636 13632
rect 4316 12544 4636 13568
rect 4316 12480 4324 12544
rect 4388 12480 4404 12544
rect 4468 12480 4484 12544
rect 4548 12480 4564 12544
rect 4628 12480 4636 12544
rect 4316 11456 4636 12480
rect 5211 12476 5277 12477
rect 5211 12412 5212 12476
rect 5276 12412 5277 12476
rect 5211 12411 5277 12412
rect 5214 12341 5274 12411
rect 5211 12340 5277 12341
rect 5211 12276 5212 12340
rect 5276 12276 5277 12340
rect 5211 12275 5277 12276
rect 4316 11392 4324 11456
rect 4388 11392 4404 11456
rect 4468 11392 4484 11456
rect 4548 11392 4564 11456
rect 4628 11392 4636 11456
rect 4316 10368 4636 11392
rect 4316 10304 4324 10368
rect 4388 10304 4404 10368
rect 4468 10304 4484 10368
rect 4548 10304 4564 10368
rect 4628 10304 4636 10368
rect 4316 9280 4636 10304
rect 5398 10029 5458 17987
rect 5395 10028 5461 10029
rect 5395 9964 5396 10028
rect 5460 9964 5461 10028
rect 5395 9963 5461 9964
rect 4316 9216 4324 9280
rect 4388 9216 4404 9280
rect 4468 9216 4484 9280
rect 4548 9216 4564 9280
rect 4628 9216 4636 9280
rect 4316 8192 4636 9216
rect 5582 8669 5642 19347
rect 5766 17373 5826 24515
rect 5950 21861 6010 30091
rect 6134 27709 6194 32403
rect 6315 31788 6381 31789
rect 6315 31724 6316 31788
rect 6380 31724 6381 31788
rect 6315 31723 6381 31724
rect 6318 30157 6378 31723
rect 6315 30156 6381 30157
rect 6315 30092 6316 30156
rect 6380 30092 6381 30156
rect 6315 30091 6381 30092
rect 6131 27708 6197 27709
rect 6131 27644 6132 27708
rect 6196 27644 6197 27708
rect 6131 27643 6197 27644
rect 6318 27570 6378 30091
rect 6502 29202 6562 32539
rect 6686 30021 6746 34310
rect 6867 34308 6868 34372
rect 6932 34308 6933 34372
rect 6867 34307 6933 34308
rect 6870 33965 6930 34307
rect 6867 33964 6933 33965
rect 6867 33900 6868 33964
rect 6932 33900 6933 33964
rect 6867 33899 6933 33900
rect 6870 32741 6930 33899
rect 6867 32740 6933 32741
rect 6867 32676 6868 32740
rect 6932 32676 6933 32740
rect 6867 32675 6933 32676
rect 6867 32332 6933 32333
rect 6867 32268 6868 32332
rect 6932 32268 6933 32332
rect 6867 32267 6933 32268
rect 6870 30429 6930 32267
rect 7054 31925 7114 34446
rect 7238 32605 7298 38795
rect 7235 32604 7301 32605
rect 7235 32540 7236 32604
rect 7300 32540 7301 32604
rect 7235 32539 7301 32540
rect 7051 31924 7117 31925
rect 7051 31860 7052 31924
rect 7116 31860 7117 31924
rect 7051 31859 7117 31860
rect 6867 30428 6933 30429
rect 6867 30364 6868 30428
rect 6932 30364 6933 30428
rect 6867 30363 6933 30364
rect 6683 30020 6749 30021
rect 6683 29956 6684 30020
rect 6748 29956 6749 30020
rect 6683 29955 6749 29956
rect 6502 29142 6746 29202
rect 6499 29068 6565 29069
rect 6499 29004 6500 29068
rect 6564 29004 6565 29068
rect 6499 29003 6565 29004
rect 6134 27510 6378 27570
rect 5947 21860 6013 21861
rect 5947 21796 5948 21860
rect 6012 21796 6013 21860
rect 5947 21795 6013 21796
rect 5947 19276 6013 19277
rect 5947 19212 5948 19276
rect 6012 19212 6013 19276
rect 5947 19211 6013 19212
rect 5763 17372 5829 17373
rect 5763 17308 5764 17372
rect 5828 17308 5829 17372
rect 5763 17307 5829 17308
rect 5766 13837 5826 17307
rect 5763 13836 5829 13837
rect 5763 13772 5764 13836
rect 5828 13772 5829 13836
rect 5763 13771 5829 13772
rect 5950 12885 6010 19211
rect 6134 17917 6194 27510
rect 6315 26076 6381 26077
rect 6315 26012 6316 26076
rect 6380 26012 6381 26076
rect 6315 26011 6381 26012
rect 6131 17916 6197 17917
rect 6131 17852 6132 17916
rect 6196 17852 6197 17916
rect 6131 17851 6197 17852
rect 6318 14517 6378 26011
rect 6502 19277 6562 29003
rect 6686 28117 6746 29142
rect 6870 28930 6930 30363
rect 7054 29205 7114 31859
rect 7422 31653 7482 40427
rect 7787 39540 7853 39541
rect 7787 39476 7788 39540
rect 7852 39476 7853 39540
rect 7787 39475 7853 39476
rect 7603 38452 7669 38453
rect 7603 38388 7604 38452
rect 7668 38388 7669 38452
rect 7603 38387 7669 38388
rect 7606 37093 7666 38387
rect 7603 37092 7669 37093
rect 7603 37028 7604 37092
rect 7668 37028 7669 37092
rect 7603 37027 7669 37028
rect 7606 35597 7666 37027
rect 7790 36141 7850 39475
rect 7971 37364 8037 37365
rect 7971 37300 7972 37364
rect 8036 37300 8037 37364
rect 7971 37299 8037 37300
rect 7787 36140 7853 36141
rect 7787 36076 7788 36140
rect 7852 36076 7853 36140
rect 7787 36075 7853 36076
rect 7603 35596 7669 35597
rect 7603 35532 7604 35596
rect 7668 35532 7669 35596
rect 7603 35531 7669 35532
rect 7787 33284 7853 33285
rect 7787 33220 7788 33284
rect 7852 33220 7853 33284
rect 7787 33219 7853 33220
rect 7603 32196 7669 32197
rect 7603 32132 7604 32196
rect 7668 32132 7669 32196
rect 7603 32131 7669 32132
rect 7419 31652 7485 31653
rect 7419 31588 7420 31652
rect 7484 31588 7485 31652
rect 7419 31587 7485 31588
rect 7422 30701 7482 31587
rect 7419 30700 7485 30701
rect 7419 30636 7420 30700
rect 7484 30636 7485 30700
rect 7419 30635 7485 30636
rect 7606 30429 7666 32131
rect 7603 30428 7669 30429
rect 7603 30364 7604 30428
rect 7668 30364 7669 30428
rect 7603 30363 7669 30364
rect 7790 30157 7850 33219
rect 7974 32061 8034 37299
rect 7971 32060 8037 32061
rect 7971 31996 7972 32060
rect 8036 31996 8037 32060
rect 7971 31995 8037 31996
rect 8158 30293 8218 43555
rect 8707 41988 8773 41989
rect 8707 41924 8708 41988
rect 8772 41924 8773 41988
rect 8707 41923 8773 41924
rect 8523 41036 8589 41037
rect 8523 40972 8524 41036
rect 8588 40972 8589 41036
rect 8523 40971 8589 40972
rect 8339 37908 8405 37909
rect 8339 37844 8340 37908
rect 8404 37844 8405 37908
rect 8339 37843 8405 37844
rect 8342 33693 8402 37843
rect 8339 33692 8405 33693
rect 8339 33628 8340 33692
rect 8404 33628 8405 33692
rect 8339 33627 8405 33628
rect 8339 32740 8405 32741
rect 8339 32676 8340 32740
rect 8404 32676 8405 32740
rect 8339 32675 8405 32676
rect 8155 30292 8221 30293
rect 8155 30228 8156 30292
rect 8220 30228 8221 30292
rect 8155 30227 8221 30228
rect 7787 30156 7853 30157
rect 7787 30092 7788 30156
rect 7852 30092 7853 30156
rect 7787 30091 7853 30092
rect 7051 29204 7117 29205
rect 7051 29140 7052 29204
rect 7116 29140 7117 29204
rect 7051 29139 7117 29140
rect 7419 28932 7485 28933
rect 6870 28870 7114 28930
rect 7054 28389 7114 28870
rect 7419 28868 7420 28932
rect 7484 28868 7485 28932
rect 7419 28867 7485 28868
rect 7971 28932 8037 28933
rect 7971 28868 7972 28932
rect 8036 28868 8037 28932
rect 7971 28867 8037 28868
rect 7051 28388 7117 28389
rect 7051 28324 7052 28388
rect 7116 28324 7117 28388
rect 7051 28323 7117 28324
rect 6683 28116 6749 28117
rect 6683 28052 6684 28116
rect 6748 28052 6749 28116
rect 6683 28051 6749 28052
rect 6867 28116 6933 28117
rect 6867 28052 6868 28116
rect 6932 28052 6933 28116
rect 6867 28051 6933 28052
rect 6683 27436 6749 27437
rect 6683 27372 6684 27436
rect 6748 27372 6749 27436
rect 6683 27371 6749 27372
rect 6686 23626 6746 27371
rect 6870 23765 6930 28051
rect 7054 26485 7114 28323
rect 7051 26484 7117 26485
rect 7051 26420 7052 26484
rect 7116 26420 7117 26484
rect 7051 26419 7117 26420
rect 7051 25668 7117 25669
rect 7051 25604 7052 25668
rect 7116 25604 7117 25668
rect 7051 25603 7117 25604
rect 6867 23764 6933 23765
rect 6867 23700 6868 23764
rect 6932 23700 6933 23764
rect 6867 23699 6933 23700
rect 6686 23566 6930 23626
rect 6683 23492 6749 23493
rect 6683 23428 6684 23492
rect 6748 23428 6749 23492
rect 6683 23427 6749 23428
rect 6499 19276 6565 19277
rect 6499 19212 6500 19276
rect 6564 19212 6565 19276
rect 6499 19211 6565 19212
rect 6686 18189 6746 23427
rect 6870 21997 6930 23566
rect 6867 21996 6933 21997
rect 6867 21932 6868 21996
rect 6932 21932 6933 21996
rect 6867 21931 6933 21932
rect 6683 18188 6749 18189
rect 6683 18124 6684 18188
rect 6748 18124 6749 18188
rect 6683 18123 6749 18124
rect 7054 17781 7114 25603
rect 7422 23765 7482 28867
rect 7787 28116 7853 28117
rect 7787 28052 7788 28116
rect 7852 28052 7853 28116
rect 7787 28051 7853 28052
rect 7603 27572 7669 27573
rect 7603 27508 7604 27572
rect 7668 27508 7669 27572
rect 7603 27507 7669 27508
rect 7419 23764 7485 23765
rect 7419 23700 7420 23764
rect 7484 23700 7485 23764
rect 7419 23699 7485 23700
rect 7422 22269 7482 23699
rect 7419 22268 7485 22269
rect 7419 22204 7420 22268
rect 7484 22204 7485 22268
rect 7419 22203 7485 22204
rect 7606 19413 7666 27507
rect 7790 20909 7850 28051
rect 7974 23357 8034 28867
rect 8155 27980 8221 27981
rect 8155 27916 8156 27980
rect 8220 27916 8221 27980
rect 8155 27915 8221 27916
rect 8158 26349 8218 27915
rect 8342 27845 8402 32675
rect 8526 30429 8586 40971
rect 8710 31789 8770 41923
rect 8891 40084 8957 40085
rect 8891 40020 8892 40084
rect 8956 40020 8957 40084
rect 8891 40019 8957 40020
rect 8707 31788 8773 31789
rect 8707 31724 8708 31788
rect 8772 31724 8773 31788
rect 8707 31723 8773 31724
rect 8707 31108 8773 31109
rect 8707 31044 8708 31108
rect 8772 31044 8773 31108
rect 8707 31043 8773 31044
rect 8523 30428 8589 30429
rect 8523 30364 8524 30428
rect 8588 30364 8589 30428
rect 8523 30363 8589 30364
rect 8523 27980 8589 27981
rect 8523 27916 8524 27980
rect 8588 27916 8589 27980
rect 8523 27915 8589 27916
rect 8339 27844 8405 27845
rect 8339 27780 8340 27844
rect 8404 27780 8405 27844
rect 8339 27779 8405 27780
rect 8526 26890 8586 27915
rect 8342 26830 8586 26890
rect 8155 26348 8221 26349
rect 8155 26284 8156 26348
rect 8220 26284 8221 26348
rect 8155 26283 8221 26284
rect 8342 26210 8402 26830
rect 8158 26150 8402 26210
rect 7971 23356 8037 23357
rect 7971 23292 7972 23356
rect 8036 23292 8037 23356
rect 7971 23291 8037 23292
rect 7971 23084 8037 23085
rect 7971 23020 7972 23084
rect 8036 23020 8037 23084
rect 7971 23019 8037 23020
rect 7974 21861 8034 23019
rect 7971 21860 8037 21861
rect 7971 21796 7972 21860
rect 8036 21796 8037 21860
rect 7971 21795 8037 21796
rect 7787 20908 7853 20909
rect 7787 20844 7788 20908
rect 7852 20844 7853 20908
rect 7787 20843 7853 20844
rect 7787 20772 7853 20773
rect 7787 20708 7788 20772
rect 7852 20708 7853 20772
rect 7787 20707 7853 20708
rect 7603 19412 7669 19413
rect 7603 19348 7604 19412
rect 7668 19348 7669 19412
rect 7603 19347 7669 19348
rect 7790 17917 7850 20707
rect 7974 19005 8034 21795
rect 8158 20093 8218 26150
rect 8339 21996 8405 21997
rect 8339 21932 8340 21996
rect 8404 21932 8405 21996
rect 8339 21931 8405 21932
rect 8155 20092 8221 20093
rect 8155 20028 8156 20092
rect 8220 20028 8221 20092
rect 8155 20027 8221 20028
rect 7971 19004 8037 19005
rect 7971 18940 7972 19004
rect 8036 18940 8037 19004
rect 7971 18939 8037 18940
rect 7787 17916 7853 17917
rect 7787 17852 7788 17916
rect 7852 17852 7853 17916
rect 7787 17851 7853 17852
rect 7051 17780 7117 17781
rect 7051 17716 7052 17780
rect 7116 17716 7117 17780
rect 7051 17715 7117 17716
rect 7419 17644 7485 17645
rect 7419 17580 7420 17644
rect 7484 17580 7485 17644
rect 7419 17579 7485 17580
rect 6683 17236 6749 17237
rect 6683 17172 6684 17236
rect 6748 17172 6749 17236
rect 6683 17171 6749 17172
rect 6686 16965 6746 17171
rect 6683 16964 6749 16965
rect 6683 16900 6684 16964
rect 6748 16900 6749 16964
rect 6683 16899 6749 16900
rect 6315 14516 6381 14517
rect 6315 14452 6316 14516
rect 6380 14452 6381 14516
rect 6315 14451 6381 14452
rect 5947 12884 6013 12885
rect 5947 12820 5948 12884
rect 6012 12820 6013 12884
rect 5947 12819 6013 12820
rect 5579 8668 5645 8669
rect 5579 8604 5580 8668
rect 5644 8604 5645 8668
rect 5579 8603 5645 8604
rect 7422 8261 7482 17579
rect 8342 16590 8402 21931
rect 8710 20090 8770 31043
rect 8894 28661 8954 40019
rect 9075 37636 9141 37637
rect 9075 37572 9076 37636
rect 9140 37572 9141 37636
rect 9075 37571 9141 37572
rect 9078 31109 9138 37571
rect 9262 33829 9322 43555
rect 9443 38724 9509 38725
rect 9443 38660 9444 38724
rect 9508 38660 9509 38724
rect 9443 38659 9509 38660
rect 9446 35325 9506 38659
rect 9443 35324 9509 35325
rect 9443 35260 9444 35324
rect 9508 35260 9509 35324
rect 9443 35259 9509 35260
rect 9259 33828 9325 33829
rect 9259 33764 9260 33828
rect 9324 33764 9325 33828
rect 9259 33763 9325 33764
rect 9259 33692 9325 33693
rect 9259 33628 9260 33692
rect 9324 33628 9325 33692
rect 9259 33627 9325 33628
rect 9075 31108 9141 31109
rect 9075 31044 9076 31108
rect 9140 31044 9141 31108
rect 9075 31043 9141 31044
rect 9262 30973 9322 33627
rect 9443 32740 9509 32741
rect 9443 32676 9444 32740
rect 9508 32676 9509 32740
rect 9443 32675 9509 32676
rect 9259 30972 9325 30973
rect 9259 30908 9260 30972
rect 9324 30908 9325 30972
rect 9259 30907 9325 30908
rect 9075 30700 9141 30701
rect 9075 30636 9076 30700
rect 9140 30636 9141 30700
rect 9075 30635 9141 30636
rect 8891 28660 8957 28661
rect 8891 28596 8892 28660
rect 8956 28596 8957 28660
rect 8891 28595 8957 28596
rect 9078 28525 9138 30635
rect 9262 30565 9322 30907
rect 9259 30564 9325 30565
rect 9259 30500 9260 30564
rect 9324 30500 9325 30564
rect 9259 30499 9325 30500
rect 9075 28524 9141 28525
rect 9075 28460 9076 28524
rect 9140 28460 9141 28524
rect 9075 28459 9141 28460
rect 8891 27572 8957 27573
rect 8891 27508 8892 27572
rect 8956 27508 8957 27572
rect 8891 27507 8957 27508
rect 8526 20030 8770 20090
rect 8526 17509 8586 20030
rect 8707 19412 8773 19413
rect 8707 19348 8708 19412
rect 8772 19348 8773 19412
rect 8707 19347 8773 19348
rect 8710 17781 8770 19347
rect 8894 17917 8954 27507
rect 9446 26077 9506 32675
rect 9630 27165 9690 43555
rect 10056 42464 10376 43024
rect 10056 42400 10064 42464
rect 10128 42400 10144 42464
rect 10208 42400 10224 42464
rect 10288 42400 10304 42464
rect 10368 42400 10376 42464
rect 9811 41716 9877 41717
rect 9811 41652 9812 41716
rect 9876 41652 9877 41716
rect 9811 41651 9877 41652
rect 9814 38861 9874 41651
rect 10056 41376 10376 42400
rect 10056 41312 10064 41376
rect 10128 41312 10144 41376
rect 10208 41312 10224 41376
rect 10288 41312 10304 41376
rect 10368 41312 10376 41376
rect 10056 40288 10376 41312
rect 10056 40224 10064 40288
rect 10128 40224 10144 40288
rect 10208 40224 10224 40288
rect 10288 40224 10304 40288
rect 10368 40224 10376 40288
rect 10056 39200 10376 40224
rect 10716 43008 11036 43024
rect 10716 42944 10724 43008
rect 10788 42944 10804 43008
rect 10868 42944 10884 43008
rect 10948 42944 10964 43008
rect 11028 42944 11036 43008
rect 10716 41920 11036 42944
rect 11467 41988 11533 41989
rect 11467 41924 11468 41988
rect 11532 41924 11533 41988
rect 11467 41923 11533 41924
rect 10716 41856 10724 41920
rect 10788 41856 10804 41920
rect 10868 41856 10884 41920
rect 10948 41856 10964 41920
rect 11028 41856 11036 41920
rect 10716 40832 11036 41856
rect 10716 40768 10724 40832
rect 10788 40768 10804 40832
rect 10868 40768 10884 40832
rect 10948 40768 10964 40832
rect 11028 40768 11036 40832
rect 10547 40220 10613 40221
rect 10547 40156 10548 40220
rect 10612 40156 10613 40220
rect 10547 40155 10613 40156
rect 10056 39136 10064 39200
rect 10128 39136 10144 39200
rect 10208 39136 10224 39200
rect 10288 39136 10304 39200
rect 10368 39136 10376 39200
rect 9811 38860 9877 38861
rect 9811 38796 9812 38860
rect 9876 38796 9877 38860
rect 9811 38795 9877 38796
rect 10056 38112 10376 39136
rect 10550 38317 10610 40155
rect 10716 39744 11036 40768
rect 11283 40084 11349 40085
rect 11283 40020 11284 40084
rect 11348 40020 11349 40084
rect 11283 40019 11349 40020
rect 10716 39680 10724 39744
rect 10788 39680 10804 39744
rect 10868 39680 10884 39744
rect 10948 39680 10964 39744
rect 11028 39680 11036 39744
rect 10716 38656 11036 39680
rect 10716 38592 10724 38656
rect 10788 38592 10804 38656
rect 10868 38592 10884 38656
rect 10948 38592 10964 38656
rect 11028 38592 11036 38656
rect 10547 38316 10613 38317
rect 10547 38252 10548 38316
rect 10612 38252 10613 38316
rect 10547 38251 10613 38252
rect 10056 38048 10064 38112
rect 10128 38048 10144 38112
rect 10208 38048 10224 38112
rect 10288 38048 10304 38112
rect 10368 38048 10376 38112
rect 9811 37908 9877 37909
rect 9811 37844 9812 37908
rect 9876 37844 9877 37908
rect 9811 37843 9877 37844
rect 9814 37229 9874 37843
rect 9811 37228 9877 37229
rect 9811 37164 9812 37228
rect 9876 37164 9877 37228
rect 9811 37163 9877 37164
rect 9814 35597 9874 37163
rect 10056 37024 10376 38048
rect 10716 37568 11036 38592
rect 11099 38316 11165 38317
rect 11099 38252 11100 38316
rect 11164 38252 11165 38316
rect 11099 38251 11165 38252
rect 10716 37504 10724 37568
rect 10788 37504 10804 37568
rect 10868 37504 10884 37568
rect 10948 37504 10964 37568
rect 11028 37504 11036 37568
rect 10547 37364 10613 37365
rect 10547 37300 10548 37364
rect 10612 37300 10613 37364
rect 10547 37299 10613 37300
rect 10056 36960 10064 37024
rect 10128 36960 10144 37024
rect 10208 36960 10224 37024
rect 10288 36960 10304 37024
rect 10368 36960 10376 37024
rect 10056 35936 10376 36960
rect 10056 35872 10064 35936
rect 10128 35872 10144 35936
rect 10208 35872 10224 35936
rect 10288 35872 10304 35936
rect 10368 35872 10376 35936
rect 9811 35596 9877 35597
rect 9811 35532 9812 35596
rect 9876 35532 9877 35596
rect 9811 35531 9877 35532
rect 9811 35324 9877 35325
rect 9811 35260 9812 35324
rect 9876 35260 9877 35324
rect 9811 35259 9877 35260
rect 9814 30293 9874 35259
rect 10056 34848 10376 35872
rect 10056 34784 10064 34848
rect 10128 34784 10144 34848
rect 10208 34784 10224 34848
rect 10288 34784 10304 34848
rect 10368 34784 10376 34848
rect 10056 33760 10376 34784
rect 10056 33696 10064 33760
rect 10128 33696 10144 33760
rect 10208 33696 10224 33760
rect 10288 33696 10304 33760
rect 10368 33696 10376 33760
rect 10056 32672 10376 33696
rect 10056 32608 10064 32672
rect 10128 32608 10144 32672
rect 10208 32608 10224 32672
rect 10288 32608 10304 32672
rect 10368 32608 10376 32672
rect 10056 31584 10376 32608
rect 10550 32197 10610 37299
rect 10716 36480 11036 37504
rect 11102 36957 11162 38251
rect 11099 36956 11165 36957
rect 11099 36892 11100 36956
rect 11164 36892 11165 36956
rect 11099 36891 11165 36892
rect 11099 36820 11165 36821
rect 11099 36756 11100 36820
rect 11164 36756 11165 36820
rect 11099 36755 11165 36756
rect 10716 36416 10724 36480
rect 10788 36416 10804 36480
rect 10868 36416 10884 36480
rect 10948 36416 10964 36480
rect 11028 36416 11036 36480
rect 10716 35392 11036 36416
rect 10716 35328 10724 35392
rect 10788 35328 10804 35392
rect 10868 35328 10884 35392
rect 10948 35328 10964 35392
rect 11028 35328 11036 35392
rect 10716 34304 11036 35328
rect 11102 35053 11162 36755
rect 11099 35052 11165 35053
rect 11099 34988 11100 35052
rect 11164 34988 11165 35052
rect 11099 34987 11165 34988
rect 10716 34240 10724 34304
rect 10788 34240 10804 34304
rect 10868 34240 10884 34304
rect 10948 34240 10964 34304
rect 11028 34240 11036 34304
rect 10716 33216 11036 34240
rect 10716 33152 10724 33216
rect 10788 33152 10804 33216
rect 10868 33152 10884 33216
rect 10948 33152 10964 33216
rect 11028 33152 11036 33216
rect 10547 32196 10613 32197
rect 10547 32132 10548 32196
rect 10612 32132 10613 32196
rect 10547 32131 10613 32132
rect 10716 32128 11036 33152
rect 10716 32064 10724 32128
rect 10788 32064 10804 32128
rect 10868 32064 10884 32128
rect 10948 32064 10964 32128
rect 11028 32064 11036 32128
rect 10547 31924 10613 31925
rect 10547 31860 10548 31924
rect 10612 31860 10613 31924
rect 10547 31859 10613 31860
rect 10056 31520 10064 31584
rect 10128 31520 10144 31584
rect 10208 31520 10224 31584
rect 10288 31520 10304 31584
rect 10368 31520 10376 31584
rect 10056 30496 10376 31520
rect 10056 30432 10064 30496
rect 10128 30432 10144 30496
rect 10208 30432 10224 30496
rect 10288 30432 10304 30496
rect 10368 30432 10376 30496
rect 9811 30292 9877 30293
rect 9811 30228 9812 30292
rect 9876 30228 9877 30292
rect 9811 30227 9877 30228
rect 10056 29408 10376 30432
rect 10550 29477 10610 31859
rect 10716 31040 11036 32064
rect 11102 31925 11162 34987
rect 11099 31924 11165 31925
rect 11099 31860 11100 31924
rect 11164 31860 11165 31924
rect 11099 31859 11165 31860
rect 11099 31652 11165 31653
rect 11099 31588 11100 31652
rect 11164 31588 11165 31652
rect 11099 31587 11165 31588
rect 10716 30976 10724 31040
rect 10788 30976 10804 31040
rect 10868 30976 10884 31040
rect 10948 30976 10964 31040
rect 11028 30976 11036 31040
rect 10716 29952 11036 30976
rect 10716 29888 10724 29952
rect 10788 29888 10804 29952
rect 10868 29888 10884 29952
rect 10948 29888 10964 29952
rect 11028 29888 11036 29952
rect 10547 29476 10613 29477
rect 10547 29412 10548 29476
rect 10612 29412 10613 29476
rect 10547 29411 10613 29412
rect 10056 29344 10064 29408
rect 10128 29344 10144 29408
rect 10208 29344 10224 29408
rect 10288 29344 10304 29408
rect 10368 29344 10376 29408
rect 10056 28320 10376 29344
rect 10056 28256 10064 28320
rect 10128 28256 10144 28320
rect 10208 28256 10224 28320
rect 10288 28256 10304 28320
rect 10368 28256 10376 28320
rect 10056 27232 10376 28256
rect 10716 28864 11036 29888
rect 10716 28800 10724 28864
rect 10788 28800 10804 28864
rect 10868 28800 10884 28864
rect 10948 28800 10964 28864
rect 11028 28800 11036 28864
rect 10716 27776 11036 28800
rect 11102 27981 11162 31587
rect 11286 29341 11346 40019
rect 11470 30293 11530 41923
rect 11651 41580 11717 41581
rect 11651 41516 11652 41580
rect 11716 41516 11717 41580
rect 11651 41515 11717 41516
rect 11654 30429 11714 41515
rect 12019 38860 12085 38861
rect 12019 38796 12020 38860
rect 12084 38796 12085 38860
rect 12019 38795 12085 38796
rect 11835 37364 11901 37365
rect 11835 37300 11836 37364
rect 11900 37300 11901 37364
rect 11835 37299 11901 37300
rect 11838 33693 11898 37299
rect 11835 33692 11901 33693
rect 11835 33628 11836 33692
rect 11900 33628 11901 33692
rect 11835 33627 11901 33628
rect 11835 33556 11901 33557
rect 11835 33492 11836 33556
rect 11900 33492 11901 33556
rect 11835 33491 11901 33492
rect 11651 30428 11717 30429
rect 11651 30364 11652 30428
rect 11716 30364 11717 30428
rect 11651 30363 11717 30364
rect 11467 30292 11533 30293
rect 11467 30228 11468 30292
rect 11532 30228 11533 30292
rect 11467 30227 11533 30228
rect 11283 29340 11349 29341
rect 11283 29276 11284 29340
rect 11348 29276 11349 29340
rect 11283 29275 11349 29276
rect 11283 28524 11349 28525
rect 11283 28460 11284 28524
rect 11348 28460 11349 28524
rect 11283 28459 11349 28460
rect 11099 27980 11165 27981
rect 11099 27916 11100 27980
rect 11164 27916 11165 27980
rect 11099 27915 11165 27916
rect 10716 27712 10724 27776
rect 10788 27712 10804 27776
rect 10868 27712 10884 27776
rect 10948 27712 10964 27776
rect 11028 27712 11036 27776
rect 10547 27436 10613 27437
rect 10547 27372 10548 27436
rect 10612 27372 10613 27436
rect 10547 27371 10613 27372
rect 10056 27168 10064 27232
rect 10128 27168 10144 27232
rect 10208 27168 10224 27232
rect 10288 27168 10304 27232
rect 10368 27168 10376 27232
rect 9627 27164 9693 27165
rect 9627 27100 9628 27164
rect 9692 27100 9693 27164
rect 9627 27099 9693 27100
rect 9627 26484 9693 26485
rect 9627 26420 9628 26484
rect 9692 26420 9693 26484
rect 9627 26419 9693 26420
rect 9443 26076 9509 26077
rect 9443 26012 9444 26076
rect 9508 26012 9509 26076
rect 9443 26011 9509 26012
rect 9259 24716 9325 24717
rect 9259 24652 9260 24716
rect 9324 24652 9325 24716
rect 9259 24651 9325 24652
rect 9075 24580 9141 24581
rect 9075 24516 9076 24580
rect 9140 24516 9141 24580
rect 9075 24515 9141 24516
rect 9078 20501 9138 24515
rect 9075 20500 9141 20501
rect 9075 20436 9076 20500
rect 9140 20436 9141 20500
rect 9075 20435 9141 20436
rect 8891 17916 8957 17917
rect 8891 17852 8892 17916
rect 8956 17852 8957 17916
rect 8891 17851 8957 17852
rect 9078 17781 9138 20435
rect 8707 17780 8773 17781
rect 8707 17716 8708 17780
rect 8772 17716 8773 17780
rect 9075 17780 9141 17781
rect 9075 17778 9076 17780
rect 8707 17715 8773 17716
rect 8894 17718 9076 17778
rect 8523 17508 8589 17509
rect 8523 17444 8524 17508
rect 8588 17444 8589 17508
rect 8523 17443 8589 17444
rect 7787 16556 7853 16557
rect 7787 16492 7788 16556
rect 7852 16492 7853 16556
rect 7787 16491 7853 16492
rect 8158 16530 8402 16590
rect 7790 13701 7850 16491
rect 7787 13700 7853 13701
rect 7787 13636 7788 13700
rect 7852 13636 7853 13700
rect 7787 13635 7853 13636
rect 8158 11117 8218 16530
rect 8894 12885 8954 17718
rect 9075 17716 9076 17718
rect 9140 17716 9141 17780
rect 9075 17715 9141 17716
rect 9075 16692 9141 16693
rect 9075 16628 9076 16692
rect 9140 16628 9141 16692
rect 9075 16627 9141 16628
rect 8891 12884 8957 12885
rect 8891 12820 8892 12884
rect 8956 12820 8957 12884
rect 8891 12819 8957 12820
rect 8155 11116 8221 11117
rect 8155 11052 8156 11116
rect 8220 11052 8221 11116
rect 8155 11051 8221 11052
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 4316 8128 4324 8192
rect 4388 8128 4404 8192
rect 4468 8128 4484 8192
rect 4548 8128 4564 8192
rect 4628 8128 4636 8192
rect 4316 7104 4636 8128
rect 9078 7445 9138 16627
rect 9262 16149 9322 24651
rect 9443 22676 9509 22677
rect 9443 22612 9444 22676
rect 9508 22612 9509 22676
rect 9443 22611 9509 22612
rect 9446 20093 9506 22611
rect 9630 20906 9690 26419
rect 9811 26348 9877 26349
rect 9811 26284 9812 26348
rect 9876 26284 9877 26348
rect 9811 26283 9877 26284
rect 9814 21997 9874 26283
rect 10056 26144 10376 27168
rect 10056 26080 10064 26144
rect 10128 26080 10144 26144
rect 10208 26080 10224 26144
rect 10288 26080 10304 26144
rect 10368 26080 10376 26144
rect 10056 25056 10376 26080
rect 10056 24992 10064 25056
rect 10128 24992 10144 25056
rect 10208 24992 10224 25056
rect 10288 24992 10304 25056
rect 10368 24992 10376 25056
rect 10056 23968 10376 24992
rect 10056 23904 10064 23968
rect 10128 23904 10144 23968
rect 10208 23904 10224 23968
rect 10288 23904 10304 23968
rect 10368 23904 10376 23968
rect 10056 22880 10376 23904
rect 10056 22816 10064 22880
rect 10128 22816 10144 22880
rect 10208 22816 10224 22880
rect 10288 22816 10304 22880
rect 10368 22816 10376 22880
rect 9811 21996 9877 21997
rect 9811 21932 9812 21996
rect 9876 21932 9877 21996
rect 9811 21931 9877 21932
rect 10056 21792 10376 22816
rect 10056 21728 10064 21792
rect 10128 21728 10144 21792
rect 10208 21728 10224 21792
rect 10288 21728 10304 21792
rect 10368 21728 10376 21792
rect 9630 20846 9874 20906
rect 9627 20772 9693 20773
rect 9627 20708 9628 20772
rect 9692 20708 9693 20772
rect 9627 20707 9693 20708
rect 9443 20092 9509 20093
rect 9443 20028 9444 20092
rect 9508 20028 9509 20092
rect 9443 20027 9509 20028
rect 9443 17916 9509 17917
rect 9443 17852 9444 17916
rect 9508 17852 9509 17916
rect 9443 17851 9509 17852
rect 9259 16148 9325 16149
rect 9259 16084 9260 16148
rect 9324 16084 9325 16148
rect 9259 16083 9325 16084
rect 9262 15333 9322 16083
rect 9259 15332 9325 15333
rect 9259 15268 9260 15332
rect 9324 15268 9325 15332
rect 9259 15267 9325 15268
rect 9446 8125 9506 17851
rect 9630 17237 9690 20707
rect 9627 17236 9693 17237
rect 9627 17172 9628 17236
rect 9692 17172 9693 17236
rect 9627 17171 9693 17172
rect 9814 16557 9874 20846
rect 10056 20704 10376 21728
rect 10550 21317 10610 27371
rect 10716 26688 11036 27712
rect 10716 26624 10724 26688
rect 10788 26624 10804 26688
rect 10868 26624 10884 26688
rect 10948 26624 10964 26688
rect 11028 26624 11036 26688
rect 10716 25600 11036 26624
rect 10716 25536 10724 25600
rect 10788 25536 10804 25600
rect 10868 25536 10884 25600
rect 10948 25536 10964 25600
rect 11028 25536 11036 25600
rect 10716 24512 11036 25536
rect 10716 24448 10724 24512
rect 10788 24448 10804 24512
rect 10868 24448 10884 24512
rect 10948 24448 10964 24512
rect 11028 24448 11036 24512
rect 10716 23424 11036 24448
rect 10716 23360 10724 23424
rect 10788 23360 10804 23424
rect 10868 23360 10884 23424
rect 10948 23360 10964 23424
rect 11028 23360 11036 23424
rect 10716 22336 11036 23360
rect 10716 22272 10724 22336
rect 10788 22272 10804 22336
rect 10868 22272 10884 22336
rect 10948 22272 10964 22336
rect 11028 22272 11036 22336
rect 10547 21316 10613 21317
rect 10547 21252 10548 21316
rect 10612 21252 10613 21316
rect 10547 21251 10613 21252
rect 10056 20640 10064 20704
rect 10128 20640 10144 20704
rect 10208 20640 10224 20704
rect 10288 20640 10304 20704
rect 10368 20640 10376 20704
rect 10056 19616 10376 20640
rect 10716 21248 11036 22272
rect 10716 21184 10724 21248
rect 10788 21184 10804 21248
rect 10868 21184 10884 21248
rect 10948 21184 10964 21248
rect 11028 21184 11036 21248
rect 10716 20160 11036 21184
rect 10716 20096 10724 20160
rect 10788 20096 10804 20160
rect 10868 20096 10884 20160
rect 10948 20096 10964 20160
rect 11028 20096 11036 20160
rect 10547 19684 10613 19685
rect 10547 19620 10548 19684
rect 10612 19620 10613 19684
rect 10547 19619 10613 19620
rect 10056 19552 10064 19616
rect 10128 19552 10144 19616
rect 10208 19552 10224 19616
rect 10288 19552 10304 19616
rect 10368 19552 10376 19616
rect 10056 18528 10376 19552
rect 10056 18464 10064 18528
rect 10128 18464 10144 18528
rect 10208 18464 10224 18528
rect 10288 18464 10304 18528
rect 10368 18464 10376 18528
rect 10056 17440 10376 18464
rect 10056 17376 10064 17440
rect 10128 17376 10144 17440
rect 10208 17376 10224 17440
rect 10288 17376 10304 17440
rect 10368 17376 10376 17440
rect 9811 16556 9877 16557
rect 9811 16492 9812 16556
rect 9876 16492 9877 16556
rect 9811 16491 9877 16492
rect 10056 16352 10376 17376
rect 10056 16288 10064 16352
rect 10128 16288 10144 16352
rect 10208 16288 10224 16352
rect 10288 16288 10304 16352
rect 10368 16288 10376 16352
rect 9811 16284 9877 16285
rect 9811 16220 9812 16284
rect 9876 16220 9877 16284
rect 9811 16219 9877 16220
rect 9814 10029 9874 16219
rect 10056 15264 10376 16288
rect 10056 15200 10064 15264
rect 10128 15200 10144 15264
rect 10208 15200 10224 15264
rect 10288 15200 10304 15264
rect 10368 15200 10376 15264
rect 10056 14176 10376 15200
rect 10056 14112 10064 14176
rect 10128 14112 10144 14176
rect 10208 14112 10224 14176
rect 10288 14112 10304 14176
rect 10368 14112 10376 14176
rect 10056 13088 10376 14112
rect 10056 13024 10064 13088
rect 10128 13024 10144 13088
rect 10208 13024 10224 13088
rect 10288 13024 10304 13088
rect 10368 13024 10376 13088
rect 10056 12000 10376 13024
rect 10550 12341 10610 19619
rect 10716 19072 11036 20096
rect 10716 19008 10724 19072
rect 10788 19008 10804 19072
rect 10868 19008 10884 19072
rect 10948 19008 10964 19072
rect 11028 19008 11036 19072
rect 10716 17984 11036 19008
rect 10716 17920 10724 17984
rect 10788 17920 10804 17984
rect 10868 17920 10884 17984
rect 10948 17920 10964 17984
rect 11028 17920 11036 17984
rect 10716 16896 11036 17920
rect 11286 17645 11346 28459
rect 11651 27708 11717 27709
rect 11651 27644 11652 27708
rect 11716 27644 11717 27708
rect 11651 27643 11717 27644
rect 11467 23492 11533 23493
rect 11467 23428 11468 23492
rect 11532 23428 11533 23492
rect 11467 23427 11533 23428
rect 11470 17781 11530 23427
rect 11467 17780 11533 17781
rect 11467 17716 11468 17780
rect 11532 17716 11533 17780
rect 11467 17715 11533 17716
rect 11283 17644 11349 17645
rect 11283 17580 11284 17644
rect 11348 17580 11349 17644
rect 11283 17579 11349 17580
rect 10716 16832 10724 16896
rect 10788 16832 10804 16896
rect 10868 16832 10884 16896
rect 10948 16832 10964 16896
rect 11028 16832 11036 16896
rect 10716 15808 11036 16832
rect 10716 15744 10724 15808
rect 10788 15744 10804 15808
rect 10868 15744 10884 15808
rect 10948 15744 10964 15808
rect 11028 15744 11036 15808
rect 10716 14720 11036 15744
rect 10716 14656 10724 14720
rect 10788 14656 10804 14720
rect 10868 14656 10884 14720
rect 10948 14656 10964 14720
rect 11028 14656 11036 14720
rect 10716 13632 11036 14656
rect 11654 13701 11714 27643
rect 11838 24989 11898 33491
rect 12022 29749 12082 38795
rect 12203 37228 12269 37229
rect 12203 37164 12204 37228
rect 12268 37164 12269 37228
rect 12203 37163 12269 37164
rect 12019 29748 12085 29749
rect 12019 29684 12020 29748
rect 12084 29684 12085 29748
rect 12019 29683 12085 29684
rect 12206 29477 12266 37163
rect 12203 29476 12269 29477
rect 12203 29412 12204 29476
rect 12268 29412 12269 29476
rect 12203 29411 12269 29412
rect 11835 24988 11901 24989
rect 11835 24924 11836 24988
rect 11900 24924 11901 24988
rect 11835 24923 11901 24924
rect 11835 23492 11901 23493
rect 11835 23428 11836 23492
rect 11900 23428 11901 23492
rect 11835 23427 11901 23428
rect 12019 23492 12085 23493
rect 12019 23428 12020 23492
rect 12084 23428 12085 23492
rect 12019 23427 12085 23428
rect 11838 15605 11898 23427
rect 12022 19413 12082 23427
rect 12571 23084 12637 23085
rect 12571 23020 12572 23084
rect 12636 23020 12637 23084
rect 12571 23019 12637 23020
rect 12019 19412 12085 19413
rect 12019 19348 12020 19412
rect 12084 19348 12085 19412
rect 12019 19347 12085 19348
rect 11835 15604 11901 15605
rect 11835 15540 11836 15604
rect 11900 15540 11901 15604
rect 11835 15539 11901 15540
rect 12574 14925 12634 23019
rect 12571 14924 12637 14925
rect 12571 14860 12572 14924
rect 12636 14860 12637 14924
rect 12571 14859 12637 14860
rect 11651 13700 11717 13701
rect 11651 13636 11652 13700
rect 11716 13636 11717 13700
rect 11651 13635 11717 13636
rect 10716 13568 10724 13632
rect 10788 13568 10804 13632
rect 10868 13568 10884 13632
rect 10948 13568 10964 13632
rect 11028 13568 11036 13632
rect 10716 12544 11036 13568
rect 10716 12480 10724 12544
rect 10788 12480 10804 12544
rect 10868 12480 10884 12544
rect 10948 12480 10964 12544
rect 11028 12480 11036 12544
rect 10547 12340 10613 12341
rect 10547 12276 10548 12340
rect 10612 12276 10613 12340
rect 10547 12275 10613 12276
rect 10056 11936 10064 12000
rect 10128 11936 10144 12000
rect 10208 11936 10224 12000
rect 10288 11936 10304 12000
rect 10368 11936 10376 12000
rect 10056 10912 10376 11936
rect 10056 10848 10064 10912
rect 10128 10848 10144 10912
rect 10208 10848 10224 10912
rect 10288 10848 10304 10912
rect 10368 10848 10376 10912
rect 9811 10028 9877 10029
rect 9811 9964 9812 10028
rect 9876 9964 9877 10028
rect 9811 9963 9877 9964
rect 10056 9824 10376 10848
rect 10056 9760 10064 9824
rect 10128 9760 10144 9824
rect 10208 9760 10224 9824
rect 10288 9760 10304 9824
rect 10368 9760 10376 9824
rect 10056 8736 10376 9760
rect 10716 11456 11036 12480
rect 11099 12476 11165 12477
rect 11099 12412 11100 12476
rect 11164 12412 11165 12476
rect 11099 12411 11165 12412
rect 10716 11392 10724 11456
rect 10788 11392 10804 11456
rect 10868 11392 10884 11456
rect 10948 11392 10964 11456
rect 11028 11392 11036 11456
rect 10716 10368 11036 11392
rect 10716 10304 10724 10368
rect 10788 10304 10804 10368
rect 10868 10304 10884 10368
rect 10948 10304 10964 10368
rect 11028 10304 11036 10368
rect 10547 9484 10613 9485
rect 10547 9420 10548 9484
rect 10612 9420 10613 9484
rect 10547 9419 10613 9420
rect 10056 8672 10064 8736
rect 10128 8672 10144 8736
rect 10208 8672 10224 8736
rect 10288 8672 10304 8736
rect 10368 8672 10376 8736
rect 9443 8124 9509 8125
rect 9443 8060 9444 8124
rect 9508 8060 9509 8124
rect 9443 8059 9509 8060
rect 10056 7648 10376 8672
rect 10056 7584 10064 7648
rect 10128 7584 10144 7648
rect 10208 7584 10224 7648
rect 10288 7584 10304 7648
rect 10368 7584 10376 7648
rect 9075 7444 9141 7445
rect 9075 7380 9076 7444
rect 9140 7380 9141 7444
rect 9075 7379 9141 7380
rect 9811 7308 9877 7309
rect 9811 7244 9812 7308
rect 9876 7244 9877 7308
rect 9811 7243 9877 7244
rect 4316 7040 4324 7104
rect 4388 7040 4404 7104
rect 4468 7040 4484 7104
rect 4548 7040 4564 7104
rect 4628 7040 4636 7104
rect 4316 6016 4636 7040
rect 4316 5952 4324 6016
rect 4388 5952 4404 6016
rect 4468 5952 4484 6016
rect 4548 5952 4564 6016
rect 4628 5952 4636 6016
rect 4316 4928 4636 5952
rect 4316 4864 4324 4928
rect 4388 4864 4404 4928
rect 4468 4864 4484 4928
rect 4548 4864 4564 4928
rect 4628 4864 4636 4928
rect 4316 3840 4636 4864
rect 4316 3776 4324 3840
rect 4388 3776 4404 3840
rect 4468 3776 4484 3840
rect 4548 3776 4564 3840
rect 4628 3776 4636 3840
rect 4316 2752 4636 3776
rect 4316 2688 4324 2752
rect 4388 2688 4404 2752
rect 4468 2688 4484 2752
rect 4548 2688 4564 2752
rect 4628 2688 4636 2752
rect 4316 1664 4636 2688
rect 9814 2549 9874 7243
rect 10056 6560 10376 7584
rect 10550 6901 10610 9419
rect 10716 9280 11036 10304
rect 11102 10029 11162 12411
rect 11099 10028 11165 10029
rect 11099 9964 11100 10028
rect 11164 9964 11165 10028
rect 11099 9963 11165 9964
rect 10716 9216 10724 9280
rect 10788 9216 10804 9280
rect 10868 9216 10884 9280
rect 10948 9216 10964 9280
rect 11028 9216 11036 9280
rect 10716 8192 11036 9216
rect 10716 8128 10724 8192
rect 10788 8128 10804 8192
rect 10868 8128 10884 8192
rect 10948 8128 10964 8192
rect 11028 8128 11036 8192
rect 10716 7104 11036 8128
rect 10716 7040 10724 7104
rect 10788 7040 10804 7104
rect 10868 7040 10884 7104
rect 10948 7040 10964 7104
rect 11028 7040 11036 7104
rect 10547 6900 10613 6901
rect 10547 6836 10548 6900
rect 10612 6836 10613 6900
rect 10547 6835 10613 6836
rect 10056 6496 10064 6560
rect 10128 6496 10144 6560
rect 10208 6496 10224 6560
rect 10288 6496 10304 6560
rect 10368 6496 10376 6560
rect 10056 5472 10376 6496
rect 10056 5408 10064 5472
rect 10128 5408 10144 5472
rect 10208 5408 10224 5472
rect 10288 5408 10304 5472
rect 10368 5408 10376 5472
rect 10056 4384 10376 5408
rect 10056 4320 10064 4384
rect 10128 4320 10144 4384
rect 10208 4320 10224 4384
rect 10288 4320 10304 4384
rect 10368 4320 10376 4384
rect 10056 3296 10376 4320
rect 10056 3232 10064 3296
rect 10128 3232 10144 3296
rect 10208 3232 10224 3296
rect 10288 3232 10304 3296
rect 10368 3232 10376 3296
rect 9811 2548 9877 2549
rect 9811 2484 9812 2548
rect 9876 2484 9877 2548
rect 9811 2483 9877 2484
rect 4316 1600 4324 1664
rect 4388 1600 4404 1664
rect 4468 1600 4484 1664
rect 4548 1600 4564 1664
rect 4628 1600 4636 1664
rect 4316 576 4636 1600
rect 4316 512 4324 576
rect 4388 512 4404 576
rect 4468 512 4484 576
rect 4548 512 4564 576
rect 4628 512 4636 576
rect 4316 496 4636 512
rect 10056 2208 10376 3232
rect 10056 2144 10064 2208
rect 10128 2144 10144 2208
rect 10208 2144 10224 2208
rect 10288 2144 10304 2208
rect 10368 2144 10376 2208
rect 10056 1120 10376 2144
rect 10056 1056 10064 1120
rect 10128 1056 10144 1120
rect 10208 1056 10224 1120
rect 10288 1056 10304 1120
rect 10368 1056 10376 1120
rect 10056 496 10376 1056
rect 10716 6016 11036 7040
rect 10716 5952 10724 6016
rect 10788 5952 10804 6016
rect 10868 5952 10884 6016
rect 10948 5952 10964 6016
rect 11028 5952 11036 6016
rect 10716 4928 11036 5952
rect 10716 4864 10724 4928
rect 10788 4864 10804 4928
rect 10868 4864 10884 4928
rect 10948 4864 10964 4928
rect 11028 4864 11036 4928
rect 10716 3840 11036 4864
rect 10716 3776 10724 3840
rect 10788 3776 10804 3840
rect 10868 3776 10884 3840
rect 10948 3776 10964 3840
rect 11028 3776 11036 3840
rect 10716 2752 11036 3776
rect 10716 2688 10724 2752
rect 10788 2688 10804 2752
rect 10868 2688 10884 2752
rect 10948 2688 10964 2752
rect 11028 2688 11036 2752
rect 10716 1664 11036 2688
rect 10716 1600 10724 1664
rect 10788 1600 10804 1664
rect 10868 1600 10884 1664
rect 10948 1600 10964 1664
rect 11028 1600 11036 1664
rect 10716 576 11036 1600
rect 10716 512 10724 576
rect 10788 512 10804 576
rect 10868 512 10884 576
rect 10948 512 10964 576
rect 11028 512 11036 576
rect 10716 496 11036 512
use sky130_fd_sc_hd__inv_2  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8096 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1762784779
transform 1 0 10948 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1762784779
transform 1 0 9384 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1762784779
transform -1 0 10396 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1762784779
transform 1 0 10672 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1762784779
transform -1 0 10672 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1762784779
transform 1 0 5888 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1762784779
transform 1 0 4416 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1762784779
transform -1 0 6164 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0863_
timestamp 1762784779
transform 1 0 8280 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1762784779
transform 1 0 5428 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1762784779
transform -1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5796 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0867_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7268 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0868_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 6072 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0869_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5428 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0870_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5520 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0871_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4876 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_2  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4784 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0873_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3680 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0874_
timestamp 1762784779
transform 1 0 3220 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0875_
timestamp 1762784779
transform 1 0 3220 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0876_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 2208 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 1762784779
transform 1 0 1472 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0878_
timestamp 1762784779
transform 1 0 828 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1762784779
transform -1 0 3128 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0880_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1656 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0881_
timestamp 1762784779
transform 1 0 1196 0 1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 1762784779
transform 1 0 11500 0 -1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0883_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 11500 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0884_
timestamp 1762784779
transform 1 0 8924 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0885_
timestamp 1762784779
transform 1 0 11592 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0886_
timestamp 1762784779
transform -1 0 12328 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8740 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0888_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 9384 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3772 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0890_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 7268 0 1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0891_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4692 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0892_
timestamp 1762784779
transform 1 0 3956 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 3496 0 -1 32096
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _0894_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 2668 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_4  _0895_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4692 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _0896_
timestamp 1762784779
transform -1 0 5704 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1762784779
transform 1 0 8740 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1762784779
transform -1 0 8188 0 1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0899_
timestamp 1762784779
transform 1 0 5704 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0900_
timestamp 1762784779
transform 1 0 5796 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0901_
timestamp 1762784779
transform 1 0 6808 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1762784779
transform 1 0 7360 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0903_
timestamp 1762784779
transform 1 0 4048 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0904_
timestamp 1762784779
transform -1 0 5704 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0905_
timestamp 1762784779
transform 1 0 8832 0 -1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1762784779
transform -1 0 5152 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1762784779
transform -1 0 4324 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0908_
timestamp 1762784779
transform -1 0 1472 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1762784779
transform -1 0 8280 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0910_
timestamp 1762784779
transform 1 0 8832 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1762784779
transform 1 0 5796 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1762784779
transform -1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0913_
timestamp 1762784779
transform 1 0 8004 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1762784779
transform 1 0 6624 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0915_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8188 0 -1 39712
box -38 -48 1234 592
use sky130_fd_sc_hd__a31o_2  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 9660 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0917_
timestamp 1762784779
transform 1 0 9936 0 1 40800
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 9016 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0919_
timestamp 1762784779
transform 1 0 8372 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0920_
timestamp 1762784779
transform -1 0 10304 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 9016 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 1762784779
transform 1 0 9476 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8280 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0924_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8004 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1762784779
transform 1 0 8004 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0926_
timestamp 1762784779
transform 1 0 8372 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6900 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0928_
timestamp 1762784779
transform 1 0 9384 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0929_
timestamp 1762784779
transform 1 0 10120 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8924 0 -1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 8372 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0932_
timestamp 1762784779
transform 1 0 7636 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0933_
timestamp 1762784779
transform 1 0 7820 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0934_
timestamp 1762784779
transform 1 0 8832 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1762784779
transform 1 0 10120 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0936_
timestamp 1762784779
transform -1 0 9936 0 1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _0937_
timestamp 1762784779
transform 1 0 8372 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0938_
timestamp 1762784779
transform -1 0 9200 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0939_
timestamp 1762784779
transform 1 0 8280 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1762784779
transform -1 0 7728 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0941_
timestamp 1762784779
transform 1 0 11868 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0942_
timestamp 1762784779
transform -1 0 9384 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0943_
timestamp 1762784779
transform 1 0 7084 0 1 34272
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2b_1  _0944_
timestamp 1762784779
transform 1 0 10028 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0945_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 9568 0 -1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _0946_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 8832 0 -1 40800
box -38 -48 2062 592
use sky130_fd_sc_hd__o311a_1  _0947_
timestamp 1762784779
transform 1 0 8096 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0948_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6532 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0949_
timestamp 1762784779
transform -1 0 9476 0 1 41888
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0950_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8832 0 -1 41888
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0951_
timestamp 1762784779
transform -1 0 7820 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0952_
timestamp 1762784779
transform -1 0 8832 0 -1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _0953_
timestamp 1762784779
transform 1 0 7176 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0954_
timestamp 1762784779
transform -1 0 7728 0 1 39712
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _0955_
timestamp 1762784779
transform 1 0 7084 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7820 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_4  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 7452 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _0958_
timestamp 1762784779
transform -1 0 3588 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0959_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 2576 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0960_
timestamp 1762784779
transform 1 0 3496 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0961_
timestamp 1762784779
transform 1 0 10488 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6256 0 1 28832
box -38 -48 1694 592
use sky130_fd_sc_hd__mux2_1  _0963_
timestamp 1762784779
transform -1 0 9200 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _0964_
timestamp 1762784779
transform 1 0 4140 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0965_
timestamp 1762784779
transform -1 0 5152 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0966_
timestamp 1762784779
transform 1 0 6808 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0967_
timestamp 1762784779
transform 1 0 4968 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0968_
timestamp 1762784779
transform 1 0 8464 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0969_
timestamp 1762784779
transform 1 0 3956 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1762784779
transform 1 0 8372 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _0971_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7728 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0972_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 6624 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0973_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4140 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0974_
timestamp 1762784779
transform -1 0 6900 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0975_
timestamp 1762784779
transform 1 0 7636 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0976_
timestamp 1762784779
transform -1 0 7268 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0977_
timestamp 1762784779
transform -1 0 8740 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1762784779
transform -1 0 8280 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _0979_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4324 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 4692 0 1 36448
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0981_
timestamp 1762784779
transform -1 0 4508 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0982_
timestamp 1762784779
transform 1 0 4324 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0983_
timestamp 1762784779
transform 1 0 7452 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0984_
timestamp 1762784779
transform 1 0 5796 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1762784779
transform -1 0 5060 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0986_
timestamp 1762784779
transform 1 0 5060 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0987_
timestamp 1762784779
transform 1 0 2668 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1762784779
transform -1 0 2668 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _0989_
timestamp 1762784779
transform -1 0 4048 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_1  _0990_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3312 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_4  _0991_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 2300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _0992_
timestamp 1762784779
transform 1 0 2208 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0993_
timestamp 1762784779
transform -1 0 3772 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0994_
timestamp 1762784779
transform 1 0 3404 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0995_
timestamp 1762784779
transform 1 0 11224 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0996_
timestamp 1762784779
transform 1 0 10396 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0997_
timestamp 1762784779
transform 1 0 10948 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1762784779
transform 1 0 11868 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0999_
timestamp 1762784779
transform 1 0 10396 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1000_
timestamp 1762784779
transform 1 0 10856 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1001_
timestamp 1762784779
transform 1 0 4784 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1002_
timestamp 1762784779
transform -1 0 5980 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1003_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 10212 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1004_
timestamp 1762784779
transform 1 0 10304 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1005_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3956 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_4  _1006_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 5704 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__xnor2_1  _1007_
timestamp 1762784779
transform -1 0 9936 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1008_
timestamp 1762784779
transform 1 0 9384 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7728 0 1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _1010_
timestamp 1762784779
transform 1 0 6992 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1011_
timestamp 1762784779
transform 1 0 7912 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1012_
timestamp 1762784779
transform 1 0 8556 0 -1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1762784779
transform -1 0 8648 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1014_
timestamp 1762784779
transform -1 0 9292 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1015_
timestamp 1762784779
transform 1 0 9108 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1016_
timestamp 1762784779
transform 1 0 8924 0 -1 29920
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 1762784779
transform 1 0 10028 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1018_
timestamp 1762784779
transform 1 0 9108 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1019_
timestamp 1762784779
transform -1 0 10396 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1020_
timestamp 1762784779
transform 1 0 9200 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1762784779
transform 1 0 9936 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1022_
timestamp 1762784779
transform 1 0 9384 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1023_
timestamp 1762784779
transform 1 0 8740 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1024_
timestamp 1762784779
transform 1 0 8096 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _1025_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3496 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1026_
timestamp 1762784779
transform 1 0 2668 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1027_
timestamp 1762784779
transform 1 0 1564 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1028_
timestamp 1762784779
transform -1 0 2116 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1029_
timestamp 1762784779
transform 1 0 2392 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1762784779
transform -1 0 6440 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1031_
timestamp 1762784779
transform 1 0 5060 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1032_
timestamp 1762784779
transform 1 0 10120 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1033_
timestamp 1762784779
transform 1 0 9660 0 -1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1034_
timestamp 1762784779
transform -1 0 10396 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1035_
timestamp 1762784779
transform -1 0 10028 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1036_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 10028 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _1037_
timestamp 1762784779
transform -1 0 10028 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1038_
timestamp 1762784779
transform 1 0 9384 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1039_
timestamp 1762784779
transform -1 0 10028 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1040_
timestamp 1762784779
transform -1 0 9384 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1041_
timestamp 1762784779
transform -1 0 7912 0 -1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__o22a_1  _1042_
timestamp 1762784779
transform 1 0 7912 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1043_
timestamp 1762784779
transform 1 0 7084 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1044_
timestamp 1762784779
transform 1 0 10028 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1762784779
transform -1 0 9108 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1046_
timestamp 1762784779
transform 1 0 9108 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1047_
timestamp 1762784779
transform 1 0 11408 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1048_
timestamp 1762784779
transform 1 0 10396 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1049_
timestamp 1762784779
transform 1 0 10948 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1050_
timestamp 1762784779
transform 1 0 11040 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1762784779
transform 1 0 10396 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1052_
timestamp 1762784779
transform -1 0 12144 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 1762784779
transform 1 0 12052 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_1  _1054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 12328 0 1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _1055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 11500 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1056_
timestamp 1762784779
transform 1 0 11500 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1057_
timestamp 1762784779
transform 1 0 10580 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1058_
timestamp 1762784779
transform 1 0 10948 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1059_
timestamp 1762784779
transform -1 0 9384 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1060_
timestamp 1762784779
transform 1 0 8648 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1762784779
transform -1 0 6992 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1062_
timestamp 1762784779
transform 1 0 6256 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1063_
timestamp 1762784779
transform 1 0 4048 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1064_
timestamp 1762784779
transform 1 0 1932 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1065_
timestamp 1762784779
transform -1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1066_
timestamp 1762784779
transform 1 0 2300 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1067_
timestamp 1762784779
transform -1 0 3956 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1068_
timestamp 1762784779
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1069_
timestamp 1762784779
transform 1 0 10028 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1070_
timestamp 1762784779
transform 1 0 9752 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1071_
timestamp 1762784779
transform -1 0 10396 0 1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1072_
timestamp 1762784779
transform 1 0 9476 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1073_
timestamp 1762784779
transform 1 0 10672 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1074_
timestamp 1762784779
transform 1 0 9660 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1075_
timestamp 1762784779
transform -1 0 10120 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1762784779
transform 1 0 9476 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1077_
timestamp 1762784779
transform 1 0 9752 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1078_
timestamp 1762784779
transform -1 0 9568 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _1079_
timestamp 1762784779
transform 1 0 5520 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1080_
timestamp 1762784779
transform 1 0 7176 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1081_
timestamp 1762784779
transform 1 0 8372 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1082_
timestamp 1762784779
transform 1 0 9108 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1083_
timestamp 1762784779
transform -1 0 10304 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1762784779
transform -1 0 11592 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1085_
timestamp 1762784779
transform 1 0 10764 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1086_
timestamp 1762784779
transform 1 0 10948 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1087_
timestamp 1762784779
transform 1 0 11040 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1088_
timestamp 1762784779
transform -1 0 10856 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1762784779
transform 1 0 11408 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 1762784779
transform -1 0 12236 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1091_
timestamp 1762784779
transform -1 0 12052 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp 1762784779
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 1762784779
transform -1 0 10580 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1094_
timestamp 1762784779
transform 1 0 11500 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1095_
timestamp 1762784779
transform 1 0 10304 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1096_
timestamp 1762784779
transform -1 0 10304 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1097_
timestamp 1762784779
transform 1 0 8280 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1098_
timestamp 1762784779
transform -1 0 3220 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1099_
timestamp 1762784779
transform -1 0 2576 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1100_
timestamp 1762784779
transform 1 0 3220 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1101_
timestamp 1762784779
transform -1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1102_
timestamp 1762784779
transform 1 0 2300 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1103_
timestamp 1762784779
transform -1 0 3404 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1104_
timestamp 1762784779
transform -1 0 3404 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1105_
timestamp 1762784779
transform -1 0 8832 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1106_
timestamp 1762784779
transform -1 0 8280 0 -1 9248
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1107_
timestamp 1762784779
transform 1 0 8372 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1108_
timestamp 1762784779
transform 1 0 9108 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1109_
timestamp 1762784779
transform 1 0 8740 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1110_
timestamp 1762784779
transform 1 0 8556 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 10672 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1112_
timestamp 1762784779
transform -1 0 10212 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1113_
timestamp 1762784779
transform -1 0 9936 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1114_
timestamp 1762784779
transform 1 0 9384 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _1115_
timestamp 1762784779
transform 1 0 5796 0 -1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1762784779
transform -1 0 5888 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1117_
timestamp 1762784779
transform 1 0 8372 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1118_
timestamp 1762784779
transform 1 0 9292 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1119_
timestamp 1762784779
transform -1 0 10488 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1762784779
transform -1 0 10120 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1121_
timestamp 1762784779
transform 1 0 10948 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1762784779
transform 1 0 9568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1123_
timestamp 1762784779
transform -1 0 11592 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1124_
timestamp 1762784779
transform -1 0 11316 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1125_
timestamp 1762784779
transform 1 0 10672 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1762784779
transform -1 0 11040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1127_
timestamp 1762784779
transform 1 0 9752 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1762784779
transform 1 0 10488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1129_
timestamp 1762784779
transform -1 0 11316 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1130_
timestamp 1762784779
transform 1 0 10948 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 1762784779
transform 1 0 10948 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1762784779
transform -1 0 11868 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1762784779
transform -1 0 10764 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1134_
timestamp 1762784779
transform 1 0 9384 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1762784779
transform 1 0 8464 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1136_
timestamp 1762784779
transform -1 0 2852 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1137_
timestamp 1762784779
transform -1 0 2668 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1138_
timestamp 1762784779
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1139_
timestamp 1762784779
transform -1 0 2024 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1140_
timestamp 1762784779
transform 1 0 2392 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1141_
timestamp 1762784779
transform -1 0 5520 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1762784779
transform -1 0 5796 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1762784779
transform 1 0 4784 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1144_
timestamp 1762784779
transform 1 0 9200 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1145_
timestamp 1762784779
transform 1 0 5244 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1146_
timestamp 1762784779
transform 1 0 7452 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1762784779
transform -1 0 7452 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1148_
timestamp 1762784779
transform -1 0 6808 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1149_
timestamp 1762784779
transform -1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1150_
timestamp 1762784779
transform -1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1762784779
transform -1 0 8556 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _1152_
timestamp 1762784779
transform 1 0 7268 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1153_
timestamp 1762784779
transform 1 0 7636 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1154_
timestamp 1762784779
transform 1 0 8740 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1155_
timestamp 1762784779
transform 1 0 6164 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_2  _1156_
timestamp 1762784779
transform 1 0 4508 0 1 27744
box -38 -48 1694 592
use sky130_fd_sc_hd__o22a_1  _1157_
timestamp 1762784779
transform 1 0 5888 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1158_
timestamp 1762784779
transform 1 0 5336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1159_
timestamp 1762784779
transform 1 0 7820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1160_
timestamp 1762784779
transform 1 0 7636 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1161_
timestamp 1762784779
transform 1 0 7084 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1162_
timestamp 1762784779
transform 1 0 9108 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1163_
timestamp 1762784779
transform 1 0 9476 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 10948 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1165_
timestamp 1762784779
transform -1 0 10396 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1166_
timestamp 1762784779
transform 1 0 8924 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1167_
timestamp 1762784779
transform 1 0 11040 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1168_
timestamp 1762784779
transform -1 0 9660 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1169_
timestamp 1762784779
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1170_
timestamp 1762784779
transform 1 0 9384 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1762784779
transform -1 0 10488 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1172_
timestamp 1762784779
transform 1 0 7636 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1173_
timestamp 1762784779
transform -1 0 8740 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1174_
timestamp 1762784779
transform 1 0 5704 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1175_
timestamp 1762784779
transform 1 0 5796 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1176_
timestamp 1762784779
transform 1 0 4232 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1177_
timestamp 1762784779
transform 1 0 1932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1178_
timestamp 1762784779
transform -1 0 2208 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1179_
timestamp 1762784779
transform 1 0 2576 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1180_
timestamp 1762784779
transform 1 0 4232 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1762784779
transform -1 0 3128 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1182_
timestamp 1762784779
transform -1 0 3496 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1183_
timestamp 1762784779
transform 1 0 7728 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1184_
timestamp 1762784779
transform 1 0 4600 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1185_
timestamp 1762784779
transform 1 0 2852 0 -1 8160
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1186_
timestamp 1762784779
transform 1 0 4508 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1187_
timestamp 1762784779
transform 1 0 5980 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1188_
timestamp 1762784779
transform -1 0 6348 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1762784779
transform -1 0 5704 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1190_
timestamp 1762784779
transform 1 0 5152 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1191_
timestamp 1762784779
transform -1 0 7268 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__mux4_2  _1192_
timestamp 1762784779
transform 1 0 4048 0 -1 28832
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1762784779
transform 1 0 4968 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1194_
timestamp 1762784779
transform 1 0 5796 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1195_
timestamp 1762784779
transform 1 0 4968 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1196_
timestamp 1762784779
transform -1 0 6716 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1762784779
transform -1 0 6440 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1198_
timestamp 1762784779
transform -1 0 6992 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1199_
timestamp 1762784779
transform 1 0 7636 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1200_
timestamp 1762784779
transform 1 0 6348 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1762784779
transform 1 0 6440 0 1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1202_
timestamp 1762784779
transform 1 0 6900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1203_
timestamp 1762784779
transform 1 0 6992 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1204_
timestamp 1762784779
transform 1 0 5612 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1762784779
transform 1 0 6624 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 1762784779
transform -1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1207_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 9844 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1208_
timestamp 1762784779
transform 1 0 6532 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1209_
timestamp 1762784779
transform 1 0 7176 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1210_
timestamp 1762784779
transform 1 0 6900 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1211_
timestamp 1762784779
transform -1 0 7360 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1212_
timestamp 1762784779
transform 1 0 6348 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1213_
timestamp 1762784779
transform -1 0 4416 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1214_
timestamp 1762784779
transform 1 0 3128 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1215_
timestamp 1762784779
transform 1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1216_
timestamp 1762784779
transform 1 0 2300 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1217_
timestamp 1762784779
transform -1 0 2024 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1218_
timestamp 1762784779
transform 1 0 3496 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1219_
timestamp 1762784779
transform -1 0 2300 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1762784779
transform -1 0 3772 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1221_
timestamp 1762784779
transform 1 0 2392 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1222_
timestamp 1762784779
transform -1 0 6808 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1223_
timestamp 1762784779
transform -1 0 5060 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _1224_
timestamp 1762784779
transform 1 0 2300 0 -1 10336
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1225_
timestamp 1762784779
transform 1 0 4048 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1226_
timestamp 1762784779
transform 1 0 5796 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 1762784779
transform -1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1228_
timestamp 1762784779
transform -1 0 5612 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 1762784779
transform -1 0 5704 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1230_
timestamp 1762784779
transform -1 0 6440 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _1231_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 5612 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1232_
timestamp 1762784779
transform -1 0 5520 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1233_
timestamp 1762784779
transform -1 0 6992 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1234_
timestamp 1762784779
transform 1 0 6072 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1235_
timestamp 1762784779
transform 1 0 4048 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1236_
timestamp 1762784779
transform 1 0 4692 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1237_
timestamp 1762784779
transform 1 0 4324 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1238_
timestamp 1762784779
transform 1 0 4968 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1762784779
transform 1 0 5612 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1240_
timestamp 1762784779
transform 1 0 5152 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1241_
timestamp 1762784779
transform -1 0 6164 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1242_
timestamp 1762784779
transform -1 0 5520 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1243_
timestamp 1762784779
transform 1 0 4876 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1762784779
transform 1 0 4876 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1245_
timestamp 1762784779
transform 1 0 5796 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1246_
timestamp 1762784779
transform -1 0 5888 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1247_
timestamp 1762784779
transform -1 0 5428 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1248_
timestamp 1762784779
transform 1 0 5336 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1249_
timestamp 1762784779
transform -1 0 5704 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1250_
timestamp 1762784779
transform 1 0 5796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1251_
timestamp 1762784779
transform 1 0 3036 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1252_
timestamp 1762784779
transform 1 0 3128 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1253_
timestamp 1762784779
transform -1 0 3680 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1254_
timestamp 1762784779
transform 1 0 1196 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _1255_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 3036 0 1 32096
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_1  _1256_
timestamp 1762784779
transform -1 0 6532 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1257_
timestamp 1762784779
transform -1 0 7084 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1258_
timestamp 1762784779
transform -1 0 7728 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1259_
timestamp 1762784779
transform 1 0 6624 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1260_
timestamp 1762784779
transform -1 0 9384 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1261_
timestamp 1762784779
transform 1 0 8188 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _1262_
timestamp 1762784779
transform 1 0 7268 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1762784779
transform -1 0 7176 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1264_
timestamp 1762784779
transform -1 0 6440 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1265_
timestamp 1762784779
transform 1 0 2392 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1762784779
transform 1 0 2116 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_4  _1267_
timestamp 1762784779
transform -1 0 2392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1268_
timestamp 1762784779
transform 1 0 6532 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1269_
timestamp 1762784779
transform 1 0 7636 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1270_
timestamp 1762784779
transform 1 0 8372 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1271_
timestamp 1762784779
transform 1 0 9476 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1272_
timestamp 1762784779
transform 1 0 11040 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 1762784779
transform 1 0 10948 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1762784779
transform 1 0 11776 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1275_
timestamp 1762784779
transform -1 0 11776 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1276_
timestamp 1762784779
transform 1 0 11132 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1277_
timestamp 1762784779
transform 1 0 11776 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1278_
timestamp 1762784779
transform -1 0 12236 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1279_
timestamp 1762784779
transform 1 0 11224 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1280_
timestamp 1762784779
transform -1 0 12052 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1281_
timestamp 1762784779
transform 1 0 9108 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1282_
timestamp 1762784779
transform 1 0 7268 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1283_
timestamp 1762784779
transform 1 0 7728 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1284_
timestamp 1762784779
transform 1 0 7176 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1285_
timestamp 1762784779
transform 1 0 3220 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1286_
timestamp 1762784779
transform 1 0 2116 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1287_
timestamp 1762784779
transform -1 0 1564 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1288_
timestamp 1762784779
transform -1 0 1932 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1289_
timestamp 1762784779
transform -1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1290_
timestamp 1762784779
transform 1 0 11224 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1291_
timestamp 1762784779
transform -1 0 12328 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1292_
timestamp 1762784779
transform 1 0 11408 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1293_
timestamp 1762784779
transform -1 0 12328 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1762784779
transform 1 0 10948 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1295_
timestamp 1762784779
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1296_
timestamp 1762784779
transform 1 0 11684 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1297_
timestamp 1762784779
transform 1 0 11408 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1298_
timestamp 1762784779
transform 1 0 11776 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1299_
timestamp 1762784779
transform 1 0 11592 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1300_
timestamp 1762784779
transform 1 0 6900 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1301_
timestamp 1762784779
transform -1 0 7452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1302_
timestamp 1762784779
transform 1 0 8372 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1303_
timestamp 1762784779
transform 1 0 7728 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1304_
timestamp 1762784779
transform 1 0 7544 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1305_
timestamp 1762784779
transform -1 0 9108 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1306_
timestamp 1762784779
transform 1 0 8372 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1307_
timestamp 1762784779
transform 1 0 7912 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1308_
timestamp 1762784779
transform 1 0 7452 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1309_
timestamp 1762784779
transform 1 0 6256 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1310_
timestamp 1762784779
transform 1 0 4048 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1311_
timestamp 1762784779
transform 1 0 920 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1312_
timestamp 1762784779
transform -1 0 2116 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1313_
timestamp 1762784779
transform -1 0 12236 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1314_
timestamp 1762784779
transform 1 0 9844 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1315_
timestamp 1762784779
transform -1 0 11592 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1316_
timestamp 1762784779
transform 1 0 10948 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1317_
timestamp 1762784779
transform -1 0 11224 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1318_
timestamp 1762784779
transform 1 0 11408 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1319_
timestamp 1762784779
transform 1 0 10488 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1320_
timestamp 1762784779
transform -1 0 11776 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1321_
timestamp 1762784779
transform 1 0 10948 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1322_
timestamp 1762784779
transform -1 0 12144 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1323_
timestamp 1762784779
transform 1 0 11592 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1324_
timestamp 1762784779
transform -1 0 7084 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1325_
timestamp 1762784779
transform 1 0 7636 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1326_
timestamp 1762784779
transform -1 0 7452 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1327_
timestamp 1762784779
transform 1 0 9200 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1328_
timestamp 1762784779
transform 1 0 10028 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _1329_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 9384 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1330_
timestamp 1762784779
transform -1 0 10028 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1331_
timestamp 1762784779
transform 1 0 8464 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1332_
timestamp 1762784779
transform -1 0 9016 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1333_
timestamp 1762784779
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1762784779
transform 1 0 4600 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1335_
timestamp 1762784779
transform 1 0 1380 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1336_
timestamp 1762784779
transform -1 0 1932 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1762784779
transform 1 0 7636 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1338_
timestamp 1762784779
transform -1 0 7912 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1339_
timestamp 1762784779
transform -1 0 9016 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1340_
timestamp 1762784779
transform -1 0 7912 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1341_
timestamp 1762784779
transform 1 0 8740 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1342_
timestamp 1762784779
transform 1 0 9200 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1343_
timestamp 1762784779
transform 1 0 9384 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1344_
timestamp 1762784779
transform 1 0 9660 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1345_
timestamp 1762784779
transform 1 0 10304 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1346_
timestamp 1762784779
transform 1 0 9568 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1762784779
transform 1 0 9108 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1348_
timestamp 1762784779
transform -1 0 11040 0 1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1762784779
transform -1 0 10856 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _1350_
timestamp 1762784779
transform -1 0 11408 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1351_
timestamp 1762784779
transform 1 0 9752 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1352_
timestamp 1762784779
transform -1 0 10856 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1353_
timestamp 1762784779
transform -1 0 8740 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1354_
timestamp 1762784779
transform 1 0 7452 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1355_
timestamp 1762784779
transform 1 0 3220 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1356_
timestamp 1762784779
transform 1 0 3404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1357_
timestamp 1762784779
transform 1 0 2484 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1358_
timestamp 1762784779
transform -1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__a31o_1  _1359_
timestamp 1762784779
transform 1 0 7084 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1360_
timestamp 1762784779
transform 1 0 9016 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1361_
timestamp 1762784779
transform 1 0 6624 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1362_
timestamp 1762784779
transform 1 0 6808 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1363_
timestamp 1762784779
transform -1 0 7728 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1364_
timestamp 1762784779
transform 1 0 6716 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1365_
timestamp 1762784779
transform 1 0 5428 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1366_
timestamp 1762784779
transform 1 0 5796 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1367_
timestamp 1762784779
transform -1 0 6348 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1368_
timestamp 1762784779
transform 1 0 10028 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1369_
timestamp 1762784779
transform 1 0 6256 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1370_
timestamp 1762784779
transform -1 0 7820 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1371_
timestamp 1762784779
transform 1 0 6900 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1372_
timestamp 1762784779
transform 1 0 5796 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1373_
timestamp 1762784779
transform -1 0 6900 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1374_
timestamp 1762784779
transform 1 0 5980 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1375_
timestamp 1762784779
transform -1 0 6900 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _1376_
timestamp 1762784779
transform 1 0 6440 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1377_
timestamp 1762784779
transform 1 0 5888 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1378_
timestamp 1762784779
transform -1 0 5244 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1379_
timestamp 1762784779
transform 1 0 4232 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1380_
timestamp 1762784779
transform 1 0 1748 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1381_
timestamp 1762784779
transform -1 0 2024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1382_
timestamp 1762784779
transform -1 0 3128 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1383_
timestamp 1762784779
transform 1 0 7360 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1384_
timestamp 1762784779
transform 1 0 3128 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1385_
timestamp 1762784779
transform 1 0 4140 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1386_
timestamp 1762784779
transform 1 0 4784 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1387_
timestamp 1762784779
transform 1 0 3864 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1388_
timestamp 1762784779
transform -1 0 4232 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1389_
timestamp 1762784779
transform 1 0 3220 0 1 544
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1390_
timestamp 1762784779
transform 1 0 3680 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1391_
timestamp 1762784779
transform 1 0 5796 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1392_
timestamp 1762784779
transform 1 0 3404 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1393_
timestamp 1762784779
transform 1 0 4692 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1394_
timestamp 1762784779
transform 1 0 4140 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1395_
timestamp 1762784779
transform 1 0 4784 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1396_
timestamp 1762784779
transform -1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1397_
timestamp 1762784779
transform 1 0 3956 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1762784779
transform 1 0 5428 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1399_
timestamp 1762784779
transform 1 0 4416 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1400_
timestamp 1762784779
transform 1 0 3680 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1401_
timestamp 1762784779
transform 1 0 3496 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1402_
timestamp 1762784779
transform -1 0 4232 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1403_
timestamp 1762784779
transform 1 0 3772 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1404_
timestamp 1762784779
transform -1 0 2576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1405_
timestamp 1762784779
transform 1 0 2300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1406_
timestamp 1762784779
transform 1 0 920 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1407_
timestamp 1762784779
transform 1 0 4232 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1408_
timestamp 1762784779
transform 1 0 2300 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1409_
timestamp 1762784779
transform 1 0 3220 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1410_
timestamp 1762784779
transform 1 0 1656 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1411_
timestamp 1762784779
transform 1 0 2300 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1412_
timestamp 1762784779
transform 1 0 2944 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1413_
timestamp 1762784779
transform 1 0 3588 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1414_
timestamp 1762784779
transform -1 0 4324 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1415_
timestamp 1762784779
transform -1 0 5060 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1416_
timestamp 1762784779
transform 1 0 3588 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1417_
timestamp 1762784779
transform 1 0 4508 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1418_
timestamp 1762784779
transform -1 0 4876 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1419_
timestamp 1762784779
transform 1 0 4324 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1420_
timestamp 1762784779
transform 1 0 3864 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1421_
timestamp 1762784779
transform 1 0 3496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1422_
timestamp 1762784779
transform -1 0 3036 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1423_
timestamp 1762784779
transform -1 0 3128 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1424_
timestamp 1762784779
transform 1 0 2024 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1425_
timestamp 1762784779
transform -1 0 2024 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1426_
timestamp 1762784779
transform -1 0 11408 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1427_
timestamp 1762784779
transform -1 0 10856 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1762784779
transform -1 0 10304 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1429_
timestamp 1762784779
transform 1 0 9752 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1430_
timestamp 1762784779
transform 1 0 11592 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1431_
timestamp 1762784779
transform 1 0 10856 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1432_
timestamp 1762784779
transform -1 0 11408 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1433_
timestamp 1762784779
transform -1 0 11592 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1434_
timestamp 1762784779
transform -1 0 10580 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1435_
timestamp 1762784779
transform 1 0 10396 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1436_
timestamp 1762784779
transform 1 0 5796 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1437_
timestamp 1762784779
transform 1 0 5980 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1438_
timestamp 1762784779
transform 1 0 7084 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1439_
timestamp 1762784779
transform 1 0 7728 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1762784779
transform -1 0 9476 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1441_
timestamp 1762784779
transform -1 0 9568 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1442_
timestamp 1762784779
transform -1 0 9752 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1443_
timestamp 1762784779
transform 1 0 6624 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1444_
timestamp 1762784779
transform 1 0 2208 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1445_
timestamp 1762784779
transform 1 0 2760 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_4  _1446_
timestamp 1762784779
transform -1 0 2208 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_1  _1447_
timestamp 1762784779
transform 1 0 9292 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1448_
timestamp 1762784779
transform -1 0 10764 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1449_
timestamp 1762784779
transform 1 0 9752 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1450_
timestamp 1762784779
transform 1 0 10028 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1451_
timestamp 1762784779
transform 1 0 9844 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1452_
timestamp 1762784779
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1453_
timestamp 1762784779
transform -1 0 12144 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp 1762784779
transform -1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1455_
timestamp 1762784779
transform 1 0 11408 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1456_
timestamp 1762784779
transform -1 0 11592 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1762784779
transform -1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1458_
timestamp 1762784779
transform -1 0 10856 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1459_
timestamp 1762784779
transform 1 0 6992 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1460_
timestamp 1762784779
transform 1 0 7452 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1461_
timestamp 1762784779
transform 1 0 7636 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1462_
timestamp 1762784779
transform 1 0 8648 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1463_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 9016 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1464_
timestamp 1762784779
transform 1 0 10304 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1465_
timestamp 1762784779
transform 1 0 8372 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1466_
timestamp 1762784779
transform 1 0 2576 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1467_
timestamp 1762784779
transform 1 0 2300 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1468_
timestamp 1762784779
transform -1 0 2208 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_4  _1469_
timestamp 1762784779
transform -1 0 2208 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1470_
timestamp 1762784779
transform 1 0 9292 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1471_
timestamp 1762784779
transform 1 0 8280 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1472_
timestamp 1762784779
transform 1 0 7636 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1473_
timestamp 1762784779
transform 1 0 8372 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1474_
timestamp 1762784779
transform -1 0 9568 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1475_
timestamp 1762784779
transform 1 0 8372 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1476_
timestamp 1762784779
transform 1 0 9016 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_2  _1477_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 10856 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1478_
timestamp 1762784779
transform 1 0 8832 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1479_
timestamp 1762784779
transform -1 0 10120 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1480_
timestamp 1762784779
transform -1 0 7728 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1481_
timestamp 1762784779
transform 1 0 7452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1762784779
transform 1 0 8464 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1483_
timestamp 1762784779
transform 1 0 8556 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1484_
timestamp 1762784779
transform 1 0 9660 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1485_
timestamp 1762784779
transform 1 0 8924 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1486_
timestamp 1762784779
transform 1 0 9108 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1487_
timestamp 1762784779
transform -1 0 6992 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1488_
timestamp 1762784779
transform 1 0 5612 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1489_
timestamp 1762784779
transform 1 0 4048 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1490_
timestamp 1762784779
transform 1 0 2392 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1491_
timestamp 1762784779
transform -1 0 2024 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1492_
timestamp 1762784779
transform 1 0 8004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1493_
timestamp 1762784779
transform 1 0 7084 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1494_
timestamp 1762784779
transform 1 0 8740 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1495_
timestamp 1762784779
transform 1 0 8372 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1496_
timestamp 1762784779
transform 1 0 8372 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1497_
timestamp 1762784779
transform -1 0 9016 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1498_
timestamp 1762784779
transform -1 0 8740 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1499_
timestamp 1762784779
transform 1 0 9016 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1500_
timestamp 1762784779
transform 1 0 7820 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1501_
timestamp 1762784779
transform 1 0 8464 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1502_
timestamp 1762784779
transform 1 0 7636 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1503_
timestamp 1762784779
transform -1 0 8280 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1504_
timestamp 1762784779
transform 1 0 6992 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1505_
timestamp 1762784779
transform 1 0 8372 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1506_
timestamp 1762784779
transform 1 0 8740 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1507_
timestamp 1762784779
transform -1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1508_
timestamp 1762784779
transform 1 0 7636 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1509_
timestamp 1762784779
transform 1 0 3220 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1510_
timestamp 1762784779
transform 1 0 4600 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1511_
timestamp 1762784779
transform 1 0 2944 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1512_
timestamp 1762784779
transform 1 0 3220 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_1  _1513_
timestamp 1762784779
transform 1 0 7820 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1514_
timestamp 1762784779
transform 1 0 4876 0 1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1762784779
transform -1 0 6164 0 1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1516_
timestamp 1762784779
transform -1 0 5060 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1517_
timestamp 1762784779
transform 1 0 5060 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1518_
timestamp 1762784779
transform 1 0 9016 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1519_
timestamp 1762784779
transform -1 0 4876 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1520_
timestamp 1762784779
transform -1 0 5520 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1521_
timestamp 1762784779
transform -1 0 6532 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1522_
timestamp 1762784779
transform 1 0 5336 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1523_
timestamp 1762784779
transform 1 0 5980 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1524_
timestamp 1762784779
transform 1 0 6532 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1525_
timestamp 1762784779
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1526_
timestamp 1762784779
transform 1 0 5612 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1527_
timestamp 1762784779
transform -1 0 7084 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1528_
timestamp 1762784779
transform 1 0 6716 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1529_
timestamp 1762784779
transform -1 0 7084 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1530_
timestamp 1762784779
transform 1 0 6256 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1762784779
transform -1 0 2944 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1532_
timestamp 1762784779
transform 1 0 2668 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1533_
timestamp 1762784779
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1534_
timestamp 1762784779
transform -1 0 3404 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _1535_
timestamp 1762784779
transform 1 0 5152 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1536_
timestamp 1762784779
transform -1 0 2392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1537_
timestamp 1762784779
transform -1 0 3128 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1538_
timestamp 1762784779
transform 1 0 3036 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1539_
timestamp 1762784779
transform -1 0 3772 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1540_
timestamp 1762784779
transform 1 0 3220 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1541_
timestamp 1762784779
transform -1 0 2576 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1762784779
transform 1 0 2760 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1543_
timestamp 1762784779
transform 1 0 3220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1544_
timestamp 1762784779
transform -1 0 4600 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1545_
timestamp 1762784779
transform 1 0 3404 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1546_
timestamp 1762784779
transform -1 0 4968 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1547_
timestamp 1762784779
transform -1 0 4692 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1548_
timestamp 1762784779
transform 1 0 6532 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1549_
timestamp 1762784779
transform -1 0 5336 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1550_
timestamp 1762784779
transform 1 0 4784 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1551_
timestamp 1762784779
transform 1 0 4876 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1552_
timestamp 1762784779
transform -1 0 5152 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1553_
timestamp 1762784779
transform 1 0 5796 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1762784779
transform 1 0 5152 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1555_
timestamp 1762784779
transform 1 0 4876 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1556_
timestamp 1762784779
transform 1 0 3864 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1557_
timestamp 1762784779
transform -1 0 1748 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1558_
timestamp 1762784779
transform -1 0 2116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__a21oi_1  _1559_
timestamp 1762784779
transform -1 0 3128 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1560_
timestamp 1762784779
transform 1 0 2576 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1561_
timestamp 1762784779
transform 1 0 2484 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1562_
timestamp 1762784779
transform -1 0 4968 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1563_
timestamp 1762784779
transform 1 0 3956 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1564_
timestamp 1762784779
transform -1 0 5704 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1565_
timestamp 1762784779
transform -1 0 5244 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1566_
timestamp 1762784779
transform 1 0 3128 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1567_
timestamp 1762784779
transform 1 0 3772 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1568_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3220 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1569_
timestamp 1762784779
transform 1 0 2760 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1570_
timestamp 1762784779
transform 1 0 3588 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1571_
timestamp 1762784779
transform -1 0 3864 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1572_
timestamp 1762784779
transform 1 0 3864 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1573_
timestamp 1762784779
transform 1 0 2024 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1574_
timestamp 1762784779
transform -1 0 2116 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_2  _1575_
timestamp 1762784779
transform -1 0 7360 0 -1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1576_
timestamp 1762784779
transform -1 0 2484 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_1  _1577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 3036 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1578_
timestamp 1762784779
transform -1 0 2576 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1579_
timestamp 1762784779
transform -1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1580_
timestamp 1762784779
transform -1 0 2668 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1581_
timestamp 1762784779
transform 1 0 2300 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1582_
timestamp 1762784779
transform -1 0 4692 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1583_
timestamp 1762784779
transform -1 0 4324 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1584_
timestamp 1762784779
transform 1 0 4324 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1585_
timestamp 1762784779
transform 1 0 4508 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1586_
timestamp 1762784779
transform 1 0 3220 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1587_
timestamp 1762784779
transform 1 0 4508 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1588_
timestamp 1762784779
transform 1 0 3956 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1762784779
transform 1 0 3220 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1590_
timestamp 1762784779
transform 1 0 3864 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1762784779
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1592_
timestamp 1762784779
transform 1 0 2484 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1593_
timestamp 1762784779
transform -1 0 4048 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1594_
timestamp 1762784779
transform 1 0 3220 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1595_
timestamp 1762784779
transform -1 0 1748 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1596_
timestamp 1762784779
transform 1 0 2300 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_4  _1597_
timestamp 1762784779
transform 1 0 920 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__xnor2_1  _1598_
timestamp 1762784779
transform -1 0 7176 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1599_
timestamp 1762784779
transform 1 0 3220 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1600_
timestamp 1762784779
transform 1 0 3220 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1601_
timestamp 1762784779
transform 1 0 3220 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1602_
timestamp 1762784779
transform -1 0 3128 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1603_
timestamp 1762784779
transform -1 0 7268 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1604_
timestamp 1762784779
transform 1 0 4508 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _1605_
timestamp 1762784779
transform -1 0 9292 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1606_
timestamp 1762784779
transform -1 0 9108 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1607_
timestamp 1762784779
transform -1 0 8280 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1608_
timestamp 1762784779
transform 1 0 9752 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1609_
timestamp 1762784779
transform -1 0 9200 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1610_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8740 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1611_
timestamp 1762784779
transform 1 0 8096 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1612_
timestamp 1762784779
transform 1 0 9108 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1613_
timestamp 1762784779
transform 1 0 3496 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1614_
timestamp 1762784779
transform -1 0 9108 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1615_
timestamp 1762784779
transform 1 0 8740 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1616_
timestamp 1762784779
transform -1 0 8280 0 1 37536
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1617_
timestamp 1762784779
transform 1 0 7176 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _1618_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5796 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1619_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 6716 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1620_
timestamp 1762784779
transform -1 0 7636 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1621_
timestamp 1762784779
transform -1 0 7176 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _1622_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6440 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1623_
timestamp 1762784779
transform -1 0 10856 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1624_
timestamp 1762784779
transform 1 0 10396 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _1625_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 11684 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1626_
timestamp 1762784779
transform -1 0 10764 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1627_
timestamp 1762784779
transform 1 0 9752 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1628_
timestamp 1762784779
transform 1 0 9660 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 1762784779
transform -1 0 12144 0 -1 36448
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1630_
timestamp 1762784779
transform 1 0 11500 0 -1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1631_
timestamp 1762784779
transform -1 0 12328 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1632_
timestamp 1762784779
transform 1 0 12052 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1633_
timestamp 1762784779
transform -1 0 12328 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1634_
timestamp 1762784779
transform -1 0 12328 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1635_
timestamp 1762784779
transform -1 0 11500 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1636_
timestamp 1762784779
transform 1 0 10948 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1637_
timestamp 1762784779
transform -1 0 7544 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1638_
timestamp 1762784779
transform -1 0 11500 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1639_
timestamp 1762784779
transform -1 0 11960 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1640_
timestamp 1762784779
transform -1 0 11868 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1641_
timestamp 1762784779
transform 1 0 10396 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1642_
timestamp 1762784779
transform 1 0 11684 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1762784779
transform 1 0 10304 0 -1 42976
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1644_
timestamp 1762784779
transform -1 0 10856 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1645_
timestamp 1762784779
transform 1 0 10396 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1646_
timestamp 1762784779
transform -1 0 10856 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1647_
timestamp 1762784779
transform 1 0 10948 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _1648_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 11500 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1649_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 11592 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1650_
timestamp 1762784779
transform 1 0 9476 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1651_
timestamp 1762784779
transform -1 0 11500 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _1652_
timestamp 1762784779
transform 1 0 9936 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1653_
timestamp 1762784779
transform -1 0 11408 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1654_
timestamp 1762784779
transform 1 0 10212 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1655_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 10948 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1656_
timestamp 1762784779
transform 1 0 6808 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1657_
timestamp 1762784779
transform 1 0 10028 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1658_
timestamp 1762784779
transform 1 0 11408 0 -1 35360
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1659_
timestamp 1762784779
transform -1 0 10028 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1660_
timestamp 1762784779
transform 1 0 9384 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1661_
timestamp 1762784779
transform 1 0 6348 0 1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1662_
timestamp 1762784779
transform -1 0 6624 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1663_
timestamp 1762784779
transform 1 0 7176 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1664_
timestamp 1762784779
transform 1 0 6256 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1665_
timestamp 1762784779
transform 1 0 6624 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1762784779
transform 1 0 6072 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1667_
timestamp 1762784779
transform 1 0 6072 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _1668_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6072 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1669_
timestamp 1762784779
transform -1 0 8280 0 1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1670_
timestamp 1762784779
transform -1 0 7360 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1671_
timestamp 1762784779
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1672_
timestamp 1762784779
transform -1 0 7728 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1673_
timestamp 1762784779
transform 1 0 5796 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1674_
timestamp 1762784779
transform -1 0 3128 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1675_
timestamp 1762784779
transform 1 0 4324 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1676_
timestamp 1762784779
transform 1 0 2484 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1677_
timestamp 1762784779
transform 1 0 5060 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_2  _1678_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 2392 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1679_
timestamp 1762784779
transform -1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1680_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 5704 0 -1 38624
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1681_
timestamp 1762784779
transform -1 0 4600 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1682_
timestamp 1762784779
transform -1 0 1656 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1683_
timestamp 1762784779
transform 1 0 4140 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1684_
timestamp 1762784779
transform 1 0 7544 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1685_
timestamp 1762784779
transform 1 0 828 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1686_
timestamp 1762784779
transform 1 0 3680 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1687_
timestamp 1762784779
transform 1 0 4784 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1688_
timestamp 1762784779
transform -1 0 8924 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1689_
timestamp 1762784779
transform 1 0 3312 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1690_
timestamp 1762784779
transform -1 0 8004 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1691_
timestamp 1762784779
transform 1 0 8372 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1692_
timestamp 1762784779
transform -1 0 5336 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1693_
timestamp 1762784779
transform 1 0 4048 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1694_
timestamp 1762784779
transform 1 0 7728 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1695_
timestamp 1762784779
transform 1 0 4324 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1696_
timestamp 1762784779
transform -1 0 8740 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1697_
timestamp 1762784779
transform -1 0 11500 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1698_
timestamp 1762784779
transform -1 0 12236 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1699_
timestamp 1762784779
transform -1 0 11224 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1700_
timestamp 1762784779
transform -1 0 12144 0 -1 29920
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1701_
timestamp 1762784779
transform -1 0 10856 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1762784779
transform 1 0 11500 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1703_
timestamp 1762784779
transform 1 0 11592 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1704_
timestamp 1762784779
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1705_
timestamp 1762784779
transform 1 0 12052 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1706_
timestamp 1762784779
transform 1 0 11040 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1707_
timestamp 1762784779
transform 1 0 11592 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1708_
timestamp 1762784779
transform 1 0 11960 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1709_
timestamp 1762784779
transform -1 0 11868 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1710_
timestamp 1762784779
transform -1 0 11500 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1711_
timestamp 1762784779
transform -1 0 10856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1712_
timestamp 1762784779
transform -1 0 12052 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1713_
timestamp 1762784779
transform -1 0 11408 0 -1 4896
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1714_
timestamp 1762784779
transform 1 0 10948 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1715_
timestamp 1762784779
transform 1 0 7728 0 -1 1632
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1716_
timestamp 1762784779
transform -1 0 8924 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1717_
timestamp 1762784779
transform 1 0 8648 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1718_
timestamp 1762784779
transform -1 0 7728 0 -1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1719_
timestamp 1762784779
transform -1 0 7728 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1720_
timestamp 1762784779
transform -1 0 7268 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1721_
timestamp 1762784779
transform 1 0 2208 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1722_
timestamp 1762784779
transform 1 0 2576 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1723_
timestamp 1762784779
transform 1 0 2300 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1724_
timestamp 1762784779
transform 1 0 1196 0 -1 3808
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1725_
timestamp 1762784779
transform -1 0 2300 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1726_
timestamp 1762784779
transform -1 0 2116 0 -1 5984
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1727_
timestamp 1762784779
transform -1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1728_
timestamp 1762784779
transform -1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _1729_
timestamp 1762784779
transform -1 0 1472 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1762784779
transform 1 0 1932 0 1 39712
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1731_
timestamp 1762784779
transform -1 0 11960 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1732_
timestamp 1762784779
transform -1 0 10028 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1733_
timestamp 1762784779
transform -1 0 12144 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1734_
timestamp 1762784779
transform 1 0 11960 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1735_
timestamp 1762784779
transform 1 0 7912 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1736_
timestamp 1762784779
transform 1 0 9476 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1737_
timestamp 1762784779
transform 1 0 8832 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1738_
timestamp 1762784779
transform 1 0 8188 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1739_
timestamp 1762784779
transform -1 0 8280 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1740_
timestamp 1762784779
transform 1 0 5152 0 -1 33184
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1741_
timestamp 1762784779
transform 1 0 6348 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _1742_
timestamp 1762784779
transform 1 0 5428 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1743_
timestamp 1762784779
transform 1 0 828 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1744_
timestamp 1762784779
transform 1 0 5244 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1762784779
transform 1 0 4784 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1746_
timestamp 1762784779
transform 1 0 3772 0 -1 34272
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1747_
timestamp 1762784779
transform 1 0 4140 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1748_
timestamp 1762784779
transform -1 0 4600 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1749_
timestamp 1762784779
transform -1 0 3772 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1750_
timestamp 1762784779
transform 1 0 4600 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1751_
timestamp 1762784779
transform 1 0 3220 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1752_
timestamp 1762784779
transform 1 0 4048 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _1753_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1656 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1754_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1656 0 -1 37536
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _1755_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1380 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1756_
timestamp 1762784779
transform 1 0 1380 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1757_
timestamp 1762784779
transform -1 0 3680 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1762784779
transform 1 0 2208 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1762784779
transform 1 0 2668 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1762784779
transform 1 0 4324 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1762784779
transform -1 0 7820 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1762_
timestamp 1762784779
transform -1 0 12328 0 1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1763_
timestamp 1762784779
transform 1 0 10764 0 1 38624
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1762784779
transform -1 0 12328 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1762784779
transform -1 0 12328 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1766_
timestamp 1762784779
transform -1 0 10856 0 -1 41888
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1767_
timestamp 1762784779
transform 1 0 10396 0 1 40800
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1762784779
transform 1 0 9292 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1762784779
transform 1 0 10856 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1770_
timestamp 1762784779
transform -1 0 12328 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1762784779
transform 1 0 9016 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1762784779
transform 1 0 4232 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1773_
timestamp 1762784779
transform 1 0 5796 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1762784779
transform 1 0 5796 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1762784779
transform 1 0 4232 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1762784779
transform 1 0 5336 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1762784779
transform 1 0 3680 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1762784779
transform 1 0 5336 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1762784779
transform 1 0 5060 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1762784779
transform 1 0 3772 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1762784779
transform 1 0 10856 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1762784779
transform -1 0 12328 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1762784779
transform 1 0 10856 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1762784779
transform 1 0 10856 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1762784779
transform 1 0 10856 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1786_
timestamp 1762784779
transform 1 0 10856 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1787_
timestamp 1762784779
transform 1 0 8372 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1788_
timestamp 1762784779
transform 1 0 6808 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1789_
timestamp 1762784779
transform 1 0 1748 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1790_
timestamp 1762784779
transform 1 0 1380 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1791_
timestamp 1762784779
transform 1 0 1104 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1792_
timestamp 1762784779
transform -1 0 2300 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1793_
timestamp 1762784779
transform -1 0 2300 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1794_
timestamp 1762784779
transform 1 0 1288 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1762784779
transform -1 0 2300 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1762784779
transform -1 0 2300 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1762784779
transform -1 0 2300 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1762784779
transform -1 0 2300 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1762784779
transform -1 0 2668 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1762784779
transform 1 0 828 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1762784779
transform 1 0 828 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1762784779
transform 1 0 828 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1762784779
transform -1 0 2300 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1804_
timestamp 1762784779
transform -1 0 2300 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1805_
timestamp 1762784779
transform 1 0 828 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1806_
timestamp 1762784779
transform -1 0 2300 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1807_
timestamp 1762784779
transform -1 0 2300 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1808_
timestamp 1762784779
transform -1 0 2300 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1809_
timestamp 1762784779
transform -1 0 2392 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1810_
timestamp 1762784779
transform -1 0 4692 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1811_
timestamp 1762784779
transform 1 0 828 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1812_
timestamp 1762784779
transform 1 0 828 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1813_
timestamp 1762784779
transform -1 0 2300 0 1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1814_
timestamp 1762784779
transform -1 0 2300 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1815_
timestamp 1762784779
transform -1 0 2300 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1816_
timestamp 1762784779
transform 1 0 1196 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1762784779
transform 1 0 1656 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1818_
timestamp 1762784779
transform 1 0 2024 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1819_
timestamp 1762784779
transform 1 0 2208 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1820_
timestamp 1762784779
transform 1 0 1564 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1821_
timestamp 1762784779
transform 1 0 2300 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1822_
timestamp 1762784779
transform 1 0 2300 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1823_
timestamp 1762784779
transform -1 0 10856 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1824_
timestamp 1762784779
transform 1 0 9016 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1825_
timestamp 1762784779
transform 1 0 10488 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1826_
timestamp 1762784779
transform 1 0 9292 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1827_
timestamp 1762784779
transform -1 0 9844 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1828_
timestamp 1762784779
transform 1 0 5980 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1829_
timestamp 1762784779
transform 1 0 3772 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1830_
timestamp 1762784779
transform 1 0 4232 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1831_
timestamp 1762784779
transform 1 0 3772 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1832_
timestamp 1762784779
transform 1 0 3680 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1833_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 1288 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1834_
timestamp 1762784779
transform -1 0 1288 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1835_
timestamp 1762784779
transform 1 0 2300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1836_
timestamp 1762784779
transform 1 0 3680 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1837_
timestamp 1762784779
transform 1 0 2300 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1838_
timestamp 1762784779
transform -1 0 1288 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1839_
timestamp 1762784779
transform -1 0 1196 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1840_
timestamp 1762784779
transform -1 0 1380 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1841_
timestamp 1762784779
transform -1 0 1196 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1842_
timestamp 1762784779
transform -1 0 1196 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1843_
timestamp 1762784779
transform -1 0 1196 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1844_
timestamp 1762784779
transform 1 0 4600 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1845_
timestamp 1762784779
transform -1 0 1196 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1846_
timestamp 1762784779
transform 1 0 4232 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1847_
timestamp 1762784779
transform -1 0 1288 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1848_
timestamp 1762784779
transform -1 0 1472 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1849_
timestamp 1762784779
transform 1 0 7912 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1850_
timestamp 1762784779
transform -1 0 1656 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1851_
timestamp 1762784779
transform 1 0 7268 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7912 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1762784779
transform -1 0 8096 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1762784779
transform -1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1762784779
transform 1 0 920 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1762784779
transform 1 0 828 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1762784779
transform -1 0 7912 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1762784779
transform 1 0 5888 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1762784779
transform -1 0 5152 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 8280 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1762784779
transform -1 0 3312 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1762784779
transform -1 0 4508 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1762784779
transform -1 0 7636 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1762784779
transform -1 0 3864 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1762784779
transform -1 0 3128 0 1 35360
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1762784779
transform -1 0 5796 0 1 38624
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1762784779
transform 1 0 10488 0 1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1762784779
transform 1 0 9016 0 -1 37536
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_8  clkload0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1472 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 2668 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload2
timestamp 1762784779
transform 1 0 5796 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1380 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1564 0 -1 36448
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_6  clkload5
timestamp 1762784779
transform 1 0 11224 0 -1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload6
timestamp 1762784779
transform 1 0 9476 0 1 37536
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  fanout10 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 7176 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout12
timestamp 1762784779
transform -1 0 7636 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout13 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6440 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 1762784779
transform -1 0 8464 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 1762784779
transform 1 0 11408 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 1762784779
transform 1 0 7728 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout17
timestamp 1762784779
transform -1 0 5796 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout18
timestamp 1762784779
transform -1 0 9384 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout19
timestamp 1762784779
transform 1 0 9660 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout20
timestamp 1762784779
transform -1 0 10948 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 1472 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout22
timestamp 1762784779
transform 1 0 1104 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout23
timestamp 1762784779
transform -1 0 2668 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 1762784779
transform 1 0 8096 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 1762784779
transform -1 0 8188 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 1762784779
transform 1 0 8556 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout27
timestamp 1762784779
transform 1 0 9936 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp 1762784779
transform 1 0 8372 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 1762784779
transform -1 0 4968 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 1762784779
transform -1 0 9568 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout31
timestamp 1762784779
transform -1 0 8096 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout32
timestamp 1762784779
transform 1 0 9752 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp 1762784779
transform -1 0 8740 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout34
timestamp 1762784779
transform 1 0 8740 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 1762784779
transform 1 0 9752 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout36
timestamp 1762784779
transform 1 0 10488 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 1762784779
transform 1 0 5796 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout38
timestamp 1762784779
transform 1 0 3864 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout39
timestamp 1762784779
transform -1 0 3772 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 1762784779
transform -1 0 3680 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 4600 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 1762784779
transform 1 0 828 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 1762784779
transform -1 0 4876 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1762784779
transform 1 0 9936 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1762784779
transform 1 0 8464 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 1762784779
transform -1 0 5428 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1762784779
transform 1 0 5336 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 1762784779
transform 1 0 6532 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout49
timestamp 1762784779
transform -1 0 3588 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout50
timestamp 1762784779
transform -1 0 4784 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 1762784779
transform -1 0 6808 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout52
timestamp 1762784779
transform 1 0 5980 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1762784779
transform 1 0 5428 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 1762784779
transform -1 0 4140 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout55
timestamp 1762784779
transform 1 0 4600 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 1762784779
transform -1 0 3128 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 1762784779
transform 1 0 7544 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout58
timestamp 1762784779
transform 1 0 3772 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout59
timestamp 1762784779
transform 1 0 6072 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1762784779
transform -1 0 8740 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout61 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5428 0 1 33184
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 1762784779
transform 1 0 7728 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout63
timestamp 1762784779
transform -1 0 6808 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout64
timestamp 1762784779
transform -1 0 7268 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout65
timestamp 1762784779
transform -1 0 7912 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 1762784779
transform 1 0 8556 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout67
timestamp 1762784779
transform -1 0 6348 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout68
timestamp 1762784779
transform -1 0 12328 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1762784779
transform 1 0 11960 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout70
timestamp 1762784779
transform -1 0 11684 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout71
timestamp 1762784779
transform 1 0 8464 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1762784779
transform -1 0 10488 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1762784779
transform 1 0 10120 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout74
timestamp 1762784779
transform -1 0 9384 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1762784779
transform 1 0 3772 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1762784779
transform 1 0 8188 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout77
timestamp 1762784779
transform 1 0 7728 0 -1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout78
timestamp 1762784779
transform 1 0 9384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout79
timestamp 1762784779
transform -1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout80
timestamp 1762784779
transform -1 0 10764 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 1762784779
transform 1 0 10212 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout82
timestamp 1762784779
transform -1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 1762784779
transform -1 0 12236 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 1762784779
transform -1 0 12144 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 1762784779
transform 1 0 11592 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout86
timestamp 1762784779
transform -1 0 12052 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 1762784779
transform 1 0 11960 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout88
timestamp 1762784779
transform -1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout89
timestamp 1762784779
transform -1 0 11868 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout90
timestamp 1762784779
transform 1 0 10948 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout91
timestamp 1762784779
transform 1 0 6532 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout92
timestamp 1762784779
transform 1 0 7176 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout93
timestamp 1762784779
transform 1 0 3772 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout94
timestamp 1762784779
transform 1 0 4140 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout95
timestamp 1762784779
transform 1 0 1196 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout96
timestamp 1762784779
transform -1 0 5704 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout97
timestamp 1762784779
transform 1 0 11960 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout98
timestamp 1762784779
transform 1 0 9108 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout99
timestamp 1762784779
transform 1 0 11960 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout100
timestamp 1762784779
transform 1 0 10304 0 1 41888
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1762784779
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40
timestamp 1762784779
transform 1 0 4232 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5336 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 5796 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63
timestamp 1762784779
transform 1 0 6348 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1762784779
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1762784779
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 8372 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_93
timestamp 1762784779
transform 1 0 9108 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99
timestamp 1762784779
transform 1 0 9660 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1762784779
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1762784779
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1762784779
transform 1 0 12052 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp 1762784779
transform 1 0 828 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 1564 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1762784779
transform 1 0 3220 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_52
timestamp 1762784779
transform 1 0 5336 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1762784779
transform 1 0 6348 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1762784779
transform 1 0 7176 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1762784779
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_125
timestamp 1762784779
transform 1 0 12052 0 -1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1762784779
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_15
timestamp 1762784779
transform 1 0 1932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1762784779
transform 1 0 2944 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1762784779
transform 1 0 4140 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_117
timestamp 1762784779
transform 1 0 11316 0 1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_125
timestamp 1762784779
transform 1 0 12052 0 1 1632
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1762784779
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1762784779
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_33
timestamp 1762784779
transform 1 0 3588 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_45
timestamp 1762784779
transform 1 0 4692 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1762784779
transform 1 0 5428 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 1762784779
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1762784779
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1762784779
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1762784779
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_125
timestamp 1762784779
transform 1 0 12052 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1762784779
transform 1 0 828 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1762784779
transform 1 0 1564 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1762784779
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_29
timestamp 1762784779
transform 1 0 3220 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_37
timestamp 1762784779
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_44
timestamp 1762784779
transform 1 0 4600 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_56
timestamp 1762784779
transform 1 0 5704 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_64
timestamp 1762784779
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_68
timestamp 1762784779
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1762784779
transform 1 0 7912 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1762784779
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1762784779
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 1762784779
transform 1 0 10580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1762784779
transform 1 0 828 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_25
timestamp 1762784779
transform 1 0 2852 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1762784779
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_57
timestamp 1762784779
transform 1 0 5796 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_65
timestamp 1762784779
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_78
timestamp 1762784779
transform 1 0 7728 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1762784779
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1762784779
transform 1 0 10120 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_125
timestamp 1762784779
transform 1 0 12052 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 828 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1762784779
transform 1 0 2852 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_29
timestamp 1762784779
transform 1 0 3220 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1762784779
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_43
timestamp 1762784779
transform 1 0 4508 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1762784779
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_80
timestamp 1762784779
transform 1 0 7912 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1762784779
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1762784779
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1762784779
transform 1 0 1932 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_23
timestamp 1762784779
transform 1 0 2668 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_32
timestamp 1762784779
transform 1 0 3496 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1762784779
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1762784779
transform 1 0 7728 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp 1762784779
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_101
timestamp 1762784779
transform 1 0 9844 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_127
timestamp 1762784779
transform 1 0 12236 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1762784779
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1762784779
transform 1 0 1932 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1762784779
transform 1 0 3220 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1762784779
transform 1 0 4048 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_48
timestamp 1762784779
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_61
timestamp 1762784779
transform 1 0 6164 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1762784779
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_96
timestamp 1762784779
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_108
timestamp 1762784779
transform 1 0 10488 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1762784779
transform 1 0 11040 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_123
timestamp 1762784779
transform 1 0 11868 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_127
timestamp 1762784779
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1762784779
transform 1 0 828 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1762784779
transform 1 0 1564 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_35
timestamp 1762784779
transform 1 0 3772 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1762784779
transform 1 0 4876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1762784779
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1762784779
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1762784779
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1762784779
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1762784779
transform 1 0 9752 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_107
timestamp 1762784779
transform 1 0 10396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1762784779
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1762784779
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_125
timestamp 1762784779
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp 1762784779
transform 1 0 2576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_36
timestamp 1762784779
transform 1 0 3864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_48
timestamp 1762784779
transform 1 0 4968 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_54
timestamp 1762784779
transform 1 0 5520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_58
timestamp 1762784779
transform 1 0 5888 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1762784779
transform 1 0 7452 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1762784779
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1762784779
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_113
timestamp 1762784779
transform 1 0 10948 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_125
timestamp 1762784779
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1762784779
transform 1 0 828 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_20
timestamp 1762784779
transform 1 0 2392 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_24
timestamp 1762784779
transform 1 0 2760 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_28
timestamp 1762784779
transform 1 0 3128 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_61
timestamp 1762784779
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_83
timestamp 1762784779
transform 1 0 8188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1762784779
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_97
timestamp 1762784779
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_120
timestamp 1762784779
transform 1 0 11592 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1762784779
transform 1 0 2852 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1762784779
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_41
timestamp 1762784779
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1762784779
transform 1 0 5152 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_58
timestamp 1762784779
transform 1 0 5888 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_62
timestamp 1762784779
transform 1 0 6256 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_74
timestamp 1762784779
transform 1 0 7360 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_96
timestamp 1762784779
transform 1 0 9384 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_108
timestamp 1762784779
transform 1 0 10488 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 1762784779
transform 1 0 2668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_49
timestamp 1762784779
transform 1 0 5060 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1762784779
transform 1 0 6256 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_68
timestamp 1762784779
transform 1 0 6808 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_75
timestamp 1762784779
transform 1 0 7452 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1762784779
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1762784779
transform 1 0 10488 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1762784779
transform 1 0 12236 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1762784779
transform 1 0 828 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_43
timestamp 1762784779
transform 1 0 4508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_68
timestamp 1762784779
transform 1 0 6808 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_74
timestamp 1762784779
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_79
timestamp 1762784779
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1762784779
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1762784779
transform 1 0 8372 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1762784779
transform 1 0 8924 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_98
timestamp 1762784779
transform 1 0 9568 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1762784779
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_125
timestamp 1762784779
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1762784779
transform 1 0 828 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_48
timestamp 1762784779
transform 1 0 4968 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_52
timestamp 1762784779
transform 1 0 5336 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_63
timestamp 1762784779
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_90
timestamp 1762784779
transform 1 0 8832 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1762784779
transform 1 0 9660 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1762784779
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1762784779
transform 1 0 828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1762784779
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_42
timestamp 1762784779
transform 1 0 4416 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1762784779
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1762784779
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_110
timestamp 1762784779
transform 1 0 10672 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1762784779
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_103
timestamp 1762784779
transform 1 0 10028 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1762784779
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_116
timestamp 1762784779
transform 1 0 11224 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_127
timestamp 1762784779
transform 1 0 12236 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1762784779
transform 1 0 828 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_17
timestamp 1762784779
transform 1 0 2116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_21
timestamp 1762784779
transform 1 0 2484 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 1762784779
transform 1 0 3220 0 1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_44
timestamp 1762784779
transform 1 0 4600 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_56
timestamp 1762784779
transform 1 0 5704 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_78
timestamp 1762784779
transform 1 0 7728 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1762784779
transform 1 0 8372 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_95
timestamp 1762784779
transform 1 0 9292 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_105
timestamp 1762784779
transform 1 0 10212 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_109
timestamp 1762784779
transform 1 0 10580 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123
timestamp 1762784779
transform 1 0 11868 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1762784779
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_23
timestamp 1762784779
transform 1 0 2668 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1762784779
transform 1 0 3772 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1762784779
transform 1 0 5428 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_64
timestamp 1762784779
transform 1 0 6440 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_71
timestamp 1762784779
transform 1 0 7084 0 -1 11424
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_82
timestamp 1762784779
transform 1 0 8096 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1762784779
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1762784779
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_120
timestamp 1762784779
transform 1 0 11592 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1762784779
transform 1 0 828 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1762784779
transform 1 0 2760 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_29
timestamp 1762784779
transform 1 0 3220 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_49
timestamp 1762784779
transform 1 0 5060 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1762784779
transform 1 0 5888 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_76
timestamp 1762784779
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1762784779
transform 1 0 8188 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_92
timestamp 1762784779
transform 1 0 9016 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_104
timestamp 1762784779
transform 1 0 10120 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_123
timestamp 1762784779
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_127
timestamp 1762784779
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1762784779
transform 1 0 828 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_8
timestamp 1762784779
transform 1 0 1288 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_21
timestamp 1762784779
transform 1 0 2484 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1762784779
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1762784779
transform 1 0 10488 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_127
timestamp 1762784779
transform 1 0 12236 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_15
timestamp 1762784779
transform 1 0 1932 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1762784779
transform 1 0 2852 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_29
timestamp 1762784779
transform 1 0 3220 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_37
timestamp 1762784779
transform 1 0 3956 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1762784779
transform 1 0 4876 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_69
timestamp 1762784779
transform 1 0 6900 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_104
timestamp 1762784779
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_116
timestamp 1762784779
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_125
timestamp 1762784779
transform 1 0 12052 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_26
timestamp 1762784779
transform 1 0 2944 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_32
timestamp 1762784779
transform 1 0 3496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_40
timestamp 1762784779
transform 1 0 4232 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1762784779
transform 1 0 4876 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1762784779
transform 1 0 5612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_57
timestamp 1762784779
transform 1 0 5796 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_63
timestamp 1762784779
transform 1 0 6348 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_70
timestamp 1762784779
transform 1 0 6992 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_82
timestamp 1762784779
transform 1 0 8096 0 -1 13600
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_94
timestamp 1762784779
transform 1 0 9200 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_106
timestamp 1762784779
transform 1 0 10304 0 -1 13600
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_116
timestamp 1762784779
transform 1 0 11224 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1762784779
transform 1 0 828 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1762784779
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1762784779
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1762784779
transform 1 0 4324 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_49
timestamp 1762784779
transform 1 0 5060 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_55
timestamp 1762784779
transform 1 0 5612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1762784779
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_69
timestamp 1762784779
transform 1 0 6900 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_81
timestamp 1762784779
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1762784779
transform 1 0 8372 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_97
timestamp 1762784779
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_105
timestamp 1762784779
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_126
timestamp 1762784779
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_34
timestamp 1762784779
transform 1 0 3680 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_44
timestamp 1762784779
transform 1 0 4600 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1762784779
transform 1 0 5520 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_71
timestamp 1762784779
transform 1 0 7084 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1762784779
transform 1 0 9384 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1762784779
transform 1 0 10672 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_126
timestamp 1762784779
transform 1 0 12144 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_19
timestamp 1762784779
transform 1 0 2300 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1762784779
transform 1 0 3036 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_33
timestamp 1762784779
transform 1 0 3588 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_44
timestamp 1762784779
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_50
timestamp 1762784779
transform 1 0 5152 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1762784779
transform 1 0 5796 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_66
timestamp 1762784779
transform 1 0 6624 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_70
timestamp 1762784779
transform 1 0 6992 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1762784779
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_126
timestamp 1762784779
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1762784779
transform 1 0 828 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_25
timestamp 1762784779
transform 1 0 2852 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_31
timestamp 1762784779
transform 1 0 3404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_41
timestamp 1762784779
transform 1 0 4324 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_47
timestamp 1762784779
transform 1 0 4876 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1762784779
transform 1 0 5244 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1762784779
transform 1 0 5612 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1762784779
transform 1 0 5796 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_65
timestamp 1762784779
transform 1 0 6532 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_71
timestamp 1762784779
transform 1 0 7084 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1762784779
transform 1 0 2300 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1762784779
transform 1 0 2944 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1762784779
transform 1 0 3220 0 1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1762784779
transform 1 0 4324 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_53
timestamp 1762784779
transform 1 0 5428 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1762784779
transform 1 0 6256 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1762784779
transform 1 0 8096 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_107
timestamp 1762784779
transform 1 0 10396 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_115
timestamp 1762784779
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1762784779
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1762784779
transform 1 0 828 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_16
timestamp 1762784779
transform 1 0 2024 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_28
timestamp 1762784779
transform 1 0 3128 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_34
timestamp 1762784779
transform 1 0 3680 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_44
timestamp 1762784779
transform 1 0 4600 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1762784779
transform 1 0 5796 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1762784779
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_86
timestamp 1762784779
transform 1 0 8464 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_93
timestamp 1762784779
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1762784779
transform 1 0 10764 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1762784779
transform 1 0 10948 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1762784779
transform 1 0 11500 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1762784779
transform 1 0 12144 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1762784779
transform 1 0 828 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_16
timestamp 1762784779
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1762784779
transform 1 0 2944 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1762784779
transform 1 0 3220 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1762784779
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_42
timestamp 1762784779
transform 1 0 4416 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_72
timestamp 1762784779
transform 1 0 7176 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_94
timestamp 1762784779
transform 1 0 9200 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_108
timestamp 1762784779
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_126
timestamp 1762784779
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_46
timestamp 1762784779
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1762784779
transform 1 0 5428 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_126
timestamp 1762784779
transform 1 0 12144 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_25
timestamp 1762784779
transform 1 0 2852 0 1 17952
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_43
timestamp 1762784779
transform 1 0 4508 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_55
timestamp 1762784779
transform 1 0 5612 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_63
timestamp 1762784779
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1762784779
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1762784779
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_92
timestamp 1762784779
transform 1 0 9016 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_97
timestamp 1762784779
transform 1 0 9476 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_105
timestamp 1762784779
transform 1 0 10212 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_109
timestamp 1762784779
transform 1 0 10580 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_117
timestamp 1762784779
transform 1 0 11316 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_125
timestamp 1762784779
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1762784779
transform 1 0 828 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_32
timestamp 1762784779
transform 1 0 3496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_36
timestamp 1762784779
transform 1 0 3864 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_33_91
timestamp 1762784779
transform 1 0 8924 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1762784779
transform 1 0 10672 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1762784779
transform 1 0 10948 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1762784779
transform 1 0 11316 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_3
timestamp 1762784779
transform 1 0 828 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_15
timestamp 1762784779
transform 1 0 1932 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_22
timestamp 1762784779
transform 1 0 2576 0 1 19040
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1762784779
transform 1 0 3220 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1762784779
transform 1 0 4324 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_53
timestamp 1762784779
transform 1 0 5428 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_94
timestamp 1762784779
transform 1 0 9200 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_98
timestamp 1762784779
transform 1 0 9568 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_113
timestamp 1762784779
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_127
timestamp 1762784779
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_3
timestamp 1762784779
transform 1 0 828 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_10
timestamp 1762784779
transform 1 0 1472 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_14
timestamp 1762784779
transform 1 0 1840 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_53
timestamp 1762784779
transform 1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_63
timestamp 1762784779
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_125
timestamp 1762784779
transform 1 0 12052 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_15
timestamp 1762784779
transform 1 0 1932 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_25
timestamp 1762784779
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_36_35
timestamp 1762784779
transform 1 0 3772 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_48
timestamp 1762784779
transform 1 0 4968 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_54
timestamp 1762784779
transform 1 0 5520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_69
timestamp 1762784779
transform 1 0 6900 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_82
timestamp 1762784779
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_107
timestamp 1762784779
transform 1 0 10396 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_124
timestamp 1762784779
transform 1 0 11960 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_19
timestamp 1762784779
transform 1 0 2300 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_37
timestamp 1762784779
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_47
timestamp 1762784779
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1762784779
transform 1 0 5612 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_61
timestamp 1762784779
transform 1 0 6164 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_70
timestamp 1762784779
transform 1 0 6992 0 -1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_79
timestamp 1762784779
transform 1 0 7820 0 -1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_91
timestamp 1762784779
transform 1 0 8924 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_103
timestamp 1762784779
transform 1 0 10028 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1762784779
transform 1 0 10764 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1762784779
transform 1 0 10948 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_121
timestamp 1762784779
transform 1 0 11684 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1762784779
transform 1 0 12236 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_3
timestamp 1762784779
transform 1 0 828 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_19
timestamp 1762784779
transform 1 0 2300 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_26
timestamp 1762784779
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_47
timestamp 1762784779
transform 1 0 4876 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_51
timestamp 1762784779
transform 1 0 5244 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_61
timestamp 1762784779
transform 1 0 6164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_69
timestamp 1762784779
transform 1 0 6900 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_75
timestamp 1762784779
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_92
timestamp 1762784779
transform 1 0 9016 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_98
timestamp 1762784779
transform 1 0 9568 0 1 21216
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_107
timestamp 1762784779
transform 1 0 10396 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_119
timestamp 1762784779
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_126
timestamp 1762784779
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_3
timestamp 1762784779
transform 1 0 828 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_6
timestamp 1762784779
transform 1 0 1104 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_48
timestamp 1762784779
transform 1 0 4968 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1762784779
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_87
timestamp 1762784779
transform 1 0 8556 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_96
timestamp 1762784779
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_127
timestamp 1762784779
transform 1 0 12236 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1762784779
transform 1 0 828 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_20
timestamp 1762784779
transform 1 0 2392 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_49
timestamp 1762784779
transform 1 0 5060 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_58
timestamp 1762784779
transform 1 0 5888 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_106
timestamp 1762784779
transform 1 0 10304 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_66
timestamp 1762784779
transform 1 0 6624 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_99
timestamp 1762784779
transform 1 0 9660 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_106
timestamp 1762784779
transform 1 0 10304 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_42_3
timestamp 1762784779
transform 1 0 828 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_45
timestamp 1762784779
transform 1 0 4692 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_78
timestamp 1762784779
transform 1 0 7728 0 1 23392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1762784779
transform 1 0 8372 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1762784779
transform 1 0 9476 0 1 23392
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_106
timestamp 1762784779
transform 1 0 10304 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_118
timestamp 1762784779
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_40
timestamp 1762784779
transform 1 0 4232 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_89
timestamp 1762784779
transform 1 0 8740 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_43_96
timestamp 1762784779
transform 1 0 9384 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1762784779
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_125
timestamp 1762784779
transform 1 0 12052 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1762784779
transform 1 0 828 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_23
timestamp 1762784779
transform 1 0 2668 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1762784779
transform 1 0 3036 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_38
timestamp 1762784779
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_88
timestamp 1762784779
transform 1 0 8648 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_119
timestamp 1762784779
transform 1 0 11500 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_27
timestamp 1762784779
transform 1 0 3036 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_33
timestamp 1762784779
transform 1 0 3588 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_45
timestamp 1762784779
transform 1 0 4692 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1762784779
transform 1 0 5244 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1762784779
transform 1 0 5612 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1762784779
transform 1 0 5796 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_65
timestamp 1762784779
transform 1 0 6532 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_92
timestamp 1762784779
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1762784779
transform 1 0 10764 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_127
timestamp 1762784779
transform 1 0 12236 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1762784779
transform 1 0 828 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_17
timestamp 1762784779
transform 1 0 2116 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_29
timestamp 1762784779
transform 1 0 3220 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_46_38
timestamp 1762784779
transform 1 0 4048 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_47
timestamp 1762784779
transform 1 0 4876 0 1 25568
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1762784779
transform 1 0 7176 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1762784779
transform 1 0 8372 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_90
timestamp 1762784779
transform 1 0 8832 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_94
timestamp 1762784779
transform 1 0 9200 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_98
timestamp 1762784779
transform 1 0 9568 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_104
timestamp 1762784779
transform 1 0 10120 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_113
timestamp 1762784779
transform 1 0 10948 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_118
timestamp 1762784779
transform 1 0 11408 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_127
timestamp 1762784779
transform 1 0 12236 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_19
timestamp 1762784779
transform 1 0 2300 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_28
timestamp 1762784779
transform 1 0 3128 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_36
timestamp 1762784779
transform 1 0 3864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_44
timestamp 1762784779
transform 1 0 4600 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1762784779
transform 1 0 5796 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_81
timestamp 1762784779
transform 1 0 8004 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_99
timestamp 1762784779
transform 1 0 9660 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1762784779
transform 1 0 10764 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1762784779
transform 1 0 10948 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_125
timestamp 1762784779
transform 1 0 12052 0 -1 26656
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1762784779
transform 1 0 1932 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1762784779
transform 1 0 3036 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_29
timestamp 1762784779
transform 1 0 3220 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_37
timestamp 1762784779
transform 1 0 3956 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_50
timestamp 1762784779
transform 1 0 5152 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_56
timestamp 1762784779
transform 1 0 5704 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_68
timestamp 1762784779
transform 1 0 6808 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_48_106
timestamp 1762784779
transform 1 0 10304 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_112
timestamp 1762784779
transform 1 0 10856 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_117
timestamp 1762784779
transform 1 0 11316 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_125
timestamp 1762784779
transform 1 0 12052 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1762784779
transform 1 0 828 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_35
timestamp 1762784779
transform 1 0 3772 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_46
timestamp 1762784779
transform 1 0 4784 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_54
timestamp 1762784779
transform 1 0 5520 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1762784779
transform 1 0 5796 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_63
timestamp 1762784779
transform 1 0 6348 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_67
timestamp 1762784779
transform 1 0 6716 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_71
timestamp 1762784779
transform 1 0 7084 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_91
timestamp 1762784779
transform 1 0 8924 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_126
timestamp 1762784779
transform 1 0 12144 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_19
timestamp 1762784779
transform 1 0 2300 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_29
timestamp 1762784779
transform 1 0 3220 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_38
timestamp 1762784779
transform 1 0 4048 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1762784779
transform 1 0 8188 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_37
timestamp 1762784779
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_57
timestamp 1762784779
transform 1 0 5796 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_74
timestamp 1762784779
transform 1 0 7360 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_106
timestamp 1762784779
transform 1 0 10304 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1762784779
transform 1 0 828 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_17
timestamp 1762784779
transform 1 0 2116 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_29
timestamp 1762784779
transform 1 0 3220 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_35
timestamp 1762784779
transform 1 0 3772 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_41
timestamp 1762784779
transform 1 0 4324 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_61
timestamp 1762784779
transform 1 0 6164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_80
timestamp 1762784779
transform 1 0 7912 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_126
timestamp 1762784779
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_3
timestamp 1762784779
transform 1 0 828 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_8
timestamp 1762784779
transform 1 0 1288 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_43
timestamp 1762784779
transform 1 0 4508 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_50
timestamp 1762784779
transform 1 0 5152 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_54
timestamp 1762784779
transform 1 0 5520 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_73
timestamp 1762784779
transform 1 0 7268 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_82
timestamp 1762784779
transform 1 0 8096 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_90
timestamp 1762784779
transform 1 0 8832 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_107
timestamp 1762784779
transform 1 0 10396 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_126
timestamp 1762784779
transform 1 0 12144 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1762784779
transform 1 0 828 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_22
timestamp 1762784779
transform 1 0 2576 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1762784779
transform 1 0 3036 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_56
timestamp 1762784779
transform 1 0 5704 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_68
timestamp 1762784779
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_54_79
timestamp 1762784779
transform 1 0 7820 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1762784779
transform 1 0 8188 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_107
timestamp 1762784779
transform 1 0 10396 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_25
timestamp 1762784779
transform 1 0 2852 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_33
timestamp 1762784779
transform 1 0 3588 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_57
timestamp 1762784779
transform 1 0 5796 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_74
timestamp 1762784779
transform 1 0 7360 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_113
timestamp 1762784779
transform 1 0 10948 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_127
timestamp 1762784779
transform 1 0 12236 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_19
timestamp 1762784779
transform 1 0 2300 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_51
timestamp 1762784779
transform 1 0 5244 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_69
timestamp 1762784779
transform 1 0 6900 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_91
timestamp 1762784779
transform 1 0 8924 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_3
timestamp 1762784779
transform 1 0 828 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_44
timestamp 1762784779
transform 1 0 4600 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1762784779
transform 1 0 5612 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1762784779
transform 1 0 10764 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1762784779
transform 1 0 3036 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_34
timestamp 1762784779
transform 1 0 3680 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_85
timestamp 1762784779
transform 1 0 8372 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1762784779
transform 1 0 5612 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_63
timestamp 1762784779
transform 1 0 6348 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_119
timestamp 1762784779
transform 1 0 11500 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_29
timestamp 1762784779
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_51
timestamp 1762784779
transform 1 0 5244 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_101
timestamp 1762784779
transform 1 0 9844 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_34
timestamp 1762784779
transform 1 0 3680 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1762784779
transform 1 0 5796 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_91
timestamp 1762784779
transform 1 0 8924 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1762784779
transform 1 0 10764 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_3
timestamp 1762784779
transform 1 0 828 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_20
timestamp 1762784779
transform 1 0 2392 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_38
timestamp 1762784779
transform 1 0 4048 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_60
timestamp 1762784779
transform 1 0 6072 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1762784779
transform 1 0 5612 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_94
timestamp 1762784779
transform 1 0 9200 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_110
timestamp 1762784779
transform 1 0 10672 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_5
timestamp 1762784779
transform 1 0 1012 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1762784779
transform 1 0 8188 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_89
timestamp 1762784779
transform 1 0 8740 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_65_39
timestamp 1762784779
transform 1 0 4140 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_94
timestamp 1762784779
transform 1 0 9200 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_103
timestamp 1762784779
transform 1 0 10028 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_126
timestamp 1762784779
transform 1 0 12144 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1762784779
transform 1 0 828 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_67_48
timestamp 1762784779
transform 1 0 4968 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_19
timestamp 1762784779
transform 1 0 2300 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_38
timestamp 1762784779
transform 1 0 4048 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_127
timestamp 1762784779
transform 1 0 12236 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_3
timestamp 1762784779
transform 1 0 828 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_29
timestamp 1762784779
transform 1 0 3220 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_77
timestamp 1762784779
transform 1 0 7636 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_70_99
timestamp 1762784779
transform 1 0 9660 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_70_110
timestamp 1762784779
transform 1 0 10672 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_7
timestamp 1762784779
transform 1 0 1196 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_18
timestamp 1762784779
transform 1 0 2208 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_47
timestamp 1762784779
transform 1 0 4876 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_69
timestamp 1762784779
transform 1 0 6900 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_89
timestamp 1762784779
transform 1 0 8740 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1762784779
transform 1 0 10764 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_91
timestamp 1762784779
transform 1 0 8924 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_106
timestamp 1762784779
transform 1 0 10304 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_3
timestamp 1762784779
transform 1 0 828 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_10
timestamp 1762784779
transform 1 0 1472 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_18
timestamp 1762784779
transform 1 0 2208 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_35
timestamp 1762784779
transform 1 0 3772 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_44
timestamp 1762784779
transform 1 0 4600 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_54
timestamp 1762784779
transform 1 0 5520 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_57
timestamp 1762784779
transform 1 0 5796 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_8
timestamp 1762784779
transform 1 0 1288 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_29
timestamp 1762784779
transform 1 0 3220 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_50
timestamp 1762784779
transform 1 0 5152 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1762784779
transform 1 0 828 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1762784779
transform 1 0 3036 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_29
timestamp 1762784779
transform 1 0 3220 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_85
timestamp 1762784779
transform 1 0 8372 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_23
timestamp 1762784779
transform 1 0 2668 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_29
timestamp 1762784779
transform 1 0 3220 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1762784779
transform 1 0 10764 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_123
timestamp 1762784779
transform 1 0 11868 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 6624 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1762784779
transform -1 0 6624 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1762784779
transform -1 0 9844 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1762784779
transform -1 0 4508 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1762784779
transform -1 0 11684 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1762784779
transform 1 0 7268 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1762784779
transform 1 0 11592 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1762784779
transform 1 0 6808 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1762784779
transform -1 0 7268 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1762784779
transform 1 0 5796 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1762784779
transform -1 0 5704 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1762784779
transform 1 0 3312 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1762784779
transform 1 0 1472 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1762784779
transform 1 0 5980 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1762784779
transform -1 0 6808 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1762784779
transform -1 0 6532 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1762784779
transform -1 0 4876 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1762784779
transform -1 0 6532 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1762784779
transform 1 0 4876 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1762784779
transform 1 0 4140 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1762784779
transform -1 0 6348 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform -1 0 6072 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1762784779
transform -1 0 3128 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1762784779
transform -1 0 8188 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1762784779
transform -1 0 10304 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1762784779
transform -1 0 3772 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1762784779
transform -1 0 5336 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1762784779
transform -1 0 3680 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1762784779
transform -1 0 10304 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1762784779
transform 1 0 4508 0 -1 42976
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  max_cap11
timestamp 1762784779
transform 1 0 8372 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_78
timestamp 1762784779
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1762784779
transform -1 0 12604 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_79
timestamp 1762784779
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1762784779
transform -1 0 12604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_80
timestamp 1762784779
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1762784779
transform -1 0 12604 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_81
timestamp 1762784779
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1762784779
transform -1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_82
timestamp 1762784779
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1762784779
transform -1 0 12604 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_83
timestamp 1762784779
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1762784779
transform -1 0 12604 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_84
timestamp 1762784779
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1762784779
transform -1 0 12604 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_85
timestamp 1762784779
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1762784779
transform -1 0 12604 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_86
timestamp 1762784779
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1762784779
transform -1 0 12604 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_87
timestamp 1762784779
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1762784779
transform -1 0 12604 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_88
timestamp 1762784779
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1762784779
transform -1 0 12604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_89
timestamp 1762784779
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1762784779
transform -1 0 12604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_90
timestamp 1762784779
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1762784779
transform -1 0 12604 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_91
timestamp 1762784779
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1762784779
transform -1 0 12604 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_92
timestamp 1762784779
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1762784779
transform -1 0 12604 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_93
timestamp 1762784779
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1762784779
transform -1 0 12604 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_94
timestamp 1762784779
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1762784779
transform -1 0 12604 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_95
timestamp 1762784779
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1762784779
transform -1 0 12604 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_96
timestamp 1762784779
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1762784779
transform -1 0 12604 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_97
timestamp 1762784779
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1762784779
transform -1 0 12604 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_98
timestamp 1762784779
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1762784779
transform -1 0 12604 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_99
timestamp 1762784779
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1762784779
transform -1 0 12604 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_100
timestamp 1762784779
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1762784779
transform -1 0 12604 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_101
timestamp 1762784779
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1762784779
transform -1 0 12604 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_102
timestamp 1762784779
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1762784779
transform -1 0 12604 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_103
timestamp 1762784779
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1762784779
transform -1 0 12604 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_104
timestamp 1762784779
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1762784779
transform -1 0 12604 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_105
timestamp 1762784779
transform 1 0 552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1762784779
transform -1 0 12604 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_106
timestamp 1762784779
transform 1 0 552 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1762784779
transform -1 0 12604 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_107
timestamp 1762784779
transform 1 0 552 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1762784779
transform -1 0 12604 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_108
timestamp 1762784779
transform 1 0 552 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1762784779
transform -1 0 12604 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_109
timestamp 1762784779
transform 1 0 552 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1762784779
transform -1 0 12604 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_110
timestamp 1762784779
transform 1 0 552 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1762784779
transform -1 0 12604 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_111
timestamp 1762784779
transform 1 0 552 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1762784779
transform -1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_112
timestamp 1762784779
transform 1 0 552 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1762784779
transform -1 0 12604 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_113
timestamp 1762784779
transform 1 0 552 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1762784779
transform -1 0 12604 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_114
timestamp 1762784779
transform 1 0 552 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1762784779
transform -1 0 12604 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_115
timestamp 1762784779
transform 1 0 552 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1762784779
transform -1 0 12604 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_116
timestamp 1762784779
transform 1 0 552 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1762784779
transform -1 0 12604 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_117
timestamp 1762784779
transform 1 0 552 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1762784779
transform -1 0 12604 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_118
timestamp 1762784779
transform 1 0 552 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1762784779
transform -1 0 12604 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_119
timestamp 1762784779
transform 1 0 552 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1762784779
transform -1 0 12604 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_120
timestamp 1762784779
transform 1 0 552 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1762784779
transform -1 0 12604 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_121
timestamp 1762784779
transform 1 0 552 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1762784779
transform -1 0 12604 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_122
timestamp 1762784779
transform 1 0 552 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1762784779
transform -1 0 12604 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_123
timestamp 1762784779
transform 1 0 552 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1762784779
transform -1 0 12604 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_124
timestamp 1762784779
transform 1 0 552 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1762784779
transform -1 0 12604 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_125
timestamp 1762784779
transform 1 0 552 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1762784779
transform -1 0 12604 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_126
timestamp 1762784779
transform 1 0 552 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1762784779
transform -1 0 12604 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_127
timestamp 1762784779
transform 1 0 552 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1762784779
transform -1 0 12604 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_128
timestamp 1762784779
transform 1 0 552 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1762784779
transform -1 0 12604 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_129
timestamp 1762784779
transform 1 0 552 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1762784779
transform -1 0 12604 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_130
timestamp 1762784779
transform 1 0 552 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1762784779
transform -1 0 12604 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_131
timestamp 1762784779
transform 1 0 552 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1762784779
transform -1 0 12604 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_132
timestamp 1762784779
transform 1 0 552 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1762784779
transform -1 0 12604 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_133
timestamp 1762784779
transform 1 0 552 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1762784779
transform -1 0 12604 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_134
timestamp 1762784779
transform 1 0 552 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1762784779
transform -1 0 12604 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_135
timestamp 1762784779
transform 1 0 552 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1762784779
transform -1 0 12604 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_136
timestamp 1762784779
transform 1 0 552 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1762784779
transform -1 0 12604 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_137
timestamp 1762784779
transform 1 0 552 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1762784779
transform -1 0 12604 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_138
timestamp 1762784779
transform 1 0 552 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1762784779
transform -1 0 12604 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_139
timestamp 1762784779
transform 1 0 552 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1762784779
transform -1 0 12604 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_140
timestamp 1762784779
transform 1 0 552 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1762784779
transform -1 0 12604 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_141
timestamp 1762784779
transform 1 0 552 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1762784779
transform -1 0 12604 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_142
timestamp 1762784779
transform 1 0 552 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1762784779
transform -1 0 12604 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_143
timestamp 1762784779
transform 1 0 552 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1762784779
transform -1 0 12604 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_144
timestamp 1762784779
transform 1 0 552 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1762784779
transform -1 0 12604 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_145
timestamp 1762784779
transform 1 0 552 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1762784779
transform -1 0 12604 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_146
timestamp 1762784779
transform 1 0 552 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1762784779
transform -1 0 12604 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Left_147
timestamp 1762784779
transform 1 0 552 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_69_Right_69
timestamp 1762784779
transform -1 0 12604 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Left_148
timestamp 1762784779
transform 1 0 552 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_70_Right_70
timestamp 1762784779
transform -1 0 12604 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Left_149
timestamp 1762784779
transform 1 0 552 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_71_Right_71
timestamp 1762784779
transform -1 0 12604 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Left_150
timestamp 1762784779
transform 1 0 552 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_72_Right_72
timestamp 1762784779
transform -1 0 12604 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Left_151
timestamp 1762784779
transform 1 0 552 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_73_Right_73
timestamp 1762784779
transform -1 0 12604 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Left_152
timestamp 1762784779
transform 1 0 552 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_74_Right_74
timestamp 1762784779
transform -1 0 12604 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Left_153
timestamp 1762784779
transform 1 0 552 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_75_Right_75
timestamp 1762784779
transform -1 0 12604 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Left_154
timestamp 1762784779
transform 1 0 552 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_76_Right_76
timestamp 1762784779
transform -1 0 12604 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Left_155
timestamp 1762784779
transform 1 0 552 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_77_Right_77
timestamp 1762784779
transform -1 0 12604 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_156 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1762784779
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_157
timestamp 1762784779
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_158
timestamp 1762784779
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_159
timestamp 1762784779
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 1762784779
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 1762784779
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_162
timestamp 1762784779
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_163
timestamp 1762784779
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_164
timestamp 1762784779
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_165
timestamp 1762784779
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_166
timestamp 1762784779
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_167
timestamp 1762784779
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_168
timestamp 1762784779
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_169
timestamp 1762784779
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_170
timestamp 1762784779
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_171
timestamp 1762784779
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_172
timestamp 1762784779
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_173
timestamp 1762784779
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_174
timestamp 1762784779
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_175
timestamp 1762784779
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_176
timestamp 1762784779
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_177
timestamp 1762784779
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_178
timestamp 1762784779
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_179
timestamp 1762784779
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_180
timestamp 1762784779
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_181
timestamp 1762784779
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_182
timestamp 1762784779
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_183
timestamp 1762784779
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_184
timestamp 1762784779
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_185
timestamp 1762784779
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_186
timestamp 1762784779
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_187
timestamp 1762784779
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_188
timestamp 1762784779
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_189
timestamp 1762784779
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_190
timestamp 1762784779
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_191
timestamp 1762784779
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_192
timestamp 1762784779
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_193
timestamp 1762784779
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_194
timestamp 1762784779
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_195
timestamp 1762784779
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_196
timestamp 1762784779
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_197
timestamp 1762784779
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_198
timestamp 1762784779
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_199
timestamp 1762784779
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_200
timestamp 1762784779
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_201
timestamp 1762784779
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_202
timestamp 1762784779
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_203
timestamp 1762784779
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_204
timestamp 1762784779
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_205
timestamp 1762784779
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_206
timestamp 1762784779
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_207
timestamp 1762784779
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_208
timestamp 1762784779
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_209
timestamp 1762784779
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_210
timestamp 1762784779
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_211
timestamp 1762784779
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_212
timestamp 1762784779
transform 1 0 5704 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_213
timestamp 1762784779
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_214
timestamp 1762784779
transform 1 0 3128 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_215
timestamp 1762784779
transform 1 0 8280 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_216
timestamp 1762784779
transform 1 0 5704 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_217
timestamp 1762784779
transform 1 0 10856 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_218
timestamp 1762784779
transform 1 0 3128 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_219
timestamp 1762784779
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_220
timestamp 1762784779
transform 1 0 5704 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_221
timestamp 1762784779
transform 1 0 10856 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_222
timestamp 1762784779
transform 1 0 3128 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_223
timestamp 1762784779
transform 1 0 8280 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_224
timestamp 1762784779
transform 1 0 5704 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_225
timestamp 1762784779
transform 1 0 10856 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1762784779
transform 1 0 3128 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1762784779
transform 1 0 8280 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1762784779
transform 1 0 5704 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1762784779
transform 1 0 10856 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_230
timestamp 1762784779
transform 1 0 3128 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_231
timestamp 1762784779
transform 1 0 8280 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_232
timestamp 1762784779
transform 1 0 5704 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_233
timestamp 1762784779
transform 1 0 10856 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_234
timestamp 1762784779
transform 1 0 3128 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_235
timestamp 1762784779
transform 1 0 8280 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_236
timestamp 1762784779
transform 1 0 5704 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_237
timestamp 1762784779
transform 1 0 10856 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_238
timestamp 1762784779
transform 1 0 3128 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_239
timestamp 1762784779
transform 1 0 8280 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_240
timestamp 1762784779
transform 1 0 5704 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_241
timestamp 1762784779
transform 1 0 10856 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_242
timestamp 1762784779
transform 1 0 3128 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_243
timestamp 1762784779
transform 1 0 8280 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_244
timestamp 1762784779
transform 1 0 5704 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_245
timestamp 1762784779
transform 1 0 10856 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_246
timestamp 1762784779
transform 1 0 3128 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_247
timestamp 1762784779
transform 1 0 8280 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_248
timestamp 1762784779
transform 1 0 5704 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_249
timestamp 1762784779
transform 1 0 10856 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_250
timestamp 1762784779
transform 1 0 3128 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_251
timestamp 1762784779
transform 1 0 8280 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_252
timestamp 1762784779
transform 1 0 5704 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_253
timestamp 1762784779
transform 1 0 10856 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_254
timestamp 1762784779
transform 1 0 3128 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_255
timestamp 1762784779
transform 1 0 8280 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_256
timestamp 1762784779
transform 1 0 5704 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_257
timestamp 1762784779
transform 1 0 10856 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_258
timestamp 1762784779
transform 1 0 3128 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_259
timestamp 1762784779
transform 1 0 8280 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_260
timestamp 1762784779
transform 1 0 5704 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_261
timestamp 1762784779
transform 1 0 10856 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_262
timestamp 1762784779
transform 1 0 3128 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_263
timestamp 1762784779
transform 1 0 8280 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_264
timestamp 1762784779
transform 1 0 5704 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_265
timestamp 1762784779
transform 1 0 10856 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_266
timestamp 1762784779
transform 1 0 3128 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_267
timestamp 1762784779
transform 1 0 8280 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_268
timestamp 1762784779
transform 1 0 5704 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_269
timestamp 1762784779
transform 1 0 10856 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_270
timestamp 1762784779
transform 1 0 3128 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_271
timestamp 1762784779
transform 1 0 8280 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_272
timestamp 1762784779
transform 1 0 5704 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_273
timestamp 1762784779
transform 1 0 10856 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_274
timestamp 1762784779
transform 1 0 3128 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_275
timestamp 1762784779
transform 1 0 8280 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_276
timestamp 1762784779
transform 1 0 5704 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_277
timestamp 1762784779
transform 1 0 10856 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_278
timestamp 1762784779
transform 1 0 3128 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_279
timestamp 1762784779
transform 1 0 8280 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_280
timestamp 1762784779
transform 1 0 5704 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_281
timestamp 1762784779
transform 1 0 10856 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_282
timestamp 1762784779
transform 1 0 3128 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_283
timestamp 1762784779
transform 1 0 8280 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_284
timestamp 1762784779
transform 1 0 5704 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_285
timestamp 1762784779
transform 1 0 10856 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_286
timestamp 1762784779
transform 1 0 3128 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_287
timestamp 1762784779
transform 1 0 8280 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_288
timestamp 1762784779
transform 1 0 5704 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_289
timestamp 1762784779
transform 1 0 10856 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_290
timestamp 1762784779
transform 1 0 3128 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_291
timestamp 1762784779
transform 1 0 8280 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_292
timestamp 1762784779
transform 1 0 5704 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_293
timestamp 1762784779
transform 1 0 10856 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_294
timestamp 1762784779
transform 1 0 3128 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_295
timestamp 1762784779
transform 1 0 8280 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_296
timestamp 1762784779
transform 1 0 5704 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_69_297
timestamp 1762784779
transform 1 0 10856 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_298
timestamp 1762784779
transform 1 0 3128 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_70_299
timestamp 1762784779
transform 1 0 8280 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_300
timestamp 1762784779
transform 1 0 5704 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_71_301
timestamp 1762784779
transform 1 0 10856 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_302
timestamp 1762784779
transform 1 0 3128 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_72_303
timestamp 1762784779
transform 1 0 8280 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_304
timestamp 1762784779
transform 1 0 5704 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_73_305
timestamp 1762784779
transform 1 0 10856 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_306
timestamp 1762784779
transform 1 0 3128 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_74_307
timestamp 1762784779
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_308
timestamp 1762784779
transform 1 0 5704 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_75_309
timestamp 1762784779
transform 1 0 10856 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_310
timestamp 1762784779
transform 1 0 3128 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_76_311
timestamp 1762784779
transform 1 0 8280 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_312
timestamp 1762784779
transform 1 0 3128 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_313
timestamp 1762784779
transform 1 0 5704 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_314
timestamp 1762784779
transform 1 0 8280 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_77_315
timestamp 1762784779
transform 1 0 10856 0 -1 42976
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 11704 400 11824 0 FreeSans 600 0 0 0 B[0]
port 1 nsew
flabel metal3 s 0 11976 400 12096 0 FreeSans 600 0 0 0 B[1]
port 2 nsew
flabel metal3 s 0 12248 400 12368 0 FreeSans 600 0 0 0 B[2]
port 3 nsew
flabel metal3 s 0 12520 400 12640 0 FreeSans 600 0 0 0 B[3]
port 4 nsew
flabel metal3 s 0 5448 400 5568 0 FreeSans 600 0 0 0 B[4]
port 5 nsew
flabel metal3 s 0 5176 400 5296 0 FreeSans 600 0 0 0 B[5]
port 6 nsew
flabel metal3 s 0 4904 400 5024 0 FreeSans 600 0 0 0 B[6]
port 7 nsew
flabel metal3 s 0 4632 400 4752 0 FreeSans 600 0 0 0 B[7]
port 8 nsew
flabel metal3 s 0 11432 400 11552 0 FreeSans 600 0 0 0 Bbias[0]
port 9 nsew
flabel metal3 s 0 11160 400 11280 0 FreeSans 600 0 0 0 Bbias[1]
port 10 nsew
flabel metal3 s 0 10888 400 11008 0 FreeSans 600 0 0 0 Bbias[2]
port 11 nsew
flabel metal3 s 0 23400 400 23520 0 FreeSans 600 0 0 0 G[0]
port 12 nsew
flabel metal3 s 0 23672 400 23792 0 FreeSans 600 0 0 0 G[1]
port 13 nsew
flabel metal3 s 0 23944 400 24064 0 FreeSans 600 0 0 0 G[2]
port 14 nsew
flabel metal3 s 0 24216 400 24336 0 FreeSans 600 0 0 0 G[3]
port 15 nsew
flabel metal3 s 0 17144 400 17264 0 FreeSans 600 0 0 0 G[4]
port 16 nsew
flabel metal3 s 0 16872 400 16992 0 FreeSans 600 0 0 0 G[5]
port 17 nsew
flabel metal3 s 0 16600 400 16720 0 FreeSans 600 0 0 0 G[6]
port 18 nsew
flabel metal3 s 0 16328 400 16448 0 FreeSans 600 0 0 0 G[7]
port 19 nsew
flabel metal3 s 0 23128 400 23248 0 FreeSans 600 0 0 0 Gbias[0]
port 20 nsew
flabel metal3 s 0 22856 400 22976 0 FreeSans 600 0 0 0 Gbias[1]
port 21 nsew
flabel metal3 s 0 22584 400 22704 0 FreeSans 600 0 0 0 Gbias[2]
port 22 nsew
flabel metal3 s 0 36184 400 36304 0 FreeSans 600 0 0 0 R[0]
port 23 nsew
flabel metal3 s 0 36456 400 36576 0 FreeSans 600 0 0 0 R[1]
port 24 nsew
flabel metal3 s 0 36728 400 36848 0 FreeSans 600 0 0 0 R[2]
port 25 nsew
flabel metal3 s 0 37000 400 37120 0 FreeSans 600 0 0 0 R[3]
port 26 nsew
flabel metal3 s 0 28840 400 28960 0 FreeSans 600 0 0 0 R[4]
port 27 nsew
flabel metal3 s 0 28568 400 28688 0 FreeSans 600 0 0 0 R[5]
port 28 nsew
flabel metal3 s 0 28296 400 28416 0 FreeSans 600 0 0 0 R[6]
port 29 nsew
flabel metal3 s 0 28024 400 28144 0 FreeSans 600 0 0 0 R[7]
port 30 nsew
flabel metal3 s 0 34824 400 34944 0 FreeSans 600 0 0 0 Rbias[0]
port 31 nsew
flabel metal3 s 0 34552 400 34672 0 FreeSans 600 0 0 0 Rbias[1]
port 32 nsew
flabel metal3 s 0 34280 400 34400 0 FreeSans 600 0 0 0 Rbias[2]
port 33 nsew
flabel metal4 s 10716 496 11036 43024 0 FreeSans 2400 90 0 0 VGND
port 34 nsew
flabel metal4 s 4316 496 4636 43024 0 FreeSans 2400 90 0 0 VGND
port 34 nsew
flabel metal4 s 10056 496 10376 43024 0 FreeSans 2400 90 0 0 VPWR
port 35 nsew
flabel metal4 s 3656 496 3976 43024 0 FreeSans 2400 90 0 0 VPWR
port 35 nsew
flabel metal2 s 9402 43500 9458 43900 0 FreeSans 280 90 0 0 clk
port 36 nsew
flabel metal2 s 9954 43500 10010 43900 0 FreeSans 280 90 0 0 ena
port 37 nsew
flabel metal2 s 8850 43500 8906 43900 0 FreeSans 280 90 0 0 rst_n
port 38 nsew
flabel metal2 s 8298 43500 8354 43900 0 FreeSans 280 90 0 0 ui_in[0]
port 39 nsew
flabel metal2 s 7746 43500 7802 43900 0 FreeSans 280 90 0 0 ui_in[1]
port 40 nsew
flabel metal2 s 7194 43500 7250 43900 0 FreeSans 280 90 0 0 ui_in[2]
port 41 nsew
flabel metal2 s 6642 43500 6698 43900 0 FreeSans 280 90 0 0 ui_in[3]
port 42 nsew
flabel metal2 s 6090 43500 6146 43900 0 FreeSans 280 90 0 0 ui_in[4]
port 43 nsew
flabel metal2 s 5538 43500 5594 43900 0 FreeSans 280 90 0 0 ui_in[5]
port 44 nsew
flabel metal2 s 4986 43500 5042 43900 0 FreeSans 280 90 0 0 ui_in[6]
port 45 nsew
flabel metal2 s 4434 43500 4490 43900 0 FreeSans 280 90 0 0 ui_in[7]
port 46 nsew
flabel metal2 s 2778 43500 2834 43900 0 FreeSans 280 90 0 0 uio_in2
port 47 nsew
flabel metal2 s 2226 43500 2282 43900 0 FreeSans 280 90 0 0 uio_in3
port 48 nsew
flabel metal2 s 1674 43500 1730 43900 0 FreeSans 280 90 0 0 uio_in4
port 49 nsew
flabel metal3 s 0 39448 400 39568 0 FreeSans 600 0 0 0 uio_out[0]
port 50 nsew
flabel metal3 s 0 39176 400 39296 0 FreeSans 600 0 0 0 uio_out[1]
port 51 nsew
flabel metal3 s 0 41624 400 41744 0 FreeSans 600 0 0 0 uo_out[0]
port 52 nsew
flabel metal3 s 0 41352 400 41472 0 FreeSans 600 0 0 0 uo_out[1]
port 53 nsew
flabel metal3 s 0 41080 400 41200 0 FreeSans 600 0 0 0 uo_out[2]
port 54 nsew
flabel metal3 s 0 40808 400 40928 0 FreeSans 600 0 0 0 uo_out[3]
port 55 nsew
flabel metal3 s 0 40536 400 40656 0 FreeSans 600 0 0 0 uo_out[4]
port 56 nsew
flabel metal3 s 0 40264 400 40384 0 FreeSans 600 0 0 0 uo_out[5]
port 57 nsew
flabel metal3 s 0 39992 400 40112 0 FreeSans 600 0 0 0 uo_out[6]
port 58 nsew
flabel metal3 s 0 39720 400 39840 0 FreeSans 600 0 0 0 uo_out[7]
port 59 nsew
<< properties >>
string FIXED_BBOX 0 0 12800 43900
string GDS_END 3756988
string GDS_FILE ../gds/controller_wrapper.gds
string GDS_START 666560
<< end >>
