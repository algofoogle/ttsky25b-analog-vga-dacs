magic
tech sky130A
timestamp 1762612625
<< nwell >>
rect 0 -4 86 243
<< pwell >>
rect 86 -4 393 243
<< nmos >>
rect 128 179 178 194
rect 128 135 178 150
rect 128 91 178 106
<< pmos >>
rect 18 177 68 192
rect 18 135 68 150
rect 18 91 68 106
<< mvnmos >>
rect 260 133 310 183
rect 260 58 310 108
<< ndiff >>
rect 128 219 159 221
rect 128 217 178 219
rect 128 200 138 217
rect 155 200 178 217
rect 128 194 178 200
rect 128 173 178 179
rect 128 156 137 173
rect 154 156 178 173
rect 128 150 178 156
rect 128 129 178 135
rect 128 112 136 129
rect 173 112 178 129
rect 128 106 178 112
rect 128 85 178 91
rect 128 68 138 85
rect 155 68 178 85
rect 128 66 178 68
rect 128 32 159 66
<< pdiff >>
rect 18 215 68 219
rect 18 198 37 215
rect 58 198 68 215
rect 18 192 68 198
rect 18 150 68 177
rect 18 129 68 135
rect 18 112 47 129
rect 64 112 68 129
rect 18 106 68 112
rect 18 84 68 91
rect 18 67 22 84
rect 39 67 68 84
rect 18 61 68 67
<< mvndiff >>
rect 260 214 310 218
rect 260 193 268 214
rect 302 193 310 214
rect 260 183 310 193
rect 260 108 310 133
rect 260 48 310 58
rect 260 28 268 48
rect 302 28 310 48
rect 260 23 310 28
<< ndiffc >>
rect 138 200 155 217
rect 137 156 154 173
rect 136 112 173 129
rect 138 68 155 85
<< pdiffc >>
rect 37 198 58 215
rect 47 112 64 129
rect 22 67 39 84
<< mvndiffc >>
rect 268 193 302 214
rect 268 28 302 48
<< psubdiff >>
rect 206 32 223 44
rect 206 2 223 15
<< nsubdiff >>
rect 18 50 68 61
rect 18 33 22 50
rect 39 33 68 50
rect 18 14 68 33
<< psubdiffcont >>
rect 206 15 223 32
<< nsubdiffcont >>
rect 22 33 39 50
<< poly >>
rect 87 204 114 212
rect 87 192 92 204
rect 5 177 18 192
rect 68 187 92 192
rect 109 194 114 204
rect 109 187 128 194
rect 68 179 128 187
rect 178 179 192 194
rect 68 177 114 179
rect 84 151 117 156
rect 84 150 92 151
rect 5 135 18 150
rect 68 135 92 150
rect 84 134 92 135
rect 109 150 117 151
rect 216 173 260 183
rect 109 135 128 150
rect 178 135 192 150
rect 216 143 221 173
rect 241 143 260 173
rect 109 134 117 135
rect 84 129 117 134
rect 216 133 260 143
rect 310 173 354 183
rect 310 143 329 173
rect 349 143 354 173
rect 310 133 354 143
rect 5 91 18 106
rect 68 98 128 106
rect 68 91 92 98
rect 87 81 92 91
rect 109 91 128 98
rect 178 91 192 106
rect 216 98 260 108
rect 109 81 114 91
rect 87 73 114 81
rect 216 68 221 98
rect 241 68 260 98
rect 216 58 260 68
rect 310 98 354 108
rect 310 68 329 98
rect 349 68 354 98
rect 310 58 354 68
<< polycont >>
rect 92 187 109 204
rect 92 134 109 151
rect 221 143 241 173
rect 329 143 349 173
rect 92 81 109 98
rect 221 68 241 98
rect 329 68 349 98
<< locali >>
rect 3 215 66 222
rect 3 198 37 215
rect 58 198 66 215
rect 92 204 109 213
rect 3 92 22 198
rect 128 200 138 217
rect 155 200 196 217
rect 92 178 109 187
rect 92 151 109 159
rect 129 156 137 173
rect 154 156 162 173
rect 39 112 47 129
rect 64 112 73 129
rect 92 126 109 134
rect 179 129 196 200
rect 260 214 310 218
rect 260 193 268 214
rect 302 193 310 214
rect 216 173 246 183
rect 324 173 354 183
rect 216 143 221 173
rect 241 143 329 173
rect 349 143 354 173
rect 216 133 354 143
rect 128 112 136 129
rect 173 112 196 129
rect 3 84 39 92
rect 3 33 22 84
rect 56 55 73 112
rect 92 98 109 107
rect 216 98 354 108
rect 216 85 221 98
rect 92 72 109 81
rect 130 68 138 85
rect 155 68 221 85
rect 241 68 329 98
rect 349 68 354 98
rect 130 67 246 68
rect 130 55 147 67
rect 216 58 246 67
rect 324 58 354 68
rect 56 38 147 55
rect 3 25 39 33
rect 200 32 223 40
rect 200 15 203 32
rect 260 28 268 48
rect 302 28 310 48
rect 200 7 223 15
<< viali >>
rect 92 187 109 204
rect 137 156 154 173
rect 92 134 109 151
rect 268 193 302 214
rect 329 143 349 173
rect 22 50 39 67
rect 92 81 109 98
rect 203 15 206 32
rect 206 15 220 32
rect 268 28 302 48
<< metal1 >>
rect 3 76 28 243
rect 170 214 310 223
rect 89 204 115 213
rect 89 187 92 204
rect 109 187 115 204
rect 89 178 115 187
rect 170 193 268 214
rect 302 193 310 214
rect 170 188 310 193
rect 170 181 208 188
rect 129 173 208 181
rect 42 151 114 160
rect 42 134 92 151
rect 109 134 114 151
rect 129 156 137 173
rect 154 156 208 173
rect 129 147 208 156
rect 42 125 114 134
rect 89 98 118 107
rect 89 81 92 98
rect 109 81 118 98
rect 3 67 42 76
rect 89 72 118 81
rect 3 50 22 67
rect 39 50 42 67
rect 3 41 42 50
rect 3 0 28 41
rect 170 40 208 147
rect 324 173 364 183
rect 324 143 329 173
rect 349 143 364 173
rect 324 133 364 143
rect 260 48 310 51
rect 170 32 223 40
rect 170 15 203 32
rect 220 15 223 32
rect 170 7 223 15
rect 260 28 268 48
rect 302 28 310 48
rect 260 7 310 28
<< labels >>
flabel metal1 178 150 203 175 0 FreeSans 64 0 0 0 VGND
port 4 nsew
flabel metal1 265 12 305 46 0 FreeSans 64 0 0 0 Iout
port 5 nsew
flabel metal1 329 138 359 178 0 FreeSans 80 0 0 0 Vbias
port 1 nsew
flabel mvndiff 265 113 305 128 0 FreeSans 80 0 0 0 SM
flabel pdiff 26 157 60 171 0 FreeSans 80 0 0 0 PUM
flabel metal1 47 130 72 155 0 FreeSans 64 0 0 0 Cn
port 7 nsew
flabel metal1 92 75 115 104 0 FreeSans 64 0 0 0 Sn
port 11 nsew
flabel metal1 12 46 37 71 0 FreeSans 64 0 0 0 VPWR
port 9 nsew
flabel locali 92 39 122 54 0 FreeSans 80 0 0 0 Ien
flabel metal1 92 181 115 210 0 FreeSans 64 0 0 0 Rn
port 12 nsew
flabel locali 130 201 136 215 0 FreeSans 80 0 0 0 PDM
<< properties >>
string FIXED_BBOX 0 0 393 232
<< end >>
