magic
tech sky130A
magscale 1 2
timestamp 1760337109
<< metal1 >>
rect 7490 11384 7530 11424
rect 7572 11384 7612 11424
rect 9138 11384 9178 11424
rect 9748 11384 9788 11424
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect -1330 10282 -1192 10750
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect -484 10542 -418 10548
rect -484 10488 -478 10542
rect -424 10488 -418 10542
rect -484 10482 -418 10488
rect -824 10448 -760 10454
rect -824 10396 -818 10448
rect -766 10396 -760 10448
rect -824 10390 -760 10396
rect -814 10276 -768 10390
rect -474 10284 -428 10482
rect 684 10282 1268 10796
rect -1470 9996 -1368 10006
rect -1470 9944 -1464 9996
rect -1412 9944 -1368 9996
rect -1470 9936 -1368 9944
rect 1434 9478 3158 9514
rect 1434 9432 1470 9478
rect 3664 9450 3700 9536
rect 4208 9472 4244 9542
rect 1312 9396 1470 9432
rect 1870 9414 3700 9450
rect 3814 9436 4244 9472
rect 4644 9500 4728 9536
rect 1312 9318 1348 9396
rect 1084 9282 1348 9318
rect 1084 9162 1120 9282
rect 1870 9162 1906 9414
rect 3814 9386 3850 9436
rect 4644 9406 4680 9500
rect 5292 9462 5328 9542
rect 5786 9464 5822 9542
rect 2656 9350 3850 9386
rect 3884 9370 4680 9406
rect 4750 9426 5328 9462
rect 5574 9428 5822 9464
rect 2656 9162 2692 9350
rect 3884 9322 3920 9370
rect 4750 9342 4786 9426
rect 5574 9398 5610 9428
rect 6382 9400 6418 9542
rect 6876 9464 6912 9542
rect 3442 9286 3920 9322
rect 4228 9306 4786 9342
rect 5014 9362 5610 9398
rect 5800 9364 6418 9400
rect 6586 9428 6912 9464
rect 3442 9162 3478 9286
rect 4228 9162 4264 9306
rect 5014 9162 5050 9362
rect 5800 9162 5836 9364
rect 6586 9162 6622 9428
rect 7392 9394 7428 9544
rect 7372 9358 7428 9394
rect 7372 9162 7408 9358
rect 8158 9162 8194 9542
rect 8594 9494 8630 9534
rect 8594 9458 8980 9494
rect 8944 9162 8980 9458
rect 9306 9360 9342 9544
rect 9678 9482 9714 9542
rect 9678 9446 10026 9482
rect 9990 9392 10026 9446
rect 10412 9460 10448 9542
rect 10764 9486 10800 9544
rect 10412 9424 10692 9460
rect 10764 9450 12124 9486
rect 10656 9398 10692 9424
rect 9306 9324 9766 9360
rect 9990 9356 10552 9392
rect 10656 9362 11338 9398
rect 9730 9162 9766 9324
rect 10516 9162 10552 9356
rect 11302 9162 11338 9362
rect 12088 9162 12124 9450
rect -2130 4230 -2090 4270
rect -2130 4148 -2090 4188
rect -2130 2582 -2090 2622
rect -2130 1972 -2090 2012
<< via1 >>
rect -1320 10750 -1202 11316
rect 694 10796 1258 11016
rect -478 10488 -424 10542
rect -818 10396 -766 10448
rect -1464 9944 -1412 9996
<< metal2 >>
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect 684 10786 1268 10796
rect -1330 10740 -1192 10750
rect -484 10542 -418 10548
rect -484 10538 -478 10542
rect -2130 10492 -478 10538
rect -484 10488 -478 10492
rect -424 10488 -418 10542
rect -484 10482 -418 10488
rect -824 10448 -760 10454
rect -824 10445 -818 10448
rect -1631 10399 -818 10445
rect -1631 10266 -1585 10399
rect -824 10396 -818 10399
rect -766 10396 -760 10448
rect -824 10390 -760 10396
rect -2130 10220 -1585 10266
rect -1470 9996 -1368 10006
rect -1470 9994 -1464 9996
rect -2130 9948 -1464 9994
rect -1470 9944 -1464 9948
rect -1412 9944 -1368 9996
rect -1470 9936 -1368 9944
rect 808 9198 886 9354
rect 0 9188 906 9198
rect 0 9118 10 9188
rect 896 9118 906 9188
rect 0 9108 906 9118
rect -44 7912 16 7952
rect -44 7448 16 7488
rect -44 6984 16 7024
rect -44 6520 16 6560
rect -44 6056 16 6096
rect -44 5592 16 5632
rect -44 5128 16 5168
rect -44 4664 16 4704
rect -44 4200 16 4240
rect -44 3736 16 3776
rect -44 3272 16 3312
rect -44 2808 16 2848
rect -44 2344 16 2384
rect -44 1880 16 1920
rect -44 1416 16 1456
<< via2 >>
rect -1320 10750 -1202 11316
rect 694 10796 1258 11016
rect 10 9118 896 9188
<< metal3 >>
rect -1330 11316 -1192 11326
rect -1330 10750 -1320 11316
rect -1202 10750 -1192 11316
rect 14268 11320 14508 11326
rect 14268 11092 14274 11320
rect 14502 11092 14508 11320
rect 684 11016 1268 11026
rect 684 10796 694 11016
rect 1258 10796 1268 11016
rect 684 10786 1268 10796
rect -1330 10740 -1192 10750
rect 0 9188 906 9198
rect 0 9118 10 9188
rect 896 9118 906 9188
rect 0 9108 906 9118
rect 14268 8742 14508 11092
rect 14268 8514 14274 8742
rect 14466 8740 14508 8742
rect 14500 8706 14508 8740
rect 14502 8514 14508 8706
rect 14268 8508 14508 8514
rect -1385 1050 -1147 1055
rect -2038 810 -2032 1050
rect -1794 1049 -1146 1050
rect -1794 811 -1385 1049
rect -1147 811 -1146 1049
rect -1794 810 -1146 811
rect -1385 805 -1147 810
<< via3 >>
rect -1320 11096 -1202 11316
rect 14274 11092 14502 11320
rect 694 10796 1258 11016
rect 10 9118 896 9188
rect 14274 8740 14466 8742
rect 14274 8706 14500 8740
rect 14274 8514 14502 8706
rect -2032 810 -1794 1050
rect -1385 811 -1147 1049
<< metal4 >>
rect -2032 11316 3228 11326
rect -2032 11096 -1320 11316
rect -1202 11096 3228 11316
rect -2032 11086 3228 11096
rect 10900 11320 14508 11326
rect 10900 11092 14274 11320
rect 14502 11092 14508 11320
rect 10900 11086 14508 11092
rect -2032 8680 -1792 11086
rect -1732 11016 3212 11026
rect -1732 10796 694 11016
rect 1258 10796 3212 11016
rect -1732 10786 3212 10796
rect 10810 10786 14828 11026
rect -1732 8680 -1492 10786
rect 0 9188 906 9198
rect 0 9118 10 9188
rect 896 9118 906 9188
rect 0 9108 906 9118
rect 14066 9108 14208 9168
rect 14466 8740 14502 8742
rect 14500 8706 14502 8740
rect 14588 8694 14828 10786
rect -2033 1050 -1793 1051
rect -2033 810 -2032 1050
rect -1794 810 -1793 1050
rect -1386 1049 -518 1050
rect -2033 809 -1793 810
rect -1732 700 -1492 950
rect -1386 811 -1385 1049
rect -1147 1000 -518 1049
rect -1147 811 370 1000
rect -1386 810 370 811
rect -758 760 370 810
rect -1732 460 202 700
rect 13022 0 13422 400
use thermo15c  thermo15c_0
timestamp 1760335364
transform 1 0 3900 0 1 16934
box -1016 -7430 7240 -5510
use array255x  XA
timestamp 1759928440
transform 1 0 60 0 1 1046
box -60 -1046 14768 8152
use thermo15  XThR
timestamp 1759723169
transform 1 0 -1114 0 1 8236
box -1016 -7616 1090 640
use vbias  XVB
timestamp 1757954071
transform 1 0 -1412 0 1 9310
box 0 0 2716 1016
<< labels >>
flabel metal4 13022 0 13422 400 0 FreeSans 1600 0 0 0 Iout
port 0 nsew
flabel metal4 -2032 11086 3228 11326 0 FreeSans 1600 0 0 0 VPWR
port 1 nsew
flabel metal4 -1732 10786 3212 11026 0 FreeSans 1600 0 0 0 VGND
port 2 nsew
flabel metal4 14066 9108 14208 9168 0 FreeSans 160 0 0 0 Vbias
port 3 nsew
flabel metal1 -2130 1972 -2090 2012 0 FreeSans 80 0 0 0 data[7]
port 1807 nsew
flabel metal1 -2130 2582 -2090 2622 0 FreeSans 80 0 0 0 data[6]
port 1806 nsew
flabel metal1 -2130 4148 -2090 4188 0 FreeSans 80 0 0 0 data[5]
port 1805 nsew
flabel metal1 -2130 4230 -2090 4270 0 FreeSans 80 0 0 0 data[4]
port 1804 nsew
flabel metal1 9748 11384 9788 11424 0 FreeSans 80 0 0 0 data[3]
port 1803 nsew
flabel metal1 9138 11384 9178 11424 0 FreeSans 80 0 0 0 data[2]
port 1802 nsew
flabel metal1 7572 11384 7612 11424 0 FreeSans 80 0 0 0 data[1]
port 1801 nsew
flabel metal1 7490 11384 7530 11424 0 FreeSans 80 0 0 0 data[0]
port 1800 nsew
flabel metal2 -2130 10492 -2084 10538 0 FreeSans 80 0 0 0 bias[0]
port 1808 nsew
flabel metal2 -2130 10220 -2084 10266 0 FreeSans 80 0 0 0 bias[1]
port 1809 nsew
flabel metal2 -2130 9948 -2084 9994 0 FreeSans 80 0 0 0 bias[2]
port 1810 nsew
<< end >>
