* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 VPWR.t1522 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1521 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1458 VPWR.t1460 VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2 VGND.t1587 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X3 VGND.t928 XThR.XTBN.Y a_n997_2667# VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR.t299 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X5 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t1712 VPWR.t1711 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X6 VGND.t291 Vbias.t6 XA.XIR[9].XIC[7].icell.SM VGND.t290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X7 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t1261 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X8 XThC.Tn[6].t7 XThC.XTBN.Y.t4 VGND.t658 VGND.t657 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X9 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1926 VGND.t1827 VGND.t1826 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X10 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t1128 VGND.t1127 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 VGND.t659 XThC.XTBN.Y.t5 XThC.Tn[5].t3 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t1032 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X13 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t1263 VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 VGND.t191 Vbias.t2 Vbias.t3 VGND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.58 as=0.725 ps=5.58 w=2.5 l=1
X15 VGND.t1276 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 XThC.Tn[12].t7 XThC.XTB5.Y VPWR.t1688 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 VGND.t293 Vbias.t7 XA.XIR[2].XIC[0].icell.SM VGND.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X18 XA.XIR[8].XIC_15.icell.PDM VPWR.t1927 VGND.t1825 VGND.t1824 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X19 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t857 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X20 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t3 VPWR.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1456 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1457 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X22 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t7 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X24 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t813 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 XA.XIR[0].XIC[4].icell.PDM VGND.t2013 VGND.t2015 VGND.t2014 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X26 VGND.t295 Vbias.t8 XA.XIR[0].XIC[13].icell.SM VGND.t294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X27 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t2072 VGND.t2071 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X28 XThR.Tn[5].t3 XThR.XTBN.Y a_n1049_5611# VPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 XThC.Tn[4].t11 XThC.XTB5.Y VGND.t2264 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X30 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t50 VGND.t585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X31 VGND.t2590 XThC.XTBN.Y.t8 XThC.Tn[2].t7 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X32 XThR.XTB2.Y XThR.XTB6.A VPWR.t1861 VPWR.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t576 VGND.t575 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X34 VGND.t1352 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t1351 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X35 VPWR.t1455 VPWR.t1453 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X36 VGND.t1823 VPWR.t1928 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t1822 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X37 VPWR.t1573 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t1572 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X38 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X39 VGND.t689 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VGND.t1821 VPWR.t1929 XA.XIR[10].XIC_15.icell.PDM VGND.t1820 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X41 VPWR.t1915 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X42 VGND.t297 Vbias.t9 XA.XIR[12].XIC[2].icell.SM VGND.t296 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X43 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1450 VPWR.t1452 VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X45 VGND.t299 Vbias.t10 XA.XIR[11].XIC_15.icell.SM VGND.t298 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X46 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t32 VGND.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X47 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t7 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X48 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X49 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t682 VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X50 VGND.t301 Vbias.t11 XA.XIR[15].XIC[3].icell.SM VGND.t300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t11 VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t1338 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t1337 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 VGND.t303 Vbias.t12 XA.XIR[14].XIC[4].icell.SM VGND.t302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X54 XThC.XTB5.Y XThC.XTB7.B VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X55 XThC.Tn[7].t3 XThC.XTBN.Y.t9 VPWR.t1889 VPWR.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X56 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t1130 VGND.t1129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X57 VGND.t2121 XThR.XTB7.Y XThR.Tn[6].t11 VGND.t2120 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X58 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t78 VPWR.t77 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X59 VPWR.t532 XThR.XTBN.Y XThR.Tn[9].t3 VPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X60 XThR.XTB7.Y XThR.XTB7.A VGND.t1064 VGND.t1063 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X61 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t1575 VPWR.t1574 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X62 VGND.t2012 VGND.t2010 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t2011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X63 VPWR.t1577 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t1576 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X64 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t1265 VGND.t1264 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X65 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t1077 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X66 VPWR.t1520 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1519 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t301 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 VPWR.t1449 VPWR.t1447 XA.XIR[2].XIC_15.icell.PUM VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X69 VGND.t305 Vbias.t13 XA.XIR[9].XIC[2].icell.SM VGND.t304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X70 a_6243_9615# XThC.XTB7.Y VPWR.t968 VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X71 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1272 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X72 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X73 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t209 VGND.t208 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 XThR.Tn[7].t3 XThR.XTBN.Y VPWR.t531 VPWR.t530 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X75 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t38 VGND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X76 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t1069 VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 a_8963_9569# XThC.XTBN.Y.t10 VGND.t2591 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X78 VGND.t1232 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t1231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X79 VGND.t1819 VPWR.t1930 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t1818 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X80 VGND.t927 XThR.XTBN.Y XThR.Tn[5].t7 VGND.t910 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X81 VGND.t1219 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t1218 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X82 VGND.t1278 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t1277 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X83 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t208 VGND.t2373 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X84 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t195 VGND.t2351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X85 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t126 VGND.t1190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X86 VGND.t307 Vbias.t14 XA.XIR[8].XIC_15.icell.SM VGND.t306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X87 VGND.t2252 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t2251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X88 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t80 VPWR.t79 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X89 VPWR.t1905 XThR.XTB6.Y a_n1049_5611# VPWR.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X90 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X91 VGND.t309 Vbias.t15 XA.XIR[1].XIC[5].icell.SM VGND.t308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X92 VGND.t1354 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t1353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X93 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1595 VPWR.t1594 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X94 VGND.t311 Vbias.t16 XA.XIR[4].XIC[6].icell.SM VGND.t310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X95 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1931 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t1817 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X96 a_n1049_7787# XThR.XTB2.Y VPWR.t1020 VPWR.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X97 VGND.t1496 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X98 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t565 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X99 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t708 VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X100 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t935 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1445 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1446 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X102 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X103 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t82 VPWR.t81 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X104 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t567 VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X105 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t569 VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t128 VPWR.t127 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X107 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t15 VGND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X108 VGND.t1317 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X109 VPWR.t611 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X110 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t1078 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t1382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X112 VPWR.t614 data[4].t0 a_n1335_4229# VPWR.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X113 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1518 VPWR.t1517 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X114 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t1131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X115 VGND.t926 XThR.XTBN.Y XThR.Tn[7].t7 VGND.t925 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X116 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X117 a_n1319_5317# XThR.XTB7.A VPWR.t691 VPWR.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X118 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X119 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t2050 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X120 VPWR.t642 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t641 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X121 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X122 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X123 XThC.Tn[9].t11 XThC.XTB2.Y VPWR.t1772 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 XA.XIR[15].XIC[4].icell.Ien VPWR.t1442 VPWR.t1444 VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X125 VGND.t2009 VGND.t2007 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t2008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X126 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1439 VPWR.t1441 VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X127 XThC.Tn[5].t2 XThC.XTBN.Y.t11 VGND.t2592 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X128 VGND.t1234 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X129 VPWR.t450 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X130 VGND.t313 Vbias.t17 XA.XIR[4].XIC[10].icell.SM VGND.t312 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X131 VPWR.t870 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t869 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X132 XThR.Tn[9].t7 XThR.XTB2.Y a_n997_3755# VGND.t947 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X133 XThC.Tn[0].t2 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t1890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X134 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1932 VGND.t1816 VGND.t1815 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X135 VGND.t315 Vbias.t18 XA.XIR[11].XIC[8].icell.SM VGND.t314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X136 XThC.Tn[5].t6 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X137 VGND.t2263 XThC.XTB5.Y XThC.Tn[4].t10 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X138 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X139 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t11 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X140 VGND.t317 Vbias.t19 XA.XIR[1].XIC[0].icell.SM VGND.t316 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X141 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t148 VGND.t1335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X142 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X143 XThC.Tn[7].t7 XThC.XTBN.Y.t14 VGND.t2594 VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X144 XThC.Tn[2].t6 XThC.XTBN.Y.t15 VGND.t2595 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X145 VGND.t1585 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t1584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X146 a_n997_1579# XThR.XTBN.Y VGND.t924 VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X147 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t1384 VGND.t1383 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X148 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t1386 VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X149 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1437 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X150 VGND.t319 Vbias.t20 XA.XIR[4].XIC[1].icell.SM VGND.t318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X151 VGND.t1340 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t1339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t133 VGND.t1226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X153 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X154 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X155 VGND.t321 Vbias.t21 XA.XIR[2].XIC[14].icell.SM VGND.t320 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X156 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t578 VGND.t577 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t1080 VGND.t1079 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t2094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X159 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X160 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t221 VGND.t2403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X161 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t760 VGND.t759 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X162 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t1519 VGND.t1518 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X163 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t925 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X164 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t872 VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X165 XA.XIR[15].XIC[0].icell.Ien VPWR.t1434 VPWR.t1436 VPWR.t1435 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X166 VGND.t1478 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t1477 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X167 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1431 VPWR.t1433 VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X168 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X169 VGND.t1144 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t1143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X170 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t1714 VPWR.t1713 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X171 VGND.t2596 XThC.XTBN.Y.t16 XThC.Tn[1].t7 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X172 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t226 VGND.t2409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X173 VPWR.t874 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X174 VGND.t323 Vbias.t22 XA.XIR[5].XIC[7].icell.SM VGND.t322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X175 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t400 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X176 XA.XIR[2].XIC_15.icell.PUM VPWR.t1429 XA.XIR[2].XIC_15.icell.Ien VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X177 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t1873 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X178 VPWR.t759 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t758 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X179 VPWR.t452 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X180 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1933 VGND.t1814 VGND.t1813 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X181 VPWR.t1428 VPWR.t1426 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1427 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VGND.t325 Vbias.t23 XA.XIR[8].XIC[8].icell.SM VGND.t324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X183 VGND.t2006 VGND.t2004 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t2005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X184 VPWR.t1891 XThC.XTBN.Y.t17 XThC.Tn[10].t11 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X185 VGND.t923 XThR.XTBN.Y XThR.Tn[3].t10 VGND.t886 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X186 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t1872 VGND.t1871 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X187 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t303 VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X188 XThR.Tn[0].t5 XThR.XTBN.Y a_n1049_8581# VPWR.t529 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X189 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t1051 VPWR.t1050 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X190 VPWR.t551 VGND.t2688 XA.XIR[0].XIC[8].icell.PUM VPWR.t550 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X191 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t141 VGND.t1301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X192 VGND.t327 Vbias.t24 XA.XIR[11].XIC[3].icell.SM VGND.t326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X193 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t2671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X194 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t2672 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t122 VGND.t1161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X196 XThC.Tn[12].t6 XThC.XTB5.Y VPWR.t1687 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X197 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X198 XThR.Tn[11].t7 XThR.XTBN.Y VPWR.t528 VPWR.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t693 VPWR.t692 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X200 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t22 VGND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X201 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t1870 VGND.t1869 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X203 VGND.t2003 VGND.t2001 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t2002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X204 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t762 VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t1388 VGND.t1387 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 VGND.t1280 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t1279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X207 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X208 XThR.Tn[2].t8 XThR.XTBN.Y VGND.t922 VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X209 VGND.t1282 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t1281 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X210 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t35 VGND.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X211 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t876 VPWR.t875 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X212 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t248 VGND.t2648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X213 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X214 VPWR.t527 XThR.XTBN.Y XThR.Tn[12].t3 VPWR.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X215 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t19 VGND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X216 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t1082 VGND.t1081 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X217 XThC.XTB7.A data[0].t0 VPWR.t283 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X218 VPWR.t761 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t760 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X219 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t401 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t329 Vbias.t25 XA.XIR[15].XIC[12].icell.SM VGND.t328 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X221 VGND.t331 Vbias.t26 XA.XIR[14].XIC[13].icell.SM VGND.t330 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X222 XA.XIR[0].XIC[13].icell.PDM VGND.t1998 VGND.t2000 VGND.t1999 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X223 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t1521 VGND.t1520 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X224 VGND.t1812 VPWR.t1934 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t1811 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X225 VGND.t1356 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X226 XThC.Tn[9].t7 XThC.XTB2.Y a_7875_9569# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X227 VGND.t2684 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t2683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t1917 VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X229 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1935 VGND.t1810 VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X230 VGND.t1358 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t1357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X231 VGND.t691 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t690 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X232 VGND.t1808 VPWR.t1936 XA.XIR[3].XIC_15.icell.PDM VGND.t1807 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X233 a_n1319_5611# XThR.XTB6.A VPWR.t1860 VPWR.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X234 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t1053 VPWR.t1052 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X235 VGND.t921 XThR.XTBN.Y a_n997_3979# VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X236 VPWR.t1892 XThC.XTBN.Y.t18 XThC.Tn[14].t3 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X237 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t81 VGND.t949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X238 VPWR.t878 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X239 VGND.t333 Vbias.t27 XA.XIR[5].XIC[2].icell.SM VGND.t332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X240 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t936 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X241 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X242 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X243 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t124 VGND.t1188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X244 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t232 VGND.t2511 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X245 VGND.t335 Vbias.t28 XA.XIR[8].XIC[3].icell.SM VGND.t334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X246 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t918 VPWR.t917 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X247 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t1868 VGND.t1867 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X248 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t305 VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X249 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t2284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X250 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t710 VPWR.t709 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X251 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t207 VGND.t2372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X252 VGND.t1248 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t1247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X253 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t1390 VGND.t1389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X254 VPWR.t53 XThR.XTB4.Y.t2 a_n1049_6699# VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VGND.t1806 VPWR.t1937 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t1805 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X256 VPWR.t553 VGND.t2689 XA.XIR[0].XIC[3].icell.PUM VPWR.t552 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X257 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t37 VGND.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X258 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t2673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X259 VPWR.t624 XThC.XTB6.Y a_5949_9615# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X260 VPWR.t1913 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t1912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X261 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X262 VPWR.t1597 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t1596 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X263 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t920 VPWR.t919 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X264 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t1132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X265 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t192 VGND.t2342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X266 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t101 VGND.t1009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X267 VGND.t1997 VGND.t1995 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X268 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X269 VGND.t1236 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t1235 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X270 VGND.t738 XThR.XTB7.B a_n1335_8107# VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X271 VPWR.t146 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t145 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X272 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t1312 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X273 VPWR.t1425 VPWR.t1423 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X274 VGND.t1238 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X275 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t148 VPWR.t147 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X276 XThC.XTB4.Y.t0 XThC.XTB7.B VPWR.t111 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X277 VGND.t1221 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t1220 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X278 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t41 VGND.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X279 VPWR.t1422 VPWR.t1420 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1421 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X280 XThR.Tn[2].t10 XThR.XTB3.Y.t3 VGND.t1170 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X281 VGND.t920 XThR.XTBN.Y a_n997_2891# VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X282 VPWR.t763 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t762 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X283 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t20 VGND.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X284 VGND.t337 Vbias.t29 XA.XIR[10].XIC[11].icell.SM VGND.t336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X285 VGND.t1994 VGND.t1992 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1993 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X286 VPWR.t1786 XThR.XTB5.Y XThR.Tn[12].t7 VPWR.t1525 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X287 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t882 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X288 VGND.t1271 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t1270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X289 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t2285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X290 VGND.t919 XThR.XTBN.Y XThR.Tn[6].t7 VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X291 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t2096 VGND.t2095 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X292 VPWR.t526 XThR.XTBN.Y XThR.Tn[9].t2 VPWR.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X293 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t1055 VPWR.t1054 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X294 XA.XIR[14].XIC_15.icell.PUM VPWR.t1418 XA.XIR[14].XIC_15.icell.Ien VPWR.t1419 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X295 VGND.t355 Vbias.t30 XA.XIR[1].XIC[14].icell.SM VGND.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X296 a_n997_715# XThR.XTBN.Y VGND.t917 VGND.t916 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t2674 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X298 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t2530 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X299 XThC.Tn[1].t6 XThC.XTBN.Y.t19 VGND.t2597 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X300 VPWR.t1599 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t1598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X301 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t28 VGND.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t937 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X303 XThR.Tn[14].t11 XThR.XTB7.Y VPWR.t1621 VPWR.t1620 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X304 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X305 XA.XIR[7].XIC_15.icell.PDM VPWR.t1938 VGND.t1804 VGND.t1803 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X306 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t85 VGND.t955 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X307 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t858 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X308 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X309 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t1866 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X310 VPWR.t1851 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X311 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t1083 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X312 VPWR.t1785 XThR.XTB5.Y a_n1049_6405# VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X313 VPWR.t1601 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1600 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X314 XThR.XTB7.B data[6].t0 VPWR.t238 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X315 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X316 VPWR.t915 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X317 VGND.t357 Vbias.t31 XA.XIR[10].XIC[9].icell.SM VGND.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X318 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t454 VPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1415 VPWR.t1417 VPWR.t1416 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X320 VGND.t1469 XThR.XTB2.Y XThR.Tn[1].t11 VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X321 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t1313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X322 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t2344 VGND.t2343 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X323 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t1002 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 XA.XIR[15].XIC[13].icell.Ien VPWR.t1412 VPWR.t1414 VPWR.t1413 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X325 VPWR.t958 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X326 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1939 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t1802 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X327 VPWR.t456 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t455 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X328 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t2531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X329 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t7 VPWR.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X330 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t113 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X331 VGND.t2598 XThC.XTBN.Y.t20 XThC.Tn[4].t3 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X332 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X333 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1410 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1411 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X334 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t245 VGND.t2551 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X335 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X336 VGND.t21 data[1].t1 a_8739_10571# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X337 XA.XIR[0].XIC[1].icell.PDM VGND.t1989 VGND.t1991 VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X338 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t202 VGND.t2365 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 VPWR.t1019 XThR.XTB2.Y XThR.Tn[9].t11 VPWR.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 VGND.t915 XThR.XTBN.Y XThR.Tn[7].t6 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X341 VGND.t1250 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t1249 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X342 VGND.t359 Vbias.t32 XA.XIR[13].XIC[5].icell.SM VGND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X343 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1940 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t1801 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X344 XThR.Tn[13].t3 XThR.XTBN.Y VPWR.t525 VPWR.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t2676 VGND.t2675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X346 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t658 VPWR.t657 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X347 VPWR.t1516 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1515 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X348 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1407 VPWR.t1409 VPWR.t1408 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X349 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t880 VPWR.t879 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X350 VPWR.t307 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t306 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X351 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t402 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X352 VGND.t361 Vbias.t33 XA.XIR[11].XIC[12].icell.SM VGND.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X353 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1404 VPWR.t1406 VPWR.t1405 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X354 VGND.t363 Vbias.t34 XA.XIR[7].XIC_15.icell.SM VGND.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X355 VPWR.t960 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t959 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X356 VGND.t1192 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t1191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X357 VGND.t2654 XThR.XTB6.Y XThR.Tn[5].t11 VGND.t2469 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X358 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t844 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X359 VGND.t365 Vbias.t35 XA.XIR[10].XIC[4].icell.SM VGND.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X360 XThR.Tn[9].t6 XThR.XTB2.Y a_n997_3755# VGND.t1299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X361 VGND.t1988 VGND.t1986 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1987 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X362 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t21 VGND.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X363 XThR.XTB6.Y XThR.XTB6.A VGND.t2548 VGND.t2547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X364 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1941 VGND.t1800 VGND.t1799 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X365 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t2503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X366 a_n997_1579# XThR.XTBN.Y VGND.t913 VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X367 VGND.t1498 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X368 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t210 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X369 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X370 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t61 VGND.t671 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X371 VPWR.t1716 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t1715 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X372 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1402 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1403 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X373 VPWR.t1057 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t1056 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X374 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t215 VGND.t2397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X375 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t1923 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X376 XA.XIR[15].XIC[6].icell.Ien VPWR.t1399 VPWR.t1401 VPWR.t1400 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X377 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1942 VGND.t1798 VGND.t1797 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X378 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t46 VGND.t561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X379 VPWR.t89 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X380 VPWR.t660 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t659 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X381 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t153 VGND.t1394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X382 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t164 VGND.t1449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X383 XA.XIR[15].XIC[9].icell.PDM VPWR.t1943 XA.XIR[15].XIC[9].icell.Ien VGND.t1796 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X384 VGND.t367 Vbias.t36 XA.XIR[13].XIC[0].icell.SM VGND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X385 VGND.t369 Vbias.t37 XA.XIR[8].XIC[12].icell.SM VGND.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X386 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t143 VGND.t1309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X387 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t130 VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X388 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t2678 VGND.t2677 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t2287 VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1944 VGND.t1795 VGND.t1794 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t2032 VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X392 VPWR.t544 XThR.XTBN.A XThR.XTBN.Y VPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X393 VPWR.t1754 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t1753 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X394 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X395 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t938 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X396 VGND.t371 Vbias.t38 XA.XIR[6].XIC[11].icell.SM VGND.t370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X397 VPWR.t1718 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t1717 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X398 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t216 VGND.t2398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X399 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t814 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X401 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1397 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X402 a_3523_10575# XThC.XTB7.B VGND.t131 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X403 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t704 VGND.t703 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t706 VGND.t705 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X405 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X406 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t1026 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X407 VPWR.t1893 XThC.XTBN.Y.t21 XThC.Tn[13].t3 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t1045 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X409 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X410 VGND.t70 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X411 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t91 VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X412 XThC.Tn[5].t11 XThC.XTB6.Y VGND.t1014 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XThC.Tn[4].t9 XThC.XTB5.Y VGND.t2262 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X414 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X415 VGND.t1793 VPWR.t1945 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t1792 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X416 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X417 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t1720 VPWR.t1719 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X418 VPWR.t19 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X419 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t1865 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X420 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t7 VGND.t2468 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X421 VPWR.t1550 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t1549 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X422 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t87 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X423 VPWR.t765 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t764 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X424 VGND.t1985 VGND.t1983 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X425 XA.XIR[15].XIC[1].icell.Ien VPWR.t1394 VPWR.t1396 VPWR.t1395 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X426 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1391 VPWR.t1393 VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X427 VGND.t1480 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t1479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X428 VGND.t1146 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t6 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 XThC.Tn[4].t2 XThC.XTBN.Y.t22 VGND.t2599 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VPWR.t922 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X432 a_n1049_5317# XThR.XTB7.Y VPWR.t1619 VPWR.t1618 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t1552 VPWR.t1551 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X434 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t23 VGND.t22 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X435 VPWR.t662 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t661 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X436 VGND.t373 Vbias.t39 XA.XIR[4].XIC[7].icell.SM VGND.t372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VPWR.t404 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t403 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X438 XThC.XTB6.Y XThC.XTB7.B VGND.t129 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X439 VPWR.t1390 VPWR.t1388 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1389 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 XA.XIR[15].XIC[4].icell.PDM VPWR.t1946 XA.XIR[15].XIC[4].icell.Ien VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X441 VPWR.t1853 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t1852 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X442 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1947 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t1790 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X443 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t3 VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X444 VGND.t375 Vbias.t40 XA.XIR[7].XIC[8].icell.SM VGND.t374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X445 VGND.t377 Vbias.t41 XA.XIR[6].XIC[9].icell.SM VGND.t376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X446 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t1047 VGND.t1046 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X447 VGND.t379 Vbias.t42 XA.XIR[3].XIC[11].icell.SM VGND.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X448 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t239 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t140 VGND.t1300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X450 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t218 VGND.t2400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X451 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X452 XThC.Tn[13].t7 XThC.XTB6.Y VPWR.t623 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X453 VGND.t663 XThC.XTBN.Y.t24 XThC.Tn[0].t7 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 XThR.Tn[3].t6 XThR.XTBN.Y a_n1049_6699# VPWR.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X456 VGND.t1194 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t1193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X457 VGND.t57 XThR.XTB4.Y.t3 XThR.Tn[3].t2 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X459 VGND.t381 Vbias.t43 XA.XIR[12].XIC[5].icell.SM VGND.t380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X460 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t1049 VGND.t1048 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t1034 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X462 VGND.t383 Vbias.t44 XA.XIR[15].XIC[6].icell.SM VGND.t382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X463 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t927 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t1422 VGND.t1421 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X465 XA.XIR[0].XIC_15.icell.PDM VPWR.t1948 VGND.t1789 VGND.t1788 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X466 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t1134 VGND.t1133 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X467 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t93 VPWR.t92 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X468 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t860 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X469 XThR.Tn[11].t2 XThR.XTB4.Y.t4 VPWR.t55 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X470 VGND.t1148 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t1147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X471 VGND.t1482 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t1481 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X472 XThC.Tn[14].t7 XThC.XTB7.Y a_10915_9569# VGND.t1410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X473 VPWR.t924 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t923 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X474 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X475 VGND.t1319 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t1318 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 VGND.t385 Vbias.t45 XA.XIR[9].XIC[5].icell.SM VGND.t384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X477 VPWR.t975 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X478 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X479 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X480 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1949 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X481 VPWR.t1387 VPWR.t1385 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X482 VGND.t387 Vbias.t46 XA.XIR[3].XIC[9].icell.SM VGND.t386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X483 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t842 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X484 VGND.t1310 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X485 VPWR.t1771 XThC.XTB2.Y XThC.Tn[9].t10 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X486 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t1756 VPWR.t1755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X487 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X488 VGND.t693 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X489 VGND.t1786 VPWR.t1950 XA.XIR[2].XIC_15.icell.PDM VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X490 VPWR.t1784 XThR.XTB5.Y XThR.Tn[12].t6 VPWR.t1527 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X491 VGND.t1500 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t1499 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X492 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t767 VPWR.t766 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X493 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t664 VPWR.t663 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X494 VGND.t389 Vbias.t47 XA.XIR[4].XIC[2].icell.SM VGND.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X495 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t579 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X496 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X497 VPWR.t1617 XThR.XTB7.Y XThR.Tn[14].t10 VPWR.t1616 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X498 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t222 VGND.t2404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X499 VGND.t391 Vbias.t48 XA.XIR[7].XIC[3].icell.SM VGND.t390 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X500 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t1051 VGND.t1050 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X501 VGND.t393 Vbias.t49 XA.XIR[6].XIC[4].icell.SM VGND.t392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X502 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t2033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X503 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X504 VGND.t395 Vbias.t50 XA.XIR[15].XIC[10].icell.SM VGND.t394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X505 XThR.Tn[8].t8 XThR.XTB1.Y.t4 a_n997_3979# VGND.t947 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X506 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t1424 VGND.t1423 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t158 VGND.t1412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X509 VGND.t1284 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X510 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1951 VGND.t1784 VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X511 VPWR.t1855 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t1854 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X512 VPWR.t1653 data[2].t0 XThC.XTB7.B VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X513 VPWR.t826 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X514 VGND.t397 Vbias.t51 XA.XIR[12].XIC[0].icell.SM VGND.t396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X515 VGND.t1583 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t1582 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X516 XThC.Tn[13].t10 XThC.XTB6.Y a_10051_9569# VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X517 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t114 VGND.t1090 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X518 XThR.Tn[4].t7 XThR.XTBN.Y a_n1049_6405# VPWR.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X519 VGND.t399 Vbias.t52 XA.XIR[15].XIC[1].icell.SM VGND.t398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X520 VGND.t401 Vbias.t53 XA.XIR[10].XIC[13].icell.SM VGND.t400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X521 XThC.Tn[8].t3 XThC.XTBN.Y.t25 VPWR.t376 VPWR.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X522 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X523 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t2035 VGND.t2034 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X524 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t900 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X525 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t61 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X526 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t1778 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X527 VGND.t1360 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1359 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X528 VGND.t242 Vbias.t54 XA.XIR[13].XIC[14].icell.SM VGND.t241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X529 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t309 VPWR.t308 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X530 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t1758 VPWR.t1757 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X531 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t90 VGND.t89 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X532 VGND.t1223 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t1222 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X533 XThC.Tn[8].t6 XThC.XTB1.Y.t4 a_7651_9569# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X534 VGND.t695 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X535 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t59 VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X536 XThC.Tn[13].t2 XThC.XTBN.Y.t26 VPWR.t378 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X537 VPWR.t555 VGND.t2690 XA.XIR[0].XIC[9].icell.PUM VPWR.t554 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X538 VGND.t1013 XThC.XTB6.Y XThC.Tn[5].t10 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X540 VGND.t244 Vbias.t55 XA.XIR[9].XIC[0].icell.SM VGND.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X541 VGND.t246 Vbias.t56 XA.XIR[0].XIC_15.icell.SM VGND.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X542 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1382 VPWR.t1384 VPWR.t1383 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X543 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t215 VGND.t214 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X544 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t217 VGND.t216 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X545 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t2036 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X546 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t602 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t251 VGND.t2655 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X548 VGND.t248 Vbias.t57 XA.XIR[3].XIC[4].icell.SM VGND.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X549 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t210 VGND.t2375 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X550 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t846 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X551 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X552 VGND.t72 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X553 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t155 VGND.t1396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X554 a_n1049_5611# XThR.XTB6.Y VPWR.t1904 VPWR.t1618 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X555 XA.XIR[13].XIC_15.icell.PUM VPWR.t1380 XA.XIR[13].XIC_15.icell.Ien VPWR.t1381 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 XThR.Tn[10].t11 XThR.XTB3.Y.t4 a_n997_2891# VGND.t2016 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X557 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1314 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X558 VGND.t2686 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t2685 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X559 VGND.t1502 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t1501 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X560 VPWR.t380 XThC.XTBN.Y.t27 XThC.Tn[7].t2 VPWR.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X561 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X562 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t1052 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X563 VPWR.t828 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t827 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X564 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t144 VGND.t1315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X565 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1378 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1379 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X566 VPWR.t1017 XThR.XTB2.Y XThR.Tn[9].t10 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X567 VPWR.t557 VGND.t2691 Vbias.t4 VPWR.t556 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X568 XThC.Tn[6].t2 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X569 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X570 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t666 VPWR.t665 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X571 VGND.t1240 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t1239 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X572 VPWR.t132 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X573 VPWR.t1857 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t1856 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X574 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X575 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1736 VPWR.t1735 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X576 VGND.t1225 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t1224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X577 XA.XIR[15].XIC_15.icell.Ien VPWR.t1375 VPWR.t1377 VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X578 VPWR.t830 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t829 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X579 VPWR.t1760 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t1759 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X580 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t5 VPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X581 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X582 XThC.Tn[0].t6 XThC.XTBN.Y.t29 VGND.t664 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X583 VPWR.t1374 VPWR.t1372 XA.XIR[9].XIC_15.icell.PUM VPWR.t1373 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X584 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t217 VGND.t2399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X585 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t741 VGND.t740 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X586 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t743 VGND.t742 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X587 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t54 VGND.t631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X588 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t3 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X589 XThR.Tn[0].t1 XThR.XTB1.Y.t5 VGND.t709 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X590 VGND.t912 XThR.XTBN.Y XThR.Tn[5].t6 VGND.t898 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X591 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t1762 VPWR.t1761 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X592 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t2119 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X593 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t92 VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X594 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t2533 VGND.t2532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X596 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t1207 VGND.t1206 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X597 VGND.t1782 VPWR.t1952 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X598 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t582 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X599 VGND.t911 XThR.XTBN.Y XThR.Tn[4].t3 VGND.t910 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X600 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t2289 VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X601 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t816 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X602 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t23 VGND.t113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X603 VGND.t1780 VPWR.t1953 XA.XIR[14].XIC_15.icell.PDM VGND.t1779 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t5 VGND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X605 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t8 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X606 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X607 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1370 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1371 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t242 VGND.t2534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X609 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t862 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X610 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t744 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X611 VGND.t74 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t529 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X613 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1738 VPWR.t1737 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X614 VGND.t1321 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VPWR.t1722 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t1721 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X616 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X617 VGND.t665 XThC.XTBN.Y.t31 a_8739_9569# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X618 VGND.t1252 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VGND.t250 Vbias.t58 XA.XIR[11].XIC[6].icell.SM VGND.t249 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X620 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1954 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t1778 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X621 VPWR.t734 bias[0].t0 Vbias.t1 VPWR.t556 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=4
X622 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t977 VPWR.t976 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X623 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t668 VPWR.t667 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X624 VGND.t1150 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t1149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X625 VGND.t1484 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t1483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X626 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1740 VPWR.t1739 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X627 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t773 VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X628 a_9827_9569# XThC.XTBN.Y.t32 VGND.t666 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X629 VPWR.t678 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t677 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X630 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X631 VPWR.t436 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X632 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1955 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X633 VGND.t252 Vbias.t59 XA.XIR[0].XIC[8].icell.SM VGND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X634 VGND.t1982 VGND.t1980 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X635 VPWR.t979 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t978 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X636 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t2345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X637 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t2291 VGND.t2290 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X638 VPWR.t1369 VPWR.t1367 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1368 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X639 XA.XIR[15].XIC[13].icell.PDM VPWR.t1956 XA.XIR[15].XIC[13].icell.Ien VGND.t1776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X640 VGND.t2206 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X641 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t27 VGND.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X642 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t746 VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X643 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t135 VGND.t1228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X644 XThR.XTB7.A data[5].t1 VPWR.t399 VPWR.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X645 VGND.t1581 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t1580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X646 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t71 VGND.t777 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X647 VPWR.t97 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X648 VGND.t254 Vbias.t60 XA.XIR[5].XIC[5].icell.SM VGND.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X649 VGND.t1216 XThC.XTBN.A XThC.XTBN.Y.t3 VGND.t1215 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t1036 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X651 VGND.t256 Vbias.t61 XA.XIR[11].XIC[10].icell.SM VGND.t255 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X652 VPWR.t433 XThR.XTB7.B XThR.XTB1.Y.t0 VPWR.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X653 VGND.t258 Vbias.t62 XA.XIR[8].XIC[6].icell.SM VGND.t257 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X654 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t6 VGND.t2467 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X655 VGND.t260 Vbias.t63 XA.XIR[12].XIC[14].icell.SM VGND.t259 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X656 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t1864 VGND.t1863 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X657 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t981 VPWR.t980 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X658 XA.XIR[14].XIC_15.icell.PDM VPWR.t1957 VGND.t1775 VGND.t1774 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X659 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1364 VPWR.t1366 VPWR.t1365 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X660 VPWR.t680 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t679 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X661 VGND.t262 Vbias.t64 XA.XIR[11].XIC[1].icell.SM VGND.t261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X662 VGND.t264 Vbias.t65 XA.XIR[7].XIC[12].icell.SM VGND.t263 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X663 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X664 VGND.t266 Vbias.t66 XA.XIR[6].XIC[13].icell.SM VGND.t265 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X665 XThC.Tn[7].t1 XThC.XTBN.Y.t33 VPWR.t382 VPWR.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X666 VGND.t737 XThR.XTB7.B a_n1335_7243# VGND.t736 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X667 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X668 VGND.t268 Vbias.t67 XA.XIR[9].XIC[14].icell.SM VGND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X669 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t748 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1958 VGND.t1773 VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[12].XIC_15.icell.PUM VPWR.t1362 XA.XIR[12].XIC_15.icell.Ien VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t6 VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X674 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t1533 VGND.t1532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X675 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X676 VGND.t2199 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t653 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X678 VGND.t1504 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t1503 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X679 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1514 VPWR.t1513 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X680 XThC.Tn[11].t9 XThC.XTB4.Y.t6 VPWR.t916 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 VGND.t1506 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t1505 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X682 VGND.t270 Vbias.t68 XA.XIR[0].XIC[3].icell.SM VGND.t269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X683 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1359 VPWR.t1361 VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X684 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t121 VGND.t1160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X685 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t42 VGND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X686 a_n997_1803# XThR.XTBN.Y VGND.t909 VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X687 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X688 XThR.Tn[3].t5 XThR.XTBN.Y a_n1049_6699# VPWR.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X689 VPWR.t63 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X690 VGND.t907 XThR.XTBN.Y XThR.Tn[3].t9 VGND.t873 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X691 VGND.t272 Vbias.t69 XA.XIR[8].XIC[10].icell.SM VGND.t271 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X692 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t832 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X693 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t832 VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X694 VGND.t1771 VPWR.t1959 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t1770 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X695 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1960 VGND.t1769 VGND.t1768 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X696 XThC.Tn[2].t2 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X697 VPWR.t1742 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t1741 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t583 VPWR.t582 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X699 VPWR.t749 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t748 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X700 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t52 VGND.t600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X701 VPWR.t99 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X702 XThR.Tn[11].t3 XThR.XTB4.Y.t5 VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X703 VGND.t274 Vbias.t70 XA.XIR[5].XIC[0].icell.SM VGND.t273 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X704 VPWR.t1358 VPWR.t1356 XA.XIR[8].XIC_15.icell.PUM VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X705 VGND.t1979 VGND.t1977 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X706 VPWR.t1770 XThC.XTB2.Y a_3773_9615# VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t1071 VPWR.t1070 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X708 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1354 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1355 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X709 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t97 VGND.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X710 VGND.t276 Vbias.t71 XA.XIR[8].XIC[1].icell.SM VGND.t275 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X711 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t1862 VGND.t1861 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X712 VGND.t278 Vbias.t72 XA.XIR[3].XIC[13].icell.SM VGND.t277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X713 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X714 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t142 VGND.t1302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X715 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t1209 VGND.t1208 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X716 VGND.t752 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X717 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t2360 VGND.t2359 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X718 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1496 VPWR.t1495 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X720 VGND.t1767 VPWR.t1961 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t1766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X721 VPWR.t1579 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t1578 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X722 VPWR.t1849 XThC.XTB6.A a_5949_10571# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X723 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t75 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 VGND.t280 Vbias.t73 XA.XIR[2].XIC[11].icell.SM VGND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X725 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t817 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X726 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t231 VGND.t2510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X727 VGND.t1076 XThR.XTB3.Y.t5 XThR.Tn[2].t9 VGND.t1075 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X728 VPWR.t585 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t584 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X729 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X731 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X732 VGND.t282 Vbias.t74 XA.XIR[14].XIC_15.icell.SM VGND.t281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X733 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t109 VGND.t1084 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X734 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t1535 VGND.t1534 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 XThC.XTBN.Y.t1 XThC.XTBN.A VPWR.t840 VPWR.t839 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X736 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X737 VGND.t76 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X738 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t834 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X739 XThR.Tn[8].t10 XThR.XTB1.Y.t7 a_n997_3979# VGND.t1299 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X740 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t1393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X741 XA.XIR[6].XIC_15.icell.PUM VPWR.t1352 XA.XIR[6].XIC_15.icell.Ien VPWR.t1353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t1196 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X743 VGND.t78 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X744 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t460 VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X745 VGND.t1765 VPWR.t1962 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t1764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X746 VGND.t2228 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t2227 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X747 VGND.t1254 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t1253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X748 VGND.t667 XThC.XTBN.Y.t35 a_9827_9569# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X749 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t70 VGND.t757 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X750 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t928 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X751 VPWR.t65 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t64 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X752 VPWR.t967 XThC.XTB7.Y XThC.Tn[14].t11 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X753 XThR.Tn[4].t6 XThR.XTBN.Y a_n1049_6405# VPWR.t523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X754 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X755 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X756 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t836 VPWR.t835 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X757 VPWR.t47 XThR.XTB4.Y.t6 a_n1049_6699# VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X758 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t1764 VPWR.t1763 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X759 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t196 VGND.t2353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X760 VPWR.t1744 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t1743 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X761 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t587 VPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X762 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t67 VPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X763 VPWR.t751 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t750 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X764 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t1069 VPWR.t1068 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X765 XA.XIR[15].XIC[1].icell.PDM VPWR.t1963 XA.XIR[15].XIC[1].icell.Ien VGND.t1763 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 VPWR.t1724 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t1723 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X767 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t1450 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X768 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1964 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t1762 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X769 VGND.t284 Vbias.t75 XA.XIR[2].XIC[9].icell.SM VGND.t283 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X770 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t1746 VPWR.t1745 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X771 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t95 VGND.t1000 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X772 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t241 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X773 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t90 VGND.t992 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X774 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t2341 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X775 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t255 VGND.t2682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X776 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t73 VGND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X777 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t2362 VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X778 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t58 VGND.t668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X779 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1512 VPWR.t1511 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X780 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t228 VGND.t2487 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X781 VPWR.t522 XThR.XTBN.Y XThR.Tn[8].t6 VPWR.t521 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X782 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t462 VPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X783 XThR.Tn[10].t0 XThR.XTB3.Y.t6 a_n997_2891# VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X784 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X785 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X786 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t110 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X787 VPWR.t1848 XThC.XTB6.A XThC.XTB2.Y VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X788 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t2348 VGND.t2347 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X789 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t431 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X790 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X791 VGND.t531 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X792 VGND.t1323 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t1322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 XThR.XTB3.Y.t2 XThR.XTB7.A VPWR.t689 VPWR.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X794 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X795 VGND.t1256 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t1255 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X796 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t774 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X797 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1965 VGND.t1761 VGND.t1760 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X798 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t2118 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X799 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X800 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t654 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X801 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t1581 VPWR.t1580 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X802 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t2367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X803 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t1748 VPWR.t1747 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X804 XThR.Tn[0].t9 XThR.XTBN.Y VGND.t906 VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X805 VPWR.t1783 XThR.XTB5.Y a_n1049_6405# VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X806 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t753 VPWR.t752 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X807 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t1451 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X808 XThC.Tn[10].t1 XThC.XTB3.Y.t4 VPWR.t612 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X809 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t2363 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X810 VPWR.t520 XThR.XTBN.Y XThR.Tn[10].t7 VPWR.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 VGND.t286 Vbias.t76 XA.XIR[2].XIC[4].icell.SM VGND.t285 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X812 VPWR.t216 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t215 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X813 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t213 VGND.t2395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X814 VPWR.t383 XThC.XTBN.Y.t36 XThC.Tn[13].t1 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X816 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t1536 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X817 VGND.t288 Vbias.t77 XA.XIR[15].XIC[7].icell.SM VGND.t287 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X818 a_3773_9615# XThC.XTB2.Y VPWR.t1769 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X819 XThC.Tn[5].t9 XThC.XTB6.Y VGND.t1012 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X820 VGND.t449 Vbias.t78 XA.XIR[14].XIC[8].icell.SM VGND.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X821 XThC.Tn[2].t8 XThC.XTB3.Y.t5 VGND.t998 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 VPWR.t1726 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t1725 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X823 VPWR.t1510 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1509 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X824 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t96 VGND.t95 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X825 VGND.t1579 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X826 VPWR.t311 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t310 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X827 VPWR.t943 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t942 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X828 VGND.t905 XThR.XTBN.Y a_n997_3755# VGND.t894 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X829 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X830 VGND.t451 Vbias.t79 XA.XIR[5].XIC[14].icell.SM VGND.t450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X831 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t48 VGND.t563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X832 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t66 VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X833 VPWR.t713 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1966 VGND.t1759 VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X835 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X836 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t1583 VPWR.t1582 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X837 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t98 VGND.t97 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X838 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t433 VGND.t432 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X839 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t929 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X840 VGND.t453 Vbias.t80 XA.XIR[1].XIC[11].icell.SM VGND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X841 VGND.t1286 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t1285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X842 XA.XIR[11].XIC_15.icell.PDM VPWR.t1967 VGND.t1757 VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X843 VGND.t455 Vbias.t81 XA.XIR[0].XIC[12].icell.SM VGND.t454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X844 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t1361 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X845 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t775 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X846 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X847 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t107 VGND.t1065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X848 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t1645 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 a_5155_9615# XThC.XTB5.Y VPWR.t1686 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X850 XA.XIR[5].XIC_15.icell.PUM VPWR.t1350 XA.XIR[5].XIC_15.icell.Ien VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X851 VPWR.t218 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t217 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X852 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t584 VGND.t583 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X853 VGND.t1198 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t1197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X854 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t343 VPWR.t342 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X855 XA.XIR[9].XIC_15.icell.PUM VPWR.t1348 XA.XIR[9].XIC_15.icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X856 VGND.t971 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t970 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X857 VPWR.t1508 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1507 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X858 VPWR.t186 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X859 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t63 VGND.t679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X860 VGND.t1755 VPWR.t1968 XA.XIR[13].XIC_15.icell.PDM VGND.t1754 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X861 VGND.t457 Vbias.t82 XA.XIR[15].XIC[2].icell.SM VGND.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X862 XThC.Tn[8].t11 XThC.XTB1.Y.t7 VPWR.t715 VPWR.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X863 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X864 VGND.t459 Vbias.t83 XA.XIR[14].XIC[3].icell.SM VGND.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X865 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t102 VGND.t1010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X866 Vbias.t5 bias[2].t0 VPWR.t1561 VPWR.t1560 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=1
X867 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t755 VPWR.t754 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X868 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t1728 VPWR.t1727 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X869 VGND.t2470 XThR.XTB5.Y XThR.Tn[4].t11 VGND.t2469 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X870 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t7 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X871 VGND.t1753 VPWR.t1969 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t1752 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X872 VPWR.t1730 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1729 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X873 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t100 VGND.t99 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t1506 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1505 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XThR.XTB5.Y XThR.XTB5.A VGND.t2681 VGND.t2547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X876 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t435 VGND.t434 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X877 VPWR.t188 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X878 VPWR.t1585 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t1584 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X879 VPWR.t945 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t944 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X881 VGND.t461 Vbias.t84 XA.XIR[1].XIC[9].icell.SM VGND.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X882 VPWR.t1347 VPWR.t1345 XA.XIR[1].XIC_15.icell.PUM VPWR.t1346 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X883 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t1125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X884 VPWR.t1344 VPWR.t1342 XA.XIR[5].XIC_15.icell.PUM VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t67 VGND.t696 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X886 XA.XIR[15].XIC_15.icell.PDM VPWR.t1970 XA.XIR[15].XIC_15.icell.Ien VGND.t1751 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X887 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t243 VGND.t2535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X888 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X889 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t1587 VPWR.t1586 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X890 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t2 VGND.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X891 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t1860 VGND.t1859 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X892 VGND.t1750 VPWR.t1971 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t1749 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t641 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X894 VPWR.t1341 VPWR.t1339 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1340 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X895 XThC.Tn[14].t6 XThC.XTB7.Y a_10915_9569# VGND.t1409 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X896 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X897 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t168 VGND.t1458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X898 a_n997_1803# XThR.XTBN.Y VGND.t904 VGND.t903 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t903 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X900 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1732 VPWR.t1731 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X901 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t3 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X903 VGND.t602 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t601 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X905 VGND.t463 Vbias.t85 XA.XIR[4].XIC[5].icell.SM VGND.t462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X906 VGND.t1288 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t1287 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X907 VPWR.t990 XThC.XTB5.A XThC.XTB1.Y.t1 VPWR.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X908 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1972 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t1748 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X909 VGND.t1290 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t1289 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X910 VGND.t465 Vbias.t86 XA.XIR[7].XIC[6].icell.SM VGND.t464 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X911 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1973 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t1747 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t2074 VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t757 VPWR.t756 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X915 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1734 VPWR.t1733 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X916 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t101 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X917 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1337 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X918 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1504 VPWR.t1503 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X919 VGND.t999 XThC.XTB3.Y.t6 XThC.Tn[2].t9 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X920 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X921 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t2 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X922 VGND.t467 Vbias.t87 XA.XIR[1].XIC[4].icell.SM VGND.t466 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X923 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t1537 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X924 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t1126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X925 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t2292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X926 a_n1319_6405# XThR.XTB5.A VPWR.t1921 VPWR.t1920 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X927 VPWR.t25 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X928 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X929 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t444 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X930 VPWR.t1336 VPWR.t1334 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X931 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t10 VGND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X932 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t571 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X933 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t717 VPWR.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X934 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t1750 VPWR.t1749 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X935 XThR.Tn[12].t2 XThR.XTBN.Y VPWR.t518 VPWR.t517 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X936 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1331 VPWR.t1333 VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X937 XThC.Tn[11].t5 XThC.XTBN.Y.t39 VPWR.t33 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X938 VGND.t1004 data[4].t2 XThR.XTB5.A VGND.t1003 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X939 XThR.XTBN.Y XThR.XTBN.A VGND.t942 VGND.t941 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X940 VGND.t469 Vbias.t88 XA.XIR[11].XIC[7].icell.SM VGND.t468 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X941 VGND.t471 Vbias.t89 XA.XIR[7].XIC[10].icell.SM VGND.t470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X942 VGND.t1113 data[3].t0 XThC.XTBN.A VGND.t1112 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X943 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t212 VGND.t2394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X944 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1974 VGND.t1746 VGND.t1745 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X945 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t1539 VGND.t1538 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X946 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t11 VGND.t2468 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X947 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X948 VGND.t473 Vbias.t90 XA.XIR[4].XIC[0].icell.SM VGND.t472 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X949 XA.XIR[10].XIC_15.icell.PDM VPWR.t1975 VGND.t1744 VGND.t1743 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X950 a_n997_2667# XThR.XTBN.Y VGND.t902 VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X951 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1329 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X952 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t170 VGND.t1470 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 VGND.t475 Vbias.t91 XA.XIR[7].XIC[1].icell.SM VGND.t474 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X955 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t2076 VGND.t2075 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X956 VGND.t477 Vbias.t92 XA.XIR[2].XIC[13].icell.SM VGND.t476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X957 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t1274 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X958 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t902 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X959 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X960 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t2563 VGND.t2562 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t51 VGND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X962 VPWR.t27 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X963 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t219 VGND.t218 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X964 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t655 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 VGND.t1426 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t1425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X966 XThC.Tn[4].t6 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X967 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t2488 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X968 VGND.t1742 VPWR.t1976 XA.XIR[12].XIC_15.icell.PDM VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X969 VPWR.t246 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t245 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X970 VPWR.t516 XThR.XTBN.Y XThR.Tn[8].t5 VPWR.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X971 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t60 VGND.t670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X972 VGND.t2240 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t2239 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X973 VGND.t1034 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t1033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X974 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X975 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t1664 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1326 VPWR.t1328 VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X977 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t5 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X978 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t1858 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X979 VGND.t479 Vbias.t93 XA.XIR[8].XIC[7].icell.SM VGND.t478 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X980 VPWR.t1685 XThC.XTB5.Y XThC.Tn[12].t5 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X981 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t99 VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X982 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1977 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t1740 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X983 VPWR.t888 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t887 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X984 VPWR.t1325 VPWR.t1323 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X985 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X986 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t947 VPWR.t946 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X987 VGND.t1976 VGND.t1974 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X988 VGND.t2230 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t2229 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X989 VGND.t901 XThR.XTBN.Y XThR.Tn[1].t3 VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X990 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t35 VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t1363 VGND.t1362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X992 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X993 VPWR.t559 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t558 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X994 VPWR.t1322 VPWR.t1320 XA.XIR[4].XIC_15.icell.PUM VPWR.t1321 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X995 VGND.t481 Vbias.t94 XA.XIR[11].XIC[2].icell.SM VGND.t480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X996 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t1752 VPWR.t1751 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X997 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t952 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X998 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t953 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X999 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t40 VGND.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1000 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t1857 VGND.t1856 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1001 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t240 VGND.t2527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1002 XThR.Tn[6].t10 XThR.XTB7.Y VGND.t2117 VGND.t2116 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_9827_9569# XThC.XTBN.Y.t41 VGND.t37 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1004 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t1906 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XThR.Tn[9].t1 XThR.XTBN.Y VPWR.t514 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t221 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t1365 VGND.t1364 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1008 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t982 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1009 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t2352 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1010 VGND.t2658 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t2657 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1011 XThC.Tn[1].t2 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1012 XThR.Tn[0].t8 XThR.XTBN.Y VGND.t900 VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 XThC.Tn[13].t9 XThC.XTB6.Y a_10051_9569# VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1014 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1015 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t16 VGND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1016 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t117 VGND.t1099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1017 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t1855 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1018 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t605 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1019 VPWR.t513 XThR.XTBN.Y XThR.Tn[10].t6 VPWR.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1020 VPWR.t71 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1021 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1022 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t2565 VGND.t2564 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t53 VGND.t617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1024 VGND.t483 Vbias.t95 XA.XIR[14].XIC[12].icell.SM VGND.t482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1025 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1317 VPWR.t1319 VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1026 VGND.t485 Vbias.t96 XA.XIR[10].XIC_15.icell.SM VGND.t484 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1027 XA.XIR[0].XIC[12].icell.PDM VGND.t1971 VGND.t1973 VGND.t1972 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1028 VGND.t80 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1029 VGND.t604 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1030 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t192 VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1031 VPWR.t966 XThC.XTB7.Y a_6243_9615# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1032 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1978 VGND.t1739 VGND.t1738 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 VGND.t606 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1034 VGND.t2232 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t2231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t589 VPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1036 VGND.t973 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t972 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t156 VGND.t1397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1038 VPWR.t561 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t560 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1039 VGND.t2201 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1040 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t1452 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1041 VGND.t1737 VPWR.t1979 XA.XIR[6].XIC_15.icell.PDM VGND.t1736 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1042 VGND.t38 XThC.XTBN.Y.t43 a_8963_9569# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1043 VGND.t487 Vbias.t97 XA.XIR[8].XIC[2].icell.SM VGND.t486 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1044 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t100 VGND.t1008 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1045 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1046 VPWR.t1067 XThR.XTB1.Y.t8 XThR.Tn[8].t11 VPWR.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1047 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1315 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1048 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t88 VGND.t965 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1049 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1050 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t118 VGND.t1107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1051 VGND.t533 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1052 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t910 VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1053 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t949 VPWR.t948 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1054 VGND.t2177 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t2176 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1055 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t1367 VGND.t1366 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1056 XThR.XTBN.A data[7].t0 VPWR.t884 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1057 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t73 VPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1058 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t1881 VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1059 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1060 VPWR.t563 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t562 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1061 VPWR.t1016 XThR.XTB2.Y a_n1049_7787# VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1062 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t1453 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1063 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t1563 VPWR.t1562 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1065 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 VPWR.t890 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t889 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1067 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t162 VGND.t1440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1068 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t78 VGND.t943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1069 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1070 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t104 VGND.t1020 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1071 XA.XIR[0].XIC[10].icell.PDM VGND.t1968 VGND.t1970 VGND.t1969 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1072 VGND.t1967 VGND.t1965 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1073 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t2053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1074 a_n1049_7493# XThR.XTBN.Y XThR.Tn[2].t4 VPWR.t511 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1075 VGND.t643 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1076 XThC.Tn[8].t10 XThC.XTB1.Y.t10 VPWR.t719 VPWR.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 VPWR.t998 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1078 VPWR.t1314 VPWR.t1312 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1313 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1079 VGND.t754 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1080 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t229 VGND.t2502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1081 XThR.Tn[0].t10 XThR.XTB1.Y.t9 VGND.t1073 VGND.t1072 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1082 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t776 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1083 VGND.t489 Vbias.t98 XA.XIR[13].XIC[11].icell.SM VGND.t488 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1084 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1085 VPWR.t1662 XThR.XTB3.Y.t8 XThR.Tn[10].t10 VPWR.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1086 VGND.t1577 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t1576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1087 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t2537 VGND.t2536 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1088 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t2539 VGND.t2538 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1089 VPWR.t1768 XThC.XTB2.Y a_3773_9615# VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 VGND.t535 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 VGND.t899 XThR.XTBN.Y XThR.Tn[4].t2 VGND.t898 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1092 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1310 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1311 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t1665 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1094 VGND.t491 Vbias.t99 XA.XIR[1].XIC[13].icell.SM VGND.t490 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1095 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t1454 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 VPWR.t36 XThC.XTBN.Y.t44 XThC.Tn[9].t3 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 VGND.t493 Vbias.t100 XA.XIR[0].XIC[6].icell.SM VGND.t492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1098 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1980 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t1735 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1099 VGND.t495 Vbias.t101 XA.XIR[4].XIC[14].icell.SM VGND.t494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1100 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t2540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1101 VGND.t40 XThC.XTBN.Y.t45 XThC.Tn[5].t1 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1102 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t2490 VGND.t2489 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1103 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1104 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t244 VGND.t2550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1105 VGND.t897 XThR.XTBN.Y a_n997_1579# VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1106 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t1634 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1107 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t1 VPWR.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1108 VGND.t2242 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t2241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1109 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1110 VGND.t1036 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t1035 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t1303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VPWR.t892 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t891 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1113 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t446 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1114 XThC.Tn[12].t10 XThC.XTB5.Y a_9827_9569# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1115 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t24 VGND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1116 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1117 VPWR.t1000 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1118 XThR.XTB6.A data[5].t2 VPWR.t886 VPWR.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1119 VGND.t2294 Vbias.t102 XA.XIR[10].XIC[8].icell.SM VGND.t2293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1120 VPWR.t1309 VPWR.t1307 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1121 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t2115 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1122 VPWR.t29 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t28 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1123 VGND.t2296 Vbias.t103 XA.XIR[13].XIC[9].icell.SM VGND.t2295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1124 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t3 VPWR.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1125 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t894 VPWR.t893 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1126 XA.XIR[15].XIC[12].icell.Ien VPWR.t1304 VPWR.t1306 VPWR.t1305 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1127 VPWR.t912 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t911 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1128 VGND.t2298 Vbias.t104 XA.XIR[0].XIC[10].icell.SM VGND.t2297 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1129 VPWR.t136 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t135 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1130 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t2541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1131 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1981 VGND.t1734 VGND.t1733 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1132 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t2055 VGND.t2054 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1133 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1134 VGND.t1964 VGND.t1962 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1963 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1135 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t2543 VGND.t2542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[3].XIC_15.icell.PDM VPWR.t1982 VGND.t1732 VGND.t1731 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1137 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t121 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1138 a_6243_9615# XThC.XTB7.Y VPWR.t965 VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1139 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1302 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1303 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1140 VGND.t2300 Vbias.t105 XA.XIR[0].XIC[1].icell.SM VGND.t2299 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1141 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t163 VGND.t1442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1142 XThC.Tn[10].t0 XThC.XTBN.Y.t47 VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1143 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t1304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1144 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t1907 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1145 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t2492 VGND.t2491 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1146 VGND.t2179 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t2178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1147 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t55 VGND.t632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1148 XA.XIR[1].XIC_15.icell.PUM VPWR.t1300 XA.XIR[1].XIC_15.icell.Ien VPWR.t1301 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XThC.Tn[10].t3 XThC.XTB3.Y.t8 a_8739_9569# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1150 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t1306 VGND.t1305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1151 VGND.t1408 XThC.XTB7.Y XThC.Tn[6].t11 VGND.t1407 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1152 VGND.t1730 VPWR.t1983 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t1729 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1153 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1984 VGND.t1728 VGND.t1727 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1154 XThR.Tn[11].t6 XThR.XTBN.Y VPWR.t510 VPWR.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1155 VGND.t2203 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t2202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1156 VPWR.t41 XThC.XTBN.Y.t48 XThC.Tn[12].t3 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 VGND.t1726 VPWR.t1985 XA.XIR[5].XIC_15.icell.PDM VGND.t1725 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 XA.XIR[15].XIC[10].icell.Ien VPWR.t1297 VPWR.t1299 VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1159 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t248 VPWR.t247 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1160 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t896 VPWR.t895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 VGND.t1724 VPWR.t1986 XA.XIR[9].XIC_15.icell.PDM VGND.t1723 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1162 VPWR.t951 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t950 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1163 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1164 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t69 VGND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1165 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1294 VPWR.t1296 VPWR.t1295 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1166 VGND.t2302 Vbias.t106 XA.XIR[6].XIC_15.icell.SM VGND.t2301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1167 VPWR.t138 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t137 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1168 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t1162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1169 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t189 VGND.t2101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1170 VGND.t2304 Vbias.t107 XA.XIR[10].XIC[3].icell.SM VGND.t2303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1171 VGND.t2234 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t2233 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1172 VGND.t2306 Vbias.t108 XA.XIR[13].XIC[4].icell.SM VGND.t2305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t1961 VGND.t1959 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1174 VGND.t2505 XThC.XTB7.A XThC.XTB7.Y VGND.t2504 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1175 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t2545 VGND.t2544 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1176 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1502 VPWR.t1501 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1177 VPWR.t914 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t913 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1178 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t10 VGND.t2467 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1179 a_n997_2667# XThR.XTBN.Y VGND.t896 VGND.t853 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 VPWR.t31 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1181 VPWR.t357 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1182 a_7875_9569# XThC.XTBN.Y.t49 VGND.t42 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1183 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t2057 VGND.t2056 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1184 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t45 VGND.t338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1185 VGND.t1575 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1186 VGND.t895 XThR.XTBN.Y a_n997_3979# VGND.t894 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1187 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t1565 VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1188 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1189 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t29 VGND.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1190 XThC.Tn[14].t2 XThC.XTBN.Y.t50 VPWR.t43 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1191 a_n1049_6699# XThR.XTB4.Y.t7 VPWR.t49 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1192 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t7 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1193 VGND.t756 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1194 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t72 VGND.t778 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1195 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t250 VPWR.t249 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1196 XThC.Tn[2].t10 XThC.XTB3.Y.t9 VGND.t1074 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1197 XThC.Tn[9].t2 XThC.XTBN.Y.t52 VPWR.t45 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1198 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t4 VGND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1199 VGND.t2308 Vbias.t109 XA.XIR[3].XIC_15.icell.SM VGND.t2307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1200 VGND.t2310 Vbias.t110 XA.XIR[12].XIC[11].icell.SM VGND.t2309 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1201 VGND.t1958 VGND.t1956 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1957 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1202 XThC.Tn[5].t0 XThC.XTBN.Y.t53 VGND.t2271 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1203 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1204 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t629 VGND.t628 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1205 VGND.t1292 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t1291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1206 XA.XIR[15].XIC[5].icell.Ien VPWR.t1291 VPWR.t1293 VPWR.t1292 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1207 VPWR.t721 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1208 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1987 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t1722 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 XThC.Tn[0].t0 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t1694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1210 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t2493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1211 VPWR.t140 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1212 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t235 VGND.t2514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1213 VPWR.t359 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1214 XThR.Tn[12].t5 XThR.XTB5.Y VPWR.t1782 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1215 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t1640 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t1635 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1217 VGND.t2312 Vbias.t111 XA.XIR[9].XIC[11].icell.SM VGND.t2311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1218 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1289 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1290 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1219 VGND.t537 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t536 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1220 XThR.Tn[6].t6 XThR.XTBN.Y VGND.t893 VGND.t892 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1221 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t2 VPWR.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1222 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t904 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1223 VGND.t891 XThR.XTBN.Y a_n997_2891# VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1224 VGND.t735 XThR.XTB7.B XThR.XTB7.Y VGND.t734 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1225 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1500 VPWR.t1499 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1226 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t1200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1227 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1228 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t2494 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1229 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t166 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1230 VPWR.t168 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1231 VGND.t1721 VPWR.t1988 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t1720 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1232 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t656 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1233 VPWR.t361 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t1411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1235 a_n997_2667# XThR.XTB4.Y.t8 XThR.Tn[11].t0 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1236 VPWR.t1288 VPWR.t1286 XA.XIR[12].XIC_15.icell.PUM VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1237 VGND.t2314 Vbias.t112 XA.XIR[12].XIC[9].icell.SM VGND.t2313 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1238 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t1002 VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1239 VGND.t1955 VGND.t1953 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1240 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1283 VPWR.t1285 VPWR.t1284 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1241 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t2028 VGND.t2027 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1242 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1280 VPWR.t1282 VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1243 VGND.t2272 XThC.XTBN.Y.t55 XThC.Tn[1].t5 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 a_n1049_6405# XThR.XTB5.Y VPWR.t1781 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1245 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t252 VPWR.t251 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1246 VPWR.t1859 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t1858 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1247 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t2058 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1248 VGND.t2316 Vbias.t113 XA.XIR[7].XIC[7].icell.SM VGND.t2315 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1249 VGND.t2318 Vbias.t114 XA.XIR[6].XIC[8].icell.SM VGND.t2317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1250 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1989 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t1719 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t1718 VPWR.t1990 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t1717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1252 VPWR.t1623 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t1622 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1253 VGND.t2320 Vbias.t115 XA.XIR[9].XIC[9].icell.SM VGND.t2319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1254 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t2569 VGND.t2568 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1255 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t125 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1256 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t197 VGND.t2354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1257 VPWR.t650 XThR.XTB1.Y.t10 XThR.Tn[8].t9 VPWR.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1258 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t243 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1259 VPWR.t508 XThR.XTBN.Y XThR.Tn[7].t2 VPWR.t507 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1260 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1278 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1261 VGND.t2379 XThC.XTB2.Y XThC.Tn[1].t11 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1262 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1276 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1263 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t2495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1264 XThC.Tn[12].t2 XThC.XTBN.Y.t56 VPWR.t1695 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t1308 VGND.t1307 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1266 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t170 VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1267 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t62 VGND.t672 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1268 VGND.t1467 XThR.XTB2.Y XThR.Tn[1].t10 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1269 XThR.Tn[1].t6 XThR.XTBN.Y a_n1049_7787# VPWR.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1270 VGND.t2322 Vbias.t116 XA.XIR[15].XIC[5].icell.SM VGND.t2321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1271 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t2571 VGND.t2570 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 VGND.t2324 Vbias.t117 XA.XIR[14].XIC[6].icell.SM VGND.t2323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1273 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t1636 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t539 VGND.t538 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1275 VGND.t2660 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1276 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t1698 VPWR.t1697 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1277 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t1625 VPWR.t1624 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1278 VGND.t1038 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t1037 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1279 VGND.t2244 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t2243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1280 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t172 VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1281 XThR.Tn[9].t9 XThR.XTB2.Y VPWR.t1015 VPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1282 XThR.Tn[7].t5 XThR.XTBN.Y VGND.t889 VGND.t888 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1283 VPWR.t711 data[1].t2 XThC.XTB6.A VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1284 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1285 VPWR.t1700 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t1699 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1286 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t363 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1287 VGND.t2326 Vbias.t118 XA.XIR[12].XIC[4].icell.SM VGND.t2325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1288 VPWR.t1275 VPWR.t1273 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1289 VGND.t2328 Vbias.t119 XA.XIR[3].XIC[8].icell.SM VGND.t2327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1290 VGND.t2273 XThC.XTBN.Y.t57 a_7875_9569# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1292 VPWR.t506 XThR.XTBN.Y XThR.Tn[13].t2 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1293 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t1835 VPWR.t1834 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1294 VPWR.t1272 VPWR.t1270 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1295 VGND.t975 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t974 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1296 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1297 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1298 VPWR.t414 XThR.XTB3.Y.t9 XThR.Tn[10].t3 VPWR.t413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1299 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t142 VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1300 VGND.t1428 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t1427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1301 XThC.Tn[3].t6 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t2253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1303 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t2254 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1304 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t898 VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1305 VGND.t2330 Vbias.t120 XA.XIR[7].XIC[2].icell.SM VGND.t2329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1306 VGND.t2332 Vbias.t121 XA.XIR[6].XIC[3].icell.SM VGND.t2331 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1307 XThR.Tn[5].t10 XThR.XTB6.Y VGND.t2653 VGND.t2465 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1308 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1309 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t2018 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1310 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t190 VGND.t2174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1311 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t254 VGND.t2679 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1312 VPWR.t431 XThR.XTB7.B XThR.XTB4.Y.t0 VPWR.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1313 VGND.t2334 Vbias.t122 XA.XIR[9].XIC[4].icell.SM VGND.t2333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1314 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t984 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t2560 VGND.t2559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 VGND.t2336 Vbias.t123 XA.XIR[14].XIC[10].icell.SM VGND.t2335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1317 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1318 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1991 VGND.t1716 VGND.t1715 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1319 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1320 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t91 VGND.t993 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1321 VGND.t2662 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t2661 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1322 VPWR.t1627 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1323 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t1702 VPWR.t1701 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1324 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t182 VGND.t2048 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1325 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t66 VGND.t682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1326 VGND.t2338 Vbias.t124 XA.XIR[15].XIC[0].icell.SM VGND.t2337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1327 VGND.t2340 Vbias.t125 XA.XIR[14].XIC[1].icell.SM VGND.t2339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1328 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t2114 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1329 VGND.t785 Vbias.t126 XA.XIR[10].XIC[12].icell.SM VGND.t784 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1330 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t131 VGND.t1212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1331 VGND.t608 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t607 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 VGND.t787 Vbias.t127 XA.XIR[13].XIC[13].icell.SM VGND.t786 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1333 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t1676 VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1334 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t541 VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1335 VGND.t645 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1336 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t1444 VGND.t1443 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1337 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1992 VGND.t1714 VGND.t1713 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1338 VGND.t977 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t976 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1339 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t1530 VPWR.t1529 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1340 VGND.t2205 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t2204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1341 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t83 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1342 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t178 VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1343 VPWR.t1704 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1344 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1345 VGND.t789 Vbias.t128 XA.XIR[3].XIC[3].icell.SM VGND.t788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1346 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t345 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1347 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t165 VGND.t1455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1348 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1349 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t39 VGND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1350 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t413 VGND.t412 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1351 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t415 VGND.t414 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t1837 VPWR.t1836 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1353 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1354 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t17 VGND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1355 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t1159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1356 VGND.t2189 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t2188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1357 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t14 VGND.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1358 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t416 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1359 VGND.t1712 VPWR.t1993 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t1711 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1360 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t2255 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1361 XThC.Tn[1].t4 XThC.XTBN.Y.t59 VGND.t2274 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1362 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t2019 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1363 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t236 VGND.t2522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1364 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1365 VPWR.t1269 VPWR.t1267 XA.XIR[15].XIC_15.icell.PUM VPWR.t1268 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1366 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1367 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t2059 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1368 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t992 VPWR.t991 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1369 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t5 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1370 VPWR.t1498 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1497 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1371 VGND.t647 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1372 XA.XIR[15].XIC[14].icell.Ien VPWR.t1264 VPWR.t1266 VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1373 VPWR.t1629 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t1628 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1374 VGND.t2086 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1375 VPWR.t196 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1376 VPWR.t1263 VPWR.t1261 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1377 XThR.Tn[13].t5 XThR.XTB6.Y a_n997_1579# VGND.t2464 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1378 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t4 VPWR.t505 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1379 VPWR.t180 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1380 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1381 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t2497 VGND.t2496 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 VGND.t791 Vbias.t129 XA.XIR[5].XIC[11].icell.SM VGND.t790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1383 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t157 VGND.t1398 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1384 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t1447 VGND.t1446 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1385 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t1862 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1386 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t182 VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1387 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t2123 VGND.t2122 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1388 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t1067 data[2].t1 XThC.XTB7.B VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t2256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1391 VGND.t887 XThR.XTBN.Y XThR.Tn[2].t7 VGND.t886 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1392 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t2499 VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1393 a_n1049_5317# XThR.XTB7.Y VPWR.t1615 VPWR.t1614 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1394 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t2020 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1395 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t238 VGND.t2524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1396 VGND.t2275 XThC.XTBN.Y.t60 XThC.Tn[4].t1 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1397 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t1637 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t419 VGND.t418 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1399 XA.XIR[2].XIC_15.icell.PDM VPWR.t1994 VGND.t1710 VGND.t1709 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1400 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t125 VGND.t1189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1401 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t1638 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1402 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t26 VGND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1404 XThR.Tn[3].t0 XThR.XTB4.Y.t9 VGND.t48 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1405 VPWR.t1494 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1493 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1406 VGND.t2181 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t2180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1407 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t254 VPWR.t253 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1408 VGND.t793 Vbias.t130 XA.XIR[11].XIC[5].icell.SM VGND.t792 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1409 VPWR.t198 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1410 VPWR.t964 XThC.XTB7.Y a_6243_9615# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1411 VPWR.t622 XThC.XTB6.Y XThC.Tn[13].t6 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1412 VPWR.t1260 VPWR.t1258 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1259 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1413 VGND.t795 Vbias.t131 XA.XIR[5].XIC[9].icell.SM VGND.t794 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1414 VGND.t10 data[1].t3 XThC.XTB5.A VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1415 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t2042 VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1416 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1831 VPWR.t1830 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1417 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t403 VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1418 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t2405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1419 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t994 VPWR.t993 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1420 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1255 VPWR.t1257 VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1421 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1631 VPWR.t1630 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 VPWR.t1554 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t1553 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1423 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t2125 VGND.t2124 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1424 VGND.t797 Vbias.t132 XA.XIR[0].XIC[7].icell.SM VGND.t796 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1425 VGND.t2277 XThC.XTBN.Y.t61 XThC.Tn[7].t6 VGND.t2276 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1426 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t2501 VGND.t2500 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1427 VPWR.t1871 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t1870 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1428 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t1448 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1429 XA.XIR[15].XIC[12].icell.PDM VPWR.t1995 XA.XIR[15].XIC[12].icell.Ien VGND.t1708 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1430 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t2044 VGND.t2043 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1431 VGND.t1952 VGND.t1950 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1432 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t123 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1433 XThR.Tn[12].t4 XThR.XTB5.Y VPWR.t1780 VPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1434 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t421 VGND.t420 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1435 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t119 VGND.t1108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1436 a_10915_9569# XThC.XTBN.Y.t62 VGND.t2279 VGND.t2278 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1437 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XThR.Tn[6].t5 XThR.XTBN.Y VGND.t836 VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1439 VPWR.t256 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t255 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1440 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t180 VGND.t2039 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1441 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1442 XThC.Tn[9].t9 XThC.XTB2.Y VPWR.t1767 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1443 VGND.t1573 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1444 VGND.t799 Vbias.t133 XA.XIR[8].XIC[5].icell.SM VGND.t798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1445 VGND.t801 Vbias.t134 XA.XIR[12].XIC[13].icell.SM VGND.t800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1446 VGND.t803 Vbias.t135 XA.XIR[15].XIC[14].icell.SM VGND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1447 a_n997_2667# XThR.XTB4.Y.t10 XThR.Tn[11].t1 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1448 VGND.t2664 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t2663 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1449 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t342 VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1450 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t2258 VGND.t2257 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t313 VPWR.t312 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1452 VGND.t1707 VPWR.t1996 XA.XIR[1].XIC_15.icell.PDM VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1453 VPWR.t1839 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1454 VPWR.t1556 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t1555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1455 VGND.t805 Vbias.t136 XA.XIR[11].XIC[0].icell.SM VGND.t804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1456 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t1706 VPWR.t1705 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1457 VGND.t807 Vbias.t137 XA.XIR[2].XIC_15.icell.SM VGND.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1458 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1252 VPWR.t1254 VPWR.t1253 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1459 VGND.t809 Vbias.t138 XA.XIR[6].XIC[12].icell.SM VGND.t808 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1460 VPWR.t1873 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1872 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1461 XA.XIR[15].XIC[10].icell.PDM VPWR.t1997 XA.XIR[15].XIC[10].icell.Ien VGND.t1705 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1462 VGND.t811 Vbias.t139 XA.XIR[5].XIC[4].icell.SM VGND.t810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1463 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 VGND.t813 Vbias.t140 XA.XIR[9].XIC[13].icell.SM VGND.t812 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1465 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t230 VGND.t2509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1466 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1467 VGND.t733 XThR.XTB7.B a_n1335_8331# VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1468 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t2046 VGND.t2045 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1470 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t405 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1471 VGND.t1054 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1472 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t178 VGND.t2037 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1473 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t1591 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1474 VPWR.t1696 XThC.XTBN.Y.t63 XThC.Tn[9].t1 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1475 XA.XIR[15].XIC_15.icell.PUM VPWR.t1250 XA.XIR[15].XIC_15.icell.Ien VPWR.t1251 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1476 a_10051_9569# XThC.XTBN.Y.t64 VGND.t2280 VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1477 VGND.t1430 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t1429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1478 VPWR.t504 XThR.XTBN.Y XThR.Tn[7].t1 VPWR.t503 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1479 VGND.t815 Vbias.t141 XA.XIR[0].XIC[2].icell.SM VGND.t814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1480 VPWR.t258 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t257 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1481 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1641 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1482 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1248 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1249 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1483 VPWR.t1532 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t1531 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1484 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t1854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1485 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t1853 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1486 XThC.Tn[11].t0 XThC.XTB4.Y.t8 VPWR.t17 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1487 VGND.t885 XThR.XTBN.Y XThR.Tn[1].t2 VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1488 XThR.Tn[1].t5 XThR.XTBN.Y a_n1049_7787# VPWR.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1489 a_7651_9569# XThC.XTBN.Y.t65 VGND.t2281 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1490 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1491 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1633 VPWR.t1632 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1492 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1493 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t1544 VPWR.t1543 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1494 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t1998 VGND.t1704 VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1495 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t176 VGND.t1555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1496 VPWR.t260 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t259 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1497 VPWR.t1708 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t1707 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1498 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t2047 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1499 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t1135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XThR.Tn[6].t9 XThR.XTB7.Y VGND.t2113 VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1501 a_n1049_5611# XThR.XTB6.Y VPWR.t1903 VPWR.t1614 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 XThR.Tn[9].t8 XThR.XTB2.Y VPWR.t1014 VPWR.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 VPWR.t1247 VPWR.t1245 XA.XIR[11].XIC_15.icell.PUM VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1504 VGND.t817 Vbias.t142 XA.XIR[8].XIC[0].icell.SM VGND.t816 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1505 VGND.t819 Vbias.t143 XA.XIR[3].XIC[12].icell.SM VGND.t818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1506 VGND.t1949 VGND.t1947 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1507 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t89 VGND.t991 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1508 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1509 XThC.Tn[4].t0 XThC.XTBN.Y.t66 VGND.t2282 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1510 VGND.t649 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t2260 VGND.t2259 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t344 VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1513 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t1908 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 VPWR.t502 XThR.XTBN.Y XThR.Tn[13].t1 VPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1515 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t2022 VGND.t2021 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1516 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1492 VPWR.t1491 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1517 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t545 VGND.t544 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1518 VPWR.t1558 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t1557 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t1702 VPWR.t1999 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t1875 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1874 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t1534 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t1533 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1642 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t82 VGND.t950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1525 VGND.t2680 XThR.XTB1.Y.t11 XThR.Tn[0].t11 VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1526 XThR.Tn[5].t5 XThR.XTBN.Y VGND.t884 VGND.t868 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t1944 VGND.t1946 VGND.t1945 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t1941 VGND.t1943 VGND.t1942 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t731 XThR.XTB7.B XThR.XTB6.Y VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t223 VGND.t2406 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1532 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t683 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1534 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t423 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1535 VGND.t2283 XThC.XTBN.Y.t67 XThC.Tn[0].t5 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1536 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t1710 VPWR.t1709 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t1546 VPWR.t1545 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1538 VGND.t2191 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t2190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t1700 VPWR.t2000 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t1699 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t2183 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t978 XThC.XTBN.Y.t68 XThC.Tn[3].t3 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t2236 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t2235 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1543 VGND.t1294 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t1293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VPWR.t1536 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t1535 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1545 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t1852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1546 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2001 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t1698 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XThC.Tn[7].t5 XThC.XTBN.Y.t69 VGND.t980 VGND.t979 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1549 VPWR.t607 XThC.XTBN.Y.t70 XThC.Tn[12].t1 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1550 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t769 VPWR.t768 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1551 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t266 VPWR.t265 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1552 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1242 VPWR.t1244 VPWR.t1243 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 VGND.t84 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t83 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1554 VGND.t722 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1555 VPWR.t1013 XThR.XTB2.Y a_n1049_7787# VPWR.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1556 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t1548 VPWR.t1547 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1557 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t2024 VGND.t2023 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t184 VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1559 VGND.t982 XThC.XTBN.Y.t71 a_10915_9569# VGND.t981 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1560 VPWR.t565 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t564 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1561 VPWR.t315 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1562 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1563 VPWR.t1490 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1489 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1564 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2002 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t1697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1565 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t996 VPWR.t995 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 XThC.Tn[11].t1 XThC.XTB4.Y.t9 a_8963_9569# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VGND.t821 Vbias.t144 XA.XIR[2].XIC[8].icell.SM VGND.t820 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1568 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t2029 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1569 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2003 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t1696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t268 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 VGND.t17 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1572 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t224 VGND.t2407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XThR.Tn[14].t3 XThR.XTBN.Y VPWR.t501 VPWR.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1574 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t220 VGND.t2402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1575 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t1773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1576 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1240 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1241 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1577 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t86 VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1578 a_7875_9569# XThC.XTBN.Y.t72 VGND.t983 VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t1571 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1580 VPWR.t1902 XThR.XTB6.Y XThR.Tn[13].t11 VPWR.t1608 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t985 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t1851 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1583 VGND.t823 Vbias.t145 XA.XIR[10].XIC[6].icell.SM VGND.t822 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1584 XA.XIR[0].XIC[3].icell.PDM VGND.t1938 VGND.t1940 VGND.t1939 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1585 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2004 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t1695 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1586 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1587 XThC.Tn[11].t10 XThC.XTB4.Y.t11 a_8963_9569# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1588 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t200 VPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1589 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t270 VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1590 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1238 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1239 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1591 XThC.Tn[0].t10 XThC.XTB1.Y.t12 VGND.t1091 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1592 VGND.t825 Vbias.t146 XA.XIR[1].XIC_15.icell.SM VGND.t824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1593 VGND.t985 XThC.XTBN.Y.t73 a_10051_9569# VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1594 VGND.t2382 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t2381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1595 VPWR.t317 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t316 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1596 VGND.t2185 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t2184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1597 XThR.XTB1.Y.t2 XThR.XTB5.A VPWR.t1919 VPWR.t1918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1598 VPWR.t567 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1599 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1600 XThR.Tn[13].t4 XThR.XTB6.Y a_n997_1579# VGND.t2463 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1601 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1602 VGND.t827 Vbias.t147 XA.XIR[11].XIC[14].icell.SM VGND.t826 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1603 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t1592 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1604 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2005 VGND.t1694 VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 VGND.t2555 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t2554 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1606 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1607 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t2549 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1608 VGND.t986 XThC.XTBN.Y.t74 a_7651_9569# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1877 VPWR.t1876 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1610 XThC.XTBN.Y.t2 XThC.XTBN.A VGND.t1214 VGND.t1213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1611 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t319 VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1612 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1235 VPWR.t1237 VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1613 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t2506 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1614 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t2507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1615 VGND.t829 Vbias.t148 XA.XIR[2].XIC[3].icell.SM VGND.t828 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1616 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t1062 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1617 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t2030 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1618 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t246 VGND.t2588 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1619 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1620 VGND.t1937 VGND.t1935 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1936 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1621 VGND.t831 Vbias.t149 XA.XIR[14].XIC[7].icell.SM VGND.t830 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1622 VGND.t2411 Vbias.t150 XA.XIR[10].XIC[10].icell.SM VGND.t2410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1623 XA.XIR[0].XIC[7].icell.PDM VGND.t1932 VGND.t1934 VGND.t1933 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1624 a_n1049_5317# XThR.XTBN.Y XThR.Tn[6].t2 VPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1625 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t1151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2006 VGND.t1692 VGND.t1691 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1627 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t694 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1628 VPWR.t609 XThC.XTBN.Y.t75 XThC.Tn[7].t0 VPWR.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 VPWR.t1488 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1487 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1630 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t1153 VGND.t1152 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 XA.XIR[15].XIC[8].icell.Ien VPWR.t1232 VPWR.t1234 VPWR.t1233 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1632 VPWR.t272 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t271 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1633 VGND.t883 XThR.XTBN.Y a_n997_1803# VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1634 VPWR.t1678 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1635 XThR.Tn[3].t8 XThR.XTBN.Y VGND.t881 VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1636 VGND.t1569 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t1568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1637 VPWR.t406 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1638 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t159 VGND.t1437 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1639 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t225 VGND.t2408 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1640 VGND.t2413 Vbias.t151 XA.XIR[10].XIC[1].icell.SM VGND.t2412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1641 VGND.t2415 Vbias.t152 XA.XIR[5].XIC[13].icell.SM VGND.t2414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1642 VPWR.t1924 XThC.XTB4.Y.t12 XThC.Tn[11].t11 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t1909 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t547 VGND.t546 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1646 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t1841 VPWR.t1840 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1647 VGND.t2088 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1648 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t1155 VGND.t1154 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 VGND.t2417 Vbias.t153 XA.XIR[8].XIC[14].icell.SM VGND.t2416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t425 VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1879 VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 VGND.t1690 VPWR.t2007 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t1689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1653 XThC.Tn[0].t4 XThC.XTBN.Y.t76 VGND.t987 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1654 VPWR.t321 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1655 VGND.t2419 Vbias.t154 XA.XIR[4].XIC[11].icell.SM VGND.t2418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1656 XThC.Tn[3].t2 XThC.XTBN.Y.t77 VGND.t988 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1657 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t84 VGND.t954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 VGND.t86 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1659 VGND.t724 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t723 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t684 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1662 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1663 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[8].XIC_15.icell.PUM VPWR.t1230 XA.XIR[8].XIC_15.icell.Ien VPWR.t1231 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t291 VPWR.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1667 VGND.t610 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1668 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t712 VGND.t711 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 VPWR.t1229 VPWR.t1227 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1228 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1670 VGND.t2238 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t2237 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1671 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t2508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1672 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t123 VGND.t1187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1673 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t262 VPWR.t261 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1674 VPWR.t1680 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1675 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1676 VGND.t2421 Vbias.t155 XA.XIR[14].XIC[2].icell.SM VGND.t2420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1677 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t906 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1678 XThC.XTB1.Y.t2 XThC.XTB5.A a_3299_10575# VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1679 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t323 VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1680 VPWR.t1486 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1485 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1681 VGND.t2370 XThR.XTB3.Y.t10 XThR.Tn[2].t11 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1682 XA.XIR[15].XIC[3].icell.Ien VPWR.t1224 VPWR.t1226 VPWR.t1225 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1683 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t1157 VGND.t1156 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1684 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t771 VPWR.t770 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1685 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t986 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1686 VPWR.t274 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1687 VGND.t2423 Vbias.t156 XA.XIR[1].XIC[8].icell.SM VGND.t2422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1688 VPWR.t798 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t797 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t626 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t625 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1691 VGND.t2425 Vbias.t157 XA.XIR[4].XIC[9].icell.SM VGND.t2424 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1692 VPWR.t741 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t740 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1693 VPWR.t408 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t108 VGND.t1066 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1695 VGND.t1931 VGND.t1929 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1930 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1696 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t194 VGND.t2350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1697 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t166 VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 VGND.t990 XThC.XTBN.Y.t78 XThC.Tn[6].t6 VGND.t989 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1699 XThC.Tn[10].t4 XThC.XTB3.Y.t11 VPWR.t695 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1700 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t239 VGND.t2525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1701 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t427 VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1702 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t1850 VGND.t1849 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1703 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t743 VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1704 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t93 VGND.t995 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1705 XThC.Tn[14].t10 XThC.XTB7.Y VPWR.t963 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t1174 VGND.t1173 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t1688 VPWR.t2008 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t1687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t749 XThC.XTB1.Y.t13 XThC.Tn[0].t8 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t8 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1711 VGND.t2557 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t2556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t1774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t33 VGND.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1715 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t186 VGND.t2060 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1716 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1717 XThR.Tn[8].t4 XThR.XTBN.Y VPWR.t500 VPWR.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1718 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t619 VGND.t618 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1719 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t621 VGND.t620 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 VGND.t2384 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t2383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t2187 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t2186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t264 VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1723 VGND.t1370 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t1369 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1724 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t202 VPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1725 VGND.t2427 Vbias.t158 XA.XIR[7].XIC[5].icell.SM VGND.t2426 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 VGND.t1296 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t1295 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1727 VGND.t2429 Vbias.t159 XA.XIR[6].XIC[6].icell.SM VGND.t2428 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t1686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y XThR.Tn[5].t1 VPWR.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t325 VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t1121 VGND.t1120 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t85 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t1848 VGND.t1847 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1734 XThR.XTBN.A data[7].t1 VGND.t1111 VGND.t1110 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1735 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t276 VPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1736 VGND.t2431 Vbias.t160 XA.XIR[1].XIC[3].icell.SM VGND.t2430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1737 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1738 XThC.Tn[14].t9 XThC.XTB7.Y VPWR.t962 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1739 VGND.t2433 Vbias.t161 XA.XIR[4].XIC[4].icell.SM VGND.t2432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1740 VPWR.t353 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t1158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t365 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t569 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2010 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t1685 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t2090 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t1137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 XThC.XTB2.Y XThC.XTB7.B VPWR.t107 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t171 VGND.t1522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1749 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1895 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t628 VPWR.t627 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t181 VGND.t2040 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1752 XThR.Tn[5].t4 XThR.XTBN.Y VGND.t880 VGND.t859 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1753 VGND.t1432 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t1431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t349 VGND.t348 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1755 VGND.t1567 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t1566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t5 XThR.XTBN.Y VPWR.t497 VPWR.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t204 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t203 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t1565 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t1564 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# XThC.XTB6.Y VPWR.t621 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t2435 Vbias.t162 XA.XIR[6].XIC[10].icell.SM VGND.t2434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t2437 Vbias.t163 XA.XIR[3].XIC[6].icell.SM VGND.t2436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t351 VGND.t350 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1763 VPWR.t696 XThC.XTB3.Y.t12 XThC.Tn[10].t5 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1764 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t623 VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1765 XThC.Tn[13].t0 XThC.XTBN.Y.t79 VPWR.t1072 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1766 XA.XIR[13].XIC_15.icell.PDM VPWR.t2011 VGND.t1684 VGND.t1683 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1767 a_n997_3755# XThR.XTBN.Y VGND.t879 VGND.t865 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1768 VGND.t2439 Vbias.t164 XA.XIR[7].XIC[0].icell.SM VGND.t2438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1769 VGND.t2441 Vbias.t165 XA.XIR[2].XIC[12].icell.SM VGND.t2440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1770 VGND.t2443 Vbias.t166 XA.XIR[6].XIC[1].icell.SM VGND.t2442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1771 VPWR.t495 XThR.XTBN.Y XThR.Tn[14].t2 VPWR.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1772 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1773 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t714 VGND.t713 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1774 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t1593 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1775 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t1123 VGND.t1122 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t13 VGND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1777 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t1864 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2012 VGND.t1682 VGND.t1681 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 VPWR.t355 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1780 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1781 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t630 VPWR.t629 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1782 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t214 VGND.t2396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1783 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1784 XThR.Tn[7].t4 XThR.XTBN.Y VGND.t878 VGND.t877 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1785 VPWR.t1223 VPWR.t1221 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1786 VGND.t1434 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t1433 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1787 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t174 VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1788 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t347 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1789 VGND.t1680 VPWR.t2013 XA.XIR[15].XIC_15.icell.PDM VGND.t1679 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1790 XThC.XTB4.Y.t1 XThC.XTB7.B VGND.t128 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1791 VPWR.t1901 XThR.XTB6.Y XThR.Tn[13].t10 VPWR.t1616 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1792 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t147 VGND.t1334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1793 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t233 VGND.t2512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1794 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1882 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1795 VGND.t2445 Vbias.t167 XA.XIR[3].XIC[10].icell.SM VGND.t2444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1796 VPWR.t776 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t775 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1797 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t2393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1798 VPWR.t134 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1799 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t278 VPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1800 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t800 VPWR.t799 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 VPWR.t616 data[4].t3 XThR.XTB7.A VPWR.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1802 VGND.t2193 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t2192 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1803 VGND.t1678 VPWR.t2014 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t1677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2015 VGND.t1676 VGND.t1675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1805 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t353 VGND.t352 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XThC.Tn[6].t5 XThC.XTBN.Y.t80 VGND.t1541 VGND.t1540 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1807 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t625 VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 VGND.t1928 VGND.t1926 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1927 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1809 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t1538 VPWR.t1537 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1810 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t410 VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 VPWR.t571 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1812 VPWR.t327 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 XThR.Tn[5].t9 XThR.XTB6.Y VGND.t2652 VGND.t2461 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1814 VPWR.t458 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1815 VPWR.t1684 XThC.XTB5.Y a_5155_9615# VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1816 VPWR.t1220 VPWR.t1218 XA.XIR[3].XIC_15.icell.PUM VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1817 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1818 VPWR.t1217 VPWR.t1215 XA.XIR[7].XIC_15.icell.PUM VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1819 VGND.t2447 Vbias.t168 XA.XIR[3].XIC[1].icell.SM VGND.t2446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1820 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t94 VGND.t996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t1910 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t10 XThR.XTB5.Y VGND.t2466 VGND.t2465 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1925 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t5 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t1176 VGND.t1175 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1826 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t227 VGND.t2458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1827 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t179 VGND.t2038 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1828 VGND.t1674 VPWR.t2016 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t1673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1829 VGND.t1542 XThC.XTBN.Y.t82 XThC.Tn[2].t5 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t1672 VPWR.t2017 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t1671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 VPWR.t438 XThC.XTB1.Y.t14 XThC.Tn[8].t9 VPWR.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1832 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t206 VGND.t2371 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1833 VGND.t2666 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t2665 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# XThC.XTBN.Y.t83 VGND.t1544 VGND.t1543 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t176 VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t930 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t145 VGND.t1324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1839 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1840 VPWR.t778 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t777 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1841 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t68 VGND.t698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1842 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t632 VPWR.t631 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1843 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1844 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1845 VGND.t2449 Vbias.t169 XA.XIR[13].XIC_15.icell.SM VGND.t2448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t802 VPWR.t801 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1847 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t2687 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1848 VGND.t2195 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t2194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 VGND.t1326 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t1325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1850 VGND.t2573 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t2572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t1540 VPWR.t1539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1852 VGND.t1056 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1853 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t227 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1854 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t127 VGND.t1199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1855 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t1021 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1856 XThR.Tn[3].t7 XThR.XTBN.Y VGND.t876 VGND.t875 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1857 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t908 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1858 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t280 VPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t804 VPWR.t803 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1213 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1214 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t252 VGND.t2656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1862 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t5 VGND.t1406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1863 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t1542 VPWR.t1541 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1864 a_4387_10575# XThC.XTB7.B VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1865 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t745 VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t412 VPWR.t411 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t573 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t150 VPWR.t149 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t1138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1871 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2018 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t1670 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t1177 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t2025 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t103 VGND.t1019 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1876 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t1086 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1877 a_10051_9569# XThC.XTBN.Y.t84 VGND.t1545 VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1878 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t137 VGND.t1230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1879 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1880 XThC.XTB1.Y.t0 XThC.XTB7.B VPWR.t106 VPWR.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1881 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t4 VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1882 VGND.t1925 VGND.t1923 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1210 VPWR.t1212 VPWR.t1211 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 a_n1049_8581# XThR.XTBN.Y XThR.Tn[0].t3 VPWR.t493 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1885 a_7651_9569# XThC.XTBN.Y.t85 VGND.t1546 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1886 VGND.t651 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1887 VPWR.t1833 XThC.XTB7.A a_6243_10571# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1888 VPWR.t1209 VPWR.t1207 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1208 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1889 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t250 VGND.t2650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1890 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t1016 VGND.t1015 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1891 VPWR.t670 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t669 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1892 XThC.Tn[10].t8 XThC.XTB3.Y.t13 a_8739_9569# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1893 VGND.t2386 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t2385 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1894 VGND.t2451 Vbias.t170 XA.XIR[1].XIC[12].icell.SM VGND.t2450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 VGND.t874 XThR.XTBN.Y XThR.Tn[2].t6 VGND.t873 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1896 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t1140 VGND.t1139 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t1142 VGND.t1141 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1898 XThR.XTB5.A data[5].t3 VGND.t946 VGND.t945 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1899 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1205 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1206 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 VGND.t2453 Vbias.t171 XA.XIR[0].XIC[5].icell.SM VGND.t2452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1901 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1902 VGND.t2455 Vbias.t172 XA.XIR[4].XIC[13].icell.SM VGND.t2454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1903 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1904 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t1023 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1905 XThR.Tn[12].t1 XThR.XTBN.Y VPWR.t492 VPWR.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 VGND.t1669 VPWR.t2019 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t1668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1907 VGND.t2457 Vbias.t173 XA.XIR[7].XIC[14].icell.SM VGND.t2456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1908 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t551 VGND.t550 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1910 XThR.Tn[12].t9 XThR.XTB5.Y a_n997_1803# VGND.t2464 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1911 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1912 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t939 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1913 XThR.Tn[3].t1 XThR.XTB4.Y.t11 VGND.t51 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1914 VGND.t872 XThR.XTBN.Y a_n997_2667# VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1915 XA.XIR[9].XIC_15.icell.PDM VPWR.t2020 VGND.t1667 VGND.t1666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1916 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t1178 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1917 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1202 VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1918 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t367 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1919 VGND.t726 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t725 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1920 VGND.t1342 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t1341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1921 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t2026 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1922 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t31 VGND.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1923 a_5155_9615# XThC.XTB5.Y VPWR.t1683 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1924 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t1124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1925 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1926 VGND.t2127 Vbias.t174 XA.XIR[10].XIC[7].icell.SM VGND.t2126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1927 VPWR.t1682 XThC.XTB5.Y XThC.Tn[12].t4 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1928 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t172 VGND.t1526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1929 VPWR.t220 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t219 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1930 XA.XIR[7].XIC_15.icell.PUM VPWR.t1200 XA.XIR[7].XIC_15.icell.Ien VPWR.t1201 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1931 VPWR.t636 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t635 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1932 VGND.t2129 Vbias.t175 XA.XIR[13].XIC[8].icell.SM VGND.t2128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1933 VPWR.t1199 VPWR.t1197 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1198 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1934 VGND.t1436 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t1435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1935 XThC.Tn[5].t4 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1936 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t766 VGND.t765 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1937 VGND.t2261 XThC.XTB5.Y XThC.Tn[4].t8 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1938 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t5 VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1939 VPWR.t723 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t722 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1940 VPWR.t634 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t633 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1941 XThC.Tn[2].t4 XThC.XTBN.Y.t87 VGND.t1547 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1942 VPWR.t747 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t746 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1943 XA.XIR[15].XIC[14].icell.PDM VPWR.t2021 XA.XIR[15].XIC[14].icell.Ien VGND.t1665 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1944 XA.XIR[15].XIC[8].icell.PDM VPWR.t2022 XA.XIR[15].XIC[8].icell.Ien VGND.t1664 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1945 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t9 VGND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1946 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1018 VGND.t1017 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1947 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t5 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1948 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t768 VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1949 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t987 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1950 VPWR.t429 XThR.XTB7.B XThR.XTB2.Y VPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1951 XThC.Tn[8].t4 XThC.XTB1.Y.t15 a_7651_9569# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1952 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t684 VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1953 VGND.t2668 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t2667 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1954 XA.XIR[6].XIC_15.icell.PDM VPWR.t2023 VGND.t1663 VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1955 VGND.t1441 XThC.XTB5.A XThC.XTB5.Y VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1956 VGND.t2131 Vbias.t176 XA.XIR[0].XIC[0].icell.SM VGND.t2130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1957 VGND.t2111 XThR.XTB7.Y XThR.Tn[6].t8 VGND.t2110 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1958 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t1241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1959 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t1588 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t1866 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1961 VGND.t2133 Vbias.t177 XA.XIR[12].XIC_15.icell.SM VGND.t2132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1962 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t130 VGND.t1211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1963 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t553 VGND.t552 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1964 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1096 VGND.t1095 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1965 VPWR.t222 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t221 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1966 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1967 XA.XIR[4].XIC_15.icell.PUM VPWR.t1195 XA.XIR[4].XIC_15.icell.Ien VPWR.t1196 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t1243 VGND.t1242 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1969 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2024 VGND.t1661 VGND.t1660 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[15].XIC[9].icell.Ien VPWR.t1192 VPWR.t1194 VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1971 VGND.t1058 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1057 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1972 XThR.Tn[9].t0 XThR.XTBN.Y VPWR.t486 VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1973 VGND.t1548 XThC.XTBN.Y.t89 a_9827_9569# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1974 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t931 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1975 VPWR.t725 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1976 VGND.t2216 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1977 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t92 VGND.t994 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1978 VGND.t1659 VPWR.t2025 XA.XIR[8].XIC_15.icell.PDM VGND.t1658 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 VPWR.t864 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t863 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1980 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t224 VPWR.t223 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1981 VGND.t2135 Vbias.t178 XA.XIR[10].XIC[2].icell.SM VGND.t2134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1982 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t56 VGND.t656 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1983 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1189 VPWR.t1191 VPWR.t1190 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1984 VGND.t2137 Vbias.t179 XA.XIR[9].XIC_15.icell.SM VGND.t2136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1985 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t2471 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1986 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1187 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1188 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1987 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t129 VGND.t1210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1988 XThC.Tn[0].t9 XThC.XTB1.Y.t16 VGND.t750 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1989 VGND.t2139 Vbias.t180 XA.XIR[13].XIC[3].icell.SM VGND.t2138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1990 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t2472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1991 VGND.t2197 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t2196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1992 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t8 VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1993 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t770 VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1994 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1484 VPWR.t1483 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1995 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t282 VPWR.t281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1996 VPWR.t727 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t726 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1997 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t686 VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1998 VGND.t1298 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t1297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1999 VPWR.t1843 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t1842 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2000 XThR.Tn[14].t1 XThR.XTBN.Y VPWR.t489 VPWR.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2001 VPWR.t850 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t849 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 VPWR.t1186 VPWR.t1184 XA.XIR[0].XIC_15.icell.PUM VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2003 VPWR.t638 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t637 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2004 XA.XIR[15].XIC[3].icell.PDM VPWR.t2026 XA.XIR[15].XIC[3].icell.Ien VGND.t1657 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2005 a_n997_3755# XThR.XTBN.Y VGND.t870 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2006 XThR.Tn[8].t2 XThR.XTB1.Y.t13 VPWR.t293 VPWR.t292 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2007 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t174 VGND.t1528 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2008 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2009 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t76 VGND.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2010 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t1845 VPWR.t1844 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2011 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1098 VGND.t1097 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2012 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t167 VGND.t1457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2013 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t47 VGND.t562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2014 a_n1049_7787# XThR.XTB2.Y VPWR.t1012 VPWR.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2015 VGND.t653 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2016 VPWR.t1788 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t1787 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2017 a_n1331_2891# data[5].t4 VGND.t207 VGND.t206 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2018 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t1790 VPWR.t1789 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2019 VPWR.t1183 VPWR.t1181 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1182 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2020 VGND.t2092 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2021 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t74 VGND.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2022 VPWR.t226 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t225 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2023 VGND.t2141 Vbias.t181 XA.XIR[15].XIC[11].icell.SM VGND.t2140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2024 XThR.XTB7.B data[6].t1 VGND.t1268 VGND.t1267 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2025 XThR.Tn[2].t3 XThR.XTBN.Y a_n1049_7493# VPWR.t487 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2026 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t589 VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2027 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t591 VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2028 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1482 VPWR.t1481 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2029 VGND.t1372 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t1371 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2030 VGND.t2143 Vbias.t182 XA.XIR[2].XIC[6].icell.SM VGND.t2142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2031 VGND.t1486 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t1485 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2027 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2033 XA.XIR[15].XIC[7].icell.PDM VPWR.t2028 XA.XIR[15].XIC[7].icell.Ien VGND.t1655 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2034 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t2473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2035 VPWR.t370 XThC.XTBN.Y.t90 XThC.Tn[8].t2 VPWR.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2036 XThR.Tn[10].t1 XThR.XTB3.Y.t12 VPWR.t144 VPWR.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2037 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t771 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2038 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t735 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2039 XThR.Tn[4].t1 XThR.XTBN.Y VGND.t869 VGND.t868 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2040 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t952 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2041 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1179 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2042 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1480 VPWR.t1479 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2043 VGND.t730 XThR.XTB7.B XThR.XTB5.Y VGND.t729 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2044 VGND.t2078 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2045 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2046 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t228 VPWR.t227 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2047 VGND.t1344 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2048 VPWR.t640 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t639 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2049 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2050 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t1846 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2051 VPWR.t1792 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t1791 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2052 VPWR.t329 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2053 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t554 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2054 VGND.t2145 Vbias.t183 XA.XIR[12].XIC[8].icell.SM VGND.t2144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2055 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2056 VPWR.t672 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t671 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2057 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t5 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2058 XThC.Tn[4].t4 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2059 VGND.t2147 Vbias.t184 XA.XIR[15].XIC[9].icell.SM VGND.t2146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2060 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t1043 VPWR.t1042 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2061 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1176 VPWR.t1178 VPWR.t1177 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2062 VGND.t1563 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t1562 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2063 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t2515 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2064 VPWR.t152 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2065 VGND.t867 XThR.XTBN.Y a_n997_1579# VGND.t849 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2066 VGND.t2149 Vbias.t185 XA.XIR[2].XIC[10].icell.SM VGND.t2148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2067 VPWR.t389 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t388 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2068 VGND.t2151 Vbias.t186 XA.XIR[6].XIC[7].icell.SM VGND.t2150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2069 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2029 VGND.t1654 VGND.t1653 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2070 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2071 VGND.t2153 Vbias.t187 XA.XIR[9].XIC[8].icell.SM VGND.t2152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2072 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2073 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1894 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2074 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t593 VGND.t592 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2075 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t9 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2076 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t65 VGND.t681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2077 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t1775 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2078 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1174 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1175 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 VGND.t2155 Vbias.t188 XA.XIR[2].XIC[1].icell.SM VGND.t2154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2080 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t185 VGND.t2052 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2081 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t1911 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2082 VGND.t2157 Vbias.t189 XA.XIR[0].XIC[14].icell.SM VGND.t2156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2083 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t1245 VGND.t1244 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2084 VGND.t2159 Vbias.t190 XA.XIR[14].XIC[5].icell.SM VGND.t2158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2085 XA.XIR[0].XIC[5].icell.PDM VGND.t1920 VGND.t1922 VGND.t1921 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2086 VPWR.t331 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2087 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t233 VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2088 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t1042 VGND.t1041 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 VGND.t2218 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2090 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t230 VPWR.t229 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2091 XThR.XTBN.Y XThR.XTBN.A VPWR.t542 VPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2092 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1045 VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2093 VPWR.t156 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2094 VGND.t2080 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t2516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2096 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t686 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2097 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t1845 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2098 VGND.t1346 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t1345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2099 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1171 VPWR.t1173 VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2100 VPWR.t391 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t390 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2101 VGND.t2161 Vbias.t191 XA.XIR[3].XIC[7].icell.SM VGND.t2160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2102 VGND.t2163 Vbias.t192 XA.XIR[12].XIC[3].icell.SM VGND.t2162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2103 XA.XIR[0].XIC_15.icell.PUM VPWR.t1169 XA.XIR[0].XIC_15.icell.Ien VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2104 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2105 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t729 VPWR.t728 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2106 VGND.t1328 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t1327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2107 VGND.t2575 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t2574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 VGND.t2165 Vbias.t193 XA.XIR[15].XIC[4].icell.SM VGND.t2164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2109 VPWR.t485 XThR.XTBN.Y XThR.Tn[11].t5 VPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2110 VGND.t1919 VGND.t1917 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1918 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2111 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t852 VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2112 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t595 VGND.t594 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2113 VPWR.t100 data[1].t4 XThC.XTB7.A VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2114 VPWR.t154 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t153 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2115 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t674 VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2116 a_8739_9569# XThC.XTBN.Y.t92 VGND.t661 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2117 VGND.t2167 Vbias.t194 XA.XIR[6].XIC[2].icell.SM VGND.t2166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2118 VGND.t940 XThR.XTBN.A XThR.XTBN.Y VGND.t939 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2119 XThC.Tn[6].t10 XThC.XTB7.Y VGND.t1405 VGND.t1404 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2120 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t3 VGND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2121 VGND.t2169 Vbias.t195 XA.XIR[9].XIC[3].icell.SM VGND.t2168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2122 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t1257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2123 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t1258 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2124 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2125 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t2518 VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2126 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1038 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2127 XThR.Tn[12].t8 XThR.XTB5.Y a_n997_1803# VGND.t2463 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2128 VGND.t1652 VPWR.t2030 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t1651 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 VGND.t2063 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t2062 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2130 VGND.t2208 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t2207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2131 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t49 VGND.t564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2132 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t203 VGND.t2366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2133 a_n997_3979# XThR.XTBN.Y VGND.t866 VGND.t865 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2134 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t43 VGND.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2135 VGND.t2171 Vbias.t196 XA.XIR[14].XIC[0].icell.SM VGND.t2170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2136 XThC.XTB7.Y XThC.XTB7.B VGND.t125 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2137 XA.XIR[0].XIC[0].icell.PDM VGND.t1914 VGND.t1916 VGND.t1915 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2138 VGND.t2173 Vbias.t197 XA.XIR[5].XIC_15.icell.SM VGND.t2172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2139 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1166 VPWR.t1168 VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2140 VGND.t137 Vbias.t198 XA.XIR[13].XIC[12].icell.SM VGND.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2141 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t780 VPWR.t779 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2142 XThC.Tn[8].t1 XThC.XTBN.Y.t93 VPWR.t372 VPWR.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2143 VGND.t1330 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t1329 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2144 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t1044 VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2145 VGND.t1060 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t1059 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2147 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t866 VPWR.t865 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2148 VGND.t139 Vbias.t199 XA.XIR[1].XIC[6].icell.SM VGND.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2149 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2031 VGND.t1650 VGND.t1649 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2150 VGND.t2220 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t2219 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2151 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t1179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2152 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t676 VPWR.t675 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2153 a_n1049_6699# XThR.XTB4.Y.t12 VPWR.t1524 VPWR.t1523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2154 VPWR.t393 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2155 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2156 VGND.t141 Vbias.t200 XA.XIR[3].XIC[2].icell.SM VGND.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2157 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t736 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2158 VGND.t143 Vbias.t201 XA.XIR[11].XIC[11].icell.SM VGND.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2159 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t782 VPWR.t781 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2160 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1164 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2161 VGND.t2388 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t2387 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2162 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t105 VGND.t1030 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2163 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1162 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2164 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t854 VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2165 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t96 VGND.t1001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2166 VGND.t1488 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t1487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2167 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2168 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2169 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t1163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2170 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t1171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2171 VGND.t1647 VPWR.t2033 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2172 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t150 VGND.t1368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2174 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2175 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2176 VGND.t428 data[1].t5 XThC.XTB6.A VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2177 VPWR.t232 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t231 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2178 VPWR.t1161 VPWR.t1159 XA.XIR[14].XIC_15.icell.PUM VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2179 a_n997_2891# XThR.XTBN.Y VGND.t864 VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2180 VGND.t1913 VGND.t1911 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2181 VGND.t655 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2182 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2183 VGND.t145 Vbias.t202 XA.XIR[1].XIC[10].icell.SM VGND.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2184 VPWR.t784 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t783 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2185 VPWR.t1158 VPWR.t1156 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2186 VGND.t2210 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2187 VPWR.t1155 VPWR.t1153 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1154 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t193 VGND.t2349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2189 VPWR.t1794 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t1793 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2190 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2034 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t1645 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2191 XThR.Tn[11].t8 XThR.XTB4.Y.t13 a_n997_2667# VGND.t2016 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2192 VGND.t147 Vbias.t203 XA.XIR[11].XIC[9].icell.SM VGND.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2193 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t557 VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2194 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t112 VGND.t1088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2195 VGND.t149 Vbias.t204 XA.XIR[8].XIC[11].icell.SM VGND.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2196 VPWR.t1681 XThC.XTB5.Y a_5155_9615# VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2197 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t1776 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2198 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t1844 VGND.t1843 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2199 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t1842 VGND.t1841 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2200 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2201 VGND.t151 Vbias.t205 XA.XIR[1].XIC[1].icell.SM VGND.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2202 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t1172 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2203 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1004 VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2204 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t236 VGND.t235 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2205 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2206 VGND.t2577 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t2576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2207 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t1260 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2208 VGND.t862 XThR.XTBN.Y XThR.Tn[0].t7 VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2209 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t559 VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2210 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t940 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2211 a_n1049_6405# XThR.XTB5.Y VPWR.t1779 VPWR.t1523 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2212 XThR.Tn[8].t7 XThR.XTB1.Y.t14 VPWR.t546 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2213 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t111 VGND.t1087 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2214 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t953 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2215 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2216 XA.XIR[5].XIC_15.icell.PDM VPWR.t2035 VGND.t1644 VGND.t1643 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2217 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t128 VGND.t1205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2218 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t1028 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2219 VGND.t1348 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 VGND.t2082 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2221 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2222 XThR.Tn[1].t9 XThR.XTB2.Y VGND.t1466 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2223 VGND.t2084 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2224 VGND.t1350 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2225 VPWR.t786 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t785 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2226 VGND.t662 XThC.XTBN.Y.t94 a_8739_9569# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2227 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t234 VPWR.t233 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2228 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t139 VGND.t1266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2229 VPWR.t1152 VPWR.t1150 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2230 XThC.Tn[1].t10 XThC.XTB2.Y VGND.t2378 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2231 VGND.t1403 XThC.XTB7.Y XThC.Tn[6].t9 VGND.t1402 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2232 VGND.t153 Vbias.t206 XA.XIR[5].XIC[8].icell.SM VGND.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2233 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2036 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2234 VPWR.t333 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2235 VPWR.t1149 VPWR.t1147 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1148 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t1 VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2237 VGND.t155 Vbias.t207 XA.XIR[8].XIC[9].icell.SM VGND.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2238 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t395 VPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2239 XThR.Tn[2].t2 XThR.XTBN.Y a_n1049_7493# VPWR.t484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2240 VGND.t1641 VPWR.t2037 XA.XIR[7].XIC_15.icell.PDM VGND.t1640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2241 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t1047 VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2242 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t1 VGND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2243 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t2520 VGND.t2519 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2244 XThR.Tn[13].t0 XThR.XTBN.Y VPWR.t483 VPWR.t482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2245 VGND.t157 Vbias.t208 XA.XIR[11].XIC[4].icell.SM VGND.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2246 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2248 VGND.t1910 VGND.t1908 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2249 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t1847 VPWR.t1846 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2250 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2251 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t1840 VGND.t1839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2252 XThR.Tn[10].t8 XThR.XTB3.Y.t13 VPWR.t652 VPWR.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2253 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t57 VGND.t660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2255 XThR.Tn[4].t0 XThR.XTBN.Y VGND.t860 VGND.t859 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2256 VPWR.t1796 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t1795 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2257 VGND.t2651 XThR.XTB6.Y XThR.Tn[5].t8 VGND.t2459 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2258 VGND.t2390 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2259 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t64 VGND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2260 VGND.t159 Vbias.t209 XA.XIR[12].XIC[12].icell.SM VGND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2261 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2262 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t173 VGND.t1527 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2263 VGND.t161 Vbias.t210 XA.XIR[15].XIC[13].icell.SM VGND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2264 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t5 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2265 VGND.t163 Vbias.t211 XA.XIR[14].XIC[14].icell.SM VGND.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2266 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t443 VGND.t442 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2267 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t1516 VGND.t1515 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2268 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2038 VGND.t1639 VGND.t1638 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2269 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t4 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2270 VGND.t2222 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t2221 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2271 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t397 VPWR.t396 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2272 VGND.t2224 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t2223 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2273 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2274 VPWR.t820 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t819 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2275 VGND.t1637 VPWR.t2039 XA.XIR[4].XIC_15.icell.PDM VGND.t1636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2276 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1144 VPWR.t1146 VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2277 VPWR.t856 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t855 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2278 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t30 VGND.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2279 VGND.t165 Vbias.t212 XA.XIR[5].XIC[3].icell.SM VGND.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2280 VGND.t167 Vbias.t213 XA.XIR[9].XIC[12].icell.SM VGND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2281 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t199 VGND.t2356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2282 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t175 VGND.t1530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2283 VGND.t1332 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t1331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2284 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2285 VGND.t169 Vbias.t214 XA.XIR[8].XIC[4].icell.SM VGND.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2286 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t1589 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t79 VGND.t944 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2288 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t1838 VGND.t1837 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 VGND.t1907 VGND.t1905 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2290 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2291 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t0 VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2292 VGND.t1635 VPWR.t2040 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t1634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2293 VGND.t1508 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1507 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2294 VPWR.t335 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2295 VPWR.t549 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2296 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t188 VGND.t2070 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2297 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2298 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t152 VGND.t1392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2299 VPWR.t1006 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2300 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t822 VPWR.t821 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2301 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t18 VGND.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2302 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2303 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t1049 VPWR.t1048 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2304 VGND.t2212 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t2211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2305 VPWR.t1798 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t1797 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2306 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2307 VPWR.t1143 VPWR.t1141 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1142 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2308 VGND.t2214 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t2213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2309 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t160 VPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2310 XThR.Tn[4].t9 XThR.XTB5.Y VGND.t2462 VGND.t2461 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2311 VPWR.t481 XThR.XTBN.Y XThR.Tn[14].t0 VPWR.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2312 VPWR.t591 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2313 XThC.Tn[13].t5 XThC.XTB6.Y VPWR.t620 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2314 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t151 VGND.t1381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2315 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t1517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2316 VGND.t1904 VGND.t1902 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2317 VGND.t1011 XThC.XTB6.Y XThC.Tn[5].t8 VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2318 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t1472 VGND.t1471 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2319 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t593 VPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2320 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t2476 VGND.t2475 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2321 VPWR.t479 XThR.XTBN.Y XThR.Tn[11].t4 VPWR.t478 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2322 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t1461 VGND.t1460 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2323 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t1836 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2324 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t77 VGND.t938 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2325 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t737 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2326 XThC.Tn[9].t4 XThC.XTB2.Y a_7875_9569# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2327 XA.XIR[4].XIC_15.icell.PDM VPWR.t2041 VGND.t1633 VGND.t1632 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2328 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t932 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 VGND.t2528 XThC.XTB6.A XThC.XTB6.Y VGND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2330 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t11 VGND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2331 VGND.t2377 XThC.XTB2.Y XThC.Tn[1].t9 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2332 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t1029 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2333 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1139 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1140 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2334 XThC.Tn[6].t0 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2335 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t204 VGND.t2368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2336 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t1413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2337 VGND.t1374 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t1373 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2338 VGND.t1115 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2339 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t1835 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2340 VPWR.t1613 XThR.XTB7.Y a_n1049_5317# VPWR.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2341 VPWR.t337 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2342 VGND.t1631 VPWR.t2042 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t1630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2343 VPWR.t619 XThC.XTB6.Y XThC.Tn[13].t4 VPWR.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2344 VPWR.t1008 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1007 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2345 a_n997_3979# XThR.XTBN.Y VGND.t858 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2346 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t788 VPWR.t787 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2347 VGND.t1901 VGND.t1899 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2348 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t1022 VPWR.t1021 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2349 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t339 VPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1136 VPWR.t1138 VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2351 VGND.t2017 XThR.XTB4.Y.t14 XThR.Tn[3].t11 VGND.t1075 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2352 a_7331_10587# data[0].t2 VPWR.t1869 VPWR.t1868 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2353 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t1 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2354 VPWR.t1478 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1477 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2355 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t2478 VGND.t2477 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2356 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1010 VPWR.t1009 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2357 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t162 VPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2358 VGND.t171 Vbias.t215 XA.XIR[2].XIC[7].icell.SM VGND.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2359 VPWR.t1 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2360 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t1473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2361 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2043 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2362 VPWR.t790 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t789 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2363 a_n1049_6699# XThR.XTBN.Y XThR.Tn[3].t3 VPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2364 XA.XIR[0].XIC[11].icell.PDM VGND.t1896 VGND.t1898 VGND.t1897 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2365 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t1777 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2366 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t113 VGND.t1089 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2367 XA.XIR[1].XIC_15.icell.PDM VPWR.t2044 VGND.t1628 VGND.t1627 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2368 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t75 VGND.t782 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2369 XThC.Tn[3].t4 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2370 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1134 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1135 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2371 XThC.XTB5.A data[0].t3 VGND.t2558 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2372 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t110 VGND.t1085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2373 VGND.t1561 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2374 VPWR.t1526 XThR.XTB4.Y.t15 XThR.Tn[11].t9 VPWR.t1525 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2375 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2376 VGND.t173 Vbias.t216 XA.XIR[10].XIC[5].icell.SM VGND.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2377 XA.XIR[0].XIC[2].icell.PDM VGND.t1893 VGND.t1895 VGND.t1894 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 VGND.t175 Vbias.t217 XA.XIR[13].XIC[6].icell.SM VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2379 VGND.t2065 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t2064 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2380 VGND.t856 XThR.XTBN.Y a_n997_715# VGND.t855 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2381 a_n997_2891# XThR.XTBN.Y VGND.t854 VGND.t853 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2382 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t238 VGND.t237 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t792 VPWR.t791 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2384 VPWR.t1806 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t1805 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2385 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t341 VPWR.t340 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2386 VPWR.t1476 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1475 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2387 VGND.t177 Vbias.t218 XA.XIR[4].XIC_15.icell.SM VGND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2388 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1131 VPWR.t1133 VPWR.t1132 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2389 VPWR.t3 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2390 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2391 VGND.t179 Vbias.t219 XA.XIR[11].XIC[13].icell.SM VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2392 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2393 XThR.Tn[11].t10 XThR.XTB4.Y.t16 a_n997_2667# VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2394 VPWR.t1130 VPWR.t1128 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1129 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2395 VGND.t1415 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t1414 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2396 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t115 VGND.t1092 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2397 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t1650 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2398 VPWR.t1766 XThC.XTB2.Y XThC.Tn[9].t8 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2399 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t1808 VPWR.t1807 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2400 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t2526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2401 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t0 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2402 VGND.t1626 VPWR.t2045 XA.XIR[0].XIC_15.icell.PDM VGND.t1625 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2403 VGND.t1510 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2404 VPWR.t374 XThC.XTBN.Y.t100 XThC.Tn[8].t0 VPWR.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2405 VGND.t181 Vbias.t220 XA.XIR[2].XIC[2].icell.SM VGND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2406 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t12 VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2407 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2408 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t1550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2409 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2410 VPWR.t236 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t235 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2411 XA.XIR[0].XIC[6].icell.PDM VGND.t1890 VGND.t1892 VGND.t1891 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2412 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t1462 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2413 a_n1049_6405# XThR.XTBN.Y XThR.Tn[4].t4 VPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2414 VGND.t183 Vbias.t221 XA.XIR[13].XIC[10].icell.SM VGND.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2415 XA.XIR[15].XIC[7].icell.Ien VPWR.t1125 VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2416 XThR.Tn[7].t0 XThR.XTBN.Y VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2417 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2046 VGND.t1624 VGND.t1623 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2418 VPWR.t794 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t793 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2419 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t25 VGND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2420 VPWR.t868 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t867 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2421 XThC.Tn[9].t0 XThC.XTBN.Y.t101 VPWR.t1689 VPWR.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2422 XThR.Tn[1].t1 XThR.XTBN.Y VGND.t852 VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2423 VPWR.t1111 VPWR.t1109 XA.XIR[13].XIC_15.icell.PUM VPWR.t1110 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2424 VGND.t2601 Vbias.t222 XA.XIR[10].XIC[0].icell.SM VGND.t2600 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2425 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t183 VGND.t2049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2426 VGND.t2603 Vbias.t223 XA.XIR[5].XIC[12].icell.SM VGND.t2602 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2427 VGND.t2605 Vbias.t224 XA.XIR[13].XIC[1].icell.SM VGND.t2604 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VGND.t2607 Vbias.t225 XA.XIR[8].XIC[13].icell.SM VGND.t2606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2429 VGND.t612 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2430 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t1567 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2431 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t1464 VGND.t1463 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2432 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t240 VGND.t239 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2433 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2047 VGND.t1622 VGND.t1621 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2434 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1074 VPWR.t1073 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2435 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t1810 VPWR.t1809 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2436 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t958 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2437 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t447 VGND.t446 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 VPWR.t1690 XThC.XTBN.Y.t102 XThC.Tn[11].t4 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2439 VPWR.t1474 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1473 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2440 VPWR.t1900 XThR.XTB6.Y a_n1049_5611# VPWR.t1612 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2441 VGND.t1620 VPWR.t2048 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1619 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2442 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t2 VGND.t46 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2443 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t1165 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2444 VPWR.t5 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2445 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t933 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2446 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t241 VGND.t2529 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2447 VGND.t2609 Vbias.t226 XA.XIR[7].XIC[11].icell.SM VGND.t2608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2448 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1123 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2449 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t1167 VGND.t1166 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2450 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t1169 VGND.t1168 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2451 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2453 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t187 VGND.t2061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2454 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t2521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2455 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t2483 VGND.t2482 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2456 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t1590 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2457 XA.XIR[15].XIC[11].icell.Ien VPWR.t1120 VPWR.t1122 VPWR.t1121 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2458 VGND.t1117 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 VGND.t1618 VPWR.t2049 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 XA.XIR[11].XIC_15.icell.PUM VPWR.t1118 XA.XIR[11].XIC_15.icell.Ien VPWR.t1119 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2461 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2462 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t1800 VPWR.t1799 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2463 VGND.t2579 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t2578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 VGND.t1616 VPWR.t2050 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XThC.Tn[2].t0 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2466 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2467 VPWR.t1818 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t1817 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2468 VPWR.t1059 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t1058 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2469 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t954 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 VGND.t728 XThR.XTB7.B XThR.XTB4.Y.t1 VGND.t727 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2471 VPWR.t1117 VPWR.t1115 XA.XIR[10].XIC_15.icell.PUM VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2472 XA.XIR[15].XIC[2].icell.Ien VPWR.t1112 VPWR.t1114 VPWR.t1113 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2473 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t595 VPWR.t594 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2474 VGND.t54 XThR.XTB1.Y.t16 XThR.Tn[0].t0 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2475 VGND.t2611 Vbias.t227 XA.XIR[1].XIC[7].icell.SM VGND.t2610 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2476 VPWR.t1668 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t1667 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2477 VPWR.t796 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t795 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2478 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t1024 VPWR.t1023 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2479 VGND.t2613 Vbias.t228 XA.XIR[4].XIC[8].icell.SM VGND.t2612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2480 VPWR.t1820 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t1819 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2481 XA.XIR[15].XIC[5].icell.PDM VPWR.t2051 XA.XIR[15].XIC[5].icell.Ien VGND.t1614 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2482 VGND.t2067 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t2066 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2483 VGND.t2615 Vbias.t229 XA.XIR[7].XIC[9].icell.SM VGND.t2614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2484 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t146 VGND.t1333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2485 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t253 VGND.t2670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2486 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1106 VPWR.t1108 VPWR.t1107 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2487 a_8739_9569# XThC.XTBN.Y.t104 VGND.t2265 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2488 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t149 VGND.t1336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2489 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t2485 VGND.t2484 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 XThC.Tn[6].t8 XThC.XTB7.Y VGND.t1401 VGND.t1400 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2491 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t1812 VPWR.t1811 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t960 VGND.t959 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2493 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t1181 VGND.t1180 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2494 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t2246 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2495 VGND.t2267 XThC.XTBN.Y.t105 XThC.Tn[7].t4 VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2496 XThC.Tn[12].t0 XThC.XTBN.Y.t106 VPWR.t1691 VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2497 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t1802 VPWR.t1801 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2498 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t1552 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2499 VGND.t1417 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t1416 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2500 VGND.t2617 Vbias.t230 XA.XIR[12].XIC[6].icell.SM VGND.t2616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2501 XThC.Tn[12].t8 XThC.XTB5.Y a_9827_9569# VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t2248 VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2503 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1896 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2504 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t955 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2505 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t6 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2506 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t1030 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2507 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1104 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1105 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2508 VGND.t2098 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t2097 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 VGND.t967 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t966 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2510 XThR.Tn[13].t9 XThR.XTB6.Y VPWR.t1899 VPWR.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2511 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t1804 VPWR.t1803 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2512 VGND.t2392 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2513 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2514 VGND.t2619 Vbias.t231 XA.XIR[6].XIC[5].icell.SM VGND.t2618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2515 VGND.t1376 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t1375 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2516 VPWR.t1670 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t1669 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2517 VGND.t1490 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t1489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2519 VGND.t2621 Vbias.t232 XA.XIR[9].XIC[6].icell.SM VGND.t2620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2520 VGND.t2268 XThC.XTBN.Y.t107 a_7875_9569# VGND.t41 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2521 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t2479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2522 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2052 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1613 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2523 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t1602 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2524 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t111 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2525 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1472 VPWR.t1471 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2526 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2527 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2528 VGND.t2623 Vbias.t233 XA.XIR[1].XIC[2].icell.SM VGND.t2622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2529 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t806 VPWR.t805 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2530 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t534 VPWR.t533 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2531 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t1183 VGND.t1182 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2532 VGND.t2625 Vbias.t234 XA.XIR[4].XIC[3].icell.SM VGND.t2624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2533 VPWR.t575 VGND.t2700 XA.XIR[0].XIC[12].icell.PUM VPWR.t574 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2534 XA.XIR[15].XIC[0].icell.PDM VPWR.t2053 XA.XIR[15].XIC[0].icell.Ien VGND.t1612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2535 a_8963_9569# XThC.XTBN.Y.t108 VGND.t2269 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2536 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t961 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2537 VGND.t614 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2538 VGND.t2627 Vbias.t235 XA.XIR[7].XIC[4].icell.SM VGND.t2626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2539 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2540 VGND.t1889 VGND.t1887 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2541 VGND.t2629 Vbias.t236 XA.XIR[12].XIC[10].icell.SM VGND.t2628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2542 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t234 VGND.t2513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2543 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t2250 VGND.t2249 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2544 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t1474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2545 VPWR.t1103 VPWR.t1101 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1102 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2546 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t237 VGND.t2523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2547 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t1476 VGND.t1475 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t1201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2550 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t1202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t417 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t416 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 VGND.t1559 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XThC.Tn[11].t3 XThC.XTBN.Y.t109 VPWR.t1692 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2554 VPWR.t597 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t596 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2555 VGND.t2631 Vbias.t237 XA.XIR[3].XIC[5].icell.SM VGND.t2630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2556 XThR.Tn[6].t1 XThR.XTBN.Y a_n1049_5317# VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2557 VGND.t2633 Vbias.t238 XA.XIR[12].XIC[1].icell.SM VGND.t2632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2558 VGND.t2635 Vbias.t239 XA.XIR[9].XIC[10].icell.SM VGND.t2634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2559 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2560 VPWR.t101 XThC.XTB4.Y.t16 XThC.Tn[11].t7 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2561 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2562 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t1568 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t1525 VGND.t1524 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2564 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2565 VGND.t2637 Vbias.t240 XA.XIR[10].XIC[14].icell.SM VGND.t2636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2566 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t930 VGND.t929 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2567 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2054 VGND.t1611 VGND.t1610 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2568 VGND.t2226 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t2225 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2569 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2570 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1470 VPWR.t1469 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2571 XA.XIR[12].XIC_15.icell.PDM VPWR.t2055 VGND.t1609 VGND.t1608 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2572 VGND.t2639 Vbias.t241 XA.XIR[6].XIC[0].icell.SM VGND.t2638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2573 VPWR.t577 VGND.t2701 XA.XIR[0].XIC[10].icell.PUM VPWR.t576 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2574 VGND.t2641 Vbias.t242 XA.XIR[9].XIC[1].icell.SM VGND.t2640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2575 VPWR.t1827 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2576 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2577 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t132 VGND.t1217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2578 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2579 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t970 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2580 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t962 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2581 VGND.t850 XThR.XTBN.Y a_n997_1803# VGND.t849 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2582 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t715 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2583 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t824 VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2584 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2585 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t205 VGND.t2369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2586 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t115 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2587 XA.XIR[10].XIC_15.icell.PUM VPWR.t1099 XA.XIR[10].XIC_15.icell.Ien VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2588 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t106 VGND.t1061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2589 a_3773_9615# XThC.XTB2.Y VPWR.t1765 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2590 VPWR.t1098 VPWR.t1096 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1097 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2591 VGND.t1512 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2592 VGND.t2581 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2593 VPWR.t419 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t418 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2594 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t738 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2595 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t136 VGND.t1229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2596 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t138 VGND.t1246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2597 VPWR.t1528 XThR.XTB4.Y.t17 XThR.Tn[11].t11 VPWR.t1527 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2598 a_n997_715# XThR.XTBN.Y VGND.t848 VGND.t847 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2599 VPWR.t51 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2600 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2601 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t808 VPWR.t807 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2602 XThR.Tn[14].t9 XThR.XTB7.Y VPWR.t1611 VPWR.t1610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2603 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t676 VGND.t675 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2604 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t536 VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2605 VGND.t2270 XThC.XTBN.Y.t110 XThC.Tn[3].t1 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2606 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t1822 VPWR.t1821 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2607 VGND.t203 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2608 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2056 VGND.t1607 VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2609 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t1203 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2610 VPWR.t421 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t420 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2611 XThC.Tn[1].t8 XThC.XTB2.Y VGND.t2376 VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2612 VPWR.t1468 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1467 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2613 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t1184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2614 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t206 VPWR.t205 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2615 VPWR.t838 XThC.XTBN.A XThC.XTBN.Y.t0 VPWR.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2616 VPWR.t644 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t643 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2617 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t931 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2618 VPWR.t11 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2619 VGND.t2643 Vbias.t243 XA.XIR[3].XIC[0].icell.SM VGND.t2642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2620 VPWR.t1095 VPWR.t1093 XA.XIR[6].XIC_15.icell.PUM VPWR.t1094 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2621 VGND.t1886 VGND.t1884 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2622 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t116 VGND.t1093 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2623 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t716 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2624 XThR.Tn[2].t0 XThR.XTB3.Y.t16 VGND.t289 VGND.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2625 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t191 VGND.t2175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2626 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t933 VGND.t932 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2627 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2628 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t161 VGND.t1439 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2629 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2630 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t718 VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2631 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t1 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2632 a_3299_10575# XThC.XTB7.B VGND.t123 VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2633 VGND.t1605 VPWR.t2057 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t1604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2634 VGND.t846 XThR.XTBN.Y XThR.Tn[6].t4 VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2635 VPWR.t579 VGND.t2702 XA.XIR[0].XIC[5].icell.PUM VPWR.t578 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2636 VGND.t2645 Vbias.t244 XA.XIR[0].XIC[11].icell.SM VGND.t2644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2637 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t934 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2638 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t80 VGND.t948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2639 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t1604 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2640 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t83 VGND.t951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2641 VPWR.t208 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t207 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2642 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t971 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2643 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t169 VGND.t1459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2644 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1090 VPWR.t1092 VPWR.t1091 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2645 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t200 VGND.t2357 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2646 VGND.t2103 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t2102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2647 VGND.t1119 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2648 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t1824 VPWR.t1823 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2649 VGND.t199 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2650 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t1204 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2651 VGND.t2583 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t2582 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VPWR.t1693 XThC.XTBN.Y.t111 XThC.Tn[10].t7 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2653 VGND.t1492 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2654 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t211 VGND.t2380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2655 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2058 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t1603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2656 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t956 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2657 VGND.t1100 XThC.XTBN.Y.t112 a_8963_9569# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2658 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t810 VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2659 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t4 VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 VPWR.t988 XThC.XTB5.A a_5155_10571# VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2661 VPWR.t961 XThC.XTB7.Y XThC.Tn[14].t8 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2662 XThR.Tn[1].t0 XThR.XTBN.Y VGND.t844 VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t1672 VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t538 VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2665 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t1826 VPWR.t1825 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2666 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t1814 VPWR.t1813 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2667 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t160 VGND.t1438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2668 VPWR.t1832 XThC.XTB7.A XThC.XTB3.Y.t2 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2669 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t210 VPWR.t209 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2670 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t1185 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2671 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2672 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t934 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2673 XThR.Tn[8].t3 XThR.XTBN.Y VPWR.t474 VPWR.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2674 VGND.t1883 VGND.t1881 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2675 VPWR.t698 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t697 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2676 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2059 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t1602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2677 XThR.Tn[5].t0 XThR.XTBN.Y a_n1049_5611# VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2678 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t9 VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2679 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t1031 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2680 VGND.t2647 Vbias.t245 XA.XIR[0].XIC[9].icell.SM VGND.t2646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2681 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2682 VPWR.t1085 VPWR.t1083 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2683 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t44 VGND.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2684 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t184 VGND.t2051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2685 a_n1049_7787# XThR.XTBN.Y XThR.Tn[1].t4 VPWR.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2686 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t1 VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2687 VPWR.t427 XThR.XTB7.B XThR.XTB3.Y.t0 VPWR.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2688 VGND.t497 Vbias.t246 XA.XIR[5].XIC[6].icell.SM VGND.t496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2689 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2060 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t1601 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2690 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1897 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2691 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t1828 VPWR.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2692 VPWR.t1829 XThC.XTB3.Y.t16 XThC.Tn[10].t9 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2693 VPWR.t730 XThC.XTBN.Y.t114 XThC.Tn[14].t1 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2694 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t700 VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2695 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t739 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2696 XA.XIR[15].XIC_15.icell.PDM VPWR.t2061 VGND.t1600 VGND.t1599 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2697 VGND.t2105 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t2104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2698 VGND.t842 XThR.XTBN.Y XThR.Tn[0].t6 VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2699 VGND.t499 Vbias.t247 XA.XIR[4].XIC[12].icell.SM VGND.t498 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2700 VGND.t2486 XThC.XTB3.Y.t17 XThC.Tn[2].t11 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2701 VGND.t501 Vbias.t248 XA.XIR[7].XIC[13].icell.SM VGND.t500 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2702 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2703 XThR.Tn[10].t4 XThR.XTBN.Y VPWR.t470 VPWR.t469 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2704 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t6 VGND.t5 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2705 VGND.t503 Vbias.t249 XA.XIR[6].XIC[14].icell.SM VGND.t502 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2706 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2062 VGND.t1598 VGND.t1597 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2707 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t117 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2708 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t1603 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2709 VPWR.t618 XThC.XTB6.Y a_5949_9615# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2710 XThR.Tn[1].t8 XThR.XTB2.Y VGND.t1465 VGND.t1072 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2711 VGND.t840 XThR.XTBN.Y a_n997_3755# VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2712 VPWR.t547 data[3].t1 XThC.XTBN.A VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2713 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t440 VPWR.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2714 XThC.Tn[3].t0 XThC.XTBN.Y.t115 VGND.t1101 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2715 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1466 VPWR.t1465 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2716 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t120 VGND.t1109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2717 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t1032 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2718 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t2480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2719 VGND.t505 Vbias.t250 XA.XIR[0].XIC[4].icell.SM VGND.t504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2720 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t209 VGND.t2374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2721 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t600 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2722 VGND.t507 Vbias.t251 XA.XIR[5].XIC[10].icell.SM VGND.t506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2723 VPWR.t385 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t384 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2724 VGND.t509 Vbias.t252 XA.XIR[13].XIC[7].icell.SM VGND.t508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2725 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t646 VPWR.t645 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2726 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2727 VPWR.t702 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t701 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2728 VPWR.t285 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t284 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2729 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t1025 VGND.t1024 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2730 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t1605 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2731 VGND.t1880 VGND.t1878 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2732 VPWR.t1076 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1075 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2733 XThR.Tn[13].t8 XThR.XTB6.Y VPWR.t1898 VPWR.t1620 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2734 VGND.t511 Vbias.t253 XA.XIR[5].XIC[1].icell.SM VGND.t510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2735 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t247 VGND.t2589 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2736 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1887 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2737 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t1559 VPWR.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2738 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t1570 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 VGND.t513 Vbias.t254 XA.XIR[3].XIC[14].icell.SM VGND.t512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2740 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t177 VGND.t1874 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2741 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t1571 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2742 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t720 VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2743 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t1833 VGND.t1832 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2744 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t1027 VGND.t1026 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2745 VPWR.t442 XThC.XTB1.Y.t18 XThC.Tn[8].t8 VPWR.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2746 VGND.t2069 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t2068 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2747 VGND.t2460 XThR.XTB5.Y XThR.Tn[4].t8 VGND.t2459 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2748 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t59 VGND.t669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2749 XThC.Tn[10].t6 XThC.XTBN.Y.t116 VPWR.t731 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2750 VGND.t1103 XThC.XTBN.Y.t117 XThC.Tn[6].t4 VGND.t1102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2751 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t2481 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2752 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t972 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2753 VPWR.t1061 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t1060 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2754 VPWR.t387 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2755 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t973 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2756 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2757 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t2669 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2758 VGND.t515 Vbias.t255 XA.XIR[15].XIC_15.icell.SM VGND.t514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2759 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2760 XA.XIR[3].XIC_15.icell.PUM VPWR.t1088 XA.XIR[3].XIC_15.icell.Ien VPWR.t1089 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t1554 VGND.t1553 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2762 VGND.t201 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2763 VGND.t1596 VPWR.t2063 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t1595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 VGND.t2585 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t2584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 VGND.t1419 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t1418 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 VGND.t2587 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t36 VGND.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2768 VPWR.t287 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t286 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2769 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t212 VPWR.t211 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2770 VPWR.t102 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2771 VPWR.t295 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2772 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t1063 VPWR.t1062 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2773 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t98 VGND.t1006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2774 XA.XIR[15].XIC[11].icell.PDM VPWR.t2064 XA.XIR[15].XIC[11].icell.Ien VGND.t1594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2775 VGND.t1593 VPWR.t2065 XA.XIR[11].XIC_15.icell.PDM VGND.t1592 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2776 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2777 VGND.t517 Vbias.t256 XA.XIR[13].XIC[2].icell.SM VGND.t516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2778 XThR.Tn[6].t0 XThR.XTBN.Y a_n1049_5317# VPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2779 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2780 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1086 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1087 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2781 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t87 VGND.t963 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2782 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t4 VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2783 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1464 VPWR.t1463 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2784 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t648 VPWR.t647 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2785 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2786 VGND.t1105 XThC.XTBN.Y.t118 a_10915_9569# VGND.t1104 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2787 VPWR.t704 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t703 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2788 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t812 VPWR.t811 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2789 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t1029 VGND.t1028 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2790 VGND.t1378 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t1377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2791 VPWR.t289 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t288 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2792 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t540 VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2793 VPWR.t297 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2794 VPWR.t581 VGND.t2703 XA.XIR[0].XIC[14].icell.PUM VPWR.t580 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2795 XA.XIR[15].XIC[2].icell.PDM VPWR.t2066 XA.XIR[15].XIC[2].icell.Ien VGND.t1591 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2796 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2797 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t219 VGND.t2401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2798 XThC.Tn[1].t0 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2799 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t249 VGND.t2649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2800 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t201 VGND.t2358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2801 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2802 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t134 VGND.t1227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2803 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t1830 VGND.t1829 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2804 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t573 VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2805 XThC.Tn[14].t0 XThC.XTBN.Y.t120 VPWR.t732 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2806 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t34 VGND.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2807 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2067 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t1590 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2808 VGND.t616 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2809 VGND.t838 XThR.XTBN.Y a_n997_715# VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2810 VPWR.t1082 VPWR.t1080 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1081 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2811 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t1065 VPWR.t1064 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2812 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t154 VGND.t1395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2813 VPWR.t599 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2814 VPWR.t1609 XThR.XTB7.Y XThR.Tn[14].t8 VPWR.t1608 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2815 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2816 VGND.t519 Vbias.t257 XA.XIR[14].XIC[11].icell.SM VGND.t518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2817 XThR.XTB6.A data[5].t5 VGND.t2553 VGND.t2552 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2818 XThR.Tn[0].t2 XThR.XTBN.Y a_n1049_8581# VPWR.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 VGND.t2107 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t2106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2820 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t636 VGND.t635 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2821 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t638 VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2822 VGND.t2109 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t2108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2823 VGND.t1557 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t1556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2824 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t214 VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2825 a_5949_9615# XThC.XTB6.Y VPWR.t617 VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2826 VGND.t1106 XThC.XTBN.Y.t121 a_10051_9569# VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2827 VGND.t1380 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t1379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2828 VGND.t521 Vbias.t258 XA.XIR[2].XIC[5].icell.SM VGND.t520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2829 VGND.t1494 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2830 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2068 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t1589 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2831 XA.XIR[15].XIC[6].icell.PDM VPWR.t2069 XA.XIR[15].XIC[6].icell.Ien VGND.t1588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2832 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t639 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2833 XA.XIR[0].XIC[9].icell.PDM VGND.t1875 VGND.t1877 VGND.t1876 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2834 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t2364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2835 VPWR.t733 XThC.XTBN.Y.t122 XThC.Tn[11].t2 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2836 VGND.t964 XThC.XTBN.Y.t123 a_7651_9569# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2837 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1462 VPWR.t1461 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2838 Vbias.t0 bias[1].t0 VPWR.t448 VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=2
X2839 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t706 VPWR.t705 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2840 XThR.Tn[2].t1 XThR.XTBN.Y VGND.t834 VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2841 VPWR.t1607 XThR.XTB7.Y a_n1049_5317# VPWR.t1606 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2842 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t10 VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2843 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2844 VGND.t969 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t968 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2845 VGND.t2100 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t2099 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2846 VPWR.t466 XThR.XTBN.Y XThR.Tn[12].t0 VPWR.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2847 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t1828 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2848 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t7 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2849 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t1186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2850 VGND.t523 Vbias.t259 XA.XIR[12].XIC[7].icell.SM VGND.t522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2851 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t198 VGND.t2355 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2852 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t7 VGND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2853 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t935 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2854 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1311 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2855 VGND.t525 Vbias.t260 XA.XIR[15].XIC[8].icell.SM VGND.t524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2856 VPWR.t1079 VPWR.t1077 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2857 VGND.t1514 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1513 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2858 VGND.t527 Vbias.t261 XA.XIR[14].XIC[9].icell.SM VGND.t526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2859 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t937 VGND.t936 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2860 VPWR.t1816 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t1815 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R1 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R2 XThR.Tn[2] XThR.Tn[2].n82 161.363
R3 XThR.Tn[2] XThR.Tn[2].n77 161.363
R4 XThR.Tn[2] XThR.Tn[2].n72 161.363
R5 XThR.Tn[2] XThR.Tn[2].n67 161.363
R6 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7 XThR.Tn[2] XThR.Tn[2].n57 161.363
R8 XThR.Tn[2] XThR.Tn[2].n52 161.363
R9 XThR.Tn[2] XThR.Tn[2].n47 161.363
R10 XThR.Tn[2] XThR.Tn[2].n42 161.363
R11 XThR.Tn[2] XThR.Tn[2].n37 161.363
R12 XThR.Tn[2] XThR.Tn[2].n32 161.363
R13 XThR.Tn[2] XThR.Tn[2].n27 161.363
R14 XThR.Tn[2] XThR.Tn[2].n22 161.363
R15 XThR.Tn[2] XThR.Tn[2].n17 161.363
R16 XThR.Tn[2] XThR.Tn[2].n12 161.363
R17 XThR.Tn[2] XThR.Tn[2].n10 161.363
R18 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R19 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R20 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R21 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R22 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R23 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R24 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R25 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R26 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R27 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R28 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R29 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R30 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R31 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R32 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R33 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R34 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R35 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R36 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R37 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R38 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R39 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R40 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R41 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R42 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R43 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R44 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R45 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R46 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R47 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R48 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R49 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R50 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R51 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R52 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R53 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R54 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R55 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R56 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R57 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R58 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R59 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R60 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R61 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R62 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R63 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R64 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R65 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R66 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R67 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R68 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R69 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R70 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R71 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R72 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R73 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R74 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R75 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R76 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R77 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R78 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R79 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R80 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R81 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R82 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R83 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R84 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R85 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R86 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R87 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R88 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R89 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R90 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R91 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R92 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R93 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R94 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R95 XThR.Tn[2].n7 XThR.Tn[2].n5 135.249
R96 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R97 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R98 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R99 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R100 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R101 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R102 XThR.Tn[2].n1 XThR.Tn[2].t4 26.5955
R103 XThR.Tn[2].n1 XThR.Tn[2].t3 26.5955
R104 XThR.Tn[2].n0 XThR.Tn[2].t5 26.5955
R105 XThR.Tn[2].n0 XThR.Tn[2].t2 26.5955
R106 XThR.Tn[2].n3 XThR.Tn[2].t7 24.9236
R107 XThR.Tn[2].n3 XThR.Tn[2].t8 24.9236
R108 XThR.Tn[2].n4 XThR.Tn[2].t6 24.9236
R109 XThR.Tn[2].n4 XThR.Tn[2].t1 24.9236
R110 XThR.Tn[2].n5 XThR.Tn[2].t9 24.9236
R111 XThR.Tn[2].n5 XThR.Tn[2].t10 24.9236
R112 XThR.Tn[2].n6 XThR.Tn[2].t11 24.9236
R113 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R114 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R115 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R116 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R117 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R118 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R119 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R120 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R121 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R122 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R123 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R124 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R125 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R126 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R127 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R128 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R129 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R130 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R131 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R132 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R133 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R134 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R135 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R136 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R137 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R138 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R139 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R140 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R141 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R142 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R143 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R144 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R145 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R146 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R147 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R148 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R149 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R150 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R151 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R152 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R153 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R154 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R155 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R156 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R157 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R158 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R159 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R160 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R161 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R162 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R163 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R164 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R165 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R166 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R167 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R168 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R169 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R170 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R171 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R172 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R173 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R174 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R175 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R176 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R177 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R178 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R179 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R180 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R181 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R182 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R183 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R184 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R185 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R186 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R187 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R188 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R189 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R190 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R191 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R192 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R193 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R194 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R195 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R196 XThR.Tn[2] XThR.Tn[2].n87 0.038
R197 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R198 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R199 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R200 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R201 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R202 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R203 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R204 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R205 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R206 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R207 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R208 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R209 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R210 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R211 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R212 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R213 VPWR.n2837 VPWR.n2823 2618.82
R214 VPWR.n2835 VPWR.n2829 2618.82
R215 VPWR.n2853 VPWR.n2823 1916.47
R216 VPWR.n2828 VPWR.n2827 1916.47
R217 VPWR.n2827 VPWR.n2821 1916.47
R218 VPWR.n2829 VPWR.n2822 1916.47
R219 VPWR.n2852 VPWR.n2824 1912.94
R220 VPWR.n2849 VPWR.n2843 1560
R221 VPWR.n2850 VPWR.n2824 1408.24
R222 VPWR.n2853 VPWR.n2852 1210.59
R223 VPWR.n2851 VPWR.n2821 1210.59
R224 VPWR.n2380 VPWR.t1225 1005.7
R225 VPWR.t1443 VPWR.n485 1005.7
R226 VPWR.t1292 VPWR.n2210 1005.7
R227 VPWR.n639 VPWR.t1400 1005.7
R228 VPWR.n2184 VPWR.t1126 1005.7
R229 VPWR.t1233 VPWR.n677 1005.7
R230 VPWR.t1193 VPWR.n2014 1005.7
R231 VPWR.n831 VPWR.t1298 1005.7
R232 VPWR.n1988 VPWR.t1121 1005.7
R233 VPWR.t1305 VPWR.n869 1005.7
R234 VPWR.n447 VPWR.t1113 1005.7
R235 VPWR.t1413 VPWR.n1818 1005.7
R236 VPWR.t1395 VPWR.n2406 1005.7
R237 VPWR.n1023 VPWR.t1265 1005.7
R238 VPWR.t1435 VPWR.n293 1005.7
R239 VPWR.n1792 VPWR.t1376 1005.7
R240 VPWR.n2591 VPWR.t1327 1005.7
R241 VPWR.n1062 VPWR.t1211 1005.7
R242 VPWR.t1842 VPWR.n2309 983.14
R243 VPWR.n2310 VPWR.t913 983.14
R244 VPWR.t1519 VPWR.n2319 983.14
R245 VPWR.n2320 VPWR.t153 983.14
R246 VPWR.t849 VPWR.n2329 983.14
R247 VPWR.n2330 VPWR.t944 983.14
R248 VPWR.t300 VPWR.n2339 983.14
R249 VPWR.n2340 VPWR.t457 983.14
R250 VPWR.t407 VPWR.n2349 983.14
R251 VPWR.n2350 VPWR.t64 983.14
R252 VPWR.t643 VPWR.n2359 983.14
R253 VPWR.n2360 VPWR.t1007 983.14
R254 VPWR.t98 VPWR.n2369 983.14
R255 VPWR.n2370 VPWR.t1549 983.14
R256 VPWR.t1058 VPWR.n2379 983.14
R257 VPWR.n542 VPWR.t921 983.14
R258 VPWR.n541 VPWR.t1667 983.14
R259 VPWR.n537 VPWR.t1497 983.14
R260 VPWR.n533 VPWR.t131 983.14
R261 VPWR.n529 VPWR.t403 983.14
R262 VPWR.n525 VPWR.t783 983.14
R263 VPWR.n521 VPWR.t195 983.14
R264 VPWR.n517 VPWR.t145 983.14
R265 VPWR.n513 VPWR.t449 983.14
R266 VPWR.n509 VPWR.t328 983.14
R267 VPWR.n505 VPWR.t997 983.14
R268 VPWR.n501 VPWR.t215 983.14
R269 VPWR.n497 VPWR.t1787 983.14
R270 VPWR.n493 VPWR.t352 983.14
R271 VPWR.n489 VPWR.t24 983.14
R272 VPWR.n2281 VPWR.t1557 983.14
R273 VPWR.n2280 VPWR.t1578 983.14
R274 VPWR.n2271 VPWR.t1473 983.14
R275 VPWR.n2270 VPWR.t320 983.14
R276 VPWR.n2261 VPWR.t1874 983.14
R277 VPWR.n2260 VPWR.t1753 983.14
R278 VPWR.n2251 VPWR.t4 983.14
R279 VPWR.n2250 VPWR.t1703 983.14
R280 VPWR.n2241 VPWR.t139 983.14
R281 VPWR.n2240 VPWR.t762 983.14
R282 VPWR.n2231 VPWR.t392 983.14
R283 VPWR.n2230 VPWR.t669 983.14
R284 VPWR.n2221 VPWR.t877 983.14
R285 VPWR.n2220 VPWR.t598 983.14
R286 VPWR.n2211 VPWR.t225 983.14
R287 VPWR.t1741 VPWR.n582 983.14
R288 VPWR.t701 VPWR.n586 983.14
R289 VPWR.t1487 VPWR.n590 983.14
R290 VPWR.t1725 VPWR.n594 983.14
R291 VPWR.t748 VPWR.n598 983.14
R292 VPWR.t793 VPWR.n602 983.14
R293 VPWR.t271 VPWR.n606 983.14
R294 VPWR.t1854 VPWR.n610 983.14
R295 VPWR.t659 VPWR.n614 983.14
R296 VPWR.t334 VPWR.n618 983.14
R297 VPWR.t1626 VPWR.n622 983.14
R298 VPWR.t889 VPWR.n626 983.14
R299 VPWR.t1795 VPWR.n630 983.14
R300 VPWR.t637 VPWR.n634 983.14
R301 VPWR.t30 VPWR.n638 983.14
R302 VPWR.t284 VPWR.n2113 983.14
R303 VPWR.n2114 VPWR.t722 983.14
R304 VPWR.t1509 VPWR.n2123 983.14
R305 VPWR.n2124 VPWR.t1815 983.14
R306 VPWR.t1075 VPWR.n2133 983.14
R307 VPWR.n2134 VPWR.t1677 983.14
R308 VPWR.t310 VPWR.n2143 983.14
R309 VPWR.n2144 VPWR.t416 983.14
R310 VPWR.t867 VPWR.n2153 983.14
R311 VPWR.n2154 VPWR.t1531 983.14
R312 VPWR.t825 VPWR.n2163 983.14
R313 VPWR.n2164 VPWR.t1596 983.14
R314 VPWR.t255 VPWR.n2173 983.14
R315 VPWR.n2174 VPWR.t356 983.14
R316 VPWR.t1715 VPWR.n2183 983.14
R317 VPWR.n734 VPWR.t633 983.14
R318 VPWR.n733 VPWR.t911 983.14
R319 VPWR.n729 VPWR.t1521 983.14
R320 VPWR.n725 VPWR.t151 983.14
R321 VPWR.n721 VPWR.t746 983.14
R322 VPWR.n717 VPWR.t942 983.14
R323 VPWR.n713 VPWR.t298 983.14
R324 VPWR.n709 VPWR.t203 983.14
R325 VPWR.n705 VPWR.t405 983.14
R326 VPWR.n701 VPWR.t62 983.14
R327 VPWR.n697 VPWR.t596 983.14
R328 VPWR.n693 VPWR.t1005 983.14
R329 VPWR.n689 VPWR.t96 983.14
R330 VPWR.n685 VPWR.t1056 983.14
R331 VPWR.n681 VPWR.t235 983.14
R332 VPWR.n2085 VPWR.t819 983.14
R333 VPWR.n2084 VPWR.t1838 983.14
R334 VPWR.n2075 VPWR.t1515 983.14
R335 VPWR.n2074 VPWR.t1805 983.14
R336 VPWR.n2065 VPWR.t855 983.14
R337 VPWR.n2064 VPWR.t950 983.14
R338 VPWR.n2055 VPWR.t306 983.14
R339 VPWR.n2054 VPWR.t155 983.14
R340 VPWR.n2045 VPWR.t863 983.14
R341 VPWR.n2044 VPWR.t70 983.14
R342 VPWR.n2035 VPWR.t1914 983.14
R343 VPWR.n2034 VPWR.t207 983.14
R344 VPWR.n2025 VPWR.t245 983.14
R345 VPWR.n2024 VPWR.t584 983.14
R346 VPWR.n2015 VPWR.t1060 983.14
R347 VPWR.t1555 VPWR.n774 983.14
R348 VPWR.t679 VPWR.n778 983.14
R349 VPWR.t1475 VPWR.n782 983.14
R350 VPWR.t316 VPWR.n786 983.14
R351 VPWR.t1872 VPWR.n790 983.14
R352 VPWR.t959 VPWR.n794 983.14
R353 VPWR.t2 VPWR.n798 983.14
R354 VPWR.t1699 VPWR.n802 983.14
R355 VPWR.t137 VPWR.n806 983.14
R356 VPWR.t760 VPWR.n810 983.14
R357 VPWR.t390 VPWR.n814 983.14
R358 VPWR.t777 VPWR.n818 983.14
R359 VPWR.t873 VPWR.n822 983.14
R360 VPWR.t386 VPWR.n826 983.14
R361 VPWR.t221 VPWR.n830 983.14
R362 VPWR.t286 VPWR.n1917 983.14
R363 VPWR.n1918 VPWR.t724 983.14
R364 VPWR.t1507 VPWR.n1927 983.14
R365 VPWR.n1928 VPWR.t1572 983.14
R366 VPWR.t294 VPWR.n1937 983.14
R367 VPWR.n1938 VPWR.t1679 983.14
R368 VPWR.t185 VPWR.n1947 983.14
R369 VPWR.n1948 VPWR.t418 983.14
R370 VPWR.t1817 VPWR.n1957 983.14
R371 VPWR.n1958 VPWR.t1533 983.14
R372 VPWR.t827 VPWR.n1967 983.14
R373 VPWR.n1968 VPWR.t1598 983.14
R374 VPWR.t257 VPWR.n1977 983.14
R375 VPWR.n1978 VPWR.t358 983.14
R376 VPWR.t1717 VPWR.n1987 983.14
R377 VPWR.n926 VPWR.t1553 983.14
R378 VPWR.n925 VPWR.t677 983.14
R379 VPWR.n921 VPWR.t1477 983.14
R380 VPWR.n917 VPWR.t314 983.14
R381 VPWR.n913 VPWR.t1870 983.14
R382 VPWR.n909 VPWR.t957 983.14
R383 VPWR.n905 VPWR.t0 983.14
R384 VPWR.n901 VPWR.t1858 983.14
R385 VPWR.n897 VPWR.t135 983.14
R386 VPWR.n893 VPWR.t758 983.14
R387 VPWR.n889 VPWR.t388 983.14
R388 VPWR.n885 VPWR.t775 983.14
R389 VPWR.n881 VPWR.t869 983.14
R390 VPWR.n877 VPWR.t384 983.14
R391 VPWR.n873 VPWR.t219 983.14
R392 VPWR.t288 VPWR.n390 983.14
R393 VPWR.t726 VPWR.n394 983.14
R394 VPWR.t1505 VPWR.n398 983.14
R395 VPWR.t1576 VPWR.n402 983.14
R396 VPWR.t296 VPWR.n406 983.14
R397 VPWR.t797 VPWR.n410 983.14
R398 VPWR.t187 VPWR.n414 983.14
R399 VPWR.t420 VPWR.n418 983.14
R400 VPWR.t1819 VPWR.n422 983.14
R401 VPWR.t1535 VPWR.n426 983.14
R402 VPWR.t829 VPWR.n430 983.14
R403 VPWR.t1600 VPWR.n434 983.14
R404 VPWR.t259 VPWR.n438 983.14
R405 VPWR.t360 VPWR.n442 983.14
R406 VPWR.t18 VPWR.n446 983.14
R407 VPWR.n1889 VPWR.t435 983.14
R408 VPWR.n1888 VPWR.t697 983.14
R409 VPWR.n1879 VPWR.t1489 983.14
R410 VPWR.n1878 VPWR.t1723 983.14
R411 VPWR.n1869 VPWR.t978 983.14
R412 VPWR.n1868 VPWR.t789 983.14
R413 VPWR.n1859 VPWR.t267 983.14
R414 VPWR.n1858 VPWR.t1852 983.14
R415 VPWR.n1849 VPWR.t455 983.14
R416 VPWR.n1848 VPWR.t332 983.14
R417 VPWR.n1839 VPWR.t1622 983.14
R418 VPWR.n1838 VPWR.t887 983.14
R419 VPWR.n1829 VPWR.t1793 983.14
R420 VPWR.n1828 VPWR.t635 983.14
R421 VPWR.n1819 VPWR.t28 983.14
R422 VPWR.n2477 VPWR.t1743 983.14
R423 VPWR.n2476 VPWR.t703 983.14
R424 VPWR.n2467 VPWR.t1485 983.14
R425 VPWR.n2466 VPWR.t1729 983.14
R426 VPWR.n2457 VPWR.t750 983.14
R427 VPWR.n2456 VPWR.t795 983.14
R428 VPWR.n2447 VPWR.t273 983.14
R429 VPWR.n2446 VPWR.t1856 983.14
R430 VPWR.n2437 VPWR.t661 983.14
R431 VPWR.n2436 VPWR.t336 983.14
R432 VPWR.n2427 VPWR.t1628 983.14
R433 VPWR.n2426 VPWR.t891 983.14
R434 VPWR.n2417 VPWR.t1797 983.14
R435 VPWR.n2416 VPWR.t639 983.14
R436 VPWR.n2407 VPWR.t167 983.14
R437 VPWR.t625 VPWR.n966 983.14
R438 VPWR.t1584 VPWR.n970 983.14
R439 VPWR.t1467 VPWR.n974 983.14
R440 VPWR.t326 VPWR.n978 983.14
R441 VPWR.t740 VPWR.n982 983.14
R442 VPWR.t1759 VPWR.n986 983.14
R443 VPWR.t10 VPWR.n990 983.14
R444 VPWR.t1707 VPWR.n994 983.14
R445 VPWR.t179 VPWR.n998 983.14
R446 VPWR.t764 VPWR.n1002 983.14
R447 VPWR.t590 VPWR.n1006 983.14
R448 VPWR.t671 VPWR.n1010 983.14
R449 VPWR.t88 VPWR.n1014 983.14
R450 VPWR.t641 VPWR.n1018 983.14
R451 VPWR.t231 VPWR.n1022 983.14
R452 VPWR.n350 VPWR.t923 983.14
R453 VPWR.n349 VPWR.t1669 983.14
R454 VPWR.n345 VPWR.t1493 983.14
R455 VPWR.n341 VPWR.t1721 983.14
R456 VPWR.n337 VPWR.t974 983.14
R457 VPWR.n333 VPWR.t785 983.14
R458 VPWR.n329 VPWR.t197 983.14
R459 VPWR.n325 VPWR.t1850 983.14
R460 VPWR.n321 VPWR.t451 983.14
R461 VPWR.n317 VPWR.t330 983.14
R462 VPWR.n313 VPWR.t999 983.14
R463 VPWR.n309 VPWR.t217 983.14
R464 VPWR.n305 VPWR.t1791 983.14
R465 VPWR.n301 VPWR.t354 983.14
R466 VPWR.n297 VPWR.t26 983.14
R467 VPWR.t1346 VPWR.n1468 983.14
R468 VPWR.t1448 VPWR.n1475 983.14
R469 VPWR.t1219 VPWR.n1481 983.14
R470 VPWR.t1321 VPWR.n1492 983.14
R471 VPWR.n1493 VPWR.t1343 983.14
R472 VPWR.t1094 VPWR.n1506 983.14
R473 VPWR.n1507 VPWR.t1216 983.14
R474 VPWR.t1357 VPWR.n1520 983.14
R475 VPWR.n1521 VPWR.t1373 983.14
R476 VPWR.n1536 VPWR.t1116 983.14
R477 VPWR.n1535 VPWR.t1246 983.14
R478 VPWR.n1761 VPWR.t1287 983.14
R479 VPWR.n1760 VPWR.t1110 983.14
R480 VPWR.n1749 VPWR.t1160 983.14
R481 VPWR.t1268 VPWR.n1791 983.14
R482 VPWR.t1274 VPWR.n2506 983.14
R483 VPWR.n2507 VPWR.t1386 983.14
R484 VPWR.t1151 VPWR.n2518 983.14
R485 VPWR.n2519 VPWR.t1259 983.14
R486 VPWR.t1271 VPWR.n2530 983.14
R487 VPWR.n2531 VPWR.t1427 983.14
R488 VPWR.t1148 VPWR.n2542 983.14
R489 VPWR.n2543 VPWR.t1308 983.14
R490 VPWR.t1324 VPWR.n2554 983.14
R491 VPWR.n2555 VPWR.t1454 983.14
R492 VPWR.t1198 VPWR.n2566 983.14
R493 VPWR.n2567 VPWR.t1228 983.14
R494 VPWR.t1078 VPWR.n2578 983.14
R495 VPWR.n2579 VPWR.t1097 983.14
R496 VPWR.t1222 VPWR.n2590 983.14
R497 VPWR.n1594 VPWR.t1157 983.14
R498 VPWR.n1593 VPWR.t1262 983.14
R499 VPWR.t1424 VPWR.n1182 983.14
R500 VPWR.t1142 VPWR.n1185 983.14
R501 VPWR.n1220 VPWR.t1154 983.14
R502 VPWR.n1219 VPWR.t1313 983.14
R503 VPWR.n1216 VPWR.t1421 983.14
R504 VPWR.n1213 VPWR.t1182 983.14
R505 VPWR.n1205 VPWR.t1208 983.14
R506 VPWR.n1202 VPWR.t1335 983.14
R507 VPWR.n1199 VPWR.t1081 983.14
R508 VPWR.n1191 VPWR.t1102 983.14
R509 VPWR.n1188 VPWR.t1340 983.14
R510 VPWR.n1740 VPWR.t1368 983.14
R511 VPWR.n1739 VPWR.t1084 983.14
R512 VPWR.n1308 VPWR.t1889 877.144
R513 VPWR.n2723 VPWR.t504 877.144
R514 VPWR.n2843 VPWR.n2822 857.648
R515 VPWR.n1122 VPWR.t1390 738.074
R516 VPWR.n99 VPWR.t1130 738.074
R517 VPWR.n290 VPWR.t567 738.074
R518 VPWR.n68 VPWR.t1199 738.074
R519 VPWR.n346 VPWR.t924 738.074
R520 VPWR.n98 VPWR.t1275 738.074
R521 VPWR.n963 VPWR.t581 738.074
R522 VPWR.n356 VPWR.t573 738.074
R523 VPWR.n357 VPWR.t1744 738.074
R524 VPWR.n318 VPWR.t1851 738.074
R525 VPWR.n75 VPWR.t1309 738.074
R526 VPWR.n971 VPWR.t1585 738.074
R527 VPWR.n369 VPWR.t274 738.074
R528 VPWR.n322 VPWR.t198 738.074
R529 VPWR.n80 VPWR.t1149 738.074
R530 VPWR.n932 VPWR.t569 738.074
R531 VPWR.n933 VPWR.t436 738.074
R532 VPWR.n936 VPWR.t698 738.074
R533 VPWR.n387 VPWR.t563 738.074
R534 VPWR.n391 VPWR.t289 738.074
R535 VPWR.n395 VPWR.t727 738.074
R536 VPWR.n365 VPWR.t751 738.074
R537 VPWR.n330 VPWR.t975 738.074
R538 VPWR.n86 VPWR.t1272 738.074
R539 VPWR.n937 VPWR.t1490 738.074
R540 VPWR.n403 VPWR.t1577 738.074
R541 VPWR.n364 VPWR.t1730 738.074
R542 VPWR.n334 VPWR.t1722 738.074
R543 VPWR.n87 VPWR.t1260 738.074
R544 VPWR.n481 VPWR.t553 738.074
R545 VPWR.n480 VPWR.t1843 738.074
R546 VPWR.n477 VPWR.t914 738.074
R547 VPWR.n476 VPWR.t1520 738.074
R548 VPWR.n472 VPWR.t850 738.074
R549 VPWR.n469 VPWR.t945 738.074
R550 VPWR.n468 VPWR.t301 738.074
R551 VPWR.n465 VPWR.t458 738.074
R552 VPWR.n464 VPWR.t408 738.074
R553 VPWR.n461 VPWR.t65 738.074
R554 VPWR.n460 VPWR.t644 738.074
R555 VPWR.n457 VPWR.t1008 738.074
R556 VPWR.n456 VPWR.t99 738.074
R557 VPWR.n453 VPWR.t1550 738.074
R558 VPWR.n452 VPWR.t1059 738.074
R559 VPWR.n473 VPWR.t154 738.074
R560 VPWR.n482 VPWR.t565 738.074
R561 VPWR.n538 VPWR.t922 738.074
R562 VPWR.n534 VPWR.t1668 738.074
R563 VPWR.n530 VPWR.t1498 738.074
R564 VPWR.n522 VPWR.t404 738.074
R565 VPWR.n518 VPWR.t784 738.074
R566 VPWR.n514 VPWR.t196 738.074
R567 VPWR.n510 VPWR.t146 738.074
R568 VPWR.n506 VPWR.t450 738.074
R569 VPWR.n502 VPWR.t329 738.074
R570 VPWR.n498 VPWR.t998 738.074
R571 VPWR.n494 VPWR.t216 738.074
R572 VPWR.n490 VPWR.t1788 738.074
R573 VPWR.n486 VPWR.t353 738.074
R574 VPWR.n483 VPWR.t25 738.074
R575 VPWR.n526 VPWR.t132 738.074
R576 VPWR.n548 VPWR.t579 738.074
R577 VPWR.n549 VPWR.t1558 738.074
R578 VPWR.n552 VPWR.t1579 738.074
R579 VPWR.n553 VPWR.t1474 738.074
R580 VPWR.n557 VPWR.t1875 738.074
R581 VPWR.n560 VPWR.t1754 738.074
R582 VPWR.n561 VPWR.t5 738.074
R583 VPWR.n564 VPWR.t1704 738.074
R584 VPWR.n565 VPWR.t140 738.074
R585 VPWR.n568 VPWR.t763 738.074
R586 VPWR.n569 VPWR.t393 738.074
R587 VPWR.n572 VPWR.t670 738.074
R588 VPWR.n573 VPWR.t878 738.074
R589 VPWR.n576 VPWR.t599 738.074
R590 VPWR.n577 VPWR.t226 738.074
R591 VPWR.n556 VPWR.t321 738.074
R592 VPWR.n579 VPWR.t571 738.074
R593 VPWR.n583 VPWR.t1742 738.074
R594 VPWR.n587 VPWR.t702 738.074
R595 VPWR.n591 VPWR.t1488 738.074
R596 VPWR.n599 VPWR.t749 738.074
R597 VPWR.n603 VPWR.t794 738.074
R598 VPWR.n607 VPWR.t272 738.074
R599 VPWR.n611 VPWR.t1855 738.074
R600 VPWR.n615 VPWR.t660 738.074
R601 VPWR.n619 VPWR.t335 738.074
R602 VPWR.n623 VPWR.t1627 738.074
R603 VPWR.n627 VPWR.t890 738.074
R604 VPWR.n631 VPWR.t1796 738.074
R605 VPWR.n635 VPWR.t638 738.074
R606 VPWR.n578 VPWR.t31 738.074
R607 VPWR.n595 VPWR.t1726 738.074
R608 VPWR.n673 VPWR.t559 738.074
R609 VPWR.n672 VPWR.t285 738.074
R610 VPWR.n669 VPWR.t723 738.074
R611 VPWR.n668 VPWR.t1510 738.074
R612 VPWR.n664 VPWR.t1076 738.074
R613 VPWR.n661 VPWR.t1678 738.074
R614 VPWR.n660 VPWR.t311 738.074
R615 VPWR.n657 VPWR.t417 738.074
R616 VPWR.n656 VPWR.t868 738.074
R617 VPWR.n653 VPWR.t1532 738.074
R618 VPWR.n652 VPWR.t826 738.074
R619 VPWR.n649 VPWR.t1597 738.074
R620 VPWR.n648 VPWR.t256 738.074
R621 VPWR.n645 VPWR.t357 738.074
R622 VPWR.n644 VPWR.t1716 738.074
R623 VPWR.n665 VPWR.t1816 738.074
R624 VPWR.n674 VPWR.t551 738.074
R625 VPWR.n730 VPWR.t634 738.074
R626 VPWR.n726 VPWR.t912 738.074
R627 VPWR.n722 VPWR.t1522 738.074
R628 VPWR.n714 VPWR.t747 738.074
R629 VPWR.n710 VPWR.t943 738.074
R630 VPWR.n706 VPWR.t299 738.074
R631 VPWR.n702 VPWR.t204 738.074
R632 VPWR.n698 VPWR.t406 738.074
R633 VPWR.n694 VPWR.t63 738.074
R634 VPWR.n690 VPWR.t597 738.074
R635 VPWR.n686 VPWR.t1006 738.074
R636 VPWR.n682 VPWR.t97 738.074
R637 VPWR.n678 VPWR.t1057 738.074
R638 VPWR.n675 VPWR.t236 738.074
R639 VPWR.n718 VPWR.t152 738.074
R640 VPWR.n740 VPWR.t555 738.074
R641 VPWR.n741 VPWR.t820 738.074
R642 VPWR.n744 VPWR.t1839 738.074
R643 VPWR.n745 VPWR.t1516 738.074
R644 VPWR.n749 VPWR.t856 738.074
R645 VPWR.n752 VPWR.t951 738.074
R646 VPWR.n753 VPWR.t307 738.074
R647 VPWR.n756 VPWR.t156 738.074
R648 VPWR.n757 VPWR.t864 738.074
R649 VPWR.n760 VPWR.t71 738.074
R650 VPWR.n761 VPWR.t1915 738.074
R651 VPWR.n764 VPWR.t208 738.074
R652 VPWR.n765 VPWR.t246 738.074
R653 VPWR.n768 VPWR.t585 738.074
R654 VPWR.n769 VPWR.t1061 738.074
R655 VPWR.n748 VPWR.t1806 738.074
R656 VPWR.n771 VPWR.t577 738.074
R657 VPWR.n775 VPWR.t1556 738.074
R658 VPWR.n779 VPWR.t680 738.074
R659 VPWR.n783 VPWR.t1476 738.074
R660 VPWR.n791 VPWR.t1873 738.074
R661 VPWR.n795 VPWR.t960 738.074
R662 VPWR.n799 VPWR.t3 738.074
R663 VPWR.n803 VPWR.t1700 738.074
R664 VPWR.n807 VPWR.t138 738.074
R665 VPWR.n811 VPWR.t761 738.074
R666 VPWR.n815 VPWR.t391 738.074
R667 VPWR.n819 VPWR.t778 738.074
R668 VPWR.n823 VPWR.t874 738.074
R669 VPWR.n827 VPWR.t387 738.074
R670 VPWR.n770 VPWR.t222 738.074
R671 VPWR.n787 VPWR.t317 738.074
R672 VPWR.n865 VPWR.t561 738.074
R673 VPWR.n864 VPWR.t287 738.074
R674 VPWR.n861 VPWR.t725 738.074
R675 VPWR.n860 VPWR.t1508 738.074
R676 VPWR.n856 VPWR.t295 738.074
R677 VPWR.n853 VPWR.t1680 738.074
R678 VPWR.n852 VPWR.t186 738.074
R679 VPWR.n849 VPWR.t419 738.074
R680 VPWR.n848 VPWR.t1818 738.074
R681 VPWR.n845 VPWR.t1534 738.074
R682 VPWR.n844 VPWR.t828 738.074
R683 VPWR.n841 VPWR.t1599 738.074
R684 VPWR.n840 VPWR.t258 738.074
R685 VPWR.n837 VPWR.t359 738.074
R686 VPWR.n836 VPWR.t1718 738.074
R687 VPWR.n857 VPWR.t1573 738.074
R688 VPWR.n866 VPWR.t575 738.074
R689 VPWR.n922 VPWR.t1554 738.074
R690 VPWR.n918 VPWR.t678 738.074
R691 VPWR.n914 VPWR.t1478 738.074
R692 VPWR.n906 VPWR.t1871 738.074
R693 VPWR.n902 VPWR.t958 738.074
R694 VPWR.n898 VPWR.t1 738.074
R695 VPWR.n894 VPWR.t1859 738.074
R696 VPWR.n890 VPWR.t136 738.074
R697 VPWR.n886 VPWR.t759 738.074
R698 VPWR.n882 VPWR.t389 738.074
R699 VPWR.n878 VPWR.t776 738.074
R700 VPWR.n874 VPWR.t870 738.074
R701 VPWR.n870 VPWR.t385 738.074
R702 VPWR.n867 VPWR.t220 738.074
R703 VPWR.n910 VPWR.t315 738.074
R704 VPWR.n940 VPWR.t1724 738.074
R705 VPWR.n979 VPWR.t327 738.074
R706 VPWR.n1179 VPWR.t1143 738.074
R707 VPWR.n399 VPWR.t1506 738.074
R708 VPWR.n361 VPWR.t1486 738.074
R709 VPWR.n338 VPWR.t1494 738.074
R710 VPWR.n92 VPWR.t1152 738.074
R711 VPWR.n975 VPWR.t1468 738.074
R712 VPWR.n1183 VPWR.t1425 738.074
R713 VPWR.n941 VPWR.t979 738.074
R714 VPWR.n983 VPWR.t741 738.074
R715 VPWR.n1217 VPWR.t1155 738.074
R716 VPWR.n407 VPWR.t297 738.074
R717 VPWR.n415 VPWR.t188 738.074
R718 VPWR.n419 VPWR.t421 738.074
R719 VPWR.n423 VPWR.t1820 738.074
R720 VPWR.n427 VPWR.t1536 738.074
R721 VPWR.n431 VPWR.t830 738.074
R722 VPWR.n435 VPWR.t1601 738.074
R723 VPWR.n439 VPWR.t260 738.074
R724 VPWR.n443 VPWR.t361 738.074
R725 VPWR.n386 VPWR.t19 738.074
R726 VPWR.n411 VPWR.t798 738.074
R727 VPWR.n368 VPWR.t796 738.074
R728 VPWR.n326 VPWR.t786 738.074
R729 VPWR.n81 VPWR.t1428 738.074
R730 VPWR.n987 VPWR.t1760 738.074
R731 VPWR.n1214 VPWR.t1314 738.074
R732 VPWR.n944 VPWR.t790 738.074
R733 VPWR.n948 VPWR.t1853 738.074
R734 VPWR.n949 VPWR.t456 738.074
R735 VPWR.n952 VPWR.t333 738.074
R736 VPWR.n953 VPWR.t1623 738.074
R737 VPWR.n956 VPWR.t888 738.074
R738 VPWR.n957 VPWR.t1794 738.074
R739 VPWR.n960 VPWR.t636 738.074
R740 VPWR.n961 VPWR.t29 738.074
R741 VPWR.n945 VPWR.t268 738.074
R742 VPWR.n991 VPWR.t11 738.074
R743 VPWR.n1206 VPWR.t1422 738.074
R744 VPWR.n360 VPWR.t704 738.074
R745 VPWR.n342 VPWR.t1670 738.074
R746 VPWR.n93 VPWR.t1387 738.074
R747 VPWR.n1180 VPWR.t1263 738.074
R748 VPWR.n995 VPWR.t1708 738.074
R749 VPWR.n1203 VPWR.t1183 738.074
R750 VPWR.n372 VPWR.t1857 738.074
R751 VPWR.n376 VPWR.t337 738.074
R752 VPWR.n377 VPWR.t1629 738.074
R753 VPWR.n380 VPWR.t892 738.074
R754 VPWR.n381 VPWR.t1798 738.074
R755 VPWR.n384 VPWR.t640 738.074
R756 VPWR.n385 VPWR.t168 738.074
R757 VPWR.n373 VPWR.t662 738.074
R758 VPWR.n314 VPWR.t452 738.074
R759 VPWR.n74 VPWR.t1325 738.074
R760 VPWR.n1200 VPWR.t1209 738.074
R761 VPWR.n999 VPWR.t180 738.074
R762 VPWR.n1003 VPWR.t765 738.074
R763 VPWR.n1007 VPWR.t591 738.074
R764 VPWR.n1011 VPWR.t672 738.074
R765 VPWR.n1015 VPWR.t89 738.074
R766 VPWR.n1019 VPWR.t642 738.074
R767 VPWR.n962 VPWR.t232 738.074
R768 VPWR.n967 VPWR.t626 738.074
R769 VPWR.n1123 VPWR.t1158 738.074
R770 VPWR.n310 VPWR.t331 738.074
R771 VPWR.n69 VPWR.t1455 738.074
R772 VPWR.n1192 VPWR.t1336 738.074
R773 VPWR.n1189 VPWR.t1082 738.074
R774 VPWR.n306 VPWR.t1000 738.074
R775 VPWR.n302 VPWR.t218 738.074
R776 VPWR.n294 VPWR.t355 738.074
R777 VPWR.n291 VPWR.t27 738.074
R778 VPWR.n298 VPWR.t1792 738.074
R779 VPWR.n1058 VPWR.t1341 738.074
R780 VPWR.n1186 VPWR.t1103 738.074
R781 VPWR.n63 VPWR.t1229 738.074
R782 VPWR.n62 VPWR.t1079 738.074
R783 VPWR.n57 VPWR.t1098 738.074
R784 VPWR.n56 VPWR.t1223 738.074
R785 VPWR.n1059 VPWR.t1369 738.074
R786 VPWR.n1061 VPWR.t1085 738.074
R787 VPWR.n2856 VPWR.n2821 702.354
R788 VPWR.n2856 VPWR.n2822 702.354
R789 VPWR.n2854 VPWR.n2853 702.354
R790 VPWR.n2854 VPWR.n2821 702.354
R791 VPWR.n2837 VPWR.n2828 702.354
R792 VPWR.n2850 VPWR.n2849 702.354
R793 VPWR.n2835 VPWR.n2828 702.354
R794 VPWR.n2815 VPWR.t1561 651.634
R795 VPWR.n2831 VPWR.t557 651.505
R796 VPWR.n2825 VPWR.t734 651.505
R797 VPWR.n2862 VPWR.t448 651.431
R798 VPWR.n1061 VPWR.t1212 646.071
R799 VPWR.n1122 VPWR.t1108 646.071
R800 VPWR.n1059 VPWR.t1361 646.071
R801 VPWR.n56 VPWR.t1328 646.071
R802 VPWR.n62 VPWR.t1452 646.071
R803 VPWR.n99 VPWR.t1237 646.071
R804 VPWR.n1053 VPWR.t95 646.071
R805 VPWR.n1231 VPWR.t1565 646.071
R806 VPWR.n298 VPWR.t1045 646.071
R807 VPWR.n290 VPWR.t1748 646.071
R808 VPWR.n306 VPWR.t896 646.071
R809 VPWR.n68 VPWR.t1191 646.071
R810 VPWR.n1153 VPWR.t771 646.071
R811 VPWR.n346 VPWR.t700 646.071
R812 VPWR.n98 VPWR.t1366 646.071
R813 VPWR.n967 VPWR.t910 646.071
R814 VPWR.n963 VPWR.t1845 646.071
R815 VPWR.n999 VPWR.t67 646.071
R816 VPWR.n373 VPWR.t538 646.071
R817 VPWR.n356 VPWR.t1563 646.071
R818 VPWR.n357 VPWR.t708 646.071
R819 VPWR.n372 VPWR.t668 646.071
R820 VPWR.n318 VPWR.t658 646.071
R821 VPWR.n75 VPWR.t1296 646.071
R822 VPWR.n971 VPWR.t1504 646.071
R823 VPWR.n369 VPWR.t200 646.071
R824 VPWR.n322 VPWR.t1702 646.071
R825 VPWR.n80 VPWR.t1168 646.071
R826 VPWR.n945 VPWR.t1706 646.071
R827 VPWR.n932 VPWR.t1750 646.071
R828 VPWR.n933 VPWR.t706 646.071
R829 VPWR.n936 VPWR.t1466 646.071
R830 VPWR.n944 VPWR.t276 646.071
R831 VPWR.n411 VPWR.t194 646.071
R832 VPWR.n387 VPWR.t920 646.071
R833 VPWR.n391 VPWR.t782 646.071
R834 VPWR.n395 VPWR.t1480 646.071
R835 VPWR.n407 VPWR.t804 646.071
R836 VPWR.n365 VPWR.t810 646.071
R837 VPWR.n330 VPWR.t792 646.071
R838 VPWR.n86 VPWR.t1409 646.071
R839 VPWR.n937 VPWR.t319 646.071
R840 VPWR.n403 VPWR.t82 646.071
R841 VPWR.n364 VPWR.t757 646.071
R842 VPWR.n334 VPWR.t981 646.071
R843 VPWR.n87 VPWR.t1254 646.071
R844 VPWR.n473 VPWR.t854 646.071
R845 VPWR.n481 VPWR.t822 646.071
R846 VPWR.n480 VPWR.t1837 646.071
R847 VPWR.n477 VPWR.t1500 646.071
R848 VPWR.n476 VPWR.t128 646.071
R849 VPWR.n472 VPWR.t949 646.071
R850 VPWR.n469 VPWR.t305 646.071
R851 VPWR.n468 VPWR.t214 646.071
R852 VPWR.n465 VPWR.t412 646.071
R853 VPWR.n464 VPWR.t73 646.071
R854 VPWR.n461 VPWR.t648 646.071
R855 VPWR.n460 VPWR.t210 646.071
R856 VPWR.n457 VPWR.t264 646.071
R857 VPWR.n456 VPWR.t587 646.071
R858 VPWR.n453 VPWR.t21 646.071
R859 VPWR.n452 VPWR.t1226 646.071
R860 VPWR.n526 VPWR.t977 646.071
R861 VPWR.n482 VPWR.t1746 646.071
R862 VPWR.n538 VPWR.t1672 646.071
R863 VPWR.n534 VPWR.t1472 646.071
R864 VPWR.n530 VPWR.t1831 646.071
R865 VPWR.n522 VPWR.t788 646.071
R866 VPWR.n518 VPWR.t266 646.071
R867 VPWR.n514 VPWR.t1698 646.071
R868 VPWR.n510 VPWR.t454 646.071
R869 VPWR.n506 VPWR.t339 646.071
R870 VPWR.n502 VPWR.t1002 646.071
R871 VPWR.n498 VPWR.t894 646.071
R872 VPWR.n494 VPWR.t872 646.071
R873 VPWR.n490 VPWR.t1043 646.071
R874 VPWR.n486 VPWR.t174 646.071
R875 VPWR.n483 VPWR.t1444 646.071
R876 VPWR.n556 VPWR.t743 646.071
R877 VPWR.n548 VPWR.t632 646.071
R878 VPWR.n549 VPWR.t1587 646.071
R879 VPWR.n552 VPWR.t1512 646.071
R880 VPWR.n553 VPWR.t1812 646.071
R881 VPWR.n557 VPWR.t1762 646.071
R882 VPWR.n560 VPWR.t13 646.071
R883 VPWR.n561 VPWR.t162 646.071
R884 VPWR.n564 VPWR.t182 646.071
R885 VPWR.n565 VPWR.t61 646.071
R886 VPWR.n568 VPWR.t593 646.071
R887 VPWR.n569 VPWR.t1004 646.071
R888 VPWR.n572 VPWR.t252 646.071
R889 VPWR.n573 VPWR.t1055 646.071
R890 VPWR.n576 VPWR.t1712 646.071
R891 VPWR.n577 VPWR.t1293 646.071
R892 VPWR.n595 VPWR.t755 646.071
R893 VPWR.n579 VPWR.t1752 646.071
R894 VPWR.n583 VPWR.t682 646.071
R895 VPWR.n587 VPWR.t1464 646.071
R896 VPWR.n591 VPWR.t323 646.071
R897 VPWR.n599 VPWR.t808 646.071
R898 VPWR.n603 VPWR.t278 646.071
R899 VPWR.n607 VPWR.t1710 646.071
R900 VPWR.n611 VPWR.t666 646.071
R901 VPWR.n615 VPWR.t536 646.071
R902 VPWR.n619 VPWR.t1633 646.071
R903 VPWR.n623 VPWR.t992 646.071
R904 VPWR.n627 VPWR.t91 646.071
R905 VPWR.n631 VPWR.t1049 646.071
R906 VPWR.n635 VPWR.t228 646.071
R907 VPWR.n578 VPWR.t1401 646.071
R908 VPWR.n665 VPWR.t78 646.071
R909 VPWR.n673 VPWR.t693 646.071
R910 VPWR.n672 VPWR.t729 646.071
R911 VPWR.n669 VPWR.t1484 646.071
R912 VPWR.n668 VPWR.t1728 646.071
R913 VPWR.n664 VPWR.t800 646.071
R914 VPWR.n661 VPWR.t190 646.071
R915 VPWR.n660 VPWR.t460 646.071
R916 VPWR.n657 VPWR.t1822 646.071
R917 VPWR.n656 VPWR.t1538 646.071
R918 VPWR.n653 VPWR.t832 646.071
R919 VPWR.n652 VPWR.t1736 646.071
R920 VPWR.n649 VPWR.t1800 646.071
R921 VPWR.n648 VPWR.t1544 646.071
R922 VPWR.n645 VPWR.t166 646.071
R923 VPWR.n644 VPWR.t1127 646.071
R924 VPWR.n718 VPWR.t852 646.071
R925 VPWR.n674 VPWR.t1847 646.071
R926 VPWR.n730 VPWR.t1835 646.071
R927 VPWR.n726 VPWR.t1502 646.071
R928 VPWR.n722 VPWR.t1575 646.071
R929 VPWR.n714 VPWR.t947 646.071
R930 VPWR.n710 VPWR.t303 646.071
R931 VPWR.n706 VPWR.t212 646.071
R932 VPWR.n702 VPWR.t410 646.071
R933 VPWR.n698 VPWR.t69 646.071
R934 VPWR.n694 VPWR.t646 646.071
R935 VPWR.n690 VPWR.t206 646.071
R936 VPWR.n686 VPWR.t262 646.071
R937 VPWR.n682 VPWR.t583 646.071
R938 VPWR.n678 VPWR.t1720 646.071
R939 VPWR.n675 VPWR.t1234 646.071
R940 VPWR.n748 VPWR.t1074 646.071
R941 VPWR.n740 VPWR.t824 646.071
R942 VPWR.n741 VPWR.t1841 646.071
R943 VPWR.n744 VPWR.t1492 646.071
R944 VPWR.n745 VPWR.t130 646.071
R945 VPWR.n749 VPWR.t1676 646.071
R946 VPWR.n752 VPWR.t309 646.071
R947 VPWR.n753 VPWR.t148 646.071
R948 VPWR.n756 VPWR.t866 646.071
R949 VPWR.n757 VPWR.t1530 646.071
R950 VPWR.n760 VPWR.t1917 646.071
R951 VPWR.n761 VPWR.t1595 646.071
R952 VPWR.n764 VPWR.t1790 646.071
R953 VPWR.n765 VPWR.t589 646.071
R954 VPWR.n768 VPWR.t23 646.071
R955 VPWR.n769 VPWR.t1194 646.071
R956 VPWR.n787 VPWR.t1879 646.071
R957 VPWR.n771 VPWR.t630 646.071
R958 VPWR.n775 VPWR.t1583 646.071
R959 VPWR.n779 VPWR.t1496 646.071
R960 VPWR.n783 VPWR.t1810 646.071
R961 VPWR.n791 VPWR.t1758 646.071
R962 VPWR.n795 VPWR.t9 646.071
R963 VPWR.n799 VPWR.t160 646.071
R964 VPWR.n803 VPWR.t178 646.071
R965 VPWR.n807 VPWR.t59 646.071
R966 VPWR.n811 VPWR.t397 646.071
R967 VPWR.n815 VPWR.t676 646.071
R968 VPWR.n819 VPWR.t250 646.071
R969 VPWR.n823 VPWR.t1053 646.071
R970 VPWR.n827 VPWR.t1065 646.071
R971 VPWR.n770 VPWR.t1299 646.071
R972 VPWR.n857 VPWR.t80 646.071
R973 VPWR.n865 VPWR.t918 646.071
R974 VPWR.n864 VPWR.t780 646.071
R975 VPWR.n861 VPWR.t1482 646.071
R976 VPWR.n860 VPWR.t1732 646.071
R977 VPWR.n856 VPWR.t802 646.071
R978 VPWR.n853 VPWR.t192 646.071
R979 VPWR.n852 VPWR.t462 646.071
R980 VPWR.n849 VPWR.t1824 646.071
R981 VPWR.n848 VPWR.t1540 646.071
R982 VPWR.n845 VPWR.t834 646.071
R983 VPWR.n844 VPWR.t1738 646.071
R984 VPWR.n841 VPWR.t1802 646.071
R985 VPWR.n840 VPWR.t1546 646.071
R986 VPWR.n837 VPWR.t170 646.071
R987 VPWR.n836 VPWR.t1122 646.071
R988 VPWR.n910 VPWR.t1877 646.071
R989 VPWR.n866 VPWR.t628 646.071
R990 VPWR.n922 VPWR.t1581 646.071
R991 VPWR.n918 VPWR.t1514 646.071
R992 VPWR.n914 VPWR.t1808 646.071
R993 VPWR.n906 VPWR.t1756 646.071
R994 VPWR.n902 VPWR.t7 646.071
R995 VPWR.n898 VPWR.t158 646.071
R996 VPWR.n894 VPWR.t142 646.071
R997 VPWR.n890 VPWR.t767 646.071
R998 VPWR.n886 VPWR.t395 646.071
R999 VPWR.n882 VPWR.t674 646.071
R1000 VPWR.n878 VPWR.t248 646.071
R1001 VPWR.n874 VPWR.t1051 646.071
R1002 VPWR.n870 VPWR.t1063 646.071
R1003 VPWR.n867 VPWR.t1306 646.071
R1004 VPWR.n940 VPWR.t753 646.071
R1005 VPWR.n979 VPWR.t745 646.071
R1006 VPWR.n1227 VPWR.t1881 646.071
R1007 VPWR.n1179 VPWR.t1138 646.071
R1008 VPWR.n399 VPWR.t1734 646.071
R1009 VPWR.n361 VPWR.t325 646.071
R1010 VPWR.n338 VPWR.t313 646.071
R1011 VPWR.n92 VPWR.t1146 646.071
R1012 VPWR.n975 VPWR.t1814 646.071
R1013 VPWR.n1485 VPWR.t150 646.071
R1014 VPWR.n1183 VPWR.t1417 646.071
R1015 VPWR.n941 VPWR.t806 646.071
R1016 VPWR.n983 VPWR.t1764 646.071
R1017 VPWR.n1173 VPWR.t812 646.071
R1018 VPWR.n1217 VPWR.t1285 646.071
R1019 VPWR.n415 VPWR.t464 646.071
R1020 VPWR.n419 VPWR.t1826 646.071
R1021 VPWR.n423 VPWR.t1542 646.071
R1022 VPWR.n427 VPWR.t836 646.071
R1023 VPWR.n431 VPWR.t1740 646.071
R1024 VPWR.n435 VPWR.t1804 646.071
R1025 VPWR.n439 VPWR.t1548 646.071
R1026 VPWR.n443 VPWR.t172 646.071
R1027 VPWR.n386 VPWR.t1114 646.071
R1028 VPWR.n368 VPWR.t280 646.071
R1029 VPWR.n326 VPWR.t270 646.071
R1030 VPWR.n81 VPWR.t1133 646.071
R1031 VPWR.n987 VPWR.t15 646.071
R1032 VPWR.n1169 VPWR.t282 646.071
R1033 VPWR.n1214 VPWR.t1393 646.071
R1034 VPWR.n948 VPWR.t664 646.071
R1035 VPWR.n949 VPWR.t534 646.071
R1036 VPWR.n952 VPWR.t1631 646.071
R1037 VPWR.n953 VPWR.t898 646.071
R1038 VPWR.n956 VPWR.t880 646.071
R1039 VPWR.n957 VPWR.t1047 646.071
R1040 VPWR.n960 VPWR.t224 646.071
R1041 VPWR.n961 VPWR.t1414 646.071
R1042 VPWR.n991 VPWR.t164 646.071
R1043 VPWR.n1163 VPWR.t202 646.071
R1044 VPWR.n1206 VPWR.t1433 646.071
R1045 VPWR.n360 VPWR.t1462 646.071
R1046 VPWR.n342 VPWR.t1470 646.071
R1047 VPWR.n93 VPWR.t1384 646.071
R1048 VPWR.n1479 VPWR.t1518 646.071
R1049 VPWR.n1180 VPWR.t1257 646.071
R1050 VPWR.n995 VPWR.t184 646.071
R1051 VPWR.n1159 VPWR.t1069 646.071
R1052 VPWR.n1203 VPWR.t1178 646.071
R1053 VPWR.n376 VPWR.t769 646.071
R1054 VPWR.n377 VPWR.t994 646.071
R1055 VPWR.n380 VPWR.t93 646.071
R1056 VPWR.n381 VPWR.t1022 646.071
R1057 VPWR.n384 VPWR.t230 646.071
R1058 VPWR.n385 VPWR.t1396 646.071
R1059 VPWR.n314 VPWR.t341 646.071
R1060 VPWR.n74 VPWR.t1406 646.071
R1061 VPWR.n1149 VPWR.t540 646.071
R1062 VPWR.n1200 VPWR.t1282 646.071
R1063 VPWR.n1003 VPWR.t595 646.071
R1064 VPWR.n1007 VPWR.t1010 646.071
R1065 VPWR.n1011 VPWR.t254 646.071
R1066 VPWR.n1015 VPWR.t1552 646.071
R1067 VPWR.n1019 VPWR.t1714 646.071
R1068 VPWR.n962 VPWR.t1266 646.071
R1069 VPWR.n1472 VPWR.t710 646.071
R1070 VPWR.n1123 VPWR.t1244 646.071
R1071 VPWR.n310 VPWR.t1625 646.071
R1072 VPWR.n69 VPWR.t1173 646.071
R1073 VPWR.n1192 VPWR.t1441 646.071
R1074 VPWR.n1049 VPWR.t996 646.071
R1075 VPWR.n1189 VPWR.t1460 646.071
R1076 VPWR.n302 VPWR.t876 646.071
R1077 VPWR.n294 VPWR.t176 646.071
R1078 VPWR.n291 VPWR.t1436 646.071
R1079 VPWR.n1058 VPWR.t1333 646.071
R1080 VPWR.n1748 VPWR.t1024 646.071
R1081 VPWR.n1036 VPWR.t234 646.071
R1082 VPWR.n1032 VPWR.t1377 646.071
R1083 VPWR.n1186 VPWR.t1204 646.071
R1084 VPWR.n63 VPWR.t1319 646.071
R1085 VPWR.n57 VPWR.t1092 646.071
R1086 VPWR.n1230 VPWR.t1186 642.13
R1087 VPWR.n1152 VPWR.t1117 642.13
R1088 VPWR.n1226 VPWR.t1322 642.13
R1089 VPWR.n1484 VPWR.t1220 642.13
R1090 VPWR.n1172 VPWR.t1344 642.13
R1091 VPWR.n1168 VPWR.t1095 642.13
R1092 VPWR.n1162 VPWR.t1217 642.13
R1093 VPWR.n1478 VPWR.t1449 642.13
R1094 VPWR.n1158 VPWR.t1358 642.13
R1095 VPWR.n1148 VPWR.t1374 642.13
R1096 VPWR.n1471 VPWR.t1347 642.13
R1097 VPWR.n1048 VPWR.t1247 642.13
R1098 VPWR.n1747 VPWR.t1111 642.13
R1099 VPWR.n1035 VPWR.t1161 642.13
R1100 VPWR.n1031 VPWR.t1269 642.13
R1101 VPWR.n1052 VPWR.t1288 642.13
R1102 VPWR.n2309 VPWR.t821 629.652
R1103 VPWR.n2310 VPWR.t1836 629.652
R1104 VPWR.n2319 VPWR.t1499 629.652
R1105 VPWR.n2320 VPWR.t127 629.652
R1106 VPWR.n2329 VPWR.t853 629.652
R1107 VPWR.n2330 VPWR.t948 629.652
R1108 VPWR.n2339 VPWR.t304 629.652
R1109 VPWR.n2340 VPWR.t213 629.652
R1110 VPWR.n2349 VPWR.t411 629.652
R1111 VPWR.n2350 VPWR.t72 629.652
R1112 VPWR.n2359 VPWR.t647 629.652
R1113 VPWR.n2360 VPWR.t209 629.652
R1114 VPWR.n2369 VPWR.t263 629.652
R1115 VPWR.n2370 VPWR.t586 629.652
R1116 VPWR.n2379 VPWR.t20 629.652
R1117 VPWR.n542 VPWR.t1745 629.652
R1118 VPWR.t1671 VPWR.n541 629.652
R1119 VPWR.t1471 VPWR.n537 629.652
R1120 VPWR.t1830 VPWR.n533 629.652
R1121 VPWR.t976 VPWR.n529 629.652
R1122 VPWR.t787 VPWR.n525 629.652
R1123 VPWR.t265 VPWR.n521 629.652
R1124 VPWR.t1697 VPWR.n517 629.652
R1125 VPWR.t453 VPWR.n513 629.652
R1126 VPWR.t338 VPWR.n509 629.652
R1127 VPWR.t1001 VPWR.n505 629.652
R1128 VPWR.t893 VPWR.n501 629.652
R1129 VPWR.t871 VPWR.n497 629.652
R1130 VPWR.t1042 VPWR.n493 629.652
R1131 VPWR.t173 VPWR.n489 629.652
R1132 VPWR.n2281 VPWR.t631 629.652
R1133 VPWR.t1586 VPWR.n2280 629.652
R1134 VPWR.n2271 VPWR.t1511 629.652
R1135 VPWR.t1811 VPWR.n2270 629.652
R1136 VPWR.n2261 VPWR.t742 629.652
R1137 VPWR.t1761 VPWR.n2260 629.652
R1138 VPWR.n2251 VPWR.t12 629.652
R1139 VPWR.t161 VPWR.n2250 629.652
R1140 VPWR.n2241 VPWR.t181 629.652
R1141 VPWR.t60 VPWR.n2240 629.652
R1142 VPWR.n2231 VPWR.t592 629.652
R1143 VPWR.t1003 VPWR.n2230 629.652
R1144 VPWR.n2221 VPWR.t251 629.652
R1145 VPWR.t1054 VPWR.n2220 629.652
R1146 VPWR.n2211 VPWR.t1711 629.652
R1147 VPWR.n582 VPWR.t1751 629.652
R1148 VPWR.n586 VPWR.t681 629.652
R1149 VPWR.n590 VPWR.t1463 629.652
R1150 VPWR.n594 VPWR.t322 629.652
R1151 VPWR.n598 VPWR.t754 629.652
R1152 VPWR.n602 VPWR.t807 629.652
R1153 VPWR.n606 VPWR.t277 629.652
R1154 VPWR.n610 VPWR.t1709 629.652
R1155 VPWR.n614 VPWR.t665 629.652
R1156 VPWR.n618 VPWR.t535 629.652
R1157 VPWR.n622 VPWR.t1632 629.652
R1158 VPWR.n626 VPWR.t991 629.652
R1159 VPWR.n630 VPWR.t90 629.652
R1160 VPWR.n634 VPWR.t1048 629.652
R1161 VPWR.n638 VPWR.t227 629.652
R1162 VPWR.n2113 VPWR.t692 629.652
R1163 VPWR.n2114 VPWR.t728 629.652
R1164 VPWR.n2123 VPWR.t1483 629.652
R1165 VPWR.n2124 VPWR.t1727 629.652
R1166 VPWR.n2133 VPWR.t77 629.652
R1167 VPWR.n2134 VPWR.t799 629.652
R1168 VPWR.n2143 VPWR.t189 629.652
R1169 VPWR.n2144 VPWR.t459 629.652
R1170 VPWR.n2153 VPWR.t1821 629.652
R1171 VPWR.n2154 VPWR.t1537 629.652
R1172 VPWR.n2163 VPWR.t831 629.652
R1173 VPWR.n2164 VPWR.t1735 629.652
R1174 VPWR.n2173 VPWR.t1799 629.652
R1175 VPWR.n2174 VPWR.t1543 629.652
R1176 VPWR.n2183 VPWR.t165 629.652
R1177 VPWR.n734 VPWR.t1846 629.652
R1178 VPWR.t1834 VPWR.n733 629.652
R1179 VPWR.t1501 VPWR.n729 629.652
R1180 VPWR.t1574 VPWR.n725 629.652
R1181 VPWR.t851 VPWR.n721 629.652
R1182 VPWR.t946 VPWR.n717 629.652
R1183 VPWR.t302 VPWR.n713 629.652
R1184 VPWR.t211 VPWR.n709 629.652
R1185 VPWR.t409 VPWR.n705 629.652
R1186 VPWR.t68 VPWR.n701 629.652
R1187 VPWR.t645 VPWR.n697 629.652
R1188 VPWR.t205 VPWR.n693 629.652
R1189 VPWR.t261 VPWR.n689 629.652
R1190 VPWR.t582 VPWR.n685 629.652
R1191 VPWR.t1719 VPWR.n681 629.652
R1192 VPWR.n2085 VPWR.t823 629.652
R1193 VPWR.t1840 VPWR.n2084 629.652
R1194 VPWR.n2075 VPWR.t1491 629.652
R1195 VPWR.t129 VPWR.n2074 629.652
R1196 VPWR.n2065 VPWR.t1073 629.652
R1197 VPWR.t1675 VPWR.n2064 629.652
R1198 VPWR.n2055 VPWR.t308 629.652
R1199 VPWR.t147 VPWR.n2054 629.652
R1200 VPWR.n2045 VPWR.t865 629.652
R1201 VPWR.t1529 VPWR.n2044 629.652
R1202 VPWR.n2035 VPWR.t1916 629.652
R1203 VPWR.t1594 VPWR.n2034 629.652
R1204 VPWR.n2025 VPWR.t1789 629.652
R1205 VPWR.t588 VPWR.n2024 629.652
R1206 VPWR.n2015 VPWR.t22 629.652
R1207 VPWR.n774 VPWR.t629 629.652
R1208 VPWR.n778 VPWR.t1582 629.652
R1209 VPWR.n782 VPWR.t1495 629.652
R1210 VPWR.n786 VPWR.t1809 629.652
R1211 VPWR.n790 VPWR.t1878 629.652
R1212 VPWR.n794 VPWR.t1757 629.652
R1213 VPWR.n798 VPWR.t8 629.652
R1214 VPWR.n802 VPWR.t159 629.652
R1215 VPWR.n806 VPWR.t177 629.652
R1216 VPWR.n810 VPWR.t58 629.652
R1217 VPWR.n814 VPWR.t396 629.652
R1218 VPWR.n818 VPWR.t675 629.652
R1219 VPWR.n822 VPWR.t249 629.652
R1220 VPWR.n826 VPWR.t1052 629.652
R1221 VPWR.n830 VPWR.t1064 629.652
R1222 VPWR.n1917 VPWR.t917 629.652
R1223 VPWR.n1918 VPWR.t779 629.652
R1224 VPWR.n1927 VPWR.t1481 629.652
R1225 VPWR.n1928 VPWR.t1731 629.652
R1226 VPWR.n1937 VPWR.t79 629.652
R1227 VPWR.n1938 VPWR.t801 629.652
R1228 VPWR.n1947 VPWR.t191 629.652
R1229 VPWR.n1948 VPWR.t461 629.652
R1230 VPWR.n1957 VPWR.t1823 629.652
R1231 VPWR.n1958 VPWR.t1539 629.652
R1232 VPWR.n1967 VPWR.t833 629.652
R1233 VPWR.n1968 VPWR.t1737 629.652
R1234 VPWR.n1977 VPWR.t1801 629.652
R1235 VPWR.n1978 VPWR.t1545 629.652
R1236 VPWR.n1987 VPWR.t169 629.652
R1237 VPWR.n926 VPWR.t627 629.652
R1238 VPWR.t1580 VPWR.n925 629.652
R1239 VPWR.t1513 VPWR.n921 629.652
R1240 VPWR.t1807 VPWR.n917 629.652
R1241 VPWR.t1876 VPWR.n913 629.652
R1242 VPWR.t1755 VPWR.n909 629.652
R1243 VPWR.t6 VPWR.n905 629.652
R1244 VPWR.t157 VPWR.n901 629.652
R1245 VPWR.t141 VPWR.n897 629.652
R1246 VPWR.t766 VPWR.n893 629.652
R1247 VPWR.t394 VPWR.n889 629.652
R1248 VPWR.t673 VPWR.n885 629.652
R1249 VPWR.t247 VPWR.n881 629.652
R1250 VPWR.t1050 VPWR.n877 629.652
R1251 VPWR.t1062 VPWR.n873 629.652
R1252 VPWR.n390 VPWR.t919 629.652
R1253 VPWR.n394 VPWR.t781 629.652
R1254 VPWR.n398 VPWR.t1479 629.652
R1255 VPWR.n402 VPWR.t1733 629.652
R1256 VPWR.n406 VPWR.t81 629.652
R1257 VPWR.n410 VPWR.t803 629.652
R1258 VPWR.n414 VPWR.t193 629.652
R1259 VPWR.n418 VPWR.t463 629.652
R1260 VPWR.n422 VPWR.t1825 629.652
R1261 VPWR.n426 VPWR.t1541 629.652
R1262 VPWR.n430 VPWR.t835 629.652
R1263 VPWR.n434 VPWR.t1739 629.652
R1264 VPWR.n438 VPWR.t1803 629.652
R1265 VPWR.n442 VPWR.t1547 629.652
R1266 VPWR.n446 VPWR.t171 629.652
R1267 VPWR.n1889 VPWR.t1749 629.652
R1268 VPWR.t705 VPWR.n1888 629.652
R1269 VPWR.n1879 VPWR.t1465 629.652
R1270 VPWR.t318 VPWR.n1878 629.652
R1271 VPWR.n1869 VPWR.t752 629.652
R1272 VPWR.t805 VPWR.n1868 629.652
R1273 VPWR.n1859 VPWR.t275 629.652
R1274 VPWR.t1705 VPWR.n1858 629.652
R1275 VPWR.n1849 VPWR.t663 629.652
R1276 VPWR.t533 VPWR.n1848 629.652
R1277 VPWR.n1839 VPWR.t1630 629.652
R1278 VPWR.t897 VPWR.n1838 629.652
R1279 VPWR.n1829 VPWR.t879 629.652
R1280 VPWR.t1046 VPWR.n1828 629.652
R1281 VPWR.n1819 VPWR.t223 629.652
R1282 VPWR.n2477 VPWR.t1562 629.652
R1283 VPWR.t707 VPWR.n2476 629.652
R1284 VPWR.n2467 VPWR.t1461 629.652
R1285 VPWR.t324 VPWR.n2466 629.652
R1286 VPWR.n2457 VPWR.t756 629.652
R1287 VPWR.t809 VPWR.n2456 629.652
R1288 VPWR.n2447 VPWR.t279 629.652
R1289 VPWR.t199 VPWR.n2446 629.652
R1290 VPWR.n2437 VPWR.t667 629.652
R1291 VPWR.t537 VPWR.n2436 629.652
R1292 VPWR.n2427 VPWR.t768 629.652
R1293 VPWR.t993 VPWR.n2426 629.652
R1294 VPWR.n2417 VPWR.t92 629.652
R1295 VPWR.t1021 VPWR.n2416 629.652
R1296 VPWR.n2407 VPWR.t229 629.652
R1297 VPWR.n966 VPWR.t1844 629.652
R1298 VPWR.n970 VPWR.t909 629.652
R1299 VPWR.n974 VPWR.t1503 629.652
R1300 VPWR.n978 VPWR.t1813 629.652
R1301 VPWR.n982 VPWR.t744 629.652
R1302 VPWR.n986 VPWR.t1763 629.652
R1303 VPWR.n990 VPWR.t14 629.652
R1304 VPWR.n994 VPWR.t163 629.652
R1305 VPWR.n998 VPWR.t183 629.652
R1306 VPWR.n1002 VPWR.t66 629.652
R1307 VPWR.n1006 VPWR.t594 629.652
R1308 VPWR.n1010 VPWR.t1009 629.652
R1309 VPWR.n1014 VPWR.t253 629.652
R1310 VPWR.n1018 VPWR.t1551 629.652
R1311 VPWR.n1022 VPWR.t1713 629.652
R1312 VPWR.n350 VPWR.t1747 629.652
R1313 VPWR.t699 VPWR.n349 629.652
R1314 VPWR.t1469 VPWR.n345 629.652
R1315 VPWR.t312 VPWR.n341 629.652
R1316 VPWR.t980 VPWR.n337 629.652
R1317 VPWR.t791 VPWR.n333 629.652
R1318 VPWR.t269 VPWR.n329 629.652
R1319 VPWR.t1701 VPWR.n325 629.652
R1320 VPWR.t657 VPWR.n321 629.652
R1321 VPWR.t340 VPWR.n317 629.652
R1322 VPWR.t1624 VPWR.n313 629.652
R1323 VPWR.t895 VPWR.n309 629.652
R1324 VPWR.t875 VPWR.n305 629.652
R1325 VPWR.t1044 VPWR.n301 629.652
R1326 VPWR.t175 VPWR.n297 629.652
R1327 VPWR.n1468 VPWR.t1564 629.652
R1328 VPWR.n1475 VPWR.t709 629.652
R1329 VPWR.n1481 VPWR.t1517 629.652
R1330 VPWR.n1492 VPWR.t149 629.652
R1331 VPWR.n1493 VPWR.t1880 629.652
R1332 VPWR.n1506 VPWR.t811 629.652
R1333 VPWR.n1507 VPWR.t281 629.652
R1334 VPWR.n1520 VPWR.t201 629.652
R1335 VPWR.n1521 VPWR.t1068 629.652
R1336 VPWR.n1536 VPWR.t539 629.652
R1337 VPWR.t770 VPWR.n1535 629.652
R1338 VPWR.n1761 VPWR.t995 629.652
R1339 VPWR.t94 VPWR.n1760 629.652
R1340 VPWR.n1749 VPWR.t1023 629.652
R1341 VPWR.n1791 VPWR.t233 629.652
R1342 VPWR.n2506 VPWR.t1236 629.652
R1343 VPWR.n2507 VPWR.t1365 629.652
R1344 VPWR.n2518 VPWR.t1383 629.652
R1345 VPWR.n2519 VPWR.t1145 629.652
R1346 VPWR.n2530 VPWR.t1253 629.652
R1347 VPWR.n2531 VPWR.t1408 629.652
R1348 VPWR.n2542 VPWR.t1132 629.652
R1349 VPWR.n2543 VPWR.t1167 629.652
R1350 VPWR.n2554 VPWR.t1295 629.652
R1351 VPWR.n2555 VPWR.t1405 629.652
R1352 VPWR.n2566 VPWR.t1172 629.652
R1353 VPWR.n2567 VPWR.t1190 629.652
R1354 VPWR.n2578 VPWR.t1318 629.652
R1355 VPWR.n2579 VPWR.t1451 629.652
R1356 VPWR.n2590 VPWR.t1091 629.652
R1357 VPWR.n1594 VPWR.t1107 629.652
R1358 VPWR.t1243 VPWR.n1593 629.652
R1359 VPWR.n1182 VPWR.t1256 629.652
R1360 VPWR.n1185 VPWR.t1416 629.652
R1361 VPWR.n1220 VPWR.t1137 629.652
R1362 VPWR.t1284 VPWR.n1219 629.652
R1363 VPWR.t1392 VPWR.n1216 629.652
R1364 VPWR.t1432 VPWR.n1213 629.652
R1365 VPWR.t1177 VPWR.n1205 629.652
R1366 VPWR.t1281 VPWR.n1202 629.652
R1367 VPWR.t1440 VPWR.n1199 629.652
R1368 VPWR.t1459 VPWR.n1191 629.652
R1369 VPWR.t1203 VPWR.n1188 629.652
R1370 VPWR.n1740 VPWR.t1332 629.652
R1371 VPWR.t1360 VPWR.n1739 629.652
R1372 VPWR.n2836 VPWR.t556 531.804
R1373 VPWR.n2855 VPWR.t556 531.804
R1374 VPWR.n2851 VPWR.n2850 504.707
R1375 VPWR.t821 VPWR.t402 486.048
R1376 VPWR.t1836 VPWR.t1651 486.048
R1377 VPWR.t1647 VPWR.t1499 486.048
R1378 VPWR.t127 VPWR.t1646 486.048
R1379 VPWR.t401 VPWR.t853 486.048
R1380 VPWR.t948 VPWR.t1866 486.048
R1381 VPWR.t1865 VPWR.t304 486.048
R1382 VPWR.t213 VPWR.t400 486.048
R1383 VPWR.t103 VPWR.t411 486.048
R1384 VPWR.t72 VPWR.t1867 486.048
R1385 VPWR.t1645 VPWR.t647 486.048
R1386 VPWR.t209 VPWR.t1644 486.048
R1387 VPWR.t1864 VPWR.t263 486.048
R1388 VPWR.t586 VPWR.t1863 486.048
R1389 VPWR.t1862 VPWR.t20 486.048
R1390 VPWR.t1225 VPWR.t1652 486.048
R1391 VPWR.t1745 VPWR.t1643 486.048
R1392 VPWR.t75 VPWR.t1671 486.048
R1393 VPWR.t738 VPWR.t1471 486.048
R1394 VPWR.t737 VPWR.t1830 486.048
R1395 VPWR.t1642 VPWR.t976 486.048
R1396 VPWR.t938 VPWR.t787 486.048
R1397 VPWR.t937 VPWR.t265 486.048
R1398 VPWR.t1641 VPWR.t1697 486.048
R1399 VPWR.t1640 VPWR.t453 486.048
R1400 VPWR.t74 VPWR.t338 486.048
R1401 VPWR.t736 VPWR.t1001 486.048
R1402 VPWR.t735 VPWR.t893 486.048
R1403 VPWR.t936 VPWR.t871 486.048
R1404 VPWR.t935 VPWR.t1042 486.048
R1405 VPWR.t739 VPWR.t173 486.048
R1406 VPWR.t76 VPWR.t1443 486.048
R1407 VPWR.t631 VPWR.t1887 486.048
R1408 VPWR.t1882 VPWR.t1586 486.048
R1409 VPWR.t1511 VPWR.t1655 486.048
R1410 VPWR.t1654 VPWR.t1811 486.048
R1411 VPWR.t742 VPWR.t1886 486.048
R1412 VPWR.t1660 VPWR.t1761 486.048
R1413 VPWR.t12 VPWR.t1659 486.048
R1414 VPWR.t1885 VPWR.t161 486.048
R1415 VPWR.t181 VPWR.t1884 486.048
R1416 VPWR.t1661 VPWR.t60 486.048
R1417 VPWR.t592 VPWR.t1923 486.048
R1418 VPWR.t1922 VPWR.t1003 486.048
R1419 VPWR.t251 VPWR.t1658 486.048
R1420 VPWR.t1657 VPWR.t1054 486.048
R1421 VPWR.t1711 VPWR.t1656 486.048
R1422 VPWR.t1883 VPWR.t1292 486.048
R1423 VPWR.t1751 VPWR.t367 486.048
R1424 VPWR.t681 VPWR.t362 486.048
R1425 VPWR.t1463 VPWR.t351 486.048
R1426 VPWR.t322 VPWR.t350 486.048
R1427 VPWR.t754 VPWR.t366 486.048
R1428 VPWR.t807 VPWR.t847 486.048
R1429 VPWR.t277 VPWR.t846 486.048
R1430 VPWR.t1709 VPWR.t365 486.048
R1431 VPWR.t665 VPWR.t364 486.048
R1432 VPWR.t535 VPWR.t848 486.048
R1433 VPWR.t1632 VPWR.t349 486.048
R1434 VPWR.t991 VPWR.t348 486.048
R1435 VPWR.t90 VPWR.t845 486.048
R1436 VPWR.t1048 VPWR.t844 486.048
R1437 VPWR.t227 VPWR.t843 486.048
R1438 VPWR.t1400 VPWR.t363 486.048
R1439 VPWR.t692 VPWR.t446 486.048
R1440 VPWR.t728 VPWR.t841 486.048
R1441 VPWR.t1648 VPWR.t1483 486.048
R1442 VPWR.t1727 VPWR.t1593 486.048
R1443 VPWR.t445 VPWR.t77 486.048
R1444 VPWR.t799 VPWR.t116 486.048
R1445 VPWR.t115 VPWR.t189 486.048
R1446 VPWR.t459 VPWR.t444 486.048
R1447 VPWR.t443 VPWR.t1821 486.048
R1448 VPWR.t1537 VPWR.t117 486.048
R1449 VPWR.t1592 VPWR.t831 486.048
R1450 VPWR.t1735 VPWR.t1591 486.048
R1451 VPWR.t114 VPWR.t1799 486.048
R1452 VPWR.t1543 VPWR.t1650 486.048
R1453 VPWR.t1649 VPWR.t165 486.048
R1454 VPWR.t1126 VPWR.t842 486.048
R1455 VPWR.t1846 VPWR.t774 486.048
R1456 VPWR.t940 VPWR.t1834 486.048
R1457 VPWR.t656 VPWR.t1501 486.048
R1458 VPWR.t655 VPWR.t1574 486.048
R1459 VPWR.t773 VPWR.t851 486.048
R1460 VPWR.t87 VPWR.t946 486.048
R1461 VPWR.t86 VPWR.t302 486.048
R1462 VPWR.t772 VPWR.t211 486.048
R1463 VPWR.t1603 VPWR.t409 486.048
R1464 VPWR.t939 VPWR.t68 486.048
R1465 VPWR.t654 VPWR.t645 486.048
R1466 VPWR.t653 VPWR.t205 486.048
R1467 VPWR.t85 VPWR.t261 486.048
R1468 VPWR.t84 VPWR.t582 486.048
R1469 VPWR.t83 VPWR.t1719 486.048
R1470 VPWR.t1602 VPWR.t1233 486.048
R1471 VPWR.t823 VPWR.t1036 486.048
R1472 VPWR.t1041 VPWR.t1840 486.048
R1473 VPWR.t1491 VPWR.t985 486.048
R1474 VPWR.t984 VPWR.t129 486.048
R1475 VPWR.t1073 VPWR.t1035 486.048
R1476 VPWR.t1039 VPWR.t1675 486.048
R1477 VPWR.t308 VPWR.t1038 486.048
R1478 VPWR.t1034 VPWR.t147 486.048
R1479 VPWR.t865 VPWR.t1033 486.048
R1480 VPWR.t1040 VPWR.t1529 486.048
R1481 VPWR.t1916 VPWR.t983 486.048
R1482 VPWR.t982 VPWR.t1594 486.048
R1483 VPWR.t1789 VPWR.t1037 486.048
R1484 VPWR.t987 VPWR.t588 486.048
R1485 VPWR.t22 VPWR.t986 486.048
R1486 VPWR.t1032 VPWR.t1193 486.048
R1487 VPWR.t629 VPWR.t1897 486.048
R1488 VPWR.t1582 VPWR.t1895 486.048
R1489 VPWR.t1495 VPWR.t119 486.048
R1490 VPWR.t1809 VPWR.t120 486.048
R1491 VPWR.t1878 VPWR.t610 486.048
R1492 VPWR.t1757 VPWR.t123 486.048
R1493 VPWR.t8 VPWR.t124 486.048
R1494 VPWR.t159 VPWR.t1896 486.048
R1495 VPWR.t177 VPWR.t126 486.048
R1496 VPWR.t58 VPWR.t122 486.048
R1497 VPWR.t396 VPWR.t113 486.048
R1498 VPWR.t675 VPWR.t112 486.048
R1499 VPWR.t249 VPWR.t125 486.048
R1500 VPWR.t1052 VPWR.t121 486.048
R1501 VPWR.t1064 VPWR.t118 486.048
R1502 VPWR.t1298 VPWR.t1894 486.048
R1503 VPWR.t917 VPWR.t1907 486.048
R1504 VPWR.t779 VPWR.t899 486.048
R1505 VPWR.t1911 VPWR.t1481 486.048
R1506 VPWR.t1731 VPWR.t1910 486.048
R1507 VPWR.t1906 VPWR.t79 486.048
R1508 VPWR.t801 VPWR.t1570 486.048
R1509 VPWR.t1569 VPWR.t191 486.048
R1510 VPWR.t461 VPWR.t902 486.048
R1511 VPWR.t901 VPWR.t1823 486.048
R1512 VPWR.t1539 VPWR.t1571 486.048
R1513 VPWR.t1909 VPWR.t833 486.048
R1514 VPWR.t1737 VPWR.t1908 486.048
R1515 VPWR.t1568 VPWR.t1801 486.048
R1516 VPWR.t1545 VPWR.t1567 486.048
R1517 VPWR.t1566 VPWR.t169 486.048
R1518 VPWR.t1121 VPWR.t900 486.048
R1519 VPWR.t627 VPWR.t956 486.048
R1520 VPWR.t1639 VPWR.t1580 486.048
R1521 VPWR.t928 VPWR.t1513 486.048
R1522 VPWR.t927 VPWR.t1807 486.048
R1523 VPWR.t955 VPWR.t1876 486.048
R1524 VPWR.t1637 VPWR.t1755 486.048
R1525 VPWR.t1636 VPWR.t6 486.048
R1526 VPWR.t954 VPWR.t157 486.048
R1527 VPWR.t953 VPWR.t141 486.048
R1528 VPWR.t1638 VPWR.t766 486.048
R1529 VPWR.t926 VPWR.t394 486.048
R1530 VPWR.t925 VPWR.t673 486.048
R1531 VPWR.t1635 VPWR.t247 486.048
R1532 VPWR.t1634 VPWR.t1050 486.048
R1533 VPWR.t929 VPWR.t1062 486.048
R1534 VPWR.t952 VPWR.t1305 486.048
R1535 VPWR.t919 VPWR.t606 486.048
R1536 VPWR.t781 VPWR.t941 486.048
R1537 VPWR.t1479 VPWR.t686 486.048
R1538 VPWR.t1733 VPWR.t685 486.048
R1539 VPWR.t81 VPWR.t605 486.048
R1540 VPWR.t803 VPWR.t972 486.048
R1541 VPWR.t193 VPWR.t971 486.048
R1542 VPWR.t463 VPWR.t604 486.048
R1543 VPWR.t1825 VPWR.t603 486.048
R1544 VPWR.t1541 VPWR.t973 486.048
R1545 VPWR.t835 VPWR.t684 486.048
R1546 VPWR.t1739 VPWR.t683 486.048
R1547 VPWR.t1803 VPWR.t970 486.048
R1548 VPWR.t1547 VPWR.t969 486.048
R1549 VPWR.t171 VPWR.t687 486.048
R1550 VPWR.t1113 VPWR.t602 486.048
R1551 VPWR.t1749 VPWR.t908 486.048
R1552 VPWR.t903 VPWR.t705 486.048
R1553 VPWR.t1465 VPWR.t1031 486.048
R1554 VPWR.t1030 VPWR.t318 486.048
R1555 VPWR.t752 VPWR.t907 486.048
R1556 VPWR.t861 VPWR.t805 486.048
R1557 VPWR.t275 VPWR.t860 486.048
R1558 VPWR.t906 VPWR.t1705 486.048
R1559 VPWR.t663 VPWR.t905 486.048
R1560 VPWR.t862 VPWR.t533 486.048
R1561 VPWR.t1630 VPWR.t1029 486.048
R1562 VPWR.t1028 VPWR.t897 486.048
R1563 VPWR.t879 VPWR.t859 486.048
R1564 VPWR.t858 VPWR.t1046 486.048
R1565 VPWR.t223 VPWR.t857 486.048
R1566 VPWR.t904 VPWR.t1413 486.048
R1567 VPWR.t1562 VPWR.t931 486.048
R1568 VPWR.t344 VPWR.t707 486.048
R1569 VPWR.t1461 VPWR.t1673 486.048
R1570 VPWR.t934 VPWR.t324 486.048
R1571 VPWR.t756 VPWR.t930 486.048
R1572 VPWR.t817 VPWR.t809 486.048
R1573 VPWR.t279 VPWR.t816 486.048
R1574 VPWR.t347 VPWR.t199 486.048
R1575 VPWR.t667 VPWR.t346 486.048
R1576 VPWR.t818 VPWR.t537 486.048
R1577 VPWR.t768 VPWR.t933 486.048
R1578 VPWR.t932 VPWR.t993 486.048
R1579 VPWR.t92 VPWR.t815 486.048
R1580 VPWR.t814 VPWR.t1021 486.048
R1581 VPWR.t229 VPWR.t1674 486.048
R1582 VPWR.t345 VPWR.t1395 486.048
R1583 VPWR.t1844 VPWR.t1025 486.048
R1584 VPWR.t909 VPWR.t1588 486.048
R1585 VPWR.t1503 VPWR.t1664 486.048
R1586 VPWR.t1813 VPWR.t1663 486.048
R1587 VPWR.t744 VPWR.t601 486.048
R1588 VPWR.t1763 VPWR.t424 486.048
R1589 VPWR.t14 VPWR.t423 486.048
R1590 VPWR.t163 VPWR.t600 486.048
R1591 VPWR.t183 VPWR.t1590 486.048
R1592 VPWR.t66 VPWR.t425 486.048
R1593 VPWR.t594 VPWR.t1027 486.048
R1594 VPWR.t1009 VPWR.t1026 486.048
R1595 VPWR.t253 VPWR.t422 486.048
R1596 VPWR.t1551 VPWR.t1666 486.048
R1597 VPWR.t1713 VPWR.t1665 486.048
R1598 VPWR.t1265 VPWR.t1589 486.048
R1599 VPWR.t1747 VPWR.t1774 486.048
R1600 VPWR.t241 VPWR.t699 486.048
R1601 VPWR.t1604 VPWR.t1469 486.048
R1602 VPWR.t1777 VPWR.t312 486.048
R1603 VPWR.t1773 VPWR.t980 486.048
R1604 VPWR.t239 VPWR.t791 486.048
R1605 VPWR.t883 VPWR.t269 486.048
R1606 VPWR.t244 VPWR.t1701 486.048
R1607 VPWR.t243 VPWR.t657 486.048
R1608 VPWR.t240 VPWR.t340 486.048
R1609 VPWR.t1776 VPWR.t1624 486.048
R1610 VPWR.t1775 VPWR.t895 486.048
R1611 VPWR.t882 VPWR.t875 486.048
R1612 VPWR.t881 VPWR.t1044 486.048
R1613 VPWR.t1605 VPWR.t175 486.048
R1614 VPWR.t242 VPWR.t1435 486.048
R1615 VPWR.t1564 VPWR.t1170 486.048
R1616 VPWR.t709 VPWR.t1301 486.048
R1617 VPWR.t1517 VPWR.t1430 486.048
R1618 VPWR.t149 VPWR.t1089 486.048
R1619 VPWR.t1880 VPWR.t1196 486.048
R1620 VPWR.t1351 VPWR.t811 486.048
R1621 VPWR.t281 VPWR.t1353 486.048
R1622 VPWR.t1201 VPWR.t201 486.048
R1623 VPWR.t1068 VPWR.t1231 486.048
R1624 VPWR.t1349 VPWR.t539 486.048
R1625 VPWR.t1100 VPWR.t770 486.048
R1626 VPWR.t1119 VPWR.t995 486.048
R1627 VPWR.t1363 VPWR.t94 486.048
R1628 VPWR.t1023 VPWR.t1381 486.048
R1629 VPWR.t1419 VPWR.t233 486.048
R1630 VPWR.t1376 VPWR.t1251 486.048
R1631 VPWR.t1236 VPWR.t1105 486.048
R1632 VPWR.t1365 VPWR.t1241 486.048
R1633 VPWR.t1371 VPWR.t1383 486.048
R1634 VPWR.t1145 VPWR.t1411 486.048
R1635 VPWR.t1135 VPWR.t1253 486.048
R1636 VPWR.t1408 VPWR.t1279 486.048
R1637 VPWR.t1303 VPWR.t1132 486.048
R1638 VPWR.t1167 VPWR.t1140 486.048
R1639 VPWR.t1175 VPWR.t1295 486.048
R1640 VPWR.t1405 VPWR.t1277 486.048
R1641 VPWR.t1438 VPWR.t1172 486.048
R1642 VPWR.t1190 VPWR.t1457 486.048
R1643 VPWR.t1311 VPWR.t1318 486.048
R1644 VPWR.t1451 VPWR.t1330 486.048
R1645 VPWR.t1355 VPWR.t1091 486.048
R1646 VPWR.t1327 VPWR.t1206 486.048
R1647 VPWR.t1107 VPWR.t1379 486.048
R1648 VPWR.t1124 VPWR.t1243 486.048
R1649 VPWR.t1256 VPWR.t1249 486.048
R1650 VPWR.t1416 VPWR.t1290 486.048
R1651 VPWR.t1137 VPWR.t1398 486.048
R1652 VPWR.t1165 VPWR.t1284 486.048
R1653 VPWR.t1180 VPWR.t1392 486.048
R1654 VPWR.t1403 VPWR.t1432 486.048
R1655 VPWR.t1446 VPWR.t1177 486.048
R1656 VPWR.t1163 VPWR.t1281 486.048
R1657 VPWR.t1316 VPWR.t1440 486.048
R1658 VPWR.t1338 VPWR.t1459 486.048
R1659 VPWR.t1188 VPWR.t1203 486.048
R1660 VPWR.t1214 VPWR.t1332 486.048
R1661 VPWR.t1239 VPWR.t1360 486.048
R1662 VPWR.t1211 VPWR.t1087 486.048
R1663 VPWR.t402 VPWR.t552 463.954
R1664 VPWR.t1651 VPWR.t1842 463.954
R1665 VPWR.t913 VPWR.t1647 463.954
R1666 VPWR.t1646 VPWR.t1519 463.954
R1667 VPWR.t153 VPWR.t401 463.954
R1668 VPWR.t1866 VPWR.t849 463.954
R1669 VPWR.t944 VPWR.t1865 463.954
R1670 VPWR.t400 VPWR.t300 463.954
R1671 VPWR.t457 VPWR.t103 463.954
R1672 VPWR.t1867 VPWR.t407 463.954
R1673 VPWR.t64 VPWR.t1645 463.954
R1674 VPWR.t1644 VPWR.t643 463.954
R1675 VPWR.t1007 VPWR.t1864 463.954
R1676 VPWR.t1863 VPWR.t98 463.954
R1677 VPWR.t1549 VPWR.t1862 463.954
R1678 VPWR.t1652 VPWR.t1058 463.954
R1679 VPWR.t1643 VPWR.t564 463.954
R1680 VPWR.t921 VPWR.t75 463.954
R1681 VPWR.t1667 VPWR.t738 463.954
R1682 VPWR.t1497 VPWR.t737 463.954
R1683 VPWR.t131 VPWR.t1642 463.954
R1684 VPWR.t403 VPWR.t938 463.954
R1685 VPWR.t783 VPWR.t937 463.954
R1686 VPWR.t195 VPWR.t1641 463.954
R1687 VPWR.t145 VPWR.t1640 463.954
R1688 VPWR.t449 VPWR.t74 463.954
R1689 VPWR.t328 VPWR.t736 463.954
R1690 VPWR.t997 VPWR.t735 463.954
R1691 VPWR.t215 VPWR.t936 463.954
R1692 VPWR.t1787 VPWR.t935 463.954
R1693 VPWR.t352 VPWR.t739 463.954
R1694 VPWR.t24 VPWR.t76 463.954
R1695 VPWR.t1887 VPWR.t578 463.954
R1696 VPWR.t1557 VPWR.t1882 463.954
R1697 VPWR.t1655 VPWR.t1578 463.954
R1698 VPWR.t1473 VPWR.t1654 463.954
R1699 VPWR.t1886 VPWR.t320 463.954
R1700 VPWR.t1874 VPWR.t1660 463.954
R1701 VPWR.t1659 VPWR.t1753 463.954
R1702 VPWR.t4 VPWR.t1885 463.954
R1703 VPWR.t1884 VPWR.t1703 463.954
R1704 VPWR.t139 VPWR.t1661 463.954
R1705 VPWR.t1923 VPWR.t762 463.954
R1706 VPWR.t392 VPWR.t1922 463.954
R1707 VPWR.t1658 VPWR.t669 463.954
R1708 VPWR.t877 VPWR.t1657 463.954
R1709 VPWR.t1656 VPWR.t598 463.954
R1710 VPWR.t225 VPWR.t1883 463.954
R1711 VPWR.t367 VPWR.t570 463.954
R1712 VPWR.t362 VPWR.t1741 463.954
R1713 VPWR.t351 VPWR.t701 463.954
R1714 VPWR.t350 VPWR.t1487 463.954
R1715 VPWR.t366 VPWR.t1725 463.954
R1716 VPWR.t847 VPWR.t748 463.954
R1717 VPWR.t846 VPWR.t793 463.954
R1718 VPWR.t365 VPWR.t271 463.954
R1719 VPWR.t364 VPWR.t1854 463.954
R1720 VPWR.t848 VPWR.t659 463.954
R1721 VPWR.t349 VPWR.t334 463.954
R1722 VPWR.t348 VPWR.t1626 463.954
R1723 VPWR.t845 VPWR.t889 463.954
R1724 VPWR.t844 VPWR.t1795 463.954
R1725 VPWR.t843 VPWR.t637 463.954
R1726 VPWR.t363 VPWR.t30 463.954
R1727 VPWR.t446 VPWR.t558 463.954
R1728 VPWR.t841 VPWR.t284 463.954
R1729 VPWR.t722 VPWR.t1648 463.954
R1730 VPWR.t1593 VPWR.t1509 463.954
R1731 VPWR.t1815 VPWR.t445 463.954
R1732 VPWR.t116 VPWR.t1075 463.954
R1733 VPWR.t1677 VPWR.t115 463.954
R1734 VPWR.t444 VPWR.t310 463.954
R1735 VPWR.t416 VPWR.t443 463.954
R1736 VPWR.t117 VPWR.t867 463.954
R1737 VPWR.t1531 VPWR.t1592 463.954
R1738 VPWR.t1591 VPWR.t825 463.954
R1739 VPWR.t1596 VPWR.t114 463.954
R1740 VPWR.t1650 VPWR.t255 463.954
R1741 VPWR.t356 VPWR.t1649 463.954
R1742 VPWR.t842 VPWR.t1715 463.954
R1743 VPWR.t774 VPWR.t550 463.954
R1744 VPWR.t633 VPWR.t940 463.954
R1745 VPWR.t911 VPWR.t656 463.954
R1746 VPWR.t1521 VPWR.t655 463.954
R1747 VPWR.t151 VPWR.t773 463.954
R1748 VPWR.t746 VPWR.t87 463.954
R1749 VPWR.t942 VPWR.t86 463.954
R1750 VPWR.t298 VPWR.t772 463.954
R1751 VPWR.t203 VPWR.t1603 463.954
R1752 VPWR.t405 VPWR.t939 463.954
R1753 VPWR.t62 VPWR.t654 463.954
R1754 VPWR.t596 VPWR.t653 463.954
R1755 VPWR.t1005 VPWR.t85 463.954
R1756 VPWR.t96 VPWR.t84 463.954
R1757 VPWR.t1056 VPWR.t83 463.954
R1758 VPWR.t235 VPWR.t1602 463.954
R1759 VPWR.t1036 VPWR.t554 463.954
R1760 VPWR.t819 VPWR.t1041 463.954
R1761 VPWR.t985 VPWR.t1838 463.954
R1762 VPWR.t1515 VPWR.t984 463.954
R1763 VPWR.t1035 VPWR.t1805 463.954
R1764 VPWR.t855 VPWR.t1039 463.954
R1765 VPWR.t1038 VPWR.t950 463.954
R1766 VPWR.t306 VPWR.t1034 463.954
R1767 VPWR.t1033 VPWR.t155 463.954
R1768 VPWR.t863 VPWR.t1040 463.954
R1769 VPWR.t983 VPWR.t70 463.954
R1770 VPWR.t1914 VPWR.t982 463.954
R1771 VPWR.t1037 VPWR.t207 463.954
R1772 VPWR.t245 VPWR.t987 463.954
R1773 VPWR.t986 VPWR.t584 463.954
R1774 VPWR.t1060 VPWR.t1032 463.954
R1775 VPWR.t1897 VPWR.t576 463.954
R1776 VPWR.t1895 VPWR.t1555 463.954
R1777 VPWR.t119 VPWR.t679 463.954
R1778 VPWR.t120 VPWR.t1475 463.954
R1779 VPWR.t610 VPWR.t316 463.954
R1780 VPWR.t123 VPWR.t1872 463.954
R1781 VPWR.t124 VPWR.t959 463.954
R1782 VPWR.t1896 VPWR.t2 463.954
R1783 VPWR.t126 VPWR.t1699 463.954
R1784 VPWR.t122 VPWR.t137 463.954
R1785 VPWR.t113 VPWR.t760 463.954
R1786 VPWR.t112 VPWR.t390 463.954
R1787 VPWR.t125 VPWR.t777 463.954
R1788 VPWR.t121 VPWR.t873 463.954
R1789 VPWR.t118 VPWR.t386 463.954
R1790 VPWR.t1894 VPWR.t221 463.954
R1791 VPWR.t1907 VPWR.t560 463.954
R1792 VPWR.t899 VPWR.t286 463.954
R1793 VPWR.t724 VPWR.t1911 463.954
R1794 VPWR.t1910 VPWR.t1507 463.954
R1795 VPWR.t1572 VPWR.t1906 463.954
R1796 VPWR.t1570 VPWR.t294 463.954
R1797 VPWR.t1679 VPWR.t1569 463.954
R1798 VPWR.t902 VPWR.t185 463.954
R1799 VPWR.t418 VPWR.t901 463.954
R1800 VPWR.t1571 VPWR.t1817 463.954
R1801 VPWR.t1533 VPWR.t1909 463.954
R1802 VPWR.t1908 VPWR.t827 463.954
R1803 VPWR.t1598 VPWR.t1568 463.954
R1804 VPWR.t1567 VPWR.t257 463.954
R1805 VPWR.t358 VPWR.t1566 463.954
R1806 VPWR.t900 VPWR.t1717 463.954
R1807 VPWR.t956 VPWR.t574 463.954
R1808 VPWR.t1553 VPWR.t1639 463.954
R1809 VPWR.t677 VPWR.t928 463.954
R1810 VPWR.t1477 VPWR.t927 463.954
R1811 VPWR.t314 VPWR.t955 463.954
R1812 VPWR.t1870 VPWR.t1637 463.954
R1813 VPWR.t957 VPWR.t1636 463.954
R1814 VPWR.t0 VPWR.t954 463.954
R1815 VPWR.t1858 VPWR.t953 463.954
R1816 VPWR.t135 VPWR.t1638 463.954
R1817 VPWR.t758 VPWR.t926 463.954
R1818 VPWR.t388 VPWR.t925 463.954
R1819 VPWR.t775 VPWR.t1635 463.954
R1820 VPWR.t869 VPWR.t1634 463.954
R1821 VPWR.t384 VPWR.t929 463.954
R1822 VPWR.t219 VPWR.t952 463.954
R1823 VPWR.t606 VPWR.t562 463.954
R1824 VPWR.t941 VPWR.t288 463.954
R1825 VPWR.t686 VPWR.t726 463.954
R1826 VPWR.t685 VPWR.t1505 463.954
R1827 VPWR.t605 VPWR.t1576 463.954
R1828 VPWR.t972 VPWR.t296 463.954
R1829 VPWR.t971 VPWR.t797 463.954
R1830 VPWR.t604 VPWR.t187 463.954
R1831 VPWR.t603 VPWR.t420 463.954
R1832 VPWR.t973 VPWR.t1819 463.954
R1833 VPWR.t684 VPWR.t1535 463.954
R1834 VPWR.t683 VPWR.t829 463.954
R1835 VPWR.t970 VPWR.t1600 463.954
R1836 VPWR.t969 VPWR.t259 463.954
R1837 VPWR.t687 VPWR.t360 463.954
R1838 VPWR.t602 VPWR.t18 463.954
R1839 VPWR.t908 VPWR.t568 463.954
R1840 VPWR.t435 VPWR.t903 463.954
R1841 VPWR.t1031 VPWR.t697 463.954
R1842 VPWR.t1489 VPWR.t1030 463.954
R1843 VPWR.t907 VPWR.t1723 463.954
R1844 VPWR.t978 VPWR.t861 463.954
R1845 VPWR.t860 VPWR.t789 463.954
R1846 VPWR.t267 VPWR.t906 463.954
R1847 VPWR.t905 VPWR.t1852 463.954
R1848 VPWR.t455 VPWR.t862 463.954
R1849 VPWR.t1029 VPWR.t332 463.954
R1850 VPWR.t1622 VPWR.t1028 463.954
R1851 VPWR.t859 VPWR.t887 463.954
R1852 VPWR.t1793 VPWR.t858 463.954
R1853 VPWR.t857 VPWR.t635 463.954
R1854 VPWR.t28 VPWR.t904 463.954
R1855 VPWR.t931 VPWR.t572 463.954
R1856 VPWR.t1743 VPWR.t344 463.954
R1857 VPWR.t1673 VPWR.t703 463.954
R1858 VPWR.t1485 VPWR.t934 463.954
R1859 VPWR.t930 VPWR.t1729 463.954
R1860 VPWR.t750 VPWR.t817 463.954
R1861 VPWR.t816 VPWR.t795 463.954
R1862 VPWR.t273 VPWR.t347 463.954
R1863 VPWR.t346 VPWR.t1856 463.954
R1864 VPWR.t661 VPWR.t818 463.954
R1865 VPWR.t933 VPWR.t336 463.954
R1866 VPWR.t1628 VPWR.t932 463.954
R1867 VPWR.t815 VPWR.t891 463.954
R1868 VPWR.t1797 VPWR.t814 463.954
R1869 VPWR.t1674 VPWR.t639 463.954
R1870 VPWR.t167 VPWR.t345 463.954
R1871 VPWR.t1025 VPWR.t580 463.954
R1872 VPWR.t1588 VPWR.t625 463.954
R1873 VPWR.t1664 VPWR.t1584 463.954
R1874 VPWR.t1663 VPWR.t1467 463.954
R1875 VPWR.t601 VPWR.t326 463.954
R1876 VPWR.t424 VPWR.t740 463.954
R1877 VPWR.t423 VPWR.t1759 463.954
R1878 VPWR.t600 VPWR.t10 463.954
R1879 VPWR.t1590 VPWR.t1707 463.954
R1880 VPWR.t425 VPWR.t179 463.954
R1881 VPWR.t1027 VPWR.t764 463.954
R1882 VPWR.t1026 VPWR.t590 463.954
R1883 VPWR.t422 VPWR.t671 463.954
R1884 VPWR.t1666 VPWR.t88 463.954
R1885 VPWR.t1665 VPWR.t641 463.954
R1886 VPWR.t1589 VPWR.t231 463.954
R1887 VPWR.t1774 VPWR.t566 463.954
R1888 VPWR.t923 VPWR.t241 463.954
R1889 VPWR.t1669 VPWR.t1604 463.954
R1890 VPWR.t1493 VPWR.t1777 463.954
R1891 VPWR.t1721 VPWR.t1773 463.954
R1892 VPWR.t974 VPWR.t239 463.954
R1893 VPWR.t785 VPWR.t883 463.954
R1894 VPWR.t197 VPWR.t244 463.954
R1895 VPWR.t1850 VPWR.t243 463.954
R1896 VPWR.t451 VPWR.t240 463.954
R1897 VPWR.t330 VPWR.t1776 463.954
R1898 VPWR.t999 VPWR.t1775 463.954
R1899 VPWR.t217 VPWR.t882 463.954
R1900 VPWR.t1791 VPWR.t881 463.954
R1901 VPWR.t354 VPWR.t1605 463.954
R1902 VPWR.t26 VPWR.t242 463.954
R1903 VPWR.t1170 VPWR.t1185 463.954
R1904 VPWR.t1301 VPWR.t1346 463.954
R1905 VPWR.t1430 VPWR.t1448 463.954
R1906 VPWR.t1089 VPWR.t1219 463.954
R1907 VPWR.t1196 VPWR.t1321 463.954
R1908 VPWR.t1343 VPWR.t1351 463.954
R1909 VPWR.t1353 VPWR.t1094 463.954
R1910 VPWR.t1216 VPWR.t1201 463.954
R1911 VPWR.t1231 VPWR.t1357 463.954
R1912 VPWR.t1373 VPWR.t1349 463.954
R1913 VPWR.t1116 VPWR.t1100 463.954
R1914 VPWR.t1246 VPWR.t1119 463.954
R1915 VPWR.t1287 VPWR.t1363 463.954
R1916 VPWR.t1381 VPWR.t1110 463.954
R1917 VPWR.t1160 VPWR.t1419 463.954
R1918 VPWR.t1251 VPWR.t1268 463.954
R1919 VPWR.t1105 VPWR.t1129 463.954
R1920 VPWR.t1241 VPWR.t1274 463.954
R1921 VPWR.t1386 VPWR.t1371 463.954
R1922 VPWR.t1411 VPWR.t1151 463.954
R1923 VPWR.t1259 VPWR.t1135 463.954
R1924 VPWR.t1279 VPWR.t1271 463.954
R1925 VPWR.t1427 VPWR.t1303 463.954
R1926 VPWR.t1140 VPWR.t1148 463.954
R1927 VPWR.t1308 VPWR.t1175 463.954
R1928 VPWR.t1277 VPWR.t1324 463.954
R1929 VPWR.t1454 VPWR.t1438 463.954
R1930 VPWR.t1457 VPWR.t1198 463.954
R1931 VPWR.t1228 VPWR.t1311 463.954
R1932 VPWR.t1330 VPWR.t1078 463.954
R1933 VPWR.t1097 VPWR.t1355 463.954
R1934 VPWR.t1206 VPWR.t1222 463.954
R1935 VPWR.t1379 VPWR.t1389 463.954
R1936 VPWR.t1157 VPWR.t1124 463.954
R1937 VPWR.t1249 VPWR.t1262 463.954
R1938 VPWR.t1290 VPWR.t1424 463.954
R1939 VPWR.t1398 VPWR.t1142 463.954
R1940 VPWR.t1154 VPWR.t1165 463.954
R1941 VPWR.t1313 VPWR.t1180 463.954
R1942 VPWR.t1421 VPWR.t1403 463.954
R1943 VPWR.t1182 VPWR.t1446 463.954
R1944 VPWR.t1208 VPWR.t1163 463.954
R1945 VPWR.t1335 VPWR.t1316 463.954
R1946 VPWR.t1081 VPWR.t1338 463.954
R1947 VPWR.t1102 VPWR.t1188 463.954
R1948 VPWR.t1340 VPWR.t1214 463.954
R1949 VPWR.t1368 VPWR.t1239 463.954
R1950 VPWR.t1087 VPWR.t1084 463.954
R1951 VPWR.n2626 VPWR.t1610 428.822
R1952 VPWR.n1595 VPWR.n1594 376.045
R1953 VPWR.n2506 VPWR.n2505 376.045
R1954 VPWR.n1468 VPWR.n1467 376.045
R1955 VPWR.n351 VPWR.n350 376.045
R1956 VPWR.n2568 VPWR.n2567 376.045
R1957 VPWR.n1535 VPWR.n1534 376.045
R1958 VPWR.n349 VPWR.n348 376.045
R1959 VPWR.n2508 VPWR.n2507 376.045
R1960 VPWR.n966 VPWR.n965 376.045
R1961 VPWR.n2478 VPWR.n2477 376.045
R1962 VPWR.n2476 VPWR.n2475 376.045
R1963 VPWR.n321 VPWR.n320 376.045
R1964 VPWR.n2554 VPWR.n2553 376.045
R1965 VPWR.n974 VPWR.n973 376.045
R1966 VPWR.n2446 VPWR.n2445 376.045
R1967 VPWR.n325 VPWR.n324 376.045
R1968 VPWR.n2544 VPWR.n2543 376.045
R1969 VPWR.n1890 VPWR.n1889 376.045
R1970 VPWR.n1888 VPWR.n1887 376.045
R1971 VPWR.n1880 VPWR.n1879 376.045
R1972 VPWR.n390 VPWR.n389 376.045
R1973 VPWR.n394 VPWR.n393 376.045
R1974 VPWR.n398 VPWR.n397 376.045
R1975 VPWR.n2456 VPWR.n2455 376.045
R1976 VPWR.n333 VPWR.n332 376.045
R1977 VPWR.n2532 VPWR.n2531 376.045
R1978 VPWR.n1878 VPWR.n1877 376.045
R1979 VPWR.n406 VPWR.n405 376.045
R1980 VPWR.n2458 VPWR.n2457 376.045
R1981 VPWR.n337 VPWR.n336 376.045
R1982 VPWR.n2530 VPWR.n2529 376.045
R1983 VPWR.n2309 VPWR.n2308 376.045
R1984 VPWR.n2311 VPWR.n2310 376.045
R1985 VPWR.n2319 VPWR.n2318 376.045
R1986 VPWR.n2321 VPWR.n2320 376.045
R1987 VPWR.n2331 VPWR.n2330 376.045
R1988 VPWR.n2339 VPWR.n2338 376.045
R1989 VPWR.n2341 VPWR.n2340 376.045
R1990 VPWR.n2349 VPWR.n2348 376.045
R1991 VPWR.n2351 VPWR.n2350 376.045
R1992 VPWR.n2359 VPWR.n2358 376.045
R1993 VPWR.n2361 VPWR.n2360 376.045
R1994 VPWR.n2369 VPWR.n2368 376.045
R1995 VPWR.n2371 VPWR.n2370 376.045
R1996 VPWR.n2379 VPWR.n2378 376.045
R1997 VPWR.n2329 VPWR.n2328 376.045
R1998 VPWR.n543 VPWR.n542 376.045
R1999 VPWR.n541 VPWR.n540 376.045
R2000 VPWR.n537 VPWR.n536 376.045
R2001 VPWR.n533 VPWR.n532 376.045
R2002 VPWR.n525 VPWR.n524 376.045
R2003 VPWR.n521 VPWR.n520 376.045
R2004 VPWR.n517 VPWR.n516 376.045
R2005 VPWR.n513 VPWR.n512 376.045
R2006 VPWR.n509 VPWR.n508 376.045
R2007 VPWR.n505 VPWR.n504 376.045
R2008 VPWR.n501 VPWR.n500 376.045
R2009 VPWR.n497 VPWR.n496 376.045
R2010 VPWR.n493 VPWR.n492 376.045
R2011 VPWR.n489 VPWR.n488 376.045
R2012 VPWR.n529 VPWR.n528 376.045
R2013 VPWR.n2282 VPWR.n2281 376.045
R2014 VPWR.n2280 VPWR.n2279 376.045
R2015 VPWR.n2272 VPWR.n2271 376.045
R2016 VPWR.n2270 VPWR.n2269 376.045
R2017 VPWR.n2260 VPWR.n2259 376.045
R2018 VPWR.n2252 VPWR.n2251 376.045
R2019 VPWR.n2250 VPWR.n2249 376.045
R2020 VPWR.n2242 VPWR.n2241 376.045
R2021 VPWR.n2240 VPWR.n2239 376.045
R2022 VPWR.n2232 VPWR.n2231 376.045
R2023 VPWR.n2230 VPWR.n2229 376.045
R2024 VPWR.n2222 VPWR.n2221 376.045
R2025 VPWR.n2220 VPWR.n2219 376.045
R2026 VPWR.n2212 VPWR.n2211 376.045
R2027 VPWR.n2262 VPWR.n2261 376.045
R2028 VPWR.n582 VPWR.n581 376.045
R2029 VPWR.n586 VPWR.n585 376.045
R2030 VPWR.n590 VPWR.n589 376.045
R2031 VPWR.n594 VPWR.n593 376.045
R2032 VPWR.n602 VPWR.n601 376.045
R2033 VPWR.n606 VPWR.n605 376.045
R2034 VPWR.n610 VPWR.n609 376.045
R2035 VPWR.n614 VPWR.n613 376.045
R2036 VPWR.n618 VPWR.n617 376.045
R2037 VPWR.n622 VPWR.n621 376.045
R2038 VPWR.n626 VPWR.n625 376.045
R2039 VPWR.n630 VPWR.n629 376.045
R2040 VPWR.n634 VPWR.n633 376.045
R2041 VPWR.n638 VPWR.n637 376.045
R2042 VPWR.n598 VPWR.n597 376.045
R2043 VPWR.n2113 VPWR.n2112 376.045
R2044 VPWR.n2115 VPWR.n2114 376.045
R2045 VPWR.n2123 VPWR.n2122 376.045
R2046 VPWR.n2125 VPWR.n2124 376.045
R2047 VPWR.n2135 VPWR.n2134 376.045
R2048 VPWR.n2143 VPWR.n2142 376.045
R2049 VPWR.n2145 VPWR.n2144 376.045
R2050 VPWR.n2153 VPWR.n2152 376.045
R2051 VPWR.n2155 VPWR.n2154 376.045
R2052 VPWR.n2163 VPWR.n2162 376.045
R2053 VPWR.n2165 VPWR.n2164 376.045
R2054 VPWR.n2173 VPWR.n2172 376.045
R2055 VPWR.n2175 VPWR.n2174 376.045
R2056 VPWR.n2183 VPWR.n2182 376.045
R2057 VPWR.n2133 VPWR.n2132 376.045
R2058 VPWR.n735 VPWR.n734 376.045
R2059 VPWR.n733 VPWR.n732 376.045
R2060 VPWR.n729 VPWR.n728 376.045
R2061 VPWR.n725 VPWR.n724 376.045
R2062 VPWR.n717 VPWR.n716 376.045
R2063 VPWR.n713 VPWR.n712 376.045
R2064 VPWR.n709 VPWR.n708 376.045
R2065 VPWR.n705 VPWR.n704 376.045
R2066 VPWR.n701 VPWR.n700 376.045
R2067 VPWR.n697 VPWR.n696 376.045
R2068 VPWR.n693 VPWR.n692 376.045
R2069 VPWR.n689 VPWR.n688 376.045
R2070 VPWR.n685 VPWR.n684 376.045
R2071 VPWR.n681 VPWR.n680 376.045
R2072 VPWR.n721 VPWR.n720 376.045
R2073 VPWR.n2086 VPWR.n2085 376.045
R2074 VPWR.n2084 VPWR.n2083 376.045
R2075 VPWR.n2076 VPWR.n2075 376.045
R2076 VPWR.n2074 VPWR.n2073 376.045
R2077 VPWR.n2064 VPWR.n2063 376.045
R2078 VPWR.n2056 VPWR.n2055 376.045
R2079 VPWR.n2054 VPWR.n2053 376.045
R2080 VPWR.n2046 VPWR.n2045 376.045
R2081 VPWR.n2044 VPWR.n2043 376.045
R2082 VPWR.n2036 VPWR.n2035 376.045
R2083 VPWR.n2034 VPWR.n2033 376.045
R2084 VPWR.n2026 VPWR.n2025 376.045
R2085 VPWR.n2024 VPWR.n2023 376.045
R2086 VPWR.n2016 VPWR.n2015 376.045
R2087 VPWR.n2066 VPWR.n2065 376.045
R2088 VPWR.n774 VPWR.n773 376.045
R2089 VPWR.n778 VPWR.n777 376.045
R2090 VPWR.n782 VPWR.n781 376.045
R2091 VPWR.n786 VPWR.n785 376.045
R2092 VPWR.n794 VPWR.n793 376.045
R2093 VPWR.n798 VPWR.n797 376.045
R2094 VPWR.n802 VPWR.n801 376.045
R2095 VPWR.n806 VPWR.n805 376.045
R2096 VPWR.n810 VPWR.n809 376.045
R2097 VPWR.n814 VPWR.n813 376.045
R2098 VPWR.n818 VPWR.n817 376.045
R2099 VPWR.n822 VPWR.n821 376.045
R2100 VPWR.n826 VPWR.n825 376.045
R2101 VPWR.n830 VPWR.n829 376.045
R2102 VPWR.n790 VPWR.n789 376.045
R2103 VPWR.n1917 VPWR.n1916 376.045
R2104 VPWR.n1919 VPWR.n1918 376.045
R2105 VPWR.n1927 VPWR.n1926 376.045
R2106 VPWR.n1929 VPWR.n1928 376.045
R2107 VPWR.n1939 VPWR.n1938 376.045
R2108 VPWR.n1947 VPWR.n1946 376.045
R2109 VPWR.n1949 VPWR.n1948 376.045
R2110 VPWR.n1957 VPWR.n1956 376.045
R2111 VPWR.n1959 VPWR.n1958 376.045
R2112 VPWR.n1967 VPWR.n1966 376.045
R2113 VPWR.n1969 VPWR.n1968 376.045
R2114 VPWR.n1977 VPWR.n1976 376.045
R2115 VPWR.n1979 VPWR.n1978 376.045
R2116 VPWR.n1987 VPWR.n1986 376.045
R2117 VPWR.n1937 VPWR.n1936 376.045
R2118 VPWR.n927 VPWR.n926 376.045
R2119 VPWR.n925 VPWR.n924 376.045
R2120 VPWR.n921 VPWR.n920 376.045
R2121 VPWR.n917 VPWR.n916 376.045
R2122 VPWR.n909 VPWR.n908 376.045
R2123 VPWR.n905 VPWR.n904 376.045
R2124 VPWR.n901 VPWR.n900 376.045
R2125 VPWR.n897 VPWR.n896 376.045
R2126 VPWR.n893 VPWR.n892 376.045
R2127 VPWR.n889 VPWR.n888 376.045
R2128 VPWR.n885 VPWR.n884 376.045
R2129 VPWR.n881 VPWR.n880 376.045
R2130 VPWR.n877 VPWR.n876 376.045
R2131 VPWR.n873 VPWR.n872 376.045
R2132 VPWR.n913 VPWR.n912 376.045
R2133 VPWR.n1870 VPWR.n1869 376.045
R2134 VPWR.n982 VPWR.n981 376.045
R2135 VPWR.n1494 VPWR.n1493 376.045
R2136 VPWR.n1221 VPWR.n1220 376.045
R2137 VPWR.n402 VPWR.n401 376.045
R2138 VPWR.n2466 VPWR.n2465 376.045
R2139 VPWR.n341 VPWR.n340 376.045
R2140 VPWR.n2520 VPWR.n2519 376.045
R2141 VPWR.n978 VPWR.n977 376.045
R2142 VPWR.n1492 VPWR.n1491 376.045
R2143 VPWR.n1185 VPWR.n1184 376.045
R2144 VPWR.n1868 VPWR.n1867 376.045
R2145 VPWR.n986 VPWR.n985 376.045
R2146 VPWR.n1506 VPWR.n1505 376.045
R2147 VPWR.n1219 VPWR.n1218 376.045
R2148 VPWR.n410 VPWR.n409 376.045
R2149 VPWR.n418 VPWR.n417 376.045
R2150 VPWR.n422 VPWR.n421 376.045
R2151 VPWR.n426 VPWR.n425 376.045
R2152 VPWR.n430 VPWR.n429 376.045
R2153 VPWR.n434 VPWR.n433 376.045
R2154 VPWR.n438 VPWR.n437 376.045
R2155 VPWR.n442 VPWR.n441 376.045
R2156 VPWR.n446 VPWR.n445 376.045
R2157 VPWR.n414 VPWR.n413 376.045
R2158 VPWR.n2448 VPWR.n2447 376.045
R2159 VPWR.n329 VPWR.n328 376.045
R2160 VPWR.n2542 VPWR.n2541 376.045
R2161 VPWR.n990 VPWR.n989 376.045
R2162 VPWR.n1508 VPWR.n1507 376.045
R2163 VPWR.n1216 VPWR.n1215 376.045
R2164 VPWR.n1860 VPWR.n1859 376.045
R2165 VPWR.n1850 VPWR.n1849 376.045
R2166 VPWR.n1848 VPWR.n1847 376.045
R2167 VPWR.n1840 VPWR.n1839 376.045
R2168 VPWR.n1838 VPWR.n1837 376.045
R2169 VPWR.n1830 VPWR.n1829 376.045
R2170 VPWR.n1828 VPWR.n1827 376.045
R2171 VPWR.n1820 VPWR.n1819 376.045
R2172 VPWR.n1858 VPWR.n1857 376.045
R2173 VPWR.n994 VPWR.n993 376.045
R2174 VPWR.n1520 VPWR.n1519 376.045
R2175 VPWR.n1213 VPWR.n1212 376.045
R2176 VPWR.n2468 VPWR.n2467 376.045
R2177 VPWR.n345 VPWR.n344 376.045
R2178 VPWR.n2518 VPWR.n2517 376.045
R2179 VPWR.n1481 VPWR.n1480 376.045
R2180 VPWR.n1182 VPWR.n1181 376.045
R2181 VPWR.n998 VPWR.n997 376.045
R2182 VPWR.n1522 VPWR.n1521 376.045
R2183 VPWR.n1205 VPWR.n1204 376.045
R2184 VPWR.n2438 VPWR.n2437 376.045
R2185 VPWR.n2428 VPWR.n2427 376.045
R2186 VPWR.n2426 VPWR.n2425 376.045
R2187 VPWR.n2418 VPWR.n2417 376.045
R2188 VPWR.n2416 VPWR.n2415 376.045
R2189 VPWR.n2408 VPWR.n2407 376.045
R2190 VPWR.n2436 VPWR.n2435 376.045
R2191 VPWR.n317 VPWR.n316 376.045
R2192 VPWR.n2556 VPWR.n2555 376.045
R2193 VPWR.n1537 VPWR.n1536 376.045
R2194 VPWR.n1202 VPWR.n1201 376.045
R2195 VPWR.n1002 VPWR.n1001 376.045
R2196 VPWR.n1006 VPWR.n1005 376.045
R2197 VPWR.n1010 VPWR.n1009 376.045
R2198 VPWR.n1014 VPWR.n1013 376.045
R2199 VPWR.n1018 VPWR.n1017 376.045
R2200 VPWR.n1022 VPWR.n1021 376.045
R2201 VPWR.n970 VPWR.n969 376.045
R2202 VPWR.n1475 VPWR.n1474 376.045
R2203 VPWR.n1593 VPWR.n1592 376.045
R2204 VPWR.n313 VPWR.n312 376.045
R2205 VPWR.n2566 VPWR.n2565 376.045
R2206 VPWR.n1199 VPWR.n1198 376.045
R2207 VPWR.n1762 VPWR.n1761 376.045
R2208 VPWR.n1191 VPWR.n1190 376.045
R2209 VPWR.n309 VPWR.n308 376.045
R2210 VPWR.n305 VPWR.n304 376.045
R2211 VPWR.n297 VPWR.n296 376.045
R2212 VPWR.n301 VPWR.n300 376.045
R2213 VPWR.n1741 VPWR.n1740 376.045
R2214 VPWR.n1750 VPWR.n1749 376.045
R2215 VPWR.n1791 VPWR.n1790 376.045
R2216 VPWR.n1760 VPWR.n1759 376.045
R2217 VPWR.n1188 VPWR.n1187 376.045
R2218 VPWR.n2578 VPWR.n2577 376.045
R2219 VPWR.n2580 VPWR.n2579 376.045
R2220 VPWR.n2590 VPWR.n2589 376.045
R2221 VPWR.n1739 VPWR.n1738 376.045
R2222 VPWR.n1339 VPWR.t1829 342.841
R2223 VPWR.n1378 VPWR.t1682 342.841
R2224 VPWR.n1415 VPWR.t967 342.841
R2225 VPWR.n2693 VPWR.t144 342.841
R2226 VPWR.n2656 VPWR.t1782 342.841
R2227 VPWR.n2599 VPWR.t1611 342.841
R2228 VPWR.n1339 VPWR.t1771 342.839
R2229 VPWR.n1378 VPWR.t101 342.839
R2230 VPWR.n1415 VPWR.t619 342.839
R2231 VPWR.n2693 VPWR.t1015 342.839
R2232 VPWR.n2656 VPWR.t55 342.839
R2233 VPWR.n2599 VPWR.t1899 342.839
R2234 VPWR.n2842 VPWR.n2824 339.212
R2235 VPWR.n1306 VPWR.t442 338.488
R2236 VPWR.n2729 VPWR.t293 338.488
R2237 VPWR.n1315 VPWR.n1314 327.377
R2238 VPWR.n1308 VPWR.n1307 327.377
R2239 VPWR.n1322 VPWR.n1321 327.377
R2240 VPWR.n1352 VPWR.n1350 327.377
R2241 VPWR.n1345 VPWR.n1343 327.377
R2242 VPWR.n1360 VPWR.n1358 327.377
R2243 VPWR.n1391 VPWR.n1389 327.377
R2244 VPWR.n1384 VPWR.n1382 327.377
R2245 VPWR.n1399 VPWR.n1397 327.377
R2246 VPWR.n1428 VPWR.n1426 327.377
R2247 VPWR.n1421 VPWR.n1419 327.377
R2248 VPWR.n1436 VPWR.n1434 327.377
R2249 VPWR.n1324 VPWR.n1323 327.375
R2250 VPWR.n1352 VPWR.n1351 327.375
R2251 VPWR.n1345 VPWR.n1344 327.375
R2252 VPWR.n1360 VPWR.n1359 327.375
R2253 VPWR.n1391 VPWR.n1390 327.375
R2254 VPWR.n1384 VPWR.n1383 327.375
R2255 VPWR.n1399 VPWR.n1398 327.375
R2256 VPWR.n1428 VPWR.n1427 327.375
R2257 VPWR.n1421 VPWR.n1420 327.375
R2258 VPWR.n1436 VPWR.n1435 327.375
R2259 VPWR.n1 VPWR 325.546
R2260 VPWR.n2667 VPWR.t143 322.262
R2261 VPWR.n2630 VPWR.t54 322.262
R2262 VPWR.n2805 VPWR.n2804 321.642
R2263 VPWR.n2722 VPWR.n2712 320.976
R2264 VPWR.n2716 VPWR.n2715 320.976
R2265 VPWR.n2710 VPWR.n2709 320.976
R2266 VPWR.n2680 VPWR.n2679 320.976
R2267 VPWR.n2686 VPWR.n2675 320.976
R2268 VPWR.n2672 VPWR.n2671 320.976
R2269 VPWR.n2643 VPWR.n2642 320.976
R2270 VPWR.n2649 VPWR.n2638 320.976
R2271 VPWR.n2635 VPWR.n2634 320.976
R2272 VPWR.n2610 VPWR.n2606 320.976
R2273 VPWR.n2614 VPWR.n2613 320.976
R2274 VPWR.n2620 VPWR.n2602 320.976
R2275 VPWR.n2727 VPWR.n2708 320.976
R2276 VPWR.n2680 VPWR.n2678 320.976
R2277 VPWR.n2686 VPWR.n2674 320.976
R2278 VPWR.n2672 VPWR.n2670 320.976
R2279 VPWR.n2643 VPWR.n2641 320.976
R2280 VPWR.n2649 VPWR.n2637 320.976
R2281 VPWR.n2635 VPWR.n2633 320.976
R2282 VPWR.n2610 VPWR.n2605 320.976
R2283 VPWR.n2614 VPWR.n2612 320.976
R2284 VPWR.n2620 VPWR.n2601 320.976
R2285 VPWR.n2801 VPWR 319.627
R2286 VPWR.n6 VPWR.n5 316.245
R2287 VPWR.n1241 VPWR.n1239 316.245
R2288 VPWR.n1264 VPWR.n1262 316.245
R2289 VPWR.n1288 VPWR.n1286 316.245
R2290 VPWR.n2784 VPWR.n2783 316.245
R2291 VPWR.n2764 VPWR.n2763 316.245
R2292 VPWR.n2745 VPWR.n2744 316.245
R2293 VPWR.n1241 VPWR.n1240 316.245
R2294 VPWR.n1264 VPWR.n1263 316.245
R2295 VPWR.n1288 VPWR.n1287 316.245
R2296 VPWR.n2784 VPWR.n2782 316.245
R2297 VPWR.n2764 VPWR.n2762 316.245
R2298 VPWR.n2745 VPWR.n2743 316.245
R2299 VPWR.n2630 VPWR.t237 313.87
R2300 VPWR.n10 VPWR.n4 310.502
R2301 VPWR.n1246 VPWR.n1238 310.502
R2302 VPWR.n1269 VPWR.n1261 310.502
R2303 VPWR.n1293 VPWR.n1285 310.502
R2304 VPWR.n2803 VPWR.n2802 310.502
R2305 VPWR.n2788 VPWR.n2787 310.502
R2306 VPWR.n2768 VPWR.n2767 310.502
R2307 VPWR.n2749 VPWR.n2748 310.502
R2308 VPWR.n1246 VPWR.n1245 310.5
R2309 VPWR.n1269 VPWR.n1268 310.5
R2310 VPWR.n1293 VPWR.n1292 310.5
R2311 VPWR.n2788 VPWR.n2786 310.5
R2312 VPWR.n2768 VPWR.n2766 310.5
R2313 VPWR.n2749 VPWR.n2747 310.5
R2314 VPWR.n2834 VPWR.n2833 279.341
R2315 VPWR.n2839 VPWR.n2838 279.341
R2316 VPWR.n1412 VPWR.t547 255.905
R2317 VPWR.n2663 VPWR.t884 255.905
R2318 VPWR.n1275 VPWR.t111 255.904
R2319 VPWR.n1412 VPWR.t1653 255.904
R2320 VPWR.n2774 VPWR.t431 255.904
R2321 VPWR.n2663 VPWR.t238 255.904
R2322 VPWR.n1303 VPWR.t840 254.019
R2323 VPWR.n2735 VPWR.t544 254.019
R2324 VPWR.n1335 VPWR.t838 252.948
R2325 VPWR.n2737 VPWR.t542 252.948
R2326 VPWR.n1373 VPWR.t711 250.722
R2327 VPWR.n2700 VPWR.t886 250.722
R2328 VPWR.n1310 VPWR.t376 249.901
R2329 VPWR.n1346 VPWR.t39 249.901
R2330 VPWR.n1385 VPWR.t1691 249.901
R2331 VPWR.n1422 VPWR.t43 249.901
R2332 VPWR.n2714 VPWR.t516 249.901
R2333 VPWR.n2677 VPWR.t513 249.901
R2334 VPWR.n2640 VPWR.t527 249.901
R2335 VPWR.n2607 VPWR.t481 249.901
R2336 VPWR.n1346 VPWR.t1689 249.901
R2337 VPWR.n1385 VPWR.t33 249.901
R2338 VPWR.n1422 VPWR.t1072 249.901
R2339 VPWR.n2677 VPWR.t526 249.901
R2340 VPWR.n2640 VPWR.t479 249.901
R2341 VPWR.n2607 VPWR.t502 249.901
R2342 VPWR.n1253 VPWR.t1832 249.363
R2343 VPWR.n1338 VPWR.t283 249.363
R2344 VPWR.n2811 VPWR.t1919 249.363
R2345 VPWR.n2795 VPWR.t689 249.363
R2346 VPWR.n2698 VPWR.t616 249.363
R2347 VPWR.n17 VPWR.t990 249.362
R2348 VPWR.n1253 VPWR.t1848 249.362
R2349 VPWR.n2795 VPWR.t1861 249.362
R2350 VPWR.t105 VPWR.t989 248.599
R2351 VPWR.t439 VPWR.t712 248.599
R2352 VPWR.t712 VPWR.t716 248.599
R2353 VPWR.t716 VPWR.t720 248.599
R2354 VPWR.t720 VPWR.t368 248.599
R2355 VPWR.t368 VPWR.t1890 248.599
R2356 VPWR.t1890 VPWR.t37 248.599
R2357 VPWR.t37 VPWR.t1694 248.599
R2358 VPWR.t371 VPWR.t373 248.599
R2359 VPWR.t373 VPWR.t375 248.599
R2360 VPWR.t529 VPWR.t505 248.599
R2361 VPWR.t493 VPWR.t529 248.599
R2362 VPWR.t467 VPWR.t493 248.599
R2363 VPWR.t290 VPWR.t467 248.599
R2364 VPWR.t50 VPWR.t290 248.599
R2365 VPWR.t1070 VPWR.t50 248.599
R2366 VPWR.t1912 VPWR.t1070 248.599
R2367 VPWR.t432 VPWR.t1918 248.599
R2368 VPWR.t473 VPWR.t515 248.599
R2369 VPWR.t521 VPWR.t473 248.599
R2370 VPWR.n15 VPWR.t106 247.394
R2371 VPWR.n1251 VPWR.t110 247.394
R2372 VPWR.n2809 VPWR.t433 247.394
R2373 VPWR.n2793 VPWR.t427 247.394
R2374 VPWR.n1251 VPWR.t107 247.394
R2375 VPWR.n2793 VPWR.t429 247.394
R2376 VPWR.n1304 VPWR.t380 244.737
R2377 VPWR.n2730 VPWR.t531 244.737
R2378 VPWR.n1374 VPWR.t100 243.886
R2379 VPWR.n2701 VPWR.t399 243.886
R2380 VPWR.n1277 VPWR.t988 243.512
R2381 VPWR.n1300 VPWR.t1833 243.512
R2382 VPWR.n1303 VPWR.t1869 243.512
R2383 VPWR.n2776 VPWR.t1921 243.512
R2384 VPWR.n2756 VPWR.t691 243.512
R2385 VPWR.n2735 VPWR.t614 243.512
R2386 VPWR.n1300 VPWR.t1849 243.512
R2387 VPWR.n2756 VPWR.t1860 243.512
R2388 VPWR.n1329 VPWR.t839 238.339
R2389 VPWR.n2705 VPWR.t543 238.339
R2390 VPWR.n2855 VPWR.t1560 237.99
R2391 VPWR.n2667 VPWR.t615 234.982
R2392 VPWR.t369 VPWR.t371 228.101
R2393 VPWR.t499 VPWR.t521 228.101
R2394 VPWR.n2801 VPWR 224.923
R2395 VPWR.n1 VPWR 219.004
R2396 VPWR.n1444 VPWR.n1443 214.613
R2397 VPWR.n1444 VPWR.n1442 214.613
R2398 VPWR.n1236 VPWR.n1235 214.326
R2399 VPWR.n1259 VPWR.n1258 214.326
R2400 VPWR.n1283 VPWR.n1282 214.326
R2401 VPWR.n1368 VPWR.n1367 214.326
R2402 VPWR.n1407 VPWR.n1406 214.326
R2403 VPWR.n1236 VPWR.n1234 214.326
R2404 VPWR.n1259 VPWR.n1257 214.326
R2405 VPWR.n1283 VPWR.n1281 214.326
R2406 VPWR.n1368 VPWR.n1366 214.326
R2407 VPWR.n1407 VPWR.n1405 214.326
R2408 VPWR.n2 VPWR.n1 213.119
R2409 VPWR.n2808 VPWR.n2801 213.119
R2410 VPWR VPWR.t105 207.166
R2411 VPWR.n2840 VPWR.n2839 204.424
R2412 VPWR.n2830 VPWR.n2817 204.424
R2413 VPWR.n2833 VPWR.n2820 204.424
R2414 VPWR.n2844 VPWR.n2841 204.048
R2415 VPWR VPWR.t1912 201.246
R2416 VPWR.t375 VPWR 189.409
R2417 VPWR.n2741 VPWR 184.63
R2418 VPWR.n1329 VPWR 182.952
R2419 VPWR.n2760 VPWR 182.952
R2420 VPWR.n2780 VPWR 181.273
R2421 VPWR.t237 VPWR 177.916
R2422 VPWR.n2848 VPWR.n2847 166.4
R2423 VPWR.n1770 VPWR.n1768 161.365
R2424 VPWR.n1041 VPWR.n1039 161.365
R2425 VPWR.n1545 VPWR.n1543 161.365
R2426 VPWR.n1550 VPWR.n1548 161.365
R2427 VPWR.n1555 VPWR.n1553 161.365
R2428 VPWR.n1560 VPWR.n1558 161.365
R2429 VPWR.n1565 VPWR.n1563 161.365
R2430 VPWR.n1570 VPWR.n1568 161.365
R2431 VPWR.n1575 VPWR.n1573 161.365
R2432 VPWR.n1580 VPWR.n1578 161.365
R2433 VPWR.n1135 VPWR.n1133 161.365
R2434 VPWR.n1460 VPWR.n1458 161.365
R2435 VPWR.n1455 VPWR.n1453 161.365
R2436 VPWR.n1775 VPWR.n1773 161.365
R2437 VPWR.n1783 VPWR.n1781 161.365
R2438 VPWR.n1779 VPWR.n1777 161.365
R2439 VPWR VPWR.n53 161.363
R2440 VPWR VPWR.n51 161.363
R2441 VPWR VPWR.n49 161.363
R2442 VPWR VPWR.n47 161.363
R2443 VPWR VPWR.n45 161.363
R2444 VPWR VPWR.n43 161.363
R2445 VPWR VPWR.n41 161.363
R2446 VPWR VPWR.n39 161.363
R2447 VPWR VPWR.n37 161.363
R2448 VPWR VPWR.n35 161.363
R2449 VPWR VPWR.n33 161.363
R2450 VPWR VPWR.n31 161.363
R2451 VPWR VPWR.n29 161.363
R2452 VPWR VPWR.n27 161.363
R2453 VPWR VPWR.n25 161.363
R2454 VPWR VPWR.n23 161.363
R2455 VPWR.n1115 VPWR.n1114 161.303
R2456 VPWR.n107 VPWR.n106 161.303
R2457 VPWR.n1120 VPWR.n1119 161.3
R2458 VPWR.n1599 VPWR.n1598 161.3
R2459 VPWR.n1602 VPWR.n1601 161.3
R2460 VPWR.n1111 VPWR.n1110 161.3
R2461 VPWR.n1126 VPWR.n1125 161.3
R2462 VPWR.n1107 VPWR.n1106 161.3
R2463 VPWR.n1612 VPWR.n1611 161.3
R2464 VPWR.n1615 VPWR.n1614 161.3
R2465 VPWR.n1618 VPWR.n1617 161.3
R2466 VPWR.n1623 VPWR.n1622 161.3
R2467 VPWR.n1626 VPWR.n1625 161.3
R2468 VPWR.n1629 VPWR.n1628 161.3
R2469 VPWR.n1101 VPWR.n1100 161.3
R2470 VPWR.n1177 VPWR.n1176 161.3
R2471 VPWR.n1097 VPWR.n1096 161.3
R2472 VPWR.n1639 VPWR.n1638 161.3
R2473 VPWR.n1642 VPWR.n1641 161.3
R2474 VPWR.n1645 VPWR.n1644 161.3
R2475 VPWR.n1650 VPWR.n1649 161.3
R2476 VPWR.n1653 VPWR.n1652 161.3
R2477 VPWR.n1656 VPWR.n1655 161.3
R2478 VPWR.n1091 VPWR.n1090 161.3
R2479 VPWR.n1209 VPWR.n1208 161.3
R2480 VPWR.n1087 VPWR.n1086 161.3
R2481 VPWR.n1666 VPWR.n1665 161.3
R2482 VPWR.n1669 VPWR.n1668 161.3
R2483 VPWR.n1672 VPWR.n1671 161.3
R2484 VPWR.n1677 VPWR.n1676 161.3
R2485 VPWR.n1680 VPWR.n1679 161.3
R2486 VPWR.n1683 VPWR.n1682 161.3
R2487 VPWR.n1081 VPWR.n1080 161.3
R2488 VPWR.n1195 VPWR.n1194 161.3
R2489 VPWR.n1077 VPWR.n1076 161.3
R2490 VPWR.n1693 VPWR.n1692 161.3
R2491 VPWR.n1696 VPWR.n1695 161.3
R2492 VPWR.n1699 VPWR.n1698 161.3
R2493 VPWR.n1704 VPWR.n1703 161.3
R2494 VPWR.n1707 VPWR.n1706 161.3
R2495 VPWR.n1710 VPWR.n1709 161.3
R2496 VPWR.n1070 VPWR.n1069 161.3
R2497 VPWR.n1719 VPWR.n1718 161.3
R2498 VPWR.n1722 VPWR.n1721 161.3
R2499 VPWR.n1717 VPWR.n1716 161.3
R2500 VPWR.n1734 VPWR.n1733 161.3
R2501 VPWR.n1117 VPWR.n1116 161.3
R2502 VPWR.n1731 VPWR.n1730 161.3
R2503 VPWR.n1065 VPWR.n1064 161.3
R2504 VPWR.n126 VPWR.n125 161.3
R2505 VPWR.n117 VPWR.n116 161.3
R2506 VPWR.n120 VPWR.n119 161.3
R2507 VPWR.n115 VPWR.n114 161.3
R2508 VPWR.n138 VPWR.n137 161.3
R2509 VPWR.n128 VPWR.n127 161.3
R2510 VPWR.n109 VPWR.n108 161.3
R2511 VPWR.n105 VPWR.n104 161.3
R2512 VPWR.n288 VPWR.n287 161.3
R2513 VPWR.n285 VPWR.n284 161.3
R2514 VPWR.n101 VPWR.n100 161.3
R2515 VPWR.n272 VPWR.n271 161.3
R2516 VPWR.n275 VPWR.n274 161.3
R2517 VPWR.n270 VPWR.n269 161.3
R2518 VPWR.n260 VPWR.n259 161.3
R2519 VPWR.n263 VPWR.n262 161.3
R2520 VPWR.n258 VPWR.n257 161.3
R2521 VPWR.n248 VPWR.n247 161.3
R2522 VPWR.n251 VPWR.n250 161.3
R2523 VPWR.n246 VPWR.n245 161.3
R2524 VPWR.n236 VPWR.n235 161.3
R2525 VPWR.n239 VPWR.n238 161.3
R2526 VPWR.n234 VPWR.n233 161.3
R2527 VPWR.n224 VPWR.n223 161.3
R2528 VPWR.n227 VPWR.n226 161.3
R2529 VPWR.n222 VPWR.n221 161.3
R2530 VPWR.n212 VPWR.n211 161.3
R2531 VPWR.n215 VPWR.n214 161.3
R2532 VPWR.n210 VPWR.n209 161.3
R2533 VPWR.n200 VPWR.n199 161.3
R2534 VPWR.n203 VPWR.n202 161.3
R2535 VPWR.n198 VPWR.n197 161.3
R2536 VPWR.n188 VPWR.n187 161.3
R2537 VPWR.n191 VPWR.n190 161.3
R2538 VPWR.n186 VPWR.n185 161.3
R2539 VPWR.n176 VPWR.n175 161.3
R2540 VPWR.n179 VPWR.n178 161.3
R2541 VPWR.n174 VPWR.n173 161.3
R2542 VPWR.n164 VPWR.n163 161.3
R2543 VPWR.n167 VPWR.n166 161.3
R2544 VPWR.n162 VPWR.n161 161.3
R2545 VPWR.n152 VPWR.n151 161.3
R2546 VPWR.n155 VPWR.n154 161.3
R2547 VPWR.n150 VPWR.n149 161.3
R2548 VPWR.n140 VPWR.n139 161.3
R2549 VPWR.n143 VPWR.n142 161.3
R2550 VPWR.n131 VPWR.n130 161.3
R2551 VPWR.n1601 VPWR.t1123 161.202
R2552 VPWR.n1106 VPWR.t1248 161.202
R2553 VPWR.n1617 VPWR.t1289 161.202
R2554 VPWR.n1628 VPWR.t1397 161.202
R2555 VPWR.n1096 VPWR.t1164 161.202
R2556 VPWR.n1644 VPWR.t1179 161.202
R2557 VPWR.n1655 VPWR.t1402 161.202
R2558 VPWR.n1086 VPWR.t1445 161.202
R2559 VPWR.n1671 VPWR.t1162 161.202
R2560 VPWR.n1682 VPWR.t1315 161.202
R2561 VPWR.n1076 VPWR.t1337 161.202
R2562 VPWR.n1698 VPWR.t1187 161.202
R2563 VPWR.n1709 VPWR.t1213 161.202
R2564 VPWR.n1721 VPWR.t1238 161.202
R2565 VPWR.n1116 VPWR.t1378 161.202
R2566 VPWR.n1730 VPWR.t1086 161.202
R2567 VPWR.n119 VPWR.t1205 161.202
R2568 VPWR.n108 VPWR.t1104 161.202
R2569 VPWR.n284 VPWR.t1240 161.202
R2570 VPWR.n274 VPWR.t1370 161.202
R2571 VPWR.n262 VPWR.t1410 161.202
R2572 VPWR.n250 VPWR.t1134 161.202
R2573 VPWR.n238 VPWR.t1278 161.202
R2574 VPWR.n226 VPWR.t1302 161.202
R2575 VPWR.n214 VPWR.t1139 161.202
R2576 VPWR.n202 VPWR.t1174 161.202
R2577 VPWR.n190 VPWR.t1276 161.202
R2578 VPWR.n178 VPWR.t1437 161.202
R2579 VPWR.n166 VPWR.t1456 161.202
R2580 VPWR.n154 VPWR.t1310 161.202
R2581 VPWR.n1768 VPWR.t1362 161.202
R2582 VPWR.n1039 VPWR.t1118 161.202
R2583 VPWR.n1543 VPWR.t1099 161.202
R2584 VPWR.n1548 VPWR.t1348 161.202
R2585 VPWR.n1553 VPWR.t1230 161.202
R2586 VPWR.n1558 VPWR.t1200 161.202
R2587 VPWR.n1563 VPWR.t1352 161.202
R2588 VPWR.n1568 VPWR.t1350 161.202
R2589 VPWR.n1573 VPWR.t1195 161.202
R2590 VPWR.n1578 VPWR.t1088 161.202
R2591 VPWR.n1133 VPWR.t1429 161.202
R2592 VPWR.n1458 VPWR.t1300 161.202
R2593 VPWR.n1453 VPWR.t1169 161.202
R2594 VPWR.n1773 VPWR.t1380 161.202
R2595 VPWR.n1781 VPWR.t1418 161.202
R2596 VPWR.n1777 VPWR.t1250 161.202
R2597 VPWR.n142 VPWR.t1329 161.202
R2598 VPWR.n130 VPWR.t1354 161.202
R2599 VPWR.n1119 VPWR.t1106 161.106
R2600 VPWR.n1110 VPWR.t1242 161.106
R2601 VPWR.n1611 VPWR.t1255 161.106
R2602 VPWR.n1622 VPWR.t1415 161.106
R2603 VPWR.n1100 VPWR.t1136 161.106
R2604 VPWR.n1638 VPWR.t1283 161.106
R2605 VPWR.n1649 VPWR.t1391 161.106
R2606 VPWR.n1090 VPWR.t1431 161.106
R2607 VPWR.n1665 VPWR.t1176 161.106
R2608 VPWR.n1676 VPWR.t1280 161.106
R2609 VPWR.n1080 VPWR.t1439 161.106
R2610 VPWR.n1692 VPWR.t1458 161.106
R2611 VPWR.n1703 VPWR.t1202 161.106
R2612 VPWR.n1069 VPWR.t1331 161.106
R2613 VPWR.n1716 VPWR.t1359 161.106
R2614 VPWR.n1064 VPWR.t1210 161.106
R2615 VPWR.n125 VPWR.t1090 161.106
R2616 VPWR.n114 VPWR.t1326 161.106
R2617 VPWR.n137 VPWR.t1450 161.106
R2618 VPWR.n104 VPWR.t1235 161.106
R2619 VPWR.n100 VPWR.t1364 161.106
R2620 VPWR.n269 VPWR.t1382 161.106
R2621 VPWR.n257 VPWR.t1144 161.106
R2622 VPWR.n245 VPWR.t1252 161.106
R2623 VPWR.n233 VPWR.t1407 161.106
R2624 VPWR.n221 VPWR.t1131 161.106
R2625 VPWR.n209 VPWR.t1166 161.106
R2626 VPWR.n197 VPWR.t1294 161.106
R2627 VPWR.n185 VPWR.t1404 161.106
R2628 VPWR.n173 VPWR.t1171 161.106
R2629 VPWR.n161 VPWR.t1189 161.106
R2630 VPWR.n149 VPWR.t1317 161.106
R2631 VPWR.n53 VPWR.t1434 161.106
R2632 VPWR.n51 VPWR.t1394 161.106
R2633 VPWR.n49 VPWR.t1112 161.106
R2634 VPWR.n47 VPWR.t1224 161.106
R2635 VPWR.n45 VPWR.t1442 161.106
R2636 VPWR.n43 VPWR.t1291 161.106
R2637 VPWR.n41 VPWR.t1399 161.106
R2638 VPWR.n39 VPWR.t1125 161.106
R2639 VPWR.n37 VPWR.t1232 161.106
R2640 VPWR.n35 VPWR.t1192 161.106
R2641 VPWR.n33 VPWR.t1297 161.106
R2642 VPWR.n31 VPWR.t1120 161.106
R2643 VPWR.n29 VPWR.t1304 161.106
R2644 VPWR.n27 VPWR.t1412 161.106
R2645 VPWR.n25 VPWR.t1264 161.106
R2646 VPWR.n23 VPWR.t1375 161.106
R2647 VPWR.n1598 VPWR.t1156 159.978
R2648 VPWR.n1125 VPWR.t1261 159.978
R2649 VPWR.n1614 VPWR.t1423 159.978
R2650 VPWR.n1625 VPWR.t1141 159.978
R2651 VPWR.n1176 VPWR.t1153 159.978
R2652 VPWR.n1641 VPWR.t1312 159.978
R2653 VPWR.n1652 VPWR.t1420 159.978
R2654 VPWR.n1208 VPWR.t1181 159.978
R2655 VPWR.n1668 VPWR.t1207 159.978
R2656 VPWR.n1679 VPWR.t1334 159.978
R2657 VPWR.n1194 VPWR.t1080 159.978
R2658 VPWR.n1695 VPWR.t1101 159.978
R2659 VPWR.n1706 VPWR.t1339 159.978
R2660 VPWR.n1718 VPWR.t1367 159.978
R2661 VPWR.n1733 VPWR.t1083 159.978
R2662 VPWR.n1114 VPWR.t1388 159.978
R2663 VPWR.n116 VPWR.t1221 159.978
R2664 VPWR.n127 VPWR.t1096 159.978
R2665 VPWR.n106 VPWR.t1128 159.978
R2666 VPWR.n287 VPWR.t1273 159.978
R2667 VPWR.n271 VPWR.t1385 159.978
R2668 VPWR.n259 VPWR.t1150 159.978
R2669 VPWR.n247 VPWR.t1258 159.978
R2670 VPWR.n235 VPWR.t1270 159.978
R2671 VPWR.n223 VPWR.t1426 159.978
R2672 VPWR.n211 VPWR.t1147 159.978
R2673 VPWR.n199 VPWR.t1307 159.978
R2674 VPWR.n187 VPWR.t1323 159.978
R2675 VPWR.n175 VPWR.t1453 159.978
R2676 VPWR.n163 VPWR.t1197 159.978
R2677 VPWR.n151 VPWR.t1227 159.978
R2678 VPWR.n1228 VPWR.t1184 159.978
R2679 VPWR.n1150 VPWR.t1115 159.978
R2680 VPWR.n1224 VPWR.t1320 159.978
R2681 VPWR.n1482 VPWR.t1218 159.978
R2682 VPWR.n1170 VPWR.t1342 159.978
R2683 VPWR.n1166 VPWR.t1093 159.978
R2684 VPWR.n1160 VPWR.t1215 159.978
R2685 VPWR.n1476 VPWR.t1447 159.978
R2686 VPWR.n1156 VPWR.t1356 159.978
R2687 VPWR.n1146 VPWR.t1372 159.978
R2688 VPWR.n1469 VPWR.t1345 159.978
R2689 VPWR.n1046 VPWR.t1245 159.978
R2690 VPWR.n1745 VPWR.t1109 159.978
R2691 VPWR.n1033 VPWR.t1159 159.978
R2692 VPWR.n1029 VPWR.t1267 159.978
R2693 VPWR.n1050 VPWR.t1286 159.978
R2694 VPWR.n139 VPWR.t1077 159.978
R2695 VPWR.n1229 VPWR.n1228 152
R2696 VPWR.n1151 VPWR.n1150 152
R2697 VPWR.n1225 VPWR.n1224 152
R2698 VPWR.n1483 VPWR.n1482 152
R2699 VPWR.n1171 VPWR.n1170 152
R2700 VPWR.n1167 VPWR.n1166 152
R2701 VPWR.n1161 VPWR.n1160 152
R2702 VPWR.n1477 VPWR.n1476 152
R2703 VPWR.n1157 VPWR.n1156 152
R2704 VPWR.n1147 VPWR.n1146 152
R2705 VPWR.n1470 VPWR.n1469 152
R2706 VPWR.n1047 VPWR.n1046 152
R2707 VPWR.n1746 VPWR.n1745 152
R2708 VPWR.n1034 VPWR.n1033 152
R2709 VPWR.n1030 VPWR.n1029 152
R2710 VPWR.n1051 VPWR.n1050 152
R2711 VPWR.n2845 VPWR.n2844 150.213
R2712 VPWR.n1601 VPWR.t2063 145.137
R2713 VPWR.n1106 VPWR.t2014 145.137
R2714 VPWR.n1617 VPWR.t2000 145.137
R2715 VPWR.n1628 VPWR.t1962 145.137
R2716 VPWR.n1096 VPWR.t2049 145.137
R2717 VPWR.n1644 VPWR.t2042 145.137
R2718 VPWR.n1655 VPWR.t1959 145.137
R2719 VPWR.n1086 VPWR.t1945 145.137
R2720 VPWR.n1671 VPWR.t2050 145.137
R2721 VPWR.n1682 VPWR.t1993 145.137
R2722 VPWR.n1076 VPWR.t1988 145.137
R2723 VPWR.n1698 VPWR.t2040 145.137
R2724 VPWR.n1709 VPWR.t2033 145.137
R2725 VPWR.n1721 VPWR.t2019 145.137
R2726 VPWR.n1116 VPWR.t1969 145.137
R2727 VPWR.n1730 VPWR.t1937 145.137
R2728 VPWR.n119 VPWR.t2048 145.137
R2729 VPWR.n108 VPWR.t1934 145.137
R2730 VPWR.n284 VPWR.t2030 145.137
R2731 VPWR.n274 VPWR.t1983 145.137
R2732 VPWR.n262 VPWR.t1971 145.137
R2733 VPWR.n250 VPWR.t1930 145.137
R2734 VPWR.n238 VPWR.t2016 145.137
R2735 VPWR.n226 VPWR.t2008 145.137
R2736 VPWR.n214 VPWR.t1928 145.137
R2737 VPWR.n202 VPWR.t2057 145.137
R2738 VPWR.n190 VPWR.t2017 145.137
R2739 VPWR.n178 VPWR.t1961 145.137
R2740 VPWR.n166 VPWR.t1952 145.137
R2741 VPWR.n154 VPWR.t2007 145.137
R2742 VPWR.n1768 VPWR.t1976 145.137
R2743 VPWR.n1039 VPWR.t2065 145.137
R2744 VPWR.n1543 VPWR.t1929 145.137
R2745 VPWR.n1548 VPWR.t1986 145.137
R2746 VPWR.n1553 VPWR.t2025 145.137
R2747 VPWR.n1558 VPWR.t2037 145.137
R2748 VPWR.n1563 VPWR.t1979 145.137
R2749 VPWR.n1568 VPWR.t1985 145.137
R2750 VPWR.n1573 VPWR.t2039 145.137
R2751 VPWR.n1578 VPWR.t1936 145.137
R2752 VPWR.n1133 VPWR.t1950 145.137
R2753 VPWR.n1458 VPWR.t1996 145.137
R2754 VPWR.n1453 VPWR.t2045 145.137
R2755 VPWR.n1773 VPWR.t1968 145.137
R2756 VPWR.n1781 VPWR.t1953 145.137
R2757 VPWR.n1777 VPWR.t2013 145.137
R2758 VPWR.n142 VPWR.t1999 145.137
R2759 VPWR.n130 VPWR.t1990 145.137
R2760 VPWR.n1119 VPWR.t2067 145.038
R2761 VPWR.n1110 VPWR.t2018 145.038
R2762 VPWR.n1611 VPWR.t2010 145.038
R2763 VPWR.n1622 VPWR.t1955 145.038
R2764 VPWR.n1100 VPWR.t2059 145.038
R2765 VPWR.n1638 VPWR.t2002 145.038
R2766 VPWR.n1649 VPWR.t1964 145.038
R2767 VPWR.n1090 VPWR.t1949 145.038
R2768 VPWR.n1665 VPWR.t2043 145.038
R2769 VPWR.n1676 VPWR.t2003 145.038
R2770 VPWR.n1080 VPWR.t1947 145.038
R2771 VPWR.n1692 VPWR.t1939 145.038
R2772 VPWR.n1703 VPWR.t2036 145.038
R2773 VPWR.n1069 VPWR.t1989 145.038
R2774 VPWR.n1716 VPWR.t1977 145.038
R2775 VPWR.n1064 VPWR.t2034 145.038
R2776 VPWR.n125 VPWR.t1940 145.038
R2777 VPWR.n114 VPWR.t2001 145.038
R2778 VPWR.n137 VPWR.t1954 145.038
R2779 VPWR.n104 VPWR.t2032 145.038
R2780 VPWR.n100 VPWR.t1987 145.038
R2781 VPWR.n269 VPWR.t1980 145.038
R2782 VPWR.n257 VPWR.t2068 145.038
R2783 VPWR.n245 VPWR.t2027 145.038
R2784 VPWR.n233 VPWR.t1972 145.038
R2785 VPWR.n221 VPWR.t1931 145.038
R2786 VPWR.n209 VPWR.t2060 145.038
R2787 VPWR.n197 VPWR.t2009 145.038
R2788 VPWR.n185 VPWR.t1973 145.038
R2789 VPWR.n173 VPWR.t2058 145.038
R2790 VPWR.n161 VPWR.t2052 145.038
R2791 VPWR.n149 VPWR.t2004 145.038
R2792 VPWR.n53 VPWR.t2053 145.038
R2793 VPWR.n51 VPWR.t1963 145.038
R2794 VPWR.n49 VPWR.t2066 145.038
R2795 VPWR.n47 VPWR.t2026 145.038
R2796 VPWR.n45 VPWR.t1946 145.038
R2797 VPWR.n43 VPWR.t2051 145.038
R2798 VPWR.n41 VPWR.t2069 145.038
R2799 VPWR.n39 VPWR.t2028 145.038
R2800 VPWR.n37 VPWR.t2022 145.038
R2801 VPWR.n35 VPWR.t1943 145.038
R2802 VPWR.n33 VPWR.t1997 145.038
R2803 VPWR.n31 VPWR.t2064 145.038
R2804 VPWR.n29 VPWR.t1995 145.038
R2805 VPWR.n27 VPWR.t1956 145.038
R2806 VPWR.n25 VPWR.t2021 145.038
R2807 VPWR.n23 VPWR.t1970 145.038
R2808 VPWR.n1598 VPWR.t1966 143.911
R2809 VPWR.n1125 VPWR.t2062 143.911
R2810 VPWR.n1614 VPWR.t2047 143.911
R2811 VPWR.n1625 VPWR.t1965 143.911
R2812 VPWR.n1176 VPWR.t1958 143.911
R2813 VPWR.n1641 VPWR.t1944 143.911
R2814 VPWR.n1652 VPWR.t2005 143.911
R2815 VPWR.n1208 VPWR.t1992 143.911
R2816 VPWR.n1668 VPWR.t1941 143.911
R2817 VPWR.n1679 VPWR.t2038 143.911
R2818 VPWR.n1194 VPWR.t2031 143.911
R2819 VPWR.n1695 VPWR.t1978 143.911
R2820 VPWR.n1706 VPWR.t1935 143.911
R2821 VPWR.n1718 VPWR.t2024 143.911
R2822 VPWR.n1733 VPWR.t1984 143.911
R2823 VPWR.n1114 VPWR.t2012 143.911
R2824 VPWR.n116 VPWR.t1951 143.911
R2825 VPWR.n127 VPWR.t1991 143.911
R2826 VPWR.n106 VPWR.t1981 143.911
R2827 VPWR.n287 VPWR.t1933 143.911
R2828 VPWR.n271 VPWR.t2029 143.911
R2829 VPWR.n259 VPWR.t2015 143.911
R2830 VPWR.n247 VPWR.t1932 143.911
R2831 VPWR.n235 VPWR.t1926 143.911
R2832 VPWR.n223 VPWR.t2056 143.911
R2833 VPWR.n211 VPWR.t1974 143.911
R2834 VPWR.n199 VPWR.t1960 143.911
R2835 VPWR.n187 VPWR.t2054 143.911
R2836 VPWR.n175 VPWR.t2006 143.911
R2837 VPWR.n163 VPWR.t1998 143.911
R2838 VPWR.n151 VPWR.t1942 143.911
R2839 VPWR.n1228 VPWR.t1948 143.911
R2840 VPWR.n1150 VPWR.t1975 143.911
R2841 VPWR.n1224 VPWR.t2041 143.911
R2842 VPWR.n1482 VPWR.t1982 143.911
R2843 VPWR.n1170 VPWR.t2035 143.911
R2844 VPWR.n1166 VPWR.t2023 143.911
R2845 VPWR.n1160 VPWR.t1938 143.911
R2846 VPWR.n1476 VPWR.t1994 143.911
R2847 VPWR.n1156 VPWR.t1927 143.911
R2848 VPWR.n1146 VPWR.t2020 143.911
R2849 VPWR.n1469 VPWR.t2044 143.911
R2850 VPWR.n1046 VPWR.t1967 143.911
R2851 VPWR.n1745 VPWR.t2011 143.911
R2852 VPWR.n1033 VPWR.t1957 143.911
R2853 VPWR.n1029 VPWR.t2061 143.911
R2854 VPWR.n1050 VPWR.t2055 143.911
R2855 VPWR.n139 VPWR.t2046 143.911
R2856 VPWR.t718 VPWR.t369 140.989
R2857 VPWR.t484 VPWR.t471 140.989
R2858 VPWR.t511 VPWR.t484 140.989
R2859 VPWR.t487 VPWR.t511 140.989
R2860 VPWR.t342 VPWR.t487 140.989
R2861 VPWR.t133 VPWR.t342 140.989
R2862 VPWR.t1011 VPWR.t133 140.989
R2863 VPWR.t548 VPWR.t1011 140.989
R2864 VPWR.t426 VPWR.t688 140.989
R2865 VPWR.t523 VPWR.t490 140.989
R2866 VPWR.t477 VPWR.t523 140.989
R2867 VPWR.t524 VPWR.t477 140.989
R2868 VPWR.t1523 VPWR.t524 140.989
R2869 VPWR.t52 VPWR.t1523 140.989
R2870 VPWR.t48 VPWR.t52 140.989
R2871 VPWR.t46 VPWR.t48 140.989
R2872 VPWR.t468 VPWR.t509 140.989
R2873 VPWR.t498 VPWR.t468 140.989
R2874 VPWR.t472 VPWR.t498 140.989
R2875 VPWR.t1614 VPWR.t472 140.989
R2876 VPWR.t1612 VPWR.t1614 140.989
R2877 VPWR.t1618 VPWR.t1612 140.989
R2878 VPWR.t1606 VPWR.t1618 140.989
R2879 VPWR.t649 VPWR.t499 140.989
R2880 VPWR.t469 VPWR.t512 140.989
R2881 VPWR.t519 VPWR.t469 140.989
R2882 VPWR.t496 VPWR.t519 140.989
R2883 VPWR.t413 VPWR.t496 140.989
R2884 VPWR.t651 VPWR.t413 140.989
R2885 VPWR.t1018 VPWR.t651 140.989
R2886 VPWR.t143 VPWR.t1018 140.989
R2887 VPWR.t491 VPWR.t478 140.989
R2888 VPWR.t465 VPWR.t491 140.989
R2889 VPWR.t517 VPWR.t465 140.989
R2890 VPWR.t1527 VPWR.t517 140.989
R2891 VPWR.t56 VPWR.t1527 140.989
R2892 VPWR.t1525 VPWR.t56 140.989
R2893 VPWR.t54 VPWR.t1525 140.989
R2894 VPWR.t488 VPWR.t480 140.989
R2895 VPWR.t494 VPWR.t488 140.989
R2896 VPWR.t482 VPWR.t494 140.989
R2897 VPWR.t1616 VPWR.t482 140.989
R2898 VPWR.t1620 VPWR.t1616 140.989
R2899 VPWR.t1608 VPWR.t1620 140.989
R2900 VPWR.t1610 VPWR.t1608 140.989
R2901 VPWR VPWR.n1442 133.312
R2902 VPWR.n2841 VPWR.n2840 129.13
R2903 VPWR.n2858 VPWR.n2819 129.13
R2904 VPWR.n2780 VPWR 127.562
R2905 VPWR.n2760 VPWR 127.562
R2906 VPWR.n2741 VPWR 127.562
R2907 VPWR VPWR.t530 125.883
R2908 VPWR.n2705 VPWR 125.883
R2909 VPWR.t428 VPWR.t690 120.849
R2910 VPWR.t1868 VPWR.t837 117.492
R2911 VPWR.t613 VPWR.t541 117.492
R2912 VPWR.t398 VPWR 115.814
R2913 VPWR VPWR.t548 114.135
R2914 VPWR VPWR.t46 114.135
R2915 VPWR VPWR.t1606 114.135
R2916 VPWR.n2859 VPWR.n2817 111.059
R2917 VPWR.t1778 VPWR 107.421
R2918 VPWR.n1330 VPWR.n1329 106.561
R2919 VPWR.n2781 VPWR.n2780 106.561
R2920 VPWR.n2761 VPWR.n2760 106.561
R2921 VPWR.n2742 VPWR.n2741 106.561
R2922 VPWR.n2706 VPWR.n2705 106.561
R2923 VPWR.n2668 VPWR.n2667 106.561
R2924 VPWR.n2631 VPWR.n2630 106.561
R2925 VPWR VPWR.t432 106.543
R2926 VPWR VPWR.n1234 104.8
R2927 VPWR VPWR.n1257 104.8
R2928 VPWR VPWR.n1281 104.8
R2929 VPWR VPWR.n1366 104.8
R2930 VPWR VPWR.n1405 104.8
R2931 VPWR.n1443 VPWR 100.883
R2932 VPWR VPWR.t439 100.624
R2933 VPWR.t447 VPWR.t1560 97.9386
R2934 VPWR.n2859 VPWR.n2858 93.3652
R2935 VPWR.n1231 VPWR.n1230 91.8492
R2936 VPWR.n1153 VPWR.n1152 91.8492
R2937 VPWR.n1227 VPWR.n1226 91.8492
R2938 VPWR.n1485 VPWR.n1484 91.8492
R2939 VPWR.n1173 VPWR.n1172 91.8492
R2940 VPWR.n1169 VPWR.n1168 91.8492
R2941 VPWR.n1163 VPWR.n1162 91.8492
R2942 VPWR.n1479 VPWR.n1478 91.8492
R2943 VPWR.n1159 VPWR.n1158 91.8492
R2944 VPWR.n1149 VPWR.n1148 91.8492
R2945 VPWR.n1472 VPWR.n1471 91.8492
R2946 VPWR.n1049 VPWR.n1048 91.8492
R2947 VPWR.n1748 VPWR.n1747 91.8492
R2948 VPWR.n1036 VPWR.n1035 91.8492
R2949 VPWR.n1032 VPWR.n1031 91.8492
R2950 VPWR.n1053 VPWR.n1052 91.8492
R2951 VPWR.n2847 VPWR.n2820 91.4829
R2952 VPWR.t447 VPWR.n2842 90.0872
R2953 VPWR.t515 VPWR 88.7855
R2954 VPWR.n1235 VPWR 79.407
R2955 VPWR.n1258 VPWR 79.407
R2956 VPWR.n1282 VPWR 79.407
R2957 VPWR.n1367 VPWR 79.407
R2958 VPWR.n1406 VPWR 79.407
R2959 VPWR.t615 VPWR.t885 78.8874
R2960 VPWR.n2840 VPWR.n2818 74.9181
R2961 VPWR.n2858 VPWR.n2818 74.9181
R2962 VPWR.n2858 VPWR.n2857 74.9181
R2963 VPWR.n2857 VPWR.n2820 74.9181
R2964 VPWR.t379 VPWR.t441 70.4952
R2965 VPWR.t441 VPWR.t381 70.4952
R2966 VPWR.t381 VPWR.t714 70.4952
R2967 VPWR.t714 VPWR.t608 70.4952
R2968 VPWR.t608 VPWR.t437 70.4952
R2969 VPWR.t437 VPWR.t1888 70.4952
R2970 VPWR.t1888 VPWR.t718 70.4952
R2971 VPWR.t503 VPWR.t649 70.4952
R2972 VPWR.t545 VPWR.t503 70.4952
R2973 VPWR.t475 VPWR.t545 70.4952
R2974 VPWR.t1066 VPWR.t475 70.4952
R2975 VPWR.t507 VPWR.t1066 70.4952
R2976 VPWR.t292 VPWR.t507 70.4952
R2977 VPWR.t530 VPWR.t292 70.4952
R2978 VPWR VPWR.t379 68.8168
R2979 VPWR.t434 VPWR.t430 68.8168
R2980 VPWR.t885 VPWR.t398 62.103
R2981 VPWR VPWR.t426 60.4245
R2982 VPWR.n2849 VPWR.n2842 59.762
R2983 VPWR.n2845 VPWR.n2819 53.8358
R2984 VPWR.t430 VPWR.t1920 52.0323
R2985 VPWR.t415 VPWR 50.3539
R2986 VPWR VPWR.t434 50.3539
R2987 VPWR VPWR.t428 50.3539
R2988 VPWR.t512 VPWR 50.3539
R2989 VPWR.t478 VPWR 50.3539
R2990 VPWR.t480 VPWR 50.3539
R2991 VPWR.n2854 VPWR.n2818 46.2505
R2992 VPWR.n2855 VPWR.n2854 46.2505
R2993 VPWR.n2835 VPWR.n2834 46.2505
R2994 VPWR.n2836 VPWR.n2835 46.2505
R2995 VPWR.n2838 VPWR.n2837 46.2505
R2996 VPWR.n2837 VPWR.n2836 46.2505
R2997 VPWR.n2844 VPWR.n2824 46.2505
R2998 VPWR.n2857 VPWR.n2856 46.2505
R2999 VPWR.n2856 VPWR.n2855 46.2505
R3000 VPWR.n2849 VPWR.n2848 46.2505
R3001 VPWR.n2846 VPWR.n2845 45.9299
R3002 VPWR.n2832 VPWR.n2830 44.8005
R3003 VPWR.n2830 VPWR.n2826 44.8005
R3004 VPWR.n2847 VPWR.n2843 37.0005
R3005 VPWR.n2843 VPWR.t1560 37.0005
R3006 VPWR.n1230 VPWR.n1229 34.7473
R3007 VPWR.n1152 VPWR.n1151 34.7473
R3008 VPWR.n1226 VPWR.n1225 34.7473
R3009 VPWR.n1484 VPWR.n1483 34.7473
R3010 VPWR.n1172 VPWR.n1171 34.7473
R3011 VPWR.n1168 VPWR.n1167 34.7473
R3012 VPWR.n1162 VPWR.n1161 34.7473
R3013 VPWR.n1478 VPWR.n1477 34.7473
R3014 VPWR.n1158 VPWR.n1157 34.7473
R3015 VPWR.n1148 VPWR.n1147 34.7473
R3016 VPWR.n1471 VPWR.n1470 34.7473
R3017 VPWR.n1048 VPWR.n1047 34.7473
R3018 VPWR.n1747 VPWR.n1746 34.7473
R3019 VPWR.n1035 VPWR.n1034 34.7473
R3020 VPWR.n1031 VPWR.n1030 34.7473
R3021 VPWR.n1052 VPWR.n1051 34.7473
R3022 VPWR.n1299 VPWR.n1298 34.6358
R3023 VPWR.n1357 VPWR.n1341 34.6358
R3024 VPWR.n1362 VPWR.n1361 34.6358
R3025 VPWR.n1396 VPWR.n1380 34.6358
R3026 VPWR.n1401 VPWR.n1400 34.6358
R3027 VPWR.n1411 VPWR.n1377 34.6358
R3028 VPWR.n1433 VPWR.n1417 34.6358
R3029 VPWR.n1438 VPWR.n1437 34.6358
R3030 VPWR.n2755 VPWR.n2754 34.6358
R3031 VPWR.n2721 VPWR.n2713 34.6358
R3032 VPWR.n2728 VPWR.n2727 34.6358
R3033 VPWR.n2685 VPWR.n2676 34.6358
R3034 VPWR.n2688 VPWR.n2687 34.6358
R3035 VPWR.n2692 VPWR.n2691 34.6358
R3036 VPWR.n2648 VPWR.n2639 34.6358
R3037 VPWR.n2651 VPWR.n2650 34.6358
R3038 VPWR.n2655 VPWR.n2654 34.6358
R3039 VPWR.n2662 VPWR.n2661 34.6358
R3040 VPWR.n2615 VPWR.n2611 34.6358
R3041 VPWR.n2619 VPWR.n2603 34.6358
R3042 VPWR.n2622 VPWR.n2621 34.6358
R3043 VPWR.n1316 VPWR.n1315 32.0005
R3044 VPWR.n1353 VPWR.n1352 32.0005
R3045 VPWR.n1392 VPWR.n1391 32.0005
R3046 VPWR.n1429 VPWR.n1428 32.0005
R3047 VPWR.n2717 VPWR.n2716 30.8711
R3048 VPWR.n2681 VPWR.n2680 30.8711
R3049 VPWR.n2644 VPWR.n2643 30.8711
R3050 VPWR.n2610 VPWR.n2609 30.8711
R3051 VPWR.n2834 VPWR.n2832 30.1181
R3052 VPWR.n2838 VPWR.n2826 30.1181
R3053 VPWR.n2848 VPWR.n2846 28.9887
R3054 VPWR.n1325 VPWR.n1324 28.2358
R3055 VPWR.n5 VPWR.t717 26.5955
R3056 VPWR.n5 VPWR.t721 26.5955
R3057 VPWR.n4 VPWR.t440 26.5955
R3058 VPWR.n4 VPWR.t713 26.5955
R3059 VPWR.n1240 VPWR.t1769 26.5955
R3060 VPWR.n1240 VPWR.t1768 26.5955
R3061 VPWR.n1239 VPWR.t1828 26.5955
R3062 VPWR.n1239 VPWR.t611 26.5955
R3063 VPWR.n1245 VPWR.t1765 26.5955
R3064 VPWR.n1245 VPWR.t1770 26.5955
R3065 VPWR.n1238 VPWR.t694 26.5955
R3066 VPWR.n1238 VPWR.t1827 26.5955
R3067 VPWR.n1263 VPWR.t813 26.5955
R3068 VPWR.n1263 VPWR.t915 26.5955
R3069 VPWR.n1262 VPWR.t1683 26.5955
R3070 VPWR.n1262 VPWR.t1681 26.5955
R3071 VPWR.n1268 VPWR.t1925 26.5955
R3072 VPWR.n1268 VPWR.t102 26.5955
R3073 VPWR.n1261 VPWR.t1686 26.5955
R3074 VPWR.n1261 VPWR.t1684 26.5955
R3075 VPWR.n1287 VPWR.t617 26.5955
R3076 VPWR.n1287 VPWR.t624 26.5955
R3077 VPWR.n1286 VPWR.t965 26.5955
R3078 VPWR.n1286 VPWR.t964 26.5955
R3079 VPWR.n1292 VPWR.t621 26.5955
R3080 VPWR.n1292 VPWR.t618 26.5955
R3081 VPWR.n1285 VPWR.t968 26.5955
R3082 VPWR.n1285 VPWR.t966 26.5955
R3083 VPWR.n1314 VPWR.t372 26.5955
R3084 VPWR.n1314 VPWR.t374 26.5955
R3085 VPWR.n1307 VPWR.t719 26.5955
R3086 VPWR.n1307 VPWR.t370 26.5955
R3087 VPWR.n1321 VPWR.t715 26.5955
R3088 VPWR.n1321 VPWR.t438 26.5955
R3089 VPWR.n1323 VPWR.t382 26.5955
R3090 VPWR.n1323 VPWR.t609 26.5955
R3091 VPWR.n1351 VPWR.t45 26.5955
R3092 VPWR.n1351 VPWR.t1696 26.5955
R3093 VPWR.n1350 VPWR.t731 26.5955
R3094 VPWR.n1350 VPWR.t1891 26.5955
R3095 VPWR.n1344 VPWR.t1772 26.5955
R3096 VPWR.n1344 VPWR.t36 26.5955
R3097 VPWR.n1343 VPWR.t695 26.5955
R3098 VPWR.n1343 VPWR.t1693 26.5955
R3099 VPWR.n1359 VPWR.t1767 26.5955
R3100 VPWR.n1359 VPWR.t1766 26.5955
R3101 VPWR.n1358 VPWR.t612 26.5955
R3102 VPWR.n1358 VPWR.t696 26.5955
R3103 VPWR.n1390 VPWR.t1692 26.5955
R3104 VPWR.n1390 VPWR.t733 26.5955
R3105 VPWR.n1389 VPWR.t1695 26.5955
R3106 VPWR.n1389 VPWR.t607 26.5955
R3107 VPWR.n1383 VPWR.t17 26.5955
R3108 VPWR.n1383 VPWR.t1690 26.5955
R3109 VPWR.n1382 VPWR.t1687 26.5955
R3110 VPWR.n1382 VPWR.t41 26.5955
R3111 VPWR.n1398 VPWR.t916 26.5955
R3112 VPWR.n1398 VPWR.t1924 26.5955
R3113 VPWR.n1397 VPWR.t1688 26.5955
R3114 VPWR.n1397 VPWR.t1685 26.5955
R3115 VPWR.n1427 VPWR.t378 26.5955
R3116 VPWR.n1427 VPWR.t383 26.5955
R3117 VPWR.n1426 VPWR.t732 26.5955
R3118 VPWR.n1426 VPWR.t1892 26.5955
R3119 VPWR.n1420 VPWR.t620 26.5955
R3120 VPWR.n1420 VPWR.t1893 26.5955
R3121 VPWR.n1419 VPWR.t962 26.5955
R3122 VPWR.n1419 VPWR.t730 26.5955
R3123 VPWR.n1435 VPWR.t623 26.5955
R3124 VPWR.n1435 VPWR.t622 26.5955
R3125 VPWR.n1434 VPWR.t963 26.5955
R3126 VPWR.n1434 VPWR.t961 26.5955
R3127 VPWR.n2802 VPWR.t1071 26.5955
R3128 VPWR.n2802 VPWR.t1913 26.5955
R3129 VPWR.n2804 VPWR.t291 26.5955
R3130 VPWR.n2804 VPWR.t51 26.5955
R3131 VPWR.n2782 VPWR.t1020 26.5955
R3132 VPWR.n2782 VPWR.t1016 26.5955
R3133 VPWR.n2783 VPWR.t343 26.5955
R3134 VPWR.n2783 VPWR.t134 26.5955
R3135 VPWR.n2786 VPWR.t1012 26.5955
R3136 VPWR.n2786 VPWR.t1013 26.5955
R3137 VPWR.n2787 VPWR.t1559 26.5955
R3138 VPWR.n2787 VPWR.t549 26.5955
R3139 VPWR.n2762 VPWR.t1524 26.5955
R3140 VPWR.n2762 VPWR.t53 26.5955
R3141 VPWR.n2763 VPWR.t1779 26.5955
R3142 VPWR.n2763 VPWR.t1785 26.5955
R3143 VPWR.n2766 VPWR.t49 26.5955
R3144 VPWR.n2766 VPWR.t47 26.5955
R3145 VPWR.n2767 VPWR.t1781 26.5955
R3146 VPWR.n2767 VPWR.t1783 26.5955
R3147 VPWR.n2743 VPWR.t1903 26.5955
R3148 VPWR.n2743 VPWR.t1900 26.5955
R3149 VPWR.n2744 VPWR.t1615 26.5955
R3150 VPWR.n2744 VPWR.t1613 26.5955
R3151 VPWR.n2747 VPWR.t1904 26.5955
R3152 VPWR.n2747 VPWR.t1905 26.5955
R3153 VPWR.n2748 VPWR.t1619 26.5955
R3154 VPWR.n2748 VPWR.t1607 26.5955
R3155 VPWR.n2708 VPWR.t476 26.5955
R3156 VPWR.n2708 VPWR.t508 26.5955
R3157 VPWR.n2712 VPWR.t500 26.5955
R3158 VPWR.n2712 VPWR.t650 26.5955
R3159 VPWR.n2715 VPWR.t474 26.5955
R3160 VPWR.n2715 VPWR.t522 26.5955
R3161 VPWR.n2709 VPWR.t546 26.5955
R3162 VPWR.n2709 VPWR.t1067 26.5955
R3163 VPWR.n2679 VPWR.t470 26.5955
R3164 VPWR.n2679 VPWR.t520 26.5955
R3165 VPWR.n2678 VPWR.t486 26.5955
R3166 VPWR.n2678 VPWR.t532 26.5955
R3167 VPWR.n2675 VPWR.t497 26.5955
R3168 VPWR.n2675 VPWR.t414 26.5955
R3169 VPWR.n2674 VPWR.t514 26.5955
R3170 VPWR.n2674 VPWR.t1017 26.5955
R3171 VPWR.n2671 VPWR.t652 26.5955
R3172 VPWR.n2671 VPWR.t1662 26.5955
R3173 VPWR.n2670 VPWR.t1014 26.5955
R3174 VPWR.n2670 VPWR.t1019 26.5955
R3175 VPWR.n2642 VPWR.t492 26.5955
R3176 VPWR.n2642 VPWR.t466 26.5955
R3177 VPWR.n2641 VPWR.t510 26.5955
R3178 VPWR.n2641 VPWR.t485 26.5955
R3179 VPWR.n2638 VPWR.t518 26.5955
R3180 VPWR.n2638 VPWR.t1784 26.5955
R3181 VPWR.n2637 VPWR.t528 26.5955
R3182 VPWR.n2637 VPWR.t1528 26.5955
R3183 VPWR.n2634 VPWR.t1780 26.5955
R3184 VPWR.n2634 VPWR.t1786 26.5955
R3185 VPWR.n2633 VPWR.t57 26.5955
R3186 VPWR.n2633 VPWR.t1526 26.5955
R3187 VPWR.n2606 VPWR.t489 26.5955
R3188 VPWR.n2606 VPWR.t495 26.5955
R3189 VPWR.n2605 VPWR.t525 26.5955
R3190 VPWR.n2605 VPWR.t506 26.5955
R3191 VPWR.n2613 VPWR.t501 26.5955
R3192 VPWR.n2613 VPWR.t1617 26.5955
R3193 VPWR.n2612 VPWR.t483 26.5955
R3194 VPWR.n2612 VPWR.t1901 26.5955
R3195 VPWR.n2602 VPWR.t1621 26.5955
R3196 VPWR.n2602 VPWR.t1609 26.5955
R3197 VPWR.n2601 VPWR.t1898 26.5955
R3198 VPWR.n2601 VPWR.t1902 26.5955
R3199 VPWR.n17 VPWR.n16 25.977
R3200 VPWR.n1253 VPWR.n1252 25.977
R3201 VPWR.n1313 VPWR.n1310 25.977
R3202 VPWR.n1349 VPWR.n1346 25.977
R3203 VPWR.n1372 VPWR.n1338 25.977
R3204 VPWR.n1388 VPWR.n1385 25.977
R3205 VPWR.n1425 VPWR.n1422 25.977
R3206 VPWR.n2811 VPWR.n2810 25.977
R3207 VPWR.n2795 VPWR.n2794 25.977
R3208 VPWR.n2717 VPWR.n2714 25.977
R3209 VPWR.n2681 VPWR.n2677 25.977
R3210 VPWR.n2699 VPWR.n2698 25.977
R3211 VPWR.n2644 VPWR.n2640 25.977
R3212 VPWR.n2609 VPWR.n2607 25.977
R3213 VPWR.n1335 VPWR.n1334 25.224
R3214 VPWR.n2737 VPWR.n2736 25.224
R3215 VPWR.n2722 VPWR.n2721 24.8476
R3216 VPWR.n2686 VPWR.n2685 24.8476
R3217 VPWR.n2649 VPWR.n2648 24.8476
R3218 VPWR.n2615 VPWR.n2614 24.8476
R3219 VPWR.n16 VPWR.n15 24.4711
R3220 VPWR.n1252 VPWR.n1251 24.4711
R3221 VPWR.n1315 VPWR.n1313 24.4711
R3222 VPWR.n1352 VPWR.n1349 24.4711
R3223 VPWR.n1391 VPWR.n1388 24.4711
R3224 VPWR.n1428 VPWR.n1425 24.4711
R3225 VPWR.n2810 VPWR.n2809 24.4711
R3226 VPWR.n2794 VPWR.n2793 24.4711
R3227 VPWR.n11 VPWR.n2 23.7181
R3228 VPWR.n1247 VPWR.n1236 23.7181
R3229 VPWR.n1270 VPWR.n1259 23.7181
R3230 VPWR.n1274 VPWR.n1259 23.7181
R3231 VPWR.n1294 VPWR.n1283 23.7181
R3232 VPWR.n1298 VPWR.n1283 23.7181
R3233 VPWR.n1330 VPWR.n1328 23.7181
R3234 VPWR.n1368 VPWR.n1365 23.7181
R3235 VPWR.n1407 VPWR.n1404 23.7181
R3236 VPWR.n1407 VPWR.n1377 23.7181
R3237 VPWR.n1444 VPWR.n1441 23.7181
R3238 VPWR.n2808 VPWR.n2807 23.7181
R3239 VPWR.n2789 VPWR.n2781 23.7181
R3240 VPWR.n2769 VPWR.n2761 23.7181
R3241 VPWR.n2773 VPWR.n2761 23.7181
R3242 VPWR.n2750 VPWR.n2742 23.7181
R3243 VPWR.n2754 VPWR.n2742 23.7181
R3244 VPWR.n2731 VPWR.n2706 23.7181
R3245 VPWR.n2694 VPWR.n2668 23.7181
R3246 VPWR.n2657 VPWR.n2631 23.7181
R3247 VPWR.n2661 VPWR.n2631 23.7181
R3248 VPWR.n2626 VPWR.n2625 23.7181
R3249 VPWR.t839 VPWR.t1868 23.4987
R3250 VPWR.t543 VPWR.t613 23.4987
R3251 VPWR.n2852 VPWR.n2841 23.1255
R3252 VPWR.n2852 VPWR.t447 23.1255
R3253 VPWR.n2851 VPWR.n2819 23.1255
R3254 VPWR.t447 VPWR.n2851 23.1255
R3255 VPWR.n11 VPWR.n10 22.9652
R3256 VPWR.n1247 VPWR.n1246 22.9652
R3257 VPWR.n1270 VPWR.n1269 22.9652
R3258 VPWR.n1294 VPWR.n1293 22.9652
R3259 VPWR.n2807 VPWR.n2803 22.9652
R3260 VPWR.n2789 VPWR.n2788 22.9652
R3261 VPWR.n2769 VPWR.n2768 22.9652
R3262 VPWR.n2750 VPWR.n2749 22.9652
R3263 VPWR.n1320 VPWR.n1308 22.2123
R3264 VPWR.n2724 VPWR.n2723 22.2123
R3265 VPWR.n10 VPWR.n3 21.4593
R3266 VPWR.n1246 VPWR.n1237 21.4593
R3267 VPWR.n1269 VPWR.n1260 21.4593
R3268 VPWR.n1293 VPWR.n1284 21.4593
R3269 VPWR.n1442 VPWR.t42 20.5957
R3270 VPWR.n1443 VPWR.t377 20.5957
R3271 VPWR.n1277 VPWR.n1276 19.9534
R3272 VPWR.n1300 VPWR.n1299 19.9534
R3273 VPWR.n1334 VPWR.n1303 19.9534
R3274 VPWR.n2776 VPWR.n2775 19.9534
R3275 VPWR.n2756 VPWR.n2755 19.9534
R3276 VPWR.n2736 VPWR.n2735 19.9534
R3277 VPWR.n2724 VPWR.n2710 18.824
R3278 VPWR.n2688 VPWR.n2672 18.824
R3279 VPWR.n2651 VPWR.n2635 18.824
R3280 VPWR.n2620 VPWR.n2619 18.824
R3281 VPWR.n1316 VPWR.n1308 18.4476
R3282 VPWR.n1353 VPWR.n1345 18.4476
R3283 VPWR.n1373 VPWR.n1372 18.4476
R3284 VPWR.n1392 VPWR.n1384 18.4476
R3285 VPWR.n1429 VPWR.n1421 18.4476
R3286 VPWR.n2700 VPWR.n2699 18.4476
R3287 VPWR.n1413 VPWR.n1412 17.5829
R3288 VPWR.n2664 VPWR.n2663 17.5829
R3289 VPWR.n6 VPWR.n3 16.9417
R3290 VPWR.n1241 VPWR.n1237 16.9417
R3291 VPWR.n1264 VPWR.n1260 16.9417
R3292 VPWR.n1288 VPWR.n1284 16.9417
R3293 VPWR.n2730 VPWR.n2729 16.5652
R3294 VPWR.n1306 VPWR.n1304 16.1887
R3295 VPWR.n1374 VPWR.n1373 16.1887
R3296 VPWR.n2701 VPWR.n2700 16.1887
R3297 VPWR.n1235 VPWR.t32 16.0935
R3298 VPWR.n1258 VPWR.t44 16.0935
R3299 VPWR.n1282 VPWR.t104 16.0935
R3300 VPWR.n1367 VPWR.t35 16.0935
R3301 VPWR.n1406 VPWR.t16 16.0935
R3302 VPWR.n1234 VPWR.t109 16.0935
R3303 VPWR.n1257 VPWR.t34 16.0935
R3304 VPWR.n1281 VPWR.t108 16.0935
R3305 VPWR.n1366 VPWR.t38 16.0935
R3306 VPWR.n1405 VPWR.t40 16.0935
R3307 VPWR.n1325 VPWR.n1306 15.8123
R3308 VPWR.n2727 VPWR.n2710 15.8123
R3309 VPWR.n2729 VPWR.n2728 15.8123
R3310 VPWR.n2691 VPWR.n2672 15.8123
R3311 VPWR.n2654 VPWR.n2635 15.8123
R3312 VPWR.n2621 VPWR.n2620 15.8123
R3313 VPWR.n1330 VPWR.n1303 13.5534
R3314 VPWR.n2735 VPWR.n2706 13.5534
R3315 VPWR.n2839 VPWR.n2823 13.2148
R3316 VPWR.n2823 VPWR.t556 13.2148
R3317 VPWR.n2827 VPWR.n2817 13.2148
R3318 VPWR.n2827 VPWR.t556 13.2148
R3319 VPWR.n2833 VPWR.n2829 13.2148
R3320 VPWR.n2829 VPWR.t556 13.2148
R3321 VPWR.n15 VPWR.n2 12.8005
R3322 VPWR.n1251 VPWR.n1236 12.8005
R3323 VPWR.n1368 VPWR.n1338 12.8005
R3324 VPWR.n2809 VPWR.n2808 12.8005
R3325 VPWR.n2793 VPWR.n2781 12.8005
R3326 VPWR.n2698 VPWR.n2668 12.8005
R3327 VPWR.n1322 VPWR.n1320 12.424
R3328 VPWR.n1360 VPWR.n1357 12.424
R3329 VPWR.n1399 VPWR.n1396 12.424
R3330 VPWR.n1436 VPWR.n1433 12.424
R3331 VPWR.n1276 VPWR.n1275 10.5417
R3332 VPWR.n1412 VPWR.n1411 10.5417
R3333 VPWR.n2775 VPWR.n2774 10.5417
R3334 VPWR.n2663 VPWR.n2662 10.5417
R3335 VPWR.n2687 VPWR.n2686 9.78874
R3336 VPWR.n2650 VPWR.n2649 9.78874
R3337 VPWR.n2614 VPWR.n2603 9.78874
R3338 VPWR.n1361 VPWR.n1360 9.41227
R3339 VPWR.n1365 VPWR.n1339 9.41227
R3340 VPWR.n1400 VPWR.n1399 9.41227
R3341 VPWR.n1404 VPWR.n1378 9.41227
R3342 VPWR.n1437 VPWR.n1436 9.41227
R3343 VPWR.n1441 VPWR.n1415 9.41227
R3344 VPWR.n2694 VPWR.n2693 9.41227
R3345 VPWR.n2657 VPWR.n2656 9.41227
R3346 VPWR.n2625 VPWR.n2599 9.41227
R3347 VPWR.n1229 VPWR 9.37021
R3348 VPWR.n1151 VPWR 9.37021
R3349 VPWR.n1225 VPWR 9.37021
R3350 VPWR.n1483 VPWR 9.37021
R3351 VPWR.n1171 VPWR 9.37021
R3352 VPWR.n1167 VPWR 9.37021
R3353 VPWR.n1161 VPWR 9.37021
R3354 VPWR.n1477 VPWR 9.37021
R3355 VPWR.n1157 VPWR 9.37021
R3356 VPWR.n1147 VPWR 9.37021
R3357 VPWR.n1470 VPWR 9.37021
R3358 VPWR.n1047 VPWR 9.37021
R3359 VPWR.n1746 VPWR 9.37021
R3360 VPWR.n1034 VPWR 9.37021
R3361 VPWR.n1030 VPWR 9.37021
R3362 VPWR.n1051 VPWR 9.37021
R3363 VPWR.n1467 VPWR.n1466 9.33404
R3364 VPWR.n352 VPWR.n351 9.33404
R3365 VPWR.n1534 VPWR.n1533 9.33404
R3366 VPWR.n348 VPWR.n347 9.33404
R3367 VPWR.n965 VPWR.n964 9.33404
R3368 VPWR.n2479 VPWR.n2478 9.33404
R3369 VPWR.n2475 VPWR.n2474 9.33404
R3370 VPWR.n320 VPWR.n319 9.33404
R3371 VPWR.n973 VPWR.n972 9.33404
R3372 VPWR.n2445 VPWR.n2444 9.33404
R3373 VPWR.n324 VPWR.n323 9.33404
R3374 VPWR.n1891 VPWR.n1890 9.33404
R3375 VPWR.n1887 VPWR.n1886 9.33404
R3376 VPWR.n1881 VPWR.n1880 9.33404
R3377 VPWR.n389 VPWR.n388 9.33404
R3378 VPWR.n393 VPWR.n392 9.33404
R3379 VPWR.n397 VPWR.n396 9.33404
R3380 VPWR.n2455 VPWR.n2454 9.33404
R3381 VPWR.n332 VPWR.n331 9.33404
R3382 VPWR.n1877 VPWR.n1876 9.33404
R3383 VPWR.n405 VPWR.n404 9.33404
R3384 VPWR.n2459 VPWR.n2458 9.33404
R3385 VPWR.n336 VPWR.n335 9.33404
R3386 VPWR.n2308 VPWR.n2307 9.33404
R3387 VPWR.n2312 VPWR.n2311 9.33404
R3388 VPWR.n2318 VPWR.n2317 9.33404
R3389 VPWR.n2322 VPWR.n2321 9.33404
R3390 VPWR.n2332 VPWR.n2331 9.33404
R3391 VPWR.n2338 VPWR.n2337 9.33404
R3392 VPWR.n2342 VPWR.n2341 9.33404
R3393 VPWR.n2348 VPWR.n2347 9.33404
R3394 VPWR.n2352 VPWR.n2351 9.33404
R3395 VPWR.n2358 VPWR.n2357 9.33404
R3396 VPWR.n2362 VPWR.n2361 9.33404
R3397 VPWR.n2368 VPWR.n2367 9.33404
R3398 VPWR.n2372 VPWR.n2371 9.33404
R3399 VPWR.n2378 VPWR.n2377 9.33404
R3400 VPWR.n2381 VPWR.n2380 9.33404
R3401 VPWR.n2328 VPWR.n2327 9.33404
R3402 VPWR.n544 VPWR.n543 9.33404
R3403 VPWR.n540 VPWR.n539 9.33404
R3404 VPWR.n536 VPWR.n535 9.33404
R3405 VPWR.n532 VPWR.n531 9.33404
R3406 VPWR.n524 VPWR.n523 9.33404
R3407 VPWR.n520 VPWR.n519 9.33404
R3408 VPWR.n516 VPWR.n515 9.33404
R3409 VPWR.n512 VPWR.n511 9.33404
R3410 VPWR.n508 VPWR.n507 9.33404
R3411 VPWR.n504 VPWR.n503 9.33404
R3412 VPWR.n500 VPWR.n499 9.33404
R3413 VPWR.n496 VPWR.n495 9.33404
R3414 VPWR.n492 VPWR.n491 9.33404
R3415 VPWR.n488 VPWR.n487 9.33404
R3416 VPWR.n485 VPWR.n484 9.33404
R3417 VPWR.n528 VPWR.n527 9.33404
R3418 VPWR.n2283 VPWR.n2282 9.33404
R3419 VPWR.n2279 VPWR.n2278 9.33404
R3420 VPWR.n2273 VPWR.n2272 9.33404
R3421 VPWR.n2269 VPWR.n2268 9.33404
R3422 VPWR.n2259 VPWR.n2258 9.33404
R3423 VPWR.n2253 VPWR.n2252 9.33404
R3424 VPWR.n2249 VPWR.n2248 9.33404
R3425 VPWR.n2243 VPWR.n2242 9.33404
R3426 VPWR.n2239 VPWR.n2238 9.33404
R3427 VPWR.n2233 VPWR.n2232 9.33404
R3428 VPWR.n2229 VPWR.n2228 9.33404
R3429 VPWR.n2223 VPWR.n2222 9.33404
R3430 VPWR.n2219 VPWR.n2218 9.33404
R3431 VPWR.n2213 VPWR.n2212 9.33404
R3432 VPWR.n2210 VPWR.n2209 9.33404
R3433 VPWR.n2263 VPWR.n2262 9.33404
R3434 VPWR.n581 VPWR.n580 9.33404
R3435 VPWR.n585 VPWR.n584 9.33404
R3436 VPWR.n589 VPWR.n588 9.33404
R3437 VPWR.n593 VPWR.n592 9.33404
R3438 VPWR.n601 VPWR.n600 9.33404
R3439 VPWR.n605 VPWR.n604 9.33404
R3440 VPWR.n609 VPWR.n608 9.33404
R3441 VPWR.n613 VPWR.n612 9.33404
R3442 VPWR.n617 VPWR.n616 9.33404
R3443 VPWR.n621 VPWR.n620 9.33404
R3444 VPWR.n625 VPWR.n624 9.33404
R3445 VPWR.n629 VPWR.n628 9.33404
R3446 VPWR.n633 VPWR.n632 9.33404
R3447 VPWR.n637 VPWR.n636 9.33404
R3448 VPWR.n640 VPWR.n639 9.33404
R3449 VPWR.n597 VPWR.n596 9.33404
R3450 VPWR.n2112 VPWR.n2111 9.33404
R3451 VPWR.n2116 VPWR.n2115 9.33404
R3452 VPWR.n2122 VPWR.n2121 9.33404
R3453 VPWR.n2126 VPWR.n2125 9.33404
R3454 VPWR.n2136 VPWR.n2135 9.33404
R3455 VPWR.n2142 VPWR.n2141 9.33404
R3456 VPWR.n2146 VPWR.n2145 9.33404
R3457 VPWR.n2152 VPWR.n2151 9.33404
R3458 VPWR.n2156 VPWR.n2155 9.33404
R3459 VPWR.n2162 VPWR.n2161 9.33404
R3460 VPWR.n2166 VPWR.n2165 9.33404
R3461 VPWR.n2172 VPWR.n2171 9.33404
R3462 VPWR.n2176 VPWR.n2175 9.33404
R3463 VPWR.n2182 VPWR.n2181 9.33404
R3464 VPWR.n2185 VPWR.n2184 9.33404
R3465 VPWR.n2132 VPWR.n2131 9.33404
R3466 VPWR.n736 VPWR.n735 9.33404
R3467 VPWR.n732 VPWR.n731 9.33404
R3468 VPWR.n728 VPWR.n727 9.33404
R3469 VPWR.n724 VPWR.n723 9.33404
R3470 VPWR.n716 VPWR.n715 9.33404
R3471 VPWR.n712 VPWR.n711 9.33404
R3472 VPWR.n708 VPWR.n707 9.33404
R3473 VPWR.n704 VPWR.n703 9.33404
R3474 VPWR.n700 VPWR.n699 9.33404
R3475 VPWR.n696 VPWR.n695 9.33404
R3476 VPWR.n692 VPWR.n691 9.33404
R3477 VPWR.n688 VPWR.n687 9.33404
R3478 VPWR.n684 VPWR.n683 9.33404
R3479 VPWR.n680 VPWR.n679 9.33404
R3480 VPWR.n677 VPWR.n676 9.33404
R3481 VPWR.n720 VPWR.n719 9.33404
R3482 VPWR.n2087 VPWR.n2086 9.33404
R3483 VPWR.n2083 VPWR.n2082 9.33404
R3484 VPWR.n2077 VPWR.n2076 9.33404
R3485 VPWR.n2073 VPWR.n2072 9.33404
R3486 VPWR.n2063 VPWR.n2062 9.33404
R3487 VPWR.n2057 VPWR.n2056 9.33404
R3488 VPWR.n2053 VPWR.n2052 9.33404
R3489 VPWR.n2047 VPWR.n2046 9.33404
R3490 VPWR.n2043 VPWR.n2042 9.33404
R3491 VPWR.n2037 VPWR.n2036 9.33404
R3492 VPWR.n2033 VPWR.n2032 9.33404
R3493 VPWR.n2027 VPWR.n2026 9.33404
R3494 VPWR.n2023 VPWR.n2022 9.33404
R3495 VPWR.n2017 VPWR.n2016 9.33404
R3496 VPWR.n2014 VPWR.n2013 9.33404
R3497 VPWR.n2067 VPWR.n2066 9.33404
R3498 VPWR.n773 VPWR.n772 9.33404
R3499 VPWR.n777 VPWR.n776 9.33404
R3500 VPWR.n781 VPWR.n780 9.33404
R3501 VPWR.n785 VPWR.n784 9.33404
R3502 VPWR.n793 VPWR.n792 9.33404
R3503 VPWR.n797 VPWR.n796 9.33404
R3504 VPWR.n801 VPWR.n800 9.33404
R3505 VPWR.n805 VPWR.n804 9.33404
R3506 VPWR.n809 VPWR.n808 9.33404
R3507 VPWR.n813 VPWR.n812 9.33404
R3508 VPWR.n817 VPWR.n816 9.33404
R3509 VPWR.n821 VPWR.n820 9.33404
R3510 VPWR.n825 VPWR.n824 9.33404
R3511 VPWR.n829 VPWR.n828 9.33404
R3512 VPWR.n832 VPWR.n831 9.33404
R3513 VPWR.n789 VPWR.n788 9.33404
R3514 VPWR.n1916 VPWR.n1915 9.33404
R3515 VPWR.n1920 VPWR.n1919 9.33404
R3516 VPWR.n1926 VPWR.n1925 9.33404
R3517 VPWR.n1930 VPWR.n1929 9.33404
R3518 VPWR.n1940 VPWR.n1939 9.33404
R3519 VPWR.n1946 VPWR.n1945 9.33404
R3520 VPWR.n1950 VPWR.n1949 9.33404
R3521 VPWR.n1956 VPWR.n1955 9.33404
R3522 VPWR.n1960 VPWR.n1959 9.33404
R3523 VPWR.n1966 VPWR.n1965 9.33404
R3524 VPWR.n1970 VPWR.n1969 9.33404
R3525 VPWR.n1976 VPWR.n1975 9.33404
R3526 VPWR.n1980 VPWR.n1979 9.33404
R3527 VPWR.n1986 VPWR.n1985 9.33404
R3528 VPWR.n1989 VPWR.n1988 9.33404
R3529 VPWR.n1936 VPWR.n1935 9.33404
R3530 VPWR.n928 VPWR.n927 9.33404
R3531 VPWR.n924 VPWR.n923 9.33404
R3532 VPWR.n920 VPWR.n919 9.33404
R3533 VPWR.n916 VPWR.n915 9.33404
R3534 VPWR.n908 VPWR.n907 9.33404
R3535 VPWR.n904 VPWR.n903 9.33404
R3536 VPWR.n900 VPWR.n899 9.33404
R3537 VPWR.n896 VPWR.n895 9.33404
R3538 VPWR.n892 VPWR.n891 9.33404
R3539 VPWR.n888 VPWR.n887 9.33404
R3540 VPWR.n884 VPWR.n883 9.33404
R3541 VPWR.n880 VPWR.n879 9.33404
R3542 VPWR.n876 VPWR.n875 9.33404
R3543 VPWR.n872 VPWR.n871 9.33404
R3544 VPWR.n869 VPWR.n868 9.33404
R3545 VPWR.n912 VPWR.n911 9.33404
R3546 VPWR.n1871 VPWR.n1870 9.33404
R3547 VPWR.n981 VPWR.n980 9.33404
R3548 VPWR.n1495 VPWR.n1494 9.33404
R3549 VPWR.n401 VPWR.n400 9.33404
R3550 VPWR.n2465 VPWR.n2464 9.33404
R3551 VPWR.n340 VPWR.n339 9.33404
R3552 VPWR.n977 VPWR.n976 9.33404
R3553 VPWR.n1491 VPWR.n1490 9.33404
R3554 VPWR.n1867 VPWR.n1866 9.33404
R3555 VPWR.n985 VPWR.n984 9.33404
R3556 VPWR.n1505 VPWR.n1504 9.33404
R3557 VPWR.n409 VPWR.n408 9.33404
R3558 VPWR.n417 VPWR.n416 9.33404
R3559 VPWR.n421 VPWR.n420 9.33404
R3560 VPWR.n425 VPWR.n424 9.33404
R3561 VPWR.n429 VPWR.n428 9.33404
R3562 VPWR.n433 VPWR.n432 9.33404
R3563 VPWR.n437 VPWR.n436 9.33404
R3564 VPWR.n441 VPWR.n440 9.33404
R3565 VPWR.n445 VPWR.n444 9.33404
R3566 VPWR.n448 VPWR.n447 9.33404
R3567 VPWR.n413 VPWR.n412 9.33404
R3568 VPWR.n2449 VPWR.n2448 9.33404
R3569 VPWR.n328 VPWR.n327 9.33404
R3570 VPWR.n989 VPWR.n988 9.33404
R3571 VPWR.n1509 VPWR.n1508 9.33404
R3572 VPWR.n1861 VPWR.n1860 9.33404
R3573 VPWR.n1851 VPWR.n1850 9.33404
R3574 VPWR.n1847 VPWR.n1846 9.33404
R3575 VPWR.n1841 VPWR.n1840 9.33404
R3576 VPWR.n1837 VPWR.n1836 9.33404
R3577 VPWR.n1831 VPWR.n1830 9.33404
R3578 VPWR.n1827 VPWR.n1826 9.33404
R3579 VPWR.n1821 VPWR.n1820 9.33404
R3580 VPWR.n1818 VPWR.n1817 9.33404
R3581 VPWR.n1857 VPWR.n1856 9.33404
R3582 VPWR.n993 VPWR.n992 9.33404
R3583 VPWR.n1519 VPWR.n1518 9.33404
R3584 VPWR.n2469 VPWR.n2468 9.33404
R3585 VPWR.n344 VPWR.n343 9.33404
R3586 VPWR.n1480 VPWR.n1130 9.33404
R3587 VPWR.n997 VPWR.n996 9.33404
R3588 VPWR.n1523 VPWR.n1522 9.33404
R3589 VPWR.n2439 VPWR.n2438 9.33404
R3590 VPWR.n2429 VPWR.n2428 9.33404
R3591 VPWR.n2425 VPWR.n2424 9.33404
R3592 VPWR.n2419 VPWR.n2418 9.33404
R3593 VPWR.n2415 VPWR.n2414 9.33404
R3594 VPWR.n2409 VPWR.n2408 9.33404
R3595 VPWR.n2406 VPWR.n2405 9.33404
R3596 VPWR.n2435 VPWR.n2434 9.33404
R3597 VPWR.n316 VPWR.n315 9.33404
R3598 VPWR.n1538 VPWR.n1537 9.33404
R3599 VPWR.n1001 VPWR.n1000 9.33404
R3600 VPWR.n1005 VPWR.n1004 9.33404
R3601 VPWR.n1009 VPWR.n1008 9.33404
R3602 VPWR.n1013 VPWR.n1012 9.33404
R3603 VPWR.n1017 VPWR.n1016 9.33404
R3604 VPWR.n1021 VPWR.n1020 9.33404
R3605 VPWR.n1024 VPWR.n1023 9.33404
R3606 VPWR.n969 VPWR.n968 9.33404
R3607 VPWR.n1474 VPWR.n1473 9.33404
R3608 VPWR.n312 VPWR.n311 9.33404
R3609 VPWR.n1763 VPWR.n1762 9.33404
R3610 VPWR.n308 VPWR.n307 9.33404
R3611 VPWR.n304 VPWR.n303 9.33404
R3612 VPWR.n296 VPWR.n295 9.33404
R3613 VPWR.n293 VPWR.n292 9.33404
R3614 VPWR.n300 VPWR.n299 9.33404
R3615 VPWR.n1751 VPWR.n1750 9.33404
R3616 VPWR.n1790 VPWR.n1789 9.33404
R3617 VPWR.n1793 VPWR.n1792 9.33404
R3618 VPWR.n1759 VPWR.n1758 9.33404
R3619 VPWR.n2714 VPWR 9.32394
R3620 VPWR.n2677 VPWR 9.32394
R3621 VPWR.n2640 VPWR 9.32394
R3622 VPWR VPWR.n2607 9.32394
R3623 VPWR.n18 VPWR.n17 9.3005
R3624 VPWR.n15 VPWR.n14 9.3005
R3625 VPWR.n13 VPWR.n2 9.3005
R3626 VPWR.n10 VPWR.n9 9.3005
R3627 VPWR.n8 VPWR.n3 9.3005
R3628 VPWR.n12 VPWR.n11 9.3005
R3629 VPWR.n16 VPWR.n0 9.3005
R3630 VPWR.n1254 VPWR.n1253 9.3005
R3631 VPWR.n1251 VPWR.n1250 9.3005
R3632 VPWR.n1249 VPWR.n1236 9.3005
R3633 VPWR.n1246 VPWR.n1244 9.3005
R3634 VPWR.n1243 VPWR.n1237 9.3005
R3635 VPWR.n1248 VPWR.n1247 9.3005
R3636 VPWR.n1252 VPWR.n1233 9.3005
R3637 VPWR.n1278 VPWR.n1277 9.3005
R3638 VPWR.n1272 VPWR.n1259 9.3005
R3639 VPWR.n1269 VPWR.n1267 9.3005
R3640 VPWR.n1266 VPWR.n1260 9.3005
R3641 VPWR.n1271 VPWR.n1270 9.3005
R3642 VPWR.n1274 VPWR.n1273 9.3005
R3643 VPWR.n1276 VPWR.n1256 9.3005
R3644 VPWR.n1301 VPWR.n1300 9.3005
R3645 VPWR.n1296 VPWR.n1283 9.3005
R3646 VPWR.n1293 VPWR.n1291 9.3005
R3647 VPWR.n1290 VPWR.n1284 9.3005
R3648 VPWR.n1295 VPWR.n1294 9.3005
R3649 VPWR.n1298 VPWR.n1297 9.3005
R3650 VPWR.n1299 VPWR.n1280 9.3005
R3651 VPWR.n1332 VPWR.n1303 9.3005
R3652 VPWR.n1331 VPWR.n1330 9.3005
R3653 VPWR.n1311 VPWR.n1310 9.3005
R3654 VPWR.n1313 VPWR.n1312 9.3005
R3655 VPWR.n1315 VPWR.n1309 9.3005
R3656 VPWR.n1317 VPWR.n1316 9.3005
R3657 VPWR.n1318 VPWR.n1308 9.3005
R3658 VPWR.n1320 VPWR.n1319 9.3005
R3659 VPWR.n1324 VPWR.n1305 9.3005
R3660 VPWR.n1326 VPWR.n1325 9.3005
R3661 VPWR.n1328 VPWR.n1327 9.3005
R3662 VPWR.n1334 VPWR.n1333 9.3005
R3663 VPWR.n1336 VPWR.n1335 9.3005
R3664 VPWR.n1375 VPWR.n1374 9.3005
R3665 VPWR.n1370 VPWR.n1338 9.3005
R3666 VPWR.n1369 VPWR.n1368 9.3005
R3667 VPWR.n1347 VPWR.n1346 9.3005
R3668 VPWR.n1349 VPWR.n1348 9.3005
R3669 VPWR.n1352 VPWR.n1342 9.3005
R3670 VPWR.n1354 VPWR.n1353 9.3005
R3671 VPWR.n1355 VPWR.n1341 9.3005
R3672 VPWR.n1357 VPWR.n1356 9.3005
R3673 VPWR.n1361 VPWR.n1340 9.3005
R3674 VPWR.n1363 VPWR.n1362 9.3005
R3675 VPWR.n1365 VPWR.n1364 9.3005
R3676 VPWR.n1372 VPWR.n1371 9.3005
R3677 VPWR.n1408 VPWR.n1407 9.3005
R3678 VPWR.n1386 VPWR.n1385 9.3005
R3679 VPWR.n1388 VPWR.n1387 9.3005
R3680 VPWR.n1391 VPWR.n1381 9.3005
R3681 VPWR.n1393 VPWR.n1392 9.3005
R3682 VPWR.n1394 VPWR.n1380 9.3005
R3683 VPWR.n1396 VPWR.n1395 9.3005
R3684 VPWR.n1400 VPWR.n1379 9.3005
R3685 VPWR.n1402 VPWR.n1401 9.3005
R3686 VPWR.n1404 VPWR.n1403 9.3005
R3687 VPWR.n1409 VPWR.n1377 9.3005
R3688 VPWR.n1411 VPWR.n1410 9.3005
R3689 VPWR.n1445 VPWR.n1444 9.3005
R3690 VPWR.n1423 VPWR.n1422 9.3005
R3691 VPWR.n1425 VPWR.n1424 9.3005
R3692 VPWR.n1428 VPWR.n1418 9.3005
R3693 VPWR.n1430 VPWR.n1429 9.3005
R3694 VPWR.n1431 VPWR.n1417 9.3005
R3695 VPWR.n1433 VPWR.n1432 9.3005
R3696 VPWR.n1437 VPWR.n1416 9.3005
R3697 VPWR.n1439 VPWR.n1438 9.3005
R3698 VPWR.n1441 VPWR.n1440 9.3005
R3699 VPWR.n2807 VPWR.n2806 9.3005
R3700 VPWR.n2808 VPWR.n2800 9.3005
R3701 VPWR.n2809 VPWR.n2799 9.3005
R3702 VPWR.n2810 VPWR.n2798 9.3005
R3703 VPWR.n2812 VPWR.n2811 9.3005
R3704 VPWR.n2796 VPWR.n2795 9.3005
R3705 VPWR.n2790 VPWR.n2789 9.3005
R3706 VPWR.n2791 VPWR.n2781 9.3005
R3707 VPWR.n2793 VPWR.n2792 9.3005
R3708 VPWR.n2794 VPWR.n2779 9.3005
R3709 VPWR.n2777 VPWR.n2776 9.3005
R3710 VPWR.n2775 VPWR.n2759 9.3005
R3711 VPWR.n2770 VPWR.n2769 9.3005
R3712 VPWR.n2771 VPWR.n2761 9.3005
R3713 VPWR.n2773 VPWR.n2772 9.3005
R3714 VPWR.n2757 VPWR.n2756 9.3005
R3715 VPWR.n2751 VPWR.n2750 9.3005
R3716 VPWR.n2752 VPWR.n2742 9.3005
R3717 VPWR.n2754 VPWR.n2753 9.3005
R3718 VPWR.n2755 VPWR.n2740 9.3005
R3719 VPWR.n2738 VPWR.n2737 9.3005
R3720 VPWR.n2718 VPWR.n2717 9.3005
R3721 VPWR.n2719 VPWR.n2713 9.3005
R3722 VPWR.n2721 VPWR.n2720 9.3005
R3723 VPWR.n2723 VPWR.n2711 9.3005
R3724 VPWR.n2725 VPWR.n2724 9.3005
R3725 VPWR.n2727 VPWR.n2726 9.3005
R3726 VPWR.n2728 VPWR.n2707 9.3005
R3727 VPWR.n2732 VPWR.n2731 9.3005
R3728 VPWR.n2733 VPWR.n2706 9.3005
R3729 VPWR.n2735 VPWR.n2734 9.3005
R3730 VPWR.n2736 VPWR.n2704 9.3005
R3731 VPWR.n2702 VPWR.n2701 9.3005
R3732 VPWR.n2682 VPWR.n2681 9.3005
R3733 VPWR.n2683 VPWR.n2676 9.3005
R3734 VPWR.n2685 VPWR.n2684 9.3005
R3735 VPWR.n2687 VPWR.n2673 9.3005
R3736 VPWR.n2689 VPWR.n2688 9.3005
R3737 VPWR.n2691 VPWR.n2690 9.3005
R3738 VPWR.n2692 VPWR.n2669 9.3005
R3739 VPWR.n2695 VPWR.n2694 9.3005
R3740 VPWR.n2696 VPWR.n2668 9.3005
R3741 VPWR.n2698 VPWR.n2697 9.3005
R3742 VPWR.n2699 VPWR.n2666 9.3005
R3743 VPWR.n2645 VPWR.n2644 9.3005
R3744 VPWR.n2646 VPWR.n2639 9.3005
R3745 VPWR.n2648 VPWR.n2647 9.3005
R3746 VPWR.n2650 VPWR.n2636 9.3005
R3747 VPWR.n2652 VPWR.n2651 9.3005
R3748 VPWR.n2654 VPWR.n2653 9.3005
R3749 VPWR.n2655 VPWR.n2632 9.3005
R3750 VPWR.n2658 VPWR.n2657 9.3005
R3751 VPWR.n2659 VPWR.n2631 9.3005
R3752 VPWR.n2661 VPWR.n2660 9.3005
R3753 VPWR.n2662 VPWR.n2629 9.3005
R3754 VPWR.n2627 VPWR.n2626 9.3005
R3755 VPWR.n2609 VPWR.n2608 9.3005
R3756 VPWR.n2611 VPWR.n2604 9.3005
R3757 VPWR.n2616 VPWR.n2615 9.3005
R3758 VPWR.n2617 VPWR.n2603 9.3005
R3759 VPWR.n2619 VPWR.n2618 9.3005
R3760 VPWR.n2621 VPWR.n2600 9.3005
R3761 VPWR.n2623 VPWR.n2622 9.3005
R3762 VPWR.n2625 VPWR.n2624 9.3005
R3763 VPWR.n2505 VPWR.n2504 9.3005
R3764 VPWR.n2569 VPWR.n2568 9.3005
R3765 VPWR.n2509 VPWR.n2508 9.3005
R3766 VPWR.n2553 VPWR.n2552 9.3005
R3767 VPWR.n2545 VPWR.n2544 9.3005
R3768 VPWR.n2533 VPWR.n2532 9.3005
R3769 VPWR.n2529 VPWR.n2528 9.3005
R3770 VPWR.n1222 VPWR.n1221 9.3005
R3771 VPWR.n2521 VPWR.n2520 9.3005
R3772 VPWR.n1184 VPWR.n1102 9.3005
R3773 VPWR.n1218 VPWR.n1094 9.3005
R3774 VPWR.n2541 VPWR.n2540 9.3005
R3775 VPWR.n1215 VPWR.n1092 9.3005
R3776 VPWR.n1212 VPWR.n1211 9.3005
R3777 VPWR.n2517 VPWR.n2516 9.3005
R3778 VPWR.n1181 VPWR.n1104 9.3005
R3779 VPWR.n1204 VPWR.n1084 9.3005
R3780 VPWR.n2557 VPWR.n2556 9.3005
R3781 VPWR.n1201 VPWR.n1082 9.3005
R3782 VPWR.n1592 VPWR.n1591 9.3005
R3783 VPWR.n2565 VPWR.n2564 9.3005
R3784 VPWR.n1198 VPWR.n1197 9.3005
R3785 VPWR.n1190 VPWR.n1074 9.3005
R3786 VPWR.n1742 VPWR.n1741 9.3005
R3787 VPWR.n1187 VPWR.n1071 9.3005
R3788 VPWR.n2577 VPWR.n2576 9.3005
R3789 VPWR.n2581 VPWR.n2580 9.3005
R3790 VPWR.n2592 VPWR.n2591 9.3005
R3791 VPWR.n2589 VPWR.n2588 9.3005
R3792 VPWR.n1738 VPWR.n1737 9.3005
R3793 VPWR.n1063 VPWR.n1062 9.3005
R3794 VPWR.n1596 VPWR.n1595 9.3005
R3795 VPWR.n1275 VPWR.n1274 8.28285
R3796 VPWR.n2774 VPWR.n2773 8.28285
R3797 VPWR.n1607 VPWR.n1109 8.25914
R3798 VPWR.n1728 VPWR.n1727 8.25914
R3799 VPWR.n281 VPWR.n113 8.25914
R3800 VPWR.n136 VPWR.n124 8.25914
R3801 VPWR.n1780 VPWR.n1779 7.91351
R3802 VPWR.n1771 VPWR.n1770 7.9105
R3803 VPWR.n1042 VPWR.n1041 7.9105
R3804 VPWR.n1546 VPWR.n1545 7.9105
R3805 VPWR.n1551 VPWR.n1550 7.9105
R3806 VPWR.n1556 VPWR.n1555 7.9105
R3807 VPWR.n1561 VPWR.n1560 7.9105
R3808 VPWR.n1566 VPWR.n1565 7.9105
R3809 VPWR.n1571 VPWR.n1570 7.9105
R3810 VPWR.n1576 VPWR.n1575 7.9105
R3811 VPWR.n1581 VPWR.n1580 7.9105
R3812 VPWR.n1136 VPWR.n1135 7.9105
R3813 VPWR.n1461 VPWR.n1460 7.9105
R3814 VPWR.n1456 VPWR.n1455 7.9105
R3815 VPWR.n1776 VPWR.n1775 7.9105
R3816 VPWR.n1784 VPWR.n1783 7.9105
R3817 VPWR.n282 VPWR.n281 7.9105
R3818 VPWR.n280 VPWR.n279 7.9105
R3819 VPWR.n268 VPWR.n267 7.9105
R3820 VPWR.n256 VPWR.n255 7.9105
R3821 VPWR.n244 VPWR.n243 7.9105
R3822 VPWR.n232 VPWR.n231 7.9105
R3823 VPWR.n220 VPWR.n219 7.9105
R3824 VPWR.n208 VPWR.n207 7.9105
R3825 VPWR.n196 VPWR.n195 7.9105
R3826 VPWR.n184 VPWR.n183 7.9105
R3827 VPWR.n172 VPWR.n171 7.9105
R3828 VPWR.n160 VPWR.n159 7.9105
R3829 VPWR.n148 VPWR.n147 7.9105
R3830 VPWR.n136 VPWR.n135 7.9105
R3831 VPWR.n1727 VPWR.n1726 7.9105
R3832 VPWR.n1715 VPWR.n1714 7.9105
R3833 VPWR.n1701 VPWR.n1068 7.9105
R3834 VPWR.n1690 VPWR.n1689 7.9105
R3835 VPWR.n1688 VPWR.n1687 7.9105
R3836 VPWR.n1674 VPWR.n1079 7.9105
R3837 VPWR.n1663 VPWR.n1662 7.9105
R3838 VPWR.n1661 VPWR.n1660 7.9105
R3839 VPWR.n1647 VPWR.n1089 7.9105
R3840 VPWR.n1636 VPWR.n1635 7.9105
R3841 VPWR.n1634 VPWR.n1633 7.9105
R3842 VPWR.n1620 VPWR.n1099 7.9105
R3843 VPWR.n1609 VPWR.n1608 7.9105
R3844 VPWR.n1607 VPWR.n1606 7.9105
R3845 VPWR.n26 VPWR.n24 7.8627
R3846 VPWR.n7 VPWR.n6 7.56315
R3847 VPWR.n1242 VPWR.n1241 7.56315
R3848 VPWR.n1265 VPWR.n1264 7.56315
R3849 VPWR.n1289 VPWR.n1288 7.56315
R3850 VPWR.n2805 VPWR.n2803 6.4511
R3851 VPWR.n2788 VPWR.n2785 6.4511
R3852 VPWR.n2768 VPWR.n2765 6.4511
R3853 VPWR.n2749 VPWR.n2746 6.4511
R3854 VPWR.n1362 VPWR.n1339 6.4005
R3855 VPWR.n1401 VPWR.n1378 6.4005
R3856 VPWR.n1438 VPWR.n1415 6.4005
R3857 VPWR.n2723 VPWR.n2722 6.4005
R3858 VPWR.n2693 VPWR.n2692 6.4005
R3859 VPWR.n2656 VPWR.n2655 6.4005
R3860 VPWR.n2622 VPWR.n2599 6.4005
R3861 VPWR.n1595 VPWR.n1122 6.04494
R3862 VPWR.n2505 VPWR.n99 6.04494
R3863 VPWR.n1467 VPWR.n1231 6.04494
R3864 VPWR.n351 VPWR.n290 6.04494
R3865 VPWR.n2568 VPWR.n68 6.04494
R3866 VPWR.n1534 VPWR.n1153 6.04494
R3867 VPWR.n348 VPWR.n346 6.04494
R3868 VPWR.n2508 VPWR.n98 6.04494
R3869 VPWR.n965 VPWR.n963 6.04494
R3870 VPWR.n2478 VPWR.n356 6.04494
R3871 VPWR.n2475 VPWR.n357 6.04494
R3872 VPWR.n320 VPWR.n318 6.04494
R3873 VPWR.n2553 VPWR.n75 6.04494
R3874 VPWR.n973 VPWR.n971 6.04494
R3875 VPWR.n2445 VPWR.n369 6.04494
R3876 VPWR.n324 VPWR.n322 6.04494
R3877 VPWR.n2544 VPWR.n80 6.04494
R3878 VPWR.n1890 VPWR.n932 6.04494
R3879 VPWR.n1887 VPWR.n933 6.04494
R3880 VPWR.n1880 VPWR.n936 6.04494
R3881 VPWR.n389 VPWR.n387 6.04494
R3882 VPWR.n393 VPWR.n391 6.04494
R3883 VPWR.n397 VPWR.n395 6.04494
R3884 VPWR.n2455 VPWR.n365 6.04494
R3885 VPWR.n332 VPWR.n330 6.04494
R3886 VPWR.n2532 VPWR.n86 6.04494
R3887 VPWR.n1877 VPWR.n937 6.04494
R3888 VPWR.n405 VPWR.n403 6.04494
R3889 VPWR.n2458 VPWR.n364 6.04494
R3890 VPWR.n336 VPWR.n334 6.04494
R3891 VPWR.n2529 VPWR.n87 6.04494
R3892 VPWR.n2308 VPWR.n481 6.04494
R3893 VPWR.n2311 VPWR.n480 6.04494
R3894 VPWR.n2318 VPWR.n477 6.04494
R3895 VPWR.n2321 VPWR.n476 6.04494
R3896 VPWR.n2331 VPWR.n472 6.04494
R3897 VPWR.n2338 VPWR.n469 6.04494
R3898 VPWR.n2341 VPWR.n468 6.04494
R3899 VPWR.n2348 VPWR.n465 6.04494
R3900 VPWR.n2351 VPWR.n464 6.04494
R3901 VPWR.n2358 VPWR.n461 6.04494
R3902 VPWR.n2361 VPWR.n460 6.04494
R3903 VPWR.n2368 VPWR.n457 6.04494
R3904 VPWR.n2371 VPWR.n456 6.04494
R3905 VPWR.n2378 VPWR.n453 6.04494
R3906 VPWR.n2380 VPWR.n452 6.04494
R3907 VPWR.n2328 VPWR.n473 6.04494
R3908 VPWR.n543 VPWR.n482 6.04494
R3909 VPWR.n540 VPWR.n538 6.04494
R3910 VPWR.n536 VPWR.n534 6.04494
R3911 VPWR.n532 VPWR.n530 6.04494
R3912 VPWR.n524 VPWR.n522 6.04494
R3913 VPWR.n520 VPWR.n518 6.04494
R3914 VPWR.n516 VPWR.n514 6.04494
R3915 VPWR.n512 VPWR.n510 6.04494
R3916 VPWR.n508 VPWR.n506 6.04494
R3917 VPWR.n504 VPWR.n502 6.04494
R3918 VPWR.n500 VPWR.n498 6.04494
R3919 VPWR.n496 VPWR.n494 6.04494
R3920 VPWR.n492 VPWR.n490 6.04494
R3921 VPWR.n488 VPWR.n486 6.04494
R3922 VPWR.n485 VPWR.n483 6.04494
R3923 VPWR.n528 VPWR.n526 6.04494
R3924 VPWR.n2282 VPWR.n548 6.04494
R3925 VPWR.n2279 VPWR.n549 6.04494
R3926 VPWR.n2272 VPWR.n552 6.04494
R3927 VPWR.n2269 VPWR.n553 6.04494
R3928 VPWR.n2259 VPWR.n557 6.04494
R3929 VPWR.n2252 VPWR.n560 6.04494
R3930 VPWR.n2249 VPWR.n561 6.04494
R3931 VPWR.n2242 VPWR.n564 6.04494
R3932 VPWR.n2239 VPWR.n565 6.04494
R3933 VPWR.n2232 VPWR.n568 6.04494
R3934 VPWR.n2229 VPWR.n569 6.04494
R3935 VPWR.n2222 VPWR.n572 6.04494
R3936 VPWR.n2219 VPWR.n573 6.04494
R3937 VPWR.n2212 VPWR.n576 6.04494
R3938 VPWR.n2210 VPWR.n577 6.04494
R3939 VPWR.n2262 VPWR.n556 6.04494
R3940 VPWR.n581 VPWR.n579 6.04494
R3941 VPWR.n585 VPWR.n583 6.04494
R3942 VPWR.n589 VPWR.n587 6.04494
R3943 VPWR.n593 VPWR.n591 6.04494
R3944 VPWR.n601 VPWR.n599 6.04494
R3945 VPWR.n605 VPWR.n603 6.04494
R3946 VPWR.n609 VPWR.n607 6.04494
R3947 VPWR.n613 VPWR.n611 6.04494
R3948 VPWR.n617 VPWR.n615 6.04494
R3949 VPWR.n621 VPWR.n619 6.04494
R3950 VPWR.n625 VPWR.n623 6.04494
R3951 VPWR.n629 VPWR.n627 6.04494
R3952 VPWR.n633 VPWR.n631 6.04494
R3953 VPWR.n637 VPWR.n635 6.04494
R3954 VPWR.n639 VPWR.n578 6.04494
R3955 VPWR.n597 VPWR.n595 6.04494
R3956 VPWR.n2112 VPWR.n673 6.04494
R3957 VPWR.n2115 VPWR.n672 6.04494
R3958 VPWR.n2122 VPWR.n669 6.04494
R3959 VPWR.n2125 VPWR.n668 6.04494
R3960 VPWR.n2135 VPWR.n664 6.04494
R3961 VPWR.n2142 VPWR.n661 6.04494
R3962 VPWR.n2145 VPWR.n660 6.04494
R3963 VPWR.n2152 VPWR.n657 6.04494
R3964 VPWR.n2155 VPWR.n656 6.04494
R3965 VPWR.n2162 VPWR.n653 6.04494
R3966 VPWR.n2165 VPWR.n652 6.04494
R3967 VPWR.n2172 VPWR.n649 6.04494
R3968 VPWR.n2175 VPWR.n648 6.04494
R3969 VPWR.n2182 VPWR.n645 6.04494
R3970 VPWR.n2184 VPWR.n644 6.04494
R3971 VPWR.n2132 VPWR.n665 6.04494
R3972 VPWR.n735 VPWR.n674 6.04494
R3973 VPWR.n732 VPWR.n730 6.04494
R3974 VPWR.n728 VPWR.n726 6.04494
R3975 VPWR.n724 VPWR.n722 6.04494
R3976 VPWR.n716 VPWR.n714 6.04494
R3977 VPWR.n712 VPWR.n710 6.04494
R3978 VPWR.n708 VPWR.n706 6.04494
R3979 VPWR.n704 VPWR.n702 6.04494
R3980 VPWR.n700 VPWR.n698 6.04494
R3981 VPWR.n696 VPWR.n694 6.04494
R3982 VPWR.n692 VPWR.n690 6.04494
R3983 VPWR.n688 VPWR.n686 6.04494
R3984 VPWR.n684 VPWR.n682 6.04494
R3985 VPWR.n680 VPWR.n678 6.04494
R3986 VPWR.n677 VPWR.n675 6.04494
R3987 VPWR.n720 VPWR.n718 6.04494
R3988 VPWR.n2086 VPWR.n740 6.04494
R3989 VPWR.n2083 VPWR.n741 6.04494
R3990 VPWR.n2076 VPWR.n744 6.04494
R3991 VPWR.n2073 VPWR.n745 6.04494
R3992 VPWR.n2063 VPWR.n749 6.04494
R3993 VPWR.n2056 VPWR.n752 6.04494
R3994 VPWR.n2053 VPWR.n753 6.04494
R3995 VPWR.n2046 VPWR.n756 6.04494
R3996 VPWR.n2043 VPWR.n757 6.04494
R3997 VPWR.n2036 VPWR.n760 6.04494
R3998 VPWR.n2033 VPWR.n761 6.04494
R3999 VPWR.n2026 VPWR.n764 6.04494
R4000 VPWR.n2023 VPWR.n765 6.04494
R4001 VPWR.n2016 VPWR.n768 6.04494
R4002 VPWR.n2014 VPWR.n769 6.04494
R4003 VPWR.n2066 VPWR.n748 6.04494
R4004 VPWR.n773 VPWR.n771 6.04494
R4005 VPWR.n777 VPWR.n775 6.04494
R4006 VPWR.n781 VPWR.n779 6.04494
R4007 VPWR.n785 VPWR.n783 6.04494
R4008 VPWR.n793 VPWR.n791 6.04494
R4009 VPWR.n797 VPWR.n795 6.04494
R4010 VPWR.n801 VPWR.n799 6.04494
R4011 VPWR.n805 VPWR.n803 6.04494
R4012 VPWR.n809 VPWR.n807 6.04494
R4013 VPWR.n813 VPWR.n811 6.04494
R4014 VPWR.n817 VPWR.n815 6.04494
R4015 VPWR.n821 VPWR.n819 6.04494
R4016 VPWR.n825 VPWR.n823 6.04494
R4017 VPWR.n829 VPWR.n827 6.04494
R4018 VPWR.n831 VPWR.n770 6.04494
R4019 VPWR.n789 VPWR.n787 6.04494
R4020 VPWR.n1916 VPWR.n865 6.04494
R4021 VPWR.n1919 VPWR.n864 6.04494
R4022 VPWR.n1926 VPWR.n861 6.04494
R4023 VPWR.n1929 VPWR.n860 6.04494
R4024 VPWR.n1939 VPWR.n856 6.04494
R4025 VPWR.n1946 VPWR.n853 6.04494
R4026 VPWR.n1949 VPWR.n852 6.04494
R4027 VPWR.n1956 VPWR.n849 6.04494
R4028 VPWR.n1959 VPWR.n848 6.04494
R4029 VPWR.n1966 VPWR.n845 6.04494
R4030 VPWR.n1969 VPWR.n844 6.04494
R4031 VPWR.n1976 VPWR.n841 6.04494
R4032 VPWR.n1979 VPWR.n840 6.04494
R4033 VPWR.n1986 VPWR.n837 6.04494
R4034 VPWR.n1988 VPWR.n836 6.04494
R4035 VPWR.n1936 VPWR.n857 6.04494
R4036 VPWR.n927 VPWR.n866 6.04494
R4037 VPWR.n924 VPWR.n922 6.04494
R4038 VPWR.n920 VPWR.n918 6.04494
R4039 VPWR.n916 VPWR.n914 6.04494
R4040 VPWR.n908 VPWR.n906 6.04494
R4041 VPWR.n904 VPWR.n902 6.04494
R4042 VPWR.n900 VPWR.n898 6.04494
R4043 VPWR.n896 VPWR.n894 6.04494
R4044 VPWR.n892 VPWR.n890 6.04494
R4045 VPWR.n888 VPWR.n886 6.04494
R4046 VPWR.n884 VPWR.n882 6.04494
R4047 VPWR.n880 VPWR.n878 6.04494
R4048 VPWR.n876 VPWR.n874 6.04494
R4049 VPWR.n872 VPWR.n870 6.04494
R4050 VPWR.n869 VPWR.n867 6.04494
R4051 VPWR.n912 VPWR.n910 6.04494
R4052 VPWR.n1870 VPWR.n940 6.04494
R4053 VPWR.n981 VPWR.n979 6.04494
R4054 VPWR.n1494 VPWR.n1227 6.04494
R4055 VPWR.n1221 VPWR.n1179 6.04494
R4056 VPWR.n401 VPWR.n399 6.04494
R4057 VPWR.n2465 VPWR.n361 6.04494
R4058 VPWR.n340 VPWR.n338 6.04494
R4059 VPWR.n2520 VPWR.n92 6.04494
R4060 VPWR.n977 VPWR.n975 6.04494
R4061 VPWR.n1491 VPWR.n1485 6.04494
R4062 VPWR.n1184 VPWR.n1183 6.04494
R4063 VPWR.n1867 VPWR.n941 6.04494
R4064 VPWR.n985 VPWR.n983 6.04494
R4065 VPWR.n1505 VPWR.n1173 6.04494
R4066 VPWR.n1218 VPWR.n1217 6.04494
R4067 VPWR.n409 VPWR.n407 6.04494
R4068 VPWR.n417 VPWR.n415 6.04494
R4069 VPWR.n421 VPWR.n419 6.04494
R4070 VPWR.n425 VPWR.n423 6.04494
R4071 VPWR.n429 VPWR.n427 6.04494
R4072 VPWR.n433 VPWR.n431 6.04494
R4073 VPWR.n437 VPWR.n435 6.04494
R4074 VPWR.n441 VPWR.n439 6.04494
R4075 VPWR.n445 VPWR.n443 6.04494
R4076 VPWR.n447 VPWR.n386 6.04494
R4077 VPWR.n413 VPWR.n411 6.04494
R4078 VPWR.n2448 VPWR.n368 6.04494
R4079 VPWR.n328 VPWR.n326 6.04494
R4080 VPWR.n2541 VPWR.n81 6.04494
R4081 VPWR.n989 VPWR.n987 6.04494
R4082 VPWR.n1508 VPWR.n1169 6.04494
R4083 VPWR.n1215 VPWR.n1214 6.04494
R4084 VPWR.n1860 VPWR.n944 6.04494
R4085 VPWR.n1850 VPWR.n948 6.04494
R4086 VPWR.n1847 VPWR.n949 6.04494
R4087 VPWR.n1840 VPWR.n952 6.04494
R4088 VPWR.n1837 VPWR.n953 6.04494
R4089 VPWR.n1830 VPWR.n956 6.04494
R4090 VPWR.n1827 VPWR.n957 6.04494
R4091 VPWR.n1820 VPWR.n960 6.04494
R4092 VPWR.n1818 VPWR.n961 6.04494
R4093 VPWR.n1857 VPWR.n945 6.04494
R4094 VPWR.n993 VPWR.n991 6.04494
R4095 VPWR.n1519 VPWR.n1163 6.04494
R4096 VPWR.n1212 VPWR.n1206 6.04494
R4097 VPWR.n2468 VPWR.n360 6.04494
R4098 VPWR.n344 VPWR.n342 6.04494
R4099 VPWR.n2517 VPWR.n93 6.04494
R4100 VPWR.n1480 VPWR.n1479 6.04494
R4101 VPWR.n1181 VPWR.n1180 6.04494
R4102 VPWR.n997 VPWR.n995 6.04494
R4103 VPWR.n1522 VPWR.n1159 6.04494
R4104 VPWR.n1204 VPWR.n1203 6.04494
R4105 VPWR.n2438 VPWR.n372 6.04494
R4106 VPWR.n2428 VPWR.n376 6.04494
R4107 VPWR.n2425 VPWR.n377 6.04494
R4108 VPWR.n2418 VPWR.n380 6.04494
R4109 VPWR.n2415 VPWR.n381 6.04494
R4110 VPWR.n2408 VPWR.n384 6.04494
R4111 VPWR.n2406 VPWR.n385 6.04494
R4112 VPWR.n2435 VPWR.n373 6.04494
R4113 VPWR.n316 VPWR.n314 6.04494
R4114 VPWR.n2556 VPWR.n74 6.04494
R4115 VPWR.n1537 VPWR.n1149 6.04494
R4116 VPWR.n1201 VPWR.n1200 6.04494
R4117 VPWR.n1001 VPWR.n999 6.04494
R4118 VPWR.n1005 VPWR.n1003 6.04494
R4119 VPWR.n1009 VPWR.n1007 6.04494
R4120 VPWR.n1013 VPWR.n1011 6.04494
R4121 VPWR.n1017 VPWR.n1015 6.04494
R4122 VPWR.n1021 VPWR.n1019 6.04494
R4123 VPWR.n1023 VPWR.n962 6.04494
R4124 VPWR.n969 VPWR.n967 6.04494
R4125 VPWR.n1474 VPWR.n1472 6.04494
R4126 VPWR.n1592 VPWR.n1123 6.04494
R4127 VPWR.n312 VPWR.n310 6.04494
R4128 VPWR.n2565 VPWR.n69 6.04494
R4129 VPWR.n1198 VPWR.n1192 6.04494
R4130 VPWR.n1762 VPWR.n1049 6.04494
R4131 VPWR.n1190 VPWR.n1189 6.04494
R4132 VPWR.n308 VPWR.n306 6.04494
R4133 VPWR.n304 VPWR.n302 6.04494
R4134 VPWR.n296 VPWR.n294 6.04494
R4135 VPWR.n293 VPWR.n291 6.04494
R4136 VPWR.n300 VPWR.n298 6.04494
R4137 VPWR.n1741 VPWR.n1058 6.04494
R4138 VPWR.n1750 VPWR.n1748 6.04494
R4139 VPWR.n1790 VPWR.n1036 6.04494
R4140 VPWR.n1792 VPWR.n1032 6.04494
R4141 VPWR.n1759 VPWR.n1053 6.04494
R4142 VPWR.n1187 VPWR.n1186 6.04494
R4143 VPWR.n2577 VPWR.n63 6.04494
R4144 VPWR.n2580 VPWR.n62 6.04494
R4145 VPWR.n2589 VPWR.n57 6.04494
R4146 VPWR.n2591 VPWR.n56 6.04494
R4147 VPWR.n1738 VPWR.n1059 6.04494
R4148 VPWR.n1062 VPWR.n1061 6.04494
R4149 VPWR.n2785 VPWR.n2784 5.39628
R4150 VPWR.n2765 VPWR.n2764 5.39628
R4151 VPWR.n2746 VPWR.n2745 5.39628
R4152 VPWR.n54 VPWR 4.72593
R4153 VPWR.n52 VPWR 4.72593
R4154 VPWR.n50 VPWR 4.72593
R4155 VPWR.n48 VPWR 4.72593
R4156 VPWR.n46 VPWR 4.72593
R4157 VPWR.n44 VPWR 4.72593
R4158 VPWR.n42 VPWR 4.72593
R4159 VPWR.n40 VPWR 4.72593
R4160 VPWR.n38 VPWR 4.72593
R4161 VPWR.n36 VPWR 4.72593
R4162 VPWR.n34 VPWR 4.72593
R4163 VPWR.n32 VPWR 4.72593
R4164 VPWR.n30 VPWR 4.72593
R4165 VPWR.n28 VPWR 4.72593
R4166 VPWR.n26 VPWR 4.72593
R4167 VPWR.n1446 VPWR.n1445 4.55954
R4168 VPWR.n2571 VPWR.n2570 4.5005
R4169 VPWR.n2511 VPWR.n2510 4.5005
R4170 VPWR.n2551 VPWR.n2550 4.5005
R4171 VPWR.n319 VPWR.n77 4.5005
R4172 VPWR.n2547 VPWR.n2546 4.5005
R4173 VPWR.n323 VPWR.n78 4.5005
R4174 VPWR.n2535 VPWR.n2534 4.5005
R4175 VPWR.n331 VPWR.n84 4.5005
R4176 VPWR.n2454 VPWR.n2453 4.5005
R4177 VPWR.n2527 VPWR.n2526 4.5005
R4178 VPWR.n335 VPWR.n89 4.5005
R4179 VPWR.n2460 VPWR.n2459 4.5005
R4180 VPWR.n1498 VPWR.n1223 4.5005
R4181 VPWR.n1497 VPWR.n1495 4.5005
R4182 VPWR.n980 VPWR.n939 4.5005
R4183 VPWR.n1872 VPWR.n1871 4.5005
R4184 VPWR.n911 VPWR.n858 4.5005
R4185 VPWR.n1935 VPWR.n1934 4.5005
R4186 VPWR.n788 VPWR.n747 4.5005
R4187 VPWR.n2068 VPWR.n2067 4.5005
R4188 VPWR.n719 VPWR.n666 4.5005
R4189 VPWR.n2131 VPWR.n2130 4.5005
R4190 VPWR.n596 VPWR.n555 4.5005
R4191 VPWR.n2264 VPWR.n2263 4.5005
R4192 VPWR.n527 VPWR.n474 4.5005
R4193 VPWR.n2327 VPWR.n2326 4.5005
R4194 VPWR.n404 VPWR.n363 4.5005
R4195 VPWR.n2523 VPWR.n2522 4.5005
R4196 VPWR.n339 VPWR.n90 4.5005
R4197 VPWR.n2464 VPWR.n2463 4.5005
R4198 VPWR.n400 VPWR.n362 4.5005
R4199 VPWR.n2323 VPWR.n2322 4.5005
R4200 VPWR.n531 VPWR.n475 4.5005
R4201 VPWR.n2268 VPWR.n2267 4.5005
R4202 VPWR.n592 VPWR.n554 4.5005
R4203 VPWR.n2127 VPWR.n2126 4.5005
R4204 VPWR.n723 VPWR.n667 4.5005
R4205 VPWR.n2072 VPWR.n2071 4.5005
R4206 VPWR.n784 VPWR.n746 4.5005
R4207 VPWR.n1931 VPWR.n1930 4.5005
R4208 VPWR.n915 VPWR.n859 4.5005
R4209 VPWR.n1488 VPWR.n1486 4.5005
R4210 VPWR.n1490 VPWR.n1489 4.5005
R4211 VPWR.n976 VPWR.n938 4.5005
R4212 VPWR.n1876 VPWR.n1875 4.5005
R4213 VPWR.n1501 VPWR.n1174 4.5005
R4214 VPWR.n1504 VPWR.n1503 4.5005
R4215 VPWR.n984 VPWR.n942 4.5005
R4216 VPWR.n1866 VPWR.n1865 4.5005
R4217 VPWR.n907 VPWR.n855 4.5005
R4218 VPWR.n1941 VPWR.n1940 4.5005
R4219 VPWR.n792 VPWR.n750 4.5005
R4220 VPWR.n2062 VPWR.n2061 4.5005
R4221 VPWR.n715 VPWR.n663 4.5005
R4222 VPWR.n2137 VPWR.n2136 4.5005
R4223 VPWR.n600 VPWR.n558 4.5005
R4224 VPWR.n2258 VPWR.n2257 4.5005
R4225 VPWR.n523 VPWR.n471 4.5005
R4226 VPWR.n2333 VPWR.n2332 4.5005
R4227 VPWR.n408 VPWR.n366 4.5005
R4228 VPWR.n2539 VPWR.n2538 4.5005
R4229 VPWR.n327 VPWR.n83 4.5005
R4230 VPWR.n2450 VPWR.n2449 4.5005
R4231 VPWR.n412 VPWR.n367 4.5005
R4232 VPWR.n2337 VPWR.n2336 4.5005
R4233 VPWR.n519 VPWR.n470 4.5005
R4234 VPWR.n2254 VPWR.n2253 4.5005
R4235 VPWR.n604 VPWR.n559 4.5005
R4236 VPWR.n2141 VPWR.n2140 4.5005
R4237 VPWR.n711 VPWR.n662 4.5005
R4238 VPWR.n2058 VPWR.n2057 4.5005
R4239 VPWR.n796 VPWR.n751 4.5005
R4240 VPWR.n1945 VPWR.n1944 4.5005
R4241 VPWR.n903 VPWR.n854 4.5005
R4242 VPWR.n1512 VPWR.n1165 4.5005
R4243 VPWR.n1511 VPWR.n1509 4.5005
R4244 VPWR.n988 VPWR.n943 4.5005
R4245 VPWR.n1862 VPWR.n1861 4.5005
R4246 VPWR.n1515 VPWR.n1164 4.5005
R4247 VPWR.n1518 VPWR.n1517 4.5005
R4248 VPWR.n992 VPWR.n946 4.5005
R4249 VPWR.n1856 VPWR.n1855 4.5005
R4250 VPWR.n899 VPWR.n851 4.5005
R4251 VPWR.n1951 VPWR.n1950 4.5005
R4252 VPWR.n800 VPWR.n754 4.5005
R4253 VPWR.n2052 VPWR.n2051 4.5005
R4254 VPWR.n707 VPWR.n659 4.5005
R4255 VPWR.n2147 VPWR.n2146 4.5005
R4256 VPWR.n608 VPWR.n562 4.5005
R4257 VPWR.n2248 VPWR.n2247 4.5005
R4258 VPWR.n515 VPWR.n467 4.5005
R4259 VPWR.n2343 VPWR.n2342 4.5005
R4260 VPWR.n416 VPWR.n370 4.5005
R4261 VPWR.n2444 VPWR.n2443 4.5005
R4262 VPWR.n2515 VPWR.n2514 4.5005
R4263 VPWR.n343 VPWR.n95 4.5005
R4264 VPWR.n2470 VPWR.n2469 4.5005
R4265 VPWR.n396 VPWR.n359 4.5005
R4266 VPWR.n2317 VPWR.n2316 4.5005
R4267 VPWR.n535 VPWR.n478 4.5005
R4268 VPWR.n2274 VPWR.n2273 4.5005
R4269 VPWR.n588 VPWR.n551 4.5005
R4270 VPWR.n2121 VPWR.n2120 4.5005
R4271 VPWR.n727 VPWR.n670 4.5005
R4272 VPWR.n2078 VPWR.n2077 4.5005
R4273 VPWR.n780 VPWR.n743 4.5005
R4274 VPWR.n1925 VPWR.n1924 4.5005
R4275 VPWR.n919 VPWR.n862 4.5005
R4276 VPWR.n1882 VPWR.n1881 4.5005
R4277 VPWR.n1586 VPWR.n1129 4.5005
R4278 VPWR.n1585 VPWR.n1130 4.5005
R4279 VPWR.n972 VPWR.n935 4.5005
R4280 VPWR.n1526 VPWR.n1155 4.5005
R4281 VPWR.n1525 VPWR.n1523 4.5005
R4282 VPWR.n996 VPWR.n947 4.5005
R4283 VPWR.n1852 VPWR.n1851 4.5005
R4284 VPWR.n895 VPWR.n850 4.5005
R4285 VPWR.n1955 VPWR.n1954 4.5005
R4286 VPWR.n804 VPWR.n755 4.5005
R4287 VPWR.n2048 VPWR.n2047 4.5005
R4288 VPWR.n703 VPWR.n658 4.5005
R4289 VPWR.n2151 VPWR.n2150 4.5005
R4290 VPWR.n612 VPWR.n563 4.5005
R4291 VPWR.n2244 VPWR.n2243 4.5005
R4292 VPWR.n511 VPWR.n466 4.5005
R4293 VPWR.n2347 VPWR.n2346 4.5005
R4294 VPWR.n420 VPWR.n371 4.5005
R4295 VPWR.n2440 VPWR.n2439 4.5005
R4296 VPWR.n2559 VPWR.n2558 4.5005
R4297 VPWR.n315 VPWR.n72 4.5005
R4298 VPWR.n2434 VPWR.n2433 4.5005
R4299 VPWR.n424 VPWR.n374 4.5005
R4300 VPWR.n2353 VPWR.n2352 4.5005
R4301 VPWR.n507 VPWR.n463 4.5005
R4302 VPWR.n2238 VPWR.n2237 4.5005
R4303 VPWR.n616 VPWR.n566 4.5005
R4304 VPWR.n2157 VPWR.n2156 4.5005
R4305 VPWR.n699 VPWR.n655 4.5005
R4306 VPWR.n2042 VPWR.n2041 4.5005
R4307 VPWR.n808 VPWR.n758 4.5005
R4308 VPWR.n1961 VPWR.n1960 4.5005
R4309 VPWR.n891 VPWR.n847 4.5005
R4310 VPWR.n1846 VPWR.n1845 4.5005
R4311 VPWR.n1145 VPWR.n1144 4.5005
R4312 VPWR.n1539 VPWR.n1538 4.5005
R4313 VPWR.n1000 VPWR.n950 4.5005
R4314 VPWR.n1590 VPWR.n1589 4.5005
R4315 VPWR.n1473 VPWR.n1128 4.5005
R4316 VPWR.n968 VPWR.n934 4.5005
R4317 VPWR.n1886 VPWR.n1885 4.5005
R4318 VPWR.n923 VPWR.n863 4.5005
R4319 VPWR.n1921 VPWR.n1920 4.5005
R4320 VPWR.n776 VPWR.n742 4.5005
R4321 VPWR.n2082 VPWR.n2081 4.5005
R4322 VPWR.n731 VPWR.n671 4.5005
R4323 VPWR.n2117 VPWR.n2116 4.5005
R4324 VPWR.n584 VPWR.n550 4.5005
R4325 VPWR.n2278 VPWR.n2277 4.5005
R4326 VPWR.n539 VPWR.n479 4.5005
R4327 VPWR.n2313 VPWR.n2312 4.5005
R4328 VPWR.n392 VPWR.n358 4.5005
R4329 VPWR.n2474 VPWR.n2473 4.5005
R4330 VPWR.n347 VPWR.n96 4.5005
R4331 VPWR.n2563 VPWR.n2562 4.5005
R4332 VPWR.n311 VPWR.n71 4.5005
R4333 VPWR.n2430 VPWR.n2429 4.5005
R4334 VPWR.n428 VPWR.n375 4.5005
R4335 VPWR.n2357 VPWR.n2356 4.5005
R4336 VPWR.n503 VPWR.n462 4.5005
R4337 VPWR.n2234 VPWR.n2233 4.5005
R4338 VPWR.n620 VPWR.n567 4.5005
R4339 VPWR.n2161 VPWR.n2160 4.5005
R4340 VPWR.n695 VPWR.n654 4.5005
R4341 VPWR.n2038 VPWR.n2037 4.5005
R4342 VPWR.n812 VPWR.n759 4.5005
R4343 VPWR.n1965 VPWR.n1964 4.5005
R4344 VPWR.n887 VPWR.n846 4.5005
R4345 VPWR.n1842 VPWR.n1841 4.5005
R4346 VPWR.n1004 VPWR.n951 4.5005
R4347 VPWR.n1531 VPWR.n1154 4.5005
R4348 VPWR.n1533 VPWR.n1532 4.5005
R4349 VPWR.n1073 VPWR.n1045 4.5005
R4350 VPWR.n1764 VPWR.n1763 4.5005
R4351 VPWR.n1008 VPWR.n954 4.5005
R4352 VPWR.n1836 VPWR.n1835 4.5005
R4353 VPWR.n883 VPWR.n843 4.5005
R4354 VPWR.n1971 VPWR.n1970 4.5005
R4355 VPWR.n816 VPWR.n762 4.5005
R4356 VPWR.n2032 VPWR.n2031 4.5005
R4357 VPWR.n691 VPWR.n651 4.5005
R4358 VPWR.n2167 VPWR.n2166 4.5005
R4359 VPWR.n624 VPWR.n570 4.5005
R4360 VPWR.n2228 VPWR.n2227 4.5005
R4361 VPWR.n499 VPWR.n459 4.5005
R4362 VPWR.n2363 VPWR.n2362 4.5005
R4363 VPWR.n432 VPWR.n378 4.5005
R4364 VPWR.n2424 VPWR.n2423 4.5005
R4365 VPWR.n307 VPWR.n66 4.5005
R4366 VPWR.n299 VPWR.n60 4.5005
R4367 VPWR.n2414 VPWR.n2413 4.5005
R4368 VPWR.n440 VPWR.n382 4.5005
R4369 VPWR.n2373 VPWR.n2372 4.5005
R4370 VPWR.n491 VPWR.n455 4.5005
R4371 VPWR.n2218 VPWR.n2217 4.5005
R4372 VPWR.n632 VPWR.n574 4.5005
R4373 VPWR.n2177 VPWR.n2176 4.5005
R4374 VPWR.n683 VPWR.n647 4.5005
R4375 VPWR.n2022 VPWR.n2021 4.5005
R4376 VPWR.n824 VPWR.n766 4.5005
R4377 VPWR.n1981 VPWR.n1980 4.5005
R4378 VPWR.n875 VPWR.n839 4.5005
R4379 VPWR.n1826 VPWR.n1825 4.5005
R4380 VPWR.n1016 VPWR.n958 4.5005
R4381 VPWR.n1753 VPWR.n1743 4.5005
R4382 VPWR.n1752 VPWR.n1751 4.5005
R4383 VPWR.n1756 VPWR.n1054 4.5005
R4384 VPWR.n1758 VPWR.n1757 4.5005
R4385 VPWR.n1012 VPWR.n955 4.5005
R4386 VPWR.n1832 VPWR.n1831 4.5005
R4387 VPWR.n879 VPWR.n842 4.5005
R4388 VPWR.n1975 VPWR.n1974 4.5005
R4389 VPWR.n820 VPWR.n763 4.5005
R4390 VPWR.n2028 VPWR.n2027 4.5005
R4391 VPWR.n687 VPWR.n650 4.5005
R4392 VPWR.n2171 VPWR.n2170 4.5005
R4393 VPWR.n628 VPWR.n571 4.5005
R4394 VPWR.n2224 VPWR.n2223 4.5005
R4395 VPWR.n495 VPWR.n458 4.5005
R4396 VPWR.n2367 VPWR.n2366 4.5005
R4397 VPWR.n436 VPWR.n379 4.5005
R4398 VPWR.n2420 VPWR.n2419 4.5005
R4399 VPWR.n303 VPWR.n65 4.5005
R4400 VPWR.n2575 VPWR.n2574 4.5005
R4401 VPWR.n2583 VPWR.n2582 4.5005
R4402 VPWR.n2587 VPWR.n2586 4.5005
R4403 VPWR.n295 VPWR.n59 4.5005
R4404 VPWR.n2410 VPWR.n2409 4.5005
R4405 VPWR.n444 VPWR.n383 4.5005
R4406 VPWR.n2377 VPWR.n2376 4.5005
R4407 VPWR.n487 VPWR.n454 4.5005
R4408 VPWR.n2214 VPWR.n2213 4.5005
R4409 VPWR.n636 VPWR.n575 4.5005
R4410 VPWR.n2181 VPWR.n2180 4.5005
R4411 VPWR.n679 VPWR.n646 4.5005
R4412 VPWR.n2018 VPWR.n2017 4.5005
R4413 VPWR.n828 VPWR.n767 4.5005
R4414 VPWR.n1985 VPWR.n1984 4.5005
R4415 VPWR.n871 VPWR.n838 4.5005
R4416 VPWR.n1822 VPWR.n1821 4.5005
R4417 VPWR.n1020 VPWR.n959 4.5005
R4418 VPWR.n1789 VPWR.n1788 4.5005
R4419 VPWR.n1736 VPWR.n1037 4.5005
R4420 VPWR.n1232 VPWR.n1121 4.5005
R4421 VPWR.n1466 VPWR.n1465 4.5005
R4422 VPWR.n964 VPWR.n931 4.5005
R4423 VPWR.n1892 VPWR.n1891 4.5005
R4424 VPWR.n929 VPWR.n928 4.5005
R4425 VPWR.n1915 VPWR.n1914 4.5005
R4426 VPWR.n772 VPWR.n739 4.5005
R4427 VPWR.n2088 VPWR.n2087 4.5005
R4428 VPWR.n737 VPWR.n736 4.5005
R4429 VPWR.n2111 VPWR.n2110 4.5005
R4430 VPWR.n580 VPWR.n547 4.5005
R4431 VPWR.n2284 VPWR.n2283 4.5005
R4432 VPWR.n545 VPWR.n544 4.5005
R4433 VPWR.n2307 VPWR.n2306 4.5005
R4434 VPWR.n388 VPWR.n355 4.5005
R4435 VPWR.n2480 VPWR.n2479 4.5005
R4436 VPWR.n353 VPWR.n352 4.5005
R4437 VPWR.n2503 VPWR.n2502 4.5005
R4438 VPWR.n2594 VPWR.n2593 4.5005
R4439 VPWR.n292 VPWR.n22 4.5005
R4440 VPWR.n2405 VPWR.n2404 4.5005
R4441 VPWR.n449 VPWR.n448 4.5005
R4442 VPWR.n2382 VPWR.n2381 4.5005
R4443 VPWR.n484 VPWR.n451 4.5005
R4444 VPWR.n2209 VPWR.n2208 4.5005
R4445 VPWR.n641 VPWR.n640 4.5005
R4446 VPWR.n2186 VPWR.n2185 4.5005
R4447 VPWR.n676 VPWR.n643 4.5005
R4448 VPWR.n2013 VPWR.n2012 4.5005
R4449 VPWR.n833 VPWR.n832 4.5005
R4450 VPWR.n1990 VPWR.n1989 4.5005
R4451 VPWR.n868 VPWR.n835 4.5005
R4452 VPWR.n1817 VPWR.n1816 4.5005
R4453 VPWR.n1025 VPWR.n1024 4.5005
R4454 VPWR.n1794 VPWR.n1793 4.5005
R4455 VPWR.n1060 VPWR.n1028 4.5005
R4456 VPWR.n2628 VPWR 4.49965
R4457 VPWR.n19 VPWR.n18 4.20017
R4458 VPWR.n1255 VPWR.n1254 4.20017
R4459 VPWR.n1279 VPWR.n1278 4.20017
R4460 VPWR.n1302 VPWR.n1301 4.20017
R4461 VPWR.n1337 VPWR.n1336 4.20017
R4462 VPWR.n1376 VPWR.n1375 4.20017
R4463 VPWR.n1414 VPWR.n1413 4.20017
R4464 VPWR.n2813 VPWR 4.14027
R4465 VPWR.n2797 VPWR 4.14027
R4466 VPWR.n2778 VPWR 4.14027
R4467 VPWR.n2758 VPWR 4.14027
R4468 VPWR.n2739 VPWR 4.14027
R4469 VPWR.n2703 VPWR 4.14027
R4470 VPWR.n2665 VPWR 4.14027
R4471 VPWR.n55 VPWR.n54 4.0005
R4472 VPWR.n2716 VPWR.n2713 3.76521
R4473 VPWR.n2680 VPWR.n2676 3.76521
R4474 VPWR.n2643 VPWR.n2639 3.76521
R4475 VPWR.n2611 VPWR.n2610 3.76521
R4476 VPWR.n1906 VPWR.n858 3.4105
R4477 VPWR.n1934 VPWR.n1933 3.4105
R4478 VPWR.n1997 VPWR.n747 3.4105
R4479 VPWR.n2069 VPWR.n2068 3.4105
R4480 VPWR.n2102 VPWR.n666 3.4105
R4481 VPWR.n2130 VPWR.n2129 3.4105
R4482 VPWR.n2193 VPWR.n555 3.4105
R4483 VPWR.n2265 VPWR.n2264 3.4105
R4484 VPWR.n2298 VPWR.n474 3.4105
R4485 VPWR.n2326 VPWR.n2325 3.4105
R4486 VPWR.n2389 VPWR.n363 3.4105
R4487 VPWR.n2388 VPWR.n362 3.4105
R4488 VPWR.n2324 VPWR.n2323 3.4105
R4489 VPWR.n2299 VPWR.n475 3.4105
R4490 VPWR.n2267 VPWR.n2266 3.4105
R4491 VPWR.n2192 VPWR.n554 3.4105
R4492 VPWR.n2128 VPWR.n2127 3.4105
R4493 VPWR.n2103 VPWR.n667 3.4105
R4494 VPWR.n2071 VPWR.n2070 3.4105
R4495 VPWR.n1996 VPWR.n746 3.4105
R4496 VPWR.n1932 VPWR.n1931 3.4105
R4497 VPWR.n1907 VPWR.n859 3.4105
R4498 VPWR.n1875 VPWR.n1874 3.4105
R4499 VPWR.n1873 VPWR.n1872 3.4105
R4500 VPWR.n1865 VPWR.n1864 3.4105
R4501 VPWR.n1905 VPWR.n855 3.4105
R4502 VPWR.n1942 VPWR.n1941 3.4105
R4503 VPWR.n1998 VPWR.n750 3.4105
R4504 VPWR.n2061 VPWR.n2060 3.4105
R4505 VPWR.n2101 VPWR.n663 3.4105
R4506 VPWR.n2138 VPWR.n2137 3.4105
R4507 VPWR.n2194 VPWR.n558 3.4105
R4508 VPWR.n2257 VPWR.n2256 3.4105
R4509 VPWR.n2297 VPWR.n471 3.4105
R4510 VPWR.n2334 VPWR.n2333 3.4105
R4511 VPWR.n2390 VPWR.n366 3.4105
R4512 VPWR.n2391 VPWR.n367 3.4105
R4513 VPWR.n2336 VPWR.n2335 3.4105
R4514 VPWR.n2296 VPWR.n470 3.4105
R4515 VPWR.n2255 VPWR.n2254 3.4105
R4516 VPWR.n2195 VPWR.n559 3.4105
R4517 VPWR.n2140 VPWR.n2139 3.4105
R4518 VPWR.n2100 VPWR.n662 3.4105
R4519 VPWR.n2059 VPWR.n2058 3.4105
R4520 VPWR.n1999 VPWR.n751 3.4105
R4521 VPWR.n1944 VPWR.n1943 3.4105
R4522 VPWR.n1904 VPWR.n854 3.4105
R4523 VPWR.n1863 VPWR.n1862 3.4105
R4524 VPWR.n1855 VPWR.n1854 3.4105
R4525 VPWR.n1903 VPWR.n851 3.4105
R4526 VPWR.n1952 VPWR.n1951 3.4105
R4527 VPWR.n2000 VPWR.n754 3.4105
R4528 VPWR.n2051 VPWR.n2050 3.4105
R4529 VPWR.n2099 VPWR.n659 3.4105
R4530 VPWR.n2148 VPWR.n2147 3.4105
R4531 VPWR.n2196 VPWR.n562 3.4105
R4532 VPWR.n2247 VPWR.n2246 3.4105
R4533 VPWR.n2295 VPWR.n467 3.4105
R4534 VPWR.n2344 VPWR.n2343 3.4105
R4535 VPWR.n2392 VPWR.n370 3.4105
R4536 VPWR.n2443 VPWR.n2442 3.4105
R4537 VPWR.n2451 VPWR.n2450 3.4105
R4538 VPWR.n2453 VPWR.n2452 3.4105
R4539 VPWR.n2461 VPWR.n2460 3.4105
R4540 VPWR.n2463 VPWR.n2462 3.4105
R4541 VPWR.n2471 VPWR.n2470 3.4105
R4542 VPWR.n2387 VPWR.n359 3.4105
R4543 VPWR.n2316 VPWR.n2315 3.4105
R4544 VPWR.n2300 VPWR.n478 3.4105
R4545 VPWR.n2275 VPWR.n2274 3.4105
R4546 VPWR.n2191 VPWR.n551 3.4105
R4547 VPWR.n2120 VPWR.n2119 3.4105
R4548 VPWR.n2104 VPWR.n670 3.4105
R4549 VPWR.n2079 VPWR.n2078 3.4105
R4550 VPWR.n1995 VPWR.n743 3.4105
R4551 VPWR.n1924 VPWR.n1923 3.4105
R4552 VPWR.n1908 VPWR.n862 3.4105
R4553 VPWR.n1883 VPWR.n1882 3.4105
R4554 VPWR.n1799 VPWR.n935 3.4105
R4555 VPWR.n1800 VPWR.n938 3.4105
R4556 VPWR.n1801 VPWR.n939 3.4105
R4557 VPWR.n1802 VPWR.n942 3.4105
R4558 VPWR.n1803 VPWR.n943 3.4105
R4559 VPWR.n1804 VPWR.n946 3.4105
R4560 VPWR.n1805 VPWR.n947 3.4105
R4561 VPWR.n1853 VPWR.n1852 3.4105
R4562 VPWR.n1902 VPWR.n850 3.4105
R4563 VPWR.n1954 VPWR.n1953 3.4105
R4564 VPWR.n2001 VPWR.n755 3.4105
R4565 VPWR.n2049 VPWR.n2048 3.4105
R4566 VPWR.n2098 VPWR.n658 3.4105
R4567 VPWR.n2150 VPWR.n2149 3.4105
R4568 VPWR.n2197 VPWR.n563 3.4105
R4569 VPWR.n2245 VPWR.n2244 3.4105
R4570 VPWR.n2294 VPWR.n466 3.4105
R4571 VPWR.n2346 VPWR.n2345 3.4105
R4572 VPWR.n2393 VPWR.n371 3.4105
R4573 VPWR.n2441 VPWR.n2440 3.4105
R4574 VPWR.n2433 VPWR.n2432 3.4105
R4575 VPWR.n2394 VPWR.n374 3.4105
R4576 VPWR.n2354 VPWR.n2353 3.4105
R4577 VPWR.n2293 VPWR.n463 3.4105
R4578 VPWR.n2237 VPWR.n2236 3.4105
R4579 VPWR.n2198 VPWR.n566 3.4105
R4580 VPWR.n2158 VPWR.n2157 3.4105
R4581 VPWR.n2097 VPWR.n655 3.4105
R4582 VPWR.n2041 VPWR.n2040 3.4105
R4583 VPWR.n2002 VPWR.n758 3.4105
R4584 VPWR.n1962 VPWR.n1961 3.4105
R4585 VPWR.n1901 VPWR.n847 3.4105
R4586 VPWR.n1845 VPWR.n1844 3.4105
R4587 VPWR.n1806 VPWR.n950 3.4105
R4588 VPWR.n1798 VPWR.n934 3.4105
R4589 VPWR.n1885 VPWR.n1884 3.4105
R4590 VPWR.n1909 VPWR.n863 3.4105
R4591 VPWR.n1922 VPWR.n1921 3.4105
R4592 VPWR.n1994 VPWR.n742 3.4105
R4593 VPWR.n2081 VPWR.n2080 3.4105
R4594 VPWR.n2105 VPWR.n671 3.4105
R4595 VPWR.n2118 VPWR.n2117 3.4105
R4596 VPWR.n2190 VPWR.n550 3.4105
R4597 VPWR.n2277 VPWR.n2276 3.4105
R4598 VPWR.n2301 VPWR.n479 3.4105
R4599 VPWR.n2314 VPWR.n2313 3.4105
R4600 VPWR.n2386 VPWR.n358 3.4105
R4601 VPWR.n2473 VPWR.n2472 3.4105
R4602 VPWR.n2497 VPWR.n96 3.4105
R4603 VPWR.n2496 VPWR.n95 3.4105
R4604 VPWR.n2495 VPWR.n90 3.4105
R4605 VPWR.n2494 VPWR.n89 3.4105
R4606 VPWR.n2493 VPWR.n84 3.4105
R4607 VPWR.n2492 VPWR.n83 3.4105
R4608 VPWR.n2491 VPWR.n78 3.4105
R4609 VPWR.n2490 VPWR.n77 3.4105
R4610 VPWR.n2489 VPWR.n72 3.4105
R4611 VPWR.n2488 VPWR.n71 3.4105
R4612 VPWR.n2431 VPWR.n2430 3.4105
R4613 VPWR.n2395 VPWR.n375 3.4105
R4614 VPWR.n2356 VPWR.n2355 3.4105
R4615 VPWR.n2292 VPWR.n462 3.4105
R4616 VPWR.n2235 VPWR.n2234 3.4105
R4617 VPWR.n2199 VPWR.n567 3.4105
R4618 VPWR.n2160 VPWR.n2159 3.4105
R4619 VPWR.n2096 VPWR.n654 3.4105
R4620 VPWR.n2039 VPWR.n2038 3.4105
R4621 VPWR.n2003 VPWR.n759 3.4105
R4622 VPWR.n1964 VPWR.n1963 3.4105
R4623 VPWR.n1900 VPWR.n846 3.4105
R4624 VPWR.n1843 VPWR.n1842 3.4105
R4625 VPWR.n1807 VPWR.n951 3.4105
R4626 VPWR.n1532 VPWR.n1143 3.4105
R4627 VPWR.n1540 VPWR.n1539 3.4105
R4628 VPWR.n1525 VPWR.n1524 3.4105
R4629 VPWR.n1517 VPWR.n1516 3.4105
R4630 VPWR.n1511 VPWR.n1510 3.4105
R4631 VPWR.n1503 VPWR.n1502 3.4105
R4632 VPWR.n1497 VPWR.n1496 3.4105
R4633 VPWR.n1489 VPWR.n1132 3.4105
R4634 VPWR.n1585 VPWR.n1584 3.4105
R4635 VPWR.n1452 VPWR.n1128 3.4105
R4636 VPWR.n1765 VPWR.n1764 3.4105
R4637 VPWR.n1808 VPWR.n954 3.4105
R4638 VPWR.n1835 VPWR.n1834 3.4105
R4639 VPWR.n1899 VPWR.n843 3.4105
R4640 VPWR.n1972 VPWR.n1971 3.4105
R4641 VPWR.n2004 VPWR.n762 3.4105
R4642 VPWR.n2031 VPWR.n2030 3.4105
R4643 VPWR.n2095 VPWR.n651 3.4105
R4644 VPWR.n2168 VPWR.n2167 3.4105
R4645 VPWR.n2200 VPWR.n570 3.4105
R4646 VPWR.n2227 VPWR.n2226 3.4105
R4647 VPWR.n2291 VPWR.n459 3.4105
R4648 VPWR.n2364 VPWR.n2363 3.4105
R4649 VPWR.n2396 VPWR.n378 3.4105
R4650 VPWR.n2423 VPWR.n2422 3.4105
R4651 VPWR.n2487 VPWR.n66 3.4105
R4652 VPWR.n2485 VPWR.n60 3.4105
R4653 VPWR.n2413 VPWR.n2412 3.4105
R4654 VPWR.n2398 VPWR.n382 3.4105
R4655 VPWR.n2374 VPWR.n2373 3.4105
R4656 VPWR.n2289 VPWR.n455 3.4105
R4657 VPWR.n2217 VPWR.n2216 3.4105
R4658 VPWR.n2202 VPWR.n574 3.4105
R4659 VPWR.n2178 VPWR.n2177 3.4105
R4660 VPWR.n2093 VPWR.n647 3.4105
R4661 VPWR.n2021 VPWR.n2020 3.4105
R4662 VPWR.n2006 VPWR.n766 3.4105
R4663 VPWR.n1982 VPWR.n1981 3.4105
R4664 VPWR.n1897 VPWR.n839 3.4105
R4665 VPWR.n1825 VPWR.n1824 3.4105
R4666 VPWR.n1810 VPWR.n958 3.4105
R4667 VPWR.n1752 VPWR.n1744 3.4105
R4668 VPWR.n1757 VPWR.n1043 3.4105
R4669 VPWR.n1809 VPWR.n955 3.4105
R4670 VPWR.n1833 VPWR.n1832 3.4105
R4671 VPWR.n1898 VPWR.n842 3.4105
R4672 VPWR.n1974 VPWR.n1973 3.4105
R4673 VPWR.n2005 VPWR.n763 3.4105
R4674 VPWR.n2029 VPWR.n2028 3.4105
R4675 VPWR.n2094 VPWR.n650 3.4105
R4676 VPWR.n2170 VPWR.n2169 3.4105
R4677 VPWR.n2201 VPWR.n571 3.4105
R4678 VPWR.n2225 VPWR.n2224 3.4105
R4679 VPWR.n2290 VPWR.n458 3.4105
R4680 VPWR.n2366 VPWR.n2365 3.4105
R4681 VPWR.n2397 VPWR.n379 3.4105
R4682 VPWR.n2421 VPWR.n2420 3.4105
R4683 VPWR.n2486 VPWR.n65 3.4105
R4684 VPWR.n2484 VPWR.n59 3.4105
R4685 VPWR.n2411 VPWR.n2410 3.4105
R4686 VPWR.n2399 VPWR.n383 3.4105
R4687 VPWR.n2376 VPWR.n2375 3.4105
R4688 VPWR.n2288 VPWR.n454 3.4105
R4689 VPWR.n2215 VPWR.n2214 3.4105
R4690 VPWR.n2203 VPWR.n575 3.4105
R4691 VPWR.n2180 VPWR.n2179 3.4105
R4692 VPWR.n2092 VPWR.n646 3.4105
R4693 VPWR.n2019 VPWR.n2018 3.4105
R4694 VPWR.n2007 VPWR.n767 3.4105
R4695 VPWR.n1984 VPWR.n1983 3.4105
R4696 VPWR.n1896 VPWR.n838 3.4105
R4697 VPWR.n1823 VPWR.n1822 3.4105
R4698 VPWR.n1811 VPWR.n959 3.4105
R4699 VPWR.n1788 VPWR.n1787 3.4105
R4700 VPWR.n1465 VPWR.n1464 3.4105
R4701 VPWR.n1797 VPWR.n931 3.4105
R4702 VPWR.n1893 VPWR.n1892 3.4105
R4703 VPWR.n1910 VPWR.n929 3.4105
R4704 VPWR.n1914 VPWR.n1913 3.4105
R4705 VPWR.n1993 VPWR.n739 3.4105
R4706 VPWR.n2089 VPWR.n2088 3.4105
R4707 VPWR.n2106 VPWR.n737 3.4105
R4708 VPWR.n2110 VPWR.n2109 3.4105
R4709 VPWR.n2189 VPWR.n547 3.4105
R4710 VPWR.n2285 VPWR.n2284 3.4105
R4711 VPWR.n2302 VPWR.n545 3.4105
R4712 VPWR.n2306 VPWR.n2305 3.4105
R4713 VPWR.n2385 VPWR.n355 3.4105
R4714 VPWR.n2481 VPWR.n2480 3.4105
R4715 VPWR.n2498 VPWR.n353 3.4105
R4716 VPWR.n2502 VPWR.n2501 3.4105
R4717 VPWR.n2512 VPWR.n2511 3.4105
R4718 VPWR.n2514 VPWR.n2513 3.4105
R4719 VPWR.n2524 VPWR.n2523 3.4105
R4720 VPWR.n2526 VPWR.n2525 3.4105
R4721 VPWR.n2536 VPWR.n2535 3.4105
R4722 VPWR.n2538 VPWR.n2537 3.4105
R4723 VPWR.n2548 VPWR.n2547 3.4105
R4724 VPWR.n2550 VPWR.n2549 3.4105
R4725 VPWR.n2560 VPWR.n2559 3.4105
R4726 VPWR.n2562 VPWR.n2561 3.4105
R4727 VPWR.n2572 VPWR.n2571 3.4105
R4728 VPWR.n2574 VPWR.n2573 3.4105
R4729 VPWR.n2584 VPWR.n2583 3.4105
R4730 VPWR.n2586 VPWR.n2585 3.4105
R4731 VPWR.n2595 VPWR.n2594 3.4105
R4732 VPWR.n2483 VPWR.n22 3.4105
R4733 VPWR.n2404 VPWR.n2403 3.4105
R4734 VPWR.n2400 VPWR.n449 3.4105
R4735 VPWR.n2383 VPWR.n2382 3.4105
R4736 VPWR.n2287 VPWR.n451 3.4105
R4737 VPWR.n2208 VPWR.n2207 3.4105
R4738 VPWR.n2204 VPWR.n641 3.4105
R4739 VPWR.n2187 VPWR.n2186 3.4105
R4740 VPWR.n2091 VPWR.n643 3.4105
R4741 VPWR.n2012 VPWR.n2011 3.4105
R4742 VPWR.n2008 VPWR.n833 3.4105
R4743 VPWR.n1991 VPWR.n1990 3.4105
R4744 VPWR.n1895 VPWR.n835 3.4105
R4745 VPWR.n1816 VPWR.n1815 3.4105
R4746 VPWR.n1812 VPWR.n1025 3.4105
R4747 VPWR.n1795 VPWR.n1794 3.4105
R4748 VPWR.n1055 VPWR.n1028 3.4105
R4749 VPWR.n1056 VPWR.n1037 3.4105
R4750 VPWR.n1754 VPWR.n1753 3.4105
R4751 VPWR.n1756 VPWR.n1755 3.4105
R4752 VPWR.n1529 VPWR.n1045 3.4105
R4753 VPWR.n1531 VPWR.n1530 3.4105
R4754 VPWR.n1528 VPWR.n1145 3.4105
R4755 VPWR.n1527 VPWR.n1526 3.4105
R4756 VPWR.n1515 VPWR.n1514 3.4105
R4757 VPWR.n1513 VPWR.n1512 3.4105
R4758 VPWR.n1501 VPWR.n1500 3.4105
R4759 VPWR.n1499 VPWR.n1498 3.4105
R4760 VPWR.n1488 VPWR.n1487 3.4105
R4761 VPWR.n1587 VPWR.n1586 3.4105
R4762 VPWR.n1589 VPWR.n1588 3.4105
R4763 VPWR.n1448 VPWR.n1232 3.4105
R4764 VPWR.n1345 VPWR.n1341 3.38874
R4765 VPWR.n1384 VPWR.n1380 3.38874
R4766 VPWR.n1421 VPWR.n1417 3.38874
R4767 VPWR.n28 VPWR.n26 3.36211
R4768 VPWR.n30 VPWR.n28 3.36211
R4769 VPWR.n32 VPWR.n30 3.36211
R4770 VPWR.n34 VPWR.n32 3.36211
R4771 VPWR.n36 VPWR.n34 3.36211
R4772 VPWR.n38 VPWR.n36 3.36211
R4773 VPWR.n40 VPWR.n38 3.36211
R4774 VPWR.n42 VPWR.n40 3.36211
R4775 VPWR.n44 VPWR.n42 3.36211
R4776 VPWR.n46 VPWR.n44 3.36211
R4777 VPWR.n48 VPWR.n46 3.36211
R4778 VPWR.n50 VPWR.n48 3.36211
R4779 VPWR.n52 VPWR.n50 3.36211
R4780 VPWR.n54 VPWR.n52 3.36211
R4781 VPWR.t837 VPWR.t415 3.35739
R4782 VPWR.t541 VPWR.t1778 3.35739
R4783 VPWR.n2571 VPWR.n66 3.28012
R4784 VPWR.n2511 VPWR.n96 3.28012
R4785 VPWR.n2550 VPWR.n77 3.28012
R4786 VPWR.n2440 VPWR.n77 3.28012
R4787 VPWR.n2547 VPWR.n78 3.28012
R4788 VPWR.n2443 VPWR.n78 3.28012
R4789 VPWR.n2535 VPWR.n84 3.28012
R4790 VPWR.n2453 VPWR.n84 3.28012
R4791 VPWR.n2453 VPWR.n366 3.28012
R4792 VPWR.n2526 VPWR.n89 3.28012
R4793 VPWR.n2460 VPWR.n89 3.28012
R4794 VPWR.n2460 VPWR.n363 3.28012
R4795 VPWR.n1498 VPWR.n1497 3.28012
R4796 VPWR.n1497 VPWR.n939 3.28012
R4797 VPWR.n1872 VPWR.n939 3.28012
R4798 VPWR.n1872 VPWR.n858 3.28012
R4799 VPWR.n1934 VPWR.n858 3.28012
R4800 VPWR.n1934 VPWR.n747 3.28012
R4801 VPWR.n2068 VPWR.n747 3.28012
R4802 VPWR.n2068 VPWR.n666 3.28012
R4803 VPWR.n2130 VPWR.n666 3.28012
R4804 VPWR.n2130 VPWR.n555 3.28012
R4805 VPWR.n2264 VPWR.n555 3.28012
R4806 VPWR.n2264 VPWR.n474 3.28012
R4807 VPWR.n2326 VPWR.n474 3.28012
R4808 VPWR.n2326 VPWR.n363 3.28012
R4809 VPWR.n2523 VPWR.n90 3.28012
R4810 VPWR.n2463 VPWR.n90 3.28012
R4811 VPWR.n2463 VPWR.n362 3.28012
R4812 VPWR.n2323 VPWR.n362 3.28012
R4813 VPWR.n2323 VPWR.n475 3.28012
R4814 VPWR.n2267 VPWR.n475 3.28012
R4815 VPWR.n2267 VPWR.n554 3.28012
R4816 VPWR.n2127 VPWR.n554 3.28012
R4817 VPWR.n2127 VPWR.n667 3.28012
R4818 VPWR.n2071 VPWR.n667 3.28012
R4819 VPWR.n2071 VPWR.n746 3.28012
R4820 VPWR.n1931 VPWR.n746 3.28012
R4821 VPWR.n1931 VPWR.n859 3.28012
R4822 VPWR.n1875 VPWR.n859 3.28012
R4823 VPWR.n1489 VPWR.n1488 3.28012
R4824 VPWR.n1489 VPWR.n938 3.28012
R4825 VPWR.n1875 VPWR.n938 3.28012
R4826 VPWR.n1503 VPWR.n1501 3.28012
R4827 VPWR.n1503 VPWR.n942 3.28012
R4828 VPWR.n1865 VPWR.n942 3.28012
R4829 VPWR.n1865 VPWR.n855 3.28012
R4830 VPWR.n1941 VPWR.n855 3.28012
R4831 VPWR.n1941 VPWR.n750 3.28012
R4832 VPWR.n2061 VPWR.n750 3.28012
R4833 VPWR.n2061 VPWR.n663 3.28012
R4834 VPWR.n2137 VPWR.n663 3.28012
R4835 VPWR.n2137 VPWR.n558 3.28012
R4836 VPWR.n2257 VPWR.n558 3.28012
R4837 VPWR.n2257 VPWR.n471 3.28012
R4838 VPWR.n2333 VPWR.n471 3.28012
R4839 VPWR.n2333 VPWR.n366 3.28012
R4840 VPWR.n2538 VPWR.n83 3.28012
R4841 VPWR.n2450 VPWR.n83 3.28012
R4842 VPWR.n2450 VPWR.n367 3.28012
R4843 VPWR.n2336 VPWR.n367 3.28012
R4844 VPWR.n2336 VPWR.n470 3.28012
R4845 VPWR.n2254 VPWR.n470 3.28012
R4846 VPWR.n2254 VPWR.n559 3.28012
R4847 VPWR.n2140 VPWR.n559 3.28012
R4848 VPWR.n2140 VPWR.n662 3.28012
R4849 VPWR.n2058 VPWR.n662 3.28012
R4850 VPWR.n2058 VPWR.n751 3.28012
R4851 VPWR.n1944 VPWR.n751 3.28012
R4852 VPWR.n1944 VPWR.n854 3.28012
R4853 VPWR.n1862 VPWR.n854 3.28012
R4854 VPWR.n1512 VPWR.n1511 3.28012
R4855 VPWR.n1511 VPWR.n943 3.28012
R4856 VPWR.n1862 VPWR.n943 3.28012
R4857 VPWR.n1517 VPWR.n1515 3.28012
R4858 VPWR.n1517 VPWR.n946 3.28012
R4859 VPWR.n1855 VPWR.n946 3.28012
R4860 VPWR.n1855 VPWR.n851 3.28012
R4861 VPWR.n1951 VPWR.n851 3.28012
R4862 VPWR.n1951 VPWR.n754 3.28012
R4863 VPWR.n2051 VPWR.n754 3.28012
R4864 VPWR.n2051 VPWR.n659 3.28012
R4865 VPWR.n2147 VPWR.n659 3.28012
R4866 VPWR.n2147 VPWR.n562 3.28012
R4867 VPWR.n2247 VPWR.n562 3.28012
R4868 VPWR.n2247 VPWR.n467 3.28012
R4869 VPWR.n2343 VPWR.n467 3.28012
R4870 VPWR.n2343 VPWR.n370 3.28012
R4871 VPWR.n2443 VPWR.n370 3.28012
R4872 VPWR.n2514 VPWR.n95 3.28012
R4873 VPWR.n2470 VPWR.n95 3.28012
R4874 VPWR.n2470 VPWR.n359 3.28012
R4875 VPWR.n2316 VPWR.n359 3.28012
R4876 VPWR.n2316 VPWR.n478 3.28012
R4877 VPWR.n2274 VPWR.n478 3.28012
R4878 VPWR.n2274 VPWR.n551 3.28012
R4879 VPWR.n2120 VPWR.n551 3.28012
R4880 VPWR.n2120 VPWR.n670 3.28012
R4881 VPWR.n2078 VPWR.n670 3.28012
R4882 VPWR.n2078 VPWR.n743 3.28012
R4883 VPWR.n1924 VPWR.n743 3.28012
R4884 VPWR.n1924 VPWR.n862 3.28012
R4885 VPWR.n1882 VPWR.n862 3.28012
R4886 VPWR.n1882 VPWR.n935 3.28012
R4887 VPWR.n1586 VPWR.n1585 3.28012
R4888 VPWR.n1585 VPWR.n935 3.28012
R4889 VPWR.n1526 VPWR.n1525 3.28012
R4890 VPWR.n1525 VPWR.n947 3.28012
R4891 VPWR.n1852 VPWR.n947 3.28012
R4892 VPWR.n1852 VPWR.n850 3.28012
R4893 VPWR.n1954 VPWR.n850 3.28012
R4894 VPWR.n1954 VPWR.n755 3.28012
R4895 VPWR.n2048 VPWR.n755 3.28012
R4896 VPWR.n2048 VPWR.n658 3.28012
R4897 VPWR.n2150 VPWR.n658 3.28012
R4898 VPWR.n2150 VPWR.n563 3.28012
R4899 VPWR.n2244 VPWR.n563 3.28012
R4900 VPWR.n2244 VPWR.n466 3.28012
R4901 VPWR.n2346 VPWR.n466 3.28012
R4902 VPWR.n2346 VPWR.n371 3.28012
R4903 VPWR.n2440 VPWR.n371 3.28012
R4904 VPWR.n2559 VPWR.n72 3.28012
R4905 VPWR.n2433 VPWR.n72 3.28012
R4906 VPWR.n2433 VPWR.n374 3.28012
R4907 VPWR.n2353 VPWR.n374 3.28012
R4908 VPWR.n2353 VPWR.n463 3.28012
R4909 VPWR.n2237 VPWR.n463 3.28012
R4910 VPWR.n2237 VPWR.n566 3.28012
R4911 VPWR.n2157 VPWR.n566 3.28012
R4912 VPWR.n2157 VPWR.n655 3.28012
R4913 VPWR.n2041 VPWR.n655 3.28012
R4914 VPWR.n2041 VPWR.n758 3.28012
R4915 VPWR.n1961 VPWR.n758 3.28012
R4916 VPWR.n1961 VPWR.n847 3.28012
R4917 VPWR.n1845 VPWR.n847 3.28012
R4918 VPWR.n1845 VPWR.n950 3.28012
R4919 VPWR.n1539 VPWR.n1145 3.28012
R4920 VPWR.n1539 VPWR.n950 3.28012
R4921 VPWR.n1589 VPWR.n1128 3.28012
R4922 VPWR.n1128 VPWR.n934 3.28012
R4923 VPWR.n1885 VPWR.n934 3.28012
R4924 VPWR.n1885 VPWR.n863 3.28012
R4925 VPWR.n1921 VPWR.n863 3.28012
R4926 VPWR.n1921 VPWR.n742 3.28012
R4927 VPWR.n2081 VPWR.n742 3.28012
R4928 VPWR.n2081 VPWR.n671 3.28012
R4929 VPWR.n2117 VPWR.n671 3.28012
R4930 VPWR.n2117 VPWR.n550 3.28012
R4931 VPWR.n2277 VPWR.n550 3.28012
R4932 VPWR.n2277 VPWR.n479 3.28012
R4933 VPWR.n2313 VPWR.n479 3.28012
R4934 VPWR.n2313 VPWR.n358 3.28012
R4935 VPWR.n2473 VPWR.n358 3.28012
R4936 VPWR.n2473 VPWR.n96 3.28012
R4937 VPWR.n2562 VPWR.n71 3.28012
R4938 VPWR.n2430 VPWR.n71 3.28012
R4939 VPWR.n2430 VPWR.n375 3.28012
R4940 VPWR.n2356 VPWR.n375 3.28012
R4941 VPWR.n2356 VPWR.n462 3.28012
R4942 VPWR.n2234 VPWR.n462 3.28012
R4943 VPWR.n2234 VPWR.n567 3.28012
R4944 VPWR.n2160 VPWR.n567 3.28012
R4945 VPWR.n2160 VPWR.n654 3.28012
R4946 VPWR.n2038 VPWR.n654 3.28012
R4947 VPWR.n2038 VPWR.n759 3.28012
R4948 VPWR.n1964 VPWR.n759 3.28012
R4949 VPWR.n1964 VPWR.n846 3.28012
R4950 VPWR.n1842 VPWR.n846 3.28012
R4951 VPWR.n1842 VPWR.n951 3.28012
R4952 VPWR.n1532 VPWR.n951 3.28012
R4953 VPWR.n1532 VPWR.n1531 3.28012
R4954 VPWR.n1764 VPWR.n1045 3.28012
R4955 VPWR.n1764 VPWR.n954 3.28012
R4956 VPWR.n1835 VPWR.n954 3.28012
R4957 VPWR.n1835 VPWR.n843 3.28012
R4958 VPWR.n1971 VPWR.n843 3.28012
R4959 VPWR.n1971 VPWR.n762 3.28012
R4960 VPWR.n2031 VPWR.n762 3.28012
R4961 VPWR.n2031 VPWR.n651 3.28012
R4962 VPWR.n2167 VPWR.n651 3.28012
R4963 VPWR.n2167 VPWR.n570 3.28012
R4964 VPWR.n2227 VPWR.n570 3.28012
R4965 VPWR.n2227 VPWR.n459 3.28012
R4966 VPWR.n2363 VPWR.n459 3.28012
R4967 VPWR.n2363 VPWR.n378 3.28012
R4968 VPWR.n2423 VPWR.n378 3.28012
R4969 VPWR.n2423 VPWR.n66 3.28012
R4970 VPWR.n2583 VPWR.n60 3.28012
R4971 VPWR.n2413 VPWR.n60 3.28012
R4972 VPWR.n2413 VPWR.n382 3.28012
R4973 VPWR.n2373 VPWR.n382 3.28012
R4974 VPWR.n2373 VPWR.n455 3.28012
R4975 VPWR.n2217 VPWR.n455 3.28012
R4976 VPWR.n2217 VPWR.n574 3.28012
R4977 VPWR.n2177 VPWR.n574 3.28012
R4978 VPWR.n2177 VPWR.n647 3.28012
R4979 VPWR.n2021 VPWR.n647 3.28012
R4980 VPWR.n2021 VPWR.n766 3.28012
R4981 VPWR.n1981 VPWR.n766 3.28012
R4982 VPWR.n1981 VPWR.n839 3.28012
R4983 VPWR.n1825 VPWR.n839 3.28012
R4984 VPWR.n1825 VPWR.n958 3.28012
R4985 VPWR.n1752 VPWR.n958 3.28012
R4986 VPWR.n1753 VPWR.n1752 3.28012
R4987 VPWR.n1757 VPWR.n1756 3.28012
R4988 VPWR.n1757 VPWR.n955 3.28012
R4989 VPWR.n1832 VPWR.n955 3.28012
R4990 VPWR.n1832 VPWR.n842 3.28012
R4991 VPWR.n1974 VPWR.n842 3.28012
R4992 VPWR.n1974 VPWR.n763 3.28012
R4993 VPWR.n2028 VPWR.n763 3.28012
R4994 VPWR.n2028 VPWR.n650 3.28012
R4995 VPWR.n2170 VPWR.n650 3.28012
R4996 VPWR.n2170 VPWR.n571 3.28012
R4997 VPWR.n2224 VPWR.n571 3.28012
R4998 VPWR.n2224 VPWR.n458 3.28012
R4999 VPWR.n2366 VPWR.n458 3.28012
R5000 VPWR.n2366 VPWR.n379 3.28012
R5001 VPWR.n2420 VPWR.n379 3.28012
R5002 VPWR.n2420 VPWR.n65 3.28012
R5003 VPWR.n2574 VPWR.n65 3.28012
R5004 VPWR.n2586 VPWR.n59 3.28012
R5005 VPWR.n2410 VPWR.n59 3.28012
R5006 VPWR.n2410 VPWR.n383 3.28012
R5007 VPWR.n2376 VPWR.n383 3.28012
R5008 VPWR.n2376 VPWR.n454 3.28012
R5009 VPWR.n2214 VPWR.n454 3.28012
R5010 VPWR.n2214 VPWR.n575 3.28012
R5011 VPWR.n2180 VPWR.n575 3.28012
R5012 VPWR.n2180 VPWR.n646 3.28012
R5013 VPWR.n2018 VPWR.n646 3.28012
R5014 VPWR.n2018 VPWR.n767 3.28012
R5015 VPWR.n1984 VPWR.n767 3.28012
R5016 VPWR.n1984 VPWR.n838 3.28012
R5017 VPWR.n1822 VPWR.n838 3.28012
R5018 VPWR.n1822 VPWR.n959 3.28012
R5019 VPWR.n1788 VPWR.n959 3.28012
R5020 VPWR.n1788 VPWR.n1037 3.28012
R5021 VPWR.n1465 VPWR.n1232 3.28012
R5022 VPWR.n1465 VPWR.n931 3.28012
R5023 VPWR.n1892 VPWR.n931 3.28012
R5024 VPWR.n1892 VPWR.n929 3.28012
R5025 VPWR.n1914 VPWR.n929 3.28012
R5026 VPWR.n1914 VPWR.n739 3.28012
R5027 VPWR.n2088 VPWR.n739 3.28012
R5028 VPWR.n2088 VPWR.n737 3.28012
R5029 VPWR.n2110 VPWR.n737 3.28012
R5030 VPWR.n2110 VPWR.n547 3.28012
R5031 VPWR.n2284 VPWR.n547 3.28012
R5032 VPWR.n2284 VPWR.n545 3.28012
R5033 VPWR.n2306 VPWR.n545 3.28012
R5034 VPWR.n2306 VPWR.n355 3.28012
R5035 VPWR.n2480 VPWR.n355 3.28012
R5036 VPWR.n2480 VPWR.n353 3.28012
R5037 VPWR.n2502 VPWR.n353 3.28012
R5038 VPWR.n2404 VPWR.n22 3.28012
R5039 VPWR.n2404 VPWR.n449 3.28012
R5040 VPWR.n2382 VPWR.n449 3.28012
R5041 VPWR.n2382 VPWR.n451 3.28012
R5042 VPWR.n2208 VPWR.n451 3.28012
R5043 VPWR.n2208 VPWR.n641 3.28012
R5044 VPWR.n2186 VPWR.n641 3.28012
R5045 VPWR.n2186 VPWR.n643 3.28012
R5046 VPWR.n2012 VPWR.n643 3.28012
R5047 VPWR.n2012 VPWR.n833 3.28012
R5048 VPWR.n1990 VPWR.n833 3.28012
R5049 VPWR.n1990 VPWR.n835 3.28012
R5050 VPWR.n1816 VPWR.n835 3.28012
R5051 VPWR.n1816 VPWR.n1025 3.28012
R5052 VPWR.n1794 VPWR.n1025 3.28012
R5053 VPWR.n1794 VPWR.n1028 3.28012
R5054 VPWR.n2594 VPWR.n22 3.26393
R5055 VPWR.n2863 VPWR 3.18182
R5056 VPWR.n2832 VPWR.n2831 3.1005
R5057 VPWR.n2826 VPWR.n2825 3.1005
R5058 VPWR.n2846 VPWR.n2815 3.1005
R5059 VPWR.n1324 VPWR.n1322 3.01226
R5060 VPWR.n1328 VPWR.n1304 2.63579
R5061 VPWR.n2731 VPWR.n2730 2.25932
R5062 VPWR.n1447 VPWR.n1446 2.06026
R5063 VPWR.n1447 VPWR.n1026 1.78803
R5064 VPWR.n2384 VPWR.n2383 1.32852
R5065 VPWR.n2287 VPWR.n450 1.32852
R5066 VPWR.n2207 VPWR.n2206 1.32852
R5067 VPWR.n2205 VPWR.n2204 1.32852
R5068 VPWR.n2188 VPWR.n2187 1.32852
R5069 VPWR.n2091 VPWR.n642 1.32852
R5070 VPWR.n2011 VPWR.n2010 1.32852
R5071 VPWR.n2009 VPWR.n2008 1.32852
R5072 VPWR.n1992 VPWR.n1991 1.32852
R5073 VPWR.n1895 VPWR.n834 1.32852
R5074 VPWR.n2401 VPWR.n2400 1.32852
R5075 VPWR.n1815 VPWR.n1814 1.32852
R5076 VPWR.n2403 VPWR.n2402 1.32852
R5077 VPWR.n1813 VPWR.n1812 1.32852
R5078 VPWR.n2483 VPWR.n21 1.32852
R5079 VPWR.n1796 VPWR.n1795 1.32852
R5080 VPWR.n2596 VPWR.n2595 1.32852
R5081 VPWR.n1055 VPWR.n1026 1.32852
R5082 VPWR.n2482 VPWR 1.25994
R5083 VPWR VPWR.n354 1.25994
R5084 VPWR VPWR.n2304 1.25994
R5085 VPWR.n2303 VPWR 1.25994
R5086 VPWR.n2286 VPWR 1.25994
R5087 VPWR VPWR.n546 1.25994
R5088 VPWR VPWR.n2108 1.25994
R5089 VPWR.n2107 VPWR 1.25994
R5090 VPWR.n2090 VPWR 1.25994
R5091 VPWR VPWR.n738 1.25994
R5092 VPWR VPWR.n1912 1.25994
R5093 VPWR.n1911 VPWR 1.25994
R5094 VPWR.n1894 VPWR 1.25994
R5095 VPWR VPWR.n930 1.25994
R5096 VPWR.n2499 VPWR 1.25994
R5097 VPWR VPWR.n1450 1.25994
R5098 VPWR VPWR.n2500 1.25994
R5099 VPWR.n1449 VPWR 1.25994
R5100 VPWR.n2597 VPWR.n2596 1.144
R5101 VPWR.n2861 VPWR.n2860 0.936724
R5102 VPWR.n2592 VPWR 0.925943
R5103 VPWR VPWR.n1063 0.925943
R5104 VPWR.n2860 VPWR.n2816 0.925245
R5105 VPWR.n2569 VPWR.n67 0.904391
R5106 VPWR.n2509 VPWR.n97 0.904391
R5107 VPWR.n2552 VPWR.n76 0.904391
R5108 VPWR.n2545 VPWR.n79 0.904391
R5109 VPWR.n2533 VPWR.n85 0.904391
R5110 VPWR.n2528 VPWR.n88 0.904391
R5111 VPWR.n1222 VPWR.n1178 0.904391
R5112 VPWR.n2521 VPWR.n91 0.904391
R5113 VPWR.n1624 VPWR.n1102 0.904391
R5114 VPWR.n1640 VPWR.n1094 0.904391
R5115 VPWR.n2540 VPWR.n82 0.904391
R5116 VPWR.n1651 VPWR.n1092 0.904391
R5117 VPWR.n1211 VPWR.n1210 0.904391
R5118 VPWR.n2516 VPWR.n94 0.904391
R5119 VPWR.n1613 VPWR.n1104 0.904391
R5120 VPWR.n1667 VPWR.n1084 0.904391
R5121 VPWR.n2557 VPWR.n73 0.904391
R5122 VPWR.n1678 VPWR.n1082 0.904391
R5123 VPWR.n1591 VPWR.n1127 0.904391
R5124 VPWR.n2564 VPWR.n70 0.904391
R5125 VPWR.n1197 VPWR.n1196 0.904391
R5126 VPWR.n1694 VPWR.n1074 0.904391
R5127 VPWR.n1742 VPWR.n1057 0.904391
R5128 VPWR.n1705 VPWR.n1071 0.904391
R5129 VPWR.n2581 VPWR.n61 0.904391
R5130 VPWR.n2588 VPWR.n58 0.904391
R5131 VPWR.n1737 VPWR.n1735 0.904391
R5132 VPWR.n1597 VPWR.n1596 0.904391
R5133 VPWR.n2504 VPWR.n289 0.904391
R5134 VPWR.n2576 VPWR.n64 0.904391
R5135 VPWR VPWR.n2863 0.812229
R5136 VPWR.n140 VPWR.n64 0.675548
R5137 VPWR.n152 VPWR.n67 0.675548
R5138 VPWR.n164 VPWR.n70 0.675548
R5139 VPWR.n176 VPWR.n73 0.675548
R5140 VPWR.n188 VPWR.n76 0.675548
R5141 VPWR.n200 VPWR.n79 0.675548
R5142 VPWR.n212 VPWR.n82 0.675548
R5143 VPWR.n224 VPWR.n85 0.675548
R5144 VPWR.n236 VPWR.n88 0.675548
R5145 VPWR.n248 VPWR.n91 0.675548
R5146 VPWR.n260 VPWR.n94 0.675548
R5147 VPWR.n272 VPWR.n97 0.675548
R5148 VPWR.n289 VPWR.n288 0.675548
R5149 VPWR.n128 VPWR.n61 0.675548
R5150 VPWR.n117 VPWR.n58 0.675548
R5151 VPWR.n1735 VPWR.n1734 0.675548
R5152 VPWR.n1719 VPWR.n1057 0.675548
R5153 VPWR.n1707 VPWR.n1705 0.675548
R5154 VPWR.n1696 VPWR.n1694 0.675548
R5155 VPWR.n1196 VPWR.n1195 0.675548
R5156 VPWR.n1680 VPWR.n1678 0.675548
R5157 VPWR.n1669 VPWR.n1667 0.675548
R5158 VPWR.n1210 VPWR.n1209 0.675548
R5159 VPWR.n1653 VPWR.n1651 0.675548
R5160 VPWR.n1642 VPWR.n1640 0.675548
R5161 VPWR.n1178 VPWR.n1177 0.675548
R5162 VPWR.n1626 VPWR.n1624 0.675548
R5163 VPWR.n1615 VPWR.n1613 0.675548
R5164 VPWR.n1127 VPWR.n1126 0.675548
R5165 VPWR.n1599 VPWR.n1597 0.675548
R5166 VPWR.n2806 VPWR.n2805 0.672385
R5167 VPWR.n2790 VPWR.n2785 0.672385
R5168 VPWR.n2770 VPWR.n2765 0.672385
R5169 VPWR.n2751 VPWR.n2746 0.672385
R5170 VPWR.n7 VPWR 0.63497
R5171 VPWR.n1242 VPWR 0.63497
R5172 VPWR.n1265 VPWR 0.63497
R5173 VPWR.n1289 VPWR 0.63497
R5174 VPWR.n24 VPWR 0.499542
R5175 VPWR.n2814 VPWR.n2813 0.442692
R5176 VPWR.n1120 VPWR.n1118 0.404056
R5177 VPWR.n144 VPWR.n138 0.404056
R5178 VPWR.n156 VPWR.n150 0.404056
R5179 VPWR.n168 VPWR.n162 0.404056
R5180 VPWR.n180 VPWR.n174 0.404056
R5181 VPWR.n192 VPWR.n186 0.404056
R5182 VPWR.n204 VPWR.n198 0.404056
R5183 VPWR.n216 VPWR.n210 0.404056
R5184 VPWR.n228 VPWR.n222 0.404056
R5185 VPWR.n240 VPWR.n234 0.404056
R5186 VPWR.n252 VPWR.n246 0.404056
R5187 VPWR.n264 VPWR.n258 0.404056
R5188 VPWR.n276 VPWR.n270 0.404056
R5189 VPWR.n283 VPWR.n101 0.404056
R5190 VPWR.n110 VPWR.n105 0.404056
R5191 VPWR.n132 VPWR.n126 0.404056
R5192 VPWR.n121 VPWR.n115 0.404056
R5193 VPWR.n1729 VPWR.n1065 0.404056
R5194 VPWR.n1723 VPWR.n1717 0.404056
R5195 VPWR.n1711 VPWR.n1070 0.404056
R5196 VPWR.n1704 VPWR.n1702 0.404056
R5197 VPWR.n1693 VPWR.n1691 0.404056
R5198 VPWR.n1684 VPWR.n1081 0.404056
R5199 VPWR.n1677 VPWR.n1675 0.404056
R5200 VPWR.n1666 VPWR.n1664 0.404056
R5201 VPWR.n1657 VPWR.n1091 0.404056
R5202 VPWR.n1650 VPWR.n1648 0.404056
R5203 VPWR.n1639 VPWR.n1637 0.404056
R5204 VPWR.n1630 VPWR.n1101 0.404056
R5205 VPWR.n1623 VPWR.n1621 0.404056
R5206 VPWR.n1612 VPWR.n1610 0.404056
R5207 VPWR.n1603 VPWR.n1111 0.404056
R5208 VPWR.n2860 VPWR.n2859 0.388
R5209 VPWR.n1608 VPWR.n1607 0.349144
R5210 VPWR.n1608 VPWR.n1099 0.349144
R5211 VPWR.n1634 VPWR.n1099 0.349144
R5212 VPWR.n1635 VPWR.n1634 0.349144
R5213 VPWR.n1635 VPWR.n1089 0.349144
R5214 VPWR.n1661 VPWR.n1089 0.349144
R5215 VPWR.n1662 VPWR.n1661 0.349144
R5216 VPWR.n1662 VPWR.n1079 0.349144
R5217 VPWR.n1688 VPWR.n1079 0.349144
R5218 VPWR.n1689 VPWR.n1688 0.349144
R5219 VPWR.n1689 VPWR.n1068 0.349144
R5220 VPWR.n1715 VPWR.n1068 0.349144
R5221 VPWR.n1727 VPWR.n1715 0.349144
R5222 VPWR.n281 VPWR.n280 0.349144
R5223 VPWR.n280 VPWR.n268 0.349144
R5224 VPWR.n268 VPWR.n256 0.349144
R5225 VPWR.n256 VPWR.n244 0.349144
R5226 VPWR.n244 VPWR.n232 0.349144
R5227 VPWR.n232 VPWR.n220 0.349144
R5228 VPWR.n220 VPWR.n208 0.349144
R5229 VPWR.n208 VPWR.n196 0.349144
R5230 VPWR.n196 VPWR.n184 0.349144
R5231 VPWR.n184 VPWR.n172 0.349144
R5232 VPWR.n172 VPWR.n160 0.349144
R5233 VPWR.n160 VPWR.n148 0.349144
R5234 VPWR.n148 VPWR.n136 0.349144
R5235 VPWR.n1462 VPWR.n1456 0.346131
R5236 VPWR.n1461 VPWR.n1457 0.346131
R5237 VPWR.n1582 VPWR.n1136 0.346131
R5238 VPWR.n1581 VPWR.n1577 0.346131
R5239 VPWR.n1576 VPWR.n1572 0.346131
R5240 VPWR.n1571 VPWR.n1567 0.346131
R5241 VPWR.n1566 VPWR.n1562 0.346131
R5242 VPWR.n1561 VPWR.n1557 0.346131
R5243 VPWR.n1556 VPWR.n1552 0.346131
R5244 VPWR.n1551 VPWR.n1547 0.346131
R5245 VPWR.n1546 VPWR.n1542 0.346131
R5246 VPWR.n1767 VPWR.n1042 0.346131
R5247 VPWR.n1784 VPWR.n1780 0.346131
R5248 VPWR.n1785 VPWR.n1776 0.346131
R5249 VPWR.n1772 VPWR.n1771 0.346131
R5250 VPWR.n2862 VPWR.n2861 0.304571
R5251 VPWR.n2594 VPWR.n55 0.300179
R5252 VPWR.n1118 VPWR.n1113 0.286958
R5253 VPWR.n145 VPWR.n144 0.286958
R5254 VPWR.n157 VPWR.n156 0.286958
R5255 VPWR.n169 VPWR.n168 0.286958
R5256 VPWR.n181 VPWR.n180 0.286958
R5257 VPWR.n193 VPWR.n192 0.286958
R5258 VPWR.n205 VPWR.n204 0.286958
R5259 VPWR.n217 VPWR.n216 0.286958
R5260 VPWR.n229 VPWR.n228 0.286958
R5261 VPWR.n241 VPWR.n240 0.286958
R5262 VPWR.n253 VPWR.n252 0.286958
R5263 VPWR.n265 VPWR.n264 0.286958
R5264 VPWR.n277 VPWR.n276 0.286958
R5265 VPWR.n283 VPWR.n102 0.286958
R5266 VPWR.n111 VPWR.n110 0.286958
R5267 VPWR.n133 VPWR.n132 0.286958
R5268 VPWR.n122 VPWR.n121 0.286958
R5269 VPWR.n1729 VPWR.n1066 0.286958
R5270 VPWR.n1724 VPWR.n1723 0.286958
R5271 VPWR.n1712 VPWR.n1711 0.286958
R5272 VPWR.n1702 VPWR.n1072 0.286958
R5273 VPWR.n1691 VPWR.n1075 0.286958
R5274 VPWR.n1685 VPWR.n1684 0.286958
R5275 VPWR.n1675 VPWR.n1083 0.286958
R5276 VPWR.n1664 VPWR.n1085 0.286958
R5277 VPWR.n1658 VPWR.n1657 0.286958
R5278 VPWR.n1648 VPWR.n1093 0.286958
R5279 VPWR.n1637 VPWR.n1095 0.286958
R5280 VPWR.n1631 VPWR.n1630 0.286958
R5281 VPWR.n1621 VPWR.n1103 0.286958
R5282 VPWR.n1610 VPWR.n1105 0.286958
R5283 VPWR.n1604 VPWR.n1603 0.286958
R5284 VPWR.n55 VPWR 0.2505
R5285 VPWR VPWR.n2481 0.249238
R5286 VPWR.n2472 VPWR 0.249238
R5287 VPWR VPWR.n2471 0.249238
R5288 VPWR.n2385 VPWR 0.249238
R5289 VPWR.n2386 VPWR 0.249238
R5290 VPWR.n2387 VPWR 0.249238
R5291 VPWR.n2388 VPWR 0.249238
R5292 VPWR.n2305 VPWR 0.249238
R5293 VPWR.n2314 VPWR 0.249238
R5294 VPWR.n2315 VPWR 0.249238
R5295 VPWR.n2324 VPWR 0.249238
R5296 VPWR.n2325 VPWR 0.249238
R5297 VPWR.n2383 VPWR 0.249238
R5298 VPWR.n2375 VPWR 0.249238
R5299 VPWR.n2374 VPWR 0.249238
R5300 VPWR.n2365 VPWR 0.249238
R5301 VPWR.n2364 VPWR 0.249238
R5302 VPWR.n2355 VPWR 0.249238
R5303 VPWR.n2354 VPWR 0.249238
R5304 VPWR.n2345 VPWR 0.249238
R5305 VPWR.n2344 VPWR 0.249238
R5306 VPWR.n2335 VPWR 0.249238
R5307 VPWR.n2334 VPWR 0.249238
R5308 VPWR VPWR.n2302 0.249238
R5309 VPWR VPWR.n2301 0.249238
R5310 VPWR VPWR.n2300 0.249238
R5311 VPWR VPWR.n2299 0.249238
R5312 VPWR VPWR.n2298 0.249238
R5313 VPWR VPWR.n2287 0.249238
R5314 VPWR VPWR.n2288 0.249238
R5315 VPWR VPWR.n2289 0.249238
R5316 VPWR VPWR.n2290 0.249238
R5317 VPWR VPWR.n2291 0.249238
R5318 VPWR VPWR.n2292 0.249238
R5319 VPWR VPWR.n2293 0.249238
R5320 VPWR VPWR.n2294 0.249238
R5321 VPWR VPWR.n2295 0.249238
R5322 VPWR VPWR.n2296 0.249238
R5323 VPWR VPWR.n2297 0.249238
R5324 VPWR VPWR.n2285 0.249238
R5325 VPWR.n2276 VPWR 0.249238
R5326 VPWR VPWR.n2275 0.249238
R5327 VPWR.n2266 VPWR 0.249238
R5328 VPWR VPWR.n2265 0.249238
R5329 VPWR.n2207 VPWR 0.249238
R5330 VPWR VPWR.n2215 0.249238
R5331 VPWR.n2216 VPWR 0.249238
R5332 VPWR VPWR.n2225 0.249238
R5333 VPWR.n2226 VPWR 0.249238
R5334 VPWR VPWR.n2235 0.249238
R5335 VPWR.n2236 VPWR 0.249238
R5336 VPWR VPWR.n2245 0.249238
R5337 VPWR.n2246 VPWR 0.249238
R5338 VPWR VPWR.n2255 0.249238
R5339 VPWR.n2256 VPWR 0.249238
R5340 VPWR.n2189 VPWR 0.249238
R5341 VPWR.n2190 VPWR 0.249238
R5342 VPWR.n2191 VPWR 0.249238
R5343 VPWR.n2192 VPWR 0.249238
R5344 VPWR.n2193 VPWR 0.249238
R5345 VPWR.n2204 VPWR 0.249238
R5346 VPWR.n2203 VPWR 0.249238
R5347 VPWR.n2202 VPWR 0.249238
R5348 VPWR.n2201 VPWR 0.249238
R5349 VPWR.n2200 VPWR 0.249238
R5350 VPWR.n2199 VPWR 0.249238
R5351 VPWR.n2198 VPWR 0.249238
R5352 VPWR.n2197 VPWR 0.249238
R5353 VPWR.n2196 VPWR 0.249238
R5354 VPWR.n2195 VPWR 0.249238
R5355 VPWR.n2194 VPWR 0.249238
R5356 VPWR.n2109 VPWR 0.249238
R5357 VPWR.n2118 VPWR 0.249238
R5358 VPWR.n2119 VPWR 0.249238
R5359 VPWR.n2128 VPWR 0.249238
R5360 VPWR.n2129 VPWR 0.249238
R5361 VPWR.n2187 VPWR 0.249238
R5362 VPWR.n2179 VPWR 0.249238
R5363 VPWR.n2178 VPWR 0.249238
R5364 VPWR.n2169 VPWR 0.249238
R5365 VPWR.n2168 VPWR 0.249238
R5366 VPWR.n2159 VPWR 0.249238
R5367 VPWR.n2158 VPWR 0.249238
R5368 VPWR.n2149 VPWR 0.249238
R5369 VPWR.n2148 VPWR 0.249238
R5370 VPWR.n2139 VPWR 0.249238
R5371 VPWR.n2138 VPWR 0.249238
R5372 VPWR VPWR.n2106 0.249238
R5373 VPWR VPWR.n2105 0.249238
R5374 VPWR VPWR.n2104 0.249238
R5375 VPWR VPWR.n2103 0.249238
R5376 VPWR VPWR.n2102 0.249238
R5377 VPWR VPWR.n2091 0.249238
R5378 VPWR VPWR.n2092 0.249238
R5379 VPWR VPWR.n2093 0.249238
R5380 VPWR VPWR.n2094 0.249238
R5381 VPWR VPWR.n2095 0.249238
R5382 VPWR VPWR.n2096 0.249238
R5383 VPWR VPWR.n2097 0.249238
R5384 VPWR VPWR.n2098 0.249238
R5385 VPWR VPWR.n2099 0.249238
R5386 VPWR VPWR.n2100 0.249238
R5387 VPWR VPWR.n2101 0.249238
R5388 VPWR VPWR.n2089 0.249238
R5389 VPWR.n2080 VPWR 0.249238
R5390 VPWR VPWR.n2079 0.249238
R5391 VPWR.n2070 VPWR 0.249238
R5392 VPWR VPWR.n2069 0.249238
R5393 VPWR.n2011 VPWR 0.249238
R5394 VPWR VPWR.n2019 0.249238
R5395 VPWR.n2020 VPWR 0.249238
R5396 VPWR VPWR.n2029 0.249238
R5397 VPWR.n2030 VPWR 0.249238
R5398 VPWR VPWR.n2039 0.249238
R5399 VPWR.n2040 VPWR 0.249238
R5400 VPWR VPWR.n2049 0.249238
R5401 VPWR.n2050 VPWR 0.249238
R5402 VPWR VPWR.n2059 0.249238
R5403 VPWR.n2060 VPWR 0.249238
R5404 VPWR.n1993 VPWR 0.249238
R5405 VPWR.n1994 VPWR 0.249238
R5406 VPWR.n1995 VPWR 0.249238
R5407 VPWR.n1996 VPWR 0.249238
R5408 VPWR.n1997 VPWR 0.249238
R5409 VPWR.n2008 VPWR 0.249238
R5410 VPWR.n2007 VPWR 0.249238
R5411 VPWR.n2006 VPWR 0.249238
R5412 VPWR.n2005 VPWR 0.249238
R5413 VPWR.n2004 VPWR 0.249238
R5414 VPWR.n2003 VPWR 0.249238
R5415 VPWR.n2002 VPWR 0.249238
R5416 VPWR.n2001 VPWR 0.249238
R5417 VPWR.n2000 VPWR 0.249238
R5418 VPWR.n1999 VPWR 0.249238
R5419 VPWR.n1998 VPWR 0.249238
R5420 VPWR.n1913 VPWR 0.249238
R5421 VPWR.n1922 VPWR 0.249238
R5422 VPWR.n1923 VPWR 0.249238
R5423 VPWR.n1932 VPWR 0.249238
R5424 VPWR.n1933 VPWR 0.249238
R5425 VPWR.n1991 VPWR 0.249238
R5426 VPWR.n1983 VPWR 0.249238
R5427 VPWR.n1982 VPWR 0.249238
R5428 VPWR.n1973 VPWR 0.249238
R5429 VPWR.n1972 VPWR 0.249238
R5430 VPWR.n1963 VPWR 0.249238
R5431 VPWR.n1962 VPWR 0.249238
R5432 VPWR.n1953 VPWR 0.249238
R5433 VPWR.n1952 VPWR 0.249238
R5434 VPWR.n1943 VPWR 0.249238
R5435 VPWR.n1942 VPWR 0.249238
R5436 VPWR VPWR.n1910 0.249238
R5437 VPWR VPWR.n1909 0.249238
R5438 VPWR VPWR.n1908 0.249238
R5439 VPWR VPWR.n1907 0.249238
R5440 VPWR VPWR.n1906 0.249238
R5441 VPWR VPWR.n1895 0.249238
R5442 VPWR VPWR.n1896 0.249238
R5443 VPWR VPWR.n1897 0.249238
R5444 VPWR VPWR.n1898 0.249238
R5445 VPWR VPWR.n1899 0.249238
R5446 VPWR VPWR.n1900 0.249238
R5447 VPWR VPWR.n1901 0.249238
R5448 VPWR VPWR.n1902 0.249238
R5449 VPWR VPWR.n1903 0.249238
R5450 VPWR VPWR.n1904 0.249238
R5451 VPWR VPWR.n1905 0.249238
R5452 VPWR.n2400 VPWR 0.249238
R5453 VPWR.n2399 VPWR 0.249238
R5454 VPWR.n2398 VPWR 0.249238
R5455 VPWR.n2397 VPWR 0.249238
R5456 VPWR.n2396 VPWR 0.249238
R5457 VPWR.n2395 VPWR 0.249238
R5458 VPWR.n2394 VPWR 0.249238
R5459 VPWR.n2393 VPWR 0.249238
R5460 VPWR.n2392 VPWR 0.249238
R5461 VPWR.n2391 VPWR 0.249238
R5462 VPWR.n2390 VPWR 0.249238
R5463 VPWR.n2389 VPWR 0.249238
R5464 VPWR VPWR.n1893 0.249238
R5465 VPWR.n1884 VPWR 0.249238
R5466 VPWR VPWR.n1883 0.249238
R5467 VPWR.n1874 VPWR 0.249238
R5468 VPWR VPWR.n1873 0.249238
R5469 VPWR.n1864 VPWR 0.249238
R5470 VPWR.n1815 VPWR 0.249238
R5471 VPWR VPWR.n1823 0.249238
R5472 VPWR.n1824 VPWR 0.249238
R5473 VPWR VPWR.n1833 0.249238
R5474 VPWR.n1834 VPWR 0.249238
R5475 VPWR VPWR.n1843 0.249238
R5476 VPWR.n1844 VPWR 0.249238
R5477 VPWR VPWR.n1853 0.249238
R5478 VPWR.n1854 VPWR 0.249238
R5479 VPWR VPWR.n1863 0.249238
R5480 VPWR.n2403 VPWR 0.249238
R5481 VPWR VPWR.n2411 0.249238
R5482 VPWR.n2412 VPWR 0.249238
R5483 VPWR VPWR.n2421 0.249238
R5484 VPWR.n2422 VPWR 0.249238
R5485 VPWR VPWR.n2431 0.249238
R5486 VPWR.n2432 VPWR 0.249238
R5487 VPWR VPWR.n2441 0.249238
R5488 VPWR.n2442 VPWR 0.249238
R5489 VPWR VPWR.n2451 0.249238
R5490 VPWR.n2452 VPWR 0.249238
R5491 VPWR VPWR.n2461 0.249238
R5492 VPWR.n2462 VPWR 0.249238
R5493 VPWR.n1797 VPWR 0.249238
R5494 VPWR.n1798 VPWR 0.249238
R5495 VPWR.n1799 VPWR 0.249238
R5496 VPWR.n1800 VPWR 0.249238
R5497 VPWR.n1801 VPWR 0.249238
R5498 VPWR.n1802 VPWR 0.249238
R5499 VPWR.n1803 VPWR 0.249238
R5500 VPWR.n1804 VPWR 0.249238
R5501 VPWR.n1805 VPWR 0.249238
R5502 VPWR.n1812 VPWR 0.249238
R5503 VPWR.n1811 VPWR 0.249238
R5504 VPWR.n1810 VPWR 0.249238
R5505 VPWR.n1809 VPWR 0.249238
R5506 VPWR.n1808 VPWR 0.249238
R5507 VPWR.n1807 VPWR 0.249238
R5508 VPWR.n1806 VPWR 0.249238
R5509 VPWR VPWR.n2498 0.249238
R5510 VPWR VPWR.n2497 0.249238
R5511 VPWR VPWR.n2496 0.249238
R5512 VPWR VPWR.n2495 0.249238
R5513 VPWR VPWR.n2494 0.249238
R5514 VPWR VPWR.n2493 0.249238
R5515 VPWR VPWR.n2492 0.249238
R5516 VPWR VPWR.n2491 0.249238
R5517 VPWR VPWR.n2490 0.249238
R5518 VPWR VPWR.n2489 0.249238
R5519 VPWR VPWR.n2488 0.249238
R5520 VPWR VPWR.n2483 0.249238
R5521 VPWR VPWR.n2484 0.249238
R5522 VPWR VPWR.n2485 0.249238
R5523 VPWR VPWR.n2486 0.249238
R5524 VPWR VPWR.n2487 0.249238
R5525 VPWR.n2501 VPWR 0.249238
R5526 VPWR.n2512 VPWR 0.249238
R5527 VPWR.n2513 VPWR 0.249238
R5528 VPWR.n2524 VPWR 0.249238
R5529 VPWR.n2525 VPWR 0.249238
R5530 VPWR.n2536 VPWR 0.249238
R5531 VPWR.n2537 VPWR 0.249238
R5532 VPWR.n2548 VPWR 0.249238
R5533 VPWR.n2549 VPWR 0.249238
R5534 VPWR.n2560 VPWR 0.249238
R5535 VPWR.n2561 VPWR 0.249238
R5536 VPWR.n2572 VPWR 0.249238
R5537 VPWR.n2573 VPWR 0.249238
R5538 VPWR.n2584 VPWR 0.249238
R5539 VPWR.n2585 VPWR 0.249238
R5540 VPWR.n2595 VPWR 0.249238
R5541 VPWR VPWR.n1055 0.249238
R5542 VPWR VPWR.n1056 0.249238
R5543 VPWR VPWR.n1754 0.249238
R5544 VPWR.n1755 VPWR 0.249238
R5545 VPWR VPWR.n1529 0.249238
R5546 VPWR.n1530 VPWR 0.249238
R5547 VPWR.n1528 VPWR 0.249238
R5548 VPWR.n1527 VPWR 0.249238
R5549 VPWR.n1514 VPWR 0.249238
R5550 VPWR.n1513 VPWR 0.249238
R5551 VPWR.n1500 VPWR 0.249238
R5552 VPWR.n1499 VPWR 0.249238
R5553 VPWR.n1487 VPWR 0.249238
R5554 VPWR VPWR.n1587 0.249238
R5555 VPWR.n1588 VPWR 0.249238
R5556 VPWR VPWR.n1448 0.249238
R5557 VPWR.n2861 VPWR.n2815 0.245065
R5558 VPWR.n2813 VPWR.n2797 0.213567
R5559 VPWR.n2797 VPWR.n2778 0.213567
R5560 VPWR.n2778 VPWR.n2758 0.213567
R5561 VPWR.n2758 VPWR.n2739 0.213567
R5562 VPWR.n2739 VPWR.n2703 0.213567
R5563 VPWR.n2703 VPWR.n2665 0.213567
R5564 VPWR.n2665 VPWR.n2628 0.213567
R5565 VPWR.n1446 VPWR.n1414 0.213567
R5566 VPWR.n1414 VPWR.n1376 0.213567
R5567 VPWR.n1376 VPWR.n1337 0.213567
R5568 VPWR.n1337 VPWR.n1302 0.213567
R5569 VPWR.n1302 VPWR.n1279 0.213567
R5570 VPWR.n1279 VPWR.n1255 0.213567
R5571 VPWR.n1255 VPWR.n19 0.213567
R5572 VPWR VPWR.n2862 0.204304
R5573 VPWR.n1449 VPWR.n1447 0.179202
R5574 VPWR.n1450 VPWR.n1449 0.154425
R5575 VPWR.n1450 VPWR.n930 0.154425
R5576 VPWR.n1894 VPWR.n930 0.154425
R5577 VPWR.n1911 VPWR.n1894 0.154425
R5578 VPWR.n1912 VPWR.n1911 0.154425
R5579 VPWR.n1912 VPWR.n738 0.154425
R5580 VPWR.n2090 VPWR.n738 0.154425
R5581 VPWR.n2107 VPWR.n2090 0.154425
R5582 VPWR.n2108 VPWR.n2107 0.154425
R5583 VPWR.n2108 VPWR.n546 0.154425
R5584 VPWR.n2286 VPWR.n546 0.154425
R5585 VPWR.n2303 VPWR.n2286 0.154425
R5586 VPWR.n2304 VPWR.n2303 0.154425
R5587 VPWR.n2304 VPWR.n354 0.154425
R5588 VPWR.n2482 VPWR.n354 0.154425
R5589 VPWR.n2499 VPWR.n2482 0.154425
R5590 VPWR.n2500 VPWR.n2499 0.154425
R5591 VPWR.n1796 VPWR.n1026 0.154425
R5592 VPWR.n1813 VPWR.n1796 0.154425
R5593 VPWR.n1814 VPWR.n1813 0.154425
R5594 VPWR.n1814 VPWR.n834 0.154425
R5595 VPWR.n1992 VPWR.n834 0.154425
R5596 VPWR.n2009 VPWR.n1992 0.154425
R5597 VPWR.n2010 VPWR.n2009 0.154425
R5598 VPWR.n2010 VPWR.n642 0.154425
R5599 VPWR.n2188 VPWR.n642 0.154425
R5600 VPWR.n2205 VPWR.n2188 0.154425
R5601 VPWR.n2206 VPWR.n2205 0.154425
R5602 VPWR.n2206 VPWR.n450 0.154425
R5603 VPWR.n2384 VPWR.n450 0.154425
R5604 VPWR.n2401 VPWR.n2384 0.154425
R5605 VPWR.n2402 VPWR.n2401 0.154425
R5606 VPWR.n2402 VPWR.n21 0.154425
R5607 VPWR.n2596 VPWR.n21 0.154425
R5608 VPWR.n8 VPWR.n7 0.147771
R5609 VPWR.n1243 VPWR.n1242 0.147771
R5610 VPWR.n1266 VPWR.n1265 0.147771
R5611 VPWR.n1290 VPWR.n1289 0.147771
R5612 VPWR.n1113 VPWR 0.135917
R5613 VPWR.n145 VPWR 0.135917
R5614 VPWR.n157 VPWR 0.135917
R5615 VPWR.n169 VPWR 0.135917
R5616 VPWR.n181 VPWR 0.135917
R5617 VPWR.n193 VPWR 0.135917
R5618 VPWR.n205 VPWR 0.135917
R5619 VPWR.n217 VPWR 0.135917
R5620 VPWR.n229 VPWR 0.135917
R5621 VPWR.n241 VPWR 0.135917
R5622 VPWR.n253 VPWR 0.135917
R5623 VPWR.n265 VPWR 0.135917
R5624 VPWR.n277 VPWR 0.135917
R5625 VPWR.n102 VPWR 0.135917
R5626 VPWR.n111 VPWR 0.135917
R5627 VPWR.n133 VPWR 0.135917
R5628 VPWR.n122 VPWR 0.135917
R5629 VPWR.n1066 VPWR 0.135917
R5630 VPWR.n1724 VPWR 0.135917
R5631 VPWR.n1712 VPWR 0.135917
R5632 VPWR.n1072 VPWR 0.135917
R5633 VPWR.n1075 VPWR 0.135917
R5634 VPWR.n1685 VPWR 0.135917
R5635 VPWR.n1083 VPWR 0.135917
R5636 VPWR.n1085 VPWR 0.135917
R5637 VPWR.n1658 VPWR 0.135917
R5638 VPWR.n1093 VPWR 0.135917
R5639 VPWR.n1095 VPWR 0.135917
R5640 VPWR.n1631 VPWR 0.135917
R5641 VPWR.n1103 VPWR 0.135917
R5642 VPWR.n1105 VPWR 0.135917
R5643 VPWR.n1604 VPWR 0.135917
R5644 VPWR.n2863 VPWR.n2814 0.127988
R5645 VPWR.n2825 VPWR.n2816 0.1255
R5646 VPWR.n2831 VPWR.n2816 0.1255
R5647 VPWR.n18 VPWR.n0 0.120292
R5648 VPWR.n14 VPWR.n0 0.120292
R5649 VPWR.n9 VPWR.n8 0.120292
R5650 VPWR.n1254 VPWR.n1233 0.120292
R5651 VPWR.n1250 VPWR.n1233 0.120292
R5652 VPWR.n1244 VPWR.n1243 0.120292
R5653 VPWR.n1278 VPWR.n1256 0.120292
R5654 VPWR.n1273 VPWR.n1256 0.120292
R5655 VPWR.n1267 VPWR.n1266 0.120292
R5656 VPWR.n1301 VPWR.n1280 0.120292
R5657 VPWR.n1297 VPWR.n1280 0.120292
R5658 VPWR.n1291 VPWR.n1290 0.120292
R5659 VPWR.n1333 VPWR.n1332 0.120292
R5660 VPWR.n1326 VPWR.n1305 0.120292
R5661 VPWR.n1319 VPWR.n1305 0.120292
R5662 VPWR.n1319 VPWR.n1318 0.120292
R5663 VPWR.n1317 VPWR.n1309 0.120292
R5664 VPWR.n1312 VPWR.n1309 0.120292
R5665 VPWR.n1312 VPWR.n1311 0.120292
R5666 VPWR.n1371 VPWR.n1370 0.120292
R5667 VPWR.n1364 VPWR.n1363 0.120292
R5668 VPWR.n1363 VPWR.n1340 0.120292
R5669 VPWR.n1356 VPWR.n1340 0.120292
R5670 VPWR.n1356 VPWR.n1355 0.120292
R5671 VPWR.n1355 VPWR.n1354 0.120292
R5672 VPWR.n1354 VPWR.n1342 0.120292
R5673 VPWR.n1348 VPWR.n1342 0.120292
R5674 VPWR.n1348 VPWR.n1347 0.120292
R5675 VPWR.n1410 VPWR.n1409 0.120292
R5676 VPWR.n1403 VPWR.n1402 0.120292
R5677 VPWR.n1402 VPWR.n1379 0.120292
R5678 VPWR.n1395 VPWR.n1379 0.120292
R5679 VPWR.n1395 VPWR.n1394 0.120292
R5680 VPWR.n1394 VPWR.n1393 0.120292
R5681 VPWR.n1393 VPWR.n1381 0.120292
R5682 VPWR.n1387 VPWR.n1381 0.120292
R5683 VPWR.n1387 VPWR.n1386 0.120292
R5684 VPWR.n1440 VPWR.n1439 0.120292
R5685 VPWR.n1439 VPWR.n1416 0.120292
R5686 VPWR.n1432 VPWR.n1416 0.120292
R5687 VPWR.n1432 VPWR.n1431 0.120292
R5688 VPWR.n1431 VPWR.n1430 0.120292
R5689 VPWR.n1430 VPWR.n1418 0.120292
R5690 VPWR.n1424 VPWR.n1418 0.120292
R5691 VPWR.n1424 VPWR.n1423 0.120292
R5692 VPWR.n2812 VPWR.n2798 0.120292
R5693 VPWR.n2796 VPWR.n2779 0.120292
R5694 VPWR.n2777 VPWR.n2759 0.120292
R5695 VPWR.n2757 VPWR.n2740 0.120292
R5696 VPWR.n2719 VPWR.n2718 0.120292
R5697 VPWR.n2720 VPWR.n2719 0.120292
R5698 VPWR.n2720 VPWR.n2711 0.120292
R5699 VPWR.n2725 VPWR.n2711 0.120292
R5700 VPWR.n2726 VPWR.n2725 0.120292
R5701 VPWR.n2726 VPWR.n2707 0.120292
R5702 VPWR.n2732 VPWR.n2707 0.120292
R5703 VPWR.n2734 VPWR.n2704 0.120292
R5704 VPWR.n2738 VPWR.n2704 0.120292
R5705 VPWR.n2683 VPWR.n2682 0.120292
R5706 VPWR.n2684 VPWR.n2683 0.120292
R5707 VPWR.n2684 VPWR.n2673 0.120292
R5708 VPWR.n2689 VPWR.n2673 0.120292
R5709 VPWR.n2690 VPWR.n2689 0.120292
R5710 VPWR.n2690 VPWR.n2669 0.120292
R5711 VPWR.n2695 VPWR.n2669 0.120292
R5712 VPWR.n2697 VPWR.n2666 0.120292
R5713 VPWR.n2702 VPWR.n2666 0.120292
R5714 VPWR.n2646 VPWR.n2645 0.120292
R5715 VPWR.n2647 VPWR.n2646 0.120292
R5716 VPWR.n2647 VPWR.n2636 0.120292
R5717 VPWR.n2652 VPWR.n2636 0.120292
R5718 VPWR.n2653 VPWR.n2652 0.120292
R5719 VPWR.n2653 VPWR.n2632 0.120292
R5720 VPWR.n2658 VPWR.n2632 0.120292
R5721 VPWR.n2660 VPWR.n2629 0.120292
R5722 VPWR.n2664 VPWR.n2629 0.120292
R5723 VPWR.n2608 VPWR.n2604 0.120292
R5724 VPWR.n2616 VPWR.n2604 0.120292
R5725 VPWR.n2617 VPWR.n2616 0.120292
R5726 VPWR.n2618 VPWR.n2617 0.120292
R5727 VPWR.n2618 VPWR.n2600 0.120292
R5728 VPWR.n2623 VPWR.n2600 0.120292
R5729 VPWR.n2624 VPWR.n2623 0.120292
R5730 VPWR.n1605 VPWR 0.118556
R5731 VPWR.n1108 VPWR 0.118556
R5732 VPWR.n1619 VPWR 0.118556
R5733 VPWR.n1632 VPWR 0.118556
R5734 VPWR.n1098 VPWR 0.118556
R5735 VPWR.n1646 VPWR 0.118556
R5736 VPWR.n1659 VPWR 0.118556
R5737 VPWR.n1088 VPWR 0.118556
R5738 VPWR.n1673 VPWR 0.118556
R5739 VPWR.n1686 VPWR 0.118556
R5740 VPWR.n1078 VPWR 0.118556
R5741 VPWR.n1700 VPWR 0.118556
R5742 VPWR.n1713 VPWR 0.118556
R5743 VPWR.n1725 VPWR 0.118556
R5744 VPWR VPWR.n1112 0.118556
R5745 VPWR.n1067 VPWR 0.118556
R5746 VPWR.n123 VPWR 0.118556
R5747 VPWR.n112 VPWR 0.118556
R5748 VPWR.n103 VPWR 0.118556
R5749 VPWR.n278 VPWR 0.118556
R5750 VPWR.n266 VPWR 0.118556
R5751 VPWR.n254 VPWR 0.118556
R5752 VPWR.n242 VPWR 0.118556
R5753 VPWR.n230 VPWR 0.118556
R5754 VPWR.n218 VPWR 0.118556
R5755 VPWR.n206 VPWR 0.118556
R5756 VPWR.n194 VPWR 0.118556
R5757 VPWR.n182 VPWR 0.118556
R5758 VPWR.n170 VPWR 0.118556
R5759 VPWR.n158 VPWR 0.118556
R5760 VPWR.n146 VPWR 0.118556
R5761 VPWR.n134 VPWR 0.118556
R5762 VPWR.n1765 VPWR.n1044 0.108238
R5763 VPWR.n1541 VPWR.n1143 0.108238
R5764 VPWR.n1540 VPWR.n1142 0.108238
R5765 VPWR.n1524 VPWR.n1141 0.108238
R5766 VPWR.n1516 VPWR.n1140 0.108238
R5767 VPWR.n1510 VPWR.n1139 0.108238
R5768 VPWR.n1502 VPWR.n1138 0.108238
R5769 VPWR.n1496 VPWR.n1137 0.108238
R5770 VPWR.n1583 VPWR.n1132 0.108238
R5771 VPWR.n1584 VPWR.n1131 0.108238
R5772 VPWR.n1463 VPWR.n1452 0.108238
R5773 VPWR.n1464 VPWR.n1451 0.108238
R5774 VPWR.n1795 VPWR.n1027 0.108238
R5775 VPWR.n1766 VPWR.n1043 0.108238
R5776 VPWR.n1744 VPWR.n1038 0.108238
R5777 VPWR.n1787 VPWR.n1786 0.108238
R5778 VPWR.n2481 VPWR 0.100405
R5779 VPWR.n2472 VPWR 0.100405
R5780 VPWR VPWR.n2385 0.100405
R5781 VPWR VPWR.n2386 0.100405
R5782 VPWR VPWR.n2387 0.100405
R5783 VPWR.n2305 VPWR 0.100405
R5784 VPWR VPWR.n2314 0.100405
R5785 VPWR.n2315 VPWR 0.100405
R5786 VPWR VPWR.n2324 0.100405
R5787 VPWR.n2375 VPWR 0.100405
R5788 VPWR VPWR.n2374 0.100405
R5789 VPWR.n2365 VPWR 0.100405
R5790 VPWR VPWR.n2364 0.100405
R5791 VPWR.n2355 VPWR 0.100405
R5792 VPWR VPWR.n2354 0.100405
R5793 VPWR.n2345 VPWR 0.100405
R5794 VPWR VPWR.n2344 0.100405
R5795 VPWR.n2335 VPWR 0.100405
R5796 VPWR VPWR.n2334 0.100405
R5797 VPWR.n2325 VPWR 0.100405
R5798 VPWR.n2302 VPWR 0.100405
R5799 VPWR.n2301 VPWR 0.100405
R5800 VPWR.n2300 VPWR 0.100405
R5801 VPWR.n2299 VPWR 0.100405
R5802 VPWR.n2288 VPWR 0.100405
R5803 VPWR.n2289 VPWR 0.100405
R5804 VPWR.n2290 VPWR 0.100405
R5805 VPWR.n2291 VPWR 0.100405
R5806 VPWR.n2292 VPWR 0.100405
R5807 VPWR.n2293 VPWR 0.100405
R5808 VPWR.n2294 VPWR 0.100405
R5809 VPWR.n2295 VPWR 0.100405
R5810 VPWR.n2296 VPWR 0.100405
R5811 VPWR.n2297 VPWR 0.100405
R5812 VPWR.n2298 VPWR 0.100405
R5813 VPWR.n2285 VPWR 0.100405
R5814 VPWR.n2276 VPWR 0.100405
R5815 VPWR.n2275 VPWR 0.100405
R5816 VPWR.n2266 VPWR 0.100405
R5817 VPWR.n2215 VPWR 0.100405
R5818 VPWR.n2216 VPWR 0.100405
R5819 VPWR.n2225 VPWR 0.100405
R5820 VPWR.n2226 VPWR 0.100405
R5821 VPWR.n2235 VPWR 0.100405
R5822 VPWR.n2236 VPWR 0.100405
R5823 VPWR.n2245 VPWR 0.100405
R5824 VPWR.n2246 VPWR 0.100405
R5825 VPWR.n2255 VPWR 0.100405
R5826 VPWR.n2256 VPWR 0.100405
R5827 VPWR.n2265 VPWR 0.100405
R5828 VPWR VPWR.n2189 0.100405
R5829 VPWR VPWR.n2190 0.100405
R5830 VPWR VPWR.n2191 0.100405
R5831 VPWR VPWR.n2192 0.100405
R5832 VPWR VPWR.n2203 0.100405
R5833 VPWR VPWR.n2202 0.100405
R5834 VPWR VPWR.n2201 0.100405
R5835 VPWR VPWR.n2200 0.100405
R5836 VPWR VPWR.n2199 0.100405
R5837 VPWR VPWR.n2198 0.100405
R5838 VPWR VPWR.n2197 0.100405
R5839 VPWR VPWR.n2196 0.100405
R5840 VPWR VPWR.n2195 0.100405
R5841 VPWR VPWR.n2194 0.100405
R5842 VPWR VPWR.n2193 0.100405
R5843 VPWR.n2109 VPWR 0.100405
R5844 VPWR VPWR.n2118 0.100405
R5845 VPWR.n2119 VPWR 0.100405
R5846 VPWR VPWR.n2128 0.100405
R5847 VPWR.n2179 VPWR 0.100405
R5848 VPWR VPWR.n2178 0.100405
R5849 VPWR.n2169 VPWR 0.100405
R5850 VPWR VPWR.n2168 0.100405
R5851 VPWR.n2159 VPWR 0.100405
R5852 VPWR VPWR.n2158 0.100405
R5853 VPWR.n2149 VPWR 0.100405
R5854 VPWR VPWR.n2148 0.100405
R5855 VPWR.n2139 VPWR 0.100405
R5856 VPWR VPWR.n2138 0.100405
R5857 VPWR.n2129 VPWR 0.100405
R5858 VPWR.n2106 VPWR 0.100405
R5859 VPWR.n2105 VPWR 0.100405
R5860 VPWR.n2104 VPWR 0.100405
R5861 VPWR.n2103 VPWR 0.100405
R5862 VPWR.n2092 VPWR 0.100405
R5863 VPWR.n2093 VPWR 0.100405
R5864 VPWR.n2094 VPWR 0.100405
R5865 VPWR.n2095 VPWR 0.100405
R5866 VPWR.n2096 VPWR 0.100405
R5867 VPWR.n2097 VPWR 0.100405
R5868 VPWR.n2098 VPWR 0.100405
R5869 VPWR.n2099 VPWR 0.100405
R5870 VPWR.n2100 VPWR 0.100405
R5871 VPWR.n2101 VPWR 0.100405
R5872 VPWR.n2102 VPWR 0.100405
R5873 VPWR.n2089 VPWR 0.100405
R5874 VPWR.n2080 VPWR 0.100405
R5875 VPWR.n2079 VPWR 0.100405
R5876 VPWR.n2070 VPWR 0.100405
R5877 VPWR.n2019 VPWR 0.100405
R5878 VPWR.n2020 VPWR 0.100405
R5879 VPWR.n2029 VPWR 0.100405
R5880 VPWR.n2030 VPWR 0.100405
R5881 VPWR.n2039 VPWR 0.100405
R5882 VPWR.n2040 VPWR 0.100405
R5883 VPWR.n2049 VPWR 0.100405
R5884 VPWR.n2050 VPWR 0.100405
R5885 VPWR.n2059 VPWR 0.100405
R5886 VPWR.n2060 VPWR 0.100405
R5887 VPWR.n2069 VPWR 0.100405
R5888 VPWR VPWR.n1993 0.100405
R5889 VPWR VPWR.n1994 0.100405
R5890 VPWR VPWR.n1995 0.100405
R5891 VPWR VPWR.n1996 0.100405
R5892 VPWR VPWR.n2007 0.100405
R5893 VPWR VPWR.n2006 0.100405
R5894 VPWR VPWR.n2005 0.100405
R5895 VPWR VPWR.n2004 0.100405
R5896 VPWR VPWR.n2003 0.100405
R5897 VPWR VPWR.n2002 0.100405
R5898 VPWR VPWR.n2001 0.100405
R5899 VPWR VPWR.n2000 0.100405
R5900 VPWR VPWR.n1999 0.100405
R5901 VPWR VPWR.n1998 0.100405
R5902 VPWR VPWR.n1997 0.100405
R5903 VPWR.n1913 VPWR 0.100405
R5904 VPWR VPWR.n1922 0.100405
R5905 VPWR.n1923 VPWR 0.100405
R5906 VPWR VPWR.n1932 0.100405
R5907 VPWR.n1983 VPWR 0.100405
R5908 VPWR VPWR.n1982 0.100405
R5909 VPWR.n1973 VPWR 0.100405
R5910 VPWR VPWR.n1972 0.100405
R5911 VPWR.n1963 VPWR 0.100405
R5912 VPWR VPWR.n1962 0.100405
R5913 VPWR.n1953 VPWR 0.100405
R5914 VPWR VPWR.n1952 0.100405
R5915 VPWR.n1943 VPWR 0.100405
R5916 VPWR VPWR.n1942 0.100405
R5917 VPWR.n1933 VPWR 0.100405
R5918 VPWR.n1910 VPWR 0.100405
R5919 VPWR.n1909 VPWR 0.100405
R5920 VPWR.n1908 VPWR 0.100405
R5921 VPWR.n1907 VPWR 0.100405
R5922 VPWR.n1896 VPWR 0.100405
R5923 VPWR.n1897 VPWR 0.100405
R5924 VPWR.n1898 VPWR 0.100405
R5925 VPWR.n1899 VPWR 0.100405
R5926 VPWR.n1900 VPWR 0.100405
R5927 VPWR.n1901 VPWR 0.100405
R5928 VPWR.n1902 VPWR 0.100405
R5929 VPWR.n1903 VPWR 0.100405
R5930 VPWR.n1904 VPWR 0.100405
R5931 VPWR.n1905 VPWR 0.100405
R5932 VPWR.n1906 VPWR 0.100405
R5933 VPWR VPWR.n2399 0.100405
R5934 VPWR VPWR.n2398 0.100405
R5935 VPWR VPWR.n2397 0.100405
R5936 VPWR VPWR.n2396 0.100405
R5937 VPWR VPWR.n2395 0.100405
R5938 VPWR VPWR.n2394 0.100405
R5939 VPWR VPWR.n2393 0.100405
R5940 VPWR VPWR.n2392 0.100405
R5941 VPWR VPWR.n2391 0.100405
R5942 VPWR VPWR.n2390 0.100405
R5943 VPWR VPWR.n2389 0.100405
R5944 VPWR VPWR.n2388 0.100405
R5945 VPWR.n1893 VPWR 0.100405
R5946 VPWR.n1884 VPWR 0.100405
R5947 VPWR.n1883 VPWR 0.100405
R5948 VPWR.n1874 VPWR 0.100405
R5949 VPWR.n1873 VPWR 0.100405
R5950 VPWR.n1823 VPWR 0.100405
R5951 VPWR.n1824 VPWR 0.100405
R5952 VPWR.n1833 VPWR 0.100405
R5953 VPWR.n1834 VPWR 0.100405
R5954 VPWR.n1843 VPWR 0.100405
R5955 VPWR.n1844 VPWR 0.100405
R5956 VPWR.n1853 VPWR 0.100405
R5957 VPWR.n1854 VPWR 0.100405
R5958 VPWR.n1863 VPWR 0.100405
R5959 VPWR.n1864 VPWR 0.100405
R5960 VPWR.n2411 VPWR 0.100405
R5961 VPWR.n2412 VPWR 0.100405
R5962 VPWR.n2421 VPWR 0.100405
R5963 VPWR.n2422 VPWR 0.100405
R5964 VPWR.n2431 VPWR 0.100405
R5965 VPWR.n2432 VPWR 0.100405
R5966 VPWR.n2441 VPWR 0.100405
R5967 VPWR.n2442 VPWR 0.100405
R5968 VPWR.n2451 VPWR 0.100405
R5969 VPWR.n2452 VPWR 0.100405
R5970 VPWR.n2461 VPWR 0.100405
R5971 VPWR.n2462 VPWR 0.100405
R5972 VPWR.n2471 VPWR 0.100405
R5973 VPWR VPWR.n1797 0.100405
R5974 VPWR VPWR.n1798 0.100405
R5975 VPWR VPWR.n1799 0.100405
R5976 VPWR VPWR.n1800 0.100405
R5977 VPWR VPWR.n1801 0.100405
R5978 VPWR VPWR.n1802 0.100405
R5979 VPWR VPWR.n1803 0.100405
R5980 VPWR VPWR.n1804 0.100405
R5981 VPWR VPWR.n1811 0.100405
R5982 VPWR VPWR.n1810 0.100405
R5983 VPWR VPWR.n1809 0.100405
R5984 VPWR VPWR.n1808 0.100405
R5985 VPWR VPWR.n1807 0.100405
R5986 VPWR VPWR.n1806 0.100405
R5987 VPWR VPWR.n1805 0.100405
R5988 VPWR.n2498 VPWR 0.100405
R5989 VPWR.n2497 VPWR 0.100405
R5990 VPWR.n2496 VPWR 0.100405
R5991 VPWR.n2495 VPWR 0.100405
R5992 VPWR.n2494 VPWR 0.100405
R5993 VPWR.n2493 VPWR 0.100405
R5994 VPWR.n2492 VPWR 0.100405
R5995 VPWR.n2491 VPWR 0.100405
R5996 VPWR.n2490 VPWR 0.100405
R5997 VPWR.n2489 VPWR 0.100405
R5998 VPWR.n2484 VPWR 0.100405
R5999 VPWR.n2485 VPWR 0.100405
R6000 VPWR.n2486 VPWR 0.100405
R6001 VPWR.n2487 VPWR 0.100405
R6002 VPWR.n2488 VPWR 0.100405
R6003 VPWR.n1143 VPWR 0.100405
R6004 VPWR VPWR.n1540 0.100405
R6005 VPWR.n1524 VPWR 0.100405
R6006 VPWR.n1516 VPWR 0.100405
R6007 VPWR.n1510 VPWR 0.100405
R6008 VPWR.n1502 VPWR 0.100405
R6009 VPWR.n1496 VPWR 0.100405
R6010 VPWR VPWR.n1132 0.100405
R6011 VPWR.n1584 VPWR 0.100405
R6012 VPWR.n1452 VPWR 0.100405
R6013 VPWR.n1464 VPWR 0.100405
R6014 VPWR.n1043 VPWR 0.100405
R6015 VPWR.n1744 VPWR 0.100405
R6016 VPWR.n1787 VPWR 0.100405
R6017 VPWR VPWR.n1765 0.100405
R6018 VPWR.n2501 VPWR 0.100405
R6019 VPWR VPWR.n2512 0.100405
R6020 VPWR.n2513 VPWR 0.100405
R6021 VPWR VPWR.n2524 0.100405
R6022 VPWR.n2525 VPWR 0.100405
R6023 VPWR VPWR.n2536 0.100405
R6024 VPWR.n2537 VPWR 0.100405
R6025 VPWR VPWR.n2548 0.100405
R6026 VPWR.n2549 VPWR 0.100405
R6027 VPWR VPWR.n2560 0.100405
R6028 VPWR.n2561 VPWR 0.100405
R6029 VPWR VPWR.n2572 0.100405
R6030 VPWR.n2573 VPWR 0.100405
R6031 VPWR VPWR.n2584 0.100405
R6032 VPWR.n2585 VPWR 0.100405
R6033 VPWR.n1056 VPWR 0.100405
R6034 VPWR.n1754 VPWR 0.100405
R6035 VPWR.n1755 VPWR 0.100405
R6036 VPWR.n1529 VPWR 0.100405
R6037 VPWR.n1530 VPWR 0.100405
R6038 VPWR VPWR.n1528 0.100405
R6039 VPWR VPWR.n1527 0.100405
R6040 VPWR.n1514 VPWR 0.100405
R6041 VPWR VPWR.n1513 0.100405
R6042 VPWR.n1500 VPWR 0.100405
R6043 VPWR VPWR.n1499 0.100405
R6044 VPWR.n1487 VPWR 0.100405
R6045 VPWR.n1587 VPWR 0.100405
R6046 VPWR.n1588 VPWR 0.100405
R6047 VPWR.n1448 VPWR 0.100405
R6048 VPWR VPWR.n2798 0.0994583
R6049 VPWR VPWR.n2779 0.0994583
R6050 VPWR VPWR.n1326 0.0981562
R6051 VPWR.n1371 VPWR 0.0981562
R6052 VPWR.n1410 VPWR 0.0981562
R6053 VPWR.n9 VPWR 0.0968542
R6054 VPWR.n1244 VPWR 0.0968542
R6055 VPWR.n1267 VPWR 0.0968542
R6056 VPWR.n1291 VPWR 0.0968542
R6057 VPWR.n1333 VPWR 0.0968542
R6058 VPWR VPWR.n2759 0.0968542
R6059 VPWR VPWR.n2740 0.0968542
R6060 VPWR.n2718 VPWR 0.0968542
R6061 VPWR.n2682 VPWR 0.0968542
R6062 VPWR.n2645 VPWR 0.0968542
R6063 VPWR.n2608 VPWR 0.0968542
R6064 VPWR VPWR.n1044 0.0945
R6065 VPWR.n1541 VPWR 0.0945
R6066 VPWR VPWR.n1142 0.0945
R6067 VPWR VPWR.n1141 0.0945
R6068 VPWR VPWR.n1140 0.0945
R6069 VPWR VPWR.n1139 0.0945
R6070 VPWR VPWR.n1138 0.0945
R6071 VPWR.n1137 VPWR 0.0945
R6072 VPWR VPWR.n1583 0.0945
R6073 VPWR VPWR.n1131 0.0945
R6074 VPWR VPWR.n1463 0.0945
R6075 VPWR.n1451 VPWR 0.0945
R6076 VPWR VPWR.n1038 0.0945
R6077 VPWR.n1786 VPWR 0.0945
R6078 VPWR VPWR.n1027 0.0945
R6079 VPWR.n1766 VPWR 0.0945
R6080 VPWR.n1117 VPWR 0.093504
R6081 VPWR.n109 VPWR 0.093504
R6082 VPWR.n143 VPWR 0.093504
R6083 VPWR.n155 VPWR 0.093504
R6084 VPWR.n167 VPWR 0.093504
R6085 VPWR.n179 VPWR 0.093504
R6086 VPWR.n191 VPWR 0.093504
R6087 VPWR.n203 VPWR 0.093504
R6088 VPWR.n215 VPWR 0.093504
R6089 VPWR.n227 VPWR 0.093504
R6090 VPWR.n239 VPWR 0.093504
R6091 VPWR.n251 VPWR 0.093504
R6092 VPWR.n263 VPWR 0.093504
R6093 VPWR.n275 VPWR 0.093504
R6094 VPWR VPWR.n285 0.093504
R6095 VPWR.n131 VPWR 0.093504
R6096 VPWR.n120 VPWR 0.093504
R6097 VPWR VPWR.n1731 0.093504
R6098 VPWR.n1722 VPWR 0.093504
R6099 VPWR.n1710 VPWR 0.093504
R6100 VPWR.n1699 VPWR 0.093504
R6101 VPWR VPWR.n1077 0.093504
R6102 VPWR.n1683 VPWR 0.093504
R6103 VPWR.n1672 VPWR 0.093504
R6104 VPWR VPWR.n1087 0.093504
R6105 VPWR.n1656 VPWR 0.093504
R6106 VPWR.n1645 VPWR 0.093504
R6107 VPWR VPWR.n1097 0.093504
R6108 VPWR.n1629 VPWR 0.093504
R6109 VPWR.n1618 VPWR 0.093504
R6110 VPWR VPWR.n1107 0.093504
R6111 VPWR.n1602 VPWR 0.093504
R6112 VPWR.n2598 VPWR 0.0849042
R6113 VPWR.n1112 VPWR.n1109 0.0845517
R6114 VPWR.n147 VPWR.n146 0.0845517
R6115 VPWR.n159 VPWR.n158 0.0845517
R6116 VPWR.n171 VPWR.n170 0.0845517
R6117 VPWR.n183 VPWR.n182 0.0845517
R6118 VPWR.n195 VPWR.n194 0.0845517
R6119 VPWR.n207 VPWR.n206 0.0845517
R6120 VPWR.n219 VPWR.n218 0.0845517
R6121 VPWR.n231 VPWR.n230 0.0845517
R6122 VPWR.n243 VPWR.n242 0.0845517
R6123 VPWR.n255 VPWR.n254 0.0845517
R6124 VPWR.n267 VPWR.n266 0.0845517
R6125 VPWR.n279 VPWR.n278 0.0845517
R6126 VPWR.n282 VPWR.n103 0.0845517
R6127 VPWR.n113 VPWR.n112 0.0845517
R6128 VPWR.n135 VPWR.n134 0.0845517
R6129 VPWR.n124 VPWR.n123 0.0845517
R6130 VPWR.n1728 VPWR.n1067 0.0845517
R6131 VPWR.n1726 VPWR.n1725 0.0845517
R6132 VPWR.n1714 VPWR.n1713 0.0845517
R6133 VPWR.n1701 VPWR.n1700 0.0845517
R6134 VPWR.n1690 VPWR.n1078 0.0845517
R6135 VPWR.n1687 VPWR.n1686 0.0845517
R6136 VPWR.n1674 VPWR.n1673 0.0845517
R6137 VPWR.n1663 VPWR.n1088 0.0845517
R6138 VPWR.n1660 VPWR.n1659 0.0845517
R6139 VPWR.n1647 VPWR.n1646 0.0845517
R6140 VPWR.n1636 VPWR.n1098 0.0845517
R6141 VPWR.n1633 VPWR.n1632 0.0845517
R6142 VPWR.n1620 VPWR.n1619 0.0845517
R6143 VPWR.n1609 VPWR.n1108 0.0845517
R6144 VPWR.n1606 VPWR.n1605 0.0845517
R6145 VPWR.n1456 VPWR.n1451 0.0740128
R6146 VPWR.n1542 VPWR.n1044 0.071
R6147 VPWR.n1547 VPWR.n1541 0.071
R6148 VPWR.n1552 VPWR.n1142 0.071
R6149 VPWR.n1557 VPWR.n1141 0.071
R6150 VPWR.n1562 VPWR.n1140 0.071
R6151 VPWR.n1567 VPWR.n1139 0.071
R6152 VPWR.n1572 VPWR.n1138 0.071
R6153 VPWR.n1577 VPWR.n1137 0.071
R6154 VPWR.n1583 VPWR.n1582 0.071
R6155 VPWR.n1457 VPWR.n1131 0.071
R6156 VPWR.n1463 VPWR.n1462 0.071
R6157 VPWR.n1772 VPWR.n1038 0.071
R6158 VPWR.n1786 VPWR.n1785 0.071
R6159 VPWR.n1780 VPWR.n1027 0.071
R6160 VPWR.n1767 VPWR.n1766 0.071
R6161 VPWR VPWR.n1115 0.0678077
R6162 VPWR VPWR.n107 0.0678077
R6163 VPWR VPWR.n141 0.0678077
R6164 VPWR VPWR.n153 0.0678077
R6165 VPWR VPWR.n165 0.0678077
R6166 VPWR VPWR.n177 0.0678077
R6167 VPWR VPWR.n189 0.0678077
R6168 VPWR VPWR.n201 0.0678077
R6169 VPWR VPWR.n213 0.0678077
R6170 VPWR VPWR.n225 0.0678077
R6171 VPWR VPWR.n237 0.0678077
R6172 VPWR VPWR.n249 0.0678077
R6173 VPWR VPWR.n261 0.0678077
R6174 VPWR VPWR.n273 0.0678077
R6175 VPWR.n286 VPWR 0.0678077
R6176 VPWR VPWR.n129 0.0678077
R6177 VPWR VPWR.n118 0.0678077
R6178 VPWR.n1732 VPWR 0.0678077
R6179 VPWR VPWR.n1720 0.0678077
R6180 VPWR VPWR.n1708 0.0678077
R6181 VPWR VPWR.n1697 0.0678077
R6182 VPWR.n1193 VPWR 0.0678077
R6183 VPWR VPWR.n1681 0.0678077
R6184 VPWR VPWR.n1670 0.0678077
R6185 VPWR.n1207 VPWR 0.0678077
R6186 VPWR VPWR.n1654 0.0678077
R6187 VPWR VPWR.n1643 0.0678077
R6188 VPWR.n1175 VPWR 0.0678077
R6189 VPWR VPWR.n1627 0.0678077
R6190 VPWR VPWR.n1616 0.0678077
R6191 VPWR.n1124 VPWR 0.0678077
R6192 VPWR VPWR.n1600 0.0678077
R6193 VPWR.n150 VPWR 0.063
R6194 VPWR.n162 VPWR 0.063
R6195 VPWR.n174 VPWR 0.063
R6196 VPWR.n186 VPWR 0.063
R6197 VPWR.n198 VPWR 0.063
R6198 VPWR.n210 VPWR 0.063
R6199 VPWR.n222 VPWR 0.063
R6200 VPWR.n234 VPWR 0.063
R6201 VPWR.n246 VPWR 0.063
R6202 VPWR.n258 VPWR 0.063
R6203 VPWR.n270 VPWR 0.063
R6204 VPWR.n101 VPWR 0.063
R6205 VPWR.n105 VPWR 0.063
R6206 VPWR.n138 VPWR 0.063
R6207 VPWR.n115 VPWR 0.063
R6208 VPWR.n126 VPWR 0.063
R6209 VPWR.n1065 VPWR 0.063
R6210 VPWR.n1717 VPWR 0.063
R6211 VPWR.n1070 VPWR 0.063
R6212 VPWR VPWR.n1704 0.063
R6213 VPWR VPWR.n1693 0.063
R6214 VPWR VPWR.n1081 0.063
R6215 VPWR VPWR.n1677 0.063
R6216 VPWR VPWR.n1666 0.063
R6217 VPWR VPWR.n1091 0.063
R6218 VPWR VPWR.n1650 0.063
R6219 VPWR VPWR.n1639 0.063
R6220 VPWR VPWR.n1101 0.063
R6221 VPWR VPWR.n1623 0.063
R6222 VPWR VPWR.n1612 0.063
R6223 VPWR VPWR.n1111 0.063
R6224 VPWR VPWR.n1120 0.063
R6225 VPWR.n1115 VPWR 0.0608448
R6226 VPWR.n107 VPWR 0.0608448
R6227 VPWR.n141 VPWR 0.0608448
R6228 VPWR.n153 VPWR 0.0608448
R6229 VPWR.n165 VPWR 0.0608448
R6230 VPWR.n177 VPWR 0.0608448
R6231 VPWR.n189 VPWR 0.0608448
R6232 VPWR.n201 VPWR 0.0608448
R6233 VPWR.n213 VPWR 0.0608448
R6234 VPWR.n225 VPWR 0.0608448
R6235 VPWR.n237 VPWR 0.0608448
R6236 VPWR.n249 VPWR 0.0608448
R6237 VPWR.n261 VPWR 0.0608448
R6238 VPWR.n273 VPWR 0.0608448
R6239 VPWR.n286 VPWR 0.0608448
R6240 VPWR.n129 VPWR 0.0608448
R6241 VPWR.n118 VPWR 0.0608448
R6242 VPWR.n1732 VPWR 0.0608448
R6243 VPWR.n1720 VPWR 0.0608448
R6244 VPWR.n1708 VPWR 0.0608448
R6245 VPWR.n1697 VPWR 0.0608448
R6246 VPWR.n1193 VPWR 0.0608448
R6247 VPWR.n1681 VPWR 0.0608448
R6248 VPWR.n1670 VPWR 0.0608448
R6249 VPWR.n1207 VPWR 0.0608448
R6250 VPWR.n1654 VPWR 0.0608448
R6251 VPWR.n1643 VPWR 0.0608448
R6252 VPWR.n1175 VPWR 0.0608448
R6253 VPWR.n1627 VPWR 0.0608448
R6254 VPWR.n1616 VPWR 0.0608448
R6255 VPWR.n1124 VPWR 0.0608448
R6256 VPWR.n1600 VPWR 0.0608448
R6257 VPWR VPWR.n13 0.0603958
R6258 VPWR VPWR.n12 0.0603958
R6259 VPWR VPWR.n1249 0.0603958
R6260 VPWR VPWR.n1248 0.0603958
R6261 VPWR VPWR.n1272 0.0603958
R6262 VPWR VPWR.n1271 0.0603958
R6263 VPWR VPWR.n1296 0.0603958
R6264 VPWR VPWR.n1295 0.0603958
R6265 VPWR.n1332 VPWR 0.0603958
R6266 VPWR VPWR.n1331 0.0603958
R6267 VPWR.n1327 VPWR 0.0603958
R6268 VPWR.n1318 VPWR 0.0603958
R6269 VPWR VPWR.n1317 0.0603958
R6270 VPWR.n1370 VPWR 0.0603958
R6271 VPWR VPWR.n1369 0.0603958
R6272 VPWR.n1364 VPWR 0.0603958
R6273 VPWR.n1409 VPWR 0.0603958
R6274 VPWR VPWR.n1408 0.0603958
R6275 VPWR.n1403 VPWR 0.0603958
R6276 VPWR.n1440 VPWR 0.0603958
R6277 VPWR VPWR.n2800 0.0603958
R6278 VPWR VPWR.n2799 0.0603958
R6279 VPWR VPWR.n2812 0.0603958
R6280 VPWR.n2791 VPWR 0.0603958
R6281 VPWR.n2792 VPWR 0.0603958
R6282 VPWR VPWR.n2796 0.0603958
R6283 VPWR.n2771 VPWR 0.0603958
R6284 VPWR.n2772 VPWR 0.0603958
R6285 VPWR VPWR.n2777 0.0603958
R6286 VPWR.n2752 VPWR 0.0603958
R6287 VPWR.n2753 VPWR 0.0603958
R6288 VPWR VPWR.n2757 0.0603958
R6289 VPWR.n2733 VPWR 0.0603958
R6290 VPWR.n2734 VPWR 0.0603958
R6291 VPWR VPWR.n2695 0.0603958
R6292 VPWR.n2696 VPWR 0.0603958
R6293 VPWR.n2697 VPWR 0.0603958
R6294 VPWR VPWR.n2658 0.0603958
R6295 VPWR.n2659 VPWR 0.0603958
R6296 VPWR.n2660 VPWR 0.0603958
R6297 VPWR.n2624 VPWR 0.0603958
R6298 VPWR.n2627 VPWR 0.0603958
R6299 VPWR.n1770 VPWR.n1769 0.0599512
R6300 VPWR.n1041 VPWR.n1040 0.0599512
R6301 VPWR.n1545 VPWR.n1544 0.0599512
R6302 VPWR.n1550 VPWR.n1549 0.0599512
R6303 VPWR.n1555 VPWR.n1554 0.0599512
R6304 VPWR.n1560 VPWR.n1559 0.0599512
R6305 VPWR.n1565 VPWR.n1564 0.0599512
R6306 VPWR.n1570 VPWR.n1569 0.0599512
R6307 VPWR.n1575 VPWR.n1574 0.0599512
R6308 VPWR.n1580 VPWR.n1579 0.0599512
R6309 VPWR.n1135 VPWR.n1134 0.0599512
R6310 VPWR.n1460 VPWR.n1459 0.0599512
R6311 VPWR.n1455 VPWR.n1454 0.0599512
R6312 VPWR.n1775 VPWR.n1774 0.0599512
R6313 VPWR.n1783 VPWR.n1782 0.0599512
R6314 VPWR.n1779 VPWR.n1778 0.0599512
R6315 VPWR.n1118 VPWR.n1117 0.0565345
R6316 VPWR.n1112 VPWR 0.0565345
R6317 VPWR.n144 VPWR.n143 0.0565345
R6318 VPWR.n146 VPWR 0.0565345
R6319 VPWR.n156 VPWR.n155 0.0565345
R6320 VPWR.n158 VPWR 0.0565345
R6321 VPWR.n168 VPWR.n167 0.0565345
R6322 VPWR.n170 VPWR 0.0565345
R6323 VPWR.n180 VPWR.n179 0.0565345
R6324 VPWR.n182 VPWR 0.0565345
R6325 VPWR.n192 VPWR.n191 0.0565345
R6326 VPWR.n194 VPWR 0.0565345
R6327 VPWR.n204 VPWR.n203 0.0565345
R6328 VPWR.n206 VPWR 0.0565345
R6329 VPWR.n216 VPWR.n215 0.0565345
R6330 VPWR.n218 VPWR 0.0565345
R6331 VPWR.n228 VPWR.n227 0.0565345
R6332 VPWR.n230 VPWR 0.0565345
R6333 VPWR.n240 VPWR.n239 0.0565345
R6334 VPWR.n242 VPWR 0.0565345
R6335 VPWR.n252 VPWR.n251 0.0565345
R6336 VPWR.n254 VPWR 0.0565345
R6337 VPWR.n264 VPWR.n263 0.0565345
R6338 VPWR.n266 VPWR 0.0565345
R6339 VPWR.n276 VPWR.n275 0.0565345
R6340 VPWR.n278 VPWR 0.0565345
R6341 VPWR.n285 VPWR.n283 0.0565345
R6342 VPWR.n103 VPWR 0.0565345
R6343 VPWR.n110 VPWR.n109 0.0565345
R6344 VPWR.n112 VPWR 0.0565345
R6345 VPWR.n132 VPWR.n131 0.0565345
R6346 VPWR.n134 VPWR 0.0565345
R6347 VPWR.n121 VPWR.n120 0.0565345
R6348 VPWR.n123 VPWR 0.0565345
R6349 VPWR.n1731 VPWR.n1729 0.0565345
R6350 VPWR.n1067 VPWR 0.0565345
R6351 VPWR.n1723 VPWR.n1722 0.0565345
R6352 VPWR.n1725 VPWR 0.0565345
R6353 VPWR.n1711 VPWR.n1710 0.0565345
R6354 VPWR.n1713 VPWR 0.0565345
R6355 VPWR.n1702 VPWR.n1699 0.0565345
R6356 VPWR.n1700 VPWR 0.0565345
R6357 VPWR.n1691 VPWR.n1077 0.0565345
R6358 VPWR.n1078 VPWR 0.0565345
R6359 VPWR.n1684 VPWR.n1683 0.0565345
R6360 VPWR.n1686 VPWR 0.0565345
R6361 VPWR.n1675 VPWR.n1672 0.0565345
R6362 VPWR.n1673 VPWR 0.0565345
R6363 VPWR.n1664 VPWR.n1087 0.0565345
R6364 VPWR.n1088 VPWR 0.0565345
R6365 VPWR.n1657 VPWR.n1656 0.0565345
R6366 VPWR.n1659 VPWR 0.0565345
R6367 VPWR.n1648 VPWR.n1645 0.0565345
R6368 VPWR.n1646 VPWR 0.0565345
R6369 VPWR.n1637 VPWR.n1097 0.0565345
R6370 VPWR.n1098 VPWR 0.0565345
R6371 VPWR.n1630 VPWR.n1629 0.0565345
R6372 VPWR.n1632 VPWR 0.0565345
R6373 VPWR.n1621 VPWR.n1618 0.0565345
R6374 VPWR.n1619 VPWR 0.0565345
R6375 VPWR.n1610 VPWR.n1107 0.0565345
R6376 VPWR.n1108 VPWR 0.0565345
R6377 VPWR.n1603 VPWR.n1602 0.0565345
R6378 VPWR.n1605 VPWR 0.0565345
R6379 VPWR.n1769 VPWR 0.0469286
R6380 VPWR.n1040 VPWR 0.0469286
R6381 VPWR.n1544 VPWR 0.0469286
R6382 VPWR.n1549 VPWR 0.0469286
R6383 VPWR.n1554 VPWR 0.0469286
R6384 VPWR.n1559 VPWR 0.0469286
R6385 VPWR.n1564 VPWR 0.0469286
R6386 VPWR.n1569 VPWR 0.0469286
R6387 VPWR.n1574 VPWR 0.0469286
R6388 VPWR.n1579 VPWR 0.0469286
R6389 VPWR.n1134 VPWR 0.0469286
R6390 VPWR.n1459 VPWR 0.0469286
R6391 VPWR.n1454 VPWR 0.0469286
R6392 VPWR.n1774 VPWR 0.0469286
R6393 VPWR.n1782 VPWR 0.0469286
R6394 VPWR.n1778 VPWR 0.0469286
R6395 VPWR.n1769 VPWR 0.0401341
R6396 VPWR.n1040 VPWR 0.0401341
R6397 VPWR.n1544 VPWR 0.0401341
R6398 VPWR.n1549 VPWR 0.0401341
R6399 VPWR.n1554 VPWR 0.0401341
R6400 VPWR.n1559 VPWR 0.0401341
R6401 VPWR.n1564 VPWR 0.0401341
R6402 VPWR.n1569 VPWR 0.0401341
R6403 VPWR.n1574 VPWR 0.0401341
R6404 VPWR.n1579 VPWR 0.0401341
R6405 VPWR.n1134 VPWR 0.0401341
R6406 VPWR.n1459 VPWR 0.0401341
R6407 VPWR.n1454 VPWR 0.0401341
R6408 VPWR.n1774 VPWR 0.0401341
R6409 VPWR.n1782 VPWR 0.0401341
R6410 VPWR.n1778 VPWR 0.0401341
R6411 VPWR.n13 VPWR 0.0382604
R6412 VPWR.n1249 VPWR 0.0382604
R6413 VPWR.n1272 VPWR 0.0382604
R6414 VPWR.n1296 VPWR 0.0382604
R6415 VPWR.n1331 VPWR 0.0382604
R6416 VPWR.n1369 VPWR 0.0382604
R6417 VPWR.n1408 VPWR 0.0382604
R6418 VPWR.n1445 VPWR 0.0382604
R6419 VPWR.n20 VPWR 0.0375125
R6420 VPWR.n20 VPWR 0.0373589
R6421 VPWR.n1118 VPWR.n1109 0.0349828
R6422 VPWR.n147 VPWR.n144 0.0349828
R6423 VPWR.n159 VPWR.n156 0.0349828
R6424 VPWR.n171 VPWR.n168 0.0349828
R6425 VPWR.n183 VPWR.n180 0.0349828
R6426 VPWR.n195 VPWR.n192 0.0349828
R6427 VPWR.n207 VPWR.n204 0.0349828
R6428 VPWR.n219 VPWR.n216 0.0349828
R6429 VPWR.n231 VPWR.n228 0.0349828
R6430 VPWR.n243 VPWR.n240 0.0349828
R6431 VPWR.n255 VPWR.n252 0.0349828
R6432 VPWR.n267 VPWR.n264 0.0349828
R6433 VPWR.n279 VPWR.n276 0.0349828
R6434 VPWR.n283 VPWR.n282 0.0349828
R6435 VPWR.n113 VPWR.n110 0.0349828
R6436 VPWR.n135 VPWR.n132 0.0349828
R6437 VPWR.n124 VPWR.n121 0.0349828
R6438 VPWR.n1729 VPWR.n1728 0.0349828
R6439 VPWR.n1726 VPWR.n1723 0.0349828
R6440 VPWR.n1714 VPWR.n1711 0.0349828
R6441 VPWR.n1702 VPWR.n1701 0.0349828
R6442 VPWR.n1691 VPWR.n1690 0.0349828
R6443 VPWR.n1687 VPWR.n1684 0.0349828
R6444 VPWR.n1675 VPWR.n1674 0.0349828
R6445 VPWR.n1664 VPWR.n1663 0.0349828
R6446 VPWR.n1660 VPWR.n1657 0.0349828
R6447 VPWR.n1648 VPWR.n1647 0.0349828
R6448 VPWR.n1637 VPWR.n1636 0.0349828
R6449 VPWR.n1633 VPWR.n1630 0.0349828
R6450 VPWR.n1621 VPWR.n1620 0.0349828
R6451 VPWR.n1610 VPWR.n1609 0.0349828
R6452 VPWR.n1606 VPWR.n1603 0.0349828
R6453 VPWR.n2504 VPWR.n2503 0.0340366
R6454 VPWR.n2570 VPWR.n2569 0.0340366
R6455 VPWR.n2510 VPWR.n2509 0.0340366
R6456 VPWR.n2552 VPWR.n2551 0.0340366
R6457 VPWR.n2546 VPWR.n2545 0.0340366
R6458 VPWR.n2534 VPWR.n2533 0.0340366
R6459 VPWR.n2528 VPWR.n2527 0.0340366
R6460 VPWR.n1223 VPWR.n1222 0.0340366
R6461 VPWR.n2522 VPWR.n2521 0.0340366
R6462 VPWR.n1486 VPWR.n1102 0.0340366
R6463 VPWR.n1174 VPWR.n1094 0.0340366
R6464 VPWR.n2540 VPWR.n2539 0.0340366
R6465 VPWR.n1165 VPWR.n1092 0.0340366
R6466 VPWR.n1211 VPWR.n1164 0.0340366
R6467 VPWR.n2516 VPWR.n2515 0.0340366
R6468 VPWR.n1129 VPWR.n1104 0.0340366
R6469 VPWR.n1155 VPWR.n1084 0.0340366
R6470 VPWR.n2558 VPWR.n2557 0.0340366
R6471 VPWR.n1144 VPWR.n1082 0.0340366
R6472 VPWR.n1591 VPWR.n1590 0.0340366
R6473 VPWR.n2564 VPWR.n2563 0.0340366
R6474 VPWR.n1197 VPWR.n1154 0.0340366
R6475 VPWR.n1074 VPWR.n1073 0.0340366
R6476 VPWR.n1743 VPWR.n1742 0.0340366
R6477 VPWR.n1071 VPWR.n1054 0.0340366
R6478 VPWR.n2576 VPWR.n2575 0.0340366
R6479 VPWR.n2582 VPWR.n2581 0.0340366
R6480 VPWR.n2593 VPWR.n2592 0.0340366
R6481 VPWR.n2588 VPWR.n2587 0.0340366
R6482 VPWR.n1737 VPWR.n1736 0.0340366
R6483 VPWR.n1063 VPWR.n1060 0.0340366
R6484 VPWR.n1596 VPWR.n1121 0.0340366
R6485 VPWR.n2628 VPWR.n2598 0.0320292
R6486 VPWR.n2800 VPWR 0.03175
R6487 VPWR VPWR.n2791 0.03175
R6488 VPWR VPWR.n2771 0.03175
R6489 VPWR VPWR.n2752 0.03175
R6490 VPWR VPWR.n2733 0.03175
R6491 VPWR VPWR.n2696 0.03175
R6492 VPWR VPWR.n2659 0.03175
R6493 VPWR VPWR.n2627 0.03175
R6494 VPWR.n2598 VPWR.n2597 0.0240975
R6495 VPWR.n2597 VPWR.n20 0.0240975
R6496 VPWR.n2814 VPWR 0.024
R6497 VPWR.n14 VPWR 0.0239375
R6498 VPWR.n12 VPWR 0.0239375
R6499 VPWR.n1250 VPWR 0.0239375
R6500 VPWR.n1248 VPWR 0.0239375
R6501 VPWR.n1271 VPWR 0.0239375
R6502 VPWR.n1295 VPWR 0.0239375
R6503 VPWR.n2753 VPWR 0.0239375
R6504 VPWR.n2503 VPWR 0.0233659
R6505 VPWR.n1466 VPWR 0.0233659
R6506 VPWR.n352 VPWR 0.0233659
R6507 VPWR.n2570 VPWR 0.0233659
R6508 VPWR.n1533 VPWR 0.0233659
R6509 VPWR.n347 VPWR 0.0233659
R6510 VPWR.n2510 VPWR 0.0233659
R6511 VPWR.n964 VPWR 0.0233659
R6512 VPWR.n2479 VPWR 0.0233659
R6513 VPWR.n2474 VPWR 0.0233659
R6514 VPWR.n319 VPWR 0.0233659
R6515 VPWR.n2551 VPWR 0.0233659
R6516 VPWR.n972 VPWR 0.0233659
R6517 VPWR.n2444 VPWR 0.0233659
R6518 VPWR.n323 VPWR 0.0233659
R6519 VPWR.n2546 VPWR 0.0233659
R6520 VPWR.n1891 VPWR 0.0233659
R6521 VPWR.n1886 VPWR 0.0233659
R6522 VPWR.n1881 VPWR 0.0233659
R6523 VPWR.n388 VPWR 0.0233659
R6524 VPWR.n392 VPWR 0.0233659
R6525 VPWR.n396 VPWR 0.0233659
R6526 VPWR.n2454 VPWR 0.0233659
R6527 VPWR.n331 VPWR 0.0233659
R6528 VPWR.n2534 VPWR 0.0233659
R6529 VPWR.n1876 VPWR 0.0233659
R6530 VPWR.n404 VPWR 0.0233659
R6531 VPWR.n2459 VPWR 0.0233659
R6532 VPWR.n335 VPWR 0.0233659
R6533 VPWR.n2527 VPWR 0.0233659
R6534 VPWR.n2307 VPWR 0.0233659
R6535 VPWR.n2312 VPWR 0.0233659
R6536 VPWR.n2317 VPWR 0.0233659
R6537 VPWR.n2322 VPWR 0.0233659
R6538 VPWR.n2332 VPWR 0.0233659
R6539 VPWR.n2337 VPWR 0.0233659
R6540 VPWR.n2342 VPWR 0.0233659
R6541 VPWR.n2347 VPWR 0.0233659
R6542 VPWR.n2352 VPWR 0.0233659
R6543 VPWR.n2357 VPWR 0.0233659
R6544 VPWR.n2362 VPWR 0.0233659
R6545 VPWR.n2367 VPWR 0.0233659
R6546 VPWR.n2372 VPWR 0.0233659
R6547 VPWR.n2377 VPWR 0.0233659
R6548 VPWR.n2381 VPWR 0.0233659
R6549 VPWR.n2327 VPWR 0.0233659
R6550 VPWR.n544 VPWR 0.0233659
R6551 VPWR.n539 VPWR 0.0233659
R6552 VPWR.n535 VPWR 0.0233659
R6553 VPWR.n531 VPWR 0.0233659
R6554 VPWR.n523 VPWR 0.0233659
R6555 VPWR.n519 VPWR 0.0233659
R6556 VPWR.n515 VPWR 0.0233659
R6557 VPWR.n511 VPWR 0.0233659
R6558 VPWR.n507 VPWR 0.0233659
R6559 VPWR.n503 VPWR 0.0233659
R6560 VPWR.n499 VPWR 0.0233659
R6561 VPWR.n495 VPWR 0.0233659
R6562 VPWR.n491 VPWR 0.0233659
R6563 VPWR.n487 VPWR 0.0233659
R6564 VPWR.n484 VPWR 0.0233659
R6565 VPWR.n527 VPWR 0.0233659
R6566 VPWR.n2283 VPWR 0.0233659
R6567 VPWR.n2278 VPWR 0.0233659
R6568 VPWR.n2273 VPWR 0.0233659
R6569 VPWR.n2268 VPWR 0.0233659
R6570 VPWR.n2258 VPWR 0.0233659
R6571 VPWR.n2253 VPWR 0.0233659
R6572 VPWR.n2248 VPWR 0.0233659
R6573 VPWR.n2243 VPWR 0.0233659
R6574 VPWR.n2238 VPWR 0.0233659
R6575 VPWR.n2233 VPWR 0.0233659
R6576 VPWR.n2228 VPWR 0.0233659
R6577 VPWR.n2223 VPWR 0.0233659
R6578 VPWR.n2218 VPWR 0.0233659
R6579 VPWR.n2213 VPWR 0.0233659
R6580 VPWR.n2209 VPWR 0.0233659
R6581 VPWR.n2263 VPWR 0.0233659
R6582 VPWR.n580 VPWR 0.0233659
R6583 VPWR.n584 VPWR 0.0233659
R6584 VPWR.n588 VPWR 0.0233659
R6585 VPWR.n592 VPWR 0.0233659
R6586 VPWR.n600 VPWR 0.0233659
R6587 VPWR.n604 VPWR 0.0233659
R6588 VPWR.n608 VPWR 0.0233659
R6589 VPWR.n612 VPWR 0.0233659
R6590 VPWR.n616 VPWR 0.0233659
R6591 VPWR.n620 VPWR 0.0233659
R6592 VPWR.n624 VPWR 0.0233659
R6593 VPWR.n628 VPWR 0.0233659
R6594 VPWR.n632 VPWR 0.0233659
R6595 VPWR.n636 VPWR 0.0233659
R6596 VPWR.n640 VPWR 0.0233659
R6597 VPWR.n596 VPWR 0.0233659
R6598 VPWR.n2111 VPWR 0.0233659
R6599 VPWR.n2116 VPWR 0.0233659
R6600 VPWR.n2121 VPWR 0.0233659
R6601 VPWR.n2126 VPWR 0.0233659
R6602 VPWR.n2136 VPWR 0.0233659
R6603 VPWR.n2141 VPWR 0.0233659
R6604 VPWR.n2146 VPWR 0.0233659
R6605 VPWR.n2151 VPWR 0.0233659
R6606 VPWR.n2156 VPWR 0.0233659
R6607 VPWR.n2161 VPWR 0.0233659
R6608 VPWR.n2166 VPWR 0.0233659
R6609 VPWR.n2171 VPWR 0.0233659
R6610 VPWR.n2176 VPWR 0.0233659
R6611 VPWR.n2181 VPWR 0.0233659
R6612 VPWR.n2185 VPWR 0.0233659
R6613 VPWR.n2131 VPWR 0.0233659
R6614 VPWR.n736 VPWR 0.0233659
R6615 VPWR.n731 VPWR 0.0233659
R6616 VPWR.n727 VPWR 0.0233659
R6617 VPWR.n723 VPWR 0.0233659
R6618 VPWR.n715 VPWR 0.0233659
R6619 VPWR.n711 VPWR 0.0233659
R6620 VPWR.n707 VPWR 0.0233659
R6621 VPWR.n703 VPWR 0.0233659
R6622 VPWR.n699 VPWR 0.0233659
R6623 VPWR.n695 VPWR 0.0233659
R6624 VPWR.n691 VPWR 0.0233659
R6625 VPWR.n687 VPWR 0.0233659
R6626 VPWR.n683 VPWR 0.0233659
R6627 VPWR.n679 VPWR 0.0233659
R6628 VPWR.n676 VPWR 0.0233659
R6629 VPWR.n719 VPWR 0.0233659
R6630 VPWR.n2087 VPWR 0.0233659
R6631 VPWR.n2082 VPWR 0.0233659
R6632 VPWR.n2077 VPWR 0.0233659
R6633 VPWR.n2072 VPWR 0.0233659
R6634 VPWR.n2062 VPWR 0.0233659
R6635 VPWR.n2057 VPWR 0.0233659
R6636 VPWR.n2052 VPWR 0.0233659
R6637 VPWR.n2047 VPWR 0.0233659
R6638 VPWR.n2042 VPWR 0.0233659
R6639 VPWR.n2037 VPWR 0.0233659
R6640 VPWR.n2032 VPWR 0.0233659
R6641 VPWR.n2027 VPWR 0.0233659
R6642 VPWR.n2022 VPWR 0.0233659
R6643 VPWR.n2017 VPWR 0.0233659
R6644 VPWR.n2013 VPWR 0.0233659
R6645 VPWR.n2067 VPWR 0.0233659
R6646 VPWR.n772 VPWR 0.0233659
R6647 VPWR.n776 VPWR 0.0233659
R6648 VPWR.n780 VPWR 0.0233659
R6649 VPWR.n784 VPWR 0.0233659
R6650 VPWR.n792 VPWR 0.0233659
R6651 VPWR.n796 VPWR 0.0233659
R6652 VPWR.n800 VPWR 0.0233659
R6653 VPWR.n804 VPWR 0.0233659
R6654 VPWR.n808 VPWR 0.0233659
R6655 VPWR.n812 VPWR 0.0233659
R6656 VPWR.n816 VPWR 0.0233659
R6657 VPWR.n820 VPWR 0.0233659
R6658 VPWR.n824 VPWR 0.0233659
R6659 VPWR.n828 VPWR 0.0233659
R6660 VPWR.n832 VPWR 0.0233659
R6661 VPWR.n788 VPWR 0.0233659
R6662 VPWR.n1915 VPWR 0.0233659
R6663 VPWR.n1920 VPWR 0.0233659
R6664 VPWR.n1925 VPWR 0.0233659
R6665 VPWR.n1930 VPWR 0.0233659
R6666 VPWR.n1940 VPWR 0.0233659
R6667 VPWR.n1945 VPWR 0.0233659
R6668 VPWR.n1950 VPWR 0.0233659
R6669 VPWR.n1955 VPWR 0.0233659
R6670 VPWR.n1960 VPWR 0.0233659
R6671 VPWR.n1965 VPWR 0.0233659
R6672 VPWR.n1970 VPWR 0.0233659
R6673 VPWR.n1975 VPWR 0.0233659
R6674 VPWR.n1980 VPWR 0.0233659
R6675 VPWR.n1985 VPWR 0.0233659
R6676 VPWR.n1989 VPWR 0.0233659
R6677 VPWR.n1935 VPWR 0.0233659
R6678 VPWR.n928 VPWR 0.0233659
R6679 VPWR.n923 VPWR 0.0233659
R6680 VPWR.n919 VPWR 0.0233659
R6681 VPWR.n915 VPWR 0.0233659
R6682 VPWR.n907 VPWR 0.0233659
R6683 VPWR.n903 VPWR 0.0233659
R6684 VPWR.n899 VPWR 0.0233659
R6685 VPWR.n895 VPWR 0.0233659
R6686 VPWR.n891 VPWR 0.0233659
R6687 VPWR.n887 VPWR 0.0233659
R6688 VPWR.n883 VPWR 0.0233659
R6689 VPWR.n879 VPWR 0.0233659
R6690 VPWR.n875 VPWR 0.0233659
R6691 VPWR.n871 VPWR 0.0233659
R6692 VPWR.n868 VPWR 0.0233659
R6693 VPWR.n911 VPWR 0.0233659
R6694 VPWR.n1871 VPWR 0.0233659
R6695 VPWR.n980 VPWR 0.0233659
R6696 VPWR.n1495 VPWR 0.0233659
R6697 VPWR.n1223 VPWR 0.0233659
R6698 VPWR.n400 VPWR 0.0233659
R6699 VPWR.n2464 VPWR 0.0233659
R6700 VPWR.n339 VPWR 0.0233659
R6701 VPWR.n2522 VPWR 0.0233659
R6702 VPWR.n976 VPWR 0.0233659
R6703 VPWR.n1490 VPWR 0.0233659
R6704 VPWR.n1486 VPWR 0.0233659
R6705 VPWR.n1866 VPWR 0.0233659
R6706 VPWR.n984 VPWR 0.0233659
R6707 VPWR.n1504 VPWR 0.0233659
R6708 VPWR.n1174 VPWR 0.0233659
R6709 VPWR.n408 VPWR 0.0233659
R6710 VPWR.n416 VPWR 0.0233659
R6711 VPWR.n420 VPWR 0.0233659
R6712 VPWR.n424 VPWR 0.0233659
R6713 VPWR.n428 VPWR 0.0233659
R6714 VPWR.n432 VPWR 0.0233659
R6715 VPWR.n436 VPWR 0.0233659
R6716 VPWR.n440 VPWR 0.0233659
R6717 VPWR.n444 VPWR 0.0233659
R6718 VPWR.n448 VPWR 0.0233659
R6719 VPWR.n412 VPWR 0.0233659
R6720 VPWR.n2449 VPWR 0.0233659
R6721 VPWR.n327 VPWR 0.0233659
R6722 VPWR.n2539 VPWR 0.0233659
R6723 VPWR.n988 VPWR 0.0233659
R6724 VPWR.n1509 VPWR 0.0233659
R6725 VPWR.n1165 VPWR 0.0233659
R6726 VPWR.n1861 VPWR 0.0233659
R6727 VPWR.n1851 VPWR 0.0233659
R6728 VPWR.n1846 VPWR 0.0233659
R6729 VPWR.n1841 VPWR 0.0233659
R6730 VPWR.n1836 VPWR 0.0233659
R6731 VPWR.n1831 VPWR 0.0233659
R6732 VPWR.n1826 VPWR 0.0233659
R6733 VPWR.n1821 VPWR 0.0233659
R6734 VPWR.n1817 VPWR 0.0233659
R6735 VPWR.n1856 VPWR 0.0233659
R6736 VPWR.n992 VPWR 0.0233659
R6737 VPWR.n1518 VPWR 0.0233659
R6738 VPWR.n1164 VPWR 0.0233659
R6739 VPWR.n2469 VPWR 0.0233659
R6740 VPWR.n343 VPWR 0.0233659
R6741 VPWR.n2515 VPWR 0.0233659
R6742 VPWR.n1130 VPWR 0.0233659
R6743 VPWR.n1129 VPWR 0.0233659
R6744 VPWR.n996 VPWR 0.0233659
R6745 VPWR.n1523 VPWR 0.0233659
R6746 VPWR.n1155 VPWR 0.0233659
R6747 VPWR.n2439 VPWR 0.0233659
R6748 VPWR.n2429 VPWR 0.0233659
R6749 VPWR.n2424 VPWR 0.0233659
R6750 VPWR.n2419 VPWR 0.0233659
R6751 VPWR.n2414 VPWR 0.0233659
R6752 VPWR.n2409 VPWR 0.0233659
R6753 VPWR.n2405 VPWR 0.0233659
R6754 VPWR.n2434 VPWR 0.0233659
R6755 VPWR.n315 VPWR 0.0233659
R6756 VPWR.n2558 VPWR 0.0233659
R6757 VPWR.n1538 VPWR 0.0233659
R6758 VPWR.n1144 VPWR 0.0233659
R6759 VPWR.n1000 VPWR 0.0233659
R6760 VPWR.n1004 VPWR 0.0233659
R6761 VPWR.n1008 VPWR 0.0233659
R6762 VPWR.n1012 VPWR 0.0233659
R6763 VPWR.n1016 VPWR 0.0233659
R6764 VPWR.n1020 VPWR 0.0233659
R6765 VPWR.n1024 VPWR 0.0233659
R6766 VPWR.n968 VPWR 0.0233659
R6767 VPWR.n1473 VPWR 0.0233659
R6768 VPWR.n1590 VPWR 0.0233659
R6769 VPWR.n311 VPWR 0.0233659
R6770 VPWR.n2563 VPWR 0.0233659
R6771 VPWR.n1154 VPWR 0.0233659
R6772 VPWR.n1763 VPWR 0.0233659
R6773 VPWR.n1073 VPWR 0.0233659
R6774 VPWR.n307 VPWR 0.0233659
R6775 VPWR.n303 VPWR 0.0233659
R6776 VPWR.n295 VPWR 0.0233659
R6777 VPWR.n292 VPWR 0.0233659
R6778 VPWR.n299 VPWR 0.0233659
R6779 VPWR.n1743 VPWR 0.0233659
R6780 VPWR.n1751 VPWR 0.0233659
R6781 VPWR.n1789 VPWR 0.0233659
R6782 VPWR.n1793 VPWR 0.0233659
R6783 VPWR.n1758 VPWR 0.0233659
R6784 VPWR.n1054 VPWR 0.0233659
R6785 VPWR.n2575 VPWR 0.0233659
R6786 VPWR.n2582 VPWR 0.0233659
R6787 VPWR.n2593 VPWR 0.0233659
R6788 VPWR.n2587 VPWR 0.0233659
R6789 VPWR.n1736 VPWR 0.0233659
R6790 VPWR.n1060 VPWR 0.0233659
R6791 VPWR.n1121 VPWR 0.0233659
R6792 VPWR.n1336 VPWR 0.0226354
R6793 VPWR.n1327 VPWR 0.0226354
R6794 VPWR.n1413 VPWR 0.0226354
R6795 VPWR.n2772 VPWR 0.0226354
R6796 VPWR VPWR.n2732 0.0226354
R6797 VPWR VPWR.n2702 0.0226354
R6798 VPWR VPWR.n2664 0.0226354
R6799 VPWR VPWR.n64 0.0220517
R6800 VPWR VPWR.n67 0.0220517
R6801 VPWR VPWR.n70 0.0220517
R6802 VPWR VPWR.n73 0.0220517
R6803 VPWR VPWR.n76 0.0220517
R6804 VPWR VPWR.n79 0.0220517
R6805 VPWR VPWR.n82 0.0220517
R6806 VPWR VPWR.n85 0.0220517
R6807 VPWR VPWR.n88 0.0220517
R6808 VPWR VPWR.n91 0.0220517
R6809 VPWR VPWR.n94 0.0220517
R6810 VPWR VPWR.n97 0.0220517
R6811 VPWR.n289 VPWR 0.0220517
R6812 VPWR VPWR.n61 0.0220517
R6813 VPWR VPWR.n58 0.0220517
R6814 VPWR.n1735 VPWR 0.0220517
R6815 VPWR VPWR.n1057 0.0220517
R6816 VPWR.n1705 VPWR 0.0220517
R6817 VPWR.n1694 VPWR 0.0220517
R6818 VPWR.n1196 VPWR 0.0220517
R6819 VPWR.n1678 VPWR 0.0220517
R6820 VPWR.n1667 VPWR 0.0220517
R6821 VPWR.n1210 VPWR 0.0220517
R6822 VPWR.n1651 VPWR 0.0220517
R6823 VPWR.n1640 VPWR 0.0220517
R6824 VPWR.n1178 VPWR 0.0220517
R6825 VPWR.n1624 VPWR 0.0220517
R6826 VPWR.n1613 VPWR 0.0220517
R6827 VPWR.n1127 VPWR 0.0220517
R6828 VPWR.n1597 VPWR 0.0220517
R6829 VPWR.n1273 VPWR 0.0213333
R6830 VPWR.n1297 VPWR 0.0213333
R6831 VPWR.n1311 VPWR 0.0213333
R6832 VPWR.n1375 VPWR 0.0213333
R6833 VPWR.n1347 VPWR 0.0213333
R6834 VPWR.n1386 VPWR 0.0213333
R6835 VPWR.n1423 VPWR 0.0213333
R6836 VPWR.n2806 VPWR 0.0213333
R6837 VPWR.n2799 VPWR 0.0213333
R6838 VPWR VPWR.n2790 0.0213333
R6839 VPWR.n2792 VPWR 0.0213333
R6840 VPWR VPWR.n2770 0.0213333
R6841 VPWR VPWR.n2751 0.0213333
R6842 VPWR VPWR.n2738 0.0213333
R6843 VPWR.n2500 VPWR 0.0196917
R6844 VPWR.n24 VPWR 0.0143889
R6845 VPWR VPWR.n19 0.0099
R6846 VPWR VPWR.n1604 0.00397222
R6847 VPWR VPWR.n1105 0.00397222
R6848 VPWR VPWR.n1103 0.00397222
R6849 VPWR VPWR.n1631 0.00397222
R6850 VPWR VPWR.n1095 0.00397222
R6851 VPWR VPWR.n1093 0.00397222
R6852 VPWR VPWR.n1658 0.00397222
R6853 VPWR VPWR.n1085 0.00397222
R6854 VPWR VPWR.n1083 0.00397222
R6855 VPWR VPWR.n1685 0.00397222
R6856 VPWR VPWR.n1075 0.00397222
R6857 VPWR VPWR.n1072 0.00397222
R6858 VPWR VPWR.n1712 0.00397222
R6859 VPWR VPWR.n1724 0.00397222
R6860 VPWR.n1113 VPWR 0.00397222
R6861 VPWR VPWR.n1066 0.00397222
R6862 VPWR VPWR.n122 0.00397222
R6863 VPWR VPWR.n111 0.00397222
R6864 VPWR VPWR.n102 0.00397222
R6865 VPWR VPWR.n277 0.00397222
R6866 VPWR VPWR.n265 0.00397222
R6867 VPWR VPWR.n253 0.00397222
R6868 VPWR VPWR.n241 0.00397222
R6869 VPWR VPWR.n229 0.00397222
R6870 VPWR VPWR.n217 0.00397222
R6871 VPWR VPWR.n205 0.00397222
R6872 VPWR VPWR.n193 0.00397222
R6873 VPWR VPWR.n181 0.00397222
R6874 VPWR VPWR.n169 0.00397222
R6875 VPWR VPWR.n157 0.00397222
R6876 VPWR VPWR.n145 0.00397222
R6877 VPWR VPWR.n133 0.00397222
R6878 VPWR.n1462 VPWR.n1461 0.00351282
R6879 VPWR.n1457 VPWR.n1136 0.00351282
R6880 VPWR.n1582 VPWR.n1581 0.00351282
R6881 VPWR.n1577 VPWR.n1576 0.00351282
R6882 VPWR.n1572 VPWR.n1571 0.00351282
R6883 VPWR.n1567 VPWR.n1566 0.00351282
R6884 VPWR.n1562 VPWR.n1561 0.00351282
R6885 VPWR.n1557 VPWR.n1556 0.00351282
R6886 VPWR.n1552 VPWR.n1551 0.00351282
R6887 VPWR.n1547 VPWR.n1546 0.00351282
R6888 VPWR.n1542 VPWR.n1042 0.00351282
R6889 VPWR.n1785 VPWR.n1784 0.00351282
R6890 VPWR.n1776 VPWR.n1772 0.00351282
R6891 VPWR.n1771 VPWR.n1767 0.00351282
R6892 VPWR.n141 VPWR.n140 0.00265517
R6893 VPWR.n153 VPWR.n152 0.00265517
R6894 VPWR.n165 VPWR.n164 0.00265517
R6895 VPWR.n177 VPWR.n176 0.00265517
R6896 VPWR.n189 VPWR.n188 0.00265517
R6897 VPWR.n201 VPWR.n200 0.00265517
R6898 VPWR.n213 VPWR.n212 0.00265517
R6899 VPWR.n225 VPWR.n224 0.00265517
R6900 VPWR.n237 VPWR.n236 0.00265517
R6901 VPWR.n249 VPWR.n248 0.00265517
R6902 VPWR.n261 VPWR.n260 0.00265517
R6903 VPWR.n273 VPWR.n272 0.00265517
R6904 VPWR.n288 VPWR.n286 0.00265517
R6905 VPWR.n129 VPWR.n128 0.00265517
R6906 VPWR.n118 VPWR.n117 0.00265517
R6907 VPWR.n1734 VPWR.n1732 0.00265517
R6908 VPWR.n1720 VPWR.n1719 0.00265517
R6909 VPWR.n1708 VPWR.n1707 0.00265517
R6910 VPWR.n1697 VPWR.n1696 0.00265517
R6911 VPWR.n1195 VPWR.n1193 0.00265517
R6912 VPWR.n1681 VPWR.n1680 0.00265517
R6913 VPWR.n1670 VPWR.n1669 0.00265517
R6914 VPWR.n1209 VPWR.n1207 0.00265517
R6915 VPWR.n1654 VPWR.n1653 0.00265517
R6916 VPWR.n1643 VPWR.n1642 0.00265517
R6917 VPWR.n1177 VPWR.n1175 0.00265517
R6918 VPWR.n1627 VPWR.n1626 0.00265517
R6919 VPWR.n1616 VPWR.n1615 0.00265517
R6920 VPWR.n1126 VPWR.n1124 0.00265517
R6921 VPWR.n1600 VPWR.n1599 0.00265517
R6922 XThC.Tn[10].n71 XThC.Tn[10].n70 256.104
R6923 XThC.Tn[10].n75 XThC.Tn[10].n74 243.679
R6924 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R6925 XThC.Tn[10].n75 XThC.Tn[10].n73 205.28
R6926 XThC.Tn[10].n71 XThC.Tn[10].n69 202.095
R6927 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R6928 XThC.Tn[10].n65 XThC.Tn[10].n63 161.365
R6929 XThC.Tn[10].n61 XThC.Tn[10].n59 161.365
R6930 XThC.Tn[10].n57 XThC.Tn[10].n55 161.365
R6931 XThC.Tn[10].n53 XThC.Tn[10].n51 161.365
R6932 XThC.Tn[10].n49 XThC.Tn[10].n47 161.365
R6933 XThC.Tn[10].n45 XThC.Tn[10].n43 161.365
R6934 XThC.Tn[10].n41 XThC.Tn[10].n39 161.365
R6935 XThC.Tn[10].n37 XThC.Tn[10].n35 161.365
R6936 XThC.Tn[10].n33 XThC.Tn[10].n31 161.365
R6937 XThC.Tn[10].n29 XThC.Tn[10].n27 161.365
R6938 XThC.Tn[10].n25 XThC.Tn[10].n23 161.365
R6939 XThC.Tn[10].n21 XThC.Tn[10].n19 161.365
R6940 XThC.Tn[10].n17 XThC.Tn[10].n15 161.365
R6941 XThC.Tn[10].n13 XThC.Tn[10].n11 161.365
R6942 XThC.Tn[10].n9 XThC.Tn[10].n7 161.365
R6943 XThC.Tn[10].n6 XThC.Tn[10].n4 161.365
R6944 XThC.Tn[10].n63 XThC.Tn[10].t42 161.202
R6945 XThC.Tn[10].n59 XThC.Tn[10].t32 161.202
R6946 XThC.Tn[10].n55 XThC.Tn[10].t19 161.202
R6947 XThC.Tn[10].n51 XThC.Tn[10].t16 161.202
R6948 XThC.Tn[10].n47 XThC.Tn[10].t40 161.202
R6949 XThC.Tn[10].n43 XThC.Tn[10].t27 161.202
R6950 XThC.Tn[10].n39 XThC.Tn[10].t26 161.202
R6951 XThC.Tn[10].n35 XThC.Tn[10].t39 161.202
R6952 XThC.Tn[10].n31 XThC.Tn[10].t37 161.202
R6953 XThC.Tn[10].n27 XThC.Tn[10].t28 161.202
R6954 XThC.Tn[10].n23 XThC.Tn[10].t15 161.202
R6955 XThC.Tn[10].n19 XThC.Tn[10].t14 161.202
R6956 XThC.Tn[10].n15 XThC.Tn[10].t25 161.202
R6957 XThC.Tn[10].n11 XThC.Tn[10].t23 161.202
R6958 XThC.Tn[10].n7 XThC.Tn[10].t21 161.202
R6959 XThC.Tn[10].n4 XThC.Tn[10].t36 161.202
R6960 XThC.Tn[10].n63 XThC.Tn[10].t13 145.137
R6961 XThC.Tn[10].n59 XThC.Tn[10].t35 145.137
R6962 XThC.Tn[10].n55 XThC.Tn[10].t22 145.137
R6963 XThC.Tn[10].n51 XThC.Tn[10].t20 145.137
R6964 XThC.Tn[10].n47 XThC.Tn[10].t12 145.137
R6965 XThC.Tn[10].n43 XThC.Tn[10].t33 145.137
R6966 XThC.Tn[10].n39 XThC.Tn[10].t31 145.137
R6967 XThC.Tn[10].n35 XThC.Tn[10].t43 145.137
R6968 XThC.Tn[10].n31 XThC.Tn[10].t41 145.137
R6969 XThC.Tn[10].n27 XThC.Tn[10].t34 145.137
R6970 XThC.Tn[10].n23 XThC.Tn[10].t18 145.137
R6971 XThC.Tn[10].n19 XThC.Tn[10].t17 145.137
R6972 XThC.Tn[10].n15 XThC.Tn[10].t30 145.137
R6973 XThC.Tn[10].n11 XThC.Tn[10].t29 145.137
R6974 XThC.Tn[10].n7 XThC.Tn[10].t24 145.137
R6975 XThC.Tn[10].n4 XThC.Tn[10].t38 145.137
R6976 XThC.Tn[10].n69 XThC.Tn[10].t5 26.5955
R6977 XThC.Tn[10].n69 XThC.Tn[10].t4 26.5955
R6978 XThC.Tn[10].n70 XThC.Tn[10].t9 26.5955
R6979 XThC.Tn[10].n70 XThC.Tn[10].t1 26.5955
R6980 XThC.Tn[10].n73 XThC.Tn[10].t7 26.5955
R6981 XThC.Tn[10].n73 XThC.Tn[10].t6 26.5955
R6982 XThC.Tn[10].n74 XThC.Tn[10].t11 26.5955
R6983 XThC.Tn[10].n74 XThC.Tn[10].t0 26.5955
R6984 XThC.Tn[10].n1 XThC.Tn[10].t10 24.9236
R6985 XThC.Tn[10].n1 XThC.Tn[10].t3 24.9236
R6986 XThC.Tn[10].n0 XThC.Tn[10].t2 24.9236
R6987 XThC.Tn[10].n0 XThC.Tn[10].t8 24.9236
R6988 XThC.Tn[10] XThC.Tn[10].n75 22.9652
R6989 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R6990 XThC.Tn[10].n72 XThC.Tn[10].n71 13.9299
R6991 XThC.Tn[10] XThC.Tn[10].n72 13.9299
R6992 XThC.Tn[10] XThC.Tn[10].n6 8.0245
R6993 XThC.Tn[10].n66 XThC.Tn[10].n65 7.9105
R6994 XThC.Tn[10].n62 XThC.Tn[10].n61 7.9105
R6995 XThC.Tn[10].n58 XThC.Tn[10].n57 7.9105
R6996 XThC.Tn[10].n54 XThC.Tn[10].n53 7.9105
R6997 XThC.Tn[10].n50 XThC.Tn[10].n49 7.9105
R6998 XThC.Tn[10].n46 XThC.Tn[10].n45 7.9105
R6999 XThC.Tn[10].n42 XThC.Tn[10].n41 7.9105
R7000 XThC.Tn[10].n38 XThC.Tn[10].n37 7.9105
R7001 XThC.Tn[10].n34 XThC.Tn[10].n33 7.9105
R7002 XThC.Tn[10].n30 XThC.Tn[10].n29 7.9105
R7003 XThC.Tn[10].n26 XThC.Tn[10].n25 7.9105
R7004 XThC.Tn[10].n22 XThC.Tn[10].n21 7.9105
R7005 XThC.Tn[10].n18 XThC.Tn[10].n17 7.9105
R7006 XThC.Tn[10].n14 XThC.Tn[10].n13 7.9105
R7007 XThC.Tn[10].n10 XThC.Tn[10].n9 7.9105
R7008 XThC.Tn[10].n68 XThC.Tn[10].n67 7.40985
R7009 XThC.Tn[10].n67 XThC.Tn[10] 4.38575
R7010 XThC.Tn[10].n72 XThC.Tn[10].n68 2.99115
R7011 XThC.Tn[10].n72 XThC.Tn[10] 2.87153
R7012 XThC.Tn[10].n3 XThC.Tn[10] 2.688
R7013 XThC.Tn[10].n68 XThC.Tn[10] 2.2734
R7014 XThC.Tn[10].n67 XThC.Tn[10].n3 0.244922
R7015 XThC.Tn[10].n10 XThC.Tn[10] 0.235138
R7016 XThC.Tn[10].n14 XThC.Tn[10] 0.235138
R7017 XThC.Tn[10].n18 XThC.Tn[10] 0.235138
R7018 XThC.Tn[10].n22 XThC.Tn[10] 0.235138
R7019 XThC.Tn[10].n26 XThC.Tn[10] 0.235138
R7020 XThC.Tn[10].n30 XThC.Tn[10] 0.235138
R7021 XThC.Tn[10].n34 XThC.Tn[10] 0.235138
R7022 XThC.Tn[10].n38 XThC.Tn[10] 0.235138
R7023 XThC.Tn[10].n42 XThC.Tn[10] 0.235138
R7024 XThC.Tn[10].n46 XThC.Tn[10] 0.235138
R7025 XThC.Tn[10].n50 XThC.Tn[10] 0.235138
R7026 XThC.Tn[10].n54 XThC.Tn[10] 0.235138
R7027 XThC.Tn[10].n58 XThC.Tn[10] 0.235138
R7028 XThC.Tn[10].n62 XThC.Tn[10] 0.235138
R7029 XThC.Tn[10].n66 XThC.Tn[10] 0.235138
R7030 XThC.Tn[10].n3 XThC.Tn[10] 0.141947
R7031 XThC.Tn[10] XThC.Tn[10].n10 0.114505
R7032 XThC.Tn[10] XThC.Tn[10].n14 0.114505
R7033 XThC.Tn[10] XThC.Tn[10].n18 0.114505
R7034 XThC.Tn[10] XThC.Tn[10].n22 0.114505
R7035 XThC.Tn[10] XThC.Tn[10].n26 0.114505
R7036 XThC.Tn[10] XThC.Tn[10].n30 0.114505
R7037 XThC.Tn[10] XThC.Tn[10].n34 0.114505
R7038 XThC.Tn[10] XThC.Tn[10].n38 0.114505
R7039 XThC.Tn[10] XThC.Tn[10].n42 0.114505
R7040 XThC.Tn[10] XThC.Tn[10].n46 0.114505
R7041 XThC.Tn[10] XThC.Tn[10].n50 0.114505
R7042 XThC.Tn[10] XThC.Tn[10].n54 0.114505
R7043 XThC.Tn[10] XThC.Tn[10].n58 0.114505
R7044 XThC.Tn[10] XThC.Tn[10].n62 0.114505
R7045 XThC.Tn[10] XThC.Tn[10].n66 0.114505
R7046 XThC.Tn[10].n65 XThC.Tn[10].n64 0.0599512
R7047 XThC.Tn[10].n61 XThC.Tn[10].n60 0.0599512
R7048 XThC.Tn[10].n57 XThC.Tn[10].n56 0.0599512
R7049 XThC.Tn[10].n53 XThC.Tn[10].n52 0.0599512
R7050 XThC.Tn[10].n49 XThC.Tn[10].n48 0.0599512
R7051 XThC.Tn[10].n45 XThC.Tn[10].n44 0.0599512
R7052 XThC.Tn[10].n41 XThC.Tn[10].n40 0.0599512
R7053 XThC.Tn[10].n37 XThC.Tn[10].n36 0.0599512
R7054 XThC.Tn[10].n33 XThC.Tn[10].n32 0.0599512
R7055 XThC.Tn[10].n29 XThC.Tn[10].n28 0.0599512
R7056 XThC.Tn[10].n25 XThC.Tn[10].n24 0.0599512
R7057 XThC.Tn[10].n21 XThC.Tn[10].n20 0.0599512
R7058 XThC.Tn[10].n17 XThC.Tn[10].n16 0.0599512
R7059 XThC.Tn[10].n13 XThC.Tn[10].n12 0.0599512
R7060 XThC.Tn[10].n9 XThC.Tn[10].n8 0.0599512
R7061 XThC.Tn[10].n6 XThC.Tn[10].n5 0.0599512
R7062 XThC.Tn[10].n64 XThC.Tn[10] 0.0469286
R7063 XThC.Tn[10].n60 XThC.Tn[10] 0.0469286
R7064 XThC.Tn[10].n56 XThC.Tn[10] 0.0469286
R7065 XThC.Tn[10].n52 XThC.Tn[10] 0.0469286
R7066 XThC.Tn[10].n48 XThC.Tn[10] 0.0469286
R7067 XThC.Tn[10].n44 XThC.Tn[10] 0.0469286
R7068 XThC.Tn[10].n40 XThC.Tn[10] 0.0469286
R7069 XThC.Tn[10].n36 XThC.Tn[10] 0.0469286
R7070 XThC.Tn[10].n32 XThC.Tn[10] 0.0469286
R7071 XThC.Tn[10].n28 XThC.Tn[10] 0.0469286
R7072 XThC.Tn[10].n24 XThC.Tn[10] 0.0469286
R7073 XThC.Tn[10].n20 XThC.Tn[10] 0.0469286
R7074 XThC.Tn[10].n16 XThC.Tn[10] 0.0469286
R7075 XThC.Tn[10].n12 XThC.Tn[10] 0.0469286
R7076 XThC.Tn[10].n8 XThC.Tn[10] 0.0469286
R7077 XThC.Tn[10].n5 XThC.Tn[10] 0.0469286
R7078 XThC.Tn[10].n64 XThC.Tn[10] 0.0401341
R7079 XThC.Tn[10].n60 XThC.Tn[10] 0.0401341
R7080 XThC.Tn[10].n56 XThC.Tn[10] 0.0401341
R7081 XThC.Tn[10].n52 XThC.Tn[10] 0.0401341
R7082 XThC.Tn[10].n48 XThC.Tn[10] 0.0401341
R7083 XThC.Tn[10].n44 XThC.Tn[10] 0.0401341
R7084 XThC.Tn[10].n40 XThC.Tn[10] 0.0401341
R7085 XThC.Tn[10].n36 XThC.Tn[10] 0.0401341
R7086 XThC.Tn[10].n32 XThC.Tn[10] 0.0401341
R7087 XThC.Tn[10].n28 XThC.Tn[10] 0.0401341
R7088 XThC.Tn[10].n24 XThC.Tn[10] 0.0401341
R7089 XThC.Tn[10].n20 XThC.Tn[10] 0.0401341
R7090 XThC.Tn[10].n16 XThC.Tn[10] 0.0401341
R7091 XThC.Tn[10].n12 XThC.Tn[10] 0.0401341
R7092 XThC.Tn[10].n8 XThC.Tn[10] 0.0401341
R7093 XThC.Tn[10].n5 XThC.Tn[10] 0.0401341
R7094 VGND.n3019 VGND.n3018 15660.6
R7095 VGND.n196 VGND.n195 13477
R7096 VGND.n3018 VGND.n7 11578
R7097 VGND.n195 VGND.n7 10429.6
R7098 VGND.n3012 VGND.n8 9309.26
R7099 VGND.n200 VGND.n199 9223.7
R7100 VGND.n198 VGND.n197 9223.7
R7101 VGND.n197 VGND.n196 9223.7
R7102 VGND.n2969 VGND.n200 9223.7
R7103 VGND.n2969 VGND.n2968 7447.41
R7104 VGND.n2249 VGND.n2248 7387.65
R7105 VGND.n2250 VGND.n2249 7387.65
R7106 VGND.n2285 VGND.n2284 7387.65
R7107 VGND.n3017 VGND.n3016 7387.65
R7108 VGND.n3016 VGND.n3015 7387.65
R7109 VGND.n3015 VGND.n3014 7387.65
R7110 VGND.n3014 VGND.n3013 7387.65
R7111 VGND.n3013 VGND.n3012 7387.65
R7112 VGND.n2351 VGND.n2285 6674.35
R7113 VGND.n1386 VGND.t1112 6324.96
R7114 VGND.n199 VGND.n198 5231.11
R7115 VGND.n1336 VGND.t1681 5168.13
R7116 VGND.n2967 VGND.n8 5074.71
R7117 VGND.n3018 VGND.n3017 5063.19
R7118 VGND.n1154 VGND.n806 4539.15
R7119 VGND VGND.n8 4240.58
R7120 VGND.t1879 VGND.t1411 4212.19
R7121 VGND.t1885 VGND.t2050 4212.19
R7122 VGND.t1900 VGND.t1311 4212.19
R7123 VGND.t1978 VGND.t1269 4212.19
R7124 VGND.t1984 VGND.t571 4212.19
R7125 VGND.t1903 VGND.t2364 4212.19
R7126 VGND.t1948 VGND.t1086 4212.19
R7127 VGND.t2367 VGND.t1993 4212.19
R7128 VGND.t111 VGND.t1912 4212.19
R7129 VGND.t2526 VGND.t1957 4212.19
R7130 VGND.t2341 VGND.t1996 4212.19
R7131 VGND.t1529 VGND.t2008 4212.19
R7132 VGND.t2503 VGND.t1924 4212.19
R7133 VGND.t2405 VGND.t1966 4212.19
R7134 VGND.n2919 VGND.n222 4077.12
R7135 VGND.n1340 VGND.n1338 3417.39
R7136 VGND.n1340 VGND.n1339 3417.39
R7137 VGND.n1388 VGND.n1387 3417.39
R7138 VGND.n2180 VGND.n504 3417.39
R7139 VGND.n503 VGND.n473 3417.39
R7140 VGND.n2353 VGND.n2352 3417.39
R7141 VGND.n2920 VGND.n2919 3331.79
R7142 VGND.n2921 VGND.n2920 3331.79
R7143 VGND.n2922 VGND.n2921 3331.79
R7144 VGND.n2923 VGND.n2922 3331.79
R7145 VGND.n2924 VGND.n2923 3331.79
R7146 VGND.n2925 VGND.n2924 3331.79
R7147 VGND.n2926 VGND.n2925 3331.79
R7148 VGND.n2927 VGND.n2926 3331.79
R7149 VGND.n2928 VGND.n2927 3331.79
R7150 VGND.n2929 VGND.n2928 3331.79
R7151 VGND.n2930 VGND.n2929 3331.79
R7152 VGND.n2931 VGND.n2930 3331.79
R7153 VGND.n2932 VGND.n2931 3331.79
R7154 VGND.n2933 VGND.n2932 3331.79
R7155 VGND.n2934 VGND.n2933 3331.79
R7156 VGND.n1339 VGND.n806 3273.91
R7157 VGND.n2181 VGND.n539 3265.22
R7158 VGND.n2934 VGND.n201 2725.63
R7159 VGND.n197 VGND.t910 2655.17
R7160 VGND.n196 VGND.t886 2655.17
R7161 VGND.n2353 VGND.n2285 2517.39
R7162 VGND.t192 VGND.n201 2334.15
R7163 VGND.t1648 VGND.n2701 2307.69
R7164 VGND.n359 VGND.t1722 2307.69
R7165 VGND.n360 VGND.t1735 2307.69
R7166 VGND.n370 VGND.t1589 2307.69
R7167 VGND.n371 VGND.t1656 2307.69
R7168 VGND.n381 VGND.t1748 2307.69
R7169 VGND.n382 VGND.t1817 2307.69
R7170 VGND.t1601 VGND.n327 2307.69
R7171 VGND.n2705 VGND.t1686 2307.69
R7172 VGND.n2728 VGND.t1747 2307.69
R7173 VGND.n2738 VGND.t1603 2307.69
R7174 VGND.t1613 VGND.n2737 2307.69
R7175 VGND.n2731 VGND.t1695 2307.69
R7176 VGND.n2776 VGND.t1778 2307.69
R7177 VGND.t1801 VGND.n2775 2307.69
R7178 VGND.n2943 VGND.t1698 2307.69
R7179 VGND.t1930 VGND.n2703 2280.49
R7180 VGND.n3020 VGND.n5 2229.43
R7181 VGND.n3020 VGND.n6 2229.43
R7182 VGND.n2348 VGND.n6 2229.43
R7183 VGND.n2348 VGND.n5 2229.43
R7184 VGND.n1338 VGND.n1337 2173.91
R7185 VGND.n2704 VGND.t2549 2132.93
R7186 VGND.n2701 VGND.t1813 2123.08
R7187 VGND.t1653 VGND.n359 2123.08
R7188 VGND.n360 VGND.t1675 2123.08
R7189 VGND.t1815 VGND.n370 2123.08
R7190 VGND.n371 VGND.t1826 2123.08
R7191 VGND.t1606 VGND.n381 2123.08
R7192 VGND.n382 VGND.t1745 2123.08
R7193 VGND.n2705 VGND.t1610 2123.08
R7194 VGND.t1691 VGND.n2728 2123.08
R7195 VGND.n2738 VGND.t1703 2123.08
R7196 VGND.n2737 VGND.t1797 2123.08
R7197 VGND.n2731 VGND.t1623 2123.08
R7198 VGND.n2776 VGND.t1715 2123.08
R7199 VGND.n2775 VGND.t1783 2123.08
R7200 VGND.n2704 VGND.t1954 2079.27
R7201 VGND.t1411 VGND.t1930 2012.2
R7202 VGND.t2050 VGND.t1879 2012.2
R7203 VGND.t1311 VGND.t1885 2012.2
R7204 VGND.t1269 VGND.t1900 2012.2
R7205 VGND.t571 VGND.t1978 2012.2
R7206 VGND.t2364 VGND.t1984 2012.2
R7207 VGND.t1086 VGND.t1903 2012.2
R7208 VGND.t2549 VGND.t1948 2012.2
R7209 VGND.t1954 VGND.t2367 2012.2
R7210 VGND.t1993 VGND.t111 2012.2
R7211 VGND.t1912 VGND.t2526 2012.2
R7212 VGND.t1957 VGND.t2341 2012.2
R7213 VGND.t1996 VGND.t1529 2012.2
R7214 VGND.t2008 VGND.t2503 2012.2
R7215 VGND.t1924 VGND.t2405 2012.2
R7216 VGND.t1966 VGND.t192 2012.2
R7217 VGND.n199 VGND 1997.7
R7218 VGND.n200 VGND 1997.7
R7219 VGND VGND.n2969 1997.7
R7220 VGND.n2968 VGND.n2944 1907.51
R7221 VGND.n2284 VGND.n2251 1831.57
R7222 VGND.n198 VGND.t845 1807.04
R7223 VGND.n2970 VGND.t1110 1785.51
R7224 VGND.n2352 VGND.n2351 1760.87
R7225 VGND.n2702 VGND.t1733 1738.46
R7226 VGND.n2250 VGND.n504 1691.3
R7227 VGND.n2351 VGND.n2350 1656.52
R7228 VGND.t947 VGND.n66 1618.39
R7229 VGND.n3011 VGND.t2016 1618.39
R7230 VGND.n2971 VGND.t2464 1618.39
R7231 VGND.n2702 VGND.n7 1604.17
R7232 VGND.n2350 VGND.n328 1517.39
R7233 VGND.n195 VGND.t861 1517.24
R7234 VGND.n2248 VGND.n540 1513.49
R7235 VGND.t1768 VGND.n2704 1507.69
R7236 VGND.n2703 VGND.n2702 1441.28
R7237 VGND.n1386 VGND.n540 1370.36
R7238 VGND.t1733 VGND.t1811 1353.85
R7239 VGND.t1811 VGND.t1648 1353.85
R7240 VGND.t1651 VGND.t1813 1353.85
R7241 VGND.t1722 VGND.t1651 1353.85
R7242 VGND.t1729 VGND.t1653 1353.85
R7243 VGND.t1735 VGND.t1729 1353.85
R7244 VGND.t1675 VGND.t1749 1353.85
R7245 VGND.t1749 VGND.t1589 1353.85
R7246 VGND.t1818 VGND.t1815 1353.85
R7247 VGND.t1656 VGND.t1818 1353.85
R7248 VGND.t1826 VGND.t1673 1353.85
R7249 VGND.t1673 VGND.t1748 1353.85
R7250 VGND.t1687 VGND.t1606 1353.85
R7251 VGND.t1817 VGND.t1687 1353.85
R7252 VGND.t1745 VGND.t1822 1353.85
R7253 VGND.t1822 VGND.t1601 1353.85
R7254 VGND.t1604 VGND.t1768 1353.85
R7255 VGND.t1686 VGND.t1604 1353.85
R7256 VGND.t1610 VGND.t1671 1353.85
R7257 VGND.t1671 VGND.t1747 1353.85
R7258 VGND.t1766 VGND.t1691 1353.85
R7259 VGND.t1603 VGND.t1766 1353.85
R7260 VGND.t1703 VGND.t1781 1353.85
R7261 VGND.t1781 VGND.t1613 1353.85
R7262 VGND.t1689 VGND.t1797 1353.85
R7263 VGND.t1695 VGND.t1689 1353.85
R7264 VGND.t1623 VGND.t1701 1353.85
R7265 VGND.t1701 VGND.t1778 1353.85
R7266 VGND.t1715 VGND.t1717 1353.85
R7267 VGND.t1717 VGND.t1801 1353.85
R7268 VGND.t1783 VGND.t1619 1353.85
R7269 VGND.t1619 VGND.t1698 1353.85
R7270 VGND.n2944 VGND.n201 1301.35
R7271 VGND.n2703 VGND.n328 1278.26
R7272 VGND.t1876 VGND.n540 1270.28
R7273 VGND.n1127 VGND.t984 1268.93
R7274 VGND.n1127 VGND.t36 1268.93
R7275 VGND.n502 VGND.t130 1253.59
R7276 VGND.t122 VGND.n502 1253.59
R7277 VGND.n2283 VGND.t14 1253.59
R7278 VGND.t126 VGND.n2283 1253.59
R7279 VGND.n538 VGND.t39 1253.59
R7280 VGND.t132 VGND.n538 1253.59
R7281 VGND.n2247 VGND.t41 1253.59
R7282 VGND.t9 VGND.n2247 1253.59
R7283 VGND.n1385 VGND.t16 1253.59
R7284 VGND.t20 VGND.n1385 1253.59
R7285 VGND.n1337 VGND.n1336 1243.48
R7286 VGND.n2251 VGND.t1921 1237.71
R7287 VGND.n66 VGND.t1003 1213.79
R7288 VGND.n2967 VGND.n2966 1198.25
R7289 VGND.n1155 VGND.n1154 1198.25
R7290 VGND.n2943 VGND.n2942 1180.79
R7291 VGND.n2936 VGND.n2935 1180.79
R7292 VGND.n2534 VGND.n208 1180.79
R7293 VGND.n2529 VGND.n209 1180.79
R7294 VGND.n2817 VGND.n210 1180.79
R7295 VGND.n1989 VGND.n211 1180.79
R7296 VGND.n1996 VGND.n212 1180.79
R7297 VGND.n2842 VGND.n213 1180.79
R7298 VGND.n1829 VGND.n214 1180.79
R7299 VGND.n1836 VGND.n215 1180.79
R7300 VGND.n2867 VGND.n216 1180.79
R7301 VGND.n1655 VGND.n217 1180.79
R7302 VGND.n1650 VGND.n218 1180.79
R7303 VGND.n2892 VGND.n219 1180.79
R7304 VGND.n1607 VGND.n220 1180.79
R7305 VGND.n2912 VGND.n221 1180.79
R7306 VGND.n1282 VGND.n222 1180.79
R7307 VGND.n2918 VGND.n2917 1180.79
R7308 VGND.n1335 VGND.n1334 1180.46
R7309 VGND.n929 VGND.n890 1180.46
R7310 VGND.n934 VGND.n933 1180.46
R7311 VGND.n939 VGND.n938 1180.46
R7312 VGND.n944 VGND.n943 1180.46
R7313 VGND.n949 VGND.n948 1180.46
R7314 VGND.n954 VGND.n953 1180.46
R7315 VGND.n959 VGND.n958 1180.46
R7316 VGND.n964 VGND.n963 1180.46
R7317 VGND.n969 VGND.n968 1180.46
R7318 VGND.n974 VGND.n973 1180.46
R7319 VGND.n979 VGND.n978 1180.46
R7320 VGND.n984 VGND.n983 1180.46
R7321 VGND.n989 VGND.n988 1180.46
R7322 VGND.n991 VGND.n990 1180.46
R7323 VGND.n1279 VGND.n1278 1180.46
R7324 VGND.n1277 VGND.n1276 1180.46
R7325 VGND.n1234 VGND.n1233 1180.46
R7326 VGND.n1239 VGND.n1238 1180.46
R7327 VGND.n1241 VGND.n1240 1180.46
R7328 VGND.n1246 VGND.n1245 1180.46
R7329 VGND.n1248 VGND.n1247 1180.46
R7330 VGND.n1220 VGND.n1219 1180.46
R7331 VGND.n1209 VGND.n1208 1180.46
R7332 VGND.n1207 VGND.n1206 1180.46
R7333 VGND.n1190 VGND.n1189 1180.46
R7334 VGND.n1188 VGND.n1187 1180.46
R7335 VGND.n1177 VGND.n1176 1180.46
R7336 VGND.n1175 VGND.n1174 1180.46
R7337 VGND.n1167 VGND.n1166 1180.46
R7338 VGND.n2775 VGND.n2774 1180.46
R7339 VGND.n2777 VGND.n2776 1180.46
R7340 VGND.n2732 VGND.n2731 1180.46
R7341 VGND.n2737 VGND.n2736 1180.46
R7342 VGND.n2739 VGND.n2738 1180.46
R7343 VGND.n2728 VGND.n2727 1180.46
R7344 VGND.n2706 VGND.n2705 1180.46
R7345 VGND.n388 VGND.n327 1180.46
R7346 VGND.n383 VGND.n382 1180.46
R7347 VGND.n381 VGND.n380 1180.46
R7348 VGND.n372 VGND.n371 1180.46
R7349 VGND.n370 VGND.n369 1180.46
R7350 VGND.n361 VGND.n360 1180.46
R7351 VGND.n359 VGND.n333 1180.46
R7352 VGND.n2701 VGND.n2700 1180.46
R7353 VGND.n2641 VGND.n2640 1180.46
R7354 VGND.n2646 VGND.n2645 1180.46
R7355 VGND.n2651 VGND.n2650 1180.46
R7356 VGND.n2656 VGND.n2655 1180.46
R7357 VGND.n2661 VGND.n2660 1180.46
R7358 VGND.n2666 VGND.n2665 1180.46
R7359 VGND.n2671 VGND.n2670 1180.46
R7360 VGND.n2673 VGND.n2672 1180.46
R7361 VGND.n2717 VGND.n2716 1180.46
R7362 VGND.n2719 VGND.n2718 1180.46
R7363 VGND.n2750 VGND.n2749 1180.46
R7364 VGND.n2757 VGND.n2756 1180.46
R7365 VGND.n2755 VGND.n2754 1180.46
R7366 VGND.n2790 VGND.n2789 1180.46
R7367 VGND.n2792 VGND.n2791 1180.46
R7368 VGND.n2345 VGND.n2344 1180.46
R7369 VGND.n2340 VGND.n2339 1180.46
R7370 VGND.n2335 VGND.n2334 1180.46
R7371 VGND.n2330 VGND.n2329 1180.46
R7372 VGND.n2325 VGND.n2324 1180.46
R7373 VGND.n2320 VGND.n2319 1180.46
R7374 VGND.n2315 VGND.n2314 1180.46
R7375 VGND.n2310 VGND.n2309 1180.46
R7376 VGND.n2305 VGND.n2304 1180.46
R7377 VGND.n2300 VGND.n2299 1180.46
R7378 VGND.n2295 VGND.n2294 1180.46
R7379 VGND.n2290 VGND.n2289 1180.46
R7380 VGND.n2545 VGND.n2544 1180.46
R7381 VGND.n2543 VGND.n2542 1180.46
R7382 VGND.n2538 VGND.n2537 1180.46
R7383 VGND.n2355 VGND.n2354 1180.46
R7384 VGND.n2379 VGND.n2378 1180.46
R7385 VGND.n2381 VGND.n2380 1180.46
R7386 VGND.n2405 VGND.n2404 1180.46
R7387 VGND.n2407 VGND.n2406 1180.46
R7388 VGND.n2431 VGND.n2430 1180.46
R7389 VGND.n2433 VGND.n2432 1180.46
R7390 VGND.n2457 VGND.n2456 1180.46
R7391 VGND.n2459 VGND.n2458 1180.46
R7392 VGND.n2483 VGND.n2482 1180.46
R7393 VGND.n2485 VGND.n2484 1180.46
R7394 VGND.n2514 VGND.n2513 1180.46
R7395 VGND.n2519 VGND.n2518 1180.46
R7396 VGND.n2524 VGND.n2523 1180.46
R7397 VGND.n2526 VGND.n2525 1180.46
R7398 VGND.n2366 VGND.n2365 1180.46
R7399 VGND.n2368 VGND.n2367 1180.46
R7400 VGND.n2392 VGND.n2391 1180.46
R7401 VGND.n2394 VGND.n2393 1180.46
R7402 VGND.n2418 VGND.n2417 1180.46
R7403 VGND.n2420 VGND.n2419 1180.46
R7404 VGND.n2444 VGND.n2443 1180.46
R7405 VGND.n2446 VGND.n2445 1180.46
R7406 VGND.n2470 VGND.n2469 1180.46
R7407 VGND.n2472 VGND.n2471 1180.46
R7408 VGND.n2496 VGND.n2495 1180.46
R7409 VGND.n2503 VGND.n2502 1180.46
R7410 VGND.n2501 VGND.n2500 1180.46
R7411 VGND.n2812 VGND.n2811 1180.46
R7412 VGND.n2814 VGND.n2813 1180.46
R7413 VGND.n1913 VGND.n1912 1180.46
R7414 VGND.n1915 VGND.n1914 1180.46
R7415 VGND.n1924 VGND.n1923 1180.46
R7416 VGND.n1926 VGND.n1925 1180.46
R7417 VGND.n1935 VGND.n1934 1180.46
R7418 VGND.n1937 VGND.n1936 1180.46
R7419 VGND.n1946 VGND.n1945 1180.46
R7420 VGND.n1948 VGND.n1947 1180.46
R7421 VGND.n1957 VGND.n1956 1180.46
R7422 VGND.n1959 VGND.n1958 1180.46
R7423 VGND.n1968 VGND.n1967 1180.46
R7424 VGND.n1970 VGND.n1969 1180.46
R7425 VGND.n1979 VGND.n1978 1180.46
R7426 VGND.n1984 VGND.n1983 1180.46
R7427 VGND.n1986 VGND.n1985 1180.46
R7428 VGND.n599 VGND.n598 1180.46
R7429 VGND.n2060 VGND.n2059 1180.46
R7430 VGND.n2058 VGND.n2057 1180.46
R7431 VGND.n2053 VGND.n2052 1180.46
R7432 VGND.n2048 VGND.n2047 1180.46
R7433 VGND.n2043 VGND.n2042 1180.46
R7434 VGND.n2038 VGND.n2037 1180.46
R7435 VGND.n2033 VGND.n2032 1180.46
R7436 VGND.n2028 VGND.n2027 1180.46
R7437 VGND.n2023 VGND.n2022 1180.46
R7438 VGND.n2018 VGND.n2017 1180.46
R7439 VGND.n2013 VGND.n2012 1180.46
R7440 VGND.n2008 VGND.n2007 1180.46
R7441 VGND.n2003 VGND.n2002 1180.46
R7442 VGND.n602 VGND.n601 1180.46
R7443 VGND.n2072 VGND.n2071 1180.46
R7444 VGND.n2077 VGND.n2076 1180.46
R7445 VGND.n2082 VGND.n2081 1180.46
R7446 VGND.n2087 VGND.n2086 1180.46
R7447 VGND.n2092 VGND.n2091 1180.46
R7448 VGND.n2097 VGND.n2096 1180.46
R7449 VGND.n2102 VGND.n2101 1180.46
R7450 VGND.n2107 VGND.n2106 1180.46
R7451 VGND.n2112 VGND.n2111 1180.46
R7452 VGND.n2117 VGND.n2116 1180.46
R7453 VGND.n2122 VGND.n2121 1180.46
R7454 VGND.n2129 VGND.n2128 1180.46
R7455 VGND.n2127 VGND.n2126 1180.46
R7456 VGND.n2837 VGND.n2836 1180.46
R7457 VGND.n2839 VGND.n2838 1180.46
R7458 VGND.n2179 VGND.n2178 1180.46
R7459 VGND.n1754 VGND.n550 1180.46
R7460 VGND.n1764 VGND.n1763 1180.46
R7461 VGND.n1766 VGND.n1765 1180.46
R7462 VGND.n1775 VGND.n1774 1180.46
R7463 VGND.n1777 VGND.n1776 1180.46
R7464 VGND.n1786 VGND.n1785 1180.46
R7465 VGND.n1788 VGND.n1787 1180.46
R7466 VGND.n1797 VGND.n1796 1180.46
R7467 VGND.n1799 VGND.n1798 1180.46
R7468 VGND.n1808 VGND.n1807 1180.46
R7469 VGND.n1810 VGND.n1809 1180.46
R7470 VGND.n1819 VGND.n1818 1180.46
R7471 VGND.n1824 VGND.n1823 1180.46
R7472 VGND.n1826 VGND.n1825 1180.46
R7473 VGND.n1681 VGND.n1680 1180.46
R7474 VGND.n1683 VGND.n1682 1180.46
R7475 VGND.n1692 VGND.n1691 1180.46
R7476 VGND.n1697 VGND.n1696 1180.46
R7477 VGND.n1702 VGND.n1701 1180.46
R7478 VGND.n1707 VGND.n1706 1180.46
R7479 VGND.n1712 VGND.n1711 1180.46
R7480 VGND.n1717 VGND.n1716 1180.46
R7481 VGND.n1722 VGND.n1721 1180.46
R7482 VGND.n1727 VGND.n1726 1180.46
R7483 VGND.n1732 VGND.n1731 1180.46
R7484 VGND.n1850 VGND.n1849 1180.46
R7485 VGND.n1848 VGND.n1847 1180.46
R7486 VGND.n1843 VGND.n1842 1180.46
R7487 VGND.n1735 VGND.n1734 1180.46
R7488 VGND.n672 VGND.n671 1180.46
R7489 VGND.n677 VGND.n676 1180.46
R7490 VGND.n682 VGND.n681 1180.46
R7491 VGND.n687 VGND.n686 1180.46
R7492 VGND.n692 VGND.n691 1180.46
R7493 VGND.n697 VGND.n696 1180.46
R7494 VGND.n702 VGND.n701 1180.46
R7495 VGND.n707 VGND.n706 1180.46
R7496 VGND.n712 VGND.n711 1180.46
R7497 VGND.n717 VGND.n716 1180.46
R7498 VGND.n722 VGND.n721 1180.46
R7499 VGND.n729 VGND.n728 1180.46
R7500 VGND.n727 VGND.n726 1180.46
R7501 VGND.n2862 VGND.n2861 1180.46
R7502 VGND.n2864 VGND.n2863 1180.46
R7503 VGND.n1355 VGND.n1354 1180.46
R7504 VGND.n877 VGND.n876 1180.46
R7505 VGND.n872 VGND.n871 1180.46
R7506 VGND.n821 VGND.n808 1180.46
R7507 VGND.n826 VGND.n825 1180.46
R7508 VGND.n831 VGND.n830 1180.46
R7509 VGND.n836 VGND.n835 1180.46
R7510 VGND.n841 VGND.n840 1180.46
R7511 VGND.n846 VGND.n845 1180.46
R7512 VGND.n851 VGND.n850 1180.46
R7513 VGND.n858 VGND.n857 1180.46
R7514 VGND.n856 VGND.n855 1180.46
R7515 VGND.n1666 VGND.n1665 1180.46
R7516 VGND.n1664 VGND.n1663 1180.46
R7517 VGND.n1659 VGND.n1658 1180.46
R7518 VGND.n1393 VGND.n1392 1180.46
R7519 VGND.n1398 VGND.n1397 1180.46
R7520 VGND.n1400 VGND.n1399 1180.46
R7521 VGND.n1493 VGND.n1492 1180.46
R7522 VGND.n1495 VGND.n1494 1180.46
R7523 VGND.n1519 VGND.n1518 1180.46
R7524 VGND.n1521 VGND.n1520 1180.46
R7525 VGND.n1545 VGND.n1544 1180.46
R7526 VGND.n1550 VGND.n1549 1180.46
R7527 VGND.n1557 VGND.n1556 1180.46
R7528 VGND.n1555 VGND.n1554 1180.46
R7529 VGND.n1635 VGND.n1634 1180.46
R7530 VGND.n1640 VGND.n1639 1180.46
R7531 VGND.n1645 VGND.n1644 1180.46
R7532 VGND.n1647 VGND.n1646 1180.46
R7533 VGND.n1413 VGND.n1412 1180.46
R7534 VGND.n1415 VGND.n1414 1180.46
R7535 VGND.n1480 VGND.n1479 1180.46
R7536 VGND.n1482 VGND.n1481 1180.46
R7537 VGND.n1506 VGND.n1505 1180.46
R7538 VGND.n1508 VGND.n1507 1180.46
R7539 VGND.n1532 VGND.n1531 1180.46
R7540 VGND.n1534 VGND.n1533 1180.46
R7541 VGND.n1569 VGND.n1568 1180.46
R7542 VGND.n1586 VGND.n1585 1180.46
R7543 VGND.n1584 VGND.n1583 1180.46
R7544 VGND.n1579 VGND.n1578 1180.46
R7545 VGND.n1574 VGND.n1573 1180.46
R7546 VGND.n2887 VGND.n2886 1180.46
R7547 VGND.n2889 VGND.n2888 1180.46
R7548 VGND.n1342 VGND.n1341 1180.46
R7549 VGND.n1426 VGND.n1425 1180.46
R7550 VGND.n1431 VGND.n1430 1180.46
R7551 VGND.n1436 VGND.n1435 1180.46
R7552 VGND.n1441 VGND.n1440 1180.46
R7553 VGND.n1446 VGND.n1445 1180.46
R7554 VGND.n1451 VGND.n1450 1180.46
R7555 VGND.n1456 VGND.n1455 1180.46
R7556 VGND.n1463 VGND.n1462 1180.46
R7557 VGND.n1461 VGND.n1460 1180.46
R7558 VGND.n1598 VGND.n1597 1180.46
R7559 VGND.n1603 VGND.n1602 1180.46
R7560 VGND.n1618 VGND.n1617 1180.46
R7561 VGND.n1616 VGND.n1615 1180.46
R7562 VGND.n1611 VGND.n1610 1180.46
R7563 VGND.n1034 VGND.n1033 1180.46
R7564 VGND.n1039 VGND.n1038 1180.46
R7565 VGND.n1099 VGND.n1098 1180.46
R7566 VGND.n1097 VGND.n1096 1180.46
R7567 VGND.n1092 VGND.n1091 1180.46
R7568 VGND.n1087 VGND.n1086 1180.46
R7569 VGND.n1082 VGND.n1081 1180.46
R7570 VGND.n1077 VGND.n1076 1180.46
R7571 VGND.n1072 VGND.n1071 1180.46
R7572 VGND.n1050 VGND.n1041 1180.46
R7573 VGND.n1055 VGND.n1054 1180.46
R7574 VGND.n1060 VGND.n1059 1180.46
R7575 VGND.n1062 VGND.n1061 1180.46
R7576 VGND.n2907 VGND.n2906 1180.46
R7577 VGND.n2909 VGND.n2908 1180.46
R7578 VGND.t1002 VGND.n3011 1180.08
R7579 VGND.n1387 VGND.n1386 1169.57
R7580 VGND.n3015 VGND.t2547 1146.36
R7581 VGND.n3017 VGND.t2546 1112.64
R7582 VGND.n3016 VGND.t1062 1112.64
R7583 VGND.n2351 VGND.n2349 1070.21
R7584 VGND.n2968 VGND 1055.35
R7585 VGND.n2251 VGND.n2250 1052.29
R7586 VGND.t657 VGND.n2181 1032.59
R7587 VGND.t2056 VGND.n2641 988.926
R7588 VGND.t1081 VGND.n2646 988.926
R7589 VGND.t1829 VGND.n2651 988.926
R7590 VGND.t2491 VGND.n2656 988.926
R7591 VGND.t2564 VGND.n2661 988.926
R7592 VGND.t2361 VGND.n2666 988.926
R7593 VGND.t552 VGND.n2671 988.926
R7594 VGND.n2672 VGND.t426 988.926
R7595 VGND.t1534 VGND.n2717 988.926
R7596 VGND.n2718 VGND.t932 988.926
R7597 VGND.t959 VGND.n2750 988.926
R7598 VGND.n2756 VGND.t1446 988.926
R7599 VGND.n2755 VGND.t91 988.926
R7600 VGND.t1471 VGND.n2790 988.926
R7601 VGND.n2791 VGND.t343 988.926
R7602 VGND.n2345 VGND.t2519 988.926
R7603 VGND.n2340 VGND.t1307 988.926
R7604 VGND.n2335 VGND.t1856 988.926
R7605 VGND.n2330 VGND.t235 988.926
R7606 VGND.n2325 VGND.t1244 988.926
R7607 VGND.n2320 VGND.t1175 988.926
R7608 VGND.n2315 VGND.t577 988.926
R7609 VGND.n2310 VGND.t719 988.926
R7610 VGND.n2305 VGND.t713 988.926
R7611 VGND.n2300 VGND.t65 988.926
R7612 VGND.n2295 VGND.t1208 988.926
R7613 VGND.n2290 VGND.t1463 988.926
R7614 VGND.n2544 VGND.t546 988.926
R7615 VGND.n2543 VGND.t2034 988.926
R7616 VGND.n2538 VGND.t1524 988.926
R7617 VGND.n2354 VGND.t2043 988.926
R7618 VGND.t1048 VGND.n2379 988.926
R7619 VGND.n2380 VGND.t1869 988.926
R7620 VGND.t2498 VGND.n2405 988.926
R7621 VGND.n2406 VGND.t2570 988.926
R7622 VGND.t1364 VGND.n2431 988.926
R7623 VGND.n2432 VGND.t558 988.926
R7624 VGND.t767 VGND.n2457 988.926
R7625 VGND.n2458 VGND.t218 988.926
R7626 VGND.t1127 VGND.n2483 988.926
R7627 VGND.n2484 VGND.t1026 988.926
R7628 VGND.t1154 VGND.n2514 988.926
R7629 VGND.t97 VGND.n2519 988.926
R7630 VGND.t673 VGND.n2524 988.926
R7631 VGND.n2525 VGND.t350 988.926
R7632 VGND.t745 VGND.n2366 988.926
R7633 VGND.n2367 VGND.t2247 988.926
R7634 VGND.t1839 VGND.n2392 988.926
R7635 VGND.n2393 VGND.t2288 988.926
R7636 VGND.t1421 VGND.n2418 988.926
R7637 VGND.n2419 VGND.t1387 988.926
R7638 VGND.t418 VGND.n2444 988.926
R7639 VGND.n2445 VGND.t2542 988.926
R7640 VGND.t759 VGND.n2470 988.926
R7641 VGND.n2471 VGND.t592 988.926
R7642 VGND.t683 VGND.n2496 988.926
R7643 VGND.n2502 VGND.t432 988.926
R7644 VGND.n2501 VGND.t1262 988.926
R7645 VGND.t622 VGND.n2812 988.926
R7646 VGND.n2813 VGND.t32 988.926
R7647 VGND.t1017 VGND.n1913 988.926
R7648 VGND.n1914 VGND.t2075 988.926
R7649 VGND.t1861 VGND.n1924 988.926
R7650 VGND.n1925 VGND.t228 988.926
R7651 VGND.t1122 VGND.n1935 988.926
R7652 VGND.n1936 VGND.t2259 988.926
R7653 VGND.t5 VGND.n1946 988.926
R7654 VGND.n1947 VGND.t239 988.926
R7655 VGND.t404 VGND.n1957 988.926
R7656 VGND.n1958 VGND.t60 988.926
R7657 VGND.t2677 VGND.n1968 988.926
R7658 VGND.n1969 VGND.t1043 988.926
R7659 VGND.t540 VGND.n1979 988.926
R7660 VGND.t1520 VGND.n1984 988.926
R7661 VGND.n1985 VGND.t442 988.926
R7662 VGND.t2054 VGND.n599 988.926
R7663 VGND.n2059 VGND.t1079 988.926
R7664 VGND.n2058 VGND.t1832 988.926
R7665 VGND.n2053 VGND.t2489 988.926
R7666 VGND.n2048 VGND.t2562 988.926
R7667 VGND.n2043 VGND.t2359 988.926
R7668 VGND.n2038 VGND.t550 988.926
R7669 VGND.n2033 VGND.t424 988.926
R7670 VGND.n2028 VGND.t1532 988.926
R7671 VGND.n2023 VGND.t929 988.926
R7672 VGND.n2018 VGND.t957 988.926
R7673 VGND.n2013 VGND.t1443 988.926
R7674 VGND.n2008 VGND.t89 988.926
R7675 VGND.n2003 VGND.t1515 988.926
R7676 VGND.n601 VGND.t341 988.926
R7677 VGND.t2045 VGND.n2072 988.926
R7678 VGND.t1050 VGND.n2077 988.926
R7679 VGND.t1867 VGND.n2082 988.926
R7680 VGND.t2500 VGND.n2087 988.926
R7681 VGND.t2559 VGND.n2092 988.926
R7682 VGND.t1366 VGND.n2097 988.926
R7683 VGND.t0 VGND.n2102 988.926
R7684 VGND.t769 VGND.n2107 988.926
R7685 VGND.t220 VGND.n2112 988.926
R7686 VGND.t1129 VGND.n2117 988.926
R7687 VGND.t1028 VGND.n2122 988.926
R7688 VGND.n2128 VGND.t1156 988.926
R7689 VGND.n2127 VGND.t99 988.926
R7690 VGND.t675 VGND.n2837 988.926
R7691 VGND.n2838 VGND.t352 988.926
R7692 VGND.n2179 VGND.t747 988.926
R7693 VGND.t2249 VGND.n1754 988.926
R7694 VGND.t1837 VGND.n1764 988.926
R7695 VGND.n1765 VGND.t2290 988.926
R7696 VGND.t1423 VGND.n1775 988.926
R7697 VGND.n1776 VGND.t1389 988.926
R7698 VGND.t420 VGND.n1786 988.926
R7699 VGND.n1787 VGND.t2544 988.926
R7700 VGND.t761 VGND.n1797 988.926
R7701 VGND.n1798 VGND.t594 988.926
R7702 VGND.t685 VGND.n1808 988.926
R7703 VGND.n1809 VGND.t434 988.926
R7704 VGND.t1264 VGND.n1819 988.926
R7705 VGND.t624 VGND.n1824 988.926
R7706 VGND.n1825 VGND.t34 988.926
R7707 VGND.t740 VGND.n1681 988.926
R7708 VGND.n1682 VGND.t1166 988.926
R7709 VGND.t1843 VGND.n1692 988.926
R7710 VGND.t214 VGND.n1697 988.926
R7711 VGND.t703 VGND.n1702 988.926
R7712 VGND.t1385 VGND.n1707 988.926
R7713 VGND.t414 VGND.n1712 988.926
R7714 VGND.t2538 VGND.n1717 988.926
R7715 VGND.t568 VGND.n1722 988.926
R7716 VGND.t590 VGND.n1727 988.926
R7717 VGND.t1141 VGND.n1732 988.926
R7718 VGND.n1849 VGND.t430 988.926
R7719 VGND.n1848 VGND.t637 988.926
R7720 VGND.n1843 VGND.t618 988.926
R7721 VGND.n1734 VGND.t30 988.926
R7722 VGND.t1015 VGND.n672 988.926
R7723 VGND.t2073 VGND.n677 988.926
R7724 VGND.t1863 VGND.n682 988.926
R7725 VGND.t226 VGND.n687 988.926
R7726 VGND.t1120 VGND.n692 988.926
R7727 VGND.t2257 VGND.n697 988.926
R7728 VGND.t3 VGND.n702 988.926
R7729 VGND.t237 VGND.n707 988.926
R7730 VGND.t402 VGND.n712 988.926
R7731 VGND.t1133 VGND.n717 988.926
R7732 VGND.t2675 VGND.n722 988.926
R7733 VGND.n728 VGND.t1041 988.926
R7734 VGND.n727 VGND.t538 988.926
R7735 VGND.t1518 VGND.n2862 988.926
R7736 VGND.n2863 VGND.t440 988.926
R7737 VGND.n1355 VGND.t1070 988.926
R7738 VGND.n877 VGND.t1097 988.926
R7739 VGND.n872 VGND.t1847 988.926
R7740 VGND.t208 VGND.n821 988.926
R7741 VGND.t572 VGND.n826 988.926
R7742 VGND.t1182 VGND.n831 988.926
R7743 VGND.t407 VGND.n836 988.926
R7744 VGND.t772 VGND.n841 988.926
R7745 VGND.t2484 VGND.n846 988.926
R7746 VGND.t2023 VGND.n851 988.926
R7747 VGND.n857 VGND.t2124 988.926
R7748 VGND.n856 VGND.t2343 988.926
R7749 VGND.n1665 VGND.t2477 988.926
R7750 VGND.n1664 VGND.t2027 988.926
R7751 VGND.n1659 VGND.t22 988.926
R7752 VGND.t2041 VGND.n1393 988.926
R7753 VGND.t1046 VGND.n1398 988.926
R7754 VGND.n1399 VGND.t1871 988.926
R7755 VGND.t2496 VGND.n1493 988.926
R7756 VGND.n1494 VGND.t2568 988.926
R7757 VGND.t1362 VGND.n1519 988.926
R7758 VGND.n1520 VGND.t556 988.926
R7759 VGND.t765 VGND.n1545 988.926
R7760 VGND.t1538 VGND.n1550 988.926
R7761 VGND.n1556 VGND.t936 988.926
R7762 VGND.n1555 VGND.t1024 988.926
R7763 VGND.t1152 VGND.n1635 988.926
R7764 VGND.t95 VGND.n1640 988.926
R7765 VGND.t1475 VGND.n1645 988.926
R7766 VGND.n1646 VGND.t348 988.926
R7767 VGND.t1068 VGND.n1413 988.926
R7768 VGND.n1414 VGND.t1095 988.926
R7769 VGND.t1849 VGND.n1480 988.926
R7770 VGND.n1481 VGND.t2071 988.926
R7771 VGND.t1553 VGND.n1506 988.926
R7772 VGND.n1507 VGND.t1180 988.926
R7773 VGND.t583 VGND.n1532 988.926
R7774 VGND.n1533 VGND.t2532 988.926
R7775 VGND.t2482 VGND.n1569 988.926
R7776 VGND.n1585 VGND.t2021 988.926
R7777 VGND.n1584 VGND.t2122 988.926
R7778 VGND.n1579 VGND.t2095 988.926
R7779 VGND.n1574 VGND.t2475 988.926
R7780 VGND.t628 VGND.n2887 988.926
R7781 VGND.n2888 VGND.t2286 988.926
R7782 VGND.n1341 VGND.t2517 988.926
R7783 VGND.t1305 VGND.n1426 988.926
R7784 VGND.t1859 VGND.n1431 988.926
R7785 VGND.t232 VGND.n1436 988.926
R7786 VGND.t1242 VGND.n1441 988.926
R7787 VGND.t1173 VGND.n1446 988.926
R7788 VGND.t575 VGND.n1451 988.926
R7789 VGND.t717 VGND.n1456 988.926
R7790 VGND.n1462 VGND.t711 988.926
R7791 VGND.n1461 VGND.t62 988.926
R7792 VGND.t1206 VGND.n1598 988.926
R7793 VGND.t1460 VGND.n1603 988.926
R7794 VGND.n1617 VGND.t544 988.926
R7795 VGND.n1616 VGND.t2031 988.926
R7796 VGND.n1611 VGND.t446 988.926
R7797 VGND.t742 VGND.n1034 988.926
R7798 VGND.t1168 VGND.n1039 988.926
R7799 VGND.n1098 VGND.t1841 988.926
R7800 VGND.n1097 VGND.t216 988.926
R7801 VGND.n1092 VGND.t705 988.926
R7802 VGND.n1087 VGND.t1383 988.926
R7803 VGND.n1082 VGND.t412 988.926
R7804 VGND.n1077 VGND.t2536 988.926
R7805 VGND.n1072 VGND.t566 988.926
R7806 VGND.t588 VGND.n1050 988.926
R7807 VGND.t1139 VGND.n1055 988.926
R7808 VGND.t2347 VGND.n1060 988.926
R7809 VGND.n1061 VGND.t635 988.926
R7810 VGND.t620 VGND.n2907 988.926
R7811 VGND.n2908 VGND.t28 988.926
R7812 VGND.n1335 VGND.t1627 988.926
R7813 VGND.t1709 VGND.n929 988.926
R7814 VGND.t1731 VGND.n934 988.926
R7815 VGND.t1632 VGND.n939 988.926
R7816 VGND.t1643 VGND.n944 988.926
R7817 VGND.t1662 VGND.n949 988.926
R7818 VGND.t1803 VGND.n954 988.926
R7819 VGND.t1824 VGND.n959 988.926
R7820 VGND.t1666 VGND.n964 988.926
R7821 VGND.t1743 VGND.n969 988.926
R7822 VGND.t1756 VGND.n974 988.926
R7823 VGND.t1608 VGND.n979 988.926
R7824 VGND.t1683 VGND.n984 988.926
R7825 VGND.t1774 VGND.n989 988.926
R7826 VGND.n990 VGND.t1599 988.926
R7827 VGND.n2248 VGND.n539 934.784
R7828 VGND.n116 VGND 927.203
R7829 VGND.n134 VGND 927.203
R7830 VGND.n2182 VGND 918.774
R7831 VGND.n194 VGND 910.346
R7832 VGND.n165 VGND 910.346
R7833 VGND.t2119 VGND.n2967 909.365
R7834 VGND.n2285 VGND.n473 900
R7835 VGND.n2641 VGND.t1555 852.769
R7836 VGND.n2646 VGND.t561 852.769
R7837 VGND.n2651 VGND.t196 852.769
R7838 VGND.n2656 VGND.t1368 852.769
R7839 VGND.n2661 VGND.t778 852.769
R7840 VGND.n2666 VGND.t187 852.769
R7841 VGND.n2671 VGND.t564 852.769
R7842 VGND.n2672 VGND.t1019 852.769
R7843 VGND.n2717 VGND.t1440 852.769
R7844 VGND.n2718 VGND.t2401 852.769
R7845 VGND.n2750 VGND.t205 852.769
R7846 VGND.n2756 VGND.t105 852.769
R7847 VGND.t1000 VGND.n2755 852.769
R7848 VGND.n2790 VGND.t1228 852.769
R7849 VGND.n2791 VGND.t1066 852.769
R7850 VGND.n2935 VGND.t2407 852.769
R7851 VGND.t600 VGND.n2345 852.769
R7852 VGND.t115 VGND.n2340 852.769
R7853 VGND.t1381 VGND.n2335 852.769
R7854 VGND.t2522 VGND.n2330 852.769
R7855 VGND.t1449 VGND.n2325 852.769
R7856 VGND.t2070 VGND.n2320 852.769
R7857 VGND.t2048 VGND.n2315 852.769
R7858 VGND.t1020 VGND.n2310 852.769
R7859 VGND.t2342 VGND.n2305 852.769
R7860 VGND.t783 VGND.n2300 852.769
R7861 VGND.t1230 VGND.n2295 852.769
R7862 VGND.t2648 VGND.n2290 852.769
R7863 VGND.n2544 VGND.t2649 852.769
R7864 VGND.t2051 VGND.n2543 852.769
R7865 VGND.t696 VGND.n2538 852.769
R7866 VGND.t780 VGND.n208 852.769
R7867 VGND.n2354 VGND.t1397 852.769
R7868 VGND.n2379 VGND.t186 852.769
R7869 VGND.n2380 VGND.t2380 852.769
R7870 VGND.n2405 VGND.t45 852.769
R7871 VGND.n2406 VGND.t757 852.769
R7872 VGND.n2431 VGND.t948 852.769
R7873 VGND.n2432 VGND.t1187 852.769
R7874 VGND.n2457 VGND.t2524 852.769
R7875 VGND.n2458 VGND.t113 852.769
R7876 VGND.n2483 VGND.t938 852.769
R7877 VGND.n2484 VGND.t1087 852.769
R7878 VGND.n2514 VGND.t1315 852.769
R7879 VGND.n2519 VGND.t118 852.769
R7880 VGND.n2524 VGND.t2403 852.769
R7881 VGND.n2525 VGND.t2514 852.769
R7882 VGND.t2550 VGND.n209 852.769
R7883 VGND.n2366 VGND.t949 852.769
R7884 VGND.n2367 VGND.t994 852.769
R7885 VGND.n2392 VGND.t1199 852.769
R7886 VGND.n2393 VGND.t1458 852.769
R7887 VGND.n2418 VGND.t1006 852.769
R7888 VGND.n2419 VGND.t1324 852.769
R7889 VGND.n2444 VGND.t679 852.769
R7890 VGND.n2445 VGND.t19 852.769
R7891 VGND.n2470 VGND.t1459 852.769
R7892 VGND.n2471 VGND.t950 852.769
R7893 VGND.n2496 VGND.t1189 852.769
R7894 VGND.n2502 VGND.t1229 852.769
R7895 VGND.t81 VGND.n2501 852.769
R7896 VGND.n2812 VGND.t1205 852.769
R7897 VGND.n2813 VGND.t2398 852.769
R7898 VGND.t955 VGND.n210 852.769
R7899 VGND.n1913 VGND.t120 852.769
R7900 VGND.n1914 VGND.t699 852.769
R7901 VGND.n1924 VGND.t1008 852.769
R7902 VGND.n1925 VGND.t1190 852.769
R7903 VGND.n1935 VGND.t656 852.769
R7904 VGND.n1936 VGND.t617 852.769
R7905 VGND.n1946 VGND.t134 852.769
R7906 VGND.n1947 VGND.t2357 852.769
R7907 VGND.n1957 VGND.t698 852.769
R7908 VGND.n1958 VGND.t1084 852.769
R7909 VGND.n1968 VGND.t2534 852.769
R7910 VGND.n1969 VGND.t2512 852.769
R7911 VGND.n1979 VGND.t2406 852.769
R7912 VGND.n1984 VGND.t116 852.769
R7913 VGND.n1985 VGND.t2061 852.769
R7914 VGND.t2368 VGND.n211 852.769
R7915 VGND.n599 VGND.t2039 852.769
R7916 VGND.n2059 VGND.t2551 852.769
R7917 VGND.t185 VGND.n2058 852.769
R7918 VGND.t13 VGND.n2053 852.769
R7919 VGND.t1442 VGND.n2048 852.769
R7920 VGND.t1301 VGND.n2043 852.769
R7921 VGND.t2052 VGND.n2038 852.769
R7922 VGND.t996 VGND.n2033 852.769
R7923 VGND.t193 VGND.n2028 852.769
R7924 VGND.t2589 VGND.n2023 852.769
R7925 VGND.t1093 VGND.n2018 852.769
R7926 VGND.t1470 VGND.n2013 852.769
R7927 VGND.t1005 VGND.n2008 852.769
R7928 VGND.t631 VGND.n2003 852.769
R7929 VGND.n601 VGND.t2408 852.769
R7930 VGND.t991 VGND.n212 852.769
R7931 VGND.n2072 VGND.t777 852.769
R7932 VGND.n2077 VGND.t1085 852.769
R7933 VGND.n2082 VGND.t680 852.769
R7934 VGND.n2087 VGND.t2679 852.769
R7935 VGND.n2092 VGND.t2365 852.769
R7936 VGND.n2097 VGND.t11 852.769
R7937 VGND.n2102 VGND.t672 852.769
R7938 VGND.n2107 VGND.t2527 852.769
R7939 VGND.n2112 VGND.t112 852.769
R7940 VGND.n2117 VGND.t58 852.769
R7941 VGND.n2122 VGND.t2038 852.769
R7942 VGND.n2128 VGND.t1226 852.769
R7943 VGND.t1874 VGND.n2127 852.769
R7944 VGND.n2837 VGND.t1439 852.769
R7945 VGND.n2838 VGND.t563 852.769
R7946 VGND.t1302 VGND.n213 852.769
R7947 VGND.t670 VGND.n2179 852.769
R7948 VGND.n1754 VGND.t1109 852.769
R7949 VGND.n1764 VGND.t1246 852.769
R7950 VGND.n1765 VGND.t954 852.769
R7951 VGND.n1775 VGND.t197 852.769
R7952 VGND.n1776 VGND.t1217 852.769
R7953 VGND.n1786 VGND.t2588 852.769
R7954 VGND.n1787 VGND.t189 852.769
R7955 VGND.n1797 VGND.t2655 852.769
R7956 VGND.n1798 VGND.t1530 852.769
R7957 VGND.n1808 VGND.t1030 852.769
R7958 VGND.n1809 VGND.t2404 852.769
R7959 VGND.n1819 VGND.t1188 852.769
R7960 VGND.n1824 VGND.t104 852.769
R7961 VGND.n1825 VGND.t2101 852.769
R7962 VGND.t1107 VGND.n214 852.769
R7963 VGND.n1681 VGND.t2409 852.769
R7964 VGND.n1682 VGND.t121 852.769
R7965 VGND.n1692 VGND.t1334 852.769
R7966 VGND.n1697 VGND.t1065 852.769
R7967 VGND.n1702 VGND.t2374 852.769
R7968 VGND.n1707 VGND.t102 852.769
R7969 VGND.n1712 VGND.t2395 852.769
R7970 VGND.n1717 VGND.t2375 852.769
R7971 VGND.n1722 VGND.t2369 852.769
R7972 VGND.n1727 VGND.t2509 852.769
R7973 VGND.n1732 VGND.t106 852.769
R7974 VGND.n1849 VGND.t2513 852.769
R7975 VGND.t944 VGND.n1848 852.769
R7976 VGND.t1001 VGND.n1843 852.769
R7977 VGND.n1734 VGND.t110 852.769
R7978 VGND.t2372 VGND.n215 852.769
R7979 VGND.n672 VGND.t1266 852.769
R7980 VGND.n677 VGND.t114 852.769
R7981 VGND.n682 VGND.t1007 852.769
R7982 VGND.n687 VGND.t585 852.769
R7983 VGND.n692 VGND.t1526 852.769
R7984 VGND.n697 VGND.t599 852.769
R7985 VGND.n702 VGND.t2355 852.769
R7986 VGND.n707 VGND.t1061 852.769
R7987 VGND.n712 VGND.t2396 852.769
R7988 VGND.n717 VGND.t43 852.769
R7989 VGND.n722 VGND.t1396 852.769
R7990 VGND.n728 VGND.t1522 852.769
R7991 VGND.t2037 VGND.n727 852.769
R7992 VGND.n2862 VGND.t103 852.769
R7993 VGND.n2863 VGND.t1092 852.769
R7994 VGND.t8 VGND.n216 852.769
R7995 VGND.t1160 VGND.n1355 852.769
R7996 VGND.t82 VGND.n877 852.769
R7997 VGND.t1392 VGND.n872 852.769
R7998 VGND.n821 VGND.t1455 852.769
R7999 VGND.n826 VGND.t671 852.769
R8000 VGND.n831 VGND.t2356 852.769
R8001 VGND.n836 VGND.t2174 852.769
R8002 VGND.n841 VGND.t965 852.769
R8003 VGND.n846 VGND.t2511 852.769
R8004 VGND.n851 VGND.t1210 852.769
R8005 VGND.n857 VGND.t2656 852.769
R8006 VGND.t1161 VGND.n856 852.769
R8007 VGND.n1665 VGND.t963 852.769
R8008 VGND.t1438 VGND.n1664 852.769
R8009 VGND.t1010 VGND.n1659 852.769
R8010 VGND.t2353 VGND.n217 852.769
R8011 VGND.n1393 VGND.t2349 852.769
R8012 VGND.n1398 VGND.t2502 852.769
R8013 VGND.n1399 VGND.t2394 852.769
R8014 VGND.n1493 VGND.t44 852.769
R8015 VGND.n1494 VGND.t2650 852.769
R8016 VGND.n1519 VGND.t59 852.769
R8017 VGND.n1520 VGND.t1395 852.769
R8018 VGND.n1545 VGND.t2523 852.769
R8019 VGND.n1550 VGND.t2040 852.769
R8020 VGND.n1556 VGND.t117 852.769
R8021 VGND.t1412 VGND.n1555 852.769
R8022 VGND.n1635 VGND.t2060 852.769
R8023 VGND.n1640 VGND.t1108 852.769
R8024 VGND.n1645 VGND.t993 852.769
R8025 VGND.n1646 VGND.t1089 852.769
R8026 VGND.t660 VGND.n218 852.769
R8027 VGND.n1413 VGND.t1394 852.769
R8028 VGND.n1414 VGND.t2366 852.769
R8029 VGND.n1480 VGND.t781 852.769
R8030 VGND.n1481 VGND.t943 852.769
R8031 VGND.n1506 VGND.t2351 852.769
R8032 VGND.n1507 VGND.t1528 852.769
R8033 VGND.n1532 VGND.t1099 852.769
R8034 VGND.n1533 VGND.t2682 852.769
R8035 VGND.n1569 VGND.t2358 852.769
R8036 VGND.n1585 VGND.t1456 852.769
R8037 VGND.t2402 VGND.n1584 852.769
R8038 VGND.t669 VGND.n1579 852.769
R8039 VGND.t1333 VGND.n1574 852.769
R8040 VGND.n2887 VGND.t782 852.769
R8041 VGND.n2888 VGND.t2399 852.769
R8042 VGND.t2400 VGND.n219 852.769
R8043 VGND.n1341 VGND.t2049 852.769
R8044 VGND.n1426 VGND.t682 852.769
R8045 VGND.n1431 VGND.t18 852.769
R8046 VGND.n1436 VGND.t1009 852.769
R8047 VGND.n1441 VGND.t204 852.769
R8048 VGND.n1446 VGND.t338 852.769
R8049 VGND.n1451 VGND.t108 852.769
R8050 VGND.n1456 VGND.t1227 852.769
R8051 VGND.n1462 VGND.t1457 852.769
R8052 VGND.t2535 VGND.n1461 852.769
R8053 VGND.n1598 VGND.t668 852.769
R8054 VGND.n1603 VGND.t1211 852.769
R8055 VGND.n1617 VGND.t2525 852.769
R8056 VGND.t956 VGND.n1616 852.769
R8057 VGND.t2175 VGND.n1611 852.769
R8058 VGND.t1336 VGND.n220 852.769
R8059 VGND.n1034 VGND.t1437 852.769
R8060 VGND.n1039 VGND.t1090 852.769
R8061 VGND.n1098 VGND.t1309 852.769
R8062 VGND.t107 VGND.n1097 852.769
R8063 VGND.t1212 VGND.n1092 852.769
R8064 VGND.t2397 VGND.n1087 852.769
R8065 VGND.t1527 VGND.n1082 852.769
R8066 VGND.t562 VGND.n1077 852.769
R8067 VGND.t119 VGND.n1072 852.769
R8068 VGND.n1050 VGND.t188 852.769
R8069 VGND.n1055 VGND.t184 852.769
R8070 VGND.n1060 VGND.t632 852.769
R8071 VGND.n1061 VGND.t12 852.769
R8072 VGND.n2907 VGND.t2487 852.769
R8073 VGND.n2908 VGND.t2458 852.769
R8074 VGND.t995 VGND.n221 852.769
R8075 VGND.t2373 VGND.n1335 852.769
R8076 VGND.n929 VGND.t2371 852.769
R8077 VGND.n934 VGND.t135 852.769
R8078 VGND.n939 VGND.t992 852.769
R8079 VGND.n944 VGND.t951 852.769
R8080 VGND.n949 VGND.t2350 852.769
R8081 VGND.n954 VGND.t2510 852.769
R8082 VGND.n959 VGND.t1300 852.769
R8083 VGND.n964 VGND.t2670 852.769
R8084 VGND.n969 VGND.t1398 852.769
R8085 VGND.n974 VGND.t2354 852.769
R8086 VGND.n979 VGND.t2529 852.769
R8087 VGND.n984 VGND.t1088 852.769
R8088 VGND.n989 VGND.t681 852.769
R8089 VGND.n990 VGND.t109 852.769
R8090 VGND.n2918 VGND.t1335 852.769
R8091 VGND.n2249 VGND 851.341
R8092 VGND.n2944 VGND.n2943 846.154
R8093 VGND.n2350 VGND.t1915 809.773
R8094 VGND.n2352 VGND.t1990 809.773
R8095 VGND.t1894 VGND.n2353 809.773
R8096 VGND.n473 VGND.t1939 809.773
R8097 VGND.t2014 VGND.n503 809.773
R8098 VGND.t1891 VGND.n504 809.773
R8099 VGND.n2180 VGND.t1933 809.773
R8100 VGND.t1945 VGND.n539 809.773
R8101 VGND.n1387 VGND.t1969 809.773
R8102 VGND.t1897 VGND.n1388 809.773
R8103 VGND.n1339 VGND.t1972 809.773
R8104 VGND.t1999 VGND.n1340 809.773
R8105 VGND.n1338 VGND.t1942 809.773
R8106 VGND.n1336 VGND.t1788 809.773
R8107 VGND.t861 VGND.t843 708.047
R8108 VGND.t843 VGND.t841 708.047
R8109 VGND.t841 VGND.t851 708.047
R8110 VGND.t851 VGND.t53 708.047
R8111 VGND.t53 VGND.t708 708.047
R8112 VGND.t708 VGND.t1468 708.047
R8113 VGND.t1468 VGND.t1072 708.047
R8114 VGND.t732 VGND.t2546 708.047
R8115 VGND.t857 VGND.t894 708.047
R8116 VGND.t894 VGND.t865 708.047
R8117 VGND.t865 VGND.t839 708.047
R8118 VGND.t839 VGND.t55 708.047
R8119 VGND.t55 VGND.t1299 708.047
R8120 VGND.t1299 VGND.t52 708.047
R8121 VGND.t52 VGND.t947 708.047
R8122 VGND.t910 VGND.t859 708.047
R8123 VGND.t859 VGND.t898 708.047
R8124 VGND.t898 VGND.t868 708.047
R8125 VGND.t868 VGND.t2469 708.047
R8126 VGND.t2469 VGND.t2465 708.047
R8127 VGND.t2465 VGND.t2459 708.047
R8128 VGND.t2459 VGND.t2461 708.047
R8129 VGND.t729 VGND.t2547 708.047
R8130 VGND.t886 VGND.t875 708.047
R8131 VGND.t875 VGND.t873 708.047
R8132 VGND.t873 VGND.t833 708.047
R8133 VGND.t833 VGND.t56 708.047
R8134 VGND.t56 VGND.t47 708.047
R8135 VGND.t47 VGND.t1075 708.047
R8136 VGND.t1075 VGND.t50 708.047
R8137 VGND.t853 VGND.t890 708.047
R8138 VGND.t890 VGND.t863 708.047
R8139 VGND.t863 VGND.t871 708.047
R8140 VGND.t871 VGND.t49 708.047
R8141 VGND.t49 VGND.t223 708.047
R8142 VGND.t223 VGND.t46 708.047
R8143 VGND.t46 VGND.t2016 708.047
R8144 VGND.t849 VGND.t903 708.047
R8145 VGND.t908 VGND.t849 708.047
R8146 VGND.t882 VGND.t908 708.047
R8147 VGND.t2467 VGND.t882 708.047
R8148 VGND.t2463 VGND.t2467 708.047
R8149 VGND.t2468 VGND.t2463 708.047
R8150 VGND.t2464 VGND.t2468 708.047
R8151 VGND.n2971 VGND.n2970 708.047
R8152 VGND.t939 VGND.t1063 691.188
R8153 VGND.t1213 VGND.t2504 691.188
R8154 VGND.t914 VGND.t892 657.471
R8155 VGND.t888 VGND.t2120 657.471
R8156 VGND.t925 VGND.t2116 657.471
R8157 VGND.t877 VGND.t2110 657.471
R8158 VGND.t2276 VGND.t1404 657.471
R8159 VGND.t979 VGND.t1402 657.471
R8160 VGND.t2266 VGND.t1400 657.471
R8161 VGND.t2593 VGND.t989 657.471
R8162 VGND.t892 VGND.t918 654.197
R8163 VGND.t989 VGND.t1540 654.197
R8164 VGND VGND.n194 640.614
R8165 VGND VGND.n134 640.614
R8166 VGND VGND.n165 640.614
R8167 VGND.n2182 VGND 640.614
R8168 VGND.n116 VGND 632.184
R8169 VGND.t536 VGND.t1313 630.62
R8170 VGND.t1164 VGND.t1270 630.62
R8171 VGND.t1845 VGND.t2387 630.62
R8172 VGND.t2488 VGND.t2385 630.62
R8173 VGND.t701 VGND.t534 630.62
R8174 VGND.t1178 VGND.t2106 630.62
R8175 VGND.t410 VGND.t2104 630.62
R8176 VGND.t775 VGND.t532 630.62
R8177 VGND.t530 VGND.t1032 630.62
R8178 VGND.t2026 VGND.t2108 630.62
R8179 VGND.t2383 VGND.t1451 630.62
R8180 VGND.t2346 VGND.t2381 630.62
R8181 VGND.t2102 VGND.t633 630.62
R8182 VGND.t2391 VGND.t2030 630.62
R8183 VGND.t340 VGND.t2389 630.62
R8184 VGND.t528 VGND.t1612 630.62
R8185 VGND.t1331 VGND.t2059 630.62
R8186 VGND.t607 VGND.t1045 630.62
R8187 VGND.t1191 VGND.t1866 630.62
R8188 VGND.t2251 VGND.t231 630.62
R8189 VGND.t1329 VGND.t2567 630.62
R8190 VGND.t603 VGND.t1382 630.62
R8191 VGND.t601 VGND.t555 630.62
R8192 VGND.t1327 VGND.t764 630.62
R8193 VGND.t1325 VGND.t1537 630.62
R8194 VGND.t605 VGND.t1131 630.62
R8195 VGND.t200 VGND.t1138 630.62
R8196 VGND.t198 VGND.t1158 630.62
R8197 VGND.t1197 VGND.t94 630.62
R8198 VGND.t1195 VGND.t677 630.62
R8199 VGND.t1193 VGND.t445 630.62
R8200 VGND.t609 VGND.t1763 630.62
R8201 VGND.t739 VGND.t1053 630.62
R8202 VGND.t1359 VGND.t2245 630.62
R8203 VGND.t1835 VGND.t1414 630.62
R8204 VGND.t1059 VGND.t2494 630.62
R8205 VGND.t707 VGND.t976 630.62
R8206 VGND.t1355 VGND.t1171 630.62
R8207 VGND.t416 VGND.t1353 630.62
R8208 VGND.t974 VGND.t2540 630.62
R8209 VGND.t570 VGND.t972 630.62
R8210 VGND.t1357 VGND.t597 630.62
R8211 VGND.t1453 VGND.t1057 630.62
R8212 VGND.t1055 VGND.t437 630.62
R8213 VGND.t639 VGND.t1351 630.62
R8214 VGND.t1022 VGND.t1418 630.62
R8215 VGND.t346 VGND.t1416 630.62
R8216 VGND.t970 VGND.t1591 630.62
R8217 VGND.t2198 VGND.t1203 630.62
R8218 VGND.t2508 VGND.t2225 630.62
R8219 VGND.t2554 VGND.t1852 630.62
R8220 VGND.t212 VGND.t2204 630.62
R8221 VGND.t694 VGND.t1551 630.62
R8222 VGND.t2255 VGND.t2221 630.62
R8223 VGND.t2219 VGND.t581 630.62
R8224 VGND.t2530 VGND.t692 630.62
R8225 VGND.t690 VGND.t1259 630.62
R8226 VGND.t2019 VGND.t2223 630.62
R8227 VGND.t2202 VGND.t2673 630.62
R8228 VGND.t2093 VGND.t2200 630.62
R8229 VGND.t2217 VGND.t2473 630.62
R8230 VGND.t2215 VGND.t626 630.62
R8231 VGND.t26 VGND.t2556 630.62
R8232 VGND.t688 VGND.t1657 630.62
R8233 VGND.t2053 VGND.t2196 630.62
R8234 VGND.t1078 VGND.t79 630.62
R8235 VGND.t1337 VGND.t1828 630.62
R8236 VGND.t587 VGND.t1118 630.62
R8237 VGND.t2194 VGND.t1126 630.62
R8238 VGND.t1185 VGND.t75 630.62
R8239 VGND.t73 VGND.t549 630.62
R8240 VGND.t423 VGND.t2192 630.62
R8241 VGND.t2190 VGND.t1531 630.62
R8242 VGND.t934 VGND.t77 630.62
R8243 VGND.t1116 VGND.t1136 630.62
R8244 VGND.t1448 VGND.t1114 630.62
R8245 VGND.t71 VGND.t88 630.62
R8246 VGND.t1473 VGND.t69 630.62
R8247 VGND.t439 VGND.t1339 630.62
R8248 VGND.t2188 VGND.t1791 630.62
R8249 VGND.t1312 VGND.t2233 630.62
R8250 VGND.t1163 VGND.t2683 630.62
R8251 VGND.t2574 VGND.t1846 630.62
R8252 VGND.t2572 VGND.t2292 630.62
R8253 VGND.t2231 VGND.t700 630.62
R8254 VGND.t2584 VGND.t1177 630.62
R8255 VGND.t2582 VGND.t409 630.62
R8256 VGND.t2229 VGND.t774 630.62
R8257 VGND.t2227 VGND.t1031 630.62
R8258 VGND.t2586 VGND.t2025 630.62
R8259 VGND.t2237 VGND.t1450 630.62
R8260 VGND.t2235 VGND.t2345 630.62
R8261 VGND.t2580 VGND.t2479 630.62
R8262 VGND.t2578 VGND.t2029 630.62
R8263 VGND.t339 VGND.t2576 630.62
R8264 VGND.t2685 VGND.t1614 630.62
R8265 VGND.t744 VGND.t648 630.62
R8266 VGND.t2246 VGND.t1239 630.62
R8267 VGND.t1834 VGND.t611 630.62
R8268 VGND.t2495 VGND.t654 630.62
R8269 VGND.t1420 VGND.t646 630.62
R8270 VGND.t1172 VGND.t1235 630.62
R8271 VGND.t417 VGND.t1233 630.62
R8272 VGND.t2541 VGND.t644 630.62
R8273 VGND.t758 VGND.t642 630.62
R8274 VGND.t598 VGND.t1237 630.62
R8275 VGND.t1454 VGND.t652 630.62
R8276 VGND.t1274 VGND.t650 630.62
R8277 VGND.t1231 VGND.t1261 630.62
R8278 VGND.t615 VGND.t1023 630.62
R8279 VGND.t347 VGND.t613 630.62
R8280 VGND.t640 VGND.t1588 630.62
R8281 VGND.t751 VGND.t1204 630.62
R8282 VGND.t1094 VGND.t202 630.62
R8283 VGND.t1851 VGND.t2087 630.62
R8284 VGND.t213 VGND.t2085 630.62
R8285 VGND.t1224 VGND.t1552 630.62
R8286 VGND.t2256 VGND.t2211 630.62
R8287 VGND.t2209 VGND.t582 630.62
R8288 VGND.t2531 VGND.t1222 630.62
R8289 VGND.t1220 VGND.t1260 630.62
R8290 VGND.t2020 VGND.t2213 630.62
R8291 VGND.t755 VGND.t2674 630.62
R8292 VGND.t2094 VGND.t753 630.62
R8293 VGND.t2207 VGND.t2474 630.62
R8294 VGND.t627 VGND.t2091 630.62
R8295 VGND.t27 VGND.t2089 630.62
R8296 VGND.t1218 VGND.t1655 630.62
R8297 VGND.t1201 VGND.t1149 630.62
R8298 VGND.t2507 VGND.t2097 630.62
R8299 VGND.t83 VGND.t1854 630.62
R8300 VGND.t211 VGND.t1037 630.62
R8301 VGND.t1549 VGND.t1147 630.62
R8302 VGND.t2253 VGND.t1347 630.62
R8303 VGND.t580 VGND.t1345 630.62
R8304 VGND.t225 VGND.t1145 630.62
R8305 VGND.t1258 VGND.t1143 630.62
R8306 VGND.t2018 VGND.t1349 630.62
R8307 VGND.t2672 VGND.t1035 630.62
R8308 VGND.t1273 VGND.t1033 630.62
R8309 VGND.t1343 VGND.t2472 630.62
R8310 VGND.t1341 VGND.t953 630.62
R8311 VGND.t24 VGND.t85 630.62
R8312 VGND.t2099 VGND.t1664 630.62
R8313 VGND.t2352 VGND.t1435 630.62
R8314 VGND.t1077 VGND.t1425 630.62
R8315 VGND.t1831 VGND.t1513 630.62
R8316 VGND.t586 VGND.t1511 630.62
R8317 VGND.t1125 VGND.t1433 630.62
R8318 VGND.t1184 VGND.t1503 630.62
R8319 VGND.t548 VGND.t1501 630.62
R8320 VGND.t422 VGND.t1431 630.62
R8321 VGND.t1039 VGND.t1429 630.62
R8322 VGND.t931 VGND.t1505 630.62
R8323 VGND.t1135 VGND.t1509 630.62
R8324 VGND.t1445 VGND.t1507 630.62
R8325 VGND.t1499 VGND.t87 630.62
R8326 VGND.t1497 VGND.t1517 630.62
R8327 VGND.t438 VGND.t1495 630.62
R8328 VGND.t1427 VGND.t1796 630.62
R8329 VGND.t1584 VGND.t2516 630.62
R8330 VGND.t1562 VGND.t1304 630.62
R8331 VGND.t1576 VGND.t1855 630.62
R8332 VGND.t2481 VGND.t1578 630.62
R8333 VGND.t1241 VGND.t1586 630.62
R8334 VGND.t1361 VGND.t1566 630.62
R8335 VGND.t574 VGND.t1568 630.62
R8336 VGND.t716 VGND.t1556 630.62
R8337 VGND.t710 VGND.t1558 630.62
R8338 VGND.t67 VGND.t1564 630.62
R8339 VGND.t962 VGND.t1580 630.62
R8340 VGND.t1582 VGND.t429 630.62
R8341 VGND.t1570 VGND.t543 630.62
R8342 VGND.t1572 VGND.t2036 630.62
R8343 VGND.t1574 VGND.t2285 630.62
R8344 VGND.t1560 VGND.t1705 630.62
R8345 VGND.t1314 VGND.t2663 630.62
R8346 VGND.t1165 VGND.t1283 630.62
R8347 VGND.t1836 VGND.t2064 630.62
R8348 VGND.t2062 VGND.t2493 630.62
R8349 VGND.t702 VGND.t2661 630.62
R8350 VGND.t1279 VGND.t1179 630.62
R8351 VGND.t411 VGND.t1277 630.62
R8352 VGND.t2659 VGND.t776 630.62
R8353 VGND.t565 VGND.t2657 630.62
R8354 VGND.t596 VGND.t1281 630.62
R8355 VGND.t2667 VGND.t1452 630.62
R8356 VGND.t2665 VGND.t436 630.62
R8357 VGND.t634 VGND.t1275 630.62
R8358 VGND.t1021 VGND.t2068 630.62
R8359 VGND.t345 VGND.t2066 630.62
R8360 VGND.t1285 VGND.t1594 630.62
R8361 VGND.t1316 VGND.t2515 630.62
R8362 VGND.t1303 VGND.t1371 630.62
R8363 VGND.t2176 VGND.t1858 630.62
R8364 VGND.t2480 VGND.t1322 630.62
R8365 VGND.t1379 VGND.t1124 630.62
R8366 VGND.t2363 VGND.t2186 630.62
R8367 VGND.t2184 VGND.t7 630.62
R8368 VGND.t715 VGND.t1377 630.62
R8369 VGND.t1375 VGND.t406 630.62
R8370 VGND.t64 VGND.t1369 630.62
R8371 VGND.t1320 VGND.t961 630.62
R8372 VGND.t1318 VGND.t1462 630.62
R8373 VGND.t2182 VGND.t542 630.62
R8374 VGND.t2180 VGND.t2033 630.62
R8375 VGND.t2284 VGND.t2178 630.62
R8376 VGND.t1373 VGND.t1708 630.62
R8377 VGND.t2058 VGND.t1487 630.62
R8378 VGND.t1291 VGND.t1083 630.62
R8379 VGND.t1873 VGND.t1247 630.62
R8380 VGND.t230 VGND.t1493 630.62
R8381 VGND.t2566 VGND.t1485 630.62
R8382 VGND.t1186 VGND.t1287 630.62
R8383 VGND.t554 VGND.t1255 630.62
R8384 VGND.t763 VGND.t1297 630.62
R8385 VGND.t1536 VGND.t1295 630.62
R8386 VGND.t1289 VGND.t935 630.62
R8387 VGND.t1491 VGND.t1137 630.62
R8388 VGND.t1151 VGND.t1489 630.62
R8389 VGND.t93 VGND.t1253 630.62
R8390 VGND.t1251 VGND.t1474 630.62
R8391 VGND.t1249 VGND.t444 630.62
R8392 VGND.t1293 VGND.t1776 630.62
R8393 VGND.t1202 VGND.t1483 630.62
R8394 VGND.t2506 VGND.t966 630.62
R8395 VGND.t1853 VGND.t721 630.62
R8396 VGND.t2243 VGND.t210 630.62
R8397 VGND.t1481 VGND.t1550 630.62
R8398 VGND.t2081 VGND.t2254 630.62
R8399 VGND.t2079 VGND.t579 630.62
R8400 VGND.t1479 VGND.t224 630.62
R8401 VGND.t1477 VGND.t1257 630.62
R8402 VGND.t68 VGND.t2083 630.62
R8403 VGND.t2671 VGND.t2241 630.62
R8404 VGND.t1272 VGND.t2239 630.62
R8405 VGND.t2471 VGND.t2077 630.62
R8406 VGND.t725 VGND.t952 630.62
R8407 VGND.t25 VGND.t723 630.62
R8408 VGND.t968 VGND.t1665 630.62
R8409 VGND.t1625 VGND.t2047 630.62
R8410 VGND.t1052 VGND.t1706 630.62
R8411 VGND.t1865 VGND.t1785 630.62
R8412 VGND.t234 VGND.t1807 630.62
R8413 VGND.t2561 VGND.t1636 630.62
R8414 VGND.t1391 VGND.t1725 630.62
R8415 VGND.t2 VGND.t1736 630.62
R8416 VGND.t771 VGND.t1640 630.62
R8417 VGND.t222 VGND.t1658 630.62
R8418 VGND.t1132 VGND.t1723 630.62
R8419 VGND.t687 VGND.t1820 630.62
R8420 VGND.t1040 VGND.t1592 630.62
R8421 VGND.t101 VGND.t1741 630.62
R8422 VGND.t678 VGND.t1754 630.62
R8423 VGND.t1523 VGND.t1779 630.62
R8424 VGND.t1679 VGND.t1751 630.62
R8425 VGND.n2704 VGND.n327 615.385
R8426 VGND.n2349 VGND.t190 602.708
R8427 VGND.n3019 VGND.t190 602.708
R8428 VGND.n3011 VGND.n3010 599.125
R8429 VGND.n194 VGND.n193 599.125
R8430 VGND.n66 VGND.n65 599.125
R8431 VGND.n117 VGND.n116 599.125
R8432 VGND.n134 VGND.n133 599.125
R8433 VGND.n165 VGND.n164 599.125
R8434 VGND.n2210 VGND.n2182 599.125
R8435 VGND.n2972 VGND.n2971 599.125
R8436 VGND VGND.t206 581.61
R8437 VGND.t1072 VGND 573.181
R8438 VGND VGND.t2112 573.181
R8439 VGND.t2461 VGND 573.181
R8440 VGND.t50 VGND 573.181
R8441 VGND.n3013 VGND 564.751
R8442 VGND.t941 VGND 564.751
R8443 VGND.n3014 VGND 564.751
R8444 VGND.n3012 VGND 556.322
R8445 VGND.t945 VGND 539.465
R8446 VGND VGND.t124 539.465
R8447 VGND.t984 VGND.n806 494.779
R8448 VGND.n1166 VGND.t1758 492.058
R8449 VGND.t1597 VGND.n1175 492.058
R8450 VGND.n1176 VGND.t1621 492.058
R8451 VGND.t1760 VGND.n1188 492.058
R8452 VGND.n1189 VGND.t1772 492.058
R8453 VGND.t1794 VGND.n1207 492.058
R8454 VGND.n1208 VGND.t1693 492.058
R8455 VGND.t1713 VGND.n1220 492.058
R8456 VGND.n1247 VGND.t1799 492.058
R8457 VGND.n1246 VGND.t1638 492.058
R8458 VGND.n1240 VGND.t1649 492.058
R8459 VGND.n1239 VGND.t1738 492.058
R8460 VGND.n1233 VGND.t1809 492.058
R8461 VGND.t1660 VGND.n1277 492.058
R8462 VGND.n1278 VGND.t1727 492.058
R8463 VGND.t835 VGND.t845 481.877
R8464 VGND.t918 VGND.t835 481.877
R8465 VGND.t1540 VGND.t1102 481.877
R8466 VGND.t1102 VGND.t657 481.877
R8467 VGND.t1112 VGND 452.382
R8468 VGND.n1166 VGND.t1162 424.312
R8469 VGND.n1175 VGND.t560 424.312
R8470 VGND.n1176 VGND.t997 424.312
R8471 VGND.n1188 VGND.t697 424.312
R8472 VGND.n1189 VGND.t194 424.312
R8473 VGND.n1207 VGND.t2669 424.312
R8474 VGND.n1208 VGND.t2393 424.312
R8475 VGND.n1220 VGND.t779 424.312
R8476 VGND.n1247 VGND.t1393 424.312
R8477 VGND.t2521 VGND.n1246 424.312
R8478 VGND.n1240 VGND.t1413 424.312
R8479 VGND.t832 VGND.n1239 424.312
R8480 VGND.n1233 VGND.t195 424.312
R8481 VGND.n1277 VGND.t630 424.312
R8482 VGND.n1278 VGND.t1159 424.312
R8483 VGND.t1200 VGND.n222 424.312
R8484 VGND.t36 VGND 419.68
R8485 VGND.n2284 VGND.n503 413.043
R8486 VGND.t1915 VGND.t2130 408.469
R8487 VGND.t316 VGND.t2056 408.469
R8488 VGND.t292 VGND.t1081 408.469
R8489 VGND.t2642 VGND.t1829 408.469
R8490 VGND.t472 VGND.t2491 408.469
R8491 VGND.t273 VGND.t2564 408.469
R8492 VGND.t2638 VGND.t2361 408.469
R8493 VGND.t2438 VGND.t552 408.469
R8494 VGND.t426 VGND.t816 408.469
R8495 VGND.t243 VGND.t1534 408.469
R8496 VGND.t932 VGND.t2600 408.469
R8497 VGND.t804 VGND.t959 408.469
R8498 VGND.t1446 VGND.t396 408.469
R8499 VGND.t91 VGND.t366 408.469
R8500 VGND.t2170 VGND.t1471 408.469
R8501 VGND.t343 VGND.t2337 408.469
R8502 VGND.t1990 VGND.t2299 408.469
R8503 VGND.t2519 VGND.t150 408.469
R8504 VGND.t1307 VGND.t2154 408.469
R8505 VGND.t1856 VGND.t2446 408.469
R8506 VGND.t235 VGND.t318 408.469
R8507 VGND.t1244 VGND.t510 408.469
R8508 VGND.t1175 VGND.t2442 408.469
R8509 VGND.t577 VGND.t474 408.469
R8510 VGND.t719 VGND.t275 408.469
R8511 VGND.t713 VGND.t2640 408.469
R8512 VGND.t65 VGND.t2412 408.469
R8513 VGND.t1208 VGND.t261 408.469
R8514 VGND.t1463 VGND.t2632 408.469
R8515 VGND.t546 VGND.t2604 408.469
R8516 VGND.t2034 VGND.t2339 408.469
R8517 VGND.t1524 VGND.t398 408.469
R8518 VGND.t814 VGND.t1894 408.469
R8519 VGND.t2043 VGND.t2622 408.469
R8520 VGND.t180 VGND.t1048 408.469
R8521 VGND.t1869 VGND.t140 408.469
R8522 VGND.t388 VGND.t2498 408.469
R8523 VGND.t2570 VGND.t332 408.469
R8524 VGND.t2166 VGND.t1364 408.469
R8525 VGND.t558 VGND.t2329 408.469
R8526 VGND.t486 VGND.t767 408.469
R8527 VGND.t218 VGND.t304 408.469
R8528 VGND.t2134 VGND.t1127 408.469
R8529 VGND.t1026 VGND.t480 408.469
R8530 VGND.t296 VGND.t1154 408.469
R8531 VGND.t516 VGND.t97 408.469
R8532 VGND.t2420 VGND.t673 408.469
R8533 VGND.t350 VGND.t456 408.469
R8534 VGND.t1939 VGND.t269 408.469
R8535 VGND.t2430 VGND.t745 408.469
R8536 VGND.t2247 VGND.t828 408.469
R8537 VGND.t788 VGND.t1839 408.469
R8538 VGND.t2288 VGND.t2624 408.469
R8539 VGND.t164 VGND.t1421 408.469
R8540 VGND.t1387 VGND.t2331 408.469
R8541 VGND.t390 VGND.t418 408.469
R8542 VGND.t2542 VGND.t334 408.469
R8543 VGND.t2168 VGND.t759 408.469
R8544 VGND.t592 VGND.t2303 408.469
R8545 VGND.t326 VGND.t683 408.469
R8546 VGND.t432 VGND.t2162 408.469
R8547 VGND.t1262 VGND.t2138 408.469
R8548 VGND.t458 VGND.t622 408.469
R8549 VGND.t32 VGND.t300 408.469
R8550 VGND.t504 VGND.t2014 408.469
R8551 VGND.t466 VGND.t1017 408.469
R8552 VGND.t2075 VGND.t285 408.469
R8553 VGND.t247 VGND.t1861 408.469
R8554 VGND.t228 VGND.t2432 408.469
R8555 VGND.t810 VGND.t1122 408.469
R8556 VGND.t2259 VGND.t392 408.469
R8557 VGND.t2626 VGND.t5 408.469
R8558 VGND.t239 VGND.t168 408.469
R8559 VGND.t2333 VGND.t404 408.469
R8560 VGND.t60 VGND.t364 408.469
R8561 VGND.t156 VGND.t2677 408.469
R8562 VGND.t1043 VGND.t2325 408.469
R8563 VGND.t2305 VGND.t540 408.469
R8564 VGND.t302 VGND.t1520 408.469
R8565 VGND.t442 VGND.t2164 408.469
R8566 VGND.t2452 VGND.t1921 408.469
R8567 VGND.t308 VGND.t2054 408.469
R8568 VGND.t1079 VGND.t520 408.469
R8569 VGND.t1832 VGND.t2630 408.469
R8570 VGND.t2489 VGND.t462 408.469
R8571 VGND.t2562 VGND.t253 408.469
R8572 VGND.t2359 VGND.t2618 408.469
R8573 VGND.t550 VGND.t2426 408.469
R8574 VGND.t424 VGND.t798 408.469
R8575 VGND.t1532 VGND.t384 408.469
R8576 VGND.t929 VGND.t172 408.469
R8577 VGND.t957 VGND.t792 408.469
R8578 VGND.t1443 VGND.t380 408.469
R8579 VGND.t89 VGND.t358 408.469
R8580 VGND.t2158 VGND.t1515 408.469
R8581 VGND.t341 VGND.t2321 408.469
R8582 VGND.t492 VGND.t1891 408.469
R8583 VGND.t138 VGND.t2045 408.469
R8584 VGND.t2142 VGND.t1050 408.469
R8585 VGND.t2436 VGND.t1867 408.469
R8586 VGND.t310 VGND.t2500 408.469
R8587 VGND.t496 VGND.t2559 408.469
R8588 VGND.t2428 VGND.t1366 408.469
R8589 VGND.t464 VGND.t0 408.469
R8590 VGND.t257 VGND.t769 408.469
R8591 VGND.t2620 VGND.t220 408.469
R8592 VGND.t822 VGND.t1129 408.469
R8593 VGND.t249 VGND.t1028 408.469
R8594 VGND.t1156 VGND.t2616 408.469
R8595 VGND.t99 VGND.t174 408.469
R8596 VGND.t2323 VGND.t675 408.469
R8597 VGND.t352 VGND.t382 408.469
R8598 VGND.t1933 VGND.t796 408.469
R8599 VGND.t2610 VGND.t747 408.469
R8600 VGND.t170 VGND.t2249 408.469
R8601 VGND.t2160 VGND.t1837 408.469
R8602 VGND.t2290 VGND.t372 408.469
R8603 VGND.t322 VGND.t1423 408.469
R8604 VGND.t1389 VGND.t2150 408.469
R8605 VGND.t2315 VGND.t420 408.469
R8606 VGND.t2544 VGND.t478 408.469
R8607 VGND.t290 VGND.t761 408.469
R8608 VGND.t594 VGND.t2126 408.469
R8609 VGND.t468 VGND.t685 408.469
R8610 VGND.t434 VGND.t522 408.469
R8611 VGND.t508 VGND.t1264 408.469
R8612 VGND.t830 VGND.t624 408.469
R8613 VGND.t34 VGND.t287 408.469
R8614 VGND.t251 VGND.t1945 408.469
R8615 VGND.t2422 VGND.t740 408.469
R8616 VGND.t1166 VGND.t820 408.469
R8617 VGND.t2327 VGND.t1843 408.469
R8618 VGND.t2612 VGND.t214 408.469
R8619 VGND.t152 VGND.t703 408.469
R8620 VGND.t2317 VGND.t1385 408.469
R8621 VGND.t374 VGND.t414 408.469
R8622 VGND.t324 VGND.t2538 408.469
R8623 VGND.t2152 VGND.t568 408.469
R8624 VGND.t2293 VGND.t590 408.469
R8625 VGND.t314 VGND.t1141 408.469
R8626 VGND.t430 VGND.t2144 408.469
R8627 VGND.t637 VGND.t2128 408.469
R8628 VGND.t448 VGND.t618 408.469
R8629 VGND.t30 VGND.t524 408.469
R8630 VGND.t2646 VGND.t1876 408.469
R8631 VGND.t460 VGND.t1015 408.469
R8632 VGND.t283 VGND.t2073 408.469
R8633 VGND.t386 VGND.t1863 408.469
R8634 VGND.t2424 VGND.t226 408.469
R8635 VGND.t794 VGND.t1120 408.469
R8636 VGND.t376 VGND.t2257 408.469
R8637 VGND.t2614 VGND.t3 408.469
R8638 VGND.t154 VGND.t237 408.469
R8639 VGND.t2319 VGND.t402 408.469
R8640 VGND.t356 VGND.t1133 408.469
R8641 VGND.t146 VGND.t2675 408.469
R8642 VGND.t1041 VGND.t2313 408.469
R8643 VGND.t538 VGND.t2295 408.469
R8644 VGND.t526 VGND.t1518 408.469
R8645 VGND.t440 VGND.t2146 408.469
R8646 VGND.t1969 VGND.t2297 408.469
R8647 VGND.t1070 VGND.t144 408.469
R8648 VGND.t1097 VGND.t2148 408.469
R8649 VGND.t2444 VGND.t1847 408.469
R8650 VGND.t312 VGND.t208 408.469
R8651 VGND.t506 VGND.t572 408.469
R8652 VGND.t2434 VGND.t1182 408.469
R8653 VGND.t470 VGND.t407 408.469
R8654 VGND.t271 VGND.t772 408.469
R8655 VGND.t2634 VGND.t2484 408.469
R8656 VGND.t2410 VGND.t2023 408.469
R8657 VGND.t2124 VGND.t255 408.469
R8658 VGND.t2343 VGND.t2628 408.469
R8659 VGND.t2477 VGND.t182 408.469
R8660 VGND.t2027 VGND.t2335 408.469
R8661 VGND.t22 VGND.t394 408.469
R8662 VGND.t2644 VGND.t1897 408.469
R8663 VGND.t452 VGND.t2041 408.469
R8664 VGND.t279 VGND.t1046 408.469
R8665 VGND.t1871 VGND.t378 408.469
R8666 VGND.t2418 VGND.t2496 408.469
R8667 VGND.t2568 VGND.t790 408.469
R8668 VGND.t370 VGND.t1362 408.469
R8669 VGND.t556 VGND.t2608 408.469
R8670 VGND.t148 VGND.t765 408.469
R8671 VGND.t2311 VGND.t1538 408.469
R8672 VGND.t936 VGND.t336 408.469
R8673 VGND.t1024 VGND.t142 408.469
R8674 VGND.t2309 VGND.t1152 408.469
R8675 VGND.t488 VGND.t95 408.469
R8676 VGND.t518 VGND.t1475 408.469
R8677 VGND.t348 VGND.t2140 408.469
R8678 VGND.t1972 VGND.t454 408.469
R8679 VGND.t2450 VGND.t1068 408.469
R8680 VGND.t1095 VGND.t2440 408.469
R8681 VGND.t818 VGND.t1849 408.469
R8682 VGND.t2071 VGND.t498 408.469
R8683 VGND.t2602 VGND.t1553 408.469
R8684 VGND.t1180 VGND.t808 408.469
R8685 VGND.t263 VGND.t583 408.469
R8686 VGND.t2532 VGND.t368 408.469
R8687 VGND.t166 VGND.t2482 408.469
R8688 VGND.t2021 VGND.t784 408.469
R8689 VGND.t2122 VGND.t360 408.469
R8690 VGND.t2095 VGND.t158 408.469
R8691 VGND.t2475 VGND.t136 408.469
R8692 VGND.t482 VGND.t628 408.469
R8693 VGND.t2286 VGND.t328 408.469
R8694 VGND.t294 VGND.t1999 408.469
R8695 VGND.t2517 VGND.t490 408.469
R8696 VGND.t476 VGND.t1305 408.469
R8697 VGND.t277 VGND.t1859 408.469
R8698 VGND.t2454 VGND.t232 408.469
R8699 VGND.t2414 VGND.t1242 408.469
R8700 VGND.t265 VGND.t1173 408.469
R8701 VGND.t500 VGND.t575 408.469
R8702 VGND.t2606 VGND.t717 408.469
R8703 VGND.t711 VGND.t812 408.469
R8704 VGND.t62 VGND.t400 408.469
R8705 VGND.t178 VGND.t1206 408.469
R8706 VGND.t800 VGND.t1460 408.469
R8707 VGND.t544 VGND.t786 408.469
R8708 VGND.t2031 VGND.t330 408.469
R8709 VGND.t446 VGND.t160 408.469
R8710 VGND.t2156 VGND.t1942 408.469
R8711 VGND.t354 VGND.t742 408.469
R8712 VGND.t320 VGND.t1168 408.469
R8713 VGND.t1841 VGND.t512 408.469
R8714 VGND.t216 VGND.t494 408.469
R8715 VGND.t705 VGND.t450 408.469
R8716 VGND.t1383 VGND.t502 408.469
R8717 VGND.t412 VGND.t2456 408.469
R8718 VGND.t2536 VGND.t2416 408.469
R8719 VGND.t267 VGND.t566 408.469
R8720 VGND.t2636 VGND.t588 408.469
R8721 VGND.t826 VGND.t1139 408.469
R8722 VGND.t259 VGND.t2347 408.469
R8723 VGND.t635 VGND.t241 408.469
R8724 VGND.t162 VGND.t620 408.469
R8725 VGND.t28 VGND.t802 408.469
R8726 VGND.t1788 VGND.t245 408.469
R8727 VGND.t824 VGND.t1627 408.469
R8728 VGND.t806 VGND.t1709 408.469
R8729 VGND.t2307 VGND.t1731 408.469
R8730 VGND.t176 VGND.t1632 408.469
R8731 VGND.t2172 VGND.t1643 408.469
R8732 VGND.t2301 VGND.t1662 408.469
R8733 VGND.t362 VGND.t1803 408.469
R8734 VGND.t306 VGND.t1824 408.469
R8735 VGND.t2136 VGND.t1666 408.469
R8736 VGND.t484 VGND.t1743 408.469
R8737 VGND.t298 VGND.t1756 408.469
R8738 VGND.t2132 VGND.t1608 408.469
R8739 VGND.t2448 VGND.t1683 408.469
R8740 VGND.t281 VGND.t1774 408.469
R8741 VGND.t1599 VGND.t514 408.469
R8742 VGND.t916 VGND.t837 397.848
R8743 VGND.t837 VGND.t847 397.848
R8744 VGND.t847 VGND.t855 397.848
R8745 VGND.t855 VGND.t2114 397.848
R8746 VGND.t2114 VGND.t2115 397.848
R8747 VGND.t2115 VGND.t2118 397.848
R8748 VGND.t2118 VGND.t2119 397.848
R8749 VGND.t727 VGND.t1062 396.17
R8750 VGND.t1267 VGND.t1002 396.17
R8751 VGND.n2935 VGND.n2934 394.137
R8752 VGND.n2933 VGND.n208 394.137
R8753 VGND.n2932 VGND.n209 394.137
R8754 VGND.n2931 VGND.n210 394.137
R8755 VGND.n2930 VGND.n211 394.137
R8756 VGND.n2929 VGND.n212 394.137
R8757 VGND.n2928 VGND.n213 394.137
R8758 VGND.n2927 VGND.n214 394.137
R8759 VGND.n2926 VGND.n215 394.137
R8760 VGND.n2925 VGND.n216 394.137
R8761 VGND.n2924 VGND.n217 394.137
R8762 VGND.n2923 VGND.n218 394.137
R8763 VGND.n2922 VGND.n219 394.137
R8764 VGND.n2921 VGND.n220 394.137
R8765 VGND.n2920 VGND.n221 394.137
R8766 VGND.n2919 VGND.n2918 394.137
R8767 VGND.n2285 VGND.t130 387.421
R8768 VGND.n2284 VGND.t14 387.421
R8769 VGND.n2250 VGND.t39 387.421
R8770 VGND.n2248 VGND.t41 387.421
R8771 VGND.n1386 VGND.t16 387.421
R8772 VGND.t1003 VGND.t2552 362.452
R8773 VGND.t2552 VGND.t945 345.594
R8774 VGND VGND.t122 328.616
R8775 VGND VGND.t126 328.616
R8776 VGND VGND.t132 328.616
R8777 VGND VGND.t9 328.616
R8778 VGND VGND.t20 328.616
R8779 VGND.t1590 VGND.t1752 313.776
R8780 VGND.t1595 VGND.t1670 313.776
R8781 VGND.t1685 VGND.t1677 313.776
R8782 VGND.t1699 VGND.t1777 313.776
R8783 VGND.t1602 VGND.t1764 313.776
R8784 VGND.t1617 VGND.t1697 313.776
R8785 VGND.t1762 VGND.t1630 313.776
R8786 VGND.t1770 VGND.t1787 313.776
R8787 VGND.t1629 VGND.t1792 313.776
R8788 VGND.t1615 VGND.t1696 313.776
R8789 VGND.t1790 VGND.t1711 313.776
R8790 VGND.t1720 VGND.t1802 313.776
R8791 VGND.t1642 VGND.t1634 313.776
R8792 VGND.t1646 VGND.t1719 313.776
R8793 VGND.t1740 VGND.t1668 313.776
R8794 VGND.t1805 VGND.t1645 313.776
R8795 VGND.t736 VGND.t727 311.877
R8796 VGND.t206 VGND.t1267 311.877
R8797 VGND VGND.t732 303.449
R8798 VGND VGND.t736 295.019
R8799 VGND.n101 VGND.t846 287.832
R8800 VGND VGND.t1407 286.591
R8801 VGND.n93 VGND.t878 282.327
R8802 VGND.n2184 VGND.t2277 282.327
R8803 VGND.n104 VGND.t915 281.13
R8804 VGND.n2189 VGND.t2594 281.13
R8805 VGND.n177 VGND.t862 280.978
R8806 VGND.n177 VGND.t901 280.978
R8807 VGND.n78 VGND.t911 280.978
R8808 VGND.n78 VGND.t927 280.978
R8809 VGND.n146 VGND.t887 280.978
R8810 VGND.n146 VGND.t923 280.978
R8811 VGND.n482 VGND.t987 280.978
R8812 VGND.n482 VGND.t2274 280.978
R8813 VGND.n2263 VGND.t2595 280.978
R8814 VGND.n2263 VGND.t1101 280.978
R8815 VGND.n518 VGND.t2282 280.978
R8816 VGND.n518 VGND.t2271 280.978
R8817 VGND.n2194 VGND.t658 280.978
R8818 VGND.t1215 VGND 278.161
R8819 VGND.n2970 VGND 271.014
R8820 VGND.n3021 VGND.n4 259.389
R8821 VGND.n2347 VGND.n4 259.389
R8822 VGND.n3022 VGND.n3 252.988
R8823 VGND VGND.t857 252.875
R8824 VGND VGND.t734 252.875
R8825 VGND VGND.t729 252.875
R8826 VGND VGND.t853 252.875
R8827 VGND.t903 VGND 252.875
R8828 VGND.n887 VGND.t246 241.393
R8829 VGND.n330 VGND.t1931 241.393
R8830 VGND.n396 VGND.t2131 241.393
R8831 VGND.n400 VGND.t2300 241.393
R8832 VGND.n469 VGND.t815 241.393
R8833 VGND.n466 VGND.t270 241.393
R8834 VGND.n625 VGND.t505 241.393
R8835 VGND.n590 VGND.t2453 241.393
R8836 VGND.n587 VGND.t493 241.393
R8837 VGND.n547 VGND.t797 241.393
R8838 VGND.n628 VGND.t252 241.393
R8839 VGND.n632 VGND.t2647 241.393
R8840 VGND.n879 VGND.t2298 241.393
R8841 VGND.n800 VGND.t2645 241.393
R8842 VGND.n797 VGND.t455 241.393
R8843 VGND.n882 VGND.t295 241.393
R8844 VGND.n1024 VGND.t2157 241.393
R8845 VGND.n1014 VGND.t1937 241.393
R8846 VGND.n1333 VGND.t825 241.284
R8847 VGND.n894 VGND.t807 241.284
R8848 VGND.n932 VGND.t2308 241.284
R8849 VGND.n937 VGND.t177 241.284
R8850 VGND.n942 VGND.t2173 241.284
R8851 VGND.n947 VGND.t2302 241.284
R8852 VGND.n952 VGND.t363 241.284
R8853 VGND.n957 VGND.t307 241.284
R8854 VGND.n962 VGND.t2137 241.284
R8855 VGND.n967 VGND.t485 241.284
R8856 VGND.n972 VGND.t299 241.284
R8857 VGND.n977 VGND.t2133 241.284
R8858 VGND.n982 VGND.t2449 241.284
R8859 VGND.n987 VGND.t282 241.284
R8860 VGND.n1280 VGND.t1976 241.284
R8861 VGND.n1275 VGND.t1928 241.284
R8862 VGND.n1232 VGND.t2012 241.284
R8863 VGND.n1237 VGND.t2006 241.284
R8864 VGND.n1225 VGND.t1964 241.284
R8865 VGND.n1244 VGND.t1919 241.284
R8866 VGND.n1001 VGND.t2003 241.284
R8867 VGND.n1218 VGND.t1961 241.284
R8868 VGND.n1210 VGND.t1952 241.284
R8869 VGND.n1205 VGND.t1910 241.284
R8870 VGND.n1009 VGND.t1988 241.284
R8871 VGND.n1186 VGND.t1982 241.284
R8872 VGND.n1178 VGND.t1907 241.284
R8873 VGND.n1173 VGND.t1889 241.284
R8874 VGND.n1168 VGND.t1883 241.284
R8875 VGND.n2773 VGND.t1967 241.284
R8876 VGND.n294 VGND.t1925 241.284
R8877 VGND.n2730 VGND.t2009 241.284
R8878 VGND.n2735 VGND.t1997 241.284
R8879 VGND.n312 VGND.t1958 241.284
R8880 VGND.n2726 VGND.t1913 241.284
R8881 VGND.n326 VGND.t1994 241.284
R8882 VGND.n387 VGND.t1955 241.284
R8883 VGND.n384 VGND.t1949 241.284
R8884 VGND.n379 VGND.t1904 241.284
R8885 VGND.n373 VGND.t1985 241.284
R8886 VGND.n368 VGND.t1979 241.284
R8887 VGND.n362 VGND.t1901 241.284
R8888 VGND.n355 VGND.t1886 241.284
R8889 VGND.n2699 VGND.t1880 241.284
R8890 VGND.n2639 VGND.t317 241.284
R8891 VGND.n2644 VGND.t293 241.284
R8892 VGND.n2649 VGND.t2643 241.284
R8893 VGND.n2654 VGND.t473 241.284
R8894 VGND.n2659 VGND.t274 241.284
R8895 VGND.n2664 VGND.t2639 241.284
R8896 VGND.n2669 VGND.t2439 241.284
R8897 VGND.n394 VGND.t817 241.284
R8898 VGND.n2715 VGND.t244 241.284
R8899 VGND.n320 VGND.t2601 241.284
R8900 VGND.n2748 VGND.t805 241.284
R8901 VGND.n304 VGND.t397 241.284
R8902 VGND.n2753 VGND.t367 241.284
R8903 VGND.n2788 VGND.t2171 241.284
R8904 VGND.n287 VGND.t2338 241.284
R8905 VGND.n2343 VGND.t151 241.284
R8906 VGND.n2338 VGND.t2155 241.284
R8907 VGND.n2333 VGND.t2447 241.284
R8908 VGND.n2328 VGND.t319 241.284
R8909 VGND.n2323 VGND.t511 241.284
R8910 VGND.n2318 VGND.t2443 241.284
R8911 VGND.n2313 VGND.t475 241.284
R8912 VGND.n2308 VGND.t276 241.284
R8913 VGND.n2303 VGND.t2641 241.284
R8914 VGND.n2298 VGND.t2413 241.284
R8915 VGND.n2293 VGND.t262 241.284
R8916 VGND.n2288 VGND.t2633 241.284
R8917 VGND.n415 VGND.t2605 241.284
R8918 VGND.n2541 VGND.t2340 241.284
R8919 VGND.n2536 VGND.t399 241.284
R8920 VGND.n472 VGND.t2623 241.284
R8921 VGND.n2377 VGND.t181 241.284
R8922 VGND.n460 VGND.t141 241.284
R8923 VGND.n2403 VGND.t389 241.284
R8924 VGND.n452 VGND.t333 241.284
R8925 VGND.n2429 VGND.t2167 241.284
R8926 VGND.n444 VGND.t2330 241.284
R8927 VGND.n2455 VGND.t487 241.284
R8928 VGND.n436 VGND.t305 241.284
R8929 VGND.n2481 VGND.t2135 241.284
R8930 VGND.n428 VGND.t481 241.284
R8931 VGND.n2512 VGND.t297 241.284
R8932 VGND.n2517 VGND.t517 241.284
R8933 VGND.n2522 VGND.t2421 241.284
R8934 VGND.n2527 VGND.t457 241.284
R8935 VGND.n2364 VGND.t2431 241.284
R8936 VGND.n464 VGND.t829 241.284
R8937 VGND.n2390 VGND.t789 241.284
R8938 VGND.n456 VGND.t2625 241.284
R8939 VGND.n2416 VGND.t165 241.284
R8940 VGND.n448 VGND.t2332 241.284
R8941 VGND.n2442 VGND.t391 241.284
R8942 VGND.n440 VGND.t335 241.284
R8943 VGND.n2468 VGND.t2169 241.284
R8944 VGND.n432 VGND.t2304 241.284
R8945 VGND.n2494 VGND.t327 241.284
R8946 VGND.n424 VGND.t2163 241.284
R8947 VGND.n2499 VGND.t2139 241.284
R8948 VGND.n2810 VGND.t459 241.284
R8949 VGND.n2815 VGND.t301 241.284
R8950 VGND.n1911 VGND.t467 241.284
R8951 VGND.n623 VGND.t286 241.284
R8952 VGND.n1922 VGND.t248 241.284
R8953 VGND.n620 VGND.t2433 241.284
R8954 VGND.n1933 VGND.t811 241.284
R8955 VGND.n617 VGND.t393 241.284
R8956 VGND.n1944 VGND.t2627 241.284
R8957 VGND.n614 VGND.t169 241.284
R8958 VGND.n1955 VGND.t2334 241.284
R8959 VGND.n611 VGND.t365 241.284
R8960 VGND.n1966 VGND.t157 241.284
R8961 VGND.n608 VGND.t2326 241.284
R8962 VGND.n1977 VGND.t2306 241.284
R8963 VGND.n1982 VGND.t303 241.284
R8964 VGND.n1987 VGND.t2165 241.284
R8965 VGND.n597 VGND.t309 241.284
R8966 VGND.n594 VGND.t521 241.284
R8967 VGND.n2056 VGND.t2631 241.284
R8968 VGND.n2051 VGND.t463 241.284
R8969 VGND.n2046 VGND.t254 241.284
R8970 VGND.n2041 VGND.t2619 241.284
R8971 VGND.n2036 VGND.t2427 241.284
R8972 VGND.n2031 VGND.t799 241.284
R8973 VGND.n2026 VGND.t385 241.284
R8974 VGND.n2021 VGND.t173 241.284
R8975 VGND.n2016 VGND.t793 241.284
R8976 VGND.n2011 VGND.t381 241.284
R8977 VGND.n2006 VGND.t359 241.284
R8978 VGND.n2001 VGND.t2159 241.284
R8979 VGND.n1994 VGND.t2322 241.284
R8980 VGND.n2070 VGND.t139 241.284
R8981 VGND.n2075 VGND.t2143 241.284
R8982 VGND.n2080 VGND.t2437 241.284
R8983 VGND.n2085 VGND.t311 241.284
R8984 VGND.n2090 VGND.t497 241.284
R8985 VGND.n2095 VGND.t2429 241.284
R8986 VGND.n2100 VGND.t465 241.284
R8987 VGND.n2105 VGND.t258 241.284
R8988 VGND.n2110 VGND.t2621 241.284
R8989 VGND.n2115 VGND.t823 241.284
R8990 VGND.n2120 VGND.t250 241.284
R8991 VGND.n585 VGND.t2617 241.284
R8992 VGND.n2125 VGND.t175 241.284
R8993 VGND.n2835 VGND.t2324 241.284
R8994 VGND.n2840 VGND.t383 241.284
R8995 VGND.n2177 VGND.t2611 241.284
R8996 VGND.n1756 VGND.t171 241.284
R8997 VGND.n1762 VGND.t2161 241.284
R8998 VGND.n1753 VGND.t373 241.284
R8999 VGND.n1773 VGND.t323 241.284
R9000 VGND.n1750 VGND.t2151 241.284
R9001 VGND.n1784 VGND.t2316 241.284
R9002 VGND.n1747 VGND.t479 241.284
R9003 VGND.n1795 VGND.t291 241.284
R9004 VGND.n1744 VGND.t2127 241.284
R9005 VGND.n1806 VGND.t469 241.284
R9006 VGND.n1741 VGND.t523 241.284
R9007 VGND.n1817 VGND.t509 241.284
R9008 VGND.n1822 VGND.t831 241.284
R9009 VGND.n1827 VGND.t288 241.284
R9010 VGND.n1679 VGND.t2423 241.284
R9011 VGND.n1676 VGND.t821 241.284
R9012 VGND.n1690 VGND.t2328 241.284
R9013 VGND.n1695 VGND.t2613 241.284
R9014 VGND.n1700 VGND.t153 241.284
R9015 VGND.n1705 VGND.t2318 241.284
R9016 VGND.n1710 VGND.t375 241.284
R9017 VGND.n1715 VGND.t325 241.284
R9018 VGND.n1720 VGND.t2153 241.284
R9019 VGND.n1725 VGND.t2294 241.284
R9020 VGND.n1730 VGND.t315 241.284
R9021 VGND.n1673 VGND.t2145 241.284
R9022 VGND.n1846 VGND.t2129 241.284
R9023 VGND.n1841 VGND.t449 241.284
R9024 VGND.n1834 VGND.t525 241.284
R9025 VGND.n670 VGND.t461 241.284
R9026 VGND.n675 VGND.t284 241.284
R9027 VGND.n680 VGND.t387 241.284
R9028 VGND.n685 VGND.t2425 241.284
R9029 VGND.n690 VGND.t795 241.284
R9030 VGND.n695 VGND.t377 241.284
R9031 VGND.n700 VGND.t2615 241.284
R9032 VGND.n705 VGND.t155 241.284
R9033 VGND.n710 VGND.t2320 241.284
R9034 VGND.n715 VGND.t357 241.284
R9035 VGND.n720 VGND.t147 241.284
R9036 VGND.n667 VGND.t2314 241.284
R9037 VGND.n725 VGND.t2296 241.284
R9038 VGND.n2860 VGND.t527 241.284
R9039 VGND.n2865 VGND.t2147 241.284
R9040 VGND.n1353 VGND.t145 241.284
R9041 VGND.n875 VGND.t2149 241.284
R9042 VGND.n870 VGND.t2445 241.284
R9043 VGND.n810 VGND.t313 241.284
R9044 VGND.n824 VGND.t507 241.284
R9045 VGND.n829 VGND.t2435 241.284
R9046 VGND.n834 VGND.t471 241.284
R9047 VGND.n839 VGND.t272 241.284
R9048 VGND.n844 VGND.t2635 241.284
R9049 VGND.n849 VGND.t2411 241.284
R9050 VGND.n820 VGND.t256 241.284
R9051 VGND.n854 VGND.t2629 241.284
R9052 VGND.n735 VGND.t183 241.284
R9053 VGND.n1662 VGND.t2336 241.284
R9054 VGND.n1657 VGND.t395 241.284
R9055 VGND.n1391 VGND.t453 241.284
R9056 VGND.n1396 VGND.t280 241.284
R9057 VGND.n805 VGND.t379 241.284
R9058 VGND.n1491 VGND.t2419 241.284
R9059 VGND.n777 VGND.t791 241.284
R9060 VGND.n1517 VGND.t371 241.284
R9061 VGND.n769 VGND.t2609 241.284
R9062 VGND.n1543 VGND.t149 241.284
R9063 VGND.n1548 VGND.t2312 241.284
R9064 VGND.n761 VGND.t337 241.284
R9065 VGND.n1553 VGND.t143 241.284
R9066 VGND.n1633 VGND.t2310 241.284
R9067 VGND.n1638 VGND.t489 241.284
R9068 VGND.n1643 VGND.t519 241.284
R9069 VGND.n1648 VGND.t2141 241.284
R9070 VGND.n1411 VGND.t2451 241.284
R9071 VGND.n795 VGND.t2441 241.284
R9072 VGND.n1478 VGND.t819 241.284
R9073 VGND.n781 VGND.t499 241.284
R9074 VGND.n1504 VGND.t2603 241.284
R9075 VGND.n773 VGND.t809 241.284
R9076 VGND.n1530 VGND.t264 241.284
R9077 VGND.n765 VGND.t369 241.284
R9078 VGND.n1567 VGND.t167 241.284
R9079 VGND.n756 VGND.t785 241.284
R9080 VGND.n1582 VGND.t361 241.284
R9081 VGND.n1577 VGND.t159 241.284
R9082 VGND.n1572 VGND.t137 241.284
R9083 VGND.n2885 VGND.t483 241.284
R9084 VGND.n2890 VGND.t329 241.284
R9085 VGND.n885 VGND.t491 241.284
R9086 VGND.n1424 VGND.t477 241.284
R9087 VGND.n1429 VGND.t278 241.284
R9088 VGND.n1434 VGND.t2455 241.284
R9089 VGND.n1439 VGND.t2415 241.284
R9090 VGND.n1444 VGND.t266 241.284
R9091 VGND.n1449 VGND.t501 241.284
R9092 VGND.n1454 VGND.t2607 241.284
R9093 VGND.n791 VGND.t813 241.284
R9094 VGND.n1459 VGND.t401 241.284
R9095 VGND.n1596 VGND.t179 241.284
R9096 VGND.n1601 VGND.t801 241.284
R9097 VGND.n750 VGND.t787 241.284
R9098 VGND.n1614 VGND.t331 241.284
R9099 VGND.n1609 VGND.t161 241.284
R9100 VGND.n1032 VGND.t355 241.284
R9101 VGND.n1037 VGND.t321 241.284
R9102 VGND.n1029 VGND.t513 241.284
R9103 VGND.n1095 VGND.t495 241.284
R9104 VGND.n1090 VGND.t451 241.284
R9105 VGND.n1085 VGND.t503 241.284
R9106 VGND.n1080 VGND.t2457 241.284
R9107 VGND.n1075 VGND.t2417 241.284
R9108 VGND.n1070 VGND.t268 241.284
R9109 VGND.n1043 VGND.t2637 241.284
R9110 VGND.n1053 VGND.t827 241.284
R9111 VGND.n1058 VGND.t260 241.284
R9112 VGND.n1049 VGND.t242 241.284
R9113 VGND.n2905 VGND.t163 241.284
R9114 VGND.n2910 VGND.t803 241.284
R9115 VGND.n928 VGND.t515 241.284
R9116 VGND.t2130 VGND.t536 222.15
R9117 VGND.t1313 VGND.t1555 222.15
R9118 VGND.t1270 VGND.t316 222.15
R9119 VGND.t561 VGND.t1164 222.15
R9120 VGND.t2387 VGND.t292 222.15
R9121 VGND.t196 VGND.t1845 222.15
R9122 VGND.t2385 VGND.t2642 222.15
R9123 VGND.t1368 VGND.t2488 222.15
R9124 VGND.t534 VGND.t472 222.15
R9125 VGND.t778 VGND.t701 222.15
R9126 VGND.t2106 VGND.t273 222.15
R9127 VGND.t187 VGND.t1178 222.15
R9128 VGND.t2104 VGND.t2638 222.15
R9129 VGND.t564 VGND.t410 222.15
R9130 VGND.t532 VGND.t2438 222.15
R9131 VGND.t1019 VGND.t775 222.15
R9132 VGND.t816 VGND.t530 222.15
R9133 VGND.t1032 VGND.t1440 222.15
R9134 VGND.t2108 VGND.t243 222.15
R9135 VGND.t2401 VGND.t2026 222.15
R9136 VGND.t2600 VGND.t2383 222.15
R9137 VGND.t1451 VGND.t205 222.15
R9138 VGND.t2381 VGND.t804 222.15
R9139 VGND.t105 VGND.t2346 222.15
R9140 VGND.t396 VGND.t2102 222.15
R9141 VGND.t633 VGND.t1000 222.15
R9142 VGND.t366 VGND.t2391 222.15
R9143 VGND.t2030 VGND.t1228 222.15
R9144 VGND.t2389 VGND.t2170 222.15
R9145 VGND.t1066 VGND.t340 222.15
R9146 VGND.t2337 VGND.t528 222.15
R9147 VGND.t1612 VGND.t2407 222.15
R9148 VGND.t2299 VGND.t1331 222.15
R9149 VGND.t2059 VGND.t600 222.15
R9150 VGND.t150 VGND.t607 222.15
R9151 VGND.t1045 VGND.t115 222.15
R9152 VGND.t2154 VGND.t1191 222.15
R9153 VGND.t1866 VGND.t1381 222.15
R9154 VGND.t2446 VGND.t2251 222.15
R9155 VGND.t231 VGND.t2522 222.15
R9156 VGND.t318 VGND.t1329 222.15
R9157 VGND.t2567 VGND.t1449 222.15
R9158 VGND.t510 VGND.t603 222.15
R9159 VGND.t1382 VGND.t2070 222.15
R9160 VGND.t2442 VGND.t601 222.15
R9161 VGND.t555 VGND.t2048 222.15
R9162 VGND.t474 VGND.t1327 222.15
R9163 VGND.t764 VGND.t1020 222.15
R9164 VGND.t275 VGND.t1325 222.15
R9165 VGND.t1537 VGND.t2342 222.15
R9166 VGND.t2640 VGND.t605 222.15
R9167 VGND.t1131 VGND.t783 222.15
R9168 VGND.t2412 VGND.t200 222.15
R9169 VGND.t1138 VGND.t1230 222.15
R9170 VGND.t261 VGND.t198 222.15
R9171 VGND.t1158 VGND.t2648 222.15
R9172 VGND.t2632 VGND.t1197 222.15
R9173 VGND.t94 VGND.t2649 222.15
R9174 VGND.t2604 VGND.t1195 222.15
R9175 VGND.t677 VGND.t2051 222.15
R9176 VGND.t2339 VGND.t1193 222.15
R9177 VGND.t445 VGND.t696 222.15
R9178 VGND.t398 VGND.t609 222.15
R9179 VGND.t1763 VGND.t780 222.15
R9180 VGND.t1053 VGND.t814 222.15
R9181 VGND.t1397 VGND.t739 222.15
R9182 VGND.t2622 VGND.t1359 222.15
R9183 VGND.t2245 VGND.t186 222.15
R9184 VGND.t1414 VGND.t180 222.15
R9185 VGND.t2380 VGND.t1835 222.15
R9186 VGND.t140 VGND.t1059 222.15
R9187 VGND.t2494 VGND.t45 222.15
R9188 VGND.t976 VGND.t388 222.15
R9189 VGND.t757 VGND.t707 222.15
R9190 VGND.t332 VGND.t1355 222.15
R9191 VGND.t1171 VGND.t948 222.15
R9192 VGND.t1353 VGND.t2166 222.15
R9193 VGND.t1187 VGND.t416 222.15
R9194 VGND.t2329 VGND.t974 222.15
R9195 VGND.t2540 VGND.t2524 222.15
R9196 VGND.t972 VGND.t486 222.15
R9197 VGND.t113 VGND.t570 222.15
R9198 VGND.t304 VGND.t1357 222.15
R9199 VGND.t597 VGND.t938 222.15
R9200 VGND.t1057 VGND.t2134 222.15
R9201 VGND.t1087 VGND.t1453 222.15
R9202 VGND.t480 VGND.t1055 222.15
R9203 VGND.t437 VGND.t1315 222.15
R9204 VGND.t1351 VGND.t296 222.15
R9205 VGND.t118 VGND.t639 222.15
R9206 VGND.t1418 VGND.t516 222.15
R9207 VGND.t2403 VGND.t1022 222.15
R9208 VGND.t1416 VGND.t2420 222.15
R9209 VGND.t2514 VGND.t346 222.15
R9210 VGND.t456 VGND.t970 222.15
R9211 VGND.t1591 VGND.t2550 222.15
R9212 VGND.t269 VGND.t2198 222.15
R9213 VGND.t1203 VGND.t949 222.15
R9214 VGND.t2225 VGND.t2430 222.15
R9215 VGND.t994 VGND.t2508 222.15
R9216 VGND.t828 VGND.t2554 222.15
R9217 VGND.t1852 VGND.t1199 222.15
R9218 VGND.t2204 VGND.t788 222.15
R9219 VGND.t1458 VGND.t212 222.15
R9220 VGND.t2624 VGND.t694 222.15
R9221 VGND.t1551 VGND.t1006 222.15
R9222 VGND.t2221 VGND.t164 222.15
R9223 VGND.t1324 VGND.t2255 222.15
R9224 VGND.t2331 VGND.t2219 222.15
R9225 VGND.t581 VGND.t679 222.15
R9226 VGND.t692 VGND.t390 222.15
R9227 VGND.t19 VGND.t2530 222.15
R9228 VGND.t334 VGND.t690 222.15
R9229 VGND.t1259 VGND.t1459 222.15
R9230 VGND.t2223 VGND.t2168 222.15
R9231 VGND.t950 VGND.t2019 222.15
R9232 VGND.t2303 VGND.t2202 222.15
R9233 VGND.t2673 VGND.t1189 222.15
R9234 VGND.t2200 VGND.t326 222.15
R9235 VGND.t1229 VGND.t2093 222.15
R9236 VGND.t2162 VGND.t2217 222.15
R9237 VGND.t2473 VGND.t81 222.15
R9238 VGND.t2138 VGND.t2215 222.15
R9239 VGND.t626 VGND.t1205 222.15
R9240 VGND.t2556 VGND.t458 222.15
R9241 VGND.t2398 VGND.t26 222.15
R9242 VGND.t300 VGND.t688 222.15
R9243 VGND.t1657 VGND.t955 222.15
R9244 VGND.t2196 VGND.t504 222.15
R9245 VGND.t120 VGND.t2053 222.15
R9246 VGND.t79 VGND.t466 222.15
R9247 VGND.t699 VGND.t1078 222.15
R9248 VGND.t285 VGND.t1337 222.15
R9249 VGND.t1828 VGND.t1008 222.15
R9250 VGND.t1118 VGND.t247 222.15
R9251 VGND.t1190 VGND.t587 222.15
R9252 VGND.t2432 VGND.t2194 222.15
R9253 VGND.t1126 VGND.t656 222.15
R9254 VGND.t75 VGND.t810 222.15
R9255 VGND.t617 VGND.t1185 222.15
R9256 VGND.t392 VGND.t73 222.15
R9257 VGND.t549 VGND.t134 222.15
R9258 VGND.t2192 VGND.t2626 222.15
R9259 VGND.t2357 VGND.t423 222.15
R9260 VGND.t168 VGND.t2190 222.15
R9261 VGND.t1531 VGND.t698 222.15
R9262 VGND.t77 VGND.t2333 222.15
R9263 VGND.t1084 VGND.t934 222.15
R9264 VGND.t364 VGND.t1116 222.15
R9265 VGND.t1136 VGND.t2534 222.15
R9266 VGND.t1114 VGND.t156 222.15
R9267 VGND.t2512 VGND.t1448 222.15
R9268 VGND.t2325 VGND.t71 222.15
R9269 VGND.t88 VGND.t2406 222.15
R9270 VGND.t69 VGND.t2305 222.15
R9271 VGND.t116 VGND.t1473 222.15
R9272 VGND.t1339 VGND.t302 222.15
R9273 VGND.t2061 VGND.t439 222.15
R9274 VGND.t2164 VGND.t2188 222.15
R9275 VGND.t1791 VGND.t2368 222.15
R9276 VGND.t2233 VGND.t2452 222.15
R9277 VGND.t2039 VGND.t1312 222.15
R9278 VGND.t2683 VGND.t308 222.15
R9279 VGND.t2551 VGND.t1163 222.15
R9280 VGND.t520 VGND.t2574 222.15
R9281 VGND.t1846 VGND.t185 222.15
R9282 VGND.t2630 VGND.t2572 222.15
R9283 VGND.t2292 VGND.t13 222.15
R9284 VGND.t462 VGND.t2231 222.15
R9285 VGND.t700 VGND.t1442 222.15
R9286 VGND.t253 VGND.t2584 222.15
R9287 VGND.t1177 VGND.t1301 222.15
R9288 VGND.t2618 VGND.t2582 222.15
R9289 VGND.t409 VGND.t2052 222.15
R9290 VGND.t2426 VGND.t2229 222.15
R9291 VGND.t774 VGND.t996 222.15
R9292 VGND.t798 VGND.t2227 222.15
R9293 VGND.t1031 VGND.t193 222.15
R9294 VGND.t384 VGND.t2586 222.15
R9295 VGND.t2025 VGND.t2589 222.15
R9296 VGND.t172 VGND.t2237 222.15
R9297 VGND.t1450 VGND.t1093 222.15
R9298 VGND.t792 VGND.t2235 222.15
R9299 VGND.t2345 VGND.t1470 222.15
R9300 VGND.t380 VGND.t2580 222.15
R9301 VGND.t2479 VGND.t1005 222.15
R9302 VGND.t358 VGND.t2578 222.15
R9303 VGND.t2029 VGND.t631 222.15
R9304 VGND.t2576 VGND.t2158 222.15
R9305 VGND.t2408 VGND.t339 222.15
R9306 VGND.t2321 VGND.t2685 222.15
R9307 VGND.t1614 VGND.t991 222.15
R9308 VGND.t648 VGND.t492 222.15
R9309 VGND.t777 VGND.t744 222.15
R9310 VGND.t1239 VGND.t138 222.15
R9311 VGND.t1085 VGND.t2246 222.15
R9312 VGND.t611 VGND.t2142 222.15
R9313 VGND.t680 VGND.t1834 222.15
R9314 VGND.t654 VGND.t2436 222.15
R9315 VGND.t2679 VGND.t2495 222.15
R9316 VGND.t646 VGND.t310 222.15
R9317 VGND.t2365 VGND.t1420 222.15
R9318 VGND.t1235 VGND.t496 222.15
R9319 VGND.t11 VGND.t1172 222.15
R9320 VGND.t1233 VGND.t2428 222.15
R9321 VGND.t672 VGND.t417 222.15
R9322 VGND.t644 VGND.t464 222.15
R9323 VGND.t2527 VGND.t2541 222.15
R9324 VGND.t642 VGND.t257 222.15
R9325 VGND.t112 VGND.t758 222.15
R9326 VGND.t1237 VGND.t2620 222.15
R9327 VGND.t58 VGND.t598 222.15
R9328 VGND.t652 VGND.t822 222.15
R9329 VGND.t2038 VGND.t1454 222.15
R9330 VGND.t650 VGND.t249 222.15
R9331 VGND.t1226 VGND.t1274 222.15
R9332 VGND.t2616 VGND.t1231 222.15
R9333 VGND.t1261 VGND.t1874 222.15
R9334 VGND.t174 VGND.t615 222.15
R9335 VGND.t1023 VGND.t1439 222.15
R9336 VGND.t613 VGND.t2323 222.15
R9337 VGND.t563 VGND.t347 222.15
R9338 VGND.t382 VGND.t640 222.15
R9339 VGND.t1588 VGND.t1302 222.15
R9340 VGND.t796 VGND.t751 222.15
R9341 VGND.t1204 VGND.t670 222.15
R9342 VGND.t202 VGND.t2610 222.15
R9343 VGND.t1109 VGND.t1094 222.15
R9344 VGND.t2087 VGND.t170 222.15
R9345 VGND.t1246 VGND.t1851 222.15
R9346 VGND.t2085 VGND.t2160 222.15
R9347 VGND.t954 VGND.t213 222.15
R9348 VGND.t372 VGND.t1224 222.15
R9349 VGND.t1552 VGND.t197 222.15
R9350 VGND.t2211 VGND.t322 222.15
R9351 VGND.t1217 VGND.t2256 222.15
R9352 VGND.t2150 VGND.t2209 222.15
R9353 VGND.t582 VGND.t2588 222.15
R9354 VGND.t1222 VGND.t2315 222.15
R9355 VGND.t189 VGND.t2531 222.15
R9356 VGND.t478 VGND.t1220 222.15
R9357 VGND.t1260 VGND.t2655 222.15
R9358 VGND.t2213 VGND.t290 222.15
R9359 VGND.t1530 VGND.t2020 222.15
R9360 VGND.t2126 VGND.t755 222.15
R9361 VGND.t2674 VGND.t1030 222.15
R9362 VGND.t753 VGND.t468 222.15
R9363 VGND.t2404 VGND.t2094 222.15
R9364 VGND.t522 VGND.t2207 222.15
R9365 VGND.t2474 VGND.t1188 222.15
R9366 VGND.t2091 VGND.t508 222.15
R9367 VGND.t104 VGND.t627 222.15
R9368 VGND.t2089 VGND.t830 222.15
R9369 VGND.t2101 VGND.t27 222.15
R9370 VGND.t287 VGND.t1218 222.15
R9371 VGND.t1655 VGND.t1107 222.15
R9372 VGND.t1149 VGND.t251 222.15
R9373 VGND.t2409 VGND.t1201 222.15
R9374 VGND.t2097 VGND.t2422 222.15
R9375 VGND.t121 VGND.t2507 222.15
R9376 VGND.t820 VGND.t83 222.15
R9377 VGND.t1854 VGND.t1334 222.15
R9378 VGND.t1037 VGND.t2327 222.15
R9379 VGND.t1065 VGND.t211 222.15
R9380 VGND.t1147 VGND.t2612 222.15
R9381 VGND.t2374 VGND.t1549 222.15
R9382 VGND.t1347 VGND.t152 222.15
R9383 VGND.t102 VGND.t2253 222.15
R9384 VGND.t1345 VGND.t2317 222.15
R9385 VGND.t2395 VGND.t580 222.15
R9386 VGND.t1145 VGND.t374 222.15
R9387 VGND.t2375 VGND.t225 222.15
R9388 VGND.t1143 VGND.t324 222.15
R9389 VGND.t2369 VGND.t1258 222.15
R9390 VGND.t1349 VGND.t2152 222.15
R9391 VGND.t2509 VGND.t2018 222.15
R9392 VGND.t1035 VGND.t2293 222.15
R9393 VGND.t106 VGND.t2672 222.15
R9394 VGND.t1033 VGND.t314 222.15
R9395 VGND.t2513 VGND.t1273 222.15
R9396 VGND.t2144 VGND.t1343 222.15
R9397 VGND.t2472 VGND.t944 222.15
R9398 VGND.t2128 VGND.t1341 222.15
R9399 VGND.t953 VGND.t1001 222.15
R9400 VGND.t85 VGND.t448 222.15
R9401 VGND.t110 VGND.t24 222.15
R9402 VGND.t524 VGND.t2099 222.15
R9403 VGND.t1664 VGND.t2372 222.15
R9404 VGND.t1435 VGND.t2646 222.15
R9405 VGND.t1266 VGND.t2352 222.15
R9406 VGND.t1425 VGND.t460 222.15
R9407 VGND.t114 VGND.t1077 222.15
R9408 VGND.t1513 VGND.t283 222.15
R9409 VGND.t1007 VGND.t1831 222.15
R9410 VGND.t1511 VGND.t386 222.15
R9411 VGND.t585 VGND.t586 222.15
R9412 VGND.t1433 VGND.t2424 222.15
R9413 VGND.t1526 VGND.t1125 222.15
R9414 VGND.t1503 VGND.t794 222.15
R9415 VGND.t599 VGND.t1184 222.15
R9416 VGND.t1501 VGND.t376 222.15
R9417 VGND.t2355 VGND.t548 222.15
R9418 VGND.t1431 VGND.t2614 222.15
R9419 VGND.t1061 VGND.t422 222.15
R9420 VGND.t1429 VGND.t154 222.15
R9421 VGND.t2396 VGND.t1039 222.15
R9422 VGND.t1505 VGND.t2319 222.15
R9423 VGND.t43 VGND.t931 222.15
R9424 VGND.t1509 VGND.t356 222.15
R9425 VGND.t1396 VGND.t1135 222.15
R9426 VGND.t1507 VGND.t146 222.15
R9427 VGND.t1522 VGND.t1445 222.15
R9428 VGND.t2313 VGND.t1499 222.15
R9429 VGND.t87 VGND.t2037 222.15
R9430 VGND.t2295 VGND.t1497 222.15
R9431 VGND.t1517 VGND.t103 222.15
R9432 VGND.t1495 VGND.t526 222.15
R9433 VGND.t1092 VGND.t438 222.15
R9434 VGND.t2146 VGND.t1427 222.15
R9435 VGND.t1796 VGND.t8 222.15
R9436 VGND.t2297 VGND.t1584 222.15
R9437 VGND.t2516 VGND.t1160 222.15
R9438 VGND.t144 VGND.t1562 222.15
R9439 VGND.t1304 VGND.t82 222.15
R9440 VGND.t2148 VGND.t1576 222.15
R9441 VGND.t1855 VGND.t1392 222.15
R9442 VGND.t1578 VGND.t2444 222.15
R9443 VGND.t1455 VGND.t2481 222.15
R9444 VGND.t1586 VGND.t312 222.15
R9445 VGND.t671 VGND.t1241 222.15
R9446 VGND.t1566 VGND.t506 222.15
R9447 VGND.t2356 VGND.t1361 222.15
R9448 VGND.t1568 VGND.t2434 222.15
R9449 VGND.t2174 VGND.t574 222.15
R9450 VGND.t1556 VGND.t470 222.15
R9451 VGND.t965 VGND.t716 222.15
R9452 VGND.t1558 VGND.t271 222.15
R9453 VGND.t2511 VGND.t710 222.15
R9454 VGND.t1564 VGND.t2634 222.15
R9455 VGND.t1210 VGND.t67 222.15
R9456 VGND.t1580 VGND.t2410 222.15
R9457 VGND.t2656 VGND.t962 222.15
R9458 VGND.t255 VGND.t1582 222.15
R9459 VGND.t429 VGND.t1161 222.15
R9460 VGND.t2628 VGND.t1570 222.15
R9461 VGND.t543 VGND.t963 222.15
R9462 VGND.t182 VGND.t1572 222.15
R9463 VGND.t2036 VGND.t1438 222.15
R9464 VGND.t2335 VGND.t1574 222.15
R9465 VGND.t2285 VGND.t1010 222.15
R9466 VGND.t394 VGND.t1560 222.15
R9467 VGND.t1705 VGND.t2353 222.15
R9468 VGND.t2663 VGND.t2644 222.15
R9469 VGND.t2349 VGND.t1314 222.15
R9470 VGND.t1283 VGND.t452 222.15
R9471 VGND.t2502 VGND.t1165 222.15
R9472 VGND.t2064 VGND.t279 222.15
R9473 VGND.t2394 VGND.t1836 222.15
R9474 VGND.t378 VGND.t2062 222.15
R9475 VGND.t2493 VGND.t44 222.15
R9476 VGND.t2661 VGND.t2418 222.15
R9477 VGND.t2650 VGND.t702 222.15
R9478 VGND.t790 VGND.t1279 222.15
R9479 VGND.t1179 VGND.t59 222.15
R9480 VGND.t1277 VGND.t370 222.15
R9481 VGND.t1395 VGND.t411 222.15
R9482 VGND.t2608 VGND.t2659 222.15
R9483 VGND.t776 VGND.t2523 222.15
R9484 VGND.t2657 VGND.t148 222.15
R9485 VGND.t2040 VGND.t565 222.15
R9486 VGND.t1281 VGND.t2311 222.15
R9487 VGND.t117 VGND.t596 222.15
R9488 VGND.t336 VGND.t2667 222.15
R9489 VGND.t1452 VGND.t1412 222.15
R9490 VGND.t142 VGND.t2665 222.15
R9491 VGND.t436 VGND.t2060 222.15
R9492 VGND.t1275 VGND.t2309 222.15
R9493 VGND.t1108 VGND.t634 222.15
R9494 VGND.t2068 VGND.t488 222.15
R9495 VGND.t993 VGND.t1021 222.15
R9496 VGND.t2066 VGND.t518 222.15
R9497 VGND.t1089 VGND.t345 222.15
R9498 VGND.t2140 VGND.t1285 222.15
R9499 VGND.t1594 VGND.t660 222.15
R9500 VGND.t454 VGND.t1316 222.15
R9501 VGND.t2515 VGND.t1394 222.15
R9502 VGND.t1371 VGND.t2450 222.15
R9503 VGND.t2366 VGND.t1303 222.15
R9504 VGND.t2440 VGND.t2176 222.15
R9505 VGND.t1858 VGND.t781 222.15
R9506 VGND.t1322 VGND.t818 222.15
R9507 VGND.t943 VGND.t2480 222.15
R9508 VGND.t498 VGND.t1379 222.15
R9509 VGND.t1124 VGND.t2351 222.15
R9510 VGND.t2186 VGND.t2602 222.15
R9511 VGND.t1528 VGND.t2363 222.15
R9512 VGND.t808 VGND.t2184 222.15
R9513 VGND.t7 VGND.t1099 222.15
R9514 VGND.t1377 VGND.t263 222.15
R9515 VGND.t2682 VGND.t715 222.15
R9516 VGND.t368 VGND.t1375 222.15
R9517 VGND.t406 VGND.t2358 222.15
R9518 VGND.t1369 VGND.t166 222.15
R9519 VGND.t1456 VGND.t64 222.15
R9520 VGND.t784 VGND.t1320 222.15
R9521 VGND.t961 VGND.t2402 222.15
R9522 VGND.t360 VGND.t1318 222.15
R9523 VGND.t1462 VGND.t669 222.15
R9524 VGND.t158 VGND.t2182 222.15
R9525 VGND.t542 VGND.t1333 222.15
R9526 VGND.t136 VGND.t2180 222.15
R9527 VGND.t2033 VGND.t782 222.15
R9528 VGND.t2178 VGND.t482 222.15
R9529 VGND.t2399 VGND.t2284 222.15
R9530 VGND.t328 VGND.t1373 222.15
R9531 VGND.t1708 VGND.t2400 222.15
R9532 VGND.t1487 VGND.t294 222.15
R9533 VGND.t2049 VGND.t2058 222.15
R9534 VGND.t490 VGND.t1291 222.15
R9535 VGND.t1083 VGND.t682 222.15
R9536 VGND.t1247 VGND.t476 222.15
R9537 VGND.t18 VGND.t1873 222.15
R9538 VGND.t1493 VGND.t277 222.15
R9539 VGND.t1009 VGND.t230 222.15
R9540 VGND.t1485 VGND.t2454 222.15
R9541 VGND.t204 VGND.t2566 222.15
R9542 VGND.t1287 VGND.t2414 222.15
R9543 VGND.t338 VGND.t1186 222.15
R9544 VGND.t1255 VGND.t265 222.15
R9545 VGND.t108 VGND.t554 222.15
R9546 VGND.t1297 VGND.t500 222.15
R9547 VGND.t1227 VGND.t763 222.15
R9548 VGND.t1295 VGND.t2606 222.15
R9549 VGND.t1457 VGND.t1536 222.15
R9550 VGND.t812 VGND.t1289 222.15
R9551 VGND.t935 VGND.t2535 222.15
R9552 VGND.t400 VGND.t1491 222.15
R9553 VGND.t1137 VGND.t668 222.15
R9554 VGND.t1489 VGND.t178 222.15
R9555 VGND.t1211 VGND.t1151 222.15
R9556 VGND.t1253 VGND.t800 222.15
R9557 VGND.t2525 VGND.t93 222.15
R9558 VGND.t786 VGND.t1251 222.15
R9559 VGND.t1474 VGND.t956 222.15
R9560 VGND.t330 VGND.t1249 222.15
R9561 VGND.t444 VGND.t2175 222.15
R9562 VGND.t160 VGND.t1293 222.15
R9563 VGND.t1776 VGND.t1336 222.15
R9564 VGND.t1483 VGND.t2156 222.15
R9565 VGND.t1437 VGND.t1202 222.15
R9566 VGND.t966 VGND.t354 222.15
R9567 VGND.t1090 VGND.t2506 222.15
R9568 VGND.t721 VGND.t320 222.15
R9569 VGND.t1309 VGND.t1853 222.15
R9570 VGND.t512 VGND.t2243 222.15
R9571 VGND.t210 VGND.t107 222.15
R9572 VGND.t494 VGND.t1481 222.15
R9573 VGND.t1550 VGND.t1212 222.15
R9574 VGND.t450 VGND.t2081 222.15
R9575 VGND.t2254 VGND.t2397 222.15
R9576 VGND.t502 VGND.t2079 222.15
R9577 VGND.t579 VGND.t1527 222.15
R9578 VGND.t2456 VGND.t1479 222.15
R9579 VGND.t224 VGND.t562 222.15
R9580 VGND.t2416 VGND.t1477 222.15
R9581 VGND.t1257 VGND.t119 222.15
R9582 VGND.t2083 VGND.t267 222.15
R9583 VGND.t188 VGND.t68 222.15
R9584 VGND.t2241 VGND.t2636 222.15
R9585 VGND.t184 VGND.t2671 222.15
R9586 VGND.t2239 VGND.t826 222.15
R9587 VGND.t632 VGND.t1272 222.15
R9588 VGND.t2077 VGND.t259 222.15
R9589 VGND.t12 VGND.t2471 222.15
R9590 VGND.t241 VGND.t725 222.15
R9591 VGND.t952 VGND.t2487 222.15
R9592 VGND.t723 VGND.t162 222.15
R9593 VGND.t2458 VGND.t25 222.15
R9594 VGND.t802 VGND.t968 222.15
R9595 VGND.t1665 VGND.t995 222.15
R9596 VGND.t245 VGND.t1625 222.15
R9597 VGND.t2047 VGND.t2373 222.15
R9598 VGND.t1706 VGND.t824 222.15
R9599 VGND.t2371 VGND.t1052 222.15
R9600 VGND.t1785 VGND.t806 222.15
R9601 VGND.t135 VGND.t1865 222.15
R9602 VGND.t1807 VGND.t2307 222.15
R9603 VGND.t992 VGND.t234 222.15
R9604 VGND.t1636 VGND.t176 222.15
R9605 VGND.t951 VGND.t2561 222.15
R9606 VGND.t1725 VGND.t2172 222.15
R9607 VGND.t2350 VGND.t1391 222.15
R9608 VGND.t1736 VGND.t2301 222.15
R9609 VGND.t2510 VGND.t2 222.15
R9610 VGND.t1640 VGND.t362 222.15
R9611 VGND.t1300 VGND.t771 222.15
R9612 VGND.t1658 VGND.t306 222.15
R9613 VGND.t2670 VGND.t222 222.15
R9614 VGND.t1723 VGND.t2136 222.15
R9615 VGND.t1398 VGND.t1132 222.15
R9616 VGND.t1820 VGND.t484 222.15
R9617 VGND.t2354 VGND.t687 222.15
R9618 VGND.t1592 VGND.t298 222.15
R9619 VGND.t2529 VGND.t1040 222.15
R9620 VGND.t1741 VGND.t2132 222.15
R9621 VGND.t1088 VGND.t101 222.15
R9622 VGND.t1754 VGND.t2448 222.15
R9623 VGND.t681 VGND.t678 222.15
R9624 VGND.t1779 VGND.t281 222.15
R9625 VGND.t109 VGND.t1523 222.15
R9626 VGND.t514 VGND.t1679 222.15
R9627 VGND.t1751 VGND.t1335 222.15
R9628 VGND.n2346 VGND.n3 218.73
R9629 VGND.n489 VGND.n487 214.365
R9630 VGND.n489 VGND.n488 214.365
R9631 VGND.n479 VGND.n477 214.365
R9632 VGND.n479 VGND.n478 214.365
R9633 VGND.n497 VGND.n495 214.365
R9634 VGND.n497 VGND.n496 214.365
R9635 VGND.n2270 VGND.n2268 214.365
R9636 VGND.n2270 VGND.n2269 214.365
R9637 VGND.n2260 VGND.n2258 214.365
R9638 VGND.n2260 VGND.n2259 214.365
R9639 VGND.n2278 VGND.n2276 214.365
R9640 VGND.n2278 VGND.n2277 214.365
R9641 VGND.n525 VGND.n523 214.365
R9642 VGND.n525 VGND.n524 214.365
R9643 VGND.n515 VGND.n513 214.365
R9644 VGND.n515 VGND.n514 214.365
R9645 VGND.n533 VGND.n531 214.365
R9646 VGND.n533 VGND.n532 214.365
R9647 VGND.n2191 VGND.n2190 214.365
R9648 VGND.n1140 VGND.n1139 213.613
R9649 VGND.n1142 VGND.n1141 213.613
R9650 VGND.n1112 VGND.n1110 213.613
R9651 VGND.n1112 VGND.n1111 213.613
R9652 VGND.n1115 VGND.n1113 213.613
R9653 VGND.n1115 VGND.n1114 213.613
R9654 VGND.n2236 VGND.n2229 213.613
R9655 VGND.n2236 VGND.n2230 213.613
R9656 VGND.n2234 VGND.n2231 213.613
R9657 VGND.n2234 VGND.n2233 213.613
R9658 VGND.n1374 VGND.n1367 213.613
R9659 VGND.n1374 VGND.n1368 213.613
R9660 VGND.n1372 VGND.n1369 213.613
R9661 VGND.n1372 VGND.n1371 213.613
R9662 VGND.n1154 VGND.t1399 211.359
R9663 VGND.n179 VGND.n175 207.965
R9664 VGND.n179 VGND.n176 207.965
R9665 VGND.n173 VGND.n171 207.965
R9666 VGND.n173 VGND.n172 207.965
R9667 VGND.n186 VGND.n169 207.965
R9668 VGND.n186 VGND.n170 207.965
R9669 VGND.n98 VGND.n97 207.965
R9670 VGND.n110 VGND.n95 207.965
R9671 VGND.n102 VGND.n100 207.965
R9672 VGND.n80 VGND.n76 207.965
R9673 VGND.n80 VGND.n77 207.965
R9674 VGND.n74 VGND.n72 207.965
R9675 VGND.n74 VGND.n73 207.965
R9676 VGND.n87 VGND.n70 207.965
R9677 VGND.n87 VGND.n71 207.965
R9678 VGND.n148 VGND.n144 207.965
R9679 VGND.n148 VGND.n145 207.965
R9680 VGND.n142 VGND.n140 207.965
R9681 VGND.n142 VGND.n141 207.965
R9682 VGND.n155 VGND.n138 207.965
R9683 VGND.n155 VGND.n139 207.965
R9684 VGND.n2188 VGND.n2187 207.965
R9685 VGND.n2205 VGND.n2185 207.965
R9686 VGND.n2981 VGND.n2979 207.213
R9687 VGND.n2981 VGND.n2980 207.213
R9688 VGND.n2985 VGND.n2976 207.213
R9689 VGND.n2985 VGND.n2977 207.213
R9690 VGND.n18 VGND.n16 207.213
R9691 VGND.n18 VGND.n17 207.213
R9692 VGND.n22 VGND.n14 207.213
R9693 VGND.n22 VGND.n15 207.213
R9694 VGND.n2951 VGND.n2950 207.213
R9695 VGND.n2955 VGND.n2949 207.213
R9696 VGND.n44 VGND.n42 207.213
R9697 VGND.n44 VGND.n43 207.213
R9698 VGND.n48 VGND.n40 207.213
R9699 VGND.n48 VGND.n41 207.213
R9700 VGND.n109 VGND.n96 207.213
R9701 VGND.n2204 VGND.n2186 207.213
R9702 VGND.t1936 VGND.t1681 203.242
R9703 VGND.t1758 VGND.t1882 203.242
R9704 VGND.t1888 VGND.t1597 203.242
R9705 VGND.t1621 VGND.t1906 203.242
R9706 VGND.t1981 VGND.t1760 203.242
R9707 VGND.t1772 VGND.t1987 203.242
R9708 VGND.t1909 VGND.t1794 203.242
R9709 VGND.t1693 VGND.t1951 203.242
R9710 VGND.t1960 VGND.t1713 203.242
R9711 VGND.t1799 VGND.t2002 203.242
R9712 VGND.t1918 VGND.t1638 203.242
R9713 VGND.t1649 VGND.t1963 203.242
R9714 VGND.t2005 VGND.t1738 203.242
R9715 VGND.t1809 VGND.t2011 203.242
R9716 VGND.t1927 VGND.t1660 203.242
R9717 VGND.t1727 VGND.t1975 203.242
R9718 VGND VGND.n332 194.419
R9719 VGND VGND.n356 194.419
R9720 VGND VGND.n363 194.419
R9721 VGND VGND.n366 194.419
R9722 VGND VGND.n374 194.419
R9723 VGND VGND.n377 194.419
R9724 VGND VGND.n385 194.419
R9725 VGND VGND.n324 194.419
R9726 VGND VGND.n313 194.419
R9727 VGND VGND.n308 194.419
R9728 VGND VGND.n310 194.419
R9729 VGND VGND.n2729 194.419
R9730 VGND VGND.n292 194.419
R9731 VGND VGND.n295 194.419
R9732 VGND VGND.n202 194.419
R9733 VGND.n887 VGND.n886 194.391
R9734 VGND.n1332 VGND.n889 194.391
R9735 VGND.n895 VGND.n893 194.391
R9736 VGND.n931 VGND.n930 194.391
R9737 VGND.n936 VGND.n935 194.391
R9738 VGND.n941 VGND.n940 194.391
R9739 VGND.n946 VGND.n945 194.391
R9740 VGND.n951 VGND.n950 194.391
R9741 VGND.n956 VGND.n955 194.391
R9742 VGND.n961 VGND.n960 194.391
R9743 VGND.n966 VGND.n965 194.391
R9744 VGND.n971 VGND.n970 194.391
R9745 VGND.n976 VGND.n975 194.391
R9746 VGND.n981 VGND.n980 194.391
R9747 VGND.n986 VGND.n985 194.391
R9748 VGND.n1281 VGND.n996 194.391
R9749 VGND.n1274 VGND.n1273 194.391
R9750 VGND.n1231 VGND.n1230 194.391
R9751 VGND.n1236 VGND.n1229 194.391
R9752 VGND.n1227 VGND.n1226 194.391
R9753 VGND.n1243 VGND.n1224 194.391
R9754 VGND.n1222 VGND.n1221 194.391
R9755 VGND.n1217 VGND.n1216 194.391
R9756 VGND.n1211 VGND.n1002 194.391
R9757 VGND.n1204 VGND.n1203 194.391
R9758 VGND.n1008 VGND.n1007 194.391
R9759 VGND.n1185 VGND.n1184 194.391
R9760 VGND.n1179 VGND.n1010 194.391
R9761 VGND.n1172 VGND.n1171 194.391
R9762 VGND.n1169 VGND.n1012 194.391
R9763 VGND.n330 VGND.n329 194.391
R9764 VGND.n396 VGND.n395 194.391
R9765 VGND.n2638 VGND.n2637 194.391
R9766 VGND.n2643 VGND.n2642 194.391
R9767 VGND.n2648 VGND.n2647 194.391
R9768 VGND.n2653 VGND.n2652 194.391
R9769 VGND.n2658 VGND.n2657 194.391
R9770 VGND.n2663 VGND.n2662 194.391
R9771 VGND.n2668 VGND.n2667 194.391
R9772 VGND.n393 VGND.n392 194.391
R9773 VGND.n2714 VGND.n2713 194.391
R9774 VGND.n319 VGND.n318 194.391
R9775 VGND.n2747 VGND.n2746 194.391
R9776 VGND.n303 VGND.n302 194.391
R9777 VGND.n2752 VGND.n2751 194.391
R9778 VGND.n2787 VGND.n2786 194.391
R9779 VGND.n286 VGND.n285 194.391
R9780 VGND.n400 VGND.n399 194.391
R9781 VGND.n2342 VGND.n2341 194.391
R9782 VGND.n2337 VGND.n2336 194.391
R9783 VGND.n2332 VGND.n2331 194.391
R9784 VGND.n2327 VGND.n2326 194.391
R9785 VGND.n2322 VGND.n2321 194.391
R9786 VGND.n2317 VGND.n2316 194.391
R9787 VGND.n2312 VGND.n2311 194.391
R9788 VGND.n2307 VGND.n2306 194.391
R9789 VGND.n2302 VGND.n2301 194.391
R9790 VGND.n2297 VGND.n2296 194.391
R9791 VGND.n2292 VGND.n2291 194.391
R9792 VGND.n2287 VGND.n2286 194.391
R9793 VGND.n414 VGND.n413 194.391
R9794 VGND.n2540 VGND.n2539 194.391
R9795 VGND.n2535 VGND.n416 194.391
R9796 VGND.n469 VGND.n468 194.391
R9797 VGND.n471 VGND.n470 194.391
R9798 VGND.n2376 VGND.n2375 194.391
R9799 VGND.n459 VGND.n458 194.391
R9800 VGND.n2402 VGND.n2401 194.391
R9801 VGND.n451 VGND.n450 194.391
R9802 VGND.n2428 VGND.n2427 194.391
R9803 VGND.n443 VGND.n442 194.391
R9804 VGND.n2454 VGND.n2453 194.391
R9805 VGND.n435 VGND.n434 194.391
R9806 VGND.n2480 VGND.n2479 194.391
R9807 VGND.n427 VGND.n426 194.391
R9808 VGND.n2511 VGND.n2510 194.391
R9809 VGND.n2516 VGND.n2515 194.391
R9810 VGND.n2521 VGND.n2520 194.391
R9811 VGND.n2528 VGND.n418 194.391
R9812 VGND.n466 VGND.n465 194.391
R9813 VGND.n2363 VGND.n2362 194.391
R9814 VGND.n463 VGND.n462 194.391
R9815 VGND.n2389 VGND.n2388 194.391
R9816 VGND.n455 VGND.n454 194.391
R9817 VGND.n2415 VGND.n2414 194.391
R9818 VGND.n447 VGND.n446 194.391
R9819 VGND.n2441 VGND.n2440 194.391
R9820 VGND.n439 VGND.n438 194.391
R9821 VGND.n2467 VGND.n2466 194.391
R9822 VGND.n431 VGND.n430 194.391
R9823 VGND.n2493 VGND.n2492 194.391
R9824 VGND.n423 VGND.n422 194.391
R9825 VGND.n2498 VGND.n2497 194.391
R9826 VGND.n2809 VGND.n2808 194.391
R9827 VGND.n2816 VGND.n276 194.391
R9828 VGND.n625 VGND.n624 194.391
R9829 VGND.n1910 VGND.n1909 194.391
R9830 VGND.n622 VGND.n621 194.391
R9831 VGND.n1921 VGND.n1920 194.391
R9832 VGND.n619 VGND.n618 194.391
R9833 VGND.n1932 VGND.n1931 194.391
R9834 VGND.n616 VGND.n615 194.391
R9835 VGND.n1943 VGND.n1942 194.391
R9836 VGND.n613 VGND.n612 194.391
R9837 VGND.n1954 VGND.n1953 194.391
R9838 VGND.n610 VGND.n609 194.391
R9839 VGND.n1965 VGND.n1964 194.391
R9840 VGND.n607 VGND.n606 194.391
R9841 VGND.n1976 VGND.n1975 194.391
R9842 VGND.n1981 VGND.n1980 194.391
R9843 VGND.n1988 VGND.n605 194.391
R9844 VGND.n590 VGND.n589 194.391
R9845 VGND.n596 VGND.n595 194.391
R9846 VGND.n593 VGND.n592 194.391
R9847 VGND.n2055 VGND.n2054 194.391
R9848 VGND.n2050 VGND.n2049 194.391
R9849 VGND.n2045 VGND.n2044 194.391
R9850 VGND.n2040 VGND.n2039 194.391
R9851 VGND.n2035 VGND.n2034 194.391
R9852 VGND.n2030 VGND.n2029 194.391
R9853 VGND.n2025 VGND.n2024 194.391
R9854 VGND.n2020 VGND.n2019 194.391
R9855 VGND.n2015 VGND.n2014 194.391
R9856 VGND.n2010 VGND.n2009 194.391
R9857 VGND.n2005 VGND.n2004 194.391
R9858 VGND.n2000 VGND.n600 194.391
R9859 VGND.n1995 VGND.n1993 194.391
R9860 VGND.n587 VGND.n586 194.391
R9861 VGND.n2069 VGND.n2068 194.391
R9862 VGND.n2074 VGND.n2073 194.391
R9863 VGND.n2079 VGND.n2078 194.391
R9864 VGND.n2084 VGND.n2083 194.391
R9865 VGND.n2089 VGND.n2088 194.391
R9866 VGND.n2094 VGND.n2093 194.391
R9867 VGND.n2099 VGND.n2098 194.391
R9868 VGND.n2104 VGND.n2103 194.391
R9869 VGND.n2109 VGND.n2108 194.391
R9870 VGND.n2114 VGND.n2113 194.391
R9871 VGND.n2119 VGND.n2118 194.391
R9872 VGND.n584 VGND.n583 194.391
R9873 VGND.n2124 VGND.n2123 194.391
R9874 VGND.n2834 VGND.n2833 194.391
R9875 VGND.n2841 VGND.n264 194.391
R9876 VGND.n547 VGND.n546 194.391
R9877 VGND.n2176 VGND.n549 194.391
R9878 VGND.n1757 VGND.n1755 194.391
R9879 VGND.n1761 VGND.n1760 194.391
R9880 VGND.n1752 VGND.n1751 194.391
R9881 VGND.n1772 VGND.n1771 194.391
R9882 VGND.n1749 VGND.n1748 194.391
R9883 VGND.n1783 VGND.n1782 194.391
R9884 VGND.n1746 VGND.n1745 194.391
R9885 VGND.n1794 VGND.n1793 194.391
R9886 VGND.n1743 VGND.n1742 194.391
R9887 VGND.n1805 VGND.n1804 194.391
R9888 VGND.n1740 VGND.n1739 194.391
R9889 VGND.n1816 VGND.n1815 194.391
R9890 VGND.n1821 VGND.n1820 194.391
R9891 VGND.n1828 VGND.n1738 194.391
R9892 VGND.n628 VGND.n627 194.391
R9893 VGND.n1678 VGND.n1677 194.391
R9894 VGND.n1675 VGND.n1674 194.391
R9895 VGND.n1689 VGND.n1688 194.391
R9896 VGND.n1694 VGND.n1693 194.391
R9897 VGND.n1699 VGND.n1698 194.391
R9898 VGND.n1704 VGND.n1703 194.391
R9899 VGND.n1709 VGND.n1708 194.391
R9900 VGND.n1714 VGND.n1713 194.391
R9901 VGND.n1719 VGND.n1718 194.391
R9902 VGND.n1724 VGND.n1723 194.391
R9903 VGND.n1729 VGND.n1728 194.391
R9904 VGND.n1672 VGND.n1671 194.391
R9905 VGND.n1845 VGND.n1844 194.391
R9906 VGND.n1840 VGND.n1733 194.391
R9907 VGND.n1835 VGND.n1833 194.391
R9908 VGND.n632 VGND.n631 194.391
R9909 VGND.n669 VGND.n668 194.391
R9910 VGND.n674 VGND.n673 194.391
R9911 VGND.n679 VGND.n678 194.391
R9912 VGND.n684 VGND.n683 194.391
R9913 VGND.n689 VGND.n688 194.391
R9914 VGND.n694 VGND.n693 194.391
R9915 VGND.n699 VGND.n698 194.391
R9916 VGND.n704 VGND.n703 194.391
R9917 VGND.n709 VGND.n708 194.391
R9918 VGND.n714 VGND.n713 194.391
R9919 VGND.n719 VGND.n718 194.391
R9920 VGND.n666 VGND.n665 194.391
R9921 VGND.n724 VGND.n723 194.391
R9922 VGND.n2859 VGND.n2858 194.391
R9923 VGND.n2866 VGND.n252 194.391
R9924 VGND.n879 VGND.n878 194.391
R9925 VGND.n1352 VGND.n1351 194.391
R9926 VGND.n874 VGND.n873 194.391
R9927 VGND.n869 VGND.n807 194.391
R9928 VGND.n811 VGND.n809 194.391
R9929 VGND.n823 VGND.n822 194.391
R9930 VGND.n828 VGND.n827 194.391
R9931 VGND.n833 VGND.n832 194.391
R9932 VGND.n838 VGND.n837 194.391
R9933 VGND.n843 VGND.n842 194.391
R9934 VGND.n848 VGND.n847 194.391
R9935 VGND.n819 VGND.n818 194.391
R9936 VGND.n853 VGND.n852 194.391
R9937 VGND.n734 VGND.n733 194.391
R9938 VGND.n1661 VGND.n1660 194.391
R9939 VGND.n1656 VGND.n736 194.391
R9940 VGND.n800 VGND.n799 194.391
R9941 VGND.n1390 VGND.n1389 194.391
R9942 VGND.n1395 VGND.n1394 194.391
R9943 VGND.n804 VGND.n803 194.391
R9944 VGND.n1490 VGND.n1489 194.391
R9945 VGND.n776 VGND.n775 194.391
R9946 VGND.n1516 VGND.n1515 194.391
R9947 VGND.n768 VGND.n767 194.391
R9948 VGND.n1542 VGND.n1541 194.391
R9949 VGND.n1547 VGND.n1546 194.391
R9950 VGND.n760 VGND.n759 194.391
R9951 VGND.n1552 VGND.n1551 194.391
R9952 VGND.n1632 VGND.n1631 194.391
R9953 VGND.n1637 VGND.n1636 194.391
R9954 VGND.n1642 VGND.n1641 194.391
R9955 VGND.n1649 VGND.n739 194.391
R9956 VGND.n797 VGND.n796 194.391
R9957 VGND.n1410 VGND.n1409 194.391
R9958 VGND.n794 VGND.n793 194.391
R9959 VGND.n1477 VGND.n1476 194.391
R9960 VGND.n780 VGND.n779 194.391
R9961 VGND.n1503 VGND.n1502 194.391
R9962 VGND.n772 VGND.n771 194.391
R9963 VGND.n1529 VGND.n1528 194.391
R9964 VGND.n764 VGND.n763 194.391
R9965 VGND.n1566 VGND.n1565 194.391
R9966 VGND.n755 VGND.n754 194.391
R9967 VGND.n1581 VGND.n1580 194.391
R9968 VGND.n1576 VGND.n1575 194.391
R9969 VGND.n1571 VGND.n1570 194.391
R9970 VGND.n2884 VGND.n2883 194.391
R9971 VGND.n2891 VGND.n239 194.391
R9972 VGND.n882 VGND.n881 194.391
R9973 VGND.n884 VGND.n883 194.391
R9974 VGND.n1423 VGND.n1422 194.391
R9975 VGND.n1428 VGND.n1427 194.391
R9976 VGND.n1433 VGND.n1432 194.391
R9977 VGND.n1438 VGND.n1437 194.391
R9978 VGND.n1443 VGND.n1442 194.391
R9979 VGND.n1448 VGND.n1447 194.391
R9980 VGND.n1453 VGND.n1452 194.391
R9981 VGND.n790 VGND.n789 194.391
R9982 VGND.n1458 VGND.n1457 194.391
R9983 VGND.n1595 VGND.n1594 194.391
R9984 VGND.n1600 VGND.n1599 194.391
R9985 VGND.n749 VGND.n748 194.391
R9986 VGND.n1613 VGND.n1612 194.391
R9987 VGND.n1608 VGND.n1604 194.391
R9988 VGND.n1024 VGND.n1023 194.391
R9989 VGND.n1031 VGND.n1030 194.391
R9990 VGND.n1036 VGND.n1035 194.391
R9991 VGND.n1028 VGND.n1027 194.391
R9992 VGND.n1094 VGND.n1093 194.391
R9993 VGND.n1089 VGND.n1088 194.391
R9994 VGND.n1084 VGND.n1083 194.391
R9995 VGND.n1079 VGND.n1078 194.391
R9996 VGND.n1074 VGND.n1073 194.391
R9997 VGND.n1069 VGND.n1040 194.391
R9998 VGND.n1044 VGND.n1042 194.391
R9999 VGND.n1052 VGND.n1051 194.391
R10000 VGND.n1057 VGND.n1056 194.391
R10001 VGND.n1048 VGND.n1047 194.391
R10002 VGND.n2904 VGND.n2903 194.391
R10003 VGND.n2911 VGND.n227 194.391
R10004 VGND.n1014 VGND.n1013 194.391
R10005 VGND.n927 VGND.n926 194.391
R10006 VGND.n2606 VGND.n2605 161.308
R10007 VGND.n2603 VGND.n2602 161.308
R10008 VGND.n2600 VGND.n2599 161.308
R10009 VGND.n2597 VGND.n2596 161.308
R10010 VGND.n2594 VGND.n2593 161.308
R10011 VGND.n2591 VGND.n2590 161.308
R10012 VGND.n2588 VGND.n2587 161.308
R10013 VGND.n2585 VGND.n2584 161.308
R10014 VGND.n2582 VGND.n2581 161.308
R10015 VGND.n2579 VGND.n2578 161.308
R10016 VGND.n2576 VGND.n2575 161.308
R10017 VGND.n2573 VGND.n2572 161.308
R10018 VGND.n2570 VGND.n2569 161.308
R10019 VGND.n2567 VGND.n2566 161.308
R10020 VGND.n2564 VGND.n2563 161.308
R10021 VGND.n2605 VGND.t2696 159.978
R10022 VGND.n2602 VGND.t2699 159.978
R10023 VGND.n2599 VGND.t2694 159.978
R10024 VGND.n2596 VGND.t2689 159.978
R10025 VGND.n2593 VGND.t2695 159.978
R10026 VGND.n2590 VGND.t2702 159.978
R10027 VGND.n2587 VGND.t2698 159.978
R10028 VGND.n2584 VGND.t2692 159.978
R10029 VGND.n2581 VGND.t2688 159.978
R10030 VGND.n2578 VGND.t2690 159.978
R10031 VGND.n2575 VGND.t2701 159.978
R10032 VGND.n2572 VGND.t2693 159.978
R10033 VGND.n2569 VGND.t2700 159.978
R10034 VGND.n2566 VGND.t2697 159.978
R10035 VGND.n2563 VGND.t2703 159.978
R10036 VGND.n123 VGND.t942 159.315
R10037 VGND.n2216 VGND.t1216 159.315
R10038 VGND.n1132 VGND.t1113 158.361
R10039 VGND.n2999 VGND.t1111 158.361
R10040 VGND.n121 VGND.t940 157.291
R10041 VGND.n544 VGND.t1214 157.291
R10042 VGND.n68 VGND.t730 156.915
R10043 VGND.n506 VGND.t133 156.915
R10044 VGND.n68 VGND.t731 156.915
R10045 VGND.n506 VGND.t129 156.915
R10046 VGND.n36 VGND.t1004 154.131
R10047 VGND.n123 VGND.t1064 154.131
R10048 VGND.n128 VGND.t2548 154.131
R10049 VGND.n128 VGND.t2681 154.131
R10050 VGND.n508 VGND.t1441 154.131
R10051 VGND.n508 VGND.t2528 154.131
R10052 VGND.n2216 VGND.t2505 154.131
R10053 VGND.n541 VGND.t2558 154.131
R10054 VGND.n3005 VGND.t1268 153.631
R10055 VGND.n60 VGND.t2553 153.631
R10056 VGND.n160 VGND.t728 153.631
R10057 VGND.n2255 VGND.t128 153.631
R10058 VGND.n2222 VGND.t428 153.631
R10059 VGND.n1360 VGND.t1067 153.631
R10060 VGND.n59 VGND.t946 152.757
R10061 VGND.n2221 VGND.t10 152.757
R10062 VGND.n92 VGND.t735 152.381
R10063 VGND.n2211 VGND.t125 152.381
R10064 VGND.n2181 VGND.n2180 152.174
R10065 VGND.n167 VGND.t738 150.922
R10066 VGND.n167 VGND.t733 150.922
R10067 VGND.n475 VGND.t131 150.922
R10068 VGND.n475 VGND.t123 150.922
R10069 VGND.n166 VGND.t1465 150.922
R10070 VGND.n67 VGND.t2652 150.922
R10071 VGND.n135 VGND.t51 150.922
R10072 VGND.n474 VGND.t2379 150.922
R10073 VGND.n2253 VGND.t1310 150.922
R10074 VGND.n505 VGND.t1011 150.922
R10075 VGND.n166 VGND.t1073 150.922
R10076 VGND.n67 VGND.t2462 150.922
R10077 VGND.n135 VGND.t1170 150.922
R10078 VGND.n474 VGND.t2206 150.922
R10079 VGND.n2253 VGND.t2486 150.922
R10080 VGND.n505 VGND.t2261 150.922
R10081 VGND.n3004 VGND.t207 147.411
R10082 VGND.n159 VGND.t737 147.411
R10083 VGND.n2254 VGND.t127 147.411
R10084 VGND.n1359 VGND.t21 147.411
R10085 VGND.n115 VGND.t2113 146.964
R10086 VGND.n545 VGND.t1408 146.964
R10087 VGND.n2605 VGND.t1914 143.911
R10088 VGND.n2602 VGND.t1989 143.911
R10089 VGND.n2599 VGND.t1893 143.911
R10090 VGND.n2596 VGND.t1938 143.911
R10091 VGND.n2593 VGND.t2013 143.911
R10092 VGND.n2590 VGND.t1920 143.911
R10093 VGND.n2587 VGND.t1890 143.911
R10094 VGND.n2584 VGND.t1932 143.911
R10095 VGND.n2581 VGND.t1944 143.911
R10096 VGND.n2578 VGND.t1875 143.911
R10097 VGND.n2575 VGND.t1968 143.911
R10098 VGND.n2572 VGND.t1896 143.911
R10099 VGND.n2569 VGND.t1971 143.911
R10100 VGND.n2566 VGND.t1998 143.911
R10101 VGND.n2563 VGND.t1941 143.911
R10102 VGND.n1388 VGND.n806 143.478
R10103 VGND VGND.t916 142.089
R10104 VGND.n1021 VGND.t1935 119.309
R10105 VGND.n994 VGND.t1974 119.309
R10106 VGND.n2630 VGND.t1929 119.309
R10107 VGND.n204 VGND.t1965 119.309
R10108 VGND.n334 VGND.t1878 119.309
R10109 VGND.n2626 VGND.t1884 119.309
R10110 VGND.n2623 VGND.t1899 119.309
R10111 VGND.n2620 VGND.t1977 119.309
R10112 VGND.n2617 VGND.t1983 119.309
R10113 VGND.n2614 VGND.t1902 119.309
R10114 VGND.n2611 VGND.t1947 119.309
R10115 VGND.n322 VGND.t1953 119.309
R10116 VGND.n315 VGND.t1992 119.309
R10117 VGND.n306 VGND.t1911 119.309
R10118 VGND.n299 VGND.t1956 119.309
R10119 VGND.n2765 VGND.t1995 119.309
R10120 VGND.n290 VGND.t2007 119.309
R10121 VGND.n297 VGND.t1923 119.309
R10122 VGND.n1018 VGND.t1881 119.309
R10123 VGND.n1015 VGND.t1887 119.309
R10124 VGND.n1180 VGND.t1905 119.309
R10125 VGND.n1006 VGND.t1980 119.309
R10126 VGND.n1004 VGND.t1986 119.309
R10127 VGND.n1195 VGND.t1908 119.309
R10128 VGND.n1212 VGND.t1950 119.309
R10129 VGND.n1000 VGND.t1959 119.309
R10130 VGND.n1253 VGND.t2001 119.309
R10131 VGND.n1256 VGND.t1917 119.309
R10132 VGND.n1259 VGND.t1962 119.309
R10133 VGND.n1262 VGND.t2004 119.309
R10134 VGND.n998 VGND.t2010 119.309
R10135 VGND.n1265 VGND.t1926 119.309
R10136 VGND.n5 VGND.n3 117.001
R10137 VGND.t190 VGND.n5 117.001
R10138 VGND.n6 VGND.n4 117.001
R10139 VGND.n328 VGND.n6 117.001
R10140 VGND.t1752 VGND.t1936 110.535
R10141 VGND.t1162 VGND.t1590 110.535
R10142 VGND.t1882 VGND.t1595 110.535
R10143 VGND.t1670 VGND.t560 110.535
R10144 VGND.t1677 VGND.t1888 110.535
R10145 VGND.t997 VGND.t1685 110.535
R10146 VGND.t1906 VGND.t1699 110.535
R10147 VGND.t1777 VGND.t697 110.535
R10148 VGND.t1764 VGND.t1981 110.535
R10149 VGND.t194 VGND.t1602 110.535
R10150 VGND.t1987 VGND.t1617 110.535
R10151 VGND.t1697 VGND.t2669 110.535
R10152 VGND.t1630 VGND.t1909 110.535
R10153 VGND.t2393 VGND.t1762 110.535
R10154 VGND.t1951 VGND.t1770 110.535
R10155 VGND.t1787 VGND.t779 110.535
R10156 VGND.t1792 VGND.t1960 110.535
R10157 VGND.t1393 VGND.t1629 110.535
R10158 VGND.t2002 VGND.t1615 110.535
R10159 VGND.t1696 VGND.t2521 110.535
R10160 VGND.t1711 VGND.t1918 110.535
R10161 VGND.t1413 VGND.t1790 110.535
R10162 VGND.t1963 VGND.t1720 110.535
R10163 VGND.t1802 VGND.t832 110.535
R10164 VGND.t1634 VGND.t2005 110.535
R10165 VGND.t195 VGND.t1642 110.535
R10166 VGND.t2011 VGND.t1646 110.535
R10167 VGND.t1719 VGND.t630 110.535
R10168 VGND.t1668 VGND.t1927 110.535
R10169 VGND.t1159 VGND.t1740 110.535
R10170 VGND.t1975 VGND.t1805 110.535
R10171 VGND.t1645 VGND.t1200 110.535
R10172 VGND.t1399 VGND.t1409 92.4699
R10173 VGND.t1409 VGND.t1406 92.4699
R10174 VGND.t1406 VGND.t1410 92.4699
R10175 VGND.t1410 VGND.t2278 92.4699
R10176 VGND.t2278 VGND.t981 92.4699
R10177 VGND.t981 VGND.t1543 92.4699
R10178 VGND.t1543 VGND.t1104 92.4699
R10179 VGND VGND.n806 80.9529
R10180 VGND VGND.n806 75.1009
R10181 VGND.n1337 VGND 74.8566
R10182 VGND.t1104 VGND 70.4533
R10183 VGND.n2285 VGND 58.8055
R10184 VGND.n2284 VGND 58.8055
R10185 VGND.n2250 VGND 58.8055
R10186 VGND.n2248 VGND 58.8055
R10187 VGND.n1386 VGND 58.8055
R10188 VGND.n2348 VGND.n2347 53.1823
R10189 VGND.n2349 VGND.n2348 53.1823
R10190 VGND.n3021 VGND.n3020 53.1823
R10191 VGND.n3020 VGND.n3019 53.1823
R10192 VGND.t2120 VGND.t914 50.5752
R10193 VGND.t2116 VGND.t888 50.5752
R10194 VGND.t2110 VGND.t925 50.5752
R10195 VGND.t2112 VGND.t877 50.5752
R10196 VGND.t1407 VGND.t2276 50.5752
R10197 VGND.t1404 VGND.t979 50.5752
R10198 VGND.t1402 VGND.t2266 50.5752
R10199 VGND.t1400 VGND.t2593 50.5752
R10200 VGND VGND.n2981 43.2063
R10201 VGND VGND.n18 43.2063
R10202 VGND VGND.n2951 43.2063
R10203 VGND VGND.n44 43.2063
R10204 VGND.n2347 VGND.n2346 40.6593
R10205 VGND.n886 VGND.t1789 34.8005
R10206 VGND.n886 VGND.t1626 34.8005
R10207 VGND.n889 VGND.t1628 34.8005
R10208 VGND.n889 VGND.t1707 34.8005
R10209 VGND.n893 VGND.t1710 34.8005
R10210 VGND.n893 VGND.t1786 34.8005
R10211 VGND.n930 VGND.t1732 34.8005
R10212 VGND.n930 VGND.t1808 34.8005
R10213 VGND.n935 VGND.t1633 34.8005
R10214 VGND.n935 VGND.t1637 34.8005
R10215 VGND.n940 VGND.t1644 34.8005
R10216 VGND.n940 VGND.t1726 34.8005
R10217 VGND.n945 VGND.t1663 34.8005
R10218 VGND.n945 VGND.t1737 34.8005
R10219 VGND.n950 VGND.t1804 34.8005
R10220 VGND.n950 VGND.t1641 34.8005
R10221 VGND.n955 VGND.t1825 34.8005
R10222 VGND.n955 VGND.t1659 34.8005
R10223 VGND.n960 VGND.t1667 34.8005
R10224 VGND.n960 VGND.t1724 34.8005
R10225 VGND.n965 VGND.t1744 34.8005
R10226 VGND.n965 VGND.t1821 34.8005
R10227 VGND.n970 VGND.t1757 34.8005
R10228 VGND.n970 VGND.t1593 34.8005
R10229 VGND.n975 VGND.t1609 34.8005
R10230 VGND.n975 VGND.t1742 34.8005
R10231 VGND.n980 VGND.t1684 34.8005
R10232 VGND.n980 VGND.t1755 34.8005
R10233 VGND.n985 VGND.t1775 34.8005
R10234 VGND.n985 VGND.t1780 34.8005
R10235 VGND.n996 VGND.t1728 34.8005
R10236 VGND.n996 VGND.t1806 34.8005
R10237 VGND.n1273 VGND.t1661 34.8005
R10238 VGND.n1273 VGND.t1669 34.8005
R10239 VGND.n1230 VGND.t1810 34.8005
R10240 VGND.n1230 VGND.t1647 34.8005
R10241 VGND.n1229 VGND.t1739 34.8005
R10242 VGND.n1229 VGND.t1635 34.8005
R10243 VGND.n1226 VGND.t1650 34.8005
R10244 VGND.n1226 VGND.t1721 34.8005
R10245 VGND.n1224 VGND.t1639 34.8005
R10246 VGND.n1224 VGND.t1712 34.8005
R10247 VGND.n1221 VGND.t1800 34.8005
R10248 VGND.n1221 VGND.t1616 34.8005
R10249 VGND.n1216 VGND.t1714 34.8005
R10250 VGND.n1216 VGND.t1793 34.8005
R10251 VGND.n1002 VGND.t1694 34.8005
R10252 VGND.n1002 VGND.t1771 34.8005
R10253 VGND.n1203 VGND.t1795 34.8005
R10254 VGND.n1203 VGND.t1631 34.8005
R10255 VGND.n1007 VGND.t1773 34.8005
R10256 VGND.n1007 VGND.t1618 34.8005
R10257 VGND.n1184 VGND.t1761 34.8005
R10258 VGND.n1184 VGND.t1765 34.8005
R10259 VGND.n1010 VGND.t1622 34.8005
R10260 VGND.n1010 VGND.t1700 34.8005
R10261 VGND.n1171 VGND.t1598 34.8005
R10262 VGND.n1171 VGND.t1678 34.8005
R10263 VGND.n1012 VGND.t1759 34.8005
R10264 VGND.n1012 VGND.t1596 34.8005
R10265 VGND.n329 VGND.t1734 34.8005
R10266 VGND.n329 VGND.t1812 34.8005
R10267 VGND.n332 VGND.t1814 34.8005
R10268 VGND.n332 VGND.t1652 34.8005
R10269 VGND.n356 VGND.t1654 34.8005
R10270 VGND.n356 VGND.t1730 34.8005
R10271 VGND.n363 VGND.t1676 34.8005
R10272 VGND.n363 VGND.t1750 34.8005
R10273 VGND.n366 VGND.t1816 34.8005
R10274 VGND.n366 VGND.t1819 34.8005
R10275 VGND.n374 VGND.t1827 34.8005
R10276 VGND.n374 VGND.t1674 34.8005
R10277 VGND.n377 VGND.t1607 34.8005
R10278 VGND.n377 VGND.t1688 34.8005
R10279 VGND.n385 VGND.t1746 34.8005
R10280 VGND.n385 VGND.t1823 34.8005
R10281 VGND.n324 VGND.t1769 34.8005
R10282 VGND.n324 VGND.t1605 34.8005
R10283 VGND.n313 VGND.t1611 34.8005
R10284 VGND.n313 VGND.t1672 34.8005
R10285 VGND.n308 VGND.t1692 34.8005
R10286 VGND.n308 VGND.t1767 34.8005
R10287 VGND.n310 VGND.t1704 34.8005
R10288 VGND.n310 VGND.t1782 34.8005
R10289 VGND.n2729 VGND.t1798 34.8005
R10290 VGND.n2729 VGND.t1690 34.8005
R10291 VGND.n292 VGND.t1624 34.8005
R10292 VGND.n292 VGND.t1702 34.8005
R10293 VGND.n295 VGND.t1716 34.8005
R10294 VGND.n295 VGND.t1718 34.8005
R10295 VGND.n202 VGND.t1784 34.8005
R10296 VGND.n202 VGND.t1620 34.8005
R10297 VGND.n395 VGND.t1916 34.8005
R10298 VGND.n395 VGND.t537 34.8005
R10299 VGND.n2637 VGND.t2057 34.8005
R10300 VGND.n2637 VGND.t1271 34.8005
R10301 VGND.n2642 VGND.t1082 34.8005
R10302 VGND.n2642 VGND.t2388 34.8005
R10303 VGND.n2647 VGND.t1830 34.8005
R10304 VGND.n2647 VGND.t2386 34.8005
R10305 VGND.n2652 VGND.t2492 34.8005
R10306 VGND.n2652 VGND.t535 34.8005
R10307 VGND.n2657 VGND.t2565 34.8005
R10308 VGND.n2657 VGND.t2107 34.8005
R10309 VGND.n2662 VGND.t2362 34.8005
R10310 VGND.n2662 VGND.t2105 34.8005
R10311 VGND.n2667 VGND.t553 34.8005
R10312 VGND.n2667 VGND.t533 34.8005
R10313 VGND.n392 VGND.t427 34.8005
R10314 VGND.n392 VGND.t531 34.8005
R10315 VGND.n2713 VGND.t1535 34.8005
R10316 VGND.n2713 VGND.t2109 34.8005
R10317 VGND.n318 VGND.t933 34.8005
R10318 VGND.n318 VGND.t2384 34.8005
R10319 VGND.n2746 VGND.t960 34.8005
R10320 VGND.n2746 VGND.t2382 34.8005
R10321 VGND.n302 VGND.t1447 34.8005
R10322 VGND.n302 VGND.t2103 34.8005
R10323 VGND.n2751 VGND.t92 34.8005
R10324 VGND.n2751 VGND.t2392 34.8005
R10325 VGND.n2786 VGND.t1472 34.8005
R10326 VGND.n2786 VGND.t2390 34.8005
R10327 VGND.n285 VGND.t344 34.8005
R10328 VGND.n285 VGND.t529 34.8005
R10329 VGND.n399 VGND.t1991 34.8005
R10330 VGND.n399 VGND.t1332 34.8005
R10331 VGND.n2341 VGND.t2520 34.8005
R10332 VGND.n2341 VGND.t608 34.8005
R10333 VGND.n2336 VGND.t1308 34.8005
R10334 VGND.n2336 VGND.t1192 34.8005
R10335 VGND.n2331 VGND.t1857 34.8005
R10336 VGND.n2331 VGND.t2252 34.8005
R10337 VGND.n2326 VGND.t236 34.8005
R10338 VGND.n2326 VGND.t1330 34.8005
R10339 VGND.n2321 VGND.t1245 34.8005
R10340 VGND.n2321 VGND.t604 34.8005
R10341 VGND.n2316 VGND.t1176 34.8005
R10342 VGND.n2316 VGND.t602 34.8005
R10343 VGND.n2311 VGND.t578 34.8005
R10344 VGND.n2311 VGND.t1328 34.8005
R10345 VGND.n2306 VGND.t720 34.8005
R10346 VGND.n2306 VGND.t1326 34.8005
R10347 VGND.n2301 VGND.t714 34.8005
R10348 VGND.n2301 VGND.t606 34.8005
R10349 VGND.n2296 VGND.t66 34.8005
R10350 VGND.n2296 VGND.t201 34.8005
R10351 VGND.n2291 VGND.t1209 34.8005
R10352 VGND.n2291 VGND.t199 34.8005
R10353 VGND.n2286 VGND.t1464 34.8005
R10354 VGND.n2286 VGND.t1198 34.8005
R10355 VGND.n413 VGND.t547 34.8005
R10356 VGND.n413 VGND.t1196 34.8005
R10357 VGND.n2539 VGND.t2035 34.8005
R10358 VGND.n2539 VGND.t1194 34.8005
R10359 VGND.n416 VGND.t1525 34.8005
R10360 VGND.n416 VGND.t610 34.8005
R10361 VGND.n468 VGND.t1895 34.8005
R10362 VGND.n468 VGND.t1054 34.8005
R10363 VGND.n470 VGND.t2044 34.8005
R10364 VGND.n470 VGND.t1360 34.8005
R10365 VGND.n2375 VGND.t1049 34.8005
R10366 VGND.n2375 VGND.t1415 34.8005
R10367 VGND.n458 VGND.t1870 34.8005
R10368 VGND.n458 VGND.t1060 34.8005
R10369 VGND.n2401 VGND.t2499 34.8005
R10370 VGND.n2401 VGND.t977 34.8005
R10371 VGND.n450 VGND.t2571 34.8005
R10372 VGND.n450 VGND.t1356 34.8005
R10373 VGND.n2427 VGND.t1365 34.8005
R10374 VGND.n2427 VGND.t1354 34.8005
R10375 VGND.n442 VGND.t559 34.8005
R10376 VGND.n442 VGND.t975 34.8005
R10377 VGND.n2453 VGND.t768 34.8005
R10378 VGND.n2453 VGND.t973 34.8005
R10379 VGND.n434 VGND.t219 34.8005
R10380 VGND.n434 VGND.t1358 34.8005
R10381 VGND.n2479 VGND.t1128 34.8005
R10382 VGND.n2479 VGND.t1058 34.8005
R10383 VGND.n426 VGND.t1027 34.8005
R10384 VGND.n426 VGND.t1056 34.8005
R10385 VGND.n2510 VGND.t1155 34.8005
R10386 VGND.n2510 VGND.t1352 34.8005
R10387 VGND.n2515 VGND.t98 34.8005
R10388 VGND.n2515 VGND.t1419 34.8005
R10389 VGND.n2520 VGND.t674 34.8005
R10390 VGND.n2520 VGND.t1417 34.8005
R10391 VGND.n418 VGND.t351 34.8005
R10392 VGND.n418 VGND.t971 34.8005
R10393 VGND.n465 VGND.t1940 34.8005
R10394 VGND.n465 VGND.t2199 34.8005
R10395 VGND.n2362 VGND.t746 34.8005
R10396 VGND.n2362 VGND.t2226 34.8005
R10397 VGND.n462 VGND.t2248 34.8005
R10398 VGND.n462 VGND.t2555 34.8005
R10399 VGND.n2388 VGND.t1840 34.8005
R10400 VGND.n2388 VGND.t2205 34.8005
R10401 VGND.n454 VGND.t2289 34.8005
R10402 VGND.n454 VGND.t695 34.8005
R10403 VGND.n2414 VGND.t1422 34.8005
R10404 VGND.n2414 VGND.t2222 34.8005
R10405 VGND.n446 VGND.t1388 34.8005
R10406 VGND.n446 VGND.t2220 34.8005
R10407 VGND.n2440 VGND.t419 34.8005
R10408 VGND.n2440 VGND.t693 34.8005
R10409 VGND.n438 VGND.t2543 34.8005
R10410 VGND.n438 VGND.t691 34.8005
R10411 VGND.n2466 VGND.t760 34.8005
R10412 VGND.n2466 VGND.t2224 34.8005
R10413 VGND.n430 VGND.t593 34.8005
R10414 VGND.n430 VGND.t2203 34.8005
R10415 VGND.n2492 VGND.t684 34.8005
R10416 VGND.n2492 VGND.t2201 34.8005
R10417 VGND.n422 VGND.t433 34.8005
R10418 VGND.n422 VGND.t2218 34.8005
R10419 VGND.n2497 VGND.t1263 34.8005
R10420 VGND.n2497 VGND.t2216 34.8005
R10421 VGND.n2808 VGND.t623 34.8005
R10422 VGND.n2808 VGND.t2557 34.8005
R10423 VGND.n276 VGND.t33 34.8005
R10424 VGND.n276 VGND.t689 34.8005
R10425 VGND.n624 VGND.t2015 34.8005
R10426 VGND.n624 VGND.t2197 34.8005
R10427 VGND.n1909 VGND.t1018 34.8005
R10428 VGND.n1909 VGND.t80 34.8005
R10429 VGND.n621 VGND.t2076 34.8005
R10430 VGND.n621 VGND.t1338 34.8005
R10431 VGND.n1920 VGND.t1862 34.8005
R10432 VGND.n1920 VGND.t1119 34.8005
R10433 VGND.n618 VGND.t229 34.8005
R10434 VGND.n618 VGND.t2195 34.8005
R10435 VGND.n1931 VGND.t1123 34.8005
R10436 VGND.n1931 VGND.t76 34.8005
R10437 VGND.n615 VGND.t2260 34.8005
R10438 VGND.n615 VGND.t74 34.8005
R10439 VGND.n1942 VGND.t6 34.8005
R10440 VGND.n1942 VGND.t2193 34.8005
R10441 VGND.n612 VGND.t240 34.8005
R10442 VGND.n612 VGND.t2191 34.8005
R10443 VGND.n1953 VGND.t405 34.8005
R10444 VGND.n1953 VGND.t78 34.8005
R10445 VGND.n609 VGND.t61 34.8005
R10446 VGND.n609 VGND.t1117 34.8005
R10447 VGND.n1964 VGND.t2678 34.8005
R10448 VGND.n1964 VGND.t1115 34.8005
R10449 VGND.n606 VGND.t1044 34.8005
R10450 VGND.n606 VGND.t72 34.8005
R10451 VGND.n1975 VGND.t541 34.8005
R10452 VGND.n1975 VGND.t70 34.8005
R10453 VGND.n1980 VGND.t1521 34.8005
R10454 VGND.n1980 VGND.t1340 34.8005
R10455 VGND.n605 VGND.t443 34.8005
R10456 VGND.n605 VGND.t2189 34.8005
R10457 VGND.n589 VGND.t1922 34.8005
R10458 VGND.n589 VGND.t2234 34.8005
R10459 VGND.n595 VGND.t2055 34.8005
R10460 VGND.n595 VGND.t2684 34.8005
R10461 VGND.n592 VGND.t1080 34.8005
R10462 VGND.n592 VGND.t2575 34.8005
R10463 VGND.n2054 VGND.t1833 34.8005
R10464 VGND.n2054 VGND.t2573 34.8005
R10465 VGND.n2049 VGND.t2490 34.8005
R10466 VGND.n2049 VGND.t2232 34.8005
R10467 VGND.n2044 VGND.t2563 34.8005
R10468 VGND.n2044 VGND.t2585 34.8005
R10469 VGND.n2039 VGND.t2360 34.8005
R10470 VGND.n2039 VGND.t2583 34.8005
R10471 VGND.n2034 VGND.t551 34.8005
R10472 VGND.n2034 VGND.t2230 34.8005
R10473 VGND.n2029 VGND.t425 34.8005
R10474 VGND.n2029 VGND.t2228 34.8005
R10475 VGND.n2024 VGND.t1533 34.8005
R10476 VGND.n2024 VGND.t2587 34.8005
R10477 VGND.n2019 VGND.t930 34.8005
R10478 VGND.n2019 VGND.t2238 34.8005
R10479 VGND.n2014 VGND.t958 34.8005
R10480 VGND.n2014 VGND.t2236 34.8005
R10481 VGND.n2009 VGND.t1444 34.8005
R10482 VGND.n2009 VGND.t2581 34.8005
R10483 VGND.n2004 VGND.t90 34.8005
R10484 VGND.n2004 VGND.t2579 34.8005
R10485 VGND.n600 VGND.t1516 34.8005
R10486 VGND.n600 VGND.t2577 34.8005
R10487 VGND.n1993 VGND.t342 34.8005
R10488 VGND.n1993 VGND.t2686 34.8005
R10489 VGND.n586 VGND.t1892 34.8005
R10490 VGND.n586 VGND.t649 34.8005
R10491 VGND.n2068 VGND.t2046 34.8005
R10492 VGND.n2068 VGND.t1240 34.8005
R10493 VGND.n2073 VGND.t1051 34.8005
R10494 VGND.n2073 VGND.t612 34.8005
R10495 VGND.n2078 VGND.t1868 34.8005
R10496 VGND.n2078 VGND.t655 34.8005
R10497 VGND.n2083 VGND.t2501 34.8005
R10498 VGND.n2083 VGND.t647 34.8005
R10499 VGND.n2088 VGND.t2560 34.8005
R10500 VGND.n2088 VGND.t1236 34.8005
R10501 VGND.n2093 VGND.t1367 34.8005
R10502 VGND.n2093 VGND.t1234 34.8005
R10503 VGND.n2098 VGND.t1 34.8005
R10504 VGND.n2098 VGND.t645 34.8005
R10505 VGND.n2103 VGND.t770 34.8005
R10506 VGND.n2103 VGND.t643 34.8005
R10507 VGND.n2108 VGND.t221 34.8005
R10508 VGND.n2108 VGND.t1238 34.8005
R10509 VGND.n2113 VGND.t1130 34.8005
R10510 VGND.n2113 VGND.t653 34.8005
R10511 VGND.n2118 VGND.t1029 34.8005
R10512 VGND.n2118 VGND.t651 34.8005
R10513 VGND.n583 VGND.t1157 34.8005
R10514 VGND.n583 VGND.t1232 34.8005
R10515 VGND.n2123 VGND.t100 34.8005
R10516 VGND.n2123 VGND.t616 34.8005
R10517 VGND.n2833 VGND.t676 34.8005
R10518 VGND.n2833 VGND.t614 34.8005
R10519 VGND.n264 VGND.t353 34.8005
R10520 VGND.n264 VGND.t641 34.8005
R10521 VGND.n546 VGND.t1934 34.8005
R10522 VGND.n546 VGND.t752 34.8005
R10523 VGND.n549 VGND.t748 34.8005
R10524 VGND.n549 VGND.t203 34.8005
R10525 VGND.n1755 VGND.t2250 34.8005
R10526 VGND.n1755 VGND.t2088 34.8005
R10527 VGND.n1760 VGND.t1838 34.8005
R10528 VGND.n1760 VGND.t2086 34.8005
R10529 VGND.n1751 VGND.t2291 34.8005
R10530 VGND.n1751 VGND.t1225 34.8005
R10531 VGND.n1771 VGND.t1424 34.8005
R10532 VGND.n1771 VGND.t2212 34.8005
R10533 VGND.n1748 VGND.t1390 34.8005
R10534 VGND.n1748 VGND.t2210 34.8005
R10535 VGND.n1782 VGND.t421 34.8005
R10536 VGND.n1782 VGND.t1223 34.8005
R10537 VGND.n1745 VGND.t2545 34.8005
R10538 VGND.n1745 VGND.t1221 34.8005
R10539 VGND.n1793 VGND.t762 34.8005
R10540 VGND.n1793 VGND.t2214 34.8005
R10541 VGND.n1742 VGND.t595 34.8005
R10542 VGND.n1742 VGND.t756 34.8005
R10543 VGND.n1804 VGND.t686 34.8005
R10544 VGND.n1804 VGND.t754 34.8005
R10545 VGND.n1739 VGND.t435 34.8005
R10546 VGND.n1739 VGND.t2208 34.8005
R10547 VGND.n1815 VGND.t1265 34.8005
R10548 VGND.n1815 VGND.t2092 34.8005
R10549 VGND.n1820 VGND.t625 34.8005
R10550 VGND.n1820 VGND.t2090 34.8005
R10551 VGND.n1738 VGND.t35 34.8005
R10552 VGND.n1738 VGND.t1219 34.8005
R10553 VGND.n627 VGND.t1946 34.8005
R10554 VGND.n627 VGND.t1150 34.8005
R10555 VGND.n1677 VGND.t741 34.8005
R10556 VGND.n1677 VGND.t2098 34.8005
R10557 VGND.n1674 VGND.t1167 34.8005
R10558 VGND.n1674 VGND.t84 34.8005
R10559 VGND.n1688 VGND.t1844 34.8005
R10560 VGND.n1688 VGND.t1038 34.8005
R10561 VGND.n1693 VGND.t215 34.8005
R10562 VGND.n1693 VGND.t1148 34.8005
R10563 VGND.n1698 VGND.t704 34.8005
R10564 VGND.n1698 VGND.t1348 34.8005
R10565 VGND.n1703 VGND.t1386 34.8005
R10566 VGND.n1703 VGND.t1346 34.8005
R10567 VGND.n1708 VGND.t415 34.8005
R10568 VGND.n1708 VGND.t1146 34.8005
R10569 VGND.n1713 VGND.t2539 34.8005
R10570 VGND.n1713 VGND.t1144 34.8005
R10571 VGND.n1718 VGND.t569 34.8005
R10572 VGND.n1718 VGND.t1350 34.8005
R10573 VGND.n1723 VGND.t591 34.8005
R10574 VGND.n1723 VGND.t1036 34.8005
R10575 VGND.n1728 VGND.t1142 34.8005
R10576 VGND.n1728 VGND.t1034 34.8005
R10577 VGND.n1671 VGND.t431 34.8005
R10578 VGND.n1671 VGND.t1344 34.8005
R10579 VGND.n1844 VGND.t638 34.8005
R10580 VGND.n1844 VGND.t1342 34.8005
R10581 VGND.n1733 VGND.t619 34.8005
R10582 VGND.n1733 VGND.t86 34.8005
R10583 VGND.n1833 VGND.t31 34.8005
R10584 VGND.n1833 VGND.t2100 34.8005
R10585 VGND.n631 VGND.t1877 34.8005
R10586 VGND.n631 VGND.t1436 34.8005
R10587 VGND.n668 VGND.t1016 34.8005
R10588 VGND.n668 VGND.t1426 34.8005
R10589 VGND.n673 VGND.t2074 34.8005
R10590 VGND.n673 VGND.t1514 34.8005
R10591 VGND.n678 VGND.t1864 34.8005
R10592 VGND.n678 VGND.t1512 34.8005
R10593 VGND.n683 VGND.t227 34.8005
R10594 VGND.n683 VGND.t1434 34.8005
R10595 VGND.n688 VGND.t1121 34.8005
R10596 VGND.n688 VGND.t1504 34.8005
R10597 VGND.n693 VGND.t2258 34.8005
R10598 VGND.n693 VGND.t1502 34.8005
R10599 VGND.n698 VGND.t4 34.8005
R10600 VGND.n698 VGND.t1432 34.8005
R10601 VGND.n703 VGND.t238 34.8005
R10602 VGND.n703 VGND.t1430 34.8005
R10603 VGND.n708 VGND.t403 34.8005
R10604 VGND.n708 VGND.t1506 34.8005
R10605 VGND.n713 VGND.t1134 34.8005
R10606 VGND.n713 VGND.t1510 34.8005
R10607 VGND.n718 VGND.t2676 34.8005
R10608 VGND.n718 VGND.t1508 34.8005
R10609 VGND.n665 VGND.t1042 34.8005
R10610 VGND.n665 VGND.t1500 34.8005
R10611 VGND.n723 VGND.t539 34.8005
R10612 VGND.n723 VGND.t1498 34.8005
R10613 VGND.n2858 VGND.t1519 34.8005
R10614 VGND.n2858 VGND.t1496 34.8005
R10615 VGND.n252 VGND.t441 34.8005
R10616 VGND.n252 VGND.t1428 34.8005
R10617 VGND.n878 VGND.t1970 34.8005
R10618 VGND.n878 VGND.t1585 34.8005
R10619 VGND.n1351 VGND.t1071 34.8005
R10620 VGND.n1351 VGND.t1563 34.8005
R10621 VGND.n873 VGND.t1098 34.8005
R10622 VGND.n873 VGND.t1577 34.8005
R10623 VGND.n807 VGND.t1848 34.8005
R10624 VGND.n807 VGND.t1579 34.8005
R10625 VGND.n809 VGND.t209 34.8005
R10626 VGND.n809 VGND.t1587 34.8005
R10627 VGND.n822 VGND.t573 34.8005
R10628 VGND.n822 VGND.t1567 34.8005
R10629 VGND.n827 VGND.t1183 34.8005
R10630 VGND.n827 VGND.t1569 34.8005
R10631 VGND.n832 VGND.t408 34.8005
R10632 VGND.n832 VGND.t1557 34.8005
R10633 VGND.n837 VGND.t773 34.8005
R10634 VGND.n837 VGND.t1559 34.8005
R10635 VGND.n842 VGND.t2485 34.8005
R10636 VGND.n842 VGND.t1565 34.8005
R10637 VGND.n847 VGND.t2024 34.8005
R10638 VGND.n847 VGND.t1581 34.8005
R10639 VGND.n818 VGND.t2125 34.8005
R10640 VGND.n818 VGND.t1583 34.8005
R10641 VGND.n852 VGND.t2344 34.8005
R10642 VGND.n852 VGND.t1571 34.8005
R10643 VGND.n733 VGND.t2478 34.8005
R10644 VGND.n733 VGND.t1573 34.8005
R10645 VGND.n1660 VGND.t2028 34.8005
R10646 VGND.n1660 VGND.t1575 34.8005
R10647 VGND.n736 VGND.t23 34.8005
R10648 VGND.n736 VGND.t1561 34.8005
R10649 VGND.n799 VGND.t1898 34.8005
R10650 VGND.n799 VGND.t2664 34.8005
R10651 VGND.n1389 VGND.t2042 34.8005
R10652 VGND.n1389 VGND.t1284 34.8005
R10653 VGND.n1394 VGND.t1047 34.8005
R10654 VGND.n1394 VGND.t2065 34.8005
R10655 VGND.n803 VGND.t1872 34.8005
R10656 VGND.n803 VGND.t2063 34.8005
R10657 VGND.n1489 VGND.t2497 34.8005
R10658 VGND.n1489 VGND.t2662 34.8005
R10659 VGND.n775 VGND.t2569 34.8005
R10660 VGND.n775 VGND.t1280 34.8005
R10661 VGND.n1515 VGND.t1363 34.8005
R10662 VGND.n1515 VGND.t1278 34.8005
R10663 VGND.n767 VGND.t557 34.8005
R10664 VGND.n767 VGND.t2660 34.8005
R10665 VGND.n1541 VGND.t766 34.8005
R10666 VGND.n1541 VGND.t2658 34.8005
R10667 VGND.n1546 VGND.t1539 34.8005
R10668 VGND.n1546 VGND.t1282 34.8005
R10669 VGND.n759 VGND.t937 34.8005
R10670 VGND.n759 VGND.t2668 34.8005
R10671 VGND.n1551 VGND.t1025 34.8005
R10672 VGND.n1551 VGND.t2666 34.8005
R10673 VGND.n1631 VGND.t1153 34.8005
R10674 VGND.n1631 VGND.t1276 34.8005
R10675 VGND.n1636 VGND.t96 34.8005
R10676 VGND.n1636 VGND.t2069 34.8005
R10677 VGND.n1641 VGND.t1476 34.8005
R10678 VGND.n1641 VGND.t2067 34.8005
R10679 VGND.n739 VGND.t349 34.8005
R10680 VGND.n739 VGND.t1286 34.8005
R10681 VGND.n796 VGND.t1973 34.8005
R10682 VGND.n796 VGND.t1317 34.8005
R10683 VGND.n1409 VGND.t1069 34.8005
R10684 VGND.n1409 VGND.t1372 34.8005
R10685 VGND.n793 VGND.t1096 34.8005
R10686 VGND.n793 VGND.t2177 34.8005
R10687 VGND.n1476 VGND.t1850 34.8005
R10688 VGND.n1476 VGND.t1323 34.8005
R10689 VGND.n779 VGND.t2072 34.8005
R10690 VGND.n779 VGND.t1380 34.8005
R10691 VGND.n1502 VGND.t1554 34.8005
R10692 VGND.n1502 VGND.t2187 34.8005
R10693 VGND.n771 VGND.t1181 34.8005
R10694 VGND.n771 VGND.t2185 34.8005
R10695 VGND.n1528 VGND.t584 34.8005
R10696 VGND.n1528 VGND.t1378 34.8005
R10697 VGND.n763 VGND.t2533 34.8005
R10698 VGND.n763 VGND.t1376 34.8005
R10699 VGND.n1565 VGND.t2483 34.8005
R10700 VGND.n1565 VGND.t1370 34.8005
R10701 VGND.n754 VGND.t2022 34.8005
R10702 VGND.n754 VGND.t1321 34.8005
R10703 VGND.n1580 VGND.t2123 34.8005
R10704 VGND.n1580 VGND.t1319 34.8005
R10705 VGND.n1575 VGND.t2096 34.8005
R10706 VGND.n1575 VGND.t2183 34.8005
R10707 VGND.n1570 VGND.t2476 34.8005
R10708 VGND.n1570 VGND.t2181 34.8005
R10709 VGND.n2883 VGND.t629 34.8005
R10710 VGND.n2883 VGND.t2179 34.8005
R10711 VGND.n239 VGND.t2287 34.8005
R10712 VGND.n239 VGND.t1374 34.8005
R10713 VGND.n881 VGND.t2000 34.8005
R10714 VGND.n881 VGND.t1488 34.8005
R10715 VGND.n883 VGND.t2518 34.8005
R10716 VGND.n883 VGND.t1292 34.8005
R10717 VGND.n1422 VGND.t1306 34.8005
R10718 VGND.n1422 VGND.t1248 34.8005
R10719 VGND.n1427 VGND.t1860 34.8005
R10720 VGND.n1427 VGND.t1494 34.8005
R10721 VGND.n1432 VGND.t233 34.8005
R10722 VGND.n1432 VGND.t1486 34.8005
R10723 VGND.n1437 VGND.t1243 34.8005
R10724 VGND.n1437 VGND.t1288 34.8005
R10725 VGND.n1442 VGND.t1174 34.8005
R10726 VGND.n1442 VGND.t1256 34.8005
R10727 VGND.n1447 VGND.t576 34.8005
R10728 VGND.n1447 VGND.t1298 34.8005
R10729 VGND.n1452 VGND.t718 34.8005
R10730 VGND.n1452 VGND.t1296 34.8005
R10731 VGND.n789 VGND.t712 34.8005
R10732 VGND.n789 VGND.t1290 34.8005
R10733 VGND.n1457 VGND.t63 34.8005
R10734 VGND.n1457 VGND.t1492 34.8005
R10735 VGND.n1594 VGND.t1207 34.8005
R10736 VGND.n1594 VGND.t1490 34.8005
R10737 VGND.n1599 VGND.t1461 34.8005
R10738 VGND.n1599 VGND.t1254 34.8005
R10739 VGND.n748 VGND.t545 34.8005
R10740 VGND.n748 VGND.t1252 34.8005
R10741 VGND.n1612 VGND.t2032 34.8005
R10742 VGND.n1612 VGND.t1250 34.8005
R10743 VGND.n1604 VGND.t447 34.8005
R10744 VGND.n1604 VGND.t1294 34.8005
R10745 VGND.n1023 VGND.t1943 34.8005
R10746 VGND.n1023 VGND.t1484 34.8005
R10747 VGND.n1030 VGND.t743 34.8005
R10748 VGND.n1030 VGND.t967 34.8005
R10749 VGND.n1035 VGND.t1169 34.8005
R10750 VGND.n1035 VGND.t722 34.8005
R10751 VGND.n1027 VGND.t1842 34.8005
R10752 VGND.n1027 VGND.t2244 34.8005
R10753 VGND.n1093 VGND.t217 34.8005
R10754 VGND.n1093 VGND.t1482 34.8005
R10755 VGND.n1088 VGND.t706 34.8005
R10756 VGND.n1088 VGND.t2082 34.8005
R10757 VGND.n1083 VGND.t1384 34.8005
R10758 VGND.n1083 VGND.t2080 34.8005
R10759 VGND.n1078 VGND.t413 34.8005
R10760 VGND.n1078 VGND.t1480 34.8005
R10761 VGND.n1073 VGND.t2537 34.8005
R10762 VGND.n1073 VGND.t1478 34.8005
R10763 VGND.n1040 VGND.t567 34.8005
R10764 VGND.n1040 VGND.t2084 34.8005
R10765 VGND.n1042 VGND.t589 34.8005
R10766 VGND.n1042 VGND.t2242 34.8005
R10767 VGND.n1051 VGND.t1140 34.8005
R10768 VGND.n1051 VGND.t2240 34.8005
R10769 VGND.n1056 VGND.t2348 34.8005
R10770 VGND.n1056 VGND.t2078 34.8005
R10771 VGND.n1047 VGND.t636 34.8005
R10772 VGND.n1047 VGND.t726 34.8005
R10773 VGND.n2903 VGND.t621 34.8005
R10774 VGND.n2903 VGND.t724 34.8005
R10775 VGND.n227 VGND.t29 34.8005
R10776 VGND.n227 VGND.t969 34.8005
R10777 VGND.n1013 VGND.t1682 34.8005
R10778 VGND.n1013 VGND.t1753 34.8005
R10779 VGND.n926 VGND.t1600 34.8005
R10780 VGND.n926 VGND.t1680 34.8005
R10781 VGND.n105 VGND.n103 34.6358
R10782 VGND.n2984 VGND.n2978 34.6358
R10783 VGND.n2987 VGND.n2986 34.6358
R10784 VGND.n2987 VGND.n2974 34.6358
R10785 VGND.n2991 VGND.n2974 34.6358
R10786 VGND.n2992 VGND.n2991 34.6358
R10787 VGND.n2993 VGND.n2992 34.6358
R10788 VGND.n21 VGND.n20 34.6358
R10789 VGND.n23 VGND.n12 34.6358
R10790 VGND.n27 VGND.n12 34.6358
R10791 VGND.n28 VGND.n27 34.6358
R10792 VGND.n29 VGND.n28 34.6358
R10793 VGND.n29 VGND.n9 34.6358
R10794 VGND.n3006 VGND.n10 34.6358
R10795 VGND.n181 VGND.n180 34.6358
R10796 VGND.n185 VGND.n184 34.6358
R10797 VGND.n2954 VGND.n2953 34.6358
R10798 VGND.n2956 VGND.n2947 34.6358
R10799 VGND.n2960 VGND.n2947 34.6358
R10800 VGND.n2961 VGND.n2960 34.6358
R10801 VGND.n2962 VGND.n2961 34.6358
R10802 VGND.n2962 VGND.n2945 34.6358
R10803 VGND.n47 VGND.n46 34.6358
R10804 VGND.n49 VGND.n38 34.6358
R10805 VGND.n53 VGND.n38 34.6358
R10806 VGND.n54 VGND.n53 34.6358
R10807 VGND.n55 VGND.n54 34.6358
R10808 VGND.n55 VGND.n35 34.6358
R10809 VGND.n109 VGND.n108 34.6358
R10810 VGND.n82 VGND.n81 34.6358
R10811 VGND.n86 VGND.n85 34.6358
R10812 VGND.n150 VGND.n149 34.6358
R10813 VGND.n154 VGND.n153 34.6358
R10814 VGND.n1153 VGND.n1135 34.6358
R10815 VGND.n1149 VGND.n1135 34.6358
R10816 VGND.n1149 VGND.n1148 34.6358
R10817 VGND.n1148 VGND.n1147 34.6358
R10818 VGND.n1147 VGND.n1137 34.6358
R10819 VGND.n1131 VGND.n1105 34.6358
R10820 VGND.n1126 VGND.n1106 34.6358
R10821 VGND.n1122 VGND.n1106 34.6358
R10822 VGND.n1122 VGND.n1121 34.6358
R10823 VGND.n1121 VGND.n1120 34.6358
R10824 VGND.n1120 VGND.n1108 34.6358
R10825 VGND.n486 VGND.n481 34.6358
R10826 VGND.n491 VGND.n490 34.6358
R10827 VGND.n2267 VGND.n2262 34.6358
R10828 VGND.n2272 VGND.n2271 34.6358
R10829 VGND.n522 VGND.n517 34.6358
R10830 VGND.n527 VGND.n526 34.6358
R10831 VGND.n2196 VGND.n2195 34.6358
R10832 VGND.n2204 VGND.n2203 34.6358
R10833 VGND.n2200 VGND.n2199 34.6358
R10834 VGND.n2243 VGND.n542 34.6358
R10835 VGND.n2243 VGND.n2242 34.6358
R10836 VGND.n2242 VGND.n2241 34.6358
R10837 VGND.n2241 VGND.n2227 34.6358
R10838 VGND.n2237 VGND.n2227 34.6358
R10839 VGND.n1361 VGND.n1356 34.6358
R10840 VGND.n1381 VGND.n1357 34.6358
R10841 VGND.n1381 VGND.n1380 34.6358
R10842 VGND.n1380 VGND.n1379 34.6358
R10843 VGND.n1379 VGND.n1365 34.6358
R10844 VGND.n1375 VGND.n1365 34.6358
R10845 VGND.n2998 VGND.n2997 34.6358
R10846 VGND.n2 VGND.t191 34.4422
R10847 VGND.n122 VGND.n121 33.1299
R10848 VGND.n2215 VGND.n544 33.1299
R10849 VGND.n111 VGND.n93 32.377
R10850 VGND.n187 VGND.n186 32.377
R10851 VGND.n111 VGND.n110 32.377
R10852 VGND.n88 VGND.n87 32.377
R10853 VGND.n156 VGND.n155 32.377
R10854 VGND.n2206 VGND.n2205 32.377
R10855 VGND.n2206 VGND.n2184 32.0005
R10856 VGND.n497 VGND.n494 30.4946
R10857 VGND.n2278 VGND.n2275 30.4946
R10858 VGND.n533 VGND.n530 30.4946
R10859 VGND.n190 VGND.n167 29.8709
R10860 VGND.n1143 VGND.n1142 28.9887
R10861 VGND.n1116 VGND.n1115 28.9887
R10862 VGND.n2235 VGND.n2234 28.9887
R10863 VGND.n1373 VGND.n1372 28.9887
R10864 VGND.n2985 VGND.n2984 27.8593
R10865 VGND.n22 VGND.n21 27.8593
R10866 VGND.n2955 VGND.n2954 27.8593
R10867 VGND.n48 VGND.n47 27.8593
R10868 VGND.n2256 VGND.n2255 27.0003
R10869 VGND.n161 VGND.n160 26.8591
R10870 VGND.n184 VGND.n173 26.3534
R10871 VGND.n108 VGND.n98 26.3534
R10872 VGND.n85 VGND.n74 26.3534
R10873 VGND.n153 VGND.n142 26.3534
R10874 VGND.n2203 VGND.n2188 26.3534
R10875 VGND.n129 VGND.n68 25.977
R10876 VGND.n498 VGND.n497 25.977
R10877 VGND.n2279 VGND.n2278 25.977
R10878 VGND.n534 VGND.n533 25.977
R10879 VGND.n509 VGND.n506 25.977
R10880 VGND.n2980 VGND.t913 24.9236
R10881 VGND.n2980 VGND.t867 24.9236
R10882 VGND.n2979 VGND.t904 24.9236
R10883 VGND.n2979 VGND.t850 24.9236
R10884 VGND.n2977 VGND.t924 24.9236
R10885 VGND.n2977 VGND.t897 24.9236
R10886 VGND.n2976 VGND.t909 24.9236
R10887 VGND.n2976 VGND.t883 24.9236
R10888 VGND.n17 VGND.t896 24.9236
R10889 VGND.n17 VGND.t928 24.9236
R10890 VGND.n16 VGND.t854 24.9236
R10891 VGND.n16 VGND.t891 24.9236
R10892 VGND.n15 VGND.t902 24.9236
R10893 VGND.n15 VGND.t872 24.9236
R10894 VGND.n14 VGND.t864 24.9236
R10895 VGND.n14 VGND.t920 24.9236
R10896 VGND.n176 VGND.t844 24.9236
R10897 VGND.n176 VGND.t885 24.9236
R10898 VGND.n175 VGND.t900 24.9236
R10899 VGND.n175 VGND.t842 24.9236
R10900 VGND.n172 VGND.t852 24.9236
R10901 VGND.n172 VGND.t1467 24.9236
R10902 VGND.n171 VGND.t906 24.9236
R10903 VGND.n171 VGND.t54 24.9236
R10904 VGND.n170 VGND.t1466 24.9236
R10905 VGND.n170 VGND.t1469 24.9236
R10906 VGND.n169 VGND.t709 24.9236
R10907 VGND.n169 VGND.t2680 24.9236
R10908 VGND.n2950 VGND.t917 24.9236
R10909 VGND.n2950 VGND.t838 24.9236
R10910 VGND.n2949 VGND.t848 24.9236
R10911 VGND.n2949 VGND.t856 24.9236
R10912 VGND.n43 VGND.t870 24.9236
R10913 VGND.n43 VGND.t905 24.9236
R10914 VGND.n42 VGND.t858 24.9236
R10915 VGND.n42 VGND.t895 24.9236
R10916 VGND.n41 VGND.t879 24.9236
R10917 VGND.n41 VGND.t840 24.9236
R10918 VGND.n40 VGND.t866 24.9236
R10919 VGND.n40 VGND.t921 24.9236
R10920 VGND.n96 VGND.t889 24.9236
R10921 VGND.n96 VGND.t926 24.9236
R10922 VGND.n97 VGND.t893 24.9236
R10923 VGND.n97 VGND.t2121 24.9236
R10924 VGND.n95 VGND.t2117 24.9236
R10925 VGND.n95 VGND.t2111 24.9236
R10926 VGND.n100 VGND.t836 24.9236
R10927 VGND.n100 VGND.t919 24.9236
R10928 VGND.n77 VGND.t880 24.9236
R10929 VGND.n77 VGND.t912 24.9236
R10930 VGND.n76 VGND.t860 24.9236
R10931 VGND.n76 VGND.t899 24.9236
R10932 VGND.n73 VGND.t884 24.9236
R10933 VGND.n73 VGND.t2654 24.9236
R10934 VGND.n72 VGND.t869 24.9236
R10935 VGND.n72 VGND.t2470 24.9236
R10936 VGND.n71 VGND.t2653 24.9236
R10937 VGND.n71 VGND.t2651 24.9236
R10938 VGND.n70 VGND.t2466 24.9236
R10939 VGND.n70 VGND.t2460 24.9236
R10940 VGND.n145 VGND.t876 24.9236
R10941 VGND.n145 VGND.t907 24.9236
R10942 VGND.n144 VGND.t922 24.9236
R10943 VGND.n144 VGND.t874 24.9236
R10944 VGND.n141 VGND.t881 24.9236
R10945 VGND.n141 VGND.t57 24.9236
R10946 VGND.n140 VGND.t834 24.9236
R10947 VGND.n140 VGND.t2370 24.9236
R10948 VGND.n139 VGND.t48 24.9236
R10949 VGND.n139 VGND.t2017 24.9236
R10950 VGND.n138 VGND.t289 24.9236
R10951 VGND.n138 VGND.t1076 24.9236
R10952 VGND.n1139 VGND.t2279 24.9236
R10953 VGND.n1139 VGND.t982 24.9236
R10954 VGND.n1141 VGND.t1544 24.9236
R10955 VGND.n1141 VGND.t1105 24.9236
R10956 VGND.n1111 VGND.t666 24.9236
R10957 VGND.n1111 VGND.t667 24.9236
R10958 VGND.n1110 VGND.t2280 24.9236
R10959 VGND.n1110 VGND.t985 24.9236
R10960 VGND.n1114 VGND.t37 24.9236
R10961 VGND.n1114 VGND.t1548 24.9236
R10962 VGND.n1113 VGND.t1545 24.9236
R10963 VGND.n1113 VGND.t1106 24.9236
R10964 VGND.n488 VGND.t664 24.9236
R10965 VGND.n488 VGND.t2283 24.9236
R10966 VGND.n487 VGND.t2597 24.9236
R10967 VGND.n487 VGND.t2272 24.9236
R10968 VGND.n478 VGND.t750 24.9236
R10969 VGND.n478 VGND.t663 24.9236
R10970 VGND.n477 VGND.t2376 24.9236
R10971 VGND.n477 VGND.t2596 24.9236
R10972 VGND.n496 VGND.t1091 24.9236
R10973 VGND.n496 VGND.t749 24.9236
R10974 VGND.n495 VGND.t2378 24.9236
R10975 VGND.n495 VGND.t2377 24.9236
R10976 VGND.n2269 VGND.t1547 24.9236
R10977 VGND.n2269 VGND.t2590 24.9236
R10978 VGND.n2268 VGND.t988 24.9236
R10979 VGND.n2268 VGND.t2270 24.9236
R10980 VGND.n2259 VGND.t1074 24.9236
R10981 VGND.n2259 VGND.t1542 24.9236
R10982 VGND.n2258 VGND.t2687 24.9236
R10983 VGND.n2258 VGND.t978 24.9236
R10984 VGND.n2277 VGND.t998 24.9236
R10985 VGND.n2277 VGND.t999 24.9236
R10986 VGND.n2276 VGND.t15 24.9236
R10987 VGND.n2276 VGND.t17 24.9236
R10988 VGND.n524 VGND.t2599 24.9236
R10989 VGND.n524 VGND.t2275 24.9236
R10990 VGND.n523 VGND.t2592 24.9236
R10991 VGND.n523 VGND.t40 24.9236
R10992 VGND.n514 VGND.t2262 24.9236
R10993 VGND.n514 VGND.t2598 24.9236
R10994 VGND.n513 VGND.t1012 24.9236
R10995 VGND.n513 VGND.t659 24.9236
R10996 VGND.n532 VGND.t2264 24.9236
R10997 VGND.n532 VGND.t2263 24.9236
R10998 VGND.n531 VGND.t1014 24.9236
R10999 VGND.n531 VGND.t1013 24.9236
R11000 VGND.n2186 VGND.t980 24.9236
R11001 VGND.n2186 VGND.t2267 24.9236
R11002 VGND.n2187 VGND.t1401 24.9236
R11003 VGND.n2187 VGND.t990 24.9236
R11004 VGND.n2185 VGND.t1405 24.9236
R11005 VGND.n2185 VGND.t1403 24.9236
R11006 VGND.n2190 VGND.t1541 24.9236
R11007 VGND.n2190 VGND.t1103 24.9236
R11008 VGND.n2230 VGND.t2281 24.9236
R11009 VGND.n2230 VGND.t986 24.9236
R11010 VGND.n2229 VGND.t42 24.9236
R11011 VGND.n2229 VGND.t2273 24.9236
R11012 VGND.n2233 VGND.t1546 24.9236
R11013 VGND.n2233 VGND.t964 24.9236
R11014 VGND.n2231 VGND.t983 24.9236
R11015 VGND.n2231 VGND.t2268 24.9236
R11016 VGND.n1368 VGND.t661 24.9236
R11017 VGND.n1368 VGND.t662 24.9236
R11018 VGND.n1367 VGND.t2269 24.9236
R11019 VGND.n1367 VGND.t1100 24.9236
R11020 VGND.n1371 VGND.t2265 24.9236
R11021 VGND.n1371 VGND.t665 24.9236
R11022 VGND.n1369 VGND.t2591 24.9236
R11023 VGND.n1369 VGND.t38 24.9236
R11024 VGND.n187 VGND.n166 24.4711
R11025 VGND.n61 VGND.n36 24.4711
R11026 VGND.n123 VGND.n122 24.4711
R11027 VGND.n88 VGND.n67 24.4711
R11028 VGND.n129 VGND.n128 24.4711
R11029 VGND.n156 VGND.n135 24.4711
R11030 VGND.n498 VGND.n474 24.4711
R11031 VGND.n2279 VGND.n2253 24.4711
R11032 VGND.n534 VGND.n505 24.4711
R11033 VGND.n509 VGND.n508 24.4711
R11034 VGND.n2216 VGND.n2215 24.4711
R11035 VGND.n2223 VGND.n541 24.4711
R11036 VGND.n164 VGND.n136 23.7181
R11037 VGND.n2993 VGND.n2972 23.7181
R11038 VGND.n3010 VGND.n9 23.7181
R11039 VGND.n3010 VGND.n10 23.7181
R11040 VGND.n2966 VGND.n2945 23.7181
R11041 VGND.n65 VGND.n35 23.7181
R11042 VGND.n1155 VGND.n1153 23.7181
R11043 VGND.n1127 VGND.n1105 23.7181
R11044 VGND.n1127 VGND.n1126 23.7181
R11045 VGND.n2283 VGND.n2252 23.7181
R11046 VGND.n2210 VGND.n545 23.7181
R11047 VGND.n2247 VGND.n542 23.7181
R11048 VGND.n1385 VGND.n1356 23.7181
R11049 VGND.n1385 VGND.n1357 23.7181
R11050 VGND.n2997 VGND.n2972 23.7181
R11051 VGND.n117 VGND.n115 23.3417
R11052 VGND.n117 VGND.n92 23.3417
R11053 VGND.n2211 VGND.n2210 23.3417
R11054 VGND.n1143 VGND.n1140 21.4593
R11055 VGND.n1116 VGND.n1112 21.4593
R11056 VGND.n2236 VGND.n2235 21.4593
R11057 VGND.n1374 VGND.n1373 21.4593
R11058 VGND.n179 VGND.n178 21.0905
R11059 VGND.n102 VGND.n101 21.0905
R11060 VGND.n80 VGND.n79 21.0905
R11061 VGND.n148 VGND.n147 21.0905
R11062 VGND.n180 VGND.n179 20.3299
R11063 VGND.n103 VGND.n102 20.3299
R11064 VGND.n81 VGND.n80 20.3299
R11065 VGND.n149 VGND.n148 20.3299
R11066 VGND.n494 VGND.n479 19.9534
R11067 VGND.n2275 VGND.n2260 19.9534
R11068 VGND.n530 VGND.n515 19.9534
R11069 VGND.n3006 VGND.n3005 19.2005
R11070 VGND.n61 VGND.n60 19.2005
R11071 VGND.n2223 VGND.n2222 19.2005
R11072 VGND.n1361 VGND.n1360 19.2005
R11073 VGND.t734 VGND.t939 16.8587
R11074 VGND.t1063 VGND.t941 16.8587
R11075 VGND.t2504 VGND.t1215 16.8587
R11076 VGND.t124 VGND.t1213 16.8587
R11077 VGND.n1133 VGND.n1132 16.077
R11078 VGND.n3000 VGND.n2999 16.077
R11079 VGND.n60 VGND.n59 15.4358
R11080 VGND.n2222 VGND.n2221 15.4358
R11081 VGND.n3005 VGND.n3004 14.6829
R11082 VGND.n160 VGND.n159 14.6829
R11083 VGND.n2255 VGND.n2254 14.6829
R11084 VGND.n1360 VGND.n1359 14.6829
R11085 VGND.n483 VGND.n482 14.5711
R11086 VGND.n2264 VGND.n2263 14.5711
R11087 VGND.n519 VGND.n518 14.5711
R11088 VGND.n2194 VGND.n2193 14.5711
R11089 VGND.n133 VGND.n68 14.3064
R11090 VGND.n538 VGND.n506 14.3064
R11091 VGND.n490 VGND.n489 13.9299
R11092 VGND.n2271 VGND.n2270 13.9299
R11093 VGND.n526 VGND.n525 13.9299
R11094 VGND.n2199 VGND.n2191 13.9299
R11095 VGND.n65 VGND.n36 13.5534
R11096 VGND.n2247 VGND.n541 13.5534
R11097 VGND.n193 VGND.n166 13.177
R11098 VGND.n133 VGND.n67 13.177
R11099 VGND.n164 VGND.n135 13.177
R11100 VGND.n502 VGND.n474 13.177
R11101 VGND.n2283 VGND.n2253 13.177
R11102 VGND.n538 VGND.n505 13.177
R11103 VGND.n193 VGND.n167 12.8005
R11104 VGND.n502 VGND.n475 12.8005
R11105 VGND.n3023 VGND.t2691 12.5645
R11106 VGND.n1132 VGND.n1131 10.5417
R11107 VGND.n2999 VGND.n2998 10.5417
R11108 VGND.n3004 VGND.n3003 10.0534
R11109 VGND.n1359 VGND.n1358 10.0534
R11110 VGND.n20 VGND.n19 9.3005
R11111 VGND.n21 VGND.n13 9.3005
R11112 VGND.n24 VGND.n23 9.3005
R11113 VGND.n25 VGND.n12 9.3005
R11114 VGND.n27 VGND.n26 9.3005
R11115 VGND.n28 VGND.n11 9.3005
R11116 VGND.n30 VGND.n29 9.3005
R11117 VGND.n31 VGND.n9 9.3005
R11118 VGND.n3008 VGND.n10 9.3005
R11119 VGND.n3007 VGND.n3006 9.3005
R11120 VGND.n3010 VGND.n3009 9.3005
R11121 VGND.n191 VGND.n167 9.3005
R11122 VGND.n180 VGND.n174 9.3005
R11123 VGND.n182 VGND.n181 9.3005
R11124 VGND.n184 VGND.n183 9.3005
R11125 VGND.n185 VGND.n168 9.3005
R11126 VGND.n188 VGND.n187 9.3005
R11127 VGND.n189 VGND.n166 9.3005
R11128 VGND.n193 VGND.n192 9.3005
R11129 VGND.n2953 VGND.n2952 9.3005
R11130 VGND.n2954 VGND.n2948 9.3005
R11131 VGND.n2957 VGND.n2956 9.3005
R11132 VGND.n2958 VGND.n2947 9.3005
R11133 VGND.n2960 VGND.n2959 9.3005
R11134 VGND.n2961 VGND.n2946 9.3005
R11135 VGND.n2963 VGND.n2962 9.3005
R11136 VGND.n2964 VGND.n2945 9.3005
R11137 VGND.n2966 VGND.n2965 9.3005
R11138 VGND.n59 VGND.n58 9.3005
R11139 VGND.n46 VGND.n45 9.3005
R11140 VGND.n47 VGND.n39 9.3005
R11141 VGND.n50 VGND.n49 9.3005
R11142 VGND.n51 VGND.n38 9.3005
R11143 VGND.n53 VGND.n52 9.3005
R11144 VGND.n54 VGND.n37 9.3005
R11145 VGND.n56 VGND.n55 9.3005
R11146 VGND.n57 VGND.n35 9.3005
R11147 VGND.n63 VGND.n36 9.3005
R11148 VGND.n62 VGND.n61 9.3005
R11149 VGND.n65 VGND.n64 9.3005
R11150 VGND.n124 VGND.n123 9.3005
R11151 VGND.n103 VGND.n99 9.3005
R11152 VGND.n106 VGND.n105 9.3005
R11153 VGND.n108 VGND.n107 9.3005
R11154 VGND.n109 VGND.n94 9.3005
R11155 VGND.n112 VGND.n111 9.3005
R11156 VGND.n114 VGND.n113 9.3005
R11157 VGND.n120 VGND.n119 9.3005
R11158 VGND.n122 VGND.n91 9.3005
R11159 VGND.n118 VGND.n117 9.3005
R11160 VGND.n128 VGND.n127 9.3005
R11161 VGND.n81 VGND.n75 9.3005
R11162 VGND.n83 VGND.n82 9.3005
R11163 VGND.n85 VGND.n84 9.3005
R11164 VGND.n86 VGND.n69 9.3005
R11165 VGND.n89 VGND.n88 9.3005
R11166 VGND.n90 VGND.n67 9.3005
R11167 VGND.n131 VGND.n68 9.3005
R11168 VGND.n130 VGND.n129 9.3005
R11169 VGND.n133 VGND.n132 9.3005
R11170 VGND.n162 VGND.n136 9.3005
R11171 VGND.n149 VGND.n143 9.3005
R11172 VGND.n151 VGND.n150 9.3005
R11173 VGND.n153 VGND.n152 9.3005
R11174 VGND.n154 VGND.n137 9.3005
R11175 VGND.n157 VGND.n156 9.3005
R11176 VGND.n158 VGND.n135 9.3005
R11177 VGND.n164 VGND.n163 9.3005
R11178 VGND.n1144 VGND.n1143 9.3005
R11179 VGND.n1145 VGND.n1137 9.3005
R11180 VGND.n1147 VGND.n1146 9.3005
R11181 VGND.n1148 VGND.n1136 9.3005
R11182 VGND.n1150 VGND.n1149 9.3005
R11183 VGND.n1151 VGND.n1135 9.3005
R11184 VGND.n1153 VGND.n1152 9.3005
R11185 VGND.n1156 VGND.n1155 9.3005
R11186 VGND.n1117 VGND.n1116 9.3005
R11187 VGND.n1118 VGND.n1108 9.3005
R11188 VGND.n1120 VGND.n1119 9.3005
R11189 VGND.n1121 VGND.n1107 9.3005
R11190 VGND.n1123 VGND.n1122 9.3005
R11191 VGND.n1124 VGND.n1106 9.3005
R11192 VGND.n1126 VGND.n1125 9.3005
R11193 VGND.n1129 VGND.n1105 9.3005
R11194 VGND.n1131 VGND.n1130 9.3005
R11195 VGND.n1128 VGND.n1127 9.3005
R11196 VGND.n500 VGND.n474 9.3005
R11197 VGND.n484 VGND.n481 9.3005
R11198 VGND.n486 VGND.n485 9.3005
R11199 VGND.n490 VGND.n480 9.3005
R11200 VGND.n492 VGND.n491 9.3005
R11201 VGND.n494 VGND.n493 9.3005
R11202 VGND.n497 VGND.n476 9.3005
R11203 VGND.n499 VGND.n498 9.3005
R11204 VGND.n502 VGND.n501 9.3005
R11205 VGND.n2281 VGND.n2253 9.3005
R11206 VGND.n2265 VGND.n2262 9.3005
R11207 VGND.n2267 VGND.n2266 9.3005
R11208 VGND.n2271 VGND.n2261 9.3005
R11209 VGND.n2273 VGND.n2272 9.3005
R11210 VGND.n2275 VGND.n2274 9.3005
R11211 VGND.n2278 VGND.n2257 9.3005
R11212 VGND.n2280 VGND.n2279 9.3005
R11213 VGND.n2256 VGND.n2252 9.3005
R11214 VGND.n2283 VGND.n2282 9.3005
R11215 VGND.n508 VGND.n507 9.3005
R11216 VGND.n511 VGND.n506 9.3005
R11217 VGND.n536 VGND.n505 9.3005
R11218 VGND.n520 VGND.n517 9.3005
R11219 VGND.n522 VGND.n521 9.3005
R11220 VGND.n526 VGND.n516 9.3005
R11221 VGND.n528 VGND.n527 9.3005
R11222 VGND.n530 VGND.n529 9.3005
R11223 VGND.n533 VGND.n512 9.3005
R11224 VGND.n535 VGND.n534 9.3005
R11225 VGND.n510 VGND.n509 9.3005
R11226 VGND.n538 VGND.n537 9.3005
R11227 VGND.n2217 VGND.n2216 9.3005
R11228 VGND.n2208 VGND.n545 9.3005
R11229 VGND.n2195 VGND.n2192 9.3005
R11230 VGND.n2197 VGND.n2196 9.3005
R11231 VGND.n2199 VGND.n2198 9.3005
R11232 VGND.n2201 VGND.n2200 9.3005
R11233 VGND.n2203 VGND.n2202 9.3005
R11234 VGND.n2204 VGND.n2183 9.3005
R11235 VGND.n2207 VGND.n2206 9.3005
R11236 VGND.n2213 VGND.n2212 9.3005
R11237 VGND.n2215 VGND.n2214 9.3005
R11238 VGND.n2210 VGND.n2209 9.3005
R11239 VGND.n2235 VGND.n2228 9.3005
R11240 VGND.n2238 VGND.n2237 9.3005
R11241 VGND.n2239 VGND.n2227 9.3005
R11242 VGND.n2241 VGND.n2240 9.3005
R11243 VGND.n2242 VGND.n2226 9.3005
R11244 VGND.n2244 VGND.n2243 9.3005
R11245 VGND.n2245 VGND.n542 9.3005
R11246 VGND.n2225 VGND.n541 9.3005
R11247 VGND.n2224 VGND.n2223 9.3005
R11248 VGND.n2221 VGND.n2220 9.3005
R11249 VGND.n2247 VGND.n2246 9.3005
R11250 VGND.n1373 VGND.n1366 9.3005
R11251 VGND.n1376 VGND.n1375 9.3005
R11252 VGND.n1377 VGND.n1365 9.3005
R11253 VGND.n1379 VGND.n1378 9.3005
R11254 VGND.n1380 VGND.n1364 9.3005
R11255 VGND.n1382 VGND.n1381 9.3005
R11256 VGND.n1383 VGND.n1357 9.3005
R11257 VGND.n1363 VGND.n1356 9.3005
R11258 VGND.n1362 VGND.n1361 9.3005
R11259 VGND.n1385 VGND.n1384 9.3005
R11260 VGND.n2982 VGND.n2978 9.3005
R11261 VGND.n2984 VGND.n2983 9.3005
R11262 VGND.n2986 VGND.n2975 9.3005
R11263 VGND.n2988 VGND.n2987 9.3005
R11264 VGND.n2989 VGND.n2974 9.3005
R11265 VGND.n2991 VGND.n2990 9.3005
R11266 VGND.n2992 VGND.n2973 9.3005
R11267 VGND.n2994 VGND.n2993 9.3005
R11268 VGND.n2995 VGND.n2972 9.3005
R11269 VGND.n2997 VGND.n2996 9.3005
R11270 VGND.n2998 VGND.n34 9.3005
R11271 VGND.n181 VGND.n173 8.28285
R11272 VGND.n82 VGND.n74 8.28285
R11273 VGND.n150 VGND.n142 8.28285
R11274 VGND.n2636 VGND.n2635 7.9105
R11275 VGND.n2693 VGND.n337 7.9105
R11276 VGND.n2692 VGND.n338 7.9105
R11277 VGND.n2687 VGND.n343 7.9105
R11278 VGND.n2686 VGND.n344 7.9105
R11279 VGND.n2681 VGND.n349 7.9105
R11280 VGND.n2680 VGND.n350 7.9105
R11281 VGND.n2675 VGND.n2674 7.9105
R11282 VGND.n2712 VGND.n2711 7.9105
R11283 VGND.n2721 VGND.n2720 7.9105
R11284 VGND.n2745 VGND.n2744 7.9105
R11285 VGND.n2759 VGND.n2758 7.9105
R11286 VGND.n2783 VGND.n288 7.9105
R11287 VGND.n2785 VGND.n2784 7.9105
R11288 VGND.n2794 VGND.n2793 7.9105
R11289 VGND.n2937 VGND.n2936 7.9105
R11290 VGND.n2559 VGND.n401 7.9105
R11291 VGND.n2558 VGND.n402 7.9105
R11292 VGND.n2557 VGND.n403 7.9105
R11293 VGND.n2556 VGND.n404 7.9105
R11294 VGND.n2555 VGND.n405 7.9105
R11295 VGND.n2554 VGND.n406 7.9105
R11296 VGND.n2553 VGND.n407 7.9105
R11297 VGND.n2552 VGND.n408 7.9105
R11298 VGND.n2551 VGND.n409 7.9105
R11299 VGND.n2550 VGND.n410 7.9105
R11300 VGND.n2549 VGND.n411 7.9105
R11301 VGND.n2548 VGND.n412 7.9105
R11302 VGND.n2547 VGND.n2546 7.9105
R11303 VGND.n2798 VGND.n282 7.9105
R11304 VGND.n2797 VGND.n283 7.9105
R11305 VGND.n2534 VGND.n2533 7.9105
R11306 VGND.n2357 VGND.n2356 7.9105
R11307 VGND.n2374 VGND.n2373 7.9105
R11308 VGND.n2383 VGND.n2382 7.9105
R11309 VGND.n2400 VGND.n2399 7.9105
R11310 VGND.n2409 VGND.n2408 7.9105
R11311 VGND.n2426 VGND.n2425 7.9105
R11312 VGND.n2435 VGND.n2434 7.9105
R11313 VGND.n2452 VGND.n2451 7.9105
R11314 VGND.n2461 VGND.n2460 7.9105
R11315 VGND.n2478 VGND.n2477 7.9105
R11316 VGND.n2487 VGND.n2486 7.9105
R11317 VGND.n2509 VGND.n2508 7.9105
R11318 VGND.n2802 VGND.n279 7.9105
R11319 VGND.n2801 VGND.n280 7.9105
R11320 VGND.n420 VGND.n419 7.9105
R11321 VGND.n2530 VGND.n2529 7.9105
R11322 VGND.n2361 VGND.n2360 7.9105
R11323 VGND.n2370 VGND.n2369 7.9105
R11324 VGND.n2387 VGND.n2386 7.9105
R11325 VGND.n2396 VGND.n2395 7.9105
R11326 VGND.n2413 VGND.n2412 7.9105
R11327 VGND.n2422 VGND.n2421 7.9105
R11328 VGND.n2439 VGND.n2438 7.9105
R11329 VGND.n2448 VGND.n2447 7.9105
R11330 VGND.n2465 VGND.n2464 7.9105
R11331 VGND.n2474 VGND.n2473 7.9105
R11332 VGND.n2491 VGND.n2490 7.9105
R11333 VGND.n2505 VGND.n2504 7.9105
R11334 VGND.n2805 VGND.n277 7.9105
R11335 VGND.n2807 VGND.n2806 7.9105
R11336 VGND.n2819 VGND.n273 7.9105
R11337 VGND.n2818 VGND.n2817 7.9105
R11338 VGND.n1908 VGND.n1907 7.9105
R11339 VGND.n1917 VGND.n1916 7.9105
R11340 VGND.n1919 VGND.n1918 7.9105
R11341 VGND.n1928 VGND.n1927 7.9105
R11342 VGND.n1930 VGND.n1929 7.9105
R11343 VGND.n1939 VGND.n1938 7.9105
R11344 VGND.n1941 VGND.n1940 7.9105
R11345 VGND.n1950 VGND.n1949 7.9105
R11346 VGND.n1952 VGND.n1951 7.9105
R11347 VGND.n1961 VGND.n1960 7.9105
R11348 VGND.n1963 VGND.n1962 7.9105
R11349 VGND.n1972 VGND.n1971 7.9105
R11350 VGND.n1974 VGND.n1973 7.9105
R11351 VGND.n2823 VGND.n270 7.9105
R11352 VGND.n2822 VGND.n271 7.9105
R11353 VGND.n1990 VGND.n1989 7.9105
R11354 VGND.n2063 VGND.n591 7.9105
R11355 VGND.n2062 VGND.n2061 7.9105
R11356 VGND.n2167 VGND.n556 7.9105
R11357 VGND.n2166 VGND.n557 7.9105
R11358 VGND.n2159 VGND.n562 7.9105
R11359 VGND.n2158 VGND.n563 7.9105
R11360 VGND.n2151 VGND.n568 7.9105
R11361 VGND.n2150 VGND.n569 7.9105
R11362 VGND.n2143 VGND.n574 7.9105
R11363 VGND.n2142 VGND.n575 7.9105
R11364 VGND.n2135 VGND.n580 7.9105
R11365 VGND.n2134 VGND.n581 7.9105
R11366 VGND.n2827 VGND.n267 7.9105
R11367 VGND.n2826 VGND.n268 7.9105
R11368 VGND.n1999 VGND.n1998 7.9105
R11369 VGND.n1997 VGND.n1996 7.9105
R11370 VGND.n2067 VGND.n2066 7.9105
R11371 VGND.n2171 VGND.n553 7.9105
R11372 VGND.n2170 VGND.n554 7.9105
R11373 VGND.n2163 VGND.n559 7.9105
R11374 VGND.n2162 VGND.n560 7.9105
R11375 VGND.n2155 VGND.n565 7.9105
R11376 VGND.n2154 VGND.n566 7.9105
R11377 VGND.n2147 VGND.n571 7.9105
R11378 VGND.n2146 VGND.n572 7.9105
R11379 VGND.n2139 VGND.n577 7.9105
R11380 VGND.n2138 VGND.n578 7.9105
R11381 VGND.n2131 VGND.n2130 7.9105
R11382 VGND.n2830 VGND.n265 7.9105
R11383 VGND.n2832 VGND.n2831 7.9105
R11384 VGND.n2844 VGND.n261 7.9105
R11385 VGND.n2843 VGND.n2842 7.9105
R11386 VGND.n1901 VGND.n548 7.9105
R11387 VGND.n2175 VGND.n2174 7.9105
R11388 VGND.n1759 VGND.n1758 7.9105
R11389 VGND.n1768 VGND.n1767 7.9105
R11390 VGND.n1770 VGND.n1769 7.9105
R11391 VGND.n1779 VGND.n1778 7.9105
R11392 VGND.n1781 VGND.n1780 7.9105
R11393 VGND.n1790 VGND.n1789 7.9105
R11394 VGND.n1792 VGND.n1791 7.9105
R11395 VGND.n1801 VGND.n1800 7.9105
R11396 VGND.n1803 VGND.n1802 7.9105
R11397 VGND.n1812 VGND.n1811 7.9105
R11398 VGND.n1814 VGND.n1813 7.9105
R11399 VGND.n2848 VGND.n258 7.9105
R11400 VGND.n2847 VGND.n259 7.9105
R11401 VGND.n1830 VGND.n1829 7.9105
R11402 VGND.n1899 VGND.n629 7.9105
R11403 VGND.n1685 VGND.n1684 7.9105
R11404 VGND.n1687 VGND.n1686 7.9105
R11405 VGND.n1884 VGND.n643 7.9105
R11406 VGND.n1883 VGND.n644 7.9105
R11407 VGND.n1876 VGND.n649 7.9105
R11408 VGND.n1875 VGND.n650 7.9105
R11409 VGND.n1868 VGND.n655 7.9105
R11410 VGND.n1867 VGND.n656 7.9105
R11411 VGND.n1860 VGND.n661 7.9105
R11412 VGND.n1859 VGND.n662 7.9105
R11413 VGND.n1852 VGND.n1851 7.9105
R11414 VGND.n2852 VGND.n255 7.9105
R11415 VGND.n2851 VGND.n256 7.9105
R11416 VGND.n1839 VGND.n1838 7.9105
R11417 VGND.n1837 VGND.n1836 7.9105
R11418 VGND.n1896 VGND.n633 7.9105
R11419 VGND.n1895 VGND.n634 7.9105
R11420 VGND.n1888 VGND.n640 7.9105
R11421 VGND.n1887 VGND.n641 7.9105
R11422 VGND.n1880 VGND.n646 7.9105
R11423 VGND.n1879 VGND.n647 7.9105
R11424 VGND.n1872 VGND.n652 7.9105
R11425 VGND.n1871 VGND.n653 7.9105
R11426 VGND.n1864 VGND.n658 7.9105
R11427 VGND.n1863 VGND.n659 7.9105
R11428 VGND.n1856 VGND.n664 7.9105
R11429 VGND.n1855 VGND.n730 7.9105
R11430 VGND.n2855 VGND.n253 7.9105
R11431 VGND.n2857 VGND.n2856 7.9105
R11432 VGND.n2869 VGND.n249 7.9105
R11433 VGND.n2868 VGND.n2867 7.9105
R11434 VGND.n1350 VGND.n1349 7.9105
R11435 VGND.n1892 VGND.n636 7.9105
R11436 VGND.n1891 VGND.n637 7.9105
R11437 VGND.n868 VGND.n867 7.9105
R11438 VGND.n866 VGND.n812 7.9105
R11439 VGND.n865 VGND.n813 7.9105
R11440 VGND.n864 VGND.n814 7.9105
R11441 VGND.n863 VGND.n815 7.9105
R11442 VGND.n862 VGND.n816 7.9105
R11443 VGND.n861 VGND.n817 7.9105
R11444 VGND.n860 VGND.n859 7.9105
R11445 VGND.n1669 VGND.n732 7.9105
R11446 VGND.n1668 VGND.n1667 7.9105
R11447 VGND.n2873 VGND.n246 7.9105
R11448 VGND.n2872 VGND.n247 7.9105
R11449 VGND.n1655 VGND.n1654 7.9105
R11450 VGND.n1404 VGND.n801 7.9105
R11451 VGND.n1403 VGND.n802 7.9105
R11452 VGND.n1402 VGND.n1401 7.9105
R11453 VGND.n1488 VGND.n1487 7.9105
R11454 VGND.n1497 VGND.n1496 7.9105
R11455 VGND.n1514 VGND.n1513 7.9105
R11456 VGND.n1523 VGND.n1522 7.9105
R11457 VGND.n1540 VGND.n1539 7.9105
R11458 VGND.n1560 VGND.n758 7.9105
R11459 VGND.n1559 VGND.n1558 7.9105
R11460 VGND.n1628 VGND.n742 7.9105
R11461 VGND.n1630 VGND.n1629 7.9105
R11462 VGND.n2877 VGND.n243 7.9105
R11463 VGND.n2876 VGND.n244 7.9105
R11464 VGND.n741 VGND.n740 7.9105
R11465 VGND.n1651 VGND.n1650 7.9105
R11466 VGND.n1408 VGND.n1407 7.9105
R11467 VGND.n1417 VGND.n1416 7.9105
R11468 VGND.n1475 VGND.n1474 7.9105
R11469 VGND.n1484 VGND.n1483 7.9105
R11470 VGND.n1501 VGND.n1500 7.9105
R11471 VGND.n1510 VGND.n1509 7.9105
R11472 VGND.n1527 VGND.n1526 7.9105
R11473 VGND.n1536 VGND.n1535 7.9105
R11474 VGND.n1564 VGND.n1563 7.9105
R11475 VGND.n1588 VGND.n1587 7.9105
R11476 VGND.n1625 VGND.n744 7.9105
R11477 VGND.n1624 VGND.n745 7.9105
R11478 VGND.n2880 VGND.n240 7.9105
R11479 VGND.n2882 VGND.n2881 7.9105
R11480 VGND.n2894 VGND.n236 7.9105
R11481 VGND.n2893 VGND.n2892 7.9105
R11482 VGND.n1344 VGND.n1343 7.9105
R11483 VGND.n1421 VGND.n1420 7.9105
R11484 VGND.n1471 VGND.n783 7.9105
R11485 VGND.n1470 VGND.n784 7.9105
R11486 VGND.n1469 VGND.n785 7.9105
R11487 VGND.n1468 VGND.n786 7.9105
R11488 VGND.n1467 VGND.n787 7.9105
R11489 VGND.n1466 VGND.n788 7.9105
R11490 VGND.n1465 VGND.n1464 7.9105
R11491 VGND.n1591 VGND.n751 7.9105
R11492 VGND.n1593 VGND.n1592 7.9105
R11493 VGND.n1621 VGND.n747 7.9105
R11494 VGND.n1620 VGND.n1619 7.9105
R11495 VGND.n2898 VGND.n231 7.9105
R11496 VGND.n2897 VGND.n232 7.9105
R11497 VGND.n1607 VGND.n1606 7.9105
R11498 VGND.n1103 VGND.n1025 7.9105
R11499 VGND.n1102 VGND.n1026 7.9105
R11500 VGND.n1101 VGND.n1100 7.9105
R11501 VGND.n1321 VGND.n899 7.9105
R11502 VGND.n1320 VGND.n900 7.9105
R11503 VGND.n1313 VGND.n905 7.9105
R11504 VGND.n1312 VGND.n906 7.9105
R11505 VGND.n1305 VGND.n911 7.9105
R11506 VGND.n1304 VGND.n912 7.9105
R11507 VGND.n1068 VGND.n1067 7.9105
R11508 VGND.n1066 VGND.n1045 7.9105
R11509 VGND.n1065 VGND.n1046 7.9105
R11510 VGND.n1064 VGND.n1063 7.9105
R11511 VGND.n2902 VGND.n2901 7.9105
R11512 VGND.n233 VGND.n228 7.9105
R11513 VGND.n2913 VGND.n2912 7.9105
R11514 VGND.n1161 VGND.n888 7.9105
R11515 VGND.n1331 VGND.n1330 7.9105
R11516 VGND.n1325 VGND.n896 7.9105
R11517 VGND.n1324 VGND.n897 7.9105
R11518 VGND.n1317 VGND.n902 7.9105
R11519 VGND.n1316 VGND.n903 7.9105
R11520 VGND.n1309 VGND.n908 7.9105
R11521 VGND.n1308 VGND.n909 7.9105
R11522 VGND.n1301 VGND.n914 7.9105
R11523 VGND.n1300 VGND.n915 7.9105
R11524 VGND.n1295 VGND.n919 7.9105
R11525 VGND.n1294 VGND.n920 7.9105
R11526 VGND.n1289 VGND.n924 7.9105
R11527 VGND.n1288 VGND.n925 7.9105
R11528 VGND.n1287 VGND.n992 7.9105
R11529 VGND.n2917 VGND.n2916 7.9105
R11530 VGND.n489 VGND.n486 7.90638
R11531 VGND.n482 VGND.n481 7.90638
R11532 VGND.n2270 VGND.n2267 7.90638
R11533 VGND.n2263 VGND.n2262 7.90638
R11534 VGND.n525 VGND.n522 7.90638
R11535 VGND.n518 VGND.n517 7.90638
R11536 VGND.n2196 VGND.n2191 7.90638
R11537 VGND.n2195 VGND.n2194 7.90638
R11538 VGND.n1142 VGND.n1138 7.4049
R11539 VGND.n1115 VGND.n1109 7.4049
R11540 VGND.n2234 VGND.n2232 7.4049
R11541 VGND.n1372 VGND.n1370 7.4049
R11542 VGND VGND.n475 7.12482
R11543 VGND.n178 VGND.n177 6.85473
R11544 VGND.n79 VGND.n78 6.85473
R11545 VGND.n147 VGND.n146 6.85473
R11546 VGND.n2986 VGND.n2985 6.77697
R11547 VGND.n23 VGND.n22 6.77697
R11548 VGND.n2956 VGND.n2955 6.77697
R11549 VGND.n49 VGND.n48 6.77697
R11550 VGND.n3022 VGND.n3021 6.4005
R11551 VGND.n104 VGND.n98 5.27109
R11552 VGND.n2189 VGND.n2188 5.27109
R11553 VGND.n2565 VGND.n2564 4.5005
R11554 VGND.n2568 VGND.n2567 4.5005
R11555 VGND.n2571 VGND.n2570 4.5005
R11556 VGND.n2574 VGND.n2573 4.5005
R11557 VGND.n2577 VGND.n2576 4.5005
R11558 VGND.n2580 VGND.n2579 4.5005
R11559 VGND.n2583 VGND.n2582 4.5005
R11560 VGND.n2586 VGND.n2585 4.5005
R11561 VGND.n2589 VGND.n2588 4.5005
R11562 VGND.n2592 VGND.n2591 4.5005
R11563 VGND.n2595 VGND.n2594 4.5005
R11564 VGND.n2598 VGND.n2597 4.5005
R11565 VGND.n2601 VGND.n2600 4.5005
R11566 VGND.n2604 VGND.n2603 4.5005
R11567 VGND.n2607 VGND.n2606 4.5005
R11568 VGND.n335 VGND.n334 4.5005
R11569 VGND.n2627 VGND.n2626 4.5005
R11570 VGND.n2624 VGND.n2623 4.5005
R11571 VGND.n2621 VGND.n2620 4.5005
R11572 VGND.n2618 VGND.n2617 4.5005
R11573 VGND.n2615 VGND.n2614 4.5005
R11574 VGND.n2612 VGND.n2611 4.5005
R11575 VGND.n323 VGND.n322 4.5005
R11576 VGND.n316 VGND.n315 4.5005
R11577 VGND.n307 VGND.n306 4.5005
R11578 VGND.n2763 VGND.n299 4.5005
R11579 VGND.n2766 VGND.n2765 4.5005
R11580 VGND.n291 VGND.n290 4.5005
R11581 VGND.n2770 VGND.n297 4.5005
R11582 VGND.n205 VGND.n204 4.5005
R11583 VGND.n2631 VGND.n2630 4.5005
R11584 VGND.n2632 VGND.n331 4.5005
R11585 VGND.n2697 VGND.n2696 4.5005
R11586 VGND.n358 VGND.n340 4.5005
R11587 VGND.n365 VGND.n341 4.5005
R11588 VGND.n354 VGND.n346 4.5005
R11589 VGND.n376 VGND.n347 4.5005
R11590 VGND.n353 VGND.n352 4.5005
R11591 VGND.n390 VGND.n389 4.5005
R11592 VGND.n2708 VGND.n2707 4.5005
R11593 VGND.n2725 VGND.n2724 4.5005
R11594 VGND.n2741 VGND.n2740 4.5005
R11595 VGND.n2762 VGND.n300 4.5005
R11596 VGND.n2733 VGND.n289 4.5005
R11597 VGND.n2779 VGND.n2778 4.5005
R11598 VGND.n2772 VGND.n2771 4.5005
R11599 VGND.n2942 VGND.n2941 4.5005
R11600 VGND.n1019 VGND.n1018 4.5005
R11601 VGND.n1016 VGND.n1015 4.5005
R11602 VGND.n1181 VGND.n1180 4.5005
R11603 VGND.n1193 VGND.n1006 4.5005
R11604 VGND.n1200 VGND.n1004 4.5005
R11605 VGND.n1197 VGND.n1195 4.5005
R11606 VGND.n1213 VGND.n1212 4.5005
R11607 VGND.n1251 VGND.n1000 4.5005
R11608 VGND.n1254 VGND.n1253 4.5005
R11609 VGND.n1257 VGND.n1256 4.5005
R11610 VGND.n1260 VGND.n1259 4.5005
R11611 VGND.n1263 VGND.n1262 4.5005
R11612 VGND.n1269 VGND.n998 4.5005
R11613 VGND.n1266 VGND.n1265 4.5005
R11614 VGND.n995 VGND.n994 4.5005
R11615 VGND.n1022 VGND.n1021 4.5005
R11616 VGND.n1165 VGND.n1164 4.5005
R11617 VGND.n1170 VGND.n891 4.5005
R11618 VGND.n1011 VGND.n892 4.5005
R11619 VGND.n1183 VGND.n1182 4.5005
R11620 VGND.n1192 VGND.n1191 4.5005
R11621 VGND.n1202 VGND.n1201 4.5005
R11622 VGND.n1196 VGND.n1003 4.5005
R11623 VGND.n1215 VGND.n1214 4.5005
R11624 VGND.n1250 VGND.n1249 4.5005
R11625 VGND.n1223 VGND.n916 4.5005
R11626 VGND.n1242 VGND.n917 4.5005
R11627 VGND.n1228 VGND.n921 4.5005
R11628 VGND.n1235 VGND.n922 4.5005
R11629 VGND.n1272 VGND.n1271 4.5005
R11630 VGND.n997 VGND.n993 4.5005
R11631 VGND.n1283 VGND.n1282 4.5005
R11632 VGND.n1157 VGND.n1156 4.41365
R11633 VGND VGND.n33 4.35375
R11634 VGND.n1134 VGND.n1133 4.05427
R11635 VGND.n507 VGND.n0 4.05427
R11636 VGND.n2218 VGND.n2217 4.05427
R11637 VGND.n2220 VGND.n2219 4.05427
R11638 VGND.n1358 VGND.n543 4.05427
R11639 VGND VGND.n3002 3.99438
R11640 VGND VGND.n32 3.99438
R11641 VGND.n125 VGND 3.99438
R11642 VGND VGND.n126 3.99438
R11643 VGND.n3001 VGND 3.99437
R11644 VGND.n1284 VGND.n223 3.77268
R11645 VGND.n2940 VGND.n206 3.77268
R11646 VGND.n1163 VGND.n1162 3.77268
R11647 VGND.n2634 VGND.n2633 3.77268
R11648 VGND.n1327 VGND.n1326 3.77268
R11649 VGND.n2691 VGND.n2690 3.77268
R11650 VGND.n1323 VGND.n898 3.77268
R11651 VGND.n2689 VGND.n2688 3.77268
R11652 VGND.n1318 VGND.n901 3.77268
R11653 VGND.n2685 VGND.n2684 3.77268
R11654 VGND.n1315 VGND.n904 3.77268
R11655 VGND.n2683 VGND.n2682 3.77268
R11656 VGND.n1310 VGND.n907 3.77268
R11657 VGND.n2679 VGND.n2678 3.77268
R11658 VGND.n1307 VGND.n910 3.77268
R11659 VGND.n2677 VGND.n2676 3.77268
R11660 VGND.n1302 VGND.n913 3.77268
R11661 VGND.n2710 VGND.n2709 3.77268
R11662 VGND.n1299 VGND.n1298 3.77268
R11663 VGND.n2723 VGND.n2722 3.77268
R11664 VGND.n1297 VGND.n1296 3.77268
R11665 VGND.n2743 VGND.n2742 3.77268
R11666 VGND.n1293 VGND.n1292 3.77268
R11667 VGND.n2761 VGND.n2760 3.77268
R11668 VGND.n1291 VGND.n1290 3.77268
R11669 VGND.n2782 VGND.n2781 3.77268
R11670 VGND.n1270 VGND.n229 3.77268
R11671 VGND.n2780 VGND.n281 3.77268
R11672 VGND.n1286 VGND.n1285 3.77268
R11673 VGND.n2795 VGND.n284 3.77268
R11674 VGND.n1329 VGND.n1328 3.77268
R11675 VGND.n2695 VGND.n2694 3.77268
R11676 VGND.n2769 VGND.n205 3.75914
R11677 VGND.n2631 VGND.n2629 3.75914
R11678 VGND.n1267 VGND.n995 3.75914
R11679 VGND.n1022 VGND.n1020 3.75914
R11680 VGND.n2771 VGND.n284 3.4105
R11681 VGND.n2780 VGND.n2779 3.4105
R11682 VGND.n2781 VGND.n289 3.4105
R11683 VGND.n2762 VGND.n2761 3.4105
R11684 VGND.n2742 VGND.n2741 3.4105
R11685 VGND.n2724 VGND.n2723 3.4105
R11686 VGND.n2709 VGND.n2708 3.4105
R11687 VGND.n2677 VGND.n390 3.4105
R11688 VGND.n2678 VGND.n352 3.4105
R11689 VGND.n2683 VGND.n347 3.4105
R11690 VGND.n2684 VGND.n346 3.4105
R11691 VGND.n2689 VGND.n341 3.4105
R11692 VGND.n2690 VGND.n340 3.4105
R11693 VGND.n2696 VGND.n2695 3.4105
R11694 VGND.n2941 VGND.n2940 3.4105
R11695 VGND.n2770 VGND.n2769 3.4105
R11696 VGND.n2768 VGND.n291 3.4105
R11697 VGND.n2767 VGND.n2766 3.4105
R11698 VGND.n2764 VGND.n2763 3.4105
R11699 VGND.n307 VGND.n298 3.4105
R11700 VGND.n2609 VGND.n316 3.4105
R11701 VGND.n2610 VGND.n323 3.4105
R11702 VGND.n2613 VGND.n2612 3.4105
R11703 VGND.n2616 VGND.n2615 3.4105
R11704 VGND.n2619 VGND.n2618 3.4105
R11705 VGND.n2622 VGND.n2621 3.4105
R11706 VGND.n2625 VGND.n2624 3.4105
R11707 VGND.n2628 VGND.n2627 3.4105
R11708 VGND.n2629 VGND.n335 3.4105
R11709 VGND.n2633 VGND.n2632 3.4105
R11710 VGND.n2937 VGND.n206 3.4105
R11711 VGND.n2635 VGND.n2634 3.4105
R11712 VGND.n2559 VGND.n397 3.4105
R11713 VGND.n2533 VGND.n2532 3.4105
R11714 VGND.n2557 VGND.n339 3.4105
R11715 VGND.n2692 VGND.n2691 3.4105
R11716 VGND.n2384 VGND.n2383 3.4105
R11717 VGND.n2358 VGND.n2357 3.4105
R11718 VGND.n2531 VGND.n2530 3.4105
R11719 VGND.n2399 VGND.n2398 3.4105
R11720 VGND.n2556 VGND.n342 3.4105
R11721 VGND.n2688 VGND.n2687 3.4105
R11722 VGND.n2397 VGND.n2396 3.4105
R11723 VGND.n2386 VGND.n2385 3.4105
R11724 VGND.n2360 VGND.n2359 3.4105
R11725 VGND.n2818 VGND.n274 3.4105
R11726 VGND.n2412 VGND.n2411 3.4105
R11727 VGND.n2410 VGND.n2409 3.4105
R11728 VGND.n2555 VGND.n345 3.4105
R11729 VGND.n2686 VGND.n2685 3.4105
R11730 VGND.n1929 VGND.n449 3.4105
R11731 VGND.n1928 VGND.n453 3.4105
R11732 VGND.n1918 VGND.n457 3.4105
R11733 VGND.n1907 VGND.n467 3.4105
R11734 VGND.n1990 VGND.n604 3.4105
R11735 VGND.n1939 VGND.n445 3.4105
R11736 VGND.n2423 VGND.n2422 3.4105
R11737 VGND.n2425 VGND.n2424 3.4105
R11738 VGND.n2554 VGND.n348 3.4105
R11739 VGND.n2682 VGND.n2681 3.4105
R11740 VGND.n2158 VGND.n2157 3.4105
R11741 VGND.n2160 VGND.n2159 3.4105
R11742 VGND.n2166 VGND.n2165 3.4105
R11743 VGND.n2168 VGND.n2167 3.4105
R11744 VGND.n2064 VGND.n2063 3.4105
R11745 VGND.n1997 VGND.n603 3.4105
R11746 VGND.n2152 VGND.n2151 3.4105
R11747 VGND.n1940 VGND.n441 3.4105
R11748 VGND.n2438 VGND.n2437 3.4105
R11749 VGND.n2436 VGND.n2435 3.4105
R11750 VGND.n2553 VGND.n351 3.4105
R11751 VGND.n2680 VGND.n2679 3.4105
R11752 VGND.n2154 VGND.n2153 3.4105
R11753 VGND.n2156 VGND.n2155 3.4105
R11754 VGND.n2162 VGND.n2161 3.4105
R11755 VGND.n2164 VGND.n2163 3.4105
R11756 VGND.n2170 VGND.n2169 3.4105
R11757 VGND.n2066 VGND.n2065 3.4105
R11758 VGND.n2843 VGND.n262 3.4105
R11759 VGND.n2148 VGND.n2147 3.4105
R11760 VGND.n2150 VGND.n2149 3.4105
R11761 VGND.n1950 VGND.n437 3.4105
R11762 VGND.n2449 VGND.n2448 3.4105
R11763 VGND.n2451 VGND.n2450 3.4105
R11764 VGND.n2552 VGND.n391 3.4105
R11765 VGND.n2676 VGND.n2675 3.4105
R11766 VGND.n1790 VGND.n570 3.4105
R11767 VGND.n1780 VGND.n567 3.4105
R11768 VGND.n1779 VGND.n564 3.4105
R11769 VGND.n1769 VGND.n561 3.4105
R11770 VGND.n1768 VGND.n558 3.4105
R11771 VGND.n1758 VGND.n555 3.4105
R11772 VGND.n1901 VGND.n588 3.4105
R11773 VGND.n1830 VGND.n1737 3.4105
R11774 VGND.n1791 VGND.n573 3.4105
R11775 VGND.n2146 VGND.n2145 3.4105
R11776 VGND.n2144 VGND.n2143 3.4105
R11777 VGND.n1951 VGND.n433 3.4105
R11778 VGND.n2464 VGND.n2463 3.4105
R11779 VGND.n2462 VGND.n2461 3.4105
R11780 VGND.n2551 VGND.n321 3.4105
R11781 VGND.n2711 VGND.n2710 3.4105
R11782 VGND.n1867 VGND.n1866 3.4105
R11783 VGND.n1869 VGND.n1868 3.4105
R11784 VGND.n1875 VGND.n1874 3.4105
R11785 VGND.n1877 VGND.n1876 3.4105
R11786 VGND.n1883 VGND.n1882 3.4105
R11787 VGND.n1885 VGND.n1884 3.4105
R11788 VGND.n1686 VGND.n639 3.4105
R11789 VGND.n1899 VGND.n1898 3.4105
R11790 VGND.n1837 VGND.n1736 3.4105
R11791 VGND.n1861 VGND.n1860 3.4105
R11792 VGND.n1801 VGND.n576 3.4105
R11793 VGND.n2140 VGND.n2139 3.4105
R11794 VGND.n2142 VGND.n2141 3.4105
R11795 VGND.n1961 VGND.n429 3.4105
R11796 VGND.n2475 VGND.n2474 3.4105
R11797 VGND.n2477 VGND.n2476 3.4105
R11798 VGND.n2550 VGND.n317 3.4105
R11799 VGND.n2722 VGND.n2721 3.4105
R11800 VGND.n1863 VGND.n1862 3.4105
R11801 VGND.n1865 VGND.n1864 3.4105
R11802 VGND.n1871 VGND.n1870 3.4105
R11803 VGND.n1873 VGND.n1872 3.4105
R11804 VGND.n1879 VGND.n1878 3.4105
R11805 VGND.n1881 VGND.n1880 3.4105
R11806 VGND.n1887 VGND.n1886 3.4105
R11807 VGND.n1889 VGND.n1888 3.4105
R11808 VGND.n1897 VGND.n1896 3.4105
R11809 VGND.n2868 VGND.n250 3.4105
R11810 VGND.n1857 VGND.n1856 3.4105
R11811 VGND.n1859 VGND.n1858 3.4105
R11812 VGND.n1802 VGND.n579 3.4105
R11813 VGND.n2138 VGND.n2137 3.4105
R11814 VGND.n2136 VGND.n2135 3.4105
R11815 VGND.n1962 VGND.n425 3.4105
R11816 VGND.n2490 VGND.n2489 3.4105
R11817 VGND.n2488 VGND.n2487 3.4105
R11818 VGND.n2549 VGND.n305 3.4105
R11819 VGND.n2744 VGND.n2743 3.4105
R11820 VGND.n860 VGND.n663 3.4105
R11821 VGND.n861 VGND.n660 3.4105
R11822 VGND.n862 VGND.n657 3.4105
R11823 VGND.n863 VGND.n654 3.4105
R11824 VGND.n864 VGND.n651 3.4105
R11825 VGND.n865 VGND.n648 3.4105
R11826 VGND.n866 VGND.n645 3.4105
R11827 VGND.n867 VGND.n642 3.4105
R11828 VGND.n1891 VGND.n1890 3.4105
R11829 VGND.n1349 VGND.n630 3.4105
R11830 VGND.n1654 VGND.n737 3.4105
R11831 VGND.n1670 VGND.n1669 3.4105
R11832 VGND.n1855 VGND.n1854 3.4105
R11833 VGND.n1853 VGND.n1852 3.4105
R11834 VGND.n1812 VGND.n582 3.4105
R11835 VGND.n2132 VGND.n2131 3.4105
R11836 VGND.n2134 VGND.n2133 3.4105
R11837 VGND.n1972 VGND.n421 3.4105
R11838 VGND.n2506 VGND.n2505 3.4105
R11839 VGND.n2508 VGND.n2507 3.4105
R11840 VGND.n2548 VGND.n301 3.4105
R11841 VGND.n2760 VGND.n2759 3.4105
R11842 VGND.n1629 VGND.n731 3.4105
R11843 VGND.n1628 VGND.n1627 3.4105
R11844 VGND.n1559 VGND.n753 3.4105
R11845 VGND.n1561 VGND.n1560 3.4105
R11846 VGND.n1539 VGND.n1538 3.4105
R11847 VGND.n1524 VGND.n1523 3.4105
R11848 VGND.n1513 VGND.n1512 3.4105
R11849 VGND.n1498 VGND.n1497 3.4105
R11850 VGND.n1487 VGND.n1486 3.4105
R11851 VGND.n1402 VGND.n638 3.4105
R11852 VGND.n1405 VGND.n1404 3.4105
R11853 VGND.n1651 VGND.n738 3.4105
R11854 VGND.n2878 VGND.n2877 3.4105
R11855 VGND.n1668 VGND.n242 3.4105
R11856 VGND.n2855 VGND.n2854 3.4105
R11857 VGND.n2853 VGND.n2852 3.4105
R11858 VGND.n1813 VGND.n254 3.4105
R11859 VGND.n2830 VGND.n2829 3.4105
R11860 VGND.n2828 VGND.n2827 3.4105
R11861 VGND.n1973 VGND.n266 3.4105
R11862 VGND.n2805 VGND.n2804 3.4105
R11863 VGND.n2803 VGND.n2802 3.4105
R11864 VGND.n2547 VGND.n278 3.4105
R11865 VGND.n2783 VGND.n2782 3.4105
R11866 VGND.n2880 VGND.n2879 3.4105
R11867 VGND.n1624 VGND.n1623 3.4105
R11868 VGND.n1626 VGND.n1625 3.4105
R11869 VGND.n1589 VGND.n1588 3.4105
R11870 VGND.n1563 VGND.n1562 3.4105
R11871 VGND.n1537 VGND.n1536 3.4105
R11872 VGND.n1526 VGND.n1525 3.4105
R11873 VGND.n1511 VGND.n1510 3.4105
R11874 VGND.n1500 VGND.n1499 3.4105
R11875 VGND.n1485 VGND.n1484 3.4105
R11876 VGND.n1474 VGND.n1473 3.4105
R11877 VGND.n1407 VGND.n1406 3.4105
R11878 VGND.n2893 VGND.n237 3.4105
R11879 VGND.n2881 VGND.n230 3.4105
R11880 VGND.n2876 VGND.n2875 3.4105
R11881 VGND.n2874 VGND.n2873 3.4105
R11882 VGND.n2856 VGND.n245 3.4105
R11883 VGND.n2851 VGND.n2850 3.4105
R11884 VGND.n2849 VGND.n2848 3.4105
R11885 VGND.n2831 VGND.n257 3.4105
R11886 VGND.n2826 VGND.n2825 3.4105
R11887 VGND.n2824 VGND.n2823 3.4105
R11888 VGND.n2806 VGND.n269 3.4105
R11889 VGND.n2801 VGND.n2800 3.4105
R11890 VGND.n2799 VGND.n2798 3.4105
R11891 VGND.n2784 VGND.n281 3.4105
R11892 VGND.n2899 VGND.n2898 3.4105
R11893 VGND.n1620 VGND.n241 3.4105
R11894 VGND.n1622 VGND.n1621 3.4105
R11895 VGND.n1592 VGND.n743 3.4105
R11896 VGND.n1591 VGND.n1590 3.4105
R11897 VGND.n1465 VGND.n757 3.4105
R11898 VGND.n1466 VGND.n762 3.4105
R11899 VGND.n1467 VGND.n766 3.4105
R11900 VGND.n1468 VGND.n770 3.4105
R11901 VGND.n1469 VGND.n774 3.4105
R11902 VGND.n1470 VGND.n778 3.4105
R11903 VGND.n1472 VGND.n1471 3.4105
R11904 VGND.n1344 VGND.n798 3.4105
R11905 VGND.n1606 VGND.n1605 3.4105
R11906 VGND.n2897 VGND.n2896 3.4105
R11907 VGND.n2895 VGND.n2894 3.4105
R11908 VGND.n740 VGND.n235 3.4105
R11909 VGND.n2872 VGND.n2871 3.4105
R11910 VGND.n2870 VGND.n2869 3.4105
R11911 VGND.n1838 VGND.n248 3.4105
R11912 VGND.n2847 VGND.n2846 3.4105
R11913 VGND.n2845 VGND.n2844 3.4105
R11914 VGND.n1998 VGND.n260 3.4105
R11915 VGND.n2822 VGND.n2821 3.4105
R11916 VGND.n2820 VGND.n2819 3.4105
R11917 VGND.n419 VGND.n272 3.4105
R11918 VGND.n2797 VGND.n2796 3.4105
R11919 VGND.n2795 VGND.n2794 3.4105
R11920 VGND.n234 VGND.n233 3.4105
R11921 VGND.n2901 VGND.n2900 3.4105
R11922 VGND.n1064 VGND.n923 3.4105
R11923 VGND.n1065 VGND.n746 3.4105
R11924 VGND.n1066 VGND.n918 3.4105
R11925 VGND.n1067 VGND.n752 3.4105
R11926 VGND.n1304 VGND.n1303 3.4105
R11927 VGND.n1306 VGND.n1305 3.4105
R11928 VGND.n1312 VGND.n1311 3.4105
R11929 VGND.n1314 VGND.n1313 3.4105
R11930 VGND.n1320 VGND.n1319 3.4105
R11931 VGND.n1322 VGND.n1321 3.4105
R11932 VGND.n1101 VGND.n782 3.4105
R11933 VGND.n1104 VGND.n1103 3.4105
R11934 VGND.n2913 VGND.n226 3.4105
R11935 VGND.n1102 VGND.n792 3.4105
R11936 VGND.n1420 VGND.n1419 3.4105
R11937 VGND.n1418 VGND.n1417 3.4105
R11938 VGND.n1403 VGND.n635 3.4105
R11939 VGND.n1893 VGND.n1892 3.4105
R11940 VGND.n1895 VGND.n1894 3.4105
R11941 VGND.n1685 VGND.n551 3.4105
R11942 VGND.n2174 VGND.n2173 3.4105
R11943 VGND.n2172 VGND.n2171 3.4105
R11944 VGND.n2062 VGND.n552 3.4105
R11945 VGND.n1917 VGND.n461 3.4105
R11946 VGND.n2371 VGND.n2370 3.4105
R11947 VGND.n2373 VGND.n2372 3.4105
R11948 VGND.n2558 VGND.n336 3.4105
R11949 VGND.n2694 VGND.n2693 3.4105
R11950 VGND.n1285 VGND.n993 3.4105
R11951 VGND.n1271 VGND.n1270 3.4105
R11952 VGND.n1291 VGND.n922 3.4105
R11953 VGND.n1292 VGND.n921 3.4105
R11954 VGND.n1297 VGND.n917 3.4105
R11955 VGND.n1298 VGND.n916 3.4105
R11956 VGND.n1250 VGND.n913 3.4105
R11957 VGND.n1214 VGND.n910 3.4105
R11958 VGND.n1196 VGND.n907 3.4105
R11959 VGND.n1201 VGND.n904 3.4105
R11960 VGND.n1192 VGND.n901 3.4105
R11961 VGND.n1182 VGND.n898 3.4105
R11962 VGND.n1327 VGND.n892 3.4105
R11963 VGND.n1328 VGND.n891 3.4105
R11964 VGND.n1284 VGND.n1283 3.4105
R11965 VGND.n1267 VGND.n1266 3.4105
R11966 VGND.n1269 VGND.n1268 3.4105
R11967 VGND.n1264 VGND.n1263 3.4105
R11968 VGND.n1261 VGND.n1260 3.4105
R11969 VGND.n1258 VGND.n1257 3.4105
R11970 VGND.n1255 VGND.n1254 3.4105
R11971 VGND.n1252 VGND.n1251 3.4105
R11972 VGND.n1213 VGND.n999 3.4105
R11973 VGND.n1198 VGND.n1197 3.4105
R11974 VGND.n1200 VGND.n1199 3.4105
R11975 VGND.n1194 VGND.n1193 3.4105
R11976 VGND.n1181 VGND.n1005 3.4105
R11977 VGND.n1017 VGND.n1016 3.4105
R11978 VGND.n1020 VGND.n1019 3.4105
R11979 VGND.n1164 VGND.n1163 3.4105
R11980 VGND.n1287 VGND.n1286 3.4105
R11981 VGND.n1288 VGND.n229 3.4105
R11982 VGND.n1290 VGND.n1289 3.4105
R11983 VGND.n1294 VGND.n1293 3.4105
R11984 VGND.n1296 VGND.n1295 3.4105
R11985 VGND.n1300 VGND.n1299 3.4105
R11986 VGND.n1302 VGND.n1301 3.4105
R11987 VGND.n1308 VGND.n1307 3.4105
R11988 VGND.n1310 VGND.n1309 3.4105
R11989 VGND.n1316 VGND.n1315 3.4105
R11990 VGND.n1318 VGND.n1317 3.4105
R11991 VGND.n1324 VGND.n1323 3.4105
R11992 VGND.n1326 VGND.n1325 3.4105
R11993 VGND.n1330 VGND.n1329 3.4105
R11994 VGND.n1162 VGND.n1161 3.4105
R11995 VGND.n2916 VGND.n223 3.4105
R11996 VGND.n105 VGND.n104 3.01226
R11997 VGND.n2200 VGND.n2189 3.01226
R11998 VGND.n2184 VGND.n545 2.63579
R11999 VGND.n2565 VGND 2.52282
R12000 VGND.n2568 VGND 2.52282
R12001 VGND.n2571 VGND 2.52282
R12002 VGND.n2574 VGND 2.52282
R12003 VGND.n2577 VGND 2.52282
R12004 VGND.n2580 VGND 2.52282
R12005 VGND.n2583 VGND 2.52282
R12006 VGND.n2586 VGND 2.52282
R12007 VGND.n2589 VGND 2.52282
R12008 VGND.n2592 VGND 2.52282
R12009 VGND.n2595 VGND 2.52282
R12010 VGND.n2598 VGND 2.52282
R12011 VGND.n2601 VGND 2.52282
R12012 VGND.n2604 VGND 2.52282
R12013 VGND.n2607 VGND 2.52282
R12014 VGND.n186 VGND.n185 2.25932
R12015 VGND.n114 VGND.n93 2.25932
R12016 VGND.n110 VGND.n109 2.25932
R12017 VGND.n87 VGND.n86 2.25932
R12018 VGND.n155 VGND.n154 2.25932
R12019 VGND.n2205 VGND.n2204 2.25932
R12020 VGND.n491 VGND.n479 1.88285
R12021 VGND.n2272 VGND.n2260 1.88285
R12022 VGND.n527 VGND.n515 1.88285
R12023 VGND.n2608 VGND 1.79514
R12024 VGND.n1158 VGND.n224 1.76378
R12025 VGND.n2608 VGND 1.57193
R12026 VGND.n2940 VGND.n2939 1.54254
R12027 VGND.n2938 VGND.n2937 1.54254
R12028 VGND.n2533 VGND.n207 1.54254
R12029 VGND.n2530 VGND.n417 1.54254
R12030 VGND.n2818 VGND.n275 1.54254
R12031 VGND.n1991 VGND.n1990 1.54254
R12032 VGND.n1997 VGND.n1992 1.54254
R12033 VGND.n2843 VGND.n263 1.54254
R12034 VGND.n1831 VGND.n1830 1.54254
R12035 VGND.n1837 VGND.n1832 1.54254
R12036 VGND.n2868 VGND.n251 1.54254
R12037 VGND.n1654 VGND.n1653 1.54254
R12038 VGND.n1652 VGND.n1651 1.54254
R12039 VGND.n2893 VGND.n238 1.54254
R12040 VGND.n1606 VGND.n225 1.54254
R12041 VGND.n2914 VGND.n2913 1.54254
R12042 VGND.n1284 VGND.n224 1.54254
R12043 VGND.n2916 VGND.n2915 1.54254
R12044 VGND.n121 VGND.n120 1.50638
R12045 VGND.n2212 VGND.n544 1.50638
R12046 VGND VGND.n2562 1.3946
R12047 VGND.n2561 VGND 1.3946
R12048 VGND.n2560 VGND 1.3946
R12049 VGND VGND.n398 1.3946
R12050 VGND.n1905 VGND 1.3946
R12051 VGND VGND.n1906 1.3946
R12052 VGND.n1904 VGND 1.3946
R12053 VGND.n1903 VGND 1.3946
R12054 VGND.n1902 VGND 1.3946
R12055 VGND.n1900 VGND 1.3946
R12056 VGND VGND.n626 1.3946
R12057 VGND VGND.n1348 1.3946
R12058 VGND.n1347 VGND 1.3946
R12059 VGND.n1346 VGND 1.3946
R12060 VGND.n1345 VGND 1.3946
R12061 VGND VGND.n880 1.3946
R12062 VGND.n1159 VGND 1.3946
R12063 VGND VGND.n1160 1.3946
R12064 VGND.n1158 VGND.n1157 1.04899
R12065 VGND.n2696 VGND.n335 1.00149
R12066 VGND.n2627 VGND.n340 1.00149
R12067 VGND.n2624 VGND.n341 1.00149
R12068 VGND.n2621 VGND.n346 1.00149
R12069 VGND.n2618 VGND.n347 1.00149
R12070 VGND.n2615 VGND.n352 1.00149
R12071 VGND.n2612 VGND.n390 1.00149
R12072 VGND.n2708 VGND.n323 1.00149
R12073 VGND.n2724 VGND.n316 1.00149
R12074 VGND.n2741 VGND.n307 1.00149
R12075 VGND.n2763 VGND.n2762 1.00149
R12076 VGND.n2766 VGND.n289 1.00149
R12077 VGND.n2779 VGND.n291 1.00149
R12078 VGND.n2771 VGND.n2770 1.00149
R12079 VGND.n2941 VGND.n205 1.00149
R12080 VGND.n1019 VGND.n891 1.00149
R12081 VGND.n1016 VGND.n892 1.00149
R12082 VGND.n1182 VGND.n1181 1.00149
R12083 VGND.n1193 VGND.n1192 1.00149
R12084 VGND.n1201 VGND.n1200 1.00149
R12085 VGND.n1197 VGND.n1196 1.00149
R12086 VGND.n1214 VGND.n1213 1.00149
R12087 VGND.n1251 VGND.n1250 1.00149
R12088 VGND.n1254 VGND.n916 1.00149
R12089 VGND.n1257 VGND.n917 1.00149
R12090 VGND.n1260 VGND.n921 1.00149
R12091 VGND.n1263 VGND.n922 1.00149
R12092 VGND.n1271 VGND.n1269 1.00149
R12093 VGND.n1266 VGND.n993 1.00149
R12094 VGND.n1283 VGND.n995 1.00149
R12095 VGND.n1164 VGND.n1022 1.00149
R12096 VGND.n2632 VGND.n2631 0.973133
R12097 VGND.n2346 VGND.n2 0.9305
R12098 VGND.n178 VGND.n174 0.929432
R12099 VGND.n101 VGND.n99 0.929432
R12100 VGND.n79 VGND.n75 0.929432
R12101 VGND.n147 VGND.n143 0.929432
R12102 VGND.n126 VGND.n1 0.916608
R12103 VGND VGND.n2565 0.839786
R12104 VGND VGND.n2568 0.839786
R12105 VGND VGND.n2571 0.839786
R12106 VGND VGND.n2574 0.839786
R12107 VGND VGND.n2577 0.839786
R12108 VGND VGND.n2580 0.839786
R12109 VGND VGND.n2583 0.839786
R12110 VGND VGND.n2586 0.839786
R12111 VGND VGND.n2589 0.839786
R12112 VGND VGND.n2592 0.839786
R12113 VGND VGND.n2595 0.839786
R12114 VGND VGND.n2598 0.839786
R12115 VGND VGND.n2601 0.839786
R12116 VGND VGND.n2604 0.839786
R12117 VGND VGND.n2607 0.839786
R12118 VGND.n3023 VGND.n3022 0.7755
R12119 VGND.n3024 VGND.n3023 0.774207
R12120 VGND.n2981 VGND.n2978 0.753441
R12121 VGND.n20 VGND.n18 0.753441
R12122 VGND.n2953 VGND.n2951 0.753441
R12123 VGND.n46 VGND.n44 0.753441
R12124 VGND.n159 VGND.n136 0.753441
R12125 VGND.n2254 VGND.n2252 0.753441
R12126 VGND.n3025 VGND 0.706681
R12127 VGND VGND.n0 0.542567
R12128 VGND.n3025 VGND.n1 0.507317
R12129 VGND.n2939 VGND.n33 0.404308
R12130 VGND.n115 VGND.n114 0.376971
R12131 VGND.n120 VGND.n92 0.376971
R12132 VGND.n1140 VGND.n1137 0.376971
R12133 VGND.n1112 VGND.n1108 0.376971
R12134 VGND.n2212 VGND.n2211 0.376971
R12135 VGND.n2237 VGND.n2236 0.376971
R12136 VGND.n1375 VGND.n1374 0.376971
R12137 VGND VGND.n3025 0.37415
R12138 VGND.n226 VGND.n223 0.362676
R12139 VGND.n1605 VGND.n226 0.362676
R12140 VGND.n1605 VGND.n237 0.362676
R12141 VGND.n738 VGND.n237 0.362676
R12142 VGND.n738 VGND.n737 0.362676
R12143 VGND.n737 VGND.n250 0.362676
R12144 VGND.n1736 VGND.n250 0.362676
R12145 VGND.n1737 VGND.n1736 0.362676
R12146 VGND.n1737 VGND.n262 0.362676
R12147 VGND.n603 VGND.n262 0.362676
R12148 VGND.n604 VGND.n603 0.362676
R12149 VGND.n604 VGND.n274 0.362676
R12150 VGND.n2531 VGND.n274 0.362676
R12151 VGND.n2532 VGND.n2531 0.362676
R12152 VGND.n2532 VGND.n206 0.362676
R12153 VGND.n1162 VGND.n1104 0.362676
R12154 VGND.n1104 VGND.n798 0.362676
R12155 VGND.n1406 VGND.n798 0.362676
R12156 VGND.n1406 VGND.n1405 0.362676
R12157 VGND.n1405 VGND.n630 0.362676
R12158 VGND.n1897 VGND.n630 0.362676
R12159 VGND.n1898 VGND.n1897 0.362676
R12160 VGND.n1898 VGND.n588 0.362676
R12161 VGND.n2065 VGND.n588 0.362676
R12162 VGND.n2065 VGND.n2064 0.362676
R12163 VGND.n2064 VGND.n467 0.362676
R12164 VGND.n2359 VGND.n467 0.362676
R12165 VGND.n2359 VGND.n2358 0.362676
R12166 VGND.n2358 VGND.n397 0.362676
R12167 VGND.n2634 VGND.n397 0.362676
R12168 VGND.n1326 VGND.n782 0.362676
R12169 VGND.n1472 VGND.n782 0.362676
R12170 VGND.n1473 VGND.n1472 0.362676
R12171 VGND.n1473 VGND.n638 0.362676
R12172 VGND.n1890 VGND.n638 0.362676
R12173 VGND.n1890 VGND.n1889 0.362676
R12174 VGND.n1889 VGND.n639 0.362676
R12175 VGND.n639 VGND.n555 0.362676
R12176 VGND.n2169 VGND.n555 0.362676
R12177 VGND.n2169 VGND.n2168 0.362676
R12178 VGND.n2168 VGND.n457 0.362676
R12179 VGND.n2385 VGND.n457 0.362676
R12180 VGND.n2385 VGND.n2384 0.362676
R12181 VGND.n2384 VGND.n339 0.362676
R12182 VGND.n2691 VGND.n339 0.362676
R12183 VGND.n1323 VGND.n1322 0.362676
R12184 VGND.n1322 VGND.n778 0.362676
R12185 VGND.n1485 VGND.n778 0.362676
R12186 VGND.n1486 VGND.n1485 0.362676
R12187 VGND.n1486 VGND.n642 0.362676
R12188 VGND.n1886 VGND.n642 0.362676
R12189 VGND.n1886 VGND.n1885 0.362676
R12190 VGND.n1885 VGND.n558 0.362676
R12191 VGND.n2164 VGND.n558 0.362676
R12192 VGND.n2165 VGND.n2164 0.362676
R12193 VGND.n2165 VGND.n453 0.362676
R12194 VGND.n2397 VGND.n453 0.362676
R12195 VGND.n2398 VGND.n2397 0.362676
R12196 VGND.n2398 VGND.n342 0.362676
R12197 VGND.n2688 VGND.n342 0.362676
R12198 VGND.n1319 VGND.n1318 0.362676
R12199 VGND.n1319 VGND.n774 0.362676
R12200 VGND.n1499 VGND.n774 0.362676
R12201 VGND.n1499 VGND.n1498 0.362676
R12202 VGND.n1498 VGND.n645 0.362676
R12203 VGND.n1881 VGND.n645 0.362676
R12204 VGND.n1882 VGND.n1881 0.362676
R12205 VGND.n1882 VGND.n561 0.362676
R12206 VGND.n2161 VGND.n561 0.362676
R12207 VGND.n2161 VGND.n2160 0.362676
R12208 VGND.n2160 VGND.n449 0.362676
R12209 VGND.n2411 VGND.n449 0.362676
R12210 VGND.n2411 VGND.n2410 0.362676
R12211 VGND.n2410 VGND.n345 0.362676
R12212 VGND.n2685 VGND.n345 0.362676
R12213 VGND.n1315 VGND.n1314 0.362676
R12214 VGND.n1314 VGND.n770 0.362676
R12215 VGND.n1511 VGND.n770 0.362676
R12216 VGND.n1512 VGND.n1511 0.362676
R12217 VGND.n1512 VGND.n648 0.362676
R12218 VGND.n1878 VGND.n648 0.362676
R12219 VGND.n1878 VGND.n1877 0.362676
R12220 VGND.n1877 VGND.n564 0.362676
R12221 VGND.n2156 VGND.n564 0.362676
R12222 VGND.n2157 VGND.n2156 0.362676
R12223 VGND.n2157 VGND.n445 0.362676
R12224 VGND.n2423 VGND.n445 0.362676
R12225 VGND.n2424 VGND.n2423 0.362676
R12226 VGND.n2424 VGND.n348 0.362676
R12227 VGND.n2682 VGND.n348 0.362676
R12228 VGND.n1311 VGND.n1310 0.362676
R12229 VGND.n1311 VGND.n766 0.362676
R12230 VGND.n1525 VGND.n766 0.362676
R12231 VGND.n1525 VGND.n1524 0.362676
R12232 VGND.n1524 VGND.n651 0.362676
R12233 VGND.n1873 VGND.n651 0.362676
R12234 VGND.n1874 VGND.n1873 0.362676
R12235 VGND.n1874 VGND.n567 0.362676
R12236 VGND.n2153 VGND.n567 0.362676
R12237 VGND.n2153 VGND.n2152 0.362676
R12238 VGND.n2152 VGND.n441 0.362676
R12239 VGND.n2437 VGND.n441 0.362676
R12240 VGND.n2437 VGND.n2436 0.362676
R12241 VGND.n2436 VGND.n351 0.362676
R12242 VGND.n2679 VGND.n351 0.362676
R12243 VGND.n1307 VGND.n1306 0.362676
R12244 VGND.n1306 VGND.n762 0.362676
R12245 VGND.n1537 VGND.n762 0.362676
R12246 VGND.n1538 VGND.n1537 0.362676
R12247 VGND.n1538 VGND.n654 0.362676
R12248 VGND.n1870 VGND.n654 0.362676
R12249 VGND.n1870 VGND.n1869 0.362676
R12250 VGND.n1869 VGND.n570 0.362676
R12251 VGND.n2148 VGND.n570 0.362676
R12252 VGND.n2149 VGND.n2148 0.362676
R12253 VGND.n2149 VGND.n437 0.362676
R12254 VGND.n2449 VGND.n437 0.362676
R12255 VGND.n2450 VGND.n2449 0.362676
R12256 VGND.n2450 VGND.n391 0.362676
R12257 VGND.n2676 VGND.n391 0.362676
R12258 VGND.n1303 VGND.n1302 0.362676
R12259 VGND.n1303 VGND.n757 0.362676
R12260 VGND.n1562 VGND.n757 0.362676
R12261 VGND.n1562 VGND.n1561 0.362676
R12262 VGND.n1561 VGND.n657 0.362676
R12263 VGND.n1865 VGND.n657 0.362676
R12264 VGND.n1866 VGND.n1865 0.362676
R12265 VGND.n1866 VGND.n573 0.362676
R12266 VGND.n2145 VGND.n573 0.362676
R12267 VGND.n2145 VGND.n2144 0.362676
R12268 VGND.n2144 VGND.n433 0.362676
R12269 VGND.n2463 VGND.n433 0.362676
R12270 VGND.n2463 VGND.n2462 0.362676
R12271 VGND.n2462 VGND.n321 0.362676
R12272 VGND.n2710 VGND.n321 0.362676
R12273 VGND.n1299 VGND.n752 0.362676
R12274 VGND.n1590 VGND.n752 0.362676
R12275 VGND.n1590 VGND.n1589 0.362676
R12276 VGND.n1589 VGND.n753 0.362676
R12277 VGND.n753 VGND.n660 0.362676
R12278 VGND.n1862 VGND.n660 0.362676
R12279 VGND.n1862 VGND.n1861 0.362676
R12280 VGND.n1861 VGND.n576 0.362676
R12281 VGND.n2140 VGND.n576 0.362676
R12282 VGND.n2141 VGND.n2140 0.362676
R12283 VGND.n2141 VGND.n429 0.362676
R12284 VGND.n2475 VGND.n429 0.362676
R12285 VGND.n2476 VGND.n2475 0.362676
R12286 VGND.n2476 VGND.n317 0.362676
R12287 VGND.n2722 VGND.n317 0.362676
R12288 VGND.n1296 VGND.n918 0.362676
R12289 VGND.n918 VGND.n743 0.362676
R12290 VGND.n1626 VGND.n743 0.362676
R12291 VGND.n1627 VGND.n1626 0.362676
R12292 VGND.n1627 VGND.n663 0.362676
R12293 VGND.n1857 VGND.n663 0.362676
R12294 VGND.n1858 VGND.n1857 0.362676
R12295 VGND.n1858 VGND.n579 0.362676
R12296 VGND.n2137 VGND.n579 0.362676
R12297 VGND.n2137 VGND.n2136 0.362676
R12298 VGND.n2136 VGND.n425 0.362676
R12299 VGND.n2489 VGND.n425 0.362676
R12300 VGND.n2489 VGND.n2488 0.362676
R12301 VGND.n2488 VGND.n305 0.362676
R12302 VGND.n2743 VGND.n305 0.362676
R12303 VGND.n1293 VGND.n746 0.362676
R12304 VGND.n1622 VGND.n746 0.362676
R12305 VGND.n1623 VGND.n1622 0.362676
R12306 VGND.n1623 VGND.n731 0.362676
R12307 VGND.n1670 VGND.n731 0.362676
R12308 VGND.n1854 VGND.n1670 0.362676
R12309 VGND.n1854 VGND.n1853 0.362676
R12310 VGND.n1853 VGND.n582 0.362676
R12311 VGND.n2132 VGND.n582 0.362676
R12312 VGND.n2133 VGND.n2132 0.362676
R12313 VGND.n2133 VGND.n421 0.362676
R12314 VGND.n2506 VGND.n421 0.362676
R12315 VGND.n2507 VGND.n2506 0.362676
R12316 VGND.n2507 VGND.n301 0.362676
R12317 VGND.n2760 VGND.n301 0.362676
R12318 VGND.n1290 VGND.n923 0.362676
R12319 VGND.n923 VGND.n241 0.362676
R12320 VGND.n2879 VGND.n241 0.362676
R12321 VGND.n2879 VGND.n2878 0.362676
R12322 VGND.n2878 VGND.n242 0.362676
R12323 VGND.n2854 VGND.n242 0.362676
R12324 VGND.n2854 VGND.n2853 0.362676
R12325 VGND.n2853 VGND.n254 0.362676
R12326 VGND.n2829 VGND.n254 0.362676
R12327 VGND.n2829 VGND.n2828 0.362676
R12328 VGND.n2828 VGND.n266 0.362676
R12329 VGND.n2804 VGND.n266 0.362676
R12330 VGND.n2804 VGND.n2803 0.362676
R12331 VGND.n2803 VGND.n278 0.362676
R12332 VGND.n2782 VGND.n278 0.362676
R12333 VGND.n2900 VGND.n229 0.362676
R12334 VGND.n2900 VGND.n2899 0.362676
R12335 VGND.n2899 VGND.n230 0.362676
R12336 VGND.n2875 VGND.n230 0.362676
R12337 VGND.n2875 VGND.n2874 0.362676
R12338 VGND.n2874 VGND.n245 0.362676
R12339 VGND.n2850 VGND.n245 0.362676
R12340 VGND.n2850 VGND.n2849 0.362676
R12341 VGND.n2849 VGND.n257 0.362676
R12342 VGND.n2825 VGND.n257 0.362676
R12343 VGND.n2825 VGND.n2824 0.362676
R12344 VGND.n2824 VGND.n269 0.362676
R12345 VGND.n2800 VGND.n269 0.362676
R12346 VGND.n2800 VGND.n2799 0.362676
R12347 VGND.n2799 VGND.n281 0.362676
R12348 VGND.n1286 VGND.n234 0.362676
R12349 VGND.n2896 VGND.n234 0.362676
R12350 VGND.n2896 VGND.n2895 0.362676
R12351 VGND.n2895 VGND.n235 0.362676
R12352 VGND.n2871 VGND.n235 0.362676
R12353 VGND.n2871 VGND.n2870 0.362676
R12354 VGND.n2870 VGND.n248 0.362676
R12355 VGND.n2846 VGND.n248 0.362676
R12356 VGND.n2846 VGND.n2845 0.362676
R12357 VGND.n2845 VGND.n260 0.362676
R12358 VGND.n2821 VGND.n260 0.362676
R12359 VGND.n2821 VGND.n2820 0.362676
R12360 VGND.n2820 VGND.n272 0.362676
R12361 VGND.n2796 VGND.n272 0.362676
R12362 VGND.n2796 VGND.n2795 0.362676
R12363 VGND.n1329 VGND.n792 0.362676
R12364 VGND.n1419 VGND.n792 0.362676
R12365 VGND.n1419 VGND.n1418 0.362676
R12366 VGND.n1418 VGND.n635 0.362676
R12367 VGND.n1893 VGND.n635 0.362676
R12368 VGND.n1894 VGND.n1893 0.362676
R12369 VGND.n1894 VGND.n551 0.362676
R12370 VGND.n2173 VGND.n551 0.362676
R12371 VGND.n2173 VGND.n2172 0.362676
R12372 VGND.n2172 VGND.n552 0.362676
R12373 VGND.n552 VGND.n461 0.362676
R12374 VGND.n2371 VGND.n461 0.362676
R12375 VGND.n2372 VGND.n2371 0.362676
R12376 VGND.n2372 VGND.n336 0.362676
R12377 VGND.n2694 VGND.n336 0.362676
R12378 VGND.n2769 VGND.n2768 0.349144
R12379 VGND.n2768 VGND.n2767 0.349144
R12380 VGND.n2767 VGND.n2764 0.349144
R12381 VGND.n2764 VGND.n298 0.349144
R12382 VGND.n2609 VGND.n298 0.349144
R12383 VGND.n2610 VGND.n2609 0.349144
R12384 VGND.n2613 VGND.n2610 0.349144
R12385 VGND.n2616 VGND.n2613 0.349144
R12386 VGND.n2619 VGND.n2616 0.349144
R12387 VGND.n2622 VGND.n2619 0.349144
R12388 VGND.n2625 VGND.n2622 0.349144
R12389 VGND.n2628 VGND.n2625 0.349144
R12390 VGND.n2629 VGND.n2628 0.349144
R12391 VGND.n1268 VGND.n1267 0.349144
R12392 VGND.n1268 VGND.n1264 0.349144
R12393 VGND.n1264 VGND.n1261 0.349144
R12394 VGND.n1261 VGND.n1258 0.349144
R12395 VGND.n1258 VGND.n1255 0.349144
R12396 VGND.n1255 VGND.n1252 0.349144
R12397 VGND.n1252 VGND.n999 0.349144
R12398 VGND.n1198 VGND.n999 0.349144
R12399 VGND.n1199 VGND.n1198 0.349144
R12400 VGND.n1199 VGND.n1194 0.349144
R12401 VGND.n1194 VGND.n1005 0.349144
R12402 VGND.n1017 VGND.n1005 0.349144
R12403 VGND.n1020 VGND.n1017 0.349144
R12404 VGND.n2700 VGND.n331 0.327628
R12405 VGND.n2697 VGND.n333 0.327628
R12406 VGND.n361 VGND.n358 0.327628
R12407 VGND.n369 VGND.n365 0.327628
R12408 VGND.n372 VGND.n354 0.327628
R12409 VGND.n380 VGND.n376 0.327628
R12410 VGND.n383 VGND.n353 0.327628
R12411 VGND.n389 VGND.n388 0.327628
R12412 VGND.n2707 VGND.n2706 0.327628
R12413 VGND.n2727 VGND.n2725 0.327628
R12414 VGND.n2740 VGND.n2739 0.327628
R12415 VGND.n2736 VGND.n300 0.327628
R12416 VGND.n2733 VGND.n2732 0.327628
R12417 VGND.n2778 VGND.n2777 0.327628
R12418 VGND.n2774 VGND.n2772 0.327628
R12419 VGND.n2793 VGND.n2792 0.327628
R12420 VGND.n2789 VGND.n2785 0.327628
R12421 VGND.n2754 VGND.n288 0.327628
R12422 VGND.n2758 VGND.n2757 0.327628
R12423 VGND.n2749 VGND.n2745 0.327628
R12424 VGND.n2720 VGND.n2719 0.327628
R12425 VGND.n2716 VGND.n2712 0.327628
R12426 VGND.n2674 VGND.n2673 0.327628
R12427 VGND.n2670 VGND.n350 0.327628
R12428 VGND.n2665 VGND.n349 0.327628
R12429 VGND.n2660 VGND.n344 0.327628
R12430 VGND.n2655 VGND.n343 0.327628
R12431 VGND.n2650 VGND.n338 0.327628
R12432 VGND.n2645 VGND.n337 0.327628
R12433 VGND.n2640 VGND.n2636 0.327628
R12434 VGND.n2537 VGND.n283 0.327628
R12435 VGND.n2542 VGND.n282 0.327628
R12436 VGND.n2546 VGND.n2545 0.327628
R12437 VGND.n2289 VGND.n412 0.327628
R12438 VGND.n2294 VGND.n411 0.327628
R12439 VGND.n2299 VGND.n410 0.327628
R12440 VGND.n2304 VGND.n409 0.327628
R12441 VGND.n2309 VGND.n408 0.327628
R12442 VGND.n2314 VGND.n407 0.327628
R12443 VGND.n2319 VGND.n406 0.327628
R12444 VGND.n2324 VGND.n405 0.327628
R12445 VGND.n2329 VGND.n404 0.327628
R12446 VGND.n2334 VGND.n403 0.327628
R12447 VGND.n2339 VGND.n402 0.327628
R12448 VGND.n2344 VGND.n401 0.327628
R12449 VGND.n2526 VGND.n420 0.327628
R12450 VGND.n2523 VGND.n280 0.327628
R12451 VGND.n2518 VGND.n279 0.327628
R12452 VGND.n2513 VGND.n2509 0.327628
R12453 VGND.n2486 VGND.n2485 0.327628
R12454 VGND.n2482 VGND.n2478 0.327628
R12455 VGND.n2460 VGND.n2459 0.327628
R12456 VGND.n2456 VGND.n2452 0.327628
R12457 VGND.n2434 VGND.n2433 0.327628
R12458 VGND.n2430 VGND.n2426 0.327628
R12459 VGND.n2408 VGND.n2407 0.327628
R12460 VGND.n2404 VGND.n2400 0.327628
R12461 VGND.n2382 VGND.n2381 0.327628
R12462 VGND.n2378 VGND.n2374 0.327628
R12463 VGND.n2356 VGND.n2355 0.327628
R12464 VGND.n2814 VGND.n273 0.327628
R12465 VGND.n2811 VGND.n2807 0.327628
R12466 VGND.n2500 VGND.n277 0.327628
R12467 VGND.n2504 VGND.n2503 0.327628
R12468 VGND.n2495 VGND.n2491 0.327628
R12469 VGND.n2473 VGND.n2472 0.327628
R12470 VGND.n2469 VGND.n2465 0.327628
R12471 VGND.n2447 VGND.n2446 0.327628
R12472 VGND.n2443 VGND.n2439 0.327628
R12473 VGND.n2421 VGND.n2420 0.327628
R12474 VGND.n2417 VGND.n2413 0.327628
R12475 VGND.n2395 VGND.n2394 0.327628
R12476 VGND.n2391 VGND.n2387 0.327628
R12477 VGND.n2369 VGND.n2368 0.327628
R12478 VGND.n2365 VGND.n2361 0.327628
R12479 VGND.n1986 VGND.n271 0.327628
R12480 VGND.n1983 VGND.n270 0.327628
R12481 VGND.n1978 VGND.n1974 0.327628
R12482 VGND.n1971 VGND.n1970 0.327628
R12483 VGND.n1967 VGND.n1963 0.327628
R12484 VGND.n1960 VGND.n1959 0.327628
R12485 VGND.n1956 VGND.n1952 0.327628
R12486 VGND.n1949 VGND.n1948 0.327628
R12487 VGND.n1945 VGND.n1941 0.327628
R12488 VGND.n1938 VGND.n1937 0.327628
R12489 VGND.n1934 VGND.n1930 0.327628
R12490 VGND.n1927 VGND.n1926 0.327628
R12491 VGND.n1923 VGND.n1919 0.327628
R12492 VGND.n1916 VGND.n1915 0.327628
R12493 VGND.n1912 VGND.n1908 0.327628
R12494 VGND.n1999 VGND.n602 0.327628
R12495 VGND.n2002 VGND.n268 0.327628
R12496 VGND.n2007 VGND.n267 0.327628
R12497 VGND.n2012 VGND.n581 0.327628
R12498 VGND.n2017 VGND.n580 0.327628
R12499 VGND.n2022 VGND.n575 0.327628
R12500 VGND.n2027 VGND.n574 0.327628
R12501 VGND.n2032 VGND.n569 0.327628
R12502 VGND.n2037 VGND.n568 0.327628
R12503 VGND.n2042 VGND.n563 0.327628
R12504 VGND.n2047 VGND.n562 0.327628
R12505 VGND.n2052 VGND.n557 0.327628
R12506 VGND.n2057 VGND.n556 0.327628
R12507 VGND.n2061 VGND.n2060 0.327628
R12508 VGND.n598 VGND.n591 0.327628
R12509 VGND.n2839 VGND.n261 0.327628
R12510 VGND.n2836 VGND.n2832 0.327628
R12511 VGND.n2126 VGND.n265 0.327628
R12512 VGND.n2130 VGND.n2129 0.327628
R12513 VGND.n2121 VGND.n578 0.327628
R12514 VGND.n2116 VGND.n577 0.327628
R12515 VGND.n2111 VGND.n572 0.327628
R12516 VGND.n2106 VGND.n571 0.327628
R12517 VGND.n2101 VGND.n566 0.327628
R12518 VGND.n2096 VGND.n565 0.327628
R12519 VGND.n2091 VGND.n560 0.327628
R12520 VGND.n2086 VGND.n559 0.327628
R12521 VGND.n2081 VGND.n554 0.327628
R12522 VGND.n2076 VGND.n553 0.327628
R12523 VGND.n2071 VGND.n2067 0.327628
R12524 VGND.n1826 VGND.n259 0.327628
R12525 VGND.n1823 VGND.n258 0.327628
R12526 VGND.n1818 VGND.n1814 0.327628
R12527 VGND.n1811 VGND.n1810 0.327628
R12528 VGND.n1807 VGND.n1803 0.327628
R12529 VGND.n1800 VGND.n1799 0.327628
R12530 VGND.n1796 VGND.n1792 0.327628
R12531 VGND.n1789 VGND.n1788 0.327628
R12532 VGND.n1785 VGND.n1781 0.327628
R12533 VGND.n1778 VGND.n1777 0.327628
R12534 VGND.n1774 VGND.n1770 0.327628
R12535 VGND.n1767 VGND.n1766 0.327628
R12536 VGND.n1763 VGND.n1759 0.327628
R12537 VGND.n2175 VGND.n550 0.327628
R12538 VGND.n2178 VGND.n548 0.327628
R12539 VGND.n1839 VGND.n1735 0.327628
R12540 VGND.n1842 VGND.n256 0.327628
R12541 VGND.n1847 VGND.n255 0.327628
R12542 VGND.n1851 VGND.n1850 0.327628
R12543 VGND.n1731 VGND.n662 0.327628
R12544 VGND.n1726 VGND.n661 0.327628
R12545 VGND.n1721 VGND.n656 0.327628
R12546 VGND.n1716 VGND.n655 0.327628
R12547 VGND.n1711 VGND.n650 0.327628
R12548 VGND.n1706 VGND.n649 0.327628
R12549 VGND.n1701 VGND.n644 0.327628
R12550 VGND.n1696 VGND.n643 0.327628
R12551 VGND.n1691 VGND.n1687 0.327628
R12552 VGND.n1684 VGND.n1683 0.327628
R12553 VGND.n1680 VGND.n629 0.327628
R12554 VGND.n2864 VGND.n249 0.327628
R12555 VGND.n2861 VGND.n2857 0.327628
R12556 VGND.n726 VGND.n253 0.327628
R12557 VGND.n730 VGND.n729 0.327628
R12558 VGND.n721 VGND.n664 0.327628
R12559 VGND.n716 VGND.n659 0.327628
R12560 VGND.n711 VGND.n658 0.327628
R12561 VGND.n706 VGND.n653 0.327628
R12562 VGND.n701 VGND.n652 0.327628
R12563 VGND.n696 VGND.n647 0.327628
R12564 VGND.n691 VGND.n646 0.327628
R12565 VGND.n686 VGND.n641 0.327628
R12566 VGND.n681 VGND.n640 0.327628
R12567 VGND.n676 VGND.n634 0.327628
R12568 VGND.n671 VGND.n633 0.327628
R12569 VGND.n1658 VGND.n247 0.327628
R12570 VGND.n1663 VGND.n246 0.327628
R12571 VGND.n1667 VGND.n1666 0.327628
R12572 VGND.n855 VGND.n732 0.327628
R12573 VGND.n859 VGND.n858 0.327628
R12574 VGND.n850 VGND.n817 0.327628
R12575 VGND.n845 VGND.n816 0.327628
R12576 VGND.n840 VGND.n815 0.327628
R12577 VGND.n835 VGND.n814 0.327628
R12578 VGND.n830 VGND.n813 0.327628
R12579 VGND.n825 VGND.n812 0.327628
R12580 VGND.n868 VGND.n808 0.327628
R12581 VGND.n871 VGND.n637 0.327628
R12582 VGND.n876 VGND.n636 0.327628
R12583 VGND.n1354 VGND.n1350 0.327628
R12584 VGND.n1647 VGND.n741 0.327628
R12585 VGND.n1644 VGND.n244 0.327628
R12586 VGND.n1639 VGND.n243 0.327628
R12587 VGND.n1634 VGND.n1630 0.327628
R12588 VGND.n1554 VGND.n742 0.327628
R12589 VGND.n1558 VGND.n1557 0.327628
R12590 VGND.n1549 VGND.n758 0.327628
R12591 VGND.n1544 VGND.n1540 0.327628
R12592 VGND.n1522 VGND.n1521 0.327628
R12593 VGND.n1518 VGND.n1514 0.327628
R12594 VGND.n1496 VGND.n1495 0.327628
R12595 VGND.n1492 VGND.n1488 0.327628
R12596 VGND.n1401 VGND.n1400 0.327628
R12597 VGND.n1397 VGND.n802 0.327628
R12598 VGND.n1392 VGND.n801 0.327628
R12599 VGND.n2889 VGND.n236 0.327628
R12600 VGND.n2886 VGND.n2882 0.327628
R12601 VGND.n1573 VGND.n240 0.327628
R12602 VGND.n1578 VGND.n745 0.327628
R12603 VGND.n1583 VGND.n744 0.327628
R12604 VGND.n1587 VGND.n1586 0.327628
R12605 VGND.n1568 VGND.n1564 0.327628
R12606 VGND.n1535 VGND.n1534 0.327628
R12607 VGND.n1531 VGND.n1527 0.327628
R12608 VGND.n1509 VGND.n1508 0.327628
R12609 VGND.n1505 VGND.n1501 0.327628
R12610 VGND.n1483 VGND.n1482 0.327628
R12611 VGND.n1479 VGND.n1475 0.327628
R12612 VGND.n1416 VGND.n1415 0.327628
R12613 VGND.n1412 VGND.n1408 0.327628
R12614 VGND.n1610 VGND.n232 0.327628
R12615 VGND.n1615 VGND.n231 0.327628
R12616 VGND.n1619 VGND.n1618 0.327628
R12617 VGND.n1602 VGND.n747 0.327628
R12618 VGND.n1597 VGND.n1593 0.327628
R12619 VGND.n1460 VGND.n751 0.327628
R12620 VGND.n1464 VGND.n1463 0.327628
R12621 VGND.n1455 VGND.n788 0.327628
R12622 VGND.n1450 VGND.n787 0.327628
R12623 VGND.n1445 VGND.n786 0.327628
R12624 VGND.n1440 VGND.n785 0.327628
R12625 VGND.n1435 VGND.n784 0.327628
R12626 VGND.n1430 VGND.n783 0.327628
R12627 VGND.n1425 VGND.n1421 0.327628
R12628 VGND.n1343 VGND.n1342 0.327628
R12629 VGND.n2909 VGND.n228 0.327628
R12630 VGND.n2906 VGND.n2902 0.327628
R12631 VGND.n1063 VGND.n1062 0.327628
R12632 VGND.n1059 VGND.n1046 0.327628
R12633 VGND.n1054 VGND.n1045 0.327628
R12634 VGND.n1068 VGND.n1041 0.327628
R12635 VGND.n1071 VGND.n912 0.327628
R12636 VGND.n1076 VGND.n911 0.327628
R12637 VGND.n1081 VGND.n906 0.327628
R12638 VGND.n1086 VGND.n905 0.327628
R12639 VGND.n1091 VGND.n900 0.327628
R12640 VGND.n1096 VGND.n899 0.327628
R12641 VGND.n1100 VGND.n1099 0.327628
R12642 VGND.n1038 VGND.n1026 0.327628
R12643 VGND.n1033 VGND.n1025 0.327628
R12644 VGND.n1167 VGND.n1165 0.327628
R12645 VGND.n1174 VGND.n1170 0.327628
R12646 VGND.n1177 VGND.n1011 0.327628
R12647 VGND.n1187 VGND.n1183 0.327628
R12648 VGND.n1191 VGND.n1190 0.327628
R12649 VGND.n1206 VGND.n1202 0.327628
R12650 VGND.n1209 VGND.n1003 0.327628
R12651 VGND.n1219 VGND.n1215 0.327628
R12652 VGND.n1249 VGND.n1248 0.327628
R12653 VGND.n1245 VGND.n1223 0.327628
R12654 VGND.n1242 VGND.n1241 0.327628
R12655 VGND.n1238 VGND.n1228 0.327628
R12656 VGND.n1235 VGND.n1234 0.327628
R12657 VGND.n1276 VGND.n1272 0.327628
R12658 VGND.n1279 VGND.n997 0.327628
R12659 VGND.n992 VGND.n991 0.327628
R12660 VGND.n988 VGND.n925 0.327628
R12661 VGND.n983 VGND.n924 0.327628
R12662 VGND.n978 VGND.n920 0.327628
R12663 VGND.n973 VGND.n919 0.327628
R12664 VGND.n968 VGND.n915 0.327628
R12665 VGND.n963 VGND.n914 0.327628
R12666 VGND.n958 VGND.n909 0.327628
R12667 VGND.n953 VGND.n908 0.327628
R12668 VGND.n948 VGND.n903 0.327628
R12669 VGND.n943 VGND.n902 0.327628
R12670 VGND.n938 VGND.n897 0.327628
R12671 VGND.n933 VGND.n896 0.327628
R12672 VGND.n1331 VGND.n890 0.327628
R12673 VGND.n1334 VGND.n888 0.327628
R12674 VGND.n126 VGND.n125 0.213567
R12675 VGND.n125 VGND.n32 0.213567
R12676 VGND.n3002 VGND.n32 0.213567
R12677 VGND.n3002 VGND.n3001 0.213567
R12678 VGND.n1157 VGND.n1134 0.213567
R12679 VGND.n1134 VGND.n543 0.213567
R12680 VGND.n2219 VGND.n543 0.213567
R12681 VGND.n2219 VGND.n2218 0.213567
R12682 VGND.n2218 VGND.n0 0.213567
R12683 VGND.n3001 VGND.n33 0.2073
R12684 VGND.n3024 VGND.n2 0.18968
R12685 VGND.n1159 VGND.n1158 0.175967
R12686 VGND.n2633 VGND 0.169807
R12687 VGND.n2695 VGND 0.169807
R12688 VGND.n2690 VGND 0.169807
R12689 VGND.n2689 VGND 0.169807
R12690 VGND.n2684 VGND 0.169807
R12691 VGND.n2683 VGND 0.169807
R12692 VGND.n2678 VGND 0.169807
R12693 VGND.n2677 VGND 0.169807
R12694 VGND.n2709 VGND 0.169807
R12695 VGND.n2723 VGND 0.169807
R12696 VGND.n2742 VGND 0.169807
R12697 VGND.n2761 VGND 0.169807
R12698 VGND.n2781 VGND 0.169807
R12699 VGND.n2780 VGND 0.169807
R12700 VGND.n284 VGND 0.169807
R12701 VGND.n2635 VGND 0.169807
R12702 VGND.n2693 VGND 0.169807
R12703 VGND.n2692 VGND 0.169807
R12704 VGND.n2687 VGND 0.169807
R12705 VGND.n2686 VGND 0.169807
R12706 VGND.n2681 VGND 0.169807
R12707 VGND.n2680 VGND 0.169807
R12708 VGND.n2675 VGND 0.169807
R12709 VGND.n2711 VGND 0.169807
R12710 VGND.n2721 VGND 0.169807
R12711 VGND.n2744 VGND 0.169807
R12712 VGND.n2759 VGND 0.169807
R12713 VGND VGND.n2783 0.169807
R12714 VGND.n2784 VGND 0.169807
R12715 VGND.n2794 VGND 0.169807
R12716 VGND.n2559 VGND 0.169807
R12717 VGND.n2558 VGND 0.169807
R12718 VGND.n2557 VGND 0.169807
R12719 VGND.n2556 VGND 0.169807
R12720 VGND.n2555 VGND 0.169807
R12721 VGND.n2554 VGND 0.169807
R12722 VGND.n2553 VGND 0.169807
R12723 VGND.n2552 VGND 0.169807
R12724 VGND.n2551 VGND 0.169807
R12725 VGND.n2550 VGND 0.169807
R12726 VGND.n2549 VGND 0.169807
R12727 VGND.n2548 VGND 0.169807
R12728 VGND.n2547 VGND 0.169807
R12729 VGND.n2798 VGND 0.169807
R12730 VGND.n2797 VGND 0.169807
R12731 VGND.n2357 VGND 0.169807
R12732 VGND.n2373 VGND 0.169807
R12733 VGND.n2383 VGND 0.169807
R12734 VGND.n2399 VGND 0.169807
R12735 VGND.n2409 VGND 0.169807
R12736 VGND.n2425 VGND 0.169807
R12737 VGND.n2435 VGND 0.169807
R12738 VGND.n2451 VGND 0.169807
R12739 VGND.n2461 VGND 0.169807
R12740 VGND.n2477 VGND 0.169807
R12741 VGND.n2487 VGND 0.169807
R12742 VGND.n2508 VGND 0.169807
R12743 VGND.n2802 VGND 0.169807
R12744 VGND.n2801 VGND 0.169807
R12745 VGND.n419 VGND 0.169807
R12746 VGND.n2360 VGND 0.169807
R12747 VGND.n2370 VGND 0.169807
R12748 VGND.n2386 VGND 0.169807
R12749 VGND.n2396 VGND 0.169807
R12750 VGND.n2412 VGND 0.169807
R12751 VGND.n2422 VGND 0.169807
R12752 VGND.n2438 VGND 0.169807
R12753 VGND.n2448 VGND 0.169807
R12754 VGND.n2464 VGND 0.169807
R12755 VGND.n2474 VGND 0.169807
R12756 VGND.n2490 VGND 0.169807
R12757 VGND.n2505 VGND 0.169807
R12758 VGND VGND.n2805 0.169807
R12759 VGND.n2806 VGND 0.169807
R12760 VGND.n2819 VGND 0.169807
R12761 VGND.n1907 VGND 0.169807
R12762 VGND VGND.n1917 0.169807
R12763 VGND.n1918 VGND 0.169807
R12764 VGND VGND.n1928 0.169807
R12765 VGND.n1929 VGND 0.169807
R12766 VGND VGND.n1939 0.169807
R12767 VGND.n1940 VGND 0.169807
R12768 VGND VGND.n1950 0.169807
R12769 VGND.n1951 VGND 0.169807
R12770 VGND VGND.n1961 0.169807
R12771 VGND.n1962 VGND 0.169807
R12772 VGND VGND.n1972 0.169807
R12773 VGND.n1973 VGND 0.169807
R12774 VGND.n2823 VGND 0.169807
R12775 VGND.n2822 VGND 0.169807
R12776 VGND.n2063 VGND 0.169807
R12777 VGND.n2062 VGND 0.169807
R12778 VGND.n2167 VGND 0.169807
R12779 VGND.n2166 VGND 0.169807
R12780 VGND.n2159 VGND 0.169807
R12781 VGND.n2158 VGND 0.169807
R12782 VGND.n2151 VGND 0.169807
R12783 VGND.n2150 VGND 0.169807
R12784 VGND.n2143 VGND 0.169807
R12785 VGND.n2142 VGND 0.169807
R12786 VGND.n2135 VGND 0.169807
R12787 VGND.n2134 VGND 0.169807
R12788 VGND.n2827 VGND 0.169807
R12789 VGND.n2826 VGND 0.169807
R12790 VGND.n1998 VGND 0.169807
R12791 VGND.n2066 VGND 0.169807
R12792 VGND.n2171 VGND 0.169807
R12793 VGND.n2170 VGND 0.169807
R12794 VGND.n2163 VGND 0.169807
R12795 VGND.n2162 VGND 0.169807
R12796 VGND.n2155 VGND 0.169807
R12797 VGND.n2154 VGND 0.169807
R12798 VGND.n2147 VGND 0.169807
R12799 VGND.n2146 VGND 0.169807
R12800 VGND.n2139 VGND 0.169807
R12801 VGND.n2138 VGND 0.169807
R12802 VGND.n2131 VGND 0.169807
R12803 VGND VGND.n2830 0.169807
R12804 VGND.n2831 VGND 0.169807
R12805 VGND.n2844 VGND 0.169807
R12806 VGND.n1901 VGND 0.169807
R12807 VGND.n2174 VGND 0.169807
R12808 VGND.n1758 VGND 0.169807
R12809 VGND VGND.n1768 0.169807
R12810 VGND.n1769 VGND 0.169807
R12811 VGND VGND.n1779 0.169807
R12812 VGND.n1780 VGND 0.169807
R12813 VGND VGND.n1790 0.169807
R12814 VGND.n1791 VGND 0.169807
R12815 VGND VGND.n1801 0.169807
R12816 VGND.n1802 VGND 0.169807
R12817 VGND VGND.n1812 0.169807
R12818 VGND.n1813 VGND 0.169807
R12819 VGND.n2848 VGND 0.169807
R12820 VGND.n2847 VGND 0.169807
R12821 VGND.n1899 VGND 0.169807
R12822 VGND VGND.n1685 0.169807
R12823 VGND.n1686 VGND 0.169807
R12824 VGND.n1884 VGND 0.169807
R12825 VGND.n1883 VGND 0.169807
R12826 VGND.n1876 VGND 0.169807
R12827 VGND.n1875 VGND 0.169807
R12828 VGND.n1868 VGND 0.169807
R12829 VGND.n1867 VGND 0.169807
R12830 VGND.n1860 VGND 0.169807
R12831 VGND.n1859 VGND 0.169807
R12832 VGND.n1852 VGND 0.169807
R12833 VGND.n2852 VGND 0.169807
R12834 VGND.n2851 VGND 0.169807
R12835 VGND.n1838 VGND 0.169807
R12836 VGND.n1896 VGND 0.169807
R12837 VGND.n1895 VGND 0.169807
R12838 VGND.n1888 VGND 0.169807
R12839 VGND.n1887 VGND 0.169807
R12840 VGND.n1880 VGND 0.169807
R12841 VGND.n1879 VGND 0.169807
R12842 VGND.n1872 VGND 0.169807
R12843 VGND.n1871 VGND 0.169807
R12844 VGND.n1864 VGND 0.169807
R12845 VGND.n1863 VGND 0.169807
R12846 VGND.n1856 VGND 0.169807
R12847 VGND.n1855 VGND 0.169807
R12848 VGND VGND.n2855 0.169807
R12849 VGND.n2856 VGND 0.169807
R12850 VGND.n2869 VGND 0.169807
R12851 VGND.n1349 VGND 0.169807
R12852 VGND.n1892 VGND 0.169807
R12853 VGND.n1891 VGND 0.169807
R12854 VGND.n867 VGND 0.169807
R12855 VGND.n866 VGND 0.169807
R12856 VGND.n865 VGND 0.169807
R12857 VGND.n864 VGND 0.169807
R12858 VGND.n863 VGND 0.169807
R12859 VGND.n862 VGND 0.169807
R12860 VGND.n861 VGND 0.169807
R12861 VGND.n860 VGND 0.169807
R12862 VGND.n1669 VGND 0.169807
R12863 VGND.n1668 VGND 0.169807
R12864 VGND.n2873 VGND 0.169807
R12865 VGND.n2872 VGND 0.169807
R12866 VGND.n1404 VGND 0.169807
R12867 VGND.n1403 VGND 0.169807
R12868 VGND.n1402 VGND 0.169807
R12869 VGND.n1487 VGND 0.169807
R12870 VGND.n1497 VGND 0.169807
R12871 VGND.n1513 VGND 0.169807
R12872 VGND.n1523 VGND 0.169807
R12873 VGND.n1539 VGND 0.169807
R12874 VGND.n1560 VGND 0.169807
R12875 VGND.n1559 VGND 0.169807
R12876 VGND VGND.n1628 0.169807
R12877 VGND.n1629 VGND 0.169807
R12878 VGND.n2877 VGND 0.169807
R12879 VGND.n2876 VGND 0.169807
R12880 VGND.n740 VGND 0.169807
R12881 VGND.n1407 VGND 0.169807
R12882 VGND.n1417 VGND 0.169807
R12883 VGND.n1474 VGND 0.169807
R12884 VGND.n1484 VGND 0.169807
R12885 VGND.n1500 VGND 0.169807
R12886 VGND.n1510 VGND 0.169807
R12887 VGND.n1526 VGND 0.169807
R12888 VGND.n1536 VGND 0.169807
R12889 VGND.n1563 VGND 0.169807
R12890 VGND.n1588 VGND 0.169807
R12891 VGND.n1625 VGND 0.169807
R12892 VGND.n1624 VGND 0.169807
R12893 VGND VGND.n2880 0.169807
R12894 VGND.n2881 VGND 0.169807
R12895 VGND.n2894 VGND 0.169807
R12896 VGND.n1344 VGND 0.169807
R12897 VGND.n1420 VGND 0.169807
R12898 VGND.n1471 VGND 0.169807
R12899 VGND.n1470 VGND 0.169807
R12900 VGND.n1469 VGND 0.169807
R12901 VGND.n1468 VGND 0.169807
R12902 VGND.n1467 VGND 0.169807
R12903 VGND.n1466 VGND 0.169807
R12904 VGND.n1465 VGND 0.169807
R12905 VGND VGND.n1591 0.169807
R12906 VGND.n1592 VGND 0.169807
R12907 VGND.n1621 VGND 0.169807
R12908 VGND.n1620 VGND 0.169807
R12909 VGND.n2898 VGND 0.169807
R12910 VGND.n2897 VGND 0.169807
R12911 VGND.n1103 VGND 0.169807
R12912 VGND.n1102 VGND 0.169807
R12913 VGND.n1101 VGND 0.169807
R12914 VGND.n1321 VGND 0.169807
R12915 VGND.n1320 VGND 0.169807
R12916 VGND.n1313 VGND 0.169807
R12917 VGND.n1312 VGND 0.169807
R12918 VGND.n1305 VGND 0.169807
R12919 VGND.n1304 VGND 0.169807
R12920 VGND.n1067 VGND 0.169807
R12921 VGND.n1066 VGND 0.169807
R12922 VGND.n1065 VGND 0.169807
R12923 VGND.n1064 VGND 0.169807
R12924 VGND.n2901 VGND 0.169807
R12925 VGND.n233 VGND 0.169807
R12926 VGND.n1163 VGND 0.169807
R12927 VGND.n1328 VGND 0.169807
R12928 VGND.n1327 VGND 0.169807
R12929 VGND VGND.n898 0.169807
R12930 VGND VGND.n901 0.169807
R12931 VGND VGND.n904 0.169807
R12932 VGND VGND.n907 0.169807
R12933 VGND VGND.n910 0.169807
R12934 VGND VGND.n913 0.169807
R12935 VGND.n1298 VGND 0.169807
R12936 VGND.n1297 VGND 0.169807
R12937 VGND.n1292 VGND 0.169807
R12938 VGND.n1291 VGND 0.169807
R12939 VGND.n1270 VGND 0.169807
R12940 VGND.n1285 VGND 0.169807
R12941 VGND.n1161 VGND 0.169807
R12942 VGND.n1330 VGND 0.169807
R12943 VGND.n1325 VGND 0.169807
R12944 VGND.n1324 VGND 0.169807
R12945 VGND.n1317 VGND 0.169807
R12946 VGND.n1316 VGND 0.169807
R12947 VGND.n1309 VGND 0.169807
R12948 VGND.n1308 VGND 0.169807
R12949 VGND.n1301 VGND 0.169807
R12950 VGND.n1300 VGND 0.169807
R12951 VGND.n1295 VGND 0.169807
R12952 VGND.n1294 VGND 0.169807
R12953 VGND.n1289 VGND 0.169807
R12954 VGND.n1288 VGND 0.169807
R12955 VGND.n1287 VGND 0.169807
R12956 VGND.n190 VGND 0.159538
R12957 VGND.n161 VGND 0.159538
R12958 VGND.n2915 VGND.n224 0.154425
R12959 VGND.n2915 VGND.n2914 0.154425
R12960 VGND.n2914 VGND.n225 0.154425
R12961 VGND.n238 VGND.n225 0.154425
R12962 VGND.n1652 VGND.n238 0.154425
R12963 VGND.n1653 VGND.n1652 0.154425
R12964 VGND.n1653 VGND.n251 0.154425
R12965 VGND.n1832 VGND.n251 0.154425
R12966 VGND.n1832 VGND.n1831 0.154425
R12967 VGND.n1831 VGND.n263 0.154425
R12968 VGND.n1992 VGND.n263 0.154425
R12969 VGND.n1992 VGND.n1991 0.154425
R12970 VGND.n1991 VGND.n275 0.154425
R12971 VGND.n417 VGND.n275 0.154425
R12972 VGND.n417 VGND.n207 0.154425
R12973 VGND.n2938 VGND.n207 0.154425
R12974 VGND.n2939 VGND.n2938 0.154425
R12975 VGND.n1160 VGND.n1159 0.154425
R12976 VGND.n1160 VGND.n880 0.154425
R12977 VGND.n1345 VGND.n880 0.154425
R12978 VGND.n1346 VGND.n1345 0.154425
R12979 VGND.n1347 VGND.n1346 0.154425
R12980 VGND.n1348 VGND.n1347 0.154425
R12981 VGND.n1348 VGND.n626 0.154425
R12982 VGND.n1900 VGND.n626 0.154425
R12983 VGND.n1902 VGND.n1900 0.154425
R12984 VGND.n1903 VGND.n1902 0.154425
R12985 VGND.n1904 VGND.n1903 0.154425
R12986 VGND.n1906 VGND.n1904 0.154425
R12987 VGND.n1906 VGND.n1905 0.154425
R12988 VGND.n1905 VGND.n398 0.154425
R12989 VGND.n2560 VGND.n398 0.154425
R12990 VGND.n2561 VGND.n2560 0.154425
R12991 VGND.n2562 VGND.n2561 0.154425
R12992 VGND.n1144 VGND.n1138 0.144904
R12993 VGND.n1117 VGND.n1109 0.144904
R12994 VGND.n2232 VGND.n2228 0.144904
R12995 VGND.n1370 VGND.n1366 0.144904
R12996 VGND.n2632 VGND.n2608 0.138284
R12997 VGND.n2700 VGND.n2699 0.13638
R12998 VGND.n355 VGND.n333 0.13638
R12999 VGND.n362 VGND.n361 0.13638
R13000 VGND.n369 VGND.n368 0.13638
R13001 VGND.n373 VGND.n372 0.13638
R13002 VGND.n380 VGND.n379 0.13638
R13003 VGND.n384 VGND.n383 0.13638
R13004 VGND.n388 VGND.n387 0.13638
R13005 VGND.n2706 VGND.n326 0.13638
R13006 VGND.n2727 VGND.n2726 0.13638
R13007 VGND.n2739 VGND.n312 0.13638
R13008 VGND.n2736 VGND.n2735 0.13638
R13009 VGND.n2732 VGND.n2730 0.13638
R13010 VGND.n2777 VGND.n294 0.13638
R13011 VGND.n2774 VGND.n2773 0.13638
R13012 VGND.n2792 VGND.n287 0.13638
R13013 VGND.n2789 VGND.n2788 0.13638
R13014 VGND.n2754 VGND.n2753 0.13638
R13015 VGND.n2757 VGND.n304 0.13638
R13016 VGND.n2749 VGND.n2748 0.13638
R13017 VGND.n2719 VGND.n320 0.13638
R13018 VGND.n2716 VGND.n2715 0.13638
R13019 VGND.n2673 VGND.n394 0.13638
R13020 VGND.n2670 VGND.n2669 0.13638
R13021 VGND.n2665 VGND.n2664 0.13638
R13022 VGND.n2660 VGND.n2659 0.13638
R13023 VGND.n2655 VGND.n2654 0.13638
R13024 VGND.n2650 VGND.n2649 0.13638
R13025 VGND.n2645 VGND.n2644 0.13638
R13026 VGND.n2640 VGND.n2639 0.13638
R13027 VGND.n2537 VGND.n2536 0.13638
R13028 VGND.n2542 VGND.n2541 0.13638
R13029 VGND.n2545 VGND.n415 0.13638
R13030 VGND.n2289 VGND.n2288 0.13638
R13031 VGND.n2294 VGND.n2293 0.13638
R13032 VGND.n2299 VGND.n2298 0.13638
R13033 VGND.n2304 VGND.n2303 0.13638
R13034 VGND.n2309 VGND.n2308 0.13638
R13035 VGND.n2314 VGND.n2313 0.13638
R13036 VGND.n2319 VGND.n2318 0.13638
R13037 VGND.n2324 VGND.n2323 0.13638
R13038 VGND.n2329 VGND.n2328 0.13638
R13039 VGND.n2334 VGND.n2333 0.13638
R13040 VGND.n2339 VGND.n2338 0.13638
R13041 VGND.n2344 VGND.n2343 0.13638
R13042 VGND.n2527 VGND.n2526 0.13638
R13043 VGND.n2523 VGND.n2522 0.13638
R13044 VGND.n2518 VGND.n2517 0.13638
R13045 VGND.n2513 VGND.n2512 0.13638
R13046 VGND.n2485 VGND.n428 0.13638
R13047 VGND.n2482 VGND.n2481 0.13638
R13048 VGND.n2459 VGND.n436 0.13638
R13049 VGND.n2456 VGND.n2455 0.13638
R13050 VGND.n2433 VGND.n444 0.13638
R13051 VGND.n2430 VGND.n2429 0.13638
R13052 VGND.n2407 VGND.n452 0.13638
R13053 VGND.n2404 VGND.n2403 0.13638
R13054 VGND.n2381 VGND.n460 0.13638
R13055 VGND.n2378 VGND.n2377 0.13638
R13056 VGND.n2355 VGND.n472 0.13638
R13057 VGND.n2815 VGND.n2814 0.13638
R13058 VGND.n2811 VGND.n2810 0.13638
R13059 VGND.n2500 VGND.n2499 0.13638
R13060 VGND.n2503 VGND.n424 0.13638
R13061 VGND.n2495 VGND.n2494 0.13638
R13062 VGND.n2472 VGND.n432 0.13638
R13063 VGND.n2469 VGND.n2468 0.13638
R13064 VGND.n2446 VGND.n440 0.13638
R13065 VGND.n2443 VGND.n2442 0.13638
R13066 VGND.n2420 VGND.n448 0.13638
R13067 VGND.n2417 VGND.n2416 0.13638
R13068 VGND.n2394 VGND.n456 0.13638
R13069 VGND.n2391 VGND.n2390 0.13638
R13070 VGND.n2368 VGND.n464 0.13638
R13071 VGND.n2365 VGND.n2364 0.13638
R13072 VGND.n1987 VGND.n1986 0.13638
R13073 VGND.n1983 VGND.n1982 0.13638
R13074 VGND.n1978 VGND.n1977 0.13638
R13075 VGND.n1970 VGND.n608 0.13638
R13076 VGND.n1967 VGND.n1966 0.13638
R13077 VGND.n1959 VGND.n611 0.13638
R13078 VGND.n1956 VGND.n1955 0.13638
R13079 VGND.n1948 VGND.n614 0.13638
R13080 VGND.n1945 VGND.n1944 0.13638
R13081 VGND.n1937 VGND.n617 0.13638
R13082 VGND.n1934 VGND.n1933 0.13638
R13083 VGND.n1926 VGND.n620 0.13638
R13084 VGND.n1923 VGND.n1922 0.13638
R13085 VGND.n1915 VGND.n623 0.13638
R13086 VGND.n1912 VGND.n1911 0.13638
R13087 VGND.n1994 VGND.n602 0.13638
R13088 VGND.n2002 VGND.n2001 0.13638
R13089 VGND.n2007 VGND.n2006 0.13638
R13090 VGND.n2012 VGND.n2011 0.13638
R13091 VGND.n2017 VGND.n2016 0.13638
R13092 VGND.n2022 VGND.n2021 0.13638
R13093 VGND.n2027 VGND.n2026 0.13638
R13094 VGND.n2032 VGND.n2031 0.13638
R13095 VGND.n2037 VGND.n2036 0.13638
R13096 VGND.n2042 VGND.n2041 0.13638
R13097 VGND.n2047 VGND.n2046 0.13638
R13098 VGND.n2052 VGND.n2051 0.13638
R13099 VGND.n2057 VGND.n2056 0.13638
R13100 VGND.n2060 VGND.n594 0.13638
R13101 VGND.n598 VGND.n597 0.13638
R13102 VGND.n2840 VGND.n2839 0.13638
R13103 VGND.n2836 VGND.n2835 0.13638
R13104 VGND.n2126 VGND.n2125 0.13638
R13105 VGND.n2129 VGND.n585 0.13638
R13106 VGND.n2121 VGND.n2120 0.13638
R13107 VGND.n2116 VGND.n2115 0.13638
R13108 VGND.n2111 VGND.n2110 0.13638
R13109 VGND.n2106 VGND.n2105 0.13638
R13110 VGND.n2101 VGND.n2100 0.13638
R13111 VGND.n2096 VGND.n2095 0.13638
R13112 VGND.n2091 VGND.n2090 0.13638
R13113 VGND.n2086 VGND.n2085 0.13638
R13114 VGND.n2081 VGND.n2080 0.13638
R13115 VGND.n2076 VGND.n2075 0.13638
R13116 VGND.n2071 VGND.n2070 0.13638
R13117 VGND.n1827 VGND.n1826 0.13638
R13118 VGND.n1823 VGND.n1822 0.13638
R13119 VGND.n1818 VGND.n1817 0.13638
R13120 VGND.n1810 VGND.n1741 0.13638
R13121 VGND.n1807 VGND.n1806 0.13638
R13122 VGND.n1799 VGND.n1744 0.13638
R13123 VGND.n1796 VGND.n1795 0.13638
R13124 VGND.n1788 VGND.n1747 0.13638
R13125 VGND.n1785 VGND.n1784 0.13638
R13126 VGND.n1777 VGND.n1750 0.13638
R13127 VGND.n1774 VGND.n1773 0.13638
R13128 VGND.n1766 VGND.n1753 0.13638
R13129 VGND.n1763 VGND.n1762 0.13638
R13130 VGND.n1756 VGND.n550 0.13638
R13131 VGND.n2178 VGND.n2177 0.13638
R13132 VGND.n1834 VGND.n1735 0.13638
R13133 VGND.n1842 VGND.n1841 0.13638
R13134 VGND.n1847 VGND.n1846 0.13638
R13135 VGND.n1850 VGND.n1673 0.13638
R13136 VGND.n1731 VGND.n1730 0.13638
R13137 VGND.n1726 VGND.n1725 0.13638
R13138 VGND.n1721 VGND.n1720 0.13638
R13139 VGND.n1716 VGND.n1715 0.13638
R13140 VGND.n1711 VGND.n1710 0.13638
R13141 VGND.n1706 VGND.n1705 0.13638
R13142 VGND.n1701 VGND.n1700 0.13638
R13143 VGND.n1696 VGND.n1695 0.13638
R13144 VGND.n1691 VGND.n1690 0.13638
R13145 VGND.n1683 VGND.n1676 0.13638
R13146 VGND.n1680 VGND.n1679 0.13638
R13147 VGND.n2865 VGND.n2864 0.13638
R13148 VGND.n2861 VGND.n2860 0.13638
R13149 VGND.n726 VGND.n725 0.13638
R13150 VGND.n729 VGND.n667 0.13638
R13151 VGND.n721 VGND.n720 0.13638
R13152 VGND.n716 VGND.n715 0.13638
R13153 VGND.n711 VGND.n710 0.13638
R13154 VGND.n706 VGND.n705 0.13638
R13155 VGND.n701 VGND.n700 0.13638
R13156 VGND.n696 VGND.n695 0.13638
R13157 VGND.n691 VGND.n690 0.13638
R13158 VGND.n686 VGND.n685 0.13638
R13159 VGND.n681 VGND.n680 0.13638
R13160 VGND.n676 VGND.n675 0.13638
R13161 VGND.n671 VGND.n670 0.13638
R13162 VGND.n1658 VGND.n1657 0.13638
R13163 VGND.n1663 VGND.n1662 0.13638
R13164 VGND.n1666 VGND.n735 0.13638
R13165 VGND.n855 VGND.n854 0.13638
R13166 VGND.n858 VGND.n820 0.13638
R13167 VGND.n850 VGND.n849 0.13638
R13168 VGND.n845 VGND.n844 0.13638
R13169 VGND.n840 VGND.n839 0.13638
R13170 VGND.n835 VGND.n834 0.13638
R13171 VGND.n830 VGND.n829 0.13638
R13172 VGND.n825 VGND.n824 0.13638
R13173 VGND.n810 VGND.n808 0.13638
R13174 VGND.n871 VGND.n870 0.13638
R13175 VGND.n876 VGND.n875 0.13638
R13176 VGND.n1354 VGND.n1353 0.13638
R13177 VGND.n1648 VGND.n1647 0.13638
R13178 VGND.n1644 VGND.n1643 0.13638
R13179 VGND.n1639 VGND.n1638 0.13638
R13180 VGND.n1634 VGND.n1633 0.13638
R13181 VGND.n1554 VGND.n1553 0.13638
R13182 VGND.n1557 VGND.n761 0.13638
R13183 VGND.n1549 VGND.n1548 0.13638
R13184 VGND.n1544 VGND.n1543 0.13638
R13185 VGND.n1521 VGND.n769 0.13638
R13186 VGND.n1518 VGND.n1517 0.13638
R13187 VGND.n1495 VGND.n777 0.13638
R13188 VGND.n1492 VGND.n1491 0.13638
R13189 VGND.n1400 VGND.n805 0.13638
R13190 VGND.n1397 VGND.n1396 0.13638
R13191 VGND.n1392 VGND.n1391 0.13638
R13192 VGND.n2890 VGND.n2889 0.13638
R13193 VGND.n2886 VGND.n2885 0.13638
R13194 VGND.n1573 VGND.n1572 0.13638
R13195 VGND.n1578 VGND.n1577 0.13638
R13196 VGND.n1583 VGND.n1582 0.13638
R13197 VGND.n1586 VGND.n756 0.13638
R13198 VGND.n1568 VGND.n1567 0.13638
R13199 VGND.n1534 VGND.n765 0.13638
R13200 VGND.n1531 VGND.n1530 0.13638
R13201 VGND.n1508 VGND.n773 0.13638
R13202 VGND.n1505 VGND.n1504 0.13638
R13203 VGND.n1482 VGND.n781 0.13638
R13204 VGND.n1479 VGND.n1478 0.13638
R13205 VGND.n1415 VGND.n795 0.13638
R13206 VGND.n1412 VGND.n1411 0.13638
R13207 VGND.n1610 VGND.n1609 0.13638
R13208 VGND.n1615 VGND.n1614 0.13638
R13209 VGND.n1618 VGND.n750 0.13638
R13210 VGND.n1602 VGND.n1601 0.13638
R13211 VGND.n1597 VGND.n1596 0.13638
R13212 VGND.n1460 VGND.n1459 0.13638
R13213 VGND.n1463 VGND.n791 0.13638
R13214 VGND.n1455 VGND.n1454 0.13638
R13215 VGND.n1450 VGND.n1449 0.13638
R13216 VGND.n1445 VGND.n1444 0.13638
R13217 VGND.n1440 VGND.n1439 0.13638
R13218 VGND.n1435 VGND.n1434 0.13638
R13219 VGND.n1430 VGND.n1429 0.13638
R13220 VGND.n1425 VGND.n1424 0.13638
R13221 VGND.n1342 VGND.n885 0.13638
R13222 VGND.n2910 VGND.n2909 0.13638
R13223 VGND.n2906 VGND.n2905 0.13638
R13224 VGND.n1062 VGND.n1049 0.13638
R13225 VGND.n1059 VGND.n1058 0.13638
R13226 VGND.n1054 VGND.n1053 0.13638
R13227 VGND.n1043 VGND.n1041 0.13638
R13228 VGND.n1071 VGND.n1070 0.13638
R13229 VGND.n1076 VGND.n1075 0.13638
R13230 VGND.n1081 VGND.n1080 0.13638
R13231 VGND.n1086 VGND.n1085 0.13638
R13232 VGND.n1091 VGND.n1090 0.13638
R13233 VGND.n1096 VGND.n1095 0.13638
R13234 VGND.n1099 VGND.n1029 0.13638
R13235 VGND.n1038 VGND.n1037 0.13638
R13236 VGND.n1033 VGND.n1032 0.13638
R13237 VGND.n1168 VGND.n1167 0.13638
R13238 VGND.n1174 VGND.n1173 0.13638
R13239 VGND.n1178 VGND.n1177 0.13638
R13240 VGND.n1187 VGND.n1186 0.13638
R13241 VGND.n1190 VGND.n1009 0.13638
R13242 VGND.n1206 VGND.n1205 0.13638
R13243 VGND.n1210 VGND.n1209 0.13638
R13244 VGND.n1219 VGND.n1218 0.13638
R13245 VGND.n1248 VGND.n1001 0.13638
R13246 VGND.n1245 VGND.n1244 0.13638
R13247 VGND.n1241 VGND.n1225 0.13638
R13248 VGND.n1238 VGND.n1237 0.13638
R13249 VGND.n1234 VGND.n1232 0.13638
R13250 VGND.n1276 VGND.n1275 0.13638
R13251 VGND.n1280 VGND.n1279 0.13638
R13252 VGND.n991 VGND.n928 0.13638
R13253 VGND.n988 VGND.n987 0.13638
R13254 VGND.n983 VGND.n982 0.13638
R13255 VGND.n978 VGND.n977 0.13638
R13256 VGND.n973 VGND.n972 0.13638
R13257 VGND.n968 VGND.n967 0.13638
R13258 VGND.n963 VGND.n962 0.13638
R13259 VGND.n958 VGND.n957 0.13638
R13260 VGND.n953 VGND.n952 0.13638
R13261 VGND.n948 VGND.n947 0.13638
R13262 VGND.n943 VGND.n942 0.13638
R13263 VGND.n938 VGND.n937 0.13638
R13264 VGND.n933 VGND.n932 0.13638
R13265 VGND.n894 VGND.n890 0.13638
R13266 VGND.n1334 VGND.n1333 0.13638
R13267 VGND VGND.n190 0.120838
R13268 VGND.n19 VGND.n13 0.120292
R13269 VGND.n24 VGND.n13 0.120292
R13270 VGND.n25 VGND.n24 0.120292
R13271 VGND.n26 VGND.n25 0.120292
R13272 VGND.n26 VGND.n11 0.120292
R13273 VGND.n30 VGND.n11 0.120292
R13274 VGND.n31 VGND.n30 0.120292
R13275 VGND.n3008 VGND.n3007 0.120292
R13276 VGND.n3007 VGND.n3003 0.120292
R13277 VGND.n182 VGND.n174 0.120292
R13278 VGND.n183 VGND.n182 0.120292
R13279 VGND.n183 VGND.n168 0.120292
R13280 VGND.n188 VGND.n168 0.120292
R13281 VGND.n189 VGND.n188 0.120292
R13282 VGND.n2952 VGND.n2948 0.120292
R13283 VGND.n2957 VGND.n2948 0.120292
R13284 VGND.n2958 VGND.n2957 0.120292
R13285 VGND.n2959 VGND.n2958 0.120292
R13286 VGND.n2959 VGND.n2946 0.120292
R13287 VGND.n2963 VGND.n2946 0.120292
R13288 VGND.n2964 VGND.n2963 0.120292
R13289 VGND.n45 VGND.n39 0.120292
R13290 VGND.n50 VGND.n39 0.120292
R13291 VGND.n51 VGND.n50 0.120292
R13292 VGND.n52 VGND.n51 0.120292
R13293 VGND.n52 VGND.n37 0.120292
R13294 VGND.n56 VGND.n37 0.120292
R13295 VGND.n57 VGND.n56 0.120292
R13296 VGND.n63 VGND.n62 0.120292
R13297 VGND.n62 VGND.n58 0.120292
R13298 VGND.n106 VGND.n99 0.120292
R13299 VGND.n107 VGND.n106 0.120292
R13300 VGND.n107 VGND.n94 0.120292
R13301 VGND.n112 VGND.n94 0.120292
R13302 VGND.n113 VGND.n112 0.120292
R13303 VGND.n124 VGND.n91 0.120292
R13304 VGND.n83 VGND.n75 0.120292
R13305 VGND.n84 VGND.n83 0.120292
R13306 VGND.n84 VGND.n69 0.120292
R13307 VGND.n89 VGND.n69 0.120292
R13308 VGND.n90 VGND.n89 0.120292
R13309 VGND.n130 VGND.n127 0.120292
R13310 VGND.n151 VGND.n143 0.120292
R13311 VGND.n152 VGND.n151 0.120292
R13312 VGND.n152 VGND.n137 0.120292
R13313 VGND.n157 VGND.n137 0.120292
R13314 VGND.n158 VGND.n157 0.120292
R13315 VGND.n1152 VGND.n1151 0.120292
R13316 VGND.n1151 VGND.n1150 0.120292
R13317 VGND.n1150 VGND.n1136 0.120292
R13318 VGND.n1146 VGND.n1136 0.120292
R13319 VGND.n1146 VGND.n1145 0.120292
R13320 VGND.n1145 VGND.n1144 0.120292
R13321 VGND.n1130 VGND.n1129 0.120292
R13322 VGND.n1125 VGND.n1124 0.120292
R13323 VGND.n1124 VGND.n1123 0.120292
R13324 VGND.n1123 VGND.n1107 0.120292
R13325 VGND.n1119 VGND.n1107 0.120292
R13326 VGND.n1119 VGND.n1118 0.120292
R13327 VGND.n1118 VGND.n1117 0.120292
R13328 VGND.n499 VGND.n476 0.120292
R13329 VGND.n493 VGND.n476 0.120292
R13330 VGND.n493 VGND.n492 0.120292
R13331 VGND.n492 VGND.n480 0.120292
R13332 VGND.n485 VGND.n480 0.120292
R13333 VGND.n485 VGND.n484 0.120292
R13334 VGND.n484 VGND.n483 0.120292
R13335 VGND.n2280 VGND.n2257 0.120292
R13336 VGND.n2274 VGND.n2257 0.120292
R13337 VGND.n2274 VGND.n2273 0.120292
R13338 VGND.n2273 VGND.n2261 0.120292
R13339 VGND.n2266 VGND.n2261 0.120292
R13340 VGND.n2266 VGND.n2265 0.120292
R13341 VGND.n2265 VGND.n2264 0.120292
R13342 VGND.n510 VGND.n507 0.120292
R13343 VGND.n511 VGND.n510 0.120292
R13344 VGND.n535 VGND.n512 0.120292
R13345 VGND.n529 VGND.n512 0.120292
R13346 VGND.n529 VGND.n528 0.120292
R13347 VGND.n528 VGND.n516 0.120292
R13348 VGND.n521 VGND.n516 0.120292
R13349 VGND.n521 VGND.n520 0.120292
R13350 VGND.n520 VGND.n519 0.120292
R13351 VGND.n2214 VGND.n2213 0.120292
R13352 VGND.n2207 VGND.n2183 0.120292
R13353 VGND.n2202 VGND.n2183 0.120292
R13354 VGND.n2202 VGND.n2201 0.120292
R13355 VGND.n2198 VGND.n2197 0.120292
R13356 VGND.n2197 VGND.n2192 0.120292
R13357 VGND.n2193 VGND.n2192 0.120292
R13358 VGND.n2225 VGND.n2224 0.120292
R13359 VGND.n2245 VGND.n2244 0.120292
R13360 VGND.n2244 VGND.n2226 0.120292
R13361 VGND.n2240 VGND.n2226 0.120292
R13362 VGND.n2240 VGND.n2239 0.120292
R13363 VGND.n2239 VGND.n2238 0.120292
R13364 VGND.n2238 VGND.n2228 0.120292
R13365 VGND.n1363 VGND.n1362 0.120292
R13366 VGND.n1383 VGND.n1382 0.120292
R13367 VGND.n1382 VGND.n1364 0.120292
R13368 VGND.n1378 VGND.n1364 0.120292
R13369 VGND.n1378 VGND.n1377 0.120292
R13370 VGND.n1377 VGND.n1376 0.120292
R13371 VGND.n1376 VGND.n1366 0.120292
R13372 VGND.n2983 VGND.n2982 0.120292
R13373 VGND.n2983 VGND.n2975 0.120292
R13374 VGND.n2988 VGND.n2975 0.120292
R13375 VGND.n2989 VGND.n2988 0.120292
R13376 VGND.n2990 VGND.n2989 0.120292
R13377 VGND.n2990 VGND.n2973 0.120292
R13378 VGND.n2994 VGND.n2973 0.120292
R13379 VGND.n2996 VGND.n34 0.120292
R13380 VGND.n3000 VGND.n34 0.120292
R13381 VGND VGND.n161 0.119536
R13382 VGND.n1138 VGND 0.117202
R13383 VGND.n1109 VGND 0.117202
R13384 VGND.n2232 VGND 0.117202
R13385 VGND.n1370 VGND 0.117202
R13386 VGND.n287 VGND.n286 0.110872
R13387 VGND.n2788 VGND.n2787 0.110872
R13388 VGND.n2753 VGND.n2752 0.110872
R13389 VGND.n304 VGND.n303 0.110872
R13390 VGND.n2748 VGND.n2747 0.110872
R13391 VGND.n320 VGND.n319 0.110872
R13392 VGND.n2715 VGND.n2714 0.110872
R13393 VGND.n394 VGND.n393 0.110872
R13394 VGND.n2669 VGND.n2668 0.110872
R13395 VGND.n2664 VGND.n2663 0.110872
R13396 VGND.n2659 VGND.n2658 0.110872
R13397 VGND.n2654 VGND.n2653 0.110872
R13398 VGND.n2649 VGND.n2648 0.110872
R13399 VGND.n2644 VGND.n2643 0.110872
R13400 VGND.n2639 VGND.n2638 0.110872
R13401 VGND.n2536 VGND.n2535 0.110872
R13402 VGND.n2541 VGND.n2540 0.110872
R13403 VGND.n415 VGND.n414 0.110872
R13404 VGND.n2288 VGND.n2287 0.110872
R13405 VGND.n2293 VGND.n2292 0.110872
R13406 VGND.n2298 VGND.n2297 0.110872
R13407 VGND.n2303 VGND.n2302 0.110872
R13408 VGND.n2308 VGND.n2307 0.110872
R13409 VGND.n2313 VGND.n2312 0.110872
R13410 VGND.n2318 VGND.n2317 0.110872
R13411 VGND.n2323 VGND.n2322 0.110872
R13412 VGND.n2328 VGND.n2327 0.110872
R13413 VGND.n2333 VGND.n2332 0.110872
R13414 VGND.n2338 VGND.n2337 0.110872
R13415 VGND.n2343 VGND.n2342 0.110872
R13416 VGND.n2528 VGND.n2527 0.110872
R13417 VGND.n2522 VGND.n2521 0.110872
R13418 VGND.n2517 VGND.n2516 0.110872
R13419 VGND.n2512 VGND.n2511 0.110872
R13420 VGND.n428 VGND.n427 0.110872
R13421 VGND.n2481 VGND.n2480 0.110872
R13422 VGND.n436 VGND.n435 0.110872
R13423 VGND.n2455 VGND.n2454 0.110872
R13424 VGND.n444 VGND.n443 0.110872
R13425 VGND.n2429 VGND.n2428 0.110872
R13426 VGND.n452 VGND.n451 0.110872
R13427 VGND.n2403 VGND.n2402 0.110872
R13428 VGND.n460 VGND.n459 0.110872
R13429 VGND.n2377 VGND.n2376 0.110872
R13430 VGND.n472 VGND.n471 0.110872
R13431 VGND.n2816 VGND.n2815 0.110872
R13432 VGND.n2810 VGND.n2809 0.110872
R13433 VGND.n2499 VGND.n2498 0.110872
R13434 VGND.n424 VGND.n423 0.110872
R13435 VGND.n2494 VGND.n2493 0.110872
R13436 VGND.n432 VGND.n431 0.110872
R13437 VGND.n2468 VGND.n2467 0.110872
R13438 VGND.n440 VGND.n439 0.110872
R13439 VGND.n2442 VGND.n2441 0.110872
R13440 VGND.n448 VGND.n447 0.110872
R13441 VGND.n2416 VGND.n2415 0.110872
R13442 VGND.n456 VGND.n455 0.110872
R13443 VGND.n2390 VGND.n2389 0.110872
R13444 VGND.n464 VGND.n463 0.110872
R13445 VGND.n2364 VGND.n2363 0.110872
R13446 VGND.n1988 VGND.n1987 0.110872
R13447 VGND.n1982 VGND.n1981 0.110872
R13448 VGND.n1977 VGND.n1976 0.110872
R13449 VGND.n608 VGND.n607 0.110872
R13450 VGND.n1966 VGND.n1965 0.110872
R13451 VGND.n611 VGND.n610 0.110872
R13452 VGND.n1955 VGND.n1954 0.110872
R13453 VGND.n614 VGND.n613 0.110872
R13454 VGND.n1944 VGND.n1943 0.110872
R13455 VGND.n617 VGND.n616 0.110872
R13456 VGND.n1933 VGND.n1932 0.110872
R13457 VGND.n620 VGND.n619 0.110872
R13458 VGND.n1922 VGND.n1921 0.110872
R13459 VGND.n623 VGND.n622 0.110872
R13460 VGND.n1911 VGND.n1910 0.110872
R13461 VGND.n1995 VGND.n1994 0.110872
R13462 VGND.n2001 VGND.n2000 0.110872
R13463 VGND.n2006 VGND.n2005 0.110872
R13464 VGND.n2011 VGND.n2010 0.110872
R13465 VGND.n2016 VGND.n2015 0.110872
R13466 VGND.n2021 VGND.n2020 0.110872
R13467 VGND.n2026 VGND.n2025 0.110872
R13468 VGND.n2031 VGND.n2030 0.110872
R13469 VGND.n2036 VGND.n2035 0.110872
R13470 VGND.n2041 VGND.n2040 0.110872
R13471 VGND.n2046 VGND.n2045 0.110872
R13472 VGND.n2051 VGND.n2050 0.110872
R13473 VGND.n2056 VGND.n2055 0.110872
R13474 VGND.n594 VGND.n593 0.110872
R13475 VGND.n597 VGND.n596 0.110872
R13476 VGND.n2841 VGND.n2840 0.110872
R13477 VGND.n2835 VGND.n2834 0.110872
R13478 VGND.n2125 VGND.n2124 0.110872
R13479 VGND.n585 VGND.n584 0.110872
R13480 VGND.n2120 VGND.n2119 0.110872
R13481 VGND.n2115 VGND.n2114 0.110872
R13482 VGND.n2110 VGND.n2109 0.110872
R13483 VGND.n2105 VGND.n2104 0.110872
R13484 VGND.n2100 VGND.n2099 0.110872
R13485 VGND.n2095 VGND.n2094 0.110872
R13486 VGND.n2090 VGND.n2089 0.110872
R13487 VGND.n2085 VGND.n2084 0.110872
R13488 VGND.n2080 VGND.n2079 0.110872
R13489 VGND.n2075 VGND.n2074 0.110872
R13490 VGND.n2070 VGND.n2069 0.110872
R13491 VGND.n1828 VGND.n1827 0.110872
R13492 VGND.n1822 VGND.n1821 0.110872
R13493 VGND.n1817 VGND.n1816 0.110872
R13494 VGND.n1741 VGND.n1740 0.110872
R13495 VGND.n1806 VGND.n1805 0.110872
R13496 VGND.n1744 VGND.n1743 0.110872
R13497 VGND.n1795 VGND.n1794 0.110872
R13498 VGND.n1747 VGND.n1746 0.110872
R13499 VGND.n1784 VGND.n1783 0.110872
R13500 VGND.n1750 VGND.n1749 0.110872
R13501 VGND.n1773 VGND.n1772 0.110872
R13502 VGND.n1753 VGND.n1752 0.110872
R13503 VGND.n1762 VGND.n1761 0.110872
R13504 VGND.n1757 VGND.n1756 0.110872
R13505 VGND.n2177 VGND.n2176 0.110872
R13506 VGND.n1835 VGND.n1834 0.110872
R13507 VGND.n1841 VGND.n1840 0.110872
R13508 VGND.n1846 VGND.n1845 0.110872
R13509 VGND.n1673 VGND.n1672 0.110872
R13510 VGND.n1730 VGND.n1729 0.110872
R13511 VGND.n1725 VGND.n1724 0.110872
R13512 VGND.n1720 VGND.n1719 0.110872
R13513 VGND.n1715 VGND.n1714 0.110872
R13514 VGND.n1710 VGND.n1709 0.110872
R13515 VGND.n1705 VGND.n1704 0.110872
R13516 VGND.n1700 VGND.n1699 0.110872
R13517 VGND.n1695 VGND.n1694 0.110872
R13518 VGND.n1690 VGND.n1689 0.110872
R13519 VGND.n1676 VGND.n1675 0.110872
R13520 VGND.n1679 VGND.n1678 0.110872
R13521 VGND.n2866 VGND.n2865 0.110872
R13522 VGND.n2860 VGND.n2859 0.110872
R13523 VGND.n725 VGND.n724 0.110872
R13524 VGND.n667 VGND.n666 0.110872
R13525 VGND.n720 VGND.n719 0.110872
R13526 VGND.n715 VGND.n714 0.110872
R13527 VGND.n710 VGND.n709 0.110872
R13528 VGND.n705 VGND.n704 0.110872
R13529 VGND.n700 VGND.n699 0.110872
R13530 VGND.n695 VGND.n694 0.110872
R13531 VGND.n690 VGND.n689 0.110872
R13532 VGND.n685 VGND.n684 0.110872
R13533 VGND.n680 VGND.n679 0.110872
R13534 VGND.n675 VGND.n674 0.110872
R13535 VGND.n670 VGND.n669 0.110872
R13536 VGND.n1657 VGND.n1656 0.110872
R13537 VGND.n1662 VGND.n1661 0.110872
R13538 VGND.n735 VGND.n734 0.110872
R13539 VGND.n854 VGND.n853 0.110872
R13540 VGND.n820 VGND.n819 0.110872
R13541 VGND.n849 VGND.n848 0.110872
R13542 VGND.n844 VGND.n843 0.110872
R13543 VGND.n839 VGND.n838 0.110872
R13544 VGND.n834 VGND.n833 0.110872
R13545 VGND.n829 VGND.n828 0.110872
R13546 VGND.n824 VGND.n823 0.110872
R13547 VGND.n811 VGND.n810 0.110872
R13548 VGND.n870 VGND.n869 0.110872
R13549 VGND.n875 VGND.n874 0.110872
R13550 VGND.n1353 VGND.n1352 0.110872
R13551 VGND.n1649 VGND.n1648 0.110872
R13552 VGND.n1643 VGND.n1642 0.110872
R13553 VGND.n1638 VGND.n1637 0.110872
R13554 VGND.n1633 VGND.n1632 0.110872
R13555 VGND.n1553 VGND.n1552 0.110872
R13556 VGND.n761 VGND.n760 0.110872
R13557 VGND.n1548 VGND.n1547 0.110872
R13558 VGND.n1543 VGND.n1542 0.110872
R13559 VGND.n769 VGND.n768 0.110872
R13560 VGND.n1517 VGND.n1516 0.110872
R13561 VGND.n777 VGND.n776 0.110872
R13562 VGND.n1491 VGND.n1490 0.110872
R13563 VGND.n805 VGND.n804 0.110872
R13564 VGND.n1396 VGND.n1395 0.110872
R13565 VGND.n1391 VGND.n1390 0.110872
R13566 VGND.n2891 VGND.n2890 0.110872
R13567 VGND.n2885 VGND.n2884 0.110872
R13568 VGND.n1572 VGND.n1571 0.110872
R13569 VGND.n1577 VGND.n1576 0.110872
R13570 VGND.n1582 VGND.n1581 0.110872
R13571 VGND.n756 VGND.n755 0.110872
R13572 VGND.n1567 VGND.n1566 0.110872
R13573 VGND.n765 VGND.n764 0.110872
R13574 VGND.n1530 VGND.n1529 0.110872
R13575 VGND.n773 VGND.n772 0.110872
R13576 VGND.n1504 VGND.n1503 0.110872
R13577 VGND.n781 VGND.n780 0.110872
R13578 VGND.n1478 VGND.n1477 0.110872
R13579 VGND.n795 VGND.n794 0.110872
R13580 VGND.n1411 VGND.n1410 0.110872
R13581 VGND.n1609 VGND.n1608 0.110872
R13582 VGND.n1614 VGND.n1613 0.110872
R13583 VGND.n750 VGND.n749 0.110872
R13584 VGND.n1601 VGND.n1600 0.110872
R13585 VGND.n1596 VGND.n1595 0.110872
R13586 VGND.n1459 VGND.n1458 0.110872
R13587 VGND.n791 VGND.n790 0.110872
R13588 VGND.n1454 VGND.n1453 0.110872
R13589 VGND.n1449 VGND.n1448 0.110872
R13590 VGND.n1444 VGND.n1443 0.110872
R13591 VGND.n1439 VGND.n1438 0.110872
R13592 VGND.n1434 VGND.n1433 0.110872
R13593 VGND.n1429 VGND.n1428 0.110872
R13594 VGND.n1424 VGND.n1423 0.110872
R13595 VGND.n885 VGND.n884 0.110872
R13596 VGND.n2911 VGND.n2910 0.110872
R13597 VGND.n2905 VGND.n2904 0.110872
R13598 VGND.n1049 VGND.n1048 0.110872
R13599 VGND.n1058 VGND.n1057 0.110872
R13600 VGND.n1053 VGND.n1052 0.110872
R13601 VGND.n1044 VGND.n1043 0.110872
R13602 VGND.n1070 VGND.n1069 0.110872
R13603 VGND.n1075 VGND.n1074 0.110872
R13604 VGND.n1080 VGND.n1079 0.110872
R13605 VGND.n1085 VGND.n1084 0.110872
R13606 VGND.n1090 VGND.n1089 0.110872
R13607 VGND.n1095 VGND.n1094 0.110872
R13608 VGND.n1029 VGND.n1028 0.110872
R13609 VGND.n1037 VGND.n1036 0.110872
R13610 VGND.n1032 VGND.n1031 0.110872
R13611 VGND.n1169 VGND.n1168 0.110872
R13612 VGND.n1173 VGND.n1172 0.110872
R13613 VGND.n1179 VGND.n1178 0.110872
R13614 VGND.n1186 VGND.n1185 0.110872
R13615 VGND.n1009 VGND.n1008 0.110872
R13616 VGND.n1205 VGND.n1204 0.110872
R13617 VGND.n1211 VGND.n1210 0.110872
R13618 VGND.n1218 VGND.n1217 0.110872
R13619 VGND.n1222 VGND.n1001 0.110872
R13620 VGND.n1244 VGND.n1243 0.110872
R13621 VGND.n1227 VGND.n1225 0.110872
R13622 VGND.n1237 VGND.n1236 0.110872
R13623 VGND.n1232 VGND.n1231 0.110872
R13624 VGND.n1275 VGND.n1274 0.110872
R13625 VGND.n1281 VGND.n1280 0.110872
R13626 VGND.n928 VGND.n927 0.110872
R13627 VGND.n987 VGND.n986 0.110872
R13628 VGND.n982 VGND.n981 0.110872
R13629 VGND.n977 VGND.n976 0.110872
R13630 VGND.n972 VGND.n971 0.110872
R13631 VGND.n967 VGND.n966 0.110872
R13632 VGND.n962 VGND.n961 0.110872
R13633 VGND.n957 VGND.n956 0.110872
R13634 VGND.n952 VGND.n951 0.110872
R13635 VGND.n947 VGND.n946 0.110872
R13636 VGND.n942 VGND.n941 0.110872
R13637 VGND.n937 VGND.n936 0.110872
R13638 VGND.n932 VGND.n931 0.110872
R13639 VGND.n895 VGND.n894 0.110872
R13640 VGND.n1333 VGND.n1332 0.110872
R13641 VGND.n1130 VGND 0.0981562
R13642 VGND.n2214 VGND 0.0981562
R13643 VGND.n1362 VGND 0.0981562
R13644 VGND.n19 VGND 0.0968542
R13645 VGND.n2952 VGND 0.0968542
R13646 VGND.n45 VGND 0.0968542
R13647 VGND VGND.n91 0.0968542
R13648 VGND VGND.n130 0.0968542
R13649 VGND VGND.n499 0.0968542
R13650 VGND VGND.n2280 0.0968542
R13651 VGND VGND.n535 0.0968542
R13652 VGND VGND.n2207 0.0968542
R13653 VGND.n2224 VGND 0.0968542
R13654 VGND.n2982 VGND 0.0968542
R13655 VGND.n2562 VGND 0.088625
R13656 VGND.n2633 VGND 0.0790114
R13657 VGND.n2695 VGND 0.0790114
R13658 VGND.n2690 VGND 0.0790114
R13659 VGND VGND.n2689 0.0790114
R13660 VGND.n2684 VGND 0.0790114
R13661 VGND VGND.n2683 0.0790114
R13662 VGND.n2678 VGND 0.0790114
R13663 VGND VGND.n2677 0.0790114
R13664 VGND.n2709 VGND 0.0790114
R13665 VGND.n2723 VGND 0.0790114
R13666 VGND.n2742 VGND 0.0790114
R13667 VGND.n2761 VGND 0.0790114
R13668 VGND.n2781 VGND 0.0790114
R13669 VGND VGND.n2780 0.0790114
R13670 VGND VGND.n284 0.0790114
R13671 VGND.n2940 VGND 0.0790114
R13672 VGND.n2635 VGND 0.0790114
R13673 VGND.n2693 VGND 0.0790114
R13674 VGND VGND.n2692 0.0790114
R13675 VGND.n2687 VGND 0.0790114
R13676 VGND VGND.n2686 0.0790114
R13677 VGND.n2681 VGND 0.0790114
R13678 VGND VGND.n2680 0.0790114
R13679 VGND.n2675 VGND 0.0790114
R13680 VGND.n2711 VGND 0.0790114
R13681 VGND.n2721 VGND 0.0790114
R13682 VGND.n2744 VGND 0.0790114
R13683 VGND.n2759 VGND 0.0790114
R13684 VGND.n2783 VGND 0.0790114
R13685 VGND.n2784 VGND 0.0790114
R13686 VGND.n2794 VGND 0.0790114
R13687 VGND.n2937 VGND 0.0790114
R13688 VGND VGND.n2559 0.0790114
R13689 VGND VGND.n2558 0.0790114
R13690 VGND VGND.n2557 0.0790114
R13691 VGND VGND.n2556 0.0790114
R13692 VGND VGND.n2555 0.0790114
R13693 VGND VGND.n2554 0.0790114
R13694 VGND VGND.n2553 0.0790114
R13695 VGND VGND.n2552 0.0790114
R13696 VGND VGND.n2551 0.0790114
R13697 VGND VGND.n2550 0.0790114
R13698 VGND VGND.n2549 0.0790114
R13699 VGND VGND.n2548 0.0790114
R13700 VGND VGND.n2547 0.0790114
R13701 VGND.n2798 VGND 0.0790114
R13702 VGND VGND.n2797 0.0790114
R13703 VGND.n2533 VGND 0.0790114
R13704 VGND.n2357 VGND 0.0790114
R13705 VGND.n2373 VGND 0.0790114
R13706 VGND.n2383 VGND 0.0790114
R13707 VGND.n2399 VGND 0.0790114
R13708 VGND.n2409 VGND 0.0790114
R13709 VGND.n2425 VGND 0.0790114
R13710 VGND.n2435 VGND 0.0790114
R13711 VGND.n2451 VGND 0.0790114
R13712 VGND.n2461 VGND 0.0790114
R13713 VGND.n2477 VGND 0.0790114
R13714 VGND.n2487 VGND 0.0790114
R13715 VGND.n2508 VGND 0.0790114
R13716 VGND.n2802 VGND 0.0790114
R13717 VGND VGND.n2801 0.0790114
R13718 VGND.n419 VGND 0.0790114
R13719 VGND.n2530 VGND 0.0790114
R13720 VGND.n2360 VGND 0.0790114
R13721 VGND.n2370 VGND 0.0790114
R13722 VGND.n2386 VGND 0.0790114
R13723 VGND.n2396 VGND 0.0790114
R13724 VGND.n2412 VGND 0.0790114
R13725 VGND.n2422 VGND 0.0790114
R13726 VGND.n2438 VGND 0.0790114
R13727 VGND.n2448 VGND 0.0790114
R13728 VGND.n2464 VGND 0.0790114
R13729 VGND.n2474 VGND 0.0790114
R13730 VGND.n2490 VGND 0.0790114
R13731 VGND.n2505 VGND 0.0790114
R13732 VGND.n2805 VGND 0.0790114
R13733 VGND.n2806 VGND 0.0790114
R13734 VGND.n2819 VGND 0.0790114
R13735 VGND VGND.n2818 0.0790114
R13736 VGND.n1907 VGND 0.0790114
R13737 VGND.n1917 VGND 0.0790114
R13738 VGND.n1918 VGND 0.0790114
R13739 VGND.n1928 VGND 0.0790114
R13740 VGND.n1929 VGND 0.0790114
R13741 VGND.n1939 VGND 0.0790114
R13742 VGND.n1940 VGND 0.0790114
R13743 VGND.n1950 VGND 0.0790114
R13744 VGND.n1951 VGND 0.0790114
R13745 VGND.n1961 VGND 0.0790114
R13746 VGND.n1962 VGND 0.0790114
R13747 VGND.n1972 VGND 0.0790114
R13748 VGND.n1973 VGND 0.0790114
R13749 VGND.n2823 VGND 0.0790114
R13750 VGND VGND.n2822 0.0790114
R13751 VGND.n1990 VGND 0.0790114
R13752 VGND.n2063 VGND 0.0790114
R13753 VGND VGND.n2062 0.0790114
R13754 VGND.n2167 VGND 0.0790114
R13755 VGND VGND.n2166 0.0790114
R13756 VGND.n2159 VGND 0.0790114
R13757 VGND VGND.n2158 0.0790114
R13758 VGND.n2151 VGND 0.0790114
R13759 VGND VGND.n2150 0.0790114
R13760 VGND.n2143 VGND 0.0790114
R13761 VGND VGND.n2142 0.0790114
R13762 VGND.n2135 VGND 0.0790114
R13763 VGND VGND.n2134 0.0790114
R13764 VGND.n2827 VGND 0.0790114
R13765 VGND VGND.n2826 0.0790114
R13766 VGND.n1998 VGND 0.0790114
R13767 VGND VGND.n1997 0.0790114
R13768 VGND.n2066 VGND 0.0790114
R13769 VGND.n2171 VGND 0.0790114
R13770 VGND VGND.n2170 0.0790114
R13771 VGND.n2163 VGND 0.0790114
R13772 VGND VGND.n2162 0.0790114
R13773 VGND.n2155 VGND 0.0790114
R13774 VGND VGND.n2154 0.0790114
R13775 VGND.n2147 VGND 0.0790114
R13776 VGND VGND.n2146 0.0790114
R13777 VGND.n2139 VGND 0.0790114
R13778 VGND VGND.n2138 0.0790114
R13779 VGND.n2131 VGND 0.0790114
R13780 VGND.n2830 VGND 0.0790114
R13781 VGND.n2831 VGND 0.0790114
R13782 VGND.n2844 VGND 0.0790114
R13783 VGND VGND.n2843 0.0790114
R13784 VGND VGND.n1901 0.0790114
R13785 VGND.n2174 VGND 0.0790114
R13786 VGND.n1758 VGND 0.0790114
R13787 VGND.n1768 VGND 0.0790114
R13788 VGND.n1769 VGND 0.0790114
R13789 VGND.n1779 VGND 0.0790114
R13790 VGND.n1780 VGND 0.0790114
R13791 VGND.n1790 VGND 0.0790114
R13792 VGND.n1791 VGND 0.0790114
R13793 VGND.n1801 VGND 0.0790114
R13794 VGND.n1802 VGND 0.0790114
R13795 VGND.n1812 VGND 0.0790114
R13796 VGND.n1813 VGND 0.0790114
R13797 VGND.n2848 VGND 0.0790114
R13798 VGND VGND.n2847 0.0790114
R13799 VGND.n1830 VGND 0.0790114
R13800 VGND VGND.n1899 0.0790114
R13801 VGND.n1685 VGND 0.0790114
R13802 VGND.n1686 VGND 0.0790114
R13803 VGND.n1884 VGND 0.0790114
R13804 VGND VGND.n1883 0.0790114
R13805 VGND.n1876 VGND 0.0790114
R13806 VGND VGND.n1875 0.0790114
R13807 VGND.n1868 VGND 0.0790114
R13808 VGND VGND.n1867 0.0790114
R13809 VGND.n1860 VGND 0.0790114
R13810 VGND VGND.n1859 0.0790114
R13811 VGND.n1852 VGND 0.0790114
R13812 VGND.n2852 VGND 0.0790114
R13813 VGND VGND.n2851 0.0790114
R13814 VGND.n1838 VGND 0.0790114
R13815 VGND VGND.n1837 0.0790114
R13816 VGND.n1896 VGND 0.0790114
R13817 VGND VGND.n1895 0.0790114
R13818 VGND.n1888 VGND 0.0790114
R13819 VGND VGND.n1887 0.0790114
R13820 VGND.n1880 VGND 0.0790114
R13821 VGND VGND.n1879 0.0790114
R13822 VGND.n1872 VGND 0.0790114
R13823 VGND VGND.n1871 0.0790114
R13824 VGND.n1864 VGND 0.0790114
R13825 VGND VGND.n1863 0.0790114
R13826 VGND.n1856 VGND 0.0790114
R13827 VGND VGND.n1855 0.0790114
R13828 VGND.n2855 VGND 0.0790114
R13829 VGND.n2856 VGND 0.0790114
R13830 VGND.n2869 VGND 0.0790114
R13831 VGND VGND.n2868 0.0790114
R13832 VGND.n1349 VGND 0.0790114
R13833 VGND.n1892 VGND 0.0790114
R13834 VGND VGND.n1891 0.0790114
R13835 VGND.n867 VGND 0.0790114
R13836 VGND VGND.n866 0.0790114
R13837 VGND VGND.n865 0.0790114
R13838 VGND VGND.n864 0.0790114
R13839 VGND VGND.n863 0.0790114
R13840 VGND VGND.n862 0.0790114
R13841 VGND VGND.n861 0.0790114
R13842 VGND VGND.n860 0.0790114
R13843 VGND.n1669 VGND 0.0790114
R13844 VGND VGND.n1668 0.0790114
R13845 VGND.n2873 VGND 0.0790114
R13846 VGND VGND.n2872 0.0790114
R13847 VGND.n1654 VGND 0.0790114
R13848 VGND.n1404 VGND 0.0790114
R13849 VGND VGND.n1403 0.0790114
R13850 VGND VGND.n1402 0.0790114
R13851 VGND.n1487 VGND 0.0790114
R13852 VGND.n1497 VGND 0.0790114
R13853 VGND.n1513 VGND 0.0790114
R13854 VGND.n1523 VGND 0.0790114
R13855 VGND.n1539 VGND 0.0790114
R13856 VGND.n1560 VGND 0.0790114
R13857 VGND VGND.n1559 0.0790114
R13858 VGND.n1628 VGND 0.0790114
R13859 VGND.n1629 VGND 0.0790114
R13860 VGND.n2877 VGND 0.0790114
R13861 VGND VGND.n2876 0.0790114
R13862 VGND.n740 VGND 0.0790114
R13863 VGND.n1651 VGND 0.0790114
R13864 VGND.n1407 VGND 0.0790114
R13865 VGND.n1417 VGND 0.0790114
R13866 VGND.n1474 VGND 0.0790114
R13867 VGND.n1484 VGND 0.0790114
R13868 VGND.n1500 VGND 0.0790114
R13869 VGND.n1510 VGND 0.0790114
R13870 VGND.n1526 VGND 0.0790114
R13871 VGND.n1536 VGND 0.0790114
R13872 VGND.n1563 VGND 0.0790114
R13873 VGND.n1588 VGND 0.0790114
R13874 VGND.n1625 VGND 0.0790114
R13875 VGND VGND.n1624 0.0790114
R13876 VGND.n2880 VGND 0.0790114
R13877 VGND.n2881 VGND 0.0790114
R13878 VGND.n2894 VGND 0.0790114
R13879 VGND VGND.n2893 0.0790114
R13880 VGND VGND.n1344 0.0790114
R13881 VGND.n1420 VGND 0.0790114
R13882 VGND.n1471 VGND 0.0790114
R13883 VGND VGND.n1470 0.0790114
R13884 VGND VGND.n1469 0.0790114
R13885 VGND VGND.n1468 0.0790114
R13886 VGND VGND.n1467 0.0790114
R13887 VGND VGND.n1466 0.0790114
R13888 VGND VGND.n1465 0.0790114
R13889 VGND.n1591 VGND 0.0790114
R13890 VGND.n1592 VGND 0.0790114
R13891 VGND.n1621 VGND 0.0790114
R13892 VGND VGND.n1620 0.0790114
R13893 VGND.n2898 VGND 0.0790114
R13894 VGND VGND.n2897 0.0790114
R13895 VGND.n1606 VGND 0.0790114
R13896 VGND.n1103 VGND 0.0790114
R13897 VGND VGND.n1102 0.0790114
R13898 VGND VGND.n1101 0.0790114
R13899 VGND.n1321 VGND 0.0790114
R13900 VGND VGND.n1320 0.0790114
R13901 VGND.n1313 VGND 0.0790114
R13902 VGND VGND.n1312 0.0790114
R13903 VGND.n1305 VGND 0.0790114
R13904 VGND VGND.n1304 0.0790114
R13905 VGND.n1067 VGND 0.0790114
R13906 VGND VGND.n1066 0.0790114
R13907 VGND VGND.n1065 0.0790114
R13908 VGND VGND.n1064 0.0790114
R13909 VGND.n2901 VGND 0.0790114
R13910 VGND.n233 VGND 0.0790114
R13911 VGND.n2913 VGND 0.0790114
R13912 VGND.n1163 VGND 0.0790114
R13913 VGND.n1328 VGND 0.0790114
R13914 VGND VGND.n1327 0.0790114
R13915 VGND.n898 VGND 0.0790114
R13916 VGND.n901 VGND 0.0790114
R13917 VGND.n904 VGND 0.0790114
R13918 VGND.n907 VGND 0.0790114
R13919 VGND.n910 VGND 0.0790114
R13920 VGND.n913 VGND 0.0790114
R13921 VGND.n1298 VGND 0.0790114
R13922 VGND VGND.n1297 0.0790114
R13923 VGND.n1292 VGND 0.0790114
R13924 VGND VGND.n1291 0.0790114
R13925 VGND.n1270 VGND 0.0790114
R13926 VGND.n1285 VGND 0.0790114
R13927 VGND VGND.n1284 0.0790114
R13928 VGND.n1161 VGND 0.0790114
R13929 VGND.n1330 VGND 0.0790114
R13930 VGND.n1325 VGND 0.0790114
R13931 VGND VGND.n1324 0.0790114
R13932 VGND.n1317 VGND 0.0790114
R13933 VGND VGND.n1316 0.0790114
R13934 VGND.n1309 VGND 0.0790114
R13935 VGND VGND.n1308 0.0790114
R13936 VGND.n1301 VGND 0.0790114
R13937 VGND VGND.n1300 0.0790114
R13938 VGND.n1295 VGND 0.0790114
R13939 VGND VGND.n1294 0.0790114
R13940 VGND.n1289 VGND 0.0790114
R13941 VGND VGND.n1288 0.0790114
R13942 VGND VGND.n1287 0.0790114
R13943 VGND.n2916 VGND 0.0790114
R13944 VGND.n2699 VGND.n2698 0.0656596
R13945 VGND.n357 VGND.n355 0.0656596
R13946 VGND.n364 VGND.n362 0.0656596
R13947 VGND.n368 VGND.n367 0.0656596
R13948 VGND.n375 VGND.n373 0.0656596
R13949 VGND.n379 VGND.n378 0.0656596
R13950 VGND.n386 VGND.n384 0.0656596
R13951 VGND.n387 VGND.n325 0.0656596
R13952 VGND.n326 VGND.n314 0.0656596
R13953 VGND.n2726 VGND.n309 0.0656596
R13954 VGND.n312 VGND.n311 0.0656596
R13955 VGND.n2735 VGND.n2734 0.0656596
R13956 VGND.n2730 VGND.n293 0.0656596
R13957 VGND.n296 VGND.n294 0.0656596
R13958 VGND.n2773 VGND.n203 0.0656596
R13959 VGND.n2606 VGND 0.063
R13960 VGND.n2603 VGND 0.063
R13961 VGND.n2600 VGND 0.063
R13962 VGND.n2597 VGND 0.063
R13963 VGND.n2594 VGND 0.063
R13964 VGND.n2591 VGND 0.063
R13965 VGND.n2588 VGND 0.063
R13966 VGND.n2585 VGND 0.063
R13967 VGND.n2582 VGND 0.063
R13968 VGND.n2579 VGND 0.063
R13969 VGND.n2576 VGND 0.063
R13970 VGND.n2573 VGND 0.063
R13971 VGND.n2570 VGND 0.063
R13972 VGND.n2567 VGND 0.063
R13973 VGND.n2564 VGND 0.063
R13974 VGND VGND.n31 0.0603958
R13975 VGND.n3009 VGND 0.0603958
R13976 VGND VGND.n3008 0.0603958
R13977 VGND.n192 VGND 0.0603958
R13978 VGND VGND.n191 0.0603958
R13979 VGND VGND.n2964 0.0603958
R13980 VGND.n2965 VGND 0.0603958
R13981 VGND VGND.n57 0.0603958
R13982 VGND.n64 VGND 0.0603958
R13983 VGND VGND.n63 0.0603958
R13984 VGND.n118 VGND 0.0603958
R13985 VGND.n119 VGND 0.0603958
R13986 VGND.n132 VGND 0.0603958
R13987 VGND VGND.n131 0.0603958
R13988 VGND.n127 VGND 0.0603958
R13989 VGND.n163 VGND 0.0603958
R13990 VGND VGND.n162 0.0603958
R13991 VGND.n1152 VGND 0.0603958
R13992 VGND.n1129 VGND 0.0603958
R13993 VGND VGND.n1128 0.0603958
R13994 VGND.n1125 VGND 0.0603958
R13995 VGND.n501 VGND 0.0603958
R13996 VGND VGND.n500 0.0603958
R13997 VGND.n483 VGND 0.0603958
R13998 VGND.n2282 VGND 0.0603958
R13999 VGND VGND.n2281 0.0603958
R14000 VGND.n2264 VGND 0.0603958
R14001 VGND.n537 VGND 0.0603958
R14002 VGND VGND.n536 0.0603958
R14003 VGND.n519 VGND 0.0603958
R14004 VGND.n2209 VGND 0.0603958
R14005 VGND VGND.n2208 0.0603958
R14006 VGND.n2201 VGND 0.0603958
R14007 VGND.n2198 VGND 0.0603958
R14008 VGND.n2193 VGND 0.0603958
R14009 VGND VGND.n2225 0.0603958
R14010 VGND.n2246 VGND 0.0603958
R14011 VGND VGND.n2245 0.0603958
R14012 VGND VGND.n1363 0.0603958
R14013 VGND.n1384 VGND 0.0603958
R14014 VGND VGND.n1383 0.0603958
R14015 VGND VGND.n2994 0.0603958
R14016 VGND.n2995 VGND 0.0603958
R14017 VGND.n2996 VGND 0.0603958
R14018 VGND.n2698 VGND 0.0574853
R14019 VGND.n357 VGND 0.0574853
R14020 VGND.n364 VGND 0.0574853
R14021 VGND.n367 VGND 0.0574853
R14022 VGND.n375 VGND 0.0574853
R14023 VGND.n378 VGND 0.0574853
R14024 VGND.n386 VGND 0.0574853
R14025 VGND.n325 VGND 0.0574853
R14026 VGND.n314 VGND 0.0574853
R14027 VGND.n309 VGND 0.0574853
R14028 VGND.n311 VGND 0.0574853
R14029 VGND.n2734 VGND 0.0574853
R14030 VGND.n293 VGND 0.0574853
R14031 VGND.n296 VGND 0.0574853
R14032 VGND.n203 VGND 0.0574853
R14033 VGND.n1021 VGND 0.0489375
R14034 VGND.n994 VGND 0.0489375
R14035 VGND.n2630 VGND 0.0489375
R14036 VGND.n204 VGND 0.0489375
R14037 VGND.n334 VGND 0.0489375
R14038 VGND.n2626 VGND 0.0489375
R14039 VGND.n2623 VGND 0.0489375
R14040 VGND.n2620 VGND 0.0489375
R14041 VGND.n2617 VGND 0.0489375
R14042 VGND.n2614 VGND 0.0489375
R14043 VGND.n2611 VGND 0.0489375
R14044 VGND.n322 VGND 0.0489375
R14045 VGND.n315 VGND 0.0489375
R14046 VGND.n306 VGND 0.0489375
R14047 VGND.n299 VGND 0.0489375
R14048 VGND.n2765 VGND 0.0489375
R14049 VGND.n290 VGND 0.0489375
R14050 VGND.n297 VGND 0.0489375
R14051 VGND.n1018 VGND 0.0489375
R14052 VGND.n1015 VGND 0.0489375
R14053 VGND.n1180 VGND 0.0489375
R14054 VGND.n1006 VGND 0.0489375
R14055 VGND.n1004 VGND 0.0489375
R14056 VGND.n1195 VGND 0.0489375
R14057 VGND.n1212 VGND 0.0489375
R14058 VGND.n1000 VGND 0.0489375
R14059 VGND.n1253 VGND 0.0489375
R14060 VGND.n1256 VGND 0.0489375
R14061 VGND.n1259 VGND 0.0489375
R14062 VGND.n1262 VGND 0.0489375
R14063 VGND.n998 VGND 0.0489375
R14064 VGND.n1265 VGND 0.0489375
R14065 VGND VGND.n330 0.037734
R14066 VGND.n286 VGND 0.037734
R14067 VGND.n2787 VGND 0.037734
R14068 VGND.n2752 VGND 0.037734
R14069 VGND.n303 VGND 0.037734
R14070 VGND.n2747 VGND 0.037734
R14071 VGND.n319 VGND 0.037734
R14072 VGND.n2714 VGND 0.037734
R14073 VGND.n393 VGND 0.037734
R14074 VGND.n2668 VGND 0.037734
R14075 VGND.n2663 VGND 0.037734
R14076 VGND.n2658 VGND 0.037734
R14077 VGND.n2653 VGND 0.037734
R14078 VGND.n2648 VGND 0.037734
R14079 VGND.n2643 VGND 0.037734
R14080 VGND.n2638 VGND 0.037734
R14081 VGND VGND.n396 0.037734
R14082 VGND.n2535 VGND 0.037734
R14083 VGND.n2540 VGND 0.037734
R14084 VGND.n414 VGND 0.037734
R14085 VGND.n2287 VGND 0.037734
R14086 VGND.n2292 VGND 0.037734
R14087 VGND.n2297 VGND 0.037734
R14088 VGND.n2302 VGND 0.037734
R14089 VGND.n2307 VGND 0.037734
R14090 VGND.n2312 VGND 0.037734
R14091 VGND.n2317 VGND 0.037734
R14092 VGND.n2322 VGND 0.037734
R14093 VGND.n2327 VGND 0.037734
R14094 VGND.n2332 VGND 0.037734
R14095 VGND.n2337 VGND 0.037734
R14096 VGND.n2342 VGND 0.037734
R14097 VGND VGND.n400 0.037734
R14098 VGND VGND.n2528 0.037734
R14099 VGND.n2521 VGND 0.037734
R14100 VGND.n2516 VGND 0.037734
R14101 VGND.n2511 VGND 0.037734
R14102 VGND.n427 VGND 0.037734
R14103 VGND.n2480 VGND 0.037734
R14104 VGND.n435 VGND 0.037734
R14105 VGND.n2454 VGND 0.037734
R14106 VGND.n443 VGND 0.037734
R14107 VGND.n2428 VGND 0.037734
R14108 VGND.n451 VGND 0.037734
R14109 VGND.n2402 VGND 0.037734
R14110 VGND.n459 VGND 0.037734
R14111 VGND.n2376 VGND 0.037734
R14112 VGND.n471 VGND 0.037734
R14113 VGND VGND.n469 0.037734
R14114 VGND VGND.n2816 0.037734
R14115 VGND.n2809 VGND 0.037734
R14116 VGND.n2498 VGND 0.037734
R14117 VGND.n423 VGND 0.037734
R14118 VGND.n2493 VGND 0.037734
R14119 VGND.n431 VGND 0.037734
R14120 VGND.n2467 VGND 0.037734
R14121 VGND.n439 VGND 0.037734
R14122 VGND.n2441 VGND 0.037734
R14123 VGND.n447 VGND 0.037734
R14124 VGND.n2415 VGND 0.037734
R14125 VGND.n455 VGND 0.037734
R14126 VGND.n2389 VGND 0.037734
R14127 VGND.n463 VGND 0.037734
R14128 VGND.n2363 VGND 0.037734
R14129 VGND VGND.n466 0.037734
R14130 VGND VGND.n1988 0.037734
R14131 VGND.n1981 VGND 0.037734
R14132 VGND.n1976 VGND 0.037734
R14133 VGND.n607 VGND 0.037734
R14134 VGND.n1965 VGND 0.037734
R14135 VGND.n610 VGND 0.037734
R14136 VGND.n1954 VGND 0.037734
R14137 VGND.n613 VGND 0.037734
R14138 VGND.n1943 VGND 0.037734
R14139 VGND.n616 VGND 0.037734
R14140 VGND.n1932 VGND 0.037734
R14141 VGND.n619 VGND 0.037734
R14142 VGND.n1921 VGND 0.037734
R14143 VGND.n622 VGND 0.037734
R14144 VGND.n1910 VGND 0.037734
R14145 VGND VGND.n625 0.037734
R14146 VGND VGND.n1995 0.037734
R14147 VGND.n2000 VGND 0.037734
R14148 VGND.n2005 VGND 0.037734
R14149 VGND.n2010 VGND 0.037734
R14150 VGND.n2015 VGND 0.037734
R14151 VGND.n2020 VGND 0.037734
R14152 VGND.n2025 VGND 0.037734
R14153 VGND.n2030 VGND 0.037734
R14154 VGND.n2035 VGND 0.037734
R14155 VGND.n2040 VGND 0.037734
R14156 VGND.n2045 VGND 0.037734
R14157 VGND.n2050 VGND 0.037734
R14158 VGND.n2055 VGND 0.037734
R14159 VGND.n593 VGND 0.037734
R14160 VGND.n596 VGND 0.037734
R14161 VGND VGND.n590 0.037734
R14162 VGND VGND.n2841 0.037734
R14163 VGND.n2834 VGND 0.037734
R14164 VGND.n2124 VGND 0.037734
R14165 VGND.n584 VGND 0.037734
R14166 VGND.n2119 VGND 0.037734
R14167 VGND.n2114 VGND 0.037734
R14168 VGND.n2109 VGND 0.037734
R14169 VGND.n2104 VGND 0.037734
R14170 VGND.n2099 VGND 0.037734
R14171 VGND.n2094 VGND 0.037734
R14172 VGND.n2089 VGND 0.037734
R14173 VGND.n2084 VGND 0.037734
R14174 VGND.n2079 VGND 0.037734
R14175 VGND.n2074 VGND 0.037734
R14176 VGND.n2069 VGND 0.037734
R14177 VGND VGND.n587 0.037734
R14178 VGND VGND.n1828 0.037734
R14179 VGND.n1821 VGND 0.037734
R14180 VGND.n1816 VGND 0.037734
R14181 VGND.n1740 VGND 0.037734
R14182 VGND.n1805 VGND 0.037734
R14183 VGND.n1743 VGND 0.037734
R14184 VGND.n1794 VGND 0.037734
R14185 VGND.n1746 VGND 0.037734
R14186 VGND.n1783 VGND 0.037734
R14187 VGND.n1749 VGND 0.037734
R14188 VGND.n1772 VGND 0.037734
R14189 VGND.n1752 VGND 0.037734
R14190 VGND.n1761 VGND 0.037734
R14191 VGND VGND.n1757 0.037734
R14192 VGND.n2176 VGND 0.037734
R14193 VGND VGND.n547 0.037734
R14194 VGND VGND.n1835 0.037734
R14195 VGND.n1840 VGND 0.037734
R14196 VGND.n1845 VGND 0.037734
R14197 VGND.n1672 VGND 0.037734
R14198 VGND.n1729 VGND 0.037734
R14199 VGND.n1724 VGND 0.037734
R14200 VGND.n1719 VGND 0.037734
R14201 VGND.n1714 VGND 0.037734
R14202 VGND.n1709 VGND 0.037734
R14203 VGND.n1704 VGND 0.037734
R14204 VGND.n1699 VGND 0.037734
R14205 VGND.n1694 VGND 0.037734
R14206 VGND.n1689 VGND 0.037734
R14207 VGND.n1675 VGND 0.037734
R14208 VGND.n1678 VGND 0.037734
R14209 VGND VGND.n628 0.037734
R14210 VGND VGND.n2866 0.037734
R14211 VGND.n2859 VGND 0.037734
R14212 VGND.n724 VGND 0.037734
R14213 VGND.n666 VGND 0.037734
R14214 VGND.n719 VGND 0.037734
R14215 VGND.n714 VGND 0.037734
R14216 VGND.n709 VGND 0.037734
R14217 VGND.n704 VGND 0.037734
R14218 VGND.n699 VGND 0.037734
R14219 VGND.n694 VGND 0.037734
R14220 VGND.n689 VGND 0.037734
R14221 VGND.n684 VGND 0.037734
R14222 VGND.n679 VGND 0.037734
R14223 VGND.n674 VGND 0.037734
R14224 VGND.n669 VGND 0.037734
R14225 VGND VGND.n632 0.037734
R14226 VGND.n1656 VGND 0.037734
R14227 VGND.n1661 VGND 0.037734
R14228 VGND.n734 VGND 0.037734
R14229 VGND.n853 VGND 0.037734
R14230 VGND.n819 VGND 0.037734
R14231 VGND.n848 VGND 0.037734
R14232 VGND.n843 VGND 0.037734
R14233 VGND.n838 VGND 0.037734
R14234 VGND.n833 VGND 0.037734
R14235 VGND.n828 VGND 0.037734
R14236 VGND.n823 VGND 0.037734
R14237 VGND VGND.n811 0.037734
R14238 VGND.n869 VGND 0.037734
R14239 VGND.n874 VGND 0.037734
R14240 VGND.n1352 VGND 0.037734
R14241 VGND VGND.n879 0.037734
R14242 VGND VGND.n1649 0.037734
R14243 VGND.n1642 VGND 0.037734
R14244 VGND.n1637 VGND 0.037734
R14245 VGND.n1632 VGND 0.037734
R14246 VGND.n1552 VGND 0.037734
R14247 VGND.n760 VGND 0.037734
R14248 VGND.n1547 VGND 0.037734
R14249 VGND.n1542 VGND 0.037734
R14250 VGND.n768 VGND 0.037734
R14251 VGND.n1516 VGND 0.037734
R14252 VGND.n776 VGND 0.037734
R14253 VGND.n1490 VGND 0.037734
R14254 VGND.n804 VGND 0.037734
R14255 VGND.n1395 VGND 0.037734
R14256 VGND.n1390 VGND 0.037734
R14257 VGND VGND.n800 0.037734
R14258 VGND VGND.n2891 0.037734
R14259 VGND.n2884 VGND 0.037734
R14260 VGND.n1571 VGND 0.037734
R14261 VGND.n1576 VGND 0.037734
R14262 VGND.n1581 VGND 0.037734
R14263 VGND.n755 VGND 0.037734
R14264 VGND.n1566 VGND 0.037734
R14265 VGND.n764 VGND 0.037734
R14266 VGND.n1529 VGND 0.037734
R14267 VGND.n772 VGND 0.037734
R14268 VGND.n1503 VGND 0.037734
R14269 VGND.n780 VGND 0.037734
R14270 VGND.n1477 VGND 0.037734
R14271 VGND.n794 VGND 0.037734
R14272 VGND.n1410 VGND 0.037734
R14273 VGND VGND.n797 0.037734
R14274 VGND.n1608 VGND 0.037734
R14275 VGND.n1613 VGND 0.037734
R14276 VGND.n749 VGND 0.037734
R14277 VGND.n1600 VGND 0.037734
R14278 VGND.n1595 VGND 0.037734
R14279 VGND.n1458 VGND 0.037734
R14280 VGND.n790 VGND 0.037734
R14281 VGND.n1453 VGND 0.037734
R14282 VGND.n1448 VGND 0.037734
R14283 VGND.n1443 VGND 0.037734
R14284 VGND.n1438 VGND 0.037734
R14285 VGND.n1433 VGND 0.037734
R14286 VGND.n1428 VGND 0.037734
R14287 VGND.n1423 VGND 0.037734
R14288 VGND.n884 VGND 0.037734
R14289 VGND VGND.n882 0.037734
R14290 VGND VGND.n2911 0.037734
R14291 VGND.n2904 VGND 0.037734
R14292 VGND.n1048 VGND 0.037734
R14293 VGND.n1057 VGND 0.037734
R14294 VGND.n1052 VGND 0.037734
R14295 VGND VGND.n1044 0.037734
R14296 VGND.n1069 VGND 0.037734
R14297 VGND.n1074 VGND 0.037734
R14298 VGND.n1079 VGND 0.037734
R14299 VGND.n1084 VGND 0.037734
R14300 VGND.n1089 VGND 0.037734
R14301 VGND.n1094 VGND 0.037734
R14302 VGND.n1028 VGND 0.037734
R14303 VGND.n1036 VGND 0.037734
R14304 VGND.n1031 VGND 0.037734
R14305 VGND VGND.n1024 0.037734
R14306 VGND VGND.n1014 0.037734
R14307 VGND VGND.n1169 0.037734
R14308 VGND.n1172 VGND 0.037734
R14309 VGND VGND.n1179 0.037734
R14310 VGND.n1185 VGND 0.037734
R14311 VGND.n1008 VGND 0.037734
R14312 VGND.n1204 VGND 0.037734
R14313 VGND VGND.n1211 0.037734
R14314 VGND.n1217 VGND 0.037734
R14315 VGND VGND.n1222 0.037734
R14316 VGND.n1243 VGND 0.037734
R14317 VGND VGND.n1227 0.037734
R14318 VGND.n1236 VGND 0.037734
R14319 VGND.n1231 VGND 0.037734
R14320 VGND.n1274 VGND 0.037734
R14321 VGND VGND.n1281 0.037734
R14322 VGND.n927 VGND 0.037734
R14323 VGND.n986 VGND 0.037734
R14324 VGND.n981 VGND 0.037734
R14325 VGND.n976 VGND 0.037734
R14326 VGND.n971 VGND 0.037734
R14327 VGND.n966 VGND 0.037734
R14328 VGND.n961 VGND 0.037734
R14329 VGND.n956 VGND 0.037734
R14330 VGND.n951 VGND 0.037734
R14331 VGND.n946 VGND 0.037734
R14332 VGND.n941 VGND 0.037734
R14333 VGND.n936 VGND 0.037734
R14334 VGND.n931 VGND 0.037734
R14335 VGND VGND.n895 0.037734
R14336 VGND.n1332 VGND 0.037734
R14337 VGND VGND.n887 0.037734
R14338 VGND.n1156 VGND 0.0343542
R14339 VGND.n1128 VGND 0.0343542
R14340 VGND.n501 VGND 0.0343542
R14341 VGND.n2282 VGND 0.0343542
R14342 VGND.n537 VGND 0.0343542
R14343 VGND.n2209 VGND 0.0343542
R14344 VGND.n2246 VGND 0.0343542
R14345 VGND.n1384 VGND 0.0343542
R14346 VGND.n3009 VGND 0.0330521
R14347 VGND.n192 VGND 0.0330521
R14348 VGND.n2965 VGND 0.0330521
R14349 VGND.n64 VGND 0.0330521
R14350 VGND VGND.n118 0.0330521
R14351 VGND.n132 VGND 0.0330521
R14352 VGND.n163 VGND 0.0330521
R14353 VGND VGND.n2995 0.0330521
R14354 VGND.n33 VGND 0.024
R14355 VGND.n1 VGND 0.024
R14356 VGND.n119 VGND 0.0239375
R14357 VGND.n131 VGND 0.0239375
R14358 VGND.n500 VGND 0.0239375
R14359 VGND.n2281 VGND 0.0239375
R14360 VGND.n536 VGND 0.0239375
R14361 VGND.n3003 VGND 0.0226354
R14362 VGND VGND.n124 0.0226354
R14363 VGND.n1133 VGND 0.0226354
R14364 VGND VGND.n2256 0.0226354
R14365 VGND.n2217 VGND 0.0226354
R14366 VGND.n2208 VGND 0.0226354
R14367 VGND.n2220 VGND 0.0226354
R14368 VGND VGND.n3000 0.0226354
R14369 VGND VGND.n189 0.0213333
R14370 VGND.n191 VGND 0.0213333
R14371 VGND.n58 VGND 0.0213333
R14372 VGND.n113 VGND 0.0213333
R14373 VGND VGND.n90 0.0213333
R14374 VGND VGND.n158 0.0213333
R14375 VGND.n162 VGND 0.0213333
R14376 VGND VGND.n511 0.0213333
R14377 VGND.n2213 VGND 0.0213333
R14378 VGND.n1358 VGND 0.0213333
R14379 VGND VGND.n3024 0.0193356
R14380 VGND.n33 VGND 0.0161667
R14381 VGND.n331 VGND 0.00980851
R14382 VGND.n2936 VGND 0.00980851
R14383 VGND.n2793 VGND 0.00980851
R14384 VGND.n2785 VGND 0.00980851
R14385 VGND VGND.n288 0.00980851
R14386 VGND.n2758 VGND 0.00980851
R14387 VGND.n2745 VGND 0.00980851
R14388 VGND.n2720 VGND 0.00980851
R14389 VGND.n2712 VGND 0.00980851
R14390 VGND.n2674 VGND 0.00980851
R14391 VGND VGND.n350 0.00980851
R14392 VGND VGND.n349 0.00980851
R14393 VGND VGND.n344 0.00980851
R14394 VGND VGND.n343 0.00980851
R14395 VGND VGND.n338 0.00980851
R14396 VGND VGND.n337 0.00980851
R14397 VGND.n2636 VGND 0.00980851
R14398 VGND VGND.n2534 0.00980851
R14399 VGND VGND.n283 0.00980851
R14400 VGND VGND.n282 0.00980851
R14401 VGND.n2546 VGND 0.00980851
R14402 VGND VGND.n412 0.00980851
R14403 VGND VGND.n411 0.00980851
R14404 VGND VGND.n410 0.00980851
R14405 VGND VGND.n409 0.00980851
R14406 VGND VGND.n408 0.00980851
R14407 VGND VGND.n407 0.00980851
R14408 VGND VGND.n406 0.00980851
R14409 VGND VGND.n405 0.00980851
R14410 VGND VGND.n404 0.00980851
R14411 VGND VGND.n403 0.00980851
R14412 VGND VGND.n402 0.00980851
R14413 VGND.n401 VGND 0.00980851
R14414 VGND.n2529 VGND 0.00980851
R14415 VGND VGND.n420 0.00980851
R14416 VGND VGND.n280 0.00980851
R14417 VGND VGND.n279 0.00980851
R14418 VGND.n2509 VGND 0.00980851
R14419 VGND.n2486 VGND 0.00980851
R14420 VGND.n2478 VGND 0.00980851
R14421 VGND.n2460 VGND 0.00980851
R14422 VGND.n2452 VGND 0.00980851
R14423 VGND.n2434 VGND 0.00980851
R14424 VGND.n2426 VGND 0.00980851
R14425 VGND.n2408 VGND 0.00980851
R14426 VGND.n2400 VGND 0.00980851
R14427 VGND.n2382 VGND 0.00980851
R14428 VGND.n2374 VGND 0.00980851
R14429 VGND.n2356 VGND 0.00980851
R14430 VGND.n2817 VGND 0.00980851
R14431 VGND VGND.n273 0.00980851
R14432 VGND.n2807 VGND 0.00980851
R14433 VGND VGND.n277 0.00980851
R14434 VGND.n2504 VGND 0.00980851
R14435 VGND.n2491 VGND 0.00980851
R14436 VGND.n2473 VGND 0.00980851
R14437 VGND.n2465 VGND 0.00980851
R14438 VGND.n2447 VGND 0.00980851
R14439 VGND.n2439 VGND 0.00980851
R14440 VGND.n2421 VGND 0.00980851
R14441 VGND.n2413 VGND 0.00980851
R14442 VGND.n2395 VGND 0.00980851
R14443 VGND.n2387 VGND 0.00980851
R14444 VGND.n2369 VGND 0.00980851
R14445 VGND.n2361 VGND 0.00980851
R14446 VGND.n1989 VGND 0.00980851
R14447 VGND VGND.n271 0.00980851
R14448 VGND VGND.n270 0.00980851
R14449 VGND.n1974 VGND 0.00980851
R14450 VGND.n1971 VGND 0.00980851
R14451 VGND.n1963 VGND 0.00980851
R14452 VGND.n1960 VGND 0.00980851
R14453 VGND.n1952 VGND 0.00980851
R14454 VGND.n1949 VGND 0.00980851
R14455 VGND.n1941 VGND 0.00980851
R14456 VGND.n1938 VGND 0.00980851
R14457 VGND.n1930 VGND 0.00980851
R14458 VGND.n1927 VGND 0.00980851
R14459 VGND.n1919 VGND 0.00980851
R14460 VGND.n1916 VGND 0.00980851
R14461 VGND.n1908 VGND 0.00980851
R14462 VGND.n1996 VGND 0.00980851
R14463 VGND VGND.n1999 0.00980851
R14464 VGND VGND.n268 0.00980851
R14465 VGND VGND.n267 0.00980851
R14466 VGND VGND.n581 0.00980851
R14467 VGND VGND.n580 0.00980851
R14468 VGND VGND.n575 0.00980851
R14469 VGND VGND.n574 0.00980851
R14470 VGND VGND.n569 0.00980851
R14471 VGND VGND.n568 0.00980851
R14472 VGND VGND.n563 0.00980851
R14473 VGND VGND.n562 0.00980851
R14474 VGND VGND.n557 0.00980851
R14475 VGND VGND.n556 0.00980851
R14476 VGND.n2061 VGND 0.00980851
R14477 VGND.n591 VGND 0.00980851
R14478 VGND.n2842 VGND 0.00980851
R14479 VGND VGND.n261 0.00980851
R14480 VGND.n2832 VGND 0.00980851
R14481 VGND VGND.n265 0.00980851
R14482 VGND.n2130 VGND 0.00980851
R14483 VGND VGND.n578 0.00980851
R14484 VGND VGND.n577 0.00980851
R14485 VGND VGND.n572 0.00980851
R14486 VGND VGND.n571 0.00980851
R14487 VGND VGND.n566 0.00980851
R14488 VGND VGND.n565 0.00980851
R14489 VGND VGND.n560 0.00980851
R14490 VGND VGND.n559 0.00980851
R14491 VGND VGND.n554 0.00980851
R14492 VGND VGND.n553 0.00980851
R14493 VGND.n2067 VGND 0.00980851
R14494 VGND.n1829 VGND 0.00980851
R14495 VGND VGND.n259 0.00980851
R14496 VGND VGND.n258 0.00980851
R14497 VGND.n1814 VGND 0.00980851
R14498 VGND.n1811 VGND 0.00980851
R14499 VGND.n1803 VGND 0.00980851
R14500 VGND.n1800 VGND 0.00980851
R14501 VGND.n1792 VGND 0.00980851
R14502 VGND.n1789 VGND 0.00980851
R14503 VGND.n1781 VGND 0.00980851
R14504 VGND.n1778 VGND 0.00980851
R14505 VGND.n1770 VGND 0.00980851
R14506 VGND.n1767 VGND 0.00980851
R14507 VGND.n1759 VGND 0.00980851
R14508 VGND VGND.n2175 0.00980851
R14509 VGND.n548 VGND 0.00980851
R14510 VGND.n1836 VGND 0.00980851
R14511 VGND VGND.n1839 0.00980851
R14512 VGND VGND.n256 0.00980851
R14513 VGND VGND.n255 0.00980851
R14514 VGND.n1851 VGND 0.00980851
R14515 VGND VGND.n662 0.00980851
R14516 VGND VGND.n661 0.00980851
R14517 VGND VGND.n656 0.00980851
R14518 VGND VGND.n655 0.00980851
R14519 VGND VGND.n650 0.00980851
R14520 VGND VGND.n649 0.00980851
R14521 VGND VGND.n644 0.00980851
R14522 VGND VGND.n643 0.00980851
R14523 VGND.n1687 VGND 0.00980851
R14524 VGND.n1684 VGND 0.00980851
R14525 VGND.n629 VGND 0.00980851
R14526 VGND.n2867 VGND 0.00980851
R14527 VGND VGND.n249 0.00980851
R14528 VGND.n2857 VGND 0.00980851
R14529 VGND VGND.n253 0.00980851
R14530 VGND.n730 VGND 0.00980851
R14531 VGND VGND.n664 0.00980851
R14532 VGND VGND.n659 0.00980851
R14533 VGND VGND.n658 0.00980851
R14534 VGND VGND.n653 0.00980851
R14535 VGND VGND.n652 0.00980851
R14536 VGND VGND.n647 0.00980851
R14537 VGND VGND.n646 0.00980851
R14538 VGND VGND.n641 0.00980851
R14539 VGND VGND.n640 0.00980851
R14540 VGND VGND.n634 0.00980851
R14541 VGND.n633 VGND 0.00980851
R14542 VGND VGND.n1655 0.00980851
R14543 VGND VGND.n247 0.00980851
R14544 VGND VGND.n246 0.00980851
R14545 VGND.n1667 VGND 0.00980851
R14546 VGND VGND.n732 0.00980851
R14547 VGND.n859 VGND 0.00980851
R14548 VGND VGND.n817 0.00980851
R14549 VGND VGND.n816 0.00980851
R14550 VGND VGND.n815 0.00980851
R14551 VGND VGND.n814 0.00980851
R14552 VGND VGND.n813 0.00980851
R14553 VGND.n812 VGND 0.00980851
R14554 VGND VGND.n868 0.00980851
R14555 VGND VGND.n637 0.00980851
R14556 VGND VGND.n636 0.00980851
R14557 VGND.n1350 VGND 0.00980851
R14558 VGND.n1650 VGND 0.00980851
R14559 VGND VGND.n741 0.00980851
R14560 VGND VGND.n244 0.00980851
R14561 VGND VGND.n243 0.00980851
R14562 VGND.n1630 VGND 0.00980851
R14563 VGND VGND.n742 0.00980851
R14564 VGND.n1558 VGND 0.00980851
R14565 VGND VGND.n758 0.00980851
R14566 VGND.n1540 VGND 0.00980851
R14567 VGND.n1522 VGND 0.00980851
R14568 VGND.n1514 VGND 0.00980851
R14569 VGND.n1496 VGND 0.00980851
R14570 VGND.n1488 VGND 0.00980851
R14571 VGND.n1401 VGND 0.00980851
R14572 VGND VGND.n802 0.00980851
R14573 VGND.n801 VGND 0.00980851
R14574 VGND.n2892 VGND 0.00980851
R14575 VGND VGND.n236 0.00980851
R14576 VGND.n2882 VGND 0.00980851
R14577 VGND VGND.n240 0.00980851
R14578 VGND VGND.n745 0.00980851
R14579 VGND VGND.n744 0.00980851
R14580 VGND.n1587 VGND 0.00980851
R14581 VGND.n1564 VGND 0.00980851
R14582 VGND.n1535 VGND 0.00980851
R14583 VGND.n1527 VGND 0.00980851
R14584 VGND.n1509 VGND 0.00980851
R14585 VGND.n1501 VGND 0.00980851
R14586 VGND.n1483 VGND 0.00980851
R14587 VGND.n1475 VGND 0.00980851
R14588 VGND.n1416 VGND 0.00980851
R14589 VGND.n1408 VGND 0.00980851
R14590 VGND VGND.n1607 0.00980851
R14591 VGND VGND.n232 0.00980851
R14592 VGND VGND.n231 0.00980851
R14593 VGND.n1619 VGND 0.00980851
R14594 VGND VGND.n747 0.00980851
R14595 VGND.n1593 VGND 0.00980851
R14596 VGND VGND.n751 0.00980851
R14597 VGND.n1464 VGND 0.00980851
R14598 VGND VGND.n788 0.00980851
R14599 VGND VGND.n787 0.00980851
R14600 VGND VGND.n786 0.00980851
R14601 VGND VGND.n785 0.00980851
R14602 VGND VGND.n784 0.00980851
R14603 VGND VGND.n783 0.00980851
R14604 VGND.n1421 VGND 0.00980851
R14605 VGND.n1343 VGND 0.00980851
R14606 VGND.n2912 VGND 0.00980851
R14607 VGND VGND.n228 0.00980851
R14608 VGND.n2902 VGND 0.00980851
R14609 VGND.n1063 VGND 0.00980851
R14610 VGND VGND.n1046 0.00980851
R14611 VGND.n1045 VGND 0.00980851
R14612 VGND VGND.n1068 0.00980851
R14613 VGND VGND.n912 0.00980851
R14614 VGND VGND.n911 0.00980851
R14615 VGND VGND.n906 0.00980851
R14616 VGND VGND.n905 0.00980851
R14617 VGND VGND.n900 0.00980851
R14618 VGND VGND.n899 0.00980851
R14619 VGND.n1100 VGND 0.00980851
R14620 VGND VGND.n1026 0.00980851
R14621 VGND.n1025 VGND 0.00980851
R14622 VGND.n1165 VGND 0.00980851
R14623 VGND.n1170 VGND 0.00980851
R14624 VGND VGND.n1011 0.00980851
R14625 VGND.n1183 VGND 0.00980851
R14626 VGND.n1191 VGND 0.00980851
R14627 VGND.n1202 VGND 0.00980851
R14628 VGND VGND.n1003 0.00980851
R14629 VGND.n1215 VGND 0.00980851
R14630 VGND.n1249 VGND 0.00980851
R14631 VGND.n1223 VGND 0.00980851
R14632 VGND VGND.n1242 0.00980851
R14633 VGND.n1228 VGND 0.00980851
R14634 VGND VGND.n1235 0.00980851
R14635 VGND.n1272 VGND 0.00980851
R14636 VGND VGND.n997 0.00980851
R14637 VGND.n1282 VGND 0.00980851
R14638 VGND.n2917 VGND 0.00980851
R14639 VGND.n992 VGND 0.00980851
R14640 VGND VGND.n925 0.00980851
R14641 VGND VGND.n924 0.00980851
R14642 VGND VGND.n920 0.00980851
R14643 VGND VGND.n919 0.00980851
R14644 VGND VGND.n915 0.00980851
R14645 VGND VGND.n914 0.00980851
R14646 VGND VGND.n909 0.00980851
R14647 VGND VGND.n908 0.00980851
R14648 VGND VGND.n903 0.00980851
R14649 VGND VGND.n902 0.00980851
R14650 VGND VGND.n897 0.00980851
R14651 VGND.n896 VGND 0.00980851
R14652 VGND VGND.n1331 0.00980851
R14653 VGND.n888 VGND 0.00980851
R14654 VGND.n2698 VGND.n2697 0.00182979
R14655 VGND.n358 VGND.n357 0.00182979
R14656 VGND.n365 VGND.n364 0.00182979
R14657 VGND.n367 VGND.n354 0.00182979
R14658 VGND.n376 VGND.n375 0.00182979
R14659 VGND.n378 VGND.n353 0.00182979
R14660 VGND.n389 VGND.n386 0.00182979
R14661 VGND.n2707 VGND.n325 0.00182979
R14662 VGND.n2725 VGND.n314 0.00182979
R14663 VGND.n2740 VGND.n309 0.00182979
R14664 VGND.n311 VGND.n300 0.00182979
R14665 VGND.n2734 VGND.n2733 0.00182979
R14666 VGND.n2778 VGND.n293 0.00182979
R14667 VGND.n2772 VGND.n296 0.00182979
R14668 VGND.n2942 VGND.n203 0.00182979
R14669 XThR.Tn[6].n2 XThR.Tn[6].n0 332.332
R14670 XThR.Tn[6].n2 XThR.Tn[6].n1 296.493
R14671 XThR.Tn[6] XThR.Tn[6].n82 161.363
R14672 XThR.Tn[6] XThR.Tn[6].n77 161.363
R14673 XThR.Tn[6] XThR.Tn[6].n72 161.363
R14674 XThR.Tn[6] XThR.Tn[6].n67 161.363
R14675 XThR.Tn[6] XThR.Tn[6].n62 161.363
R14676 XThR.Tn[6] XThR.Tn[6].n57 161.363
R14677 XThR.Tn[6] XThR.Tn[6].n52 161.363
R14678 XThR.Tn[6] XThR.Tn[6].n47 161.363
R14679 XThR.Tn[6] XThR.Tn[6].n42 161.363
R14680 XThR.Tn[6] XThR.Tn[6].n37 161.363
R14681 XThR.Tn[6] XThR.Tn[6].n32 161.363
R14682 XThR.Tn[6] XThR.Tn[6].n27 161.363
R14683 XThR.Tn[6] XThR.Tn[6].n22 161.363
R14684 XThR.Tn[6] XThR.Tn[6].n17 161.363
R14685 XThR.Tn[6] XThR.Tn[6].n12 161.363
R14686 XThR.Tn[6] XThR.Tn[6].n10 161.363
R14687 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R14688 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R14689 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R14690 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R14691 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R14692 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R14693 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R14694 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R14695 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R14696 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R14697 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R14698 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R14699 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R14700 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R14701 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R14702 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R14703 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R14704 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R14705 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R14706 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R14707 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R14708 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R14709 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R14710 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R14711 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R14712 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R14713 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R14714 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R14715 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R14716 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R14717 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R14718 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R14719 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R14720 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R14721 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R14722 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R14723 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R14724 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R14725 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R14726 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R14727 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R14728 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R14729 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R14730 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R14731 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R14732 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R14733 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R14734 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R14735 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R14736 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R14737 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R14738 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R14739 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R14740 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R14741 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R14742 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R14743 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R14744 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R14745 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R14746 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R14747 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R14748 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R14749 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R14750 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R14751 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R14752 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R14753 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R14754 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R14755 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R14756 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R14757 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R14758 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R14759 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R14760 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R14761 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R14762 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R14763 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R14764 XThR.Tn[6].n5 XThR.Tn[6].n3 135.249
R14765 XThR.Tn[6].n5 XThR.Tn[6].n4 98.982
R14766 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R14767 XThR.Tn[6].n9 XThR.Tn[6].n8 98.982
R14768 XThR.Tn[6].n7 XThR.Tn[6].n5 36.2672
R14769 XThR.Tn[6].n9 XThR.Tn[6].n7 36.2672
R14770 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R14771 XThR.Tn[6].n0 XThR.Tn[6].t2 26.5955
R14772 XThR.Tn[6].n0 XThR.Tn[6].t1 26.5955
R14773 XThR.Tn[6].n1 XThR.Tn[6].t3 26.5955
R14774 XThR.Tn[6].n1 XThR.Tn[6].t0 26.5955
R14775 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R14776 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R14777 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R14778 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R14779 XThR.Tn[6].n6 XThR.Tn[6].t7 24.9236
R14780 XThR.Tn[6].n6 XThR.Tn[6].t6 24.9236
R14781 XThR.Tn[6].n8 XThR.Tn[6].t4 24.9236
R14782 XThR.Tn[6].n8 XThR.Tn[6].t5 24.9236
R14783 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R14784 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R14785 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R14786 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R14787 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R14788 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R14789 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R14790 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R14791 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R14792 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R14793 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R14794 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R14795 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R14796 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R14797 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R14798 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R14799 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R14800 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R14801 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R14802 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R14803 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R14804 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R14805 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R14806 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R14807 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R14808 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R14809 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R14810 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R14811 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R14812 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R14813 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R14814 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R14815 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R14816 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R14817 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R14818 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R14819 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R14820 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R14821 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R14822 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R14823 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R14824 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R14825 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R14826 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R14827 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R14828 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R14829 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R14830 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R14831 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R14832 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R14833 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R14834 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R14835 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R14836 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R14837 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R14838 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R14839 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R14840 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R14841 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R14842 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R14843 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R14844 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R14845 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R14846 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R14847 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R14848 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R14849 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R14850 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R14851 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R14852 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R14853 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R14854 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R14855 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R14856 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R14857 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R14858 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R14859 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R14860 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R14861 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R14862 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R14863 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R14864 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R14865 XThR.Tn[6] XThR.Tn[6].n87 0.038
R14866 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R14867 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R14868 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R14869 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R14870 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R14871 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R14872 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R14873 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R14874 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R14875 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R14876 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R14877 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R14878 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R14879 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R14880 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R14881 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R14882 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R14883 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R14884 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R14885 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R14886 XThR.Tn[14].n87 XThR.Tn[14].n85 202.095
R14887 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R14888 XThR.Tn[14] XThR.Tn[14].n78 161.363
R14889 XThR.Tn[14] XThR.Tn[14].n73 161.363
R14890 XThR.Tn[14] XThR.Tn[14].n68 161.363
R14891 XThR.Tn[14] XThR.Tn[14].n63 161.363
R14892 XThR.Tn[14] XThR.Tn[14].n58 161.363
R14893 XThR.Tn[14] XThR.Tn[14].n53 161.363
R14894 XThR.Tn[14] XThR.Tn[14].n48 161.363
R14895 XThR.Tn[14] XThR.Tn[14].n43 161.363
R14896 XThR.Tn[14] XThR.Tn[14].n38 161.363
R14897 XThR.Tn[14] XThR.Tn[14].n33 161.363
R14898 XThR.Tn[14] XThR.Tn[14].n28 161.363
R14899 XThR.Tn[14] XThR.Tn[14].n23 161.363
R14900 XThR.Tn[14] XThR.Tn[14].n18 161.363
R14901 XThR.Tn[14] XThR.Tn[14].n13 161.363
R14902 XThR.Tn[14] XThR.Tn[14].n8 161.363
R14903 XThR.Tn[14] XThR.Tn[14].n6 161.363
R14904 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R14905 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R14906 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R14907 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R14908 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R14909 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R14910 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R14911 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R14912 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R14913 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R14914 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R14915 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R14916 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R14917 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R14918 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R14919 XThR.Tn[14].n78 XThR.Tn[14].t51 161.106
R14920 XThR.Tn[14].n73 XThR.Tn[14].t58 161.106
R14921 XThR.Tn[14].n68 XThR.Tn[14].t39 161.106
R14922 XThR.Tn[14].n63 XThR.Tn[14].t22 161.106
R14923 XThR.Tn[14].n58 XThR.Tn[14].t49 161.106
R14924 XThR.Tn[14].n53 XThR.Tn[14].t12 161.106
R14925 XThR.Tn[14].n48 XThR.Tn[14].t56 161.106
R14926 XThR.Tn[14].n43 XThR.Tn[14].t36 161.106
R14927 XThR.Tn[14].n38 XThR.Tn[14].t19 161.106
R14928 XThR.Tn[14].n33 XThR.Tn[14].t25 161.106
R14929 XThR.Tn[14].n28 XThR.Tn[14].t73 161.106
R14930 XThR.Tn[14].n23 XThR.Tn[14].t38 161.106
R14931 XThR.Tn[14].n18 XThR.Tn[14].t72 161.106
R14932 XThR.Tn[14].n13 XThR.Tn[14].t54 161.106
R14933 XThR.Tn[14].n8 XThR.Tn[14].t13 161.106
R14934 XThR.Tn[14].n6 XThR.Tn[14].t62 161.106
R14935 XThR.Tn[14].n79 XThR.Tn[14].t32 159.978
R14936 XThR.Tn[14].n74 XThR.Tn[14].t37 159.978
R14937 XThR.Tn[14].n69 XThR.Tn[14].t20 159.978
R14938 XThR.Tn[14].n64 XThR.Tn[14].t68 159.978
R14939 XThR.Tn[14].n59 XThR.Tn[14].t30 159.978
R14940 XThR.Tn[14].n54 XThR.Tn[14].t55 159.978
R14941 XThR.Tn[14].n49 XThR.Tn[14].t35 159.978
R14942 XThR.Tn[14].n44 XThR.Tn[14].t16 159.978
R14943 XThR.Tn[14].n39 XThR.Tn[14].t66 159.978
R14944 XThR.Tn[14].n34 XThR.Tn[14].t71 159.978
R14945 XThR.Tn[14].n29 XThR.Tn[14].t53 159.978
R14946 XThR.Tn[14].n24 XThR.Tn[14].t18 159.978
R14947 XThR.Tn[14].n19 XThR.Tn[14].t52 159.978
R14948 XThR.Tn[14].n14 XThR.Tn[14].t34 159.978
R14949 XThR.Tn[14].n9 XThR.Tn[14].t60 159.978
R14950 XThR.Tn[14].n78 XThR.Tn[14].t41 145.038
R14951 XThR.Tn[14].n73 XThR.Tn[14].t65 145.038
R14952 XThR.Tn[14].n68 XThR.Tn[14].t45 145.038
R14953 XThR.Tn[14].n63 XThR.Tn[14].t26 145.038
R14954 XThR.Tn[14].n58 XThR.Tn[14].t59 145.038
R14955 XThR.Tn[14].n53 XThR.Tn[14].t40 145.038
R14956 XThR.Tn[14].n48 XThR.Tn[14].t46 145.038
R14957 XThR.Tn[14].n43 XThR.Tn[14].t27 145.038
R14958 XThR.Tn[14].n38 XThR.Tn[14].t23 145.038
R14959 XThR.Tn[14].n33 XThR.Tn[14].t57 145.038
R14960 XThR.Tn[14].n28 XThR.Tn[14].t15 145.038
R14961 XThR.Tn[14].n23 XThR.Tn[14].t44 145.038
R14962 XThR.Tn[14].n18 XThR.Tn[14].t14 145.038
R14963 XThR.Tn[14].n13 XThR.Tn[14].t64 145.038
R14964 XThR.Tn[14].n8 XThR.Tn[14].t24 145.038
R14965 XThR.Tn[14].n6 XThR.Tn[14].t69 145.038
R14966 XThR.Tn[14].n79 XThR.Tn[14].t43 143.911
R14967 XThR.Tn[14].n74 XThR.Tn[14].t70 143.911
R14968 XThR.Tn[14].n69 XThR.Tn[14].t48 143.911
R14969 XThR.Tn[14].n64 XThR.Tn[14].t31 143.911
R14970 XThR.Tn[14].n59 XThR.Tn[14].t63 143.911
R14971 XThR.Tn[14].n54 XThR.Tn[14].t42 143.911
R14972 XThR.Tn[14].n49 XThR.Tn[14].t50 143.911
R14973 XThR.Tn[14].n44 XThR.Tn[14].t33 143.911
R14974 XThR.Tn[14].n39 XThR.Tn[14].t29 143.911
R14975 XThR.Tn[14].n34 XThR.Tn[14].t61 143.911
R14976 XThR.Tn[14].n29 XThR.Tn[14].t21 143.911
R14977 XThR.Tn[14].n24 XThR.Tn[14].t47 143.911
R14978 XThR.Tn[14].n19 XThR.Tn[14].t17 143.911
R14979 XThR.Tn[14].n14 XThR.Tn[14].t67 143.911
R14980 XThR.Tn[14].n9 XThR.Tn[14].t28 143.911
R14981 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R14982 XThR.Tn[14].n0 XThR.Tn[14].t0 26.5955
R14983 XThR.Tn[14].n0 XThR.Tn[14].t1 26.5955
R14984 XThR.Tn[14].n85 XThR.Tn[14].t10 26.5955
R14985 XThR.Tn[14].n85 XThR.Tn[14].t11 26.5955
R14986 XThR.Tn[14].n86 XThR.Tn[14].t8 26.5955
R14987 XThR.Tn[14].n86 XThR.Tn[14].t9 26.5955
R14988 XThR.Tn[14].n1 XThR.Tn[14].t2 26.5955
R14989 XThR.Tn[14].n1 XThR.Tn[14].t3 26.5955
R14990 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R14991 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R14992 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R14993 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R14994 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R14995 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R14996 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R14997 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R14998 XThR.Tn[14] XThR.Tn[14].n7 5.34038
R14999 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R15000 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R15001 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R15002 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R15003 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R15004 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R15005 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R15006 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R15007 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R15008 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R15009 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R15010 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R15011 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R15012 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R15013 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R15014 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R15015 XThR.Tn[14].n12 XThR.Tn[14] 2.52282
R15016 XThR.Tn[14].n17 XThR.Tn[14] 2.52282
R15017 XThR.Tn[14].n22 XThR.Tn[14] 2.52282
R15018 XThR.Tn[14].n27 XThR.Tn[14] 2.52282
R15019 XThR.Tn[14].n32 XThR.Tn[14] 2.52282
R15020 XThR.Tn[14].n37 XThR.Tn[14] 2.52282
R15021 XThR.Tn[14].n42 XThR.Tn[14] 2.52282
R15022 XThR.Tn[14].n47 XThR.Tn[14] 2.52282
R15023 XThR.Tn[14].n52 XThR.Tn[14] 2.52282
R15024 XThR.Tn[14].n57 XThR.Tn[14] 2.52282
R15025 XThR.Tn[14].n62 XThR.Tn[14] 2.52282
R15026 XThR.Tn[14].n67 XThR.Tn[14] 2.52282
R15027 XThR.Tn[14].n72 XThR.Tn[14] 2.52282
R15028 XThR.Tn[14].n77 XThR.Tn[14] 2.52282
R15029 XThR.Tn[14].n82 XThR.Tn[14] 2.52282
R15030 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R15031 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R15032 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R15033 XThR.Tn[14].n80 XThR.Tn[14] 1.08677
R15034 XThR.Tn[14].n75 XThR.Tn[14] 1.08677
R15035 XThR.Tn[14].n70 XThR.Tn[14] 1.08677
R15036 XThR.Tn[14].n65 XThR.Tn[14] 1.08677
R15037 XThR.Tn[14].n60 XThR.Tn[14] 1.08677
R15038 XThR.Tn[14].n55 XThR.Tn[14] 1.08677
R15039 XThR.Tn[14].n50 XThR.Tn[14] 1.08677
R15040 XThR.Tn[14].n45 XThR.Tn[14] 1.08677
R15041 XThR.Tn[14].n40 XThR.Tn[14] 1.08677
R15042 XThR.Tn[14].n35 XThR.Tn[14] 1.08677
R15043 XThR.Tn[14].n30 XThR.Tn[14] 1.08677
R15044 XThR.Tn[14].n25 XThR.Tn[14] 1.08677
R15045 XThR.Tn[14].n20 XThR.Tn[14] 1.08677
R15046 XThR.Tn[14].n15 XThR.Tn[14] 1.08677
R15047 XThR.Tn[14].n10 XThR.Tn[14] 1.08677
R15048 XThR.Tn[14] XThR.Tn[14].n12 0.839786
R15049 XThR.Tn[14] XThR.Tn[14].n17 0.839786
R15050 XThR.Tn[14] XThR.Tn[14].n22 0.839786
R15051 XThR.Tn[14] XThR.Tn[14].n27 0.839786
R15052 XThR.Tn[14] XThR.Tn[14].n32 0.839786
R15053 XThR.Tn[14] XThR.Tn[14].n37 0.839786
R15054 XThR.Tn[14] XThR.Tn[14].n42 0.839786
R15055 XThR.Tn[14] XThR.Tn[14].n47 0.839786
R15056 XThR.Tn[14] XThR.Tn[14].n52 0.839786
R15057 XThR.Tn[14] XThR.Tn[14].n57 0.839786
R15058 XThR.Tn[14] XThR.Tn[14].n62 0.839786
R15059 XThR.Tn[14] XThR.Tn[14].n67 0.839786
R15060 XThR.Tn[14] XThR.Tn[14].n72 0.839786
R15061 XThR.Tn[14] XThR.Tn[14].n77 0.839786
R15062 XThR.Tn[14] XThR.Tn[14].n82 0.839786
R15063 XThR.Tn[14].n7 XThR.Tn[14] 0.499542
R15064 XThR.Tn[14].n81 XThR.Tn[14] 0.063
R15065 XThR.Tn[14].n76 XThR.Tn[14] 0.063
R15066 XThR.Tn[14].n71 XThR.Tn[14] 0.063
R15067 XThR.Tn[14].n66 XThR.Tn[14] 0.063
R15068 XThR.Tn[14].n61 XThR.Tn[14] 0.063
R15069 XThR.Tn[14].n56 XThR.Tn[14] 0.063
R15070 XThR.Tn[14].n51 XThR.Tn[14] 0.063
R15071 XThR.Tn[14].n46 XThR.Tn[14] 0.063
R15072 XThR.Tn[14].n41 XThR.Tn[14] 0.063
R15073 XThR.Tn[14].n36 XThR.Tn[14] 0.063
R15074 XThR.Tn[14].n31 XThR.Tn[14] 0.063
R15075 XThR.Tn[14].n26 XThR.Tn[14] 0.063
R15076 XThR.Tn[14].n21 XThR.Tn[14] 0.063
R15077 XThR.Tn[14].n16 XThR.Tn[14] 0.063
R15078 XThR.Tn[14].n11 XThR.Tn[14] 0.063
R15079 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R15080 XThR.Tn[14] XThR.Tn[14].n83 0.038
R15081 XThR.Tn[14].n7 XThR.Tn[14] 0.0143889
R15082 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00771154
R15083 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00771154
R15084 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00771154
R15085 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00771154
R15086 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00771154
R15087 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00771154
R15088 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00771154
R15089 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00771154
R15090 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00771154
R15091 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00771154
R15092 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00771154
R15093 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00771154
R15094 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00771154
R15095 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00771154
R15096 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00771154
R15097 Vbias.n992 Vbias.t0 651.571
R15098 Vbias.n992 Vbias.t1 651.571
R15099 Vbias.n993 Vbias.t5 651.571
R15100 Vbias.n993 Vbias.t4 651.571
R15101 Vbias.n332 Vbias.t255 119.309
R15102 Vbias.n378 Vbias.t189 119.309
R15103 Vbias.n379 Vbias.t56 119.309
R15104 Vbias.n329 Vbias.t210 119.309
R15105 Vbias.n287 Vbias.t81 119.309
R15106 Vbias.n279 Vbias.t181 119.309
R15107 Vbias.n283 Vbias.t104 119.309
R15108 Vbias.n275 Vbias.t184 119.309
R15109 Vbias.n189 Vbias.t59 119.309
R15110 Vbias.n144 Vbias.t77 119.309
R15111 Vbias.n184 Vbias.t100 119.309
R15112 Vbias.n140 Vbias.t116 119.309
R15113 Vbias.n673 Vbias.t250 119.309
R15114 Vbias.n97 Vbias.t11 119.309
R15115 Vbias.n5 Vbias.t141 119.309
R15116 Vbias.n52 Vbias.t52 119.309
R15117 Vbias.n53 Vbias.t124 119.309
R15118 Vbias.n49 Vbias.t196 119.309
R15119 Vbias.n435 Vbias.t74 119.309
R15120 Vbias.n338 Vbias.t211 119.309
R15121 Vbias.n328 Vbias.t26 119.309
R15122 Vbias.n326 Vbias.t95 119.309
R15123 Vbias.n572 Vbias.t257 119.309
R15124 Vbias.n273 Vbias.t123 119.309
R15125 Vbias.n271 Vbias.t261 119.309
R15126 Vbias.n192 Vbias.t78 119.309
R15127 Vbias.n145 Vbias.t149 119.309
R15128 Vbias.n147 Vbias.t117 119.309
R15129 Vbias.n784 Vbias.t190 119.309
R15130 Vbias.n100 Vbias.t12 119.309
R15131 Vbias.n98 Vbias.t83 119.309
R15132 Vbias.n92 Vbias.t155 119.309
R15133 Vbias.n51 Vbias.t125 119.309
R15134 Vbias.n48 Vbias.t36 119.309
R15135 Vbias.n432 Vbias.t169 119.309
R15136 Vbias.n341 Vbias.t54 119.309
R15137 Vbias.n321 Vbias.t127 119.309
R15138 Vbias.n323 Vbias.t198 119.309
R15139 Vbias.n569 Vbias.t98 119.309
R15140 Vbias.n268 Vbias.t221 119.309
R15141 Vbias.n270 Vbias.t103 119.309
R15142 Vbias.n195 Vbias.t175 119.309
R15143 Vbias.n150 Vbias.t252 119.309
R15144 Vbias.n148 Vbias.t217 119.309
R15145 Vbias.n787 Vbias.t32 119.309
R15146 Vbias.n101 Vbias.t108 119.309
R15147 Vbias.n103 Vbias.t180 119.309
R15148 Vbias.n89 Vbias.t256 119.309
R15149 Vbias.n46 Vbias.t224 119.309
R15150 Vbias.n43 Vbias.t51 119.309
R15151 Vbias.n429 Vbias.t177 119.309
R15152 Vbias.n344 Vbias.t63 119.309
R15153 Vbias.n320 Vbias.t134 119.309
R15154 Vbias.n318 Vbias.t209 119.309
R15155 Vbias.n566 Vbias.t110 119.309
R15156 Vbias.n267 Vbias.t236 119.309
R15157 Vbias.n265 Vbias.t112 119.309
R15158 Vbias.n198 Vbias.t183 119.309
R15159 Vbias.n151 Vbias.t259 119.309
R15160 Vbias.n153 Vbias.t230 119.309
R15161 Vbias.n790 Vbias.t43 119.309
R15162 Vbias.n106 Vbias.t118 119.309
R15163 Vbias.n104 Vbias.t192 119.309
R15164 Vbias.n86 Vbias.t9 119.309
R15165 Vbias.n45 Vbias.t238 119.309
R15166 Vbias.n42 Vbias.t136 119.309
R15167 Vbias.n426 Vbias.t10 119.309
R15168 Vbias.n347 Vbias.t147 119.309
R15169 Vbias.n315 Vbias.t219 119.309
R15170 Vbias.n317 Vbias.t33 119.309
R15171 Vbias.n563 Vbias.t201 119.309
R15172 Vbias.n262 Vbias.t61 119.309
R15173 Vbias.n264 Vbias.t203 119.309
R15174 Vbias.n201 Vbias.t18 119.309
R15175 Vbias.n156 Vbias.t88 119.309
R15176 Vbias.n154 Vbias.t58 119.309
R15177 Vbias.n793 Vbias.t130 119.309
R15178 Vbias.n107 Vbias.t208 119.309
R15179 Vbias.n109 Vbias.t24 119.309
R15180 Vbias.n83 Vbias.t94 119.309
R15181 Vbias.n40 Vbias.t64 119.309
R15182 Vbias.n37 Vbias.t222 119.309
R15183 Vbias.n423 Vbias.t96 119.309
R15184 Vbias.n350 Vbias.t240 119.309
R15185 Vbias.n314 Vbias.t53 119.309
R15186 Vbias.n312 Vbias.t126 119.309
R15187 Vbias.n560 Vbias.t29 119.309
R15188 Vbias.n261 Vbias.t150 119.309
R15189 Vbias.n259 Vbias.t31 119.309
R15190 Vbias.n204 Vbias.t102 119.309
R15191 Vbias.n157 Vbias.t174 119.309
R15192 Vbias.n159 Vbias.t145 119.309
R15193 Vbias.n796 Vbias.t216 119.309
R15194 Vbias.n112 Vbias.t35 119.309
R15195 Vbias.n110 Vbias.t107 119.309
R15196 Vbias.n80 Vbias.t178 119.309
R15197 Vbias.n39 Vbias.t151 119.309
R15198 Vbias.n36 Vbias.t55 119.309
R15199 Vbias.n420 Vbias.t179 119.309
R15200 Vbias.n353 Vbias.t67 119.309
R15201 Vbias.n309 Vbias.t140 119.309
R15202 Vbias.n311 Vbias.t213 119.309
R15203 Vbias.n557 Vbias.t111 119.309
R15204 Vbias.n256 Vbias.t239 119.309
R15205 Vbias.n258 Vbias.t115 119.309
R15206 Vbias.n207 Vbias.t187 119.309
R15207 Vbias.n162 Vbias.t6 119.309
R15208 Vbias.n160 Vbias.t232 119.309
R15209 Vbias.n799 Vbias.t45 119.309
R15210 Vbias.n113 Vbias.t122 119.309
R15211 Vbias.n115 Vbias.t195 119.309
R15212 Vbias.n77 Vbias.t13 119.309
R15213 Vbias.n34 Vbias.t242 119.309
R15214 Vbias.n31 Vbias.t142 119.309
R15215 Vbias.n417 Vbias.t14 119.309
R15216 Vbias.n356 Vbias.t153 119.309
R15217 Vbias.n308 Vbias.t225 119.309
R15218 Vbias.n306 Vbias.t37 119.309
R15219 Vbias.n554 Vbias.t204 119.309
R15220 Vbias.n255 Vbias.t69 119.309
R15221 Vbias.n253 Vbias.t207 119.309
R15222 Vbias.n210 Vbias.t23 119.309
R15223 Vbias.n163 Vbias.t93 119.309
R15224 Vbias.n165 Vbias.t62 119.309
R15225 Vbias.n802 Vbias.t133 119.309
R15226 Vbias.n118 Vbias.t214 119.309
R15227 Vbias.n116 Vbias.t28 119.309
R15228 Vbias.n74 Vbias.t97 119.309
R15229 Vbias.n33 Vbias.t71 119.309
R15230 Vbias.n30 Vbias.t164 119.309
R15231 Vbias.n414 Vbias.t34 119.309
R15232 Vbias.n359 Vbias.t173 119.309
R15233 Vbias.n303 Vbias.t248 119.309
R15234 Vbias.n305 Vbias.t65 119.309
R15235 Vbias.n551 Vbias.t226 119.309
R15236 Vbias.n250 Vbias.t89 119.309
R15237 Vbias.n252 Vbias.t229 119.309
R15238 Vbias.n213 Vbias.t40 119.309
R15239 Vbias.n168 Vbias.t113 119.309
R15240 Vbias.n166 Vbias.t86 119.309
R15241 Vbias.n805 Vbias.t158 119.309
R15242 Vbias.n119 Vbias.t235 119.309
R15243 Vbias.n121 Vbias.t48 119.309
R15244 Vbias.n71 Vbias.t120 119.309
R15245 Vbias.n28 Vbias.t91 119.309
R15246 Vbias.n25 Vbias.t241 119.309
R15247 Vbias.n411 Vbias.t106 119.309
R15248 Vbias.n362 Vbias.t249 119.309
R15249 Vbias.n302 Vbias.t66 119.309
R15250 Vbias.n300 Vbias.t138 119.309
R15251 Vbias.n548 Vbias.t38 119.309
R15252 Vbias.n249 Vbias.t162 119.309
R15253 Vbias.n247 Vbias.t41 119.309
R15254 Vbias.n216 Vbias.t114 119.309
R15255 Vbias.n169 Vbias.t186 119.309
R15256 Vbias.n171 Vbias.t159 119.309
R15257 Vbias.n808 Vbias.t231 119.309
R15258 Vbias.n124 Vbias.t49 119.309
R15259 Vbias.n122 Vbias.t121 119.309
R15260 Vbias.n68 Vbias.t194 119.309
R15261 Vbias.n27 Vbias.t166 119.309
R15262 Vbias.n24 Vbias.t70 119.309
R15263 Vbias.n408 Vbias.t197 119.309
R15264 Vbias.n365 Vbias.t79 119.309
R15265 Vbias.n297 Vbias.t152 119.309
R15266 Vbias.n299 Vbias.t223 119.309
R15267 Vbias.n545 Vbias.t129 119.309
R15268 Vbias.n244 Vbias.t251 119.309
R15269 Vbias.n246 Vbias.t131 119.309
R15270 Vbias.n219 Vbias.t206 119.309
R15271 Vbias.n174 Vbias.t22 119.309
R15272 Vbias.n172 Vbias.t246 119.309
R15273 Vbias.n811 Vbias.t60 119.309
R15274 Vbias.n125 Vbias.t139 119.309
R15275 Vbias.n127 Vbias.t212 119.309
R15276 Vbias.n65 Vbias.t27 119.309
R15277 Vbias.n22 Vbias.t253 119.309
R15278 Vbias.n19 Vbias.t90 119.309
R15279 Vbias.n405 Vbias.t218 119.309
R15280 Vbias.n368 Vbias.t101 119.309
R15281 Vbias.n296 Vbias.t172 119.309
R15282 Vbias.n294 Vbias.t247 119.309
R15283 Vbias.n542 Vbias.t154 119.309
R15284 Vbias.n243 Vbias.t17 119.309
R15285 Vbias.n241 Vbias.t157 119.309
R15286 Vbias.n222 Vbias.t228 119.309
R15287 Vbias.n175 Vbias.t39 119.309
R15288 Vbias.n177 Vbias.t16 119.309
R15289 Vbias.n814 Vbias.t85 119.309
R15290 Vbias.n130 Vbias.t161 119.309
R15291 Vbias.n128 Vbias.t234 119.309
R15292 Vbias.n62 Vbias.t47 119.309
R15293 Vbias.n21 Vbias.t20 119.309
R15294 Vbias.n18 Vbias.t243 119.309
R15295 Vbias.n402 Vbias.t109 119.309
R15296 Vbias.n371 Vbias.t254 119.309
R15297 Vbias.n291 Vbias.t72 119.309
R15298 Vbias.n293 Vbias.t143 119.309
R15299 Vbias.n539 Vbias.t42 119.309
R15300 Vbias.n238 Vbias.t167 119.309
R15301 Vbias.n240 Vbias.t46 119.309
R15302 Vbias.n225 Vbias.t119 119.309
R15303 Vbias.n180 Vbias.t191 119.309
R15304 Vbias.n178 Vbias.t163 119.309
R15305 Vbias.n817 Vbias.t237 119.309
R15306 Vbias.n131 Vbias.t57 119.309
R15307 Vbias.n133 Vbias.t128 119.309
R15308 Vbias.n59 Vbias.t200 119.309
R15309 Vbias.n16 Vbias.t168 119.309
R15310 Vbias.n11 Vbias.t7 119.309
R15311 Vbias.n399 Vbias.t137 119.309
R15312 Vbias.n374 Vbias.t21 119.309
R15313 Vbias.n290 Vbias.t92 119.309
R15314 Vbias.n288 Vbias.t165 119.309
R15315 Vbias.n536 Vbias.t73 119.309
R15316 Vbias.n237 Vbias.t185 119.309
R15317 Vbias.n235 Vbias.t75 119.309
R15318 Vbias.n228 Vbias.t144 119.309
R15319 Vbias.n181 Vbias.t215 119.309
R15320 Vbias.n183 Vbias.t182 119.309
R15321 Vbias.n820 Vbias.t258 119.309
R15322 Vbias.n136 Vbias.t76 119.309
R15323 Vbias.n134 Vbias.t148 119.309
R15324 Vbias.n56 Vbias.t220 119.309
R15325 Vbias.n13 Vbias.t188 119.309
R15326 Vbias.n10 Vbias.t19 119.309
R15327 Vbias.n333 Vbias.t146 119.309
R15328 Vbias.n334 Vbias.t30 119.309
R15329 Vbias.n336 Vbias.t99 119.309
R15330 Vbias.n520 Vbias.t170 119.309
R15331 Vbias.n280 Vbias.t80 119.309
R15332 Vbias.n282 Vbias.t202 119.309
R15333 Vbias.n657 Vbias.t84 119.309
R15334 Vbias.n231 Vbias.t156 119.309
R15335 Vbias.n233 Vbias.t227 119.309
R15336 Vbias.n698 Vbias.t199 119.309
R15337 Vbias.n139 Vbias.t15 119.309
R15338 Vbias.n137 Vbias.t87 119.309
R15339 Vbias.n666 Vbias.t160 119.309
R15340 Vbias.n6 Vbias.t233 119.309
R15341 Vbias.n8 Vbias.t205 119.309
R15342 Vbias.n1 Vbias.t176 119.309
R15343 Vbias.n2 Vbias.t105 119.309
R15344 Vbias.n55 Vbias.t82 119.309
R15345 Vbias.n669 Vbias.t68 119.309
R15346 Vbias.n901 Vbias.t193 119.309
R15347 Vbias.n678 Vbias.t171 119.309
R15348 Vbias.n141 Vbias.t44 119.309
R15349 Vbias.n186 Vbias.t132 119.309
R15350 Vbias.n190 Vbias.t260 119.309
R15351 Vbias.n660 Vbias.t245 119.309
R15352 Vbias.n274 Vbias.t50 119.309
R15353 Vbias.n284 Vbias.t244 119.309
R15354 Vbias.n324 Vbias.t25 119.309
R15355 Vbias.n390 Vbias.t8 119.309
R15356 Vbias.n330 Vbias.t135 119.309
R15357 Vbias.n995 Vbias.t2 77.1775
R15358 Vbias.n995 Vbias.t3 34.3847
R15359 Vbias.n994 Vbias.n992 4.78773
R15360 Vbias.n994 Vbias.n993 4.78773
R15361 Vbias.n381 Vbias.n379 4.5005
R15362 Vbias.n436 Vbias.n435 4.5005
R15363 Vbias.n339 Vbias.n338 4.5005
R15364 Vbias.n443 Vbias.n328 4.5005
R15365 Vbias.n446 Vbias.n326 4.5005
R15366 Vbias.n573 Vbias.n572 4.5005
R15367 Vbias.n580 Vbias.n273 4.5005
R15368 Vbias.n583 Vbias.n271 4.5005
R15369 Vbias.n193 Vbias.n192 4.5005
R15370 Vbias.n777 Vbias.n145 4.5005
R15371 Vbias.n774 Vbias.n147 4.5005
R15372 Vbias.n785 Vbias.n784 4.5005
R15373 Vbias.n904 Vbias.n100 4.5005
R15374 Vbias.n907 Vbias.n98 4.5005
R15375 Vbias.n93 Vbias.n92 4.5005
R15376 Vbias.n915 Vbias.n51 4.5005
R15377 Vbias.n917 Vbias.n49 4.5005
R15378 Vbias.n433 Vbias.n432 4.5005
R15379 Vbias.n342 Vbias.n341 4.5005
R15380 Vbias.n452 Vbias.n321 4.5005
R15381 Vbias.n449 Vbias.n323 4.5005
R15382 Vbias.n570 Vbias.n569 4.5005
R15383 Vbias.n589 Vbias.n268 4.5005
R15384 Vbias.n586 Vbias.n270 4.5005
R15385 Vbias.n196 Vbias.n195 4.5005
R15386 Vbias.n768 Vbias.n150 4.5005
R15387 Vbias.n771 Vbias.n148 4.5005
R15388 Vbias.n788 Vbias.n787 4.5005
R15389 Vbias.n899 Vbias.n101 4.5005
R15390 Vbias.n896 Vbias.n103 4.5005
R15391 Vbias.n90 Vbias.n89 4.5005
R15392 Vbias.n922 Vbias.n46 4.5005
R15393 Vbias.n920 Vbias.n48 4.5005
R15394 Vbias.n430 Vbias.n429 4.5005
R15395 Vbias.n345 Vbias.n344 4.5005
R15396 Vbias.n455 Vbias.n320 4.5005
R15397 Vbias.n458 Vbias.n318 4.5005
R15398 Vbias.n567 Vbias.n566 4.5005
R15399 Vbias.n592 Vbias.n267 4.5005
R15400 Vbias.n595 Vbias.n265 4.5005
R15401 Vbias.n199 Vbias.n198 4.5005
R15402 Vbias.n765 Vbias.n151 4.5005
R15403 Vbias.n762 Vbias.n153 4.5005
R15404 Vbias.n791 Vbias.n790 4.5005
R15405 Vbias.n890 Vbias.n106 4.5005
R15406 Vbias.n893 Vbias.n104 4.5005
R15407 Vbias.n87 Vbias.n86 4.5005
R15408 Vbias.n925 Vbias.n45 4.5005
R15409 Vbias.n927 Vbias.n43 4.5005
R15410 Vbias.n427 Vbias.n426 4.5005
R15411 Vbias.n348 Vbias.n347 4.5005
R15412 Vbias.n464 Vbias.n315 4.5005
R15413 Vbias.n461 Vbias.n317 4.5005
R15414 Vbias.n564 Vbias.n563 4.5005
R15415 Vbias.n601 Vbias.n262 4.5005
R15416 Vbias.n598 Vbias.n264 4.5005
R15417 Vbias.n202 Vbias.n201 4.5005
R15418 Vbias.n756 Vbias.n156 4.5005
R15419 Vbias.n759 Vbias.n154 4.5005
R15420 Vbias.n794 Vbias.n793 4.5005
R15421 Vbias.n887 Vbias.n107 4.5005
R15422 Vbias.n884 Vbias.n109 4.5005
R15423 Vbias.n84 Vbias.n83 4.5005
R15424 Vbias.n932 Vbias.n40 4.5005
R15425 Vbias.n930 Vbias.n42 4.5005
R15426 Vbias.n424 Vbias.n423 4.5005
R15427 Vbias.n351 Vbias.n350 4.5005
R15428 Vbias.n467 Vbias.n314 4.5005
R15429 Vbias.n470 Vbias.n312 4.5005
R15430 Vbias.n561 Vbias.n560 4.5005
R15431 Vbias.n604 Vbias.n261 4.5005
R15432 Vbias.n607 Vbias.n259 4.5005
R15433 Vbias.n205 Vbias.n204 4.5005
R15434 Vbias.n753 Vbias.n157 4.5005
R15435 Vbias.n750 Vbias.n159 4.5005
R15436 Vbias.n797 Vbias.n796 4.5005
R15437 Vbias.n878 Vbias.n112 4.5005
R15438 Vbias.n881 Vbias.n110 4.5005
R15439 Vbias.n81 Vbias.n80 4.5005
R15440 Vbias.n935 Vbias.n39 4.5005
R15441 Vbias.n937 Vbias.n37 4.5005
R15442 Vbias.n421 Vbias.n420 4.5005
R15443 Vbias.n354 Vbias.n353 4.5005
R15444 Vbias.n476 Vbias.n309 4.5005
R15445 Vbias.n473 Vbias.n311 4.5005
R15446 Vbias.n558 Vbias.n557 4.5005
R15447 Vbias.n613 Vbias.n256 4.5005
R15448 Vbias.n610 Vbias.n258 4.5005
R15449 Vbias.n208 Vbias.n207 4.5005
R15450 Vbias.n744 Vbias.n162 4.5005
R15451 Vbias.n747 Vbias.n160 4.5005
R15452 Vbias.n800 Vbias.n799 4.5005
R15453 Vbias.n875 Vbias.n113 4.5005
R15454 Vbias.n872 Vbias.n115 4.5005
R15455 Vbias.n78 Vbias.n77 4.5005
R15456 Vbias.n942 Vbias.n34 4.5005
R15457 Vbias.n940 Vbias.n36 4.5005
R15458 Vbias.n418 Vbias.n417 4.5005
R15459 Vbias.n357 Vbias.n356 4.5005
R15460 Vbias.n479 Vbias.n308 4.5005
R15461 Vbias.n482 Vbias.n306 4.5005
R15462 Vbias.n555 Vbias.n554 4.5005
R15463 Vbias.n616 Vbias.n255 4.5005
R15464 Vbias.n619 Vbias.n253 4.5005
R15465 Vbias.n211 Vbias.n210 4.5005
R15466 Vbias.n741 Vbias.n163 4.5005
R15467 Vbias.n738 Vbias.n165 4.5005
R15468 Vbias.n803 Vbias.n802 4.5005
R15469 Vbias.n866 Vbias.n118 4.5005
R15470 Vbias.n869 Vbias.n116 4.5005
R15471 Vbias.n75 Vbias.n74 4.5005
R15472 Vbias.n945 Vbias.n33 4.5005
R15473 Vbias.n947 Vbias.n31 4.5005
R15474 Vbias.n415 Vbias.n414 4.5005
R15475 Vbias.n360 Vbias.n359 4.5005
R15476 Vbias.n488 Vbias.n303 4.5005
R15477 Vbias.n485 Vbias.n305 4.5005
R15478 Vbias.n552 Vbias.n551 4.5005
R15479 Vbias.n625 Vbias.n250 4.5005
R15480 Vbias.n622 Vbias.n252 4.5005
R15481 Vbias.n214 Vbias.n213 4.5005
R15482 Vbias.n732 Vbias.n168 4.5005
R15483 Vbias.n735 Vbias.n166 4.5005
R15484 Vbias.n806 Vbias.n805 4.5005
R15485 Vbias.n863 Vbias.n119 4.5005
R15486 Vbias.n860 Vbias.n121 4.5005
R15487 Vbias.n72 Vbias.n71 4.5005
R15488 Vbias.n952 Vbias.n28 4.5005
R15489 Vbias.n950 Vbias.n30 4.5005
R15490 Vbias.n412 Vbias.n411 4.5005
R15491 Vbias.n363 Vbias.n362 4.5005
R15492 Vbias.n491 Vbias.n302 4.5005
R15493 Vbias.n494 Vbias.n300 4.5005
R15494 Vbias.n549 Vbias.n548 4.5005
R15495 Vbias.n628 Vbias.n249 4.5005
R15496 Vbias.n631 Vbias.n247 4.5005
R15497 Vbias.n217 Vbias.n216 4.5005
R15498 Vbias.n729 Vbias.n169 4.5005
R15499 Vbias.n726 Vbias.n171 4.5005
R15500 Vbias.n809 Vbias.n808 4.5005
R15501 Vbias.n854 Vbias.n124 4.5005
R15502 Vbias.n857 Vbias.n122 4.5005
R15503 Vbias.n69 Vbias.n68 4.5005
R15504 Vbias.n955 Vbias.n27 4.5005
R15505 Vbias.n957 Vbias.n25 4.5005
R15506 Vbias.n409 Vbias.n408 4.5005
R15507 Vbias.n366 Vbias.n365 4.5005
R15508 Vbias.n500 Vbias.n297 4.5005
R15509 Vbias.n497 Vbias.n299 4.5005
R15510 Vbias.n546 Vbias.n545 4.5005
R15511 Vbias.n637 Vbias.n244 4.5005
R15512 Vbias.n634 Vbias.n246 4.5005
R15513 Vbias.n220 Vbias.n219 4.5005
R15514 Vbias.n720 Vbias.n174 4.5005
R15515 Vbias.n723 Vbias.n172 4.5005
R15516 Vbias.n812 Vbias.n811 4.5005
R15517 Vbias.n851 Vbias.n125 4.5005
R15518 Vbias.n848 Vbias.n127 4.5005
R15519 Vbias.n66 Vbias.n65 4.5005
R15520 Vbias.n962 Vbias.n22 4.5005
R15521 Vbias.n960 Vbias.n24 4.5005
R15522 Vbias.n406 Vbias.n405 4.5005
R15523 Vbias.n369 Vbias.n368 4.5005
R15524 Vbias.n503 Vbias.n296 4.5005
R15525 Vbias.n506 Vbias.n294 4.5005
R15526 Vbias.n543 Vbias.n542 4.5005
R15527 Vbias.n640 Vbias.n243 4.5005
R15528 Vbias.n643 Vbias.n241 4.5005
R15529 Vbias.n223 Vbias.n222 4.5005
R15530 Vbias.n717 Vbias.n175 4.5005
R15531 Vbias.n714 Vbias.n177 4.5005
R15532 Vbias.n815 Vbias.n814 4.5005
R15533 Vbias.n842 Vbias.n130 4.5005
R15534 Vbias.n845 Vbias.n128 4.5005
R15535 Vbias.n63 Vbias.n62 4.5005
R15536 Vbias.n965 Vbias.n21 4.5005
R15537 Vbias.n967 Vbias.n19 4.5005
R15538 Vbias.n403 Vbias.n402 4.5005
R15539 Vbias.n372 Vbias.n371 4.5005
R15540 Vbias.n512 Vbias.n291 4.5005
R15541 Vbias.n509 Vbias.n293 4.5005
R15542 Vbias.n540 Vbias.n539 4.5005
R15543 Vbias.n649 Vbias.n238 4.5005
R15544 Vbias.n646 Vbias.n240 4.5005
R15545 Vbias.n226 Vbias.n225 4.5005
R15546 Vbias.n708 Vbias.n180 4.5005
R15547 Vbias.n711 Vbias.n178 4.5005
R15548 Vbias.n818 Vbias.n817 4.5005
R15549 Vbias.n839 Vbias.n131 4.5005
R15550 Vbias.n836 Vbias.n133 4.5005
R15551 Vbias.n60 Vbias.n59 4.5005
R15552 Vbias.n972 Vbias.n16 4.5005
R15553 Vbias.n970 Vbias.n18 4.5005
R15554 Vbias.n400 Vbias.n399 4.5005
R15555 Vbias.n375 Vbias.n374 4.5005
R15556 Vbias.n515 Vbias.n290 4.5005
R15557 Vbias.n518 Vbias.n288 4.5005
R15558 Vbias.n537 Vbias.n536 4.5005
R15559 Vbias.n652 Vbias.n237 4.5005
R15560 Vbias.n655 Vbias.n235 4.5005
R15561 Vbias.n229 Vbias.n228 4.5005
R15562 Vbias.n705 Vbias.n181 4.5005
R15563 Vbias.n702 Vbias.n183 4.5005
R15564 Vbias.n821 Vbias.n820 4.5005
R15565 Vbias.n830 Vbias.n136 4.5005
R15566 Vbias.n833 Vbias.n134 4.5005
R15567 Vbias.n57 Vbias.n56 4.5005
R15568 Vbias.n975 Vbias.n13 4.5005
R15569 Vbias.n977 Vbias.n11 4.5005
R15570 Vbias.n397 Vbias.n333 4.5005
R15571 Vbias.n335 Vbias.n334 4.5005
R15572 Vbias.n394 Vbias.n336 4.5005
R15573 Vbias.n521 Vbias.n520 4.5005
R15574 Vbias.n534 Vbias.n280 4.5005
R15575 Vbias.n531 Vbias.n282 4.5005
R15576 Vbias.n658 Vbias.n657 4.5005
R15577 Vbias.n689 Vbias.n231 4.5005
R15578 Vbias.n686 Vbias.n233 4.5005
R15579 Vbias.n699 Vbias.n698 4.5005
R15580 Vbias.n824 Vbias.n139 4.5005
R15581 Vbias.n827 Vbias.n137 4.5005
R15582 Vbias.n667 Vbias.n666 4.5005
R15583 Vbias.n983 Vbias.n6 4.5005
R15584 Vbias.n9 Vbias.n8 4.5005
R15585 Vbias.n980 Vbias.n10 4.5005
R15586 Vbias.n989 Vbias.n1 4.5005
R15587 Vbias.n54 Vbias.n53 4.5005
R15588 Vbias.n913 Vbias.n52 4.5005
R15589 Vbias.n3 Vbias.n2 4.5005
R15590 Vbias.n986 Vbias.n5 4.5005
R15591 Vbias.n95 Vbias.n55 4.5005
R15592 Vbias.n909 Vbias.n97 4.5005
R15593 Vbias.n670 Vbias.n669 4.5005
R15594 Vbias.n675 Vbias.n673 4.5005
R15595 Vbias.n902 Vbias.n901 4.5005
R15596 Vbias.n783 Vbias.n140 4.5005
R15597 Vbias.n679 Vbias.n678 4.5005
R15598 Vbias.n696 Vbias.n184 4.5005
R15599 Vbias.n142 Vbias.n141 4.5005
R15600 Vbias.n779 Vbias.n144 4.5005
R15601 Vbias.n187 Vbias.n186 4.5005
R15602 Vbias.n692 Vbias.n189 4.5005
R15603 Vbias.n191 Vbias.n190 4.5005
R15604 Vbias.n276 Vbias.n275 4.5005
R15605 Vbias.n661 Vbias.n660 4.5005
R15606 Vbias.n528 Vbias.n283 4.5005
R15607 Vbias.n578 Vbias.n274 4.5005
R15608 Vbias.n575 Vbias.n279 4.5005
R15609 Vbias.n285 Vbias.n284 4.5005
R15610 Vbias.n524 Vbias.n287 4.5005
R15611 Vbias.n325 Vbias.n324 4.5005
R15612 Vbias.n441 Vbias.n329 4.5005
R15613 Vbias.n391 Vbias.n390 4.5005
R15614 Vbias.n383 Vbias.n378 4.5005
R15615 Vbias.n331 Vbias.n330 4.5005
R15616 Vbias.n438 Vbias.n332 4.5005
R15617 Vbias.n54 Vbias 3.50727
R15618 Vbias Vbias.n913 3.50727
R15619 Vbias.n95 Vbias 3.50727
R15620 Vbias.n909 Vbias 3.50727
R15621 Vbias Vbias.n902 3.50727
R15622 Vbias Vbias.n783 3.50727
R15623 Vbias Vbias.n142 3.50727
R15624 Vbias.n779 Vbias 3.50727
R15625 Vbias Vbias.n191 3.50727
R15626 Vbias.n276 Vbias 3.50727
R15627 Vbias Vbias.n578 3.50727
R15628 Vbias.n575 Vbias 3.50727
R15629 Vbias Vbias.n325 3.50727
R15630 Vbias Vbias.n441 3.50727
R15631 Vbias Vbias.n331 3.50727
R15632 Vbias.n438 Vbias 3.50727
R15633 Vbias.n990 Vbias.n989 3.4105
R15634 Vbias.n980 Vbias.n979 3.4105
R15635 Vbias.n978 Vbias.n977 3.4105
R15636 Vbias.n970 Vbias.n969 3.4105
R15637 Vbias.n968 Vbias.n967 3.4105
R15638 Vbias.n960 Vbias.n959 3.4105
R15639 Vbias.n958 Vbias.n957 3.4105
R15640 Vbias.n950 Vbias.n949 3.4105
R15641 Vbias.n948 Vbias.n947 3.4105
R15642 Vbias.n940 Vbias.n939 3.4105
R15643 Vbias.n938 Vbias.n937 3.4105
R15644 Vbias.n930 Vbias.n929 3.4105
R15645 Vbias.n928 Vbias.n927 3.4105
R15646 Vbias.n920 Vbias.n919 3.4105
R15647 Vbias.n918 Vbias.n917 3.4105
R15648 Vbias.n915 Vbias.n914 3.4105
R15649 Vbias.n923 Vbias.n922 3.4105
R15650 Vbias.n925 Vbias.n924 3.4105
R15651 Vbias.n933 Vbias.n932 3.4105
R15652 Vbias.n935 Vbias.n934 3.4105
R15653 Vbias.n943 Vbias.n942 3.4105
R15654 Vbias.n945 Vbias.n944 3.4105
R15655 Vbias.n953 Vbias.n952 3.4105
R15656 Vbias.n955 Vbias.n954 3.4105
R15657 Vbias.n963 Vbias.n962 3.4105
R15658 Vbias.n965 Vbias.n964 3.4105
R15659 Vbias.n973 Vbias.n972 3.4105
R15660 Vbias.n975 Vbias.n974 3.4105
R15661 Vbias.n15 Vbias.n9 3.4105
R15662 Vbias.n14 Vbias.n3 3.4105
R15663 Vbias.n986 Vbias.n985 3.4105
R15664 Vbias.n984 Vbias.n983 3.4105
R15665 Vbias.n58 Vbias.n57 3.4105
R15666 Vbias.n61 Vbias.n60 3.4105
R15667 Vbias.n64 Vbias.n63 3.4105
R15668 Vbias.n67 Vbias.n66 3.4105
R15669 Vbias.n70 Vbias.n69 3.4105
R15670 Vbias.n73 Vbias.n72 3.4105
R15671 Vbias.n76 Vbias.n75 3.4105
R15672 Vbias.n79 Vbias.n78 3.4105
R15673 Vbias.n82 Vbias.n81 3.4105
R15674 Vbias.n85 Vbias.n84 3.4105
R15675 Vbias.n88 Vbias.n87 3.4105
R15676 Vbias.n91 Vbias.n90 3.4105
R15677 Vbias.n94 Vbias.n93 3.4105
R15678 Vbias.n908 Vbias.n907 3.4105
R15679 Vbias.n896 Vbias.n895 3.4105
R15680 Vbias.n894 Vbias.n893 3.4105
R15681 Vbias.n884 Vbias.n883 3.4105
R15682 Vbias.n882 Vbias.n881 3.4105
R15683 Vbias.n872 Vbias.n871 3.4105
R15684 Vbias.n870 Vbias.n869 3.4105
R15685 Vbias.n860 Vbias.n859 3.4105
R15686 Vbias.n858 Vbias.n857 3.4105
R15687 Vbias.n848 Vbias.n847 3.4105
R15688 Vbias.n846 Vbias.n845 3.4105
R15689 Vbias.n836 Vbias.n835 3.4105
R15690 Vbias.n834 Vbias.n833 3.4105
R15691 Vbias.n668 Vbias.n667 3.4105
R15692 Vbias.n671 Vbias.n670 3.4105
R15693 Vbias.n676 Vbias.n675 3.4105
R15694 Vbias.n828 Vbias.n827 3.4105
R15695 Vbias.n830 Vbias.n829 3.4105
R15696 Vbias.n840 Vbias.n839 3.4105
R15697 Vbias.n842 Vbias.n841 3.4105
R15698 Vbias.n852 Vbias.n851 3.4105
R15699 Vbias.n854 Vbias.n853 3.4105
R15700 Vbias.n864 Vbias.n863 3.4105
R15701 Vbias.n866 Vbias.n865 3.4105
R15702 Vbias.n876 Vbias.n875 3.4105
R15703 Vbias.n878 Vbias.n877 3.4105
R15704 Vbias.n888 Vbias.n887 3.4105
R15705 Vbias.n890 Vbias.n889 3.4105
R15706 Vbias.n900 Vbias.n899 3.4105
R15707 Vbias.n904 Vbias.n903 3.4105
R15708 Vbias.n786 Vbias.n785 3.4105
R15709 Vbias.n789 Vbias.n788 3.4105
R15710 Vbias.n792 Vbias.n791 3.4105
R15711 Vbias.n795 Vbias.n794 3.4105
R15712 Vbias.n798 Vbias.n797 3.4105
R15713 Vbias.n801 Vbias.n800 3.4105
R15714 Vbias.n804 Vbias.n803 3.4105
R15715 Vbias.n807 Vbias.n806 3.4105
R15716 Vbias.n810 Vbias.n809 3.4105
R15717 Vbias.n813 Vbias.n812 3.4105
R15718 Vbias.n816 Vbias.n815 3.4105
R15719 Vbias.n819 Vbias.n818 3.4105
R15720 Vbias.n822 Vbias.n821 3.4105
R15721 Vbias.n824 Vbias.n823 3.4105
R15722 Vbias.n680 Vbias.n679 3.4105
R15723 Vbias.n697 Vbias.n696 3.4105
R15724 Vbias.n700 Vbias.n699 3.4105
R15725 Vbias.n702 Vbias.n701 3.4105
R15726 Vbias.n712 Vbias.n711 3.4105
R15727 Vbias.n714 Vbias.n713 3.4105
R15728 Vbias.n724 Vbias.n723 3.4105
R15729 Vbias.n726 Vbias.n725 3.4105
R15730 Vbias.n736 Vbias.n735 3.4105
R15731 Vbias.n738 Vbias.n737 3.4105
R15732 Vbias.n748 Vbias.n747 3.4105
R15733 Vbias.n750 Vbias.n749 3.4105
R15734 Vbias.n760 Vbias.n759 3.4105
R15735 Vbias.n762 Vbias.n761 3.4105
R15736 Vbias.n772 Vbias.n771 3.4105
R15737 Vbias.n774 Vbias.n773 3.4105
R15738 Vbias.n778 Vbias.n777 3.4105
R15739 Vbias.n768 Vbias.n767 3.4105
R15740 Vbias.n766 Vbias.n765 3.4105
R15741 Vbias.n756 Vbias.n755 3.4105
R15742 Vbias.n754 Vbias.n753 3.4105
R15743 Vbias.n744 Vbias.n743 3.4105
R15744 Vbias.n742 Vbias.n741 3.4105
R15745 Vbias.n732 Vbias.n731 3.4105
R15746 Vbias.n730 Vbias.n729 3.4105
R15747 Vbias.n720 Vbias.n719 3.4105
R15748 Vbias.n718 Vbias.n717 3.4105
R15749 Vbias.n708 Vbias.n707 3.4105
R15750 Vbias.n706 Vbias.n705 3.4105
R15751 Vbias.n686 Vbias.n685 3.4105
R15752 Vbias.n684 Vbias.n187 3.4105
R15753 Vbias.n692 Vbias.n691 3.4105
R15754 Vbias.n690 Vbias.n689 3.4105
R15755 Vbias.n230 Vbias.n229 3.4105
R15756 Vbias.n227 Vbias.n226 3.4105
R15757 Vbias.n224 Vbias.n223 3.4105
R15758 Vbias.n221 Vbias.n220 3.4105
R15759 Vbias.n218 Vbias.n217 3.4105
R15760 Vbias.n215 Vbias.n214 3.4105
R15761 Vbias.n212 Vbias.n211 3.4105
R15762 Vbias.n209 Vbias.n208 3.4105
R15763 Vbias.n206 Vbias.n205 3.4105
R15764 Vbias.n203 Vbias.n202 3.4105
R15765 Vbias.n200 Vbias.n199 3.4105
R15766 Vbias.n197 Vbias.n196 3.4105
R15767 Vbias.n194 Vbias.n193 3.4105
R15768 Vbias.n584 Vbias.n583 3.4105
R15769 Vbias.n586 Vbias.n585 3.4105
R15770 Vbias.n596 Vbias.n595 3.4105
R15771 Vbias.n598 Vbias.n597 3.4105
R15772 Vbias.n608 Vbias.n607 3.4105
R15773 Vbias.n610 Vbias.n609 3.4105
R15774 Vbias.n620 Vbias.n619 3.4105
R15775 Vbias.n622 Vbias.n621 3.4105
R15776 Vbias.n632 Vbias.n631 3.4105
R15777 Vbias.n634 Vbias.n633 3.4105
R15778 Vbias.n644 Vbias.n643 3.4105
R15779 Vbias.n646 Vbias.n645 3.4105
R15780 Vbias.n656 Vbias.n655 3.4105
R15781 Vbias.n659 Vbias.n658 3.4105
R15782 Vbias.n662 Vbias.n661 3.4105
R15783 Vbias.n529 Vbias.n528 3.4105
R15784 Vbias.n531 Vbias.n530 3.4105
R15785 Vbias.n652 Vbias.n651 3.4105
R15786 Vbias.n650 Vbias.n649 3.4105
R15787 Vbias.n640 Vbias.n639 3.4105
R15788 Vbias.n638 Vbias.n637 3.4105
R15789 Vbias.n628 Vbias.n627 3.4105
R15790 Vbias.n626 Vbias.n625 3.4105
R15791 Vbias.n616 Vbias.n615 3.4105
R15792 Vbias.n614 Vbias.n613 3.4105
R15793 Vbias.n604 Vbias.n603 3.4105
R15794 Vbias.n602 Vbias.n601 3.4105
R15795 Vbias.n592 Vbias.n591 3.4105
R15796 Vbias.n590 Vbias.n589 3.4105
R15797 Vbias.n580 Vbias.n579 3.4105
R15798 Vbias.n574 Vbias.n573 3.4105
R15799 Vbias.n571 Vbias.n570 3.4105
R15800 Vbias.n568 Vbias.n567 3.4105
R15801 Vbias.n565 Vbias.n564 3.4105
R15802 Vbias.n562 Vbias.n561 3.4105
R15803 Vbias.n559 Vbias.n558 3.4105
R15804 Vbias.n556 Vbias.n555 3.4105
R15805 Vbias.n553 Vbias.n552 3.4105
R15806 Vbias.n550 Vbias.n549 3.4105
R15807 Vbias.n547 Vbias.n546 3.4105
R15808 Vbias.n544 Vbias.n543 3.4105
R15809 Vbias.n541 Vbias.n540 3.4105
R15810 Vbias.n538 Vbias.n537 3.4105
R15811 Vbias.n535 Vbias.n534 3.4105
R15812 Vbias.n386 Vbias.n285 3.4105
R15813 Vbias.n524 Vbias.n523 3.4105
R15814 Vbias.n522 Vbias.n521 3.4105
R15815 Vbias.n519 Vbias.n518 3.4105
R15816 Vbias.n509 Vbias.n508 3.4105
R15817 Vbias.n507 Vbias.n506 3.4105
R15818 Vbias.n497 Vbias.n496 3.4105
R15819 Vbias.n495 Vbias.n494 3.4105
R15820 Vbias.n485 Vbias.n484 3.4105
R15821 Vbias.n483 Vbias.n482 3.4105
R15822 Vbias.n473 Vbias.n472 3.4105
R15823 Vbias.n471 Vbias.n470 3.4105
R15824 Vbias.n461 Vbias.n460 3.4105
R15825 Vbias.n459 Vbias.n458 3.4105
R15826 Vbias.n449 Vbias.n448 3.4105
R15827 Vbias.n447 Vbias.n446 3.4105
R15828 Vbias.n443 Vbias.n442 3.4105
R15829 Vbias.n453 Vbias.n452 3.4105
R15830 Vbias.n455 Vbias.n454 3.4105
R15831 Vbias.n465 Vbias.n464 3.4105
R15832 Vbias.n467 Vbias.n466 3.4105
R15833 Vbias.n477 Vbias.n476 3.4105
R15834 Vbias.n479 Vbias.n478 3.4105
R15835 Vbias.n489 Vbias.n488 3.4105
R15836 Vbias.n491 Vbias.n490 3.4105
R15837 Vbias.n501 Vbias.n500 3.4105
R15838 Vbias.n503 Vbias.n502 3.4105
R15839 Vbias.n513 Vbias.n512 3.4105
R15840 Vbias.n515 Vbias.n514 3.4105
R15841 Vbias.n394 Vbias.n393 3.4105
R15842 Vbias.n392 Vbias.n391 3.4105
R15843 Vbias.n384 Vbias.n383 3.4105
R15844 Vbias.n377 Vbias.n335 3.4105
R15845 Vbias.n376 Vbias.n375 3.4105
R15846 Vbias.n373 Vbias.n372 3.4105
R15847 Vbias.n370 Vbias.n369 3.4105
R15848 Vbias.n367 Vbias.n366 3.4105
R15849 Vbias.n364 Vbias.n363 3.4105
R15850 Vbias.n361 Vbias.n360 3.4105
R15851 Vbias.n358 Vbias.n357 3.4105
R15852 Vbias.n355 Vbias.n354 3.4105
R15853 Vbias.n352 Vbias.n351 3.4105
R15854 Vbias.n349 Vbias.n348 3.4105
R15855 Vbias.n346 Vbias.n345 3.4105
R15856 Vbias.n343 Vbias.n342 3.4105
R15857 Vbias.n340 Vbias.n339 3.4105
R15858 Vbias.n437 Vbias.n436 3.4105
R15859 Vbias.n434 Vbias.n433 3.4105
R15860 Vbias.n431 Vbias.n430 3.4105
R15861 Vbias.n428 Vbias.n427 3.4105
R15862 Vbias.n425 Vbias.n424 3.4105
R15863 Vbias.n422 Vbias.n421 3.4105
R15864 Vbias.n419 Vbias.n418 3.4105
R15865 Vbias.n416 Vbias.n415 3.4105
R15866 Vbias.n413 Vbias.n412 3.4105
R15867 Vbias.n410 Vbias.n409 3.4105
R15868 Vbias.n407 Vbias.n406 3.4105
R15869 Vbias.n404 Vbias.n403 3.4105
R15870 Vbias.n401 Vbias.n400 3.4105
R15871 Vbias.n398 Vbias.n397 3.4105
R15872 Vbias.n381 Vbias.n380 3.4105
R15873 Vbias.n382 Vbias.n381 2.9408
R15874 Vbias.n436 Vbias.n327 2.9408
R15875 Vbias.n917 Vbias.n916 2.9408
R15876 Vbias.n433 Vbias.n322 2.9408
R15877 Vbias.n921 Vbias.n920 2.9408
R15878 Vbias.n430 Vbias.n319 2.9408
R15879 Vbias.n927 Vbias.n926 2.9408
R15880 Vbias.n427 Vbias.n316 2.9408
R15881 Vbias.n931 Vbias.n930 2.9408
R15882 Vbias.n424 Vbias.n313 2.9408
R15883 Vbias.n937 Vbias.n936 2.9408
R15884 Vbias.n421 Vbias.n310 2.9408
R15885 Vbias.n941 Vbias.n940 2.9408
R15886 Vbias.n418 Vbias.n307 2.9408
R15887 Vbias.n947 Vbias.n946 2.9408
R15888 Vbias.n415 Vbias.n304 2.9408
R15889 Vbias.n951 Vbias.n950 2.9408
R15890 Vbias.n412 Vbias.n301 2.9408
R15891 Vbias.n957 Vbias.n956 2.9408
R15892 Vbias.n409 Vbias.n298 2.9408
R15893 Vbias.n961 Vbias.n960 2.9408
R15894 Vbias.n406 Vbias.n295 2.9408
R15895 Vbias.n967 Vbias.n966 2.9408
R15896 Vbias.n403 Vbias.n292 2.9408
R15897 Vbias.n971 Vbias.n970 2.9408
R15898 Vbias.n400 Vbias.n289 2.9408
R15899 Vbias.n977 Vbias.n976 2.9408
R15900 Vbias.n397 Vbias.n396 2.9408
R15901 Vbias.n981 Vbias.n980 2.9408
R15902 Vbias.n989 Vbias.n988 2.9408
R15903 Vbias.n912 Vbias.n54 2.9408
R15904 Vbias.n439 Vbias.n438 2.9408
R15905 Vbias.n444 Vbias.n327 2.76612
R15906 Vbias.n445 Vbias.n444 2.76612
R15907 Vbias.n445 Vbias.n272 2.76612
R15908 Vbias.n581 Vbias.n272 2.76612
R15909 Vbias.n582 Vbias.n581 2.76612
R15910 Vbias.n582 Vbias.n146 2.76612
R15911 Vbias.n776 Vbias.n146 2.76612
R15912 Vbias.n776 Vbias.n775 2.76612
R15913 Vbias.n775 Vbias.n99 2.76612
R15914 Vbias.n905 Vbias.n99 2.76612
R15915 Vbias.n906 Vbias.n905 2.76612
R15916 Vbias.n906 Vbias.n50 2.76612
R15917 Vbias.n916 Vbias.n50 2.76612
R15918 Vbias.n451 Vbias.n322 2.76612
R15919 Vbias.n451 Vbias.n450 2.76612
R15920 Vbias.n450 Vbias.n269 2.76612
R15921 Vbias.n588 Vbias.n269 2.76612
R15922 Vbias.n588 Vbias.n587 2.76612
R15923 Vbias.n587 Vbias.n149 2.76612
R15924 Vbias.n769 Vbias.n149 2.76612
R15925 Vbias.n770 Vbias.n769 2.76612
R15926 Vbias.n770 Vbias.n102 2.76612
R15927 Vbias.n898 Vbias.n102 2.76612
R15928 Vbias.n898 Vbias.n897 2.76612
R15929 Vbias.n897 Vbias.n47 2.76612
R15930 Vbias.n921 Vbias.n47 2.76612
R15931 Vbias.n456 Vbias.n319 2.76612
R15932 Vbias.n457 Vbias.n456 2.76612
R15933 Vbias.n457 Vbias.n266 2.76612
R15934 Vbias.n593 Vbias.n266 2.76612
R15935 Vbias.n594 Vbias.n593 2.76612
R15936 Vbias.n594 Vbias.n152 2.76612
R15937 Vbias.n764 Vbias.n152 2.76612
R15938 Vbias.n764 Vbias.n763 2.76612
R15939 Vbias.n763 Vbias.n105 2.76612
R15940 Vbias.n891 Vbias.n105 2.76612
R15941 Vbias.n892 Vbias.n891 2.76612
R15942 Vbias.n892 Vbias.n44 2.76612
R15943 Vbias.n926 Vbias.n44 2.76612
R15944 Vbias.n463 Vbias.n316 2.76612
R15945 Vbias.n463 Vbias.n462 2.76612
R15946 Vbias.n462 Vbias.n263 2.76612
R15947 Vbias.n600 Vbias.n263 2.76612
R15948 Vbias.n600 Vbias.n599 2.76612
R15949 Vbias.n599 Vbias.n155 2.76612
R15950 Vbias.n757 Vbias.n155 2.76612
R15951 Vbias.n758 Vbias.n757 2.76612
R15952 Vbias.n758 Vbias.n108 2.76612
R15953 Vbias.n886 Vbias.n108 2.76612
R15954 Vbias.n886 Vbias.n885 2.76612
R15955 Vbias.n885 Vbias.n41 2.76612
R15956 Vbias.n931 Vbias.n41 2.76612
R15957 Vbias.n468 Vbias.n313 2.76612
R15958 Vbias.n469 Vbias.n468 2.76612
R15959 Vbias.n469 Vbias.n260 2.76612
R15960 Vbias.n605 Vbias.n260 2.76612
R15961 Vbias.n606 Vbias.n605 2.76612
R15962 Vbias.n606 Vbias.n158 2.76612
R15963 Vbias.n752 Vbias.n158 2.76612
R15964 Vbias.n752 Vbias.n751 2.76612
R15965 Vbias.n751 Vbias.n111 2.76612
R15966 Vbias.n879 Vbias.n111 2.76612
R15967 Vbias.n880 Vbias.n879 2.76612
R15968 Vbias.n880 Vbias.n38 2.76612
R15969 Vbias.n936 Vbias.n38 2.76612
R15970 Vbias.n475 Vbias.n310 2.76612
R15971 Vbias.n475 Vbias.n474 2.76612
R15972 Vbias.n474 Vbias.n257 2.76612
R15973 Vbias.n612 Vbias.n257 2.76612
R15974 Vbias.n612 Vbias.n611 2.76612
R15975 Vbias.n611 Vbias.n161 2.76612
R15976 Vbias.n745 Vbias.n161 2.76612
R15977 Vbias.n746 Vbias.n745 2.76612
R15978 Vbias.n746 Vbias.n114 2.76612
R15979 Vbias.n874 Vbias.n114 2.76612
R15980 Vbias.n874 Vbias.n873 2.76612
R15981 Vbias.n873 Vbias.n35 2.76612
R15982 Vbias.n941 Vbias.n35 2.76612
R15983 Vbias.n480 Vbias.n307 2.76612
R15984 Vbias.n481 Vbias.n480 2.76612
R15985 Vbias.n481 Vbias.n254 2.76612
R15986 Vbias.n617 Vbias.n254 2.76612
R15987 Vbias.n618 Vbias.n617 2.76612
R15988 Vbias.n618 Vbias.n164 2.76612
R15989 Vbias.n740 Vbias.n164 2.76612
R15990 Vbias.n740 Vbias.n739 2.76612
R15991 Vbias.n739 Vbias.n117 2.76612
R15992 Vbias.n867 Vbias.n117 2.76612
R15993 Vbias.n868 Vbias.n867 2.76612
R15994 Vbias.n868 Vbias.n32 2.76612
R15995 Vbias.n946 Vbias.n32 2.76612
R15996 Vbias.n487 Vbias.n304 2.76612
R15997 Vbias.n487 Vbias.n486 2.76612
R15998 Vbias.n486 Vbias.n251 2.76612
R15999 Vbias.n624 Vbias.n251 2.76612
R16000 Vbias.n624 Vbias.n623 2.76612
R16001 Vbias.n623 Vbias.n167 2.76612
R16002 Vbias.n733 Vbias.n167 2.76612
R16003 Vbias.n734 Vbias.n733 2.76612
R16004 Vbias.n734 Vbias.n120 2.76612
R16005 Vbias.n862 Vbias.n120 2.76612
R16006 Vbias.n862 Vbias.n861 2.76612
R16007 Vbias.n861 Vbias.n29 2.76612
R16008 Vbias.n951 Vbias.n29 2.76612
R16009 Vbias.n492 Vbias.n301 2.76612
R16010 Vbias.n493 Vbias.n492 2.76612
R16011 Vbias.n493 Vbias.n248 2.76612
R16012 Vbias.n629 Vbias.n248 2.76612
R16013 Vbias.n630 Vbias.n629 2.76612
R16014 Vbias.n630 Vbias.n170 2.76612
R16015 Vbias.n728 Vbias.n170 2.76612
R16016 Vbias.n728 Vbias.n727 2.76612
R16017 Vbias.n727 Vbias.n123 2.76612
R16018 Vbias.n855 Vbias.n123 2.76612
R16019 Vbias.n856 Vbias.n855 2.76612
R16020 Vbias.n856 Vbias.n26 2.76612
R16021 Vbias.n956 Vbias.n26 2.76612
R16022 Vbias.n499 Vbias.n298 2.76612
R16023 Vbias.n499 Vbias.n498 2.76612
R16024 Vbias.n498 Vbias.n245 2.76612
R16025 Vbias.n636 Vbias.n245 2.76612
R16026 Vbias.n636 Vbias.n635 2.76612
R16027 Vbias.n635 Vbias.n173 2.76612
R16028 Vbias.n721 Vbias.n173 2.76612
R16029 Vbias.n722 Vbias.n721 2.76612
R16030 Vbias.n722 Vbias.n126 2.76612
R16031 Vbias.n850 Vbias.n126 2.76612
R16032 Vbias.n850 Vbias.n849 2.76612
R16033 Vbias.n849 Vbias.n23 2.76612
R16034 Vbias.n961 Vbias.n23 2.76612
R16035 Vbias.n504 Vbias.n295 2.76612
R16036 Vbias.n505 Vbias.n504 2.76612
R16037 Vbias.n505 Vbias.n242 2.76612
R16038 Vbias.n641 Vbias.n242 2.76612
R16039 Vbias.n642 Vbias.n641 2.76612
R16040 Vbias.n642 Vbias.n176 2.76612
R16041 Vbias.n716 Vbias.n176 2.76612
R16042 Vbias.n716 Vbias.n715 2.76612
R16043 Vbias.n715 Vbias.n129 2.76612
R16044 Vbias.n843 Vbias.n129 2.76612
R16045 Vbias.n844 Vbias.n843 2.76612
R16046 Vbias.n844 Vbias.n20 2.76612
R16047 Vbias.n966 Vbias.n20 2.76612
R16048 Vbias.n511 Vbias.n292 2.76612
R16049 Vbias.n511 Vbias.n510 2.76612
R16050 Vbias.n510 Vbias.n239 2.76612
R16051 Vbias.n648 Vbias.n239 2.76612
R16052 Vbias.n648 Vbias.n647 2.76612
R16053 Vbias.n647 Vbias.n179 2.76612
R16054 Vbias.n709 Vbias.n179 2.76612
R16055 Vbias.n710 Vbias.n709 2.76612
R16056 Vbias.n710 Vbias.n132 2.76612
R16057 Vbias.n838 Vbias.n132 2.76612
R16058 Vbias.n838 Vbias.n837 2.76612
R16059 Vbias.n837 Vbias.n17 2.76612
R16060 Vbias.n971 Vbias.n17 2.76612
R16061 Vbias.n516 Vbias.n289 2.76612
R16062 Vbias.n517 Vbias.n516 2.76612
R16063 Vbias.n517 Vbias.n236 2.76612
R16064 Vbias.n653 Vbias.n236 2.76612
R16065 Vbias.n654 Vbias.n653 2.76612
R16066 Vbias.n654 Vbias.n182 2.76612
R16067 Vbias.n704 Vbias.n182 2.76612
R16068 Vbias.n704 Vbias.n703 2.76612
R16069 Vbias.n703 Vbias.n135 2.76612
R16070 Vbias.n831 Vbias.n135 2.76612
R16071 Vbias.n832 Vbias.n831 2.76612
R16072 Vbias.n832 Vbias.n12 2.76612
R16073 Vbias.n976 Vbias.n12 2.76612
R16074 Vbias.n396 Vbias.n395 2.76612
R16075 Vbias.n395 Vbias.n281 2.76612
R16076 Vbias.n533 Vbias.n281 2.76612
R16077 Vbias.n533 Vbias.n532 2.76612
R16078 Vbias.n532 Vbias.n232 2.76612
R16079 Vbias.n688 Vbias.n232 2.76612
R16080 Vbias.n688 Vbias.n687 2.76612
R16081 Vbias.n687 Vbias.n138 2.76612
R16082 Vbias.n825 Vbias.n138 2.76612
R16083 Vbias.n826 Vbias.n825 2.76612
R16084 Vbias.n826 Vbias.n7 2.76612
R16085 Vbias.n982 Vbias.n7 2.76612
R16086 Vbias.n982 Vbias.n981 2.76612
R16087 Vbias.n912 Vbias.n911 2.76612
R16088 Vbias.n988 Vbias.n987 2.76612
R16089 Vbias.n987 Vbias.n4 2.76612
R16090 Vbias.n911 Vbias.n910 2.76612
R16091 Vbias.n910 Vbias.n96 2.76612
R16092 Vbias.n674 Vbias.n4 2.76612
R16093 Vbias.n674 Vbias.n185 2.76612
R16094 Vbias.n782 Vbias.n96 2.76612
R16095 Vbias.n782 Vbias.n781 2.76612
R16096 Vbias.n695 Vbias.n185 2.76612
R16097 Vbias.n695 Vbias.n694 2.76612
R16098 Vbias.n781 Vbias.n780 2.76612
R16099 Vbias.n780 Vbias.n143 2.76612
R16100 Vbias.n694 Vbias.n693 2.76612
R16101 Vbias.n693 Vbias.n188 2.76612
R16102 Vbias.n277 Vbias.n143 2.76612
R16103 Vbias.n577 Vbias.n277 2.76612
R16104 Vbias.n527 Vbias.n188 2.76612
R16105 Vbias.n527 Vbias.n526 2.76612
R16106 Vbias.n577 Vbias.n576 2.76612
R16107 Vbias.n576 Vbias.n278 2.76612
R16108 Vbias.n526 Vbias.n525 2.76612
R16109 Vbias.n525 Vbias.n286 2.76612
R16110 Vbias.n440 Vbias.n278 2.76612
R16111 Vbias.n440 Vbias.n439 2.76612
R16112 Vbias.n382 Vbias.n286 2.76612
R16113 Vbias.n996 Vbias.n994 2.09636
R16114 Vbias Vbias.n337 1.6647
R16115 Vbias Vbias.n389 1.6647
R16116 Vbias.n387 Vbias 1.6647
R16117 Vbias.n663 Vbias 1.6647
R16118 Vbias Vbias.n683 1.6647
R16119 Vbias.n681 Vbias 1.6647
R16120 Vbias.n672 Vbias 1.6647
R16121 Vbias Vbias.n0 1.6647
R16122 Vbias.n991 Vbias 1.6647
R16123 Vbias.n665 Vbias 1.6647
R16124 Vbias.n677 Vbias 1.6647
R16125 Vbias.n682 Vbias 1.6647
R16126 Vbias.n664 Vbias 1.6647
R16127 Vbias Vbias.n234 1.6647
R16128 Vbias.n388 Vbias 1.6647
R16129 Vbias.n385 Vbias 1.6647
R16130 Vbias.n997 Vbias 1.34721
R16131 Vbias Vbias.n996 0.752103
R16132 Vbias.n997 Vbias.n991 0.5692
R16133 Vbias.n996 Vbias.n995 0.515506
R16134 Vbias.n385 Vbias.n337 0.410967
R16135 Vbias.n389 Vbias.n385 0.410967
R16136 Vbias.n389 Vbias.n388 0.410967
R16137 Vbias.n388 Vbias.n387 0.410967
R16138 Vbias.n387 Vbias.n234 0.410967
R16139 Vbias.n663 Vbias.n234 0.410967
R16140 Vbias.n664 Vbias.n663 0.410967
R16141 Vbias.n683 Vbias.n664 0.410967
R16142 Vbias.n683 Vbias.n682 0.410967
R16143 Vbias.n682 Vbias.n681 0.410967
R16144 Vbias.n681 Vbias.n677 0.410967
R16145 Vbias.n677 Vbias.n672 0.410967
R16146 Vbias.n672 Vbias.n665 0.410967
R16147 Vbias.n665 Vbias.n0 0.410967
R16148 Vbias.n991 Vbias.n0 0.410967
R16149 Vbias.n337 Vbias 0.383811
R16150 Vbias.n990 Vbias 0.252372
R16151 Vbias.n979 Vbias 0.252372
R16152 Vbias.n978 Vbias 0.252372
R16153 Vbias.n969 Vbias 0.252372
R16154 Vbias.n968 Vbias 0.252372
R16155 Vbias.n959 Vbias 0.252372
R16156 Vbias.n958 Vbias 0.252372
R16157 Vbias.n949 Vbias 0.252372
R16158 Vbias.n948 Vbias 0.252372
R16159 Vbias.n939 Vbias 0.252372
R16160 Vbias.n938 Vbias 0.252372
R16161 Vbias.n929 Vbias 0.252372
R16162 Vbias.n928 Vbias 0.252372
R16163 Vbias.n919 Vbias 0.252372
R16164 Vbias.n918 Vbias 0.252372
R16165 Vbias.n914 Vbias 0.252372
R16166 Vbias.n923 Vbias 0.252372
R16167 Vbias.n924 Vbias 0.252372
R16168 Vbias.n933 Vbias 0.252372
R16169 Vbias.n934 Vbias 0.252372
R16170 Vbias.n943 Vbias 0.252372
R16171 Vbias.n944 Vbias 0.252372
R16172 Vbias.n953 Vbias 0.252372
R16173 Vbias.n954 Vbias 0.252372
R16174 Vbias.n963 Vbias 0.252372
R16175 Vbias.n964 Vbias 0.252372
R16176 Vbias.n973 Vbias 0.252372
R16177 Vbias.n974 Vbias 0.252372
R16178 Vbias Vbias.n15 0.252372
R16179 Vbias Vbias.n14 0.252372
R16180 Vbias.n985 Vbias 0.252372
R16181 Vbias.n984 Vbias 0.252372
R16182 Vbias Vbias.n58 0.252372
R16183 Vbias Vbias.n61 0.252372
R16184 Vbias Vbias.n64 0.252372
R16185 Vbias Vbias.n67 0.252372
R16186 Vbias Vbias.n70 0.252372
R16187 Vbias Vbias.n73 0.252372
R16188 Vbias Vbias.n76 0.252372
R16189 Vbias Vbias.n79 0.252372
R16190 Vbias Vbias.n82 0.252372
R16191 Vbias Vbias.n85 0.252372
R16192 Vbias Vbias.n88 0.252372
R16193 Vbias Vbias.n91 0.252372
R16194 Vbias Vbias.n94 0.252372
R16195 Vbias Vbias.n908 0.252372
R16196 Vbias.n895 Vbias 0.252372
R16197 Vbias Vbias.n894 0.252372
R16198 Vbias.n883 Vbias 0.252372
R16199 Vbias Vbias.n882 0.252372
R16200 Vbias.n871 Vbias 0.252372
R16201 Vbias Vbias.n870 0.252372
R16202 Vbias.n859 Vbias 0.252372
R16203 Vbias Vbias.n858 0.252372
R16204 Vbias.n847 Vbias 0.252372
R16205 Vbias Vbias.n846 0.252372
R16206 Vbias.n835 Vbias 0.252372
R16207 Vbias Vbias.n834 0.252372
R16208 Vbias.n668 Vbias 0.252372
R16209 Vbias.n671 Vbias 0.252372
R16210 Vbias.n676 Vbias 0.252372
R16211 Vbias Vbias.n828 0.252372
R16212 Vbias.n829 Vbias 0.252372
R16213 Vbias Vbias.n840 0.252372
R16214 Vbias.n841 Vbias 0.252372
R16215 Vbias Vbias.n852 0.252372
R16216 Vbias.n853 Vbias 0.252372
R16217 Vbias Vbias.n864 0.252372
R16218 Vbias.n865 Vbias 0.252372
R16219 Vbias Vbias.n876 0.252372
R16220 Vbias.n877 Vbias 0.252372
R16221 Vbias Vbias.n888 0.252372
R16222 Vbias.n889 Vbias 0.252372
R16223 Vbias Vbias.n900 0.252372
R16224 Vbias.n903 Vbias 0.252372
R16225 Vbias.n786 Vbias 0.252372
R16226 Vbias.n789 Vbias 0.252372
R16227 Vbias.n792 Vbias 0.252372
R16228 Vbias.n795 Vbias 0.252372
R16229 Vbias.n798 Vbias 0.252372
R16230 Vbias.n801 Vbias 0.252372
R16231 Vbias.n804 Vbias 0.252372
R16232 Vbias.n807 Vbias 0.252372
R16233 Vbias.n810 Vbias 0.252372
R16234 Vbias.n813 Vbias 0.252372
R16235 Vbias.n816 Vbias 0.252372
R16236 Vbias.n819 Vbias 0.252372
R16237 Vbias.n822 Vbias 0.252372
R16238 Vbias.n823 Vbias 0.252372
R16239 Vbias.n680 Vbias 0.252372
R16240 Vbias Vbias.n697 0.252372
R16241 Vbias Vbias.n700 0.252372
R16242 Vbias.n701 Vbias 0.252372
R16243 Vbias Vbias.n712 0.252372
R16244 Vbias.n713 Vbias 0.252372
R16245 Vbias Vbias.n724 0.252372
R16246 Vbias.n725 Vbias 0.252372
R16247 Vbias Vbias.n736 0.252372
R16248 Vbias.n737 Vbias 0.252372
R16249 Vbias Vbias.n748 0.252372
R16250 Vbias.n749 Vbias 0.252372
R16251 Vbias Vbias.n760 0.252372
R16252 Vbias.n761 Vbias 0.252372
R16253 Vbias Vbias.n772 0.252372
R16254 Vbias.n773 Vbias 0.252372
R16255 Vbias Vbias.n778 0.252372
R16256 Vbias.n767 Vbias 0.252372
R16257 Vbias Vbias.n766 0.252372
R16258 Vbias.n755 Vbias 0.252372
R16259 Vbias Vbias.n754 0.252372
R16260 Vbias.n743 Vbias 0.252372
R16261 Vbias Vbias.n742 0.252372
R16262 Vbias.n731 Vbias 0.252372
R16263 Vbias Vbias.n730 0.252372
R16264 Vbias.n719 Vbias 0.252372
R16265 Vbias Vbias.n718 0.252372
R16266 Vbias.n707 Vbias 0.252372
R16267 Vbias Vbias.n706 0.252372
R16268 Vbias.n685 Vbias 0.252372
R16269 Vbias Vbias.n684 0.252372
R16270 Vbias.n691 Vbias 0.252372
R16271 Vbias.n690 Vbias 0.252372
R16272 Vbias.n230 Vbias 0.252372
R16273 Vbias.n227 Vbias 0.252372
R16274 Vbias.n224 Vbias 0.252372
R16275 Vbias.n221 Vbias 0.252372
R16276 Vbias.n218 Vbias 0.252372
R16277 Vbias.n215 Vbias 0.252372
R16278 Vbias.n212 Vbias 0.252372
R16279 Vbias.n209 Vbias 0.252372
R16280 Vbias.n206 Vbias 0.252372
R16281 Vbias.n203 Vbias 0.252372
R16282 Vbias.n200 Vbias 0.252372
R16283 Vbias.n197 Vbias 0.252372
R16284 Vbias.n194 Vbias 0.252372
R16285 Vbias.n584 Vbias 0.252372
R16286 Vbias.n585 Vbias 0.252372
R16287 Vbias.n596 Vbias 0.252372
R16288 Vbias.n597 Vbias 0.252372
R16289 Vbias.n608 Vbias 0.252372
R16290 Vbias.n609 Vbias 0.252372
R16291 Vbias.n620 Vbias 0.252372
R16292 Vbias.n621 Vbias 0.252372
R16293 Vbias.n632 Vbias 0.252372
R16294 Vbias.n633 Vbias 0.252372
R16295 Vbias.n644 Vbias 0.252372
R16296 Vbias.n645 Vbias 0.252372
R16297 Vbias.n656 Vbias 0.252372
R16298 Vbias.n659 Vbias 0.252372
R16299 Vbias.n662 Vbias 0.252372
R16300 Vbias Vbias.n529 0.252372
R16301 Vbias.n530 Vbias 0.252372
R16302 Vbias.n651 Vbias 0.252372
R16303 Vbias.n650 Vbias 0.252372
R16304 Vbias.n639 Vbias 0.252372
R16305 Vbias.n638 Vbias 0.252372
R16306 Vbias.n627 Vbias 0.252372
R16307 Vbias.n626 Vbias 0.252372
R16308 Vbias.n615 Vbias 0.252372
R16309 Vbias.n614 Vbias 0.252372
R16310 Vbias.n603 Vbias 0.252372
R16311 Vbias.n602 Vbias 0.252372
R16312 Vbias.n591 Vbias 0.252372
R16313 Vbias.n590 Vbias 0.252372
R16314 Vbias.n579 Vbias 0.252372
R16315 Vbias Vbias.n574 0.252372
R16316 Vbias Vbias.n571 0.252372
R16317 Vbias Vbias.n568 0.252372
R16318 Vbias Vbias.n565 0.252372
R16319 Vbias Vbias.n562 0.252372
R16320 Vbias Vbias.n559 0.252372
R16321 Vbias Vbias.n556 0.252372
R16322 Vbias Vbias.n553 0.252372
R16323 Vbias Vbias.n550 0.252372
R16324 Vbias Vbias.n547 0.252372
R16325 Vbias Vbias.n544 0.252372
R16326 Vbias Vbias.n541 0.252372
R16327 Vbias Vbias.n538 0.252372
R16328 Vbias Vbias.n535 0.252372
R16329 Vbias.n386 Vbias 0.252372
R16330 Vbias.n523 Vbias 0.252372
R16331 Vbias.n522 Vbias 0.252372
R16332 Vbias.n519 Vbias 0.252372
R16333 Vbias.n508 Vbias 0.252372
R16334 Vbias.n507 Vbias 0.252372
R16335 Vbias.n496 Vbias 0.252372
R16336 Vbias.n495 Vbias 0.252372
R16337 Vbias.n484 Vbias 0.252372
R16338 Vbias.n483 Vbias 0.252372
R16339 Vbias.n472 Vbias 0.252372
R16340 Vbias.n471 Vbias 0.252372
R16341 Vbias.n460 Vbias 0.252372
R16342 Vbias.n459 Vbias 0.252372
R16343 Vbias.n448 Vbias 0.252372
R16344 Vbias.n447 Vbias 0.252372
R16345 Vbias.n442 Vbias 0.252372
R16346 Vbias.n453 Vbias 0.252372
R16347 Vbias.n454 Vbias 0.252372
R16348 Vbias.n465 Vbias 0.252372
R16349 Vbias.n466 Vbias 0.252372
R16350 Vbias.n477 Vbias 0.252372
R16351 Vbias.n478 Vbias 0.252372
R16352 Vbias.n489 Vbias 0.252372
R16353 Vbias.n490 Vbias 0.252372
R16354 Vbias.n501 Vbias 0.252372
R16355 Vbias.n502 Vbias 0.252372
R16356 Vbias.n513 Vbias 0.252372
R16357 Vbias.n514 Vbias 0.252372
R16358 Vbias.n393 Vbias 0.252372
R16359 Vbias Vbias.n392 0.252372
R16360 Vbias.n384 Vbias 0.252372
R16361 Vbias.n377 Vbias 0.252372
R16362 Vbias.n376 Vbias 0.252372
R16363 Vbias.n373 Vbias 0.252372
R16364 Vbias.n370 Vbias 0.252372
R16365 Vbias.n367 Vbias 0.252372
R16366 Vbias.n364 Vbias 0.252372
R16367 Vbias.n361 Vbias 0.252372
R16368 Vbias.n358 Vbias 0.252372
R16369 Vbias.n355 Vbias 0.252372
R16370 Vbias.n352 Vbias 0.252372
R16371 Vbias.n349 Vbias 0.252372
R16372 Vbias.n346 Vbias 0.252372
R16373 Vbias.n343 Vbias 0.252372
R16374 Vbias.n340 Vbias 0.252372
R16375 Vbias Vbias.n437 0.252372
R16376 Vbias Vbias.n434 0.252372
R16377 Vbias Vbias.n431 0.252372
R16378 Vbias Vbias.n428 0.252372
R16379 Vbias Vbias.n425 0.252372
R16380 Vbias Vbias.n422 0.252372
R16381 Vbias Vbias.n419 0.252372
R16382 Vbias Vbias.n416 0.252372
R16383 Vbias Vbias.n413 0.252372
R16384 Vbias Vbias.n410 0.252372
R16385 Vbias Vbias.n407 0.252372
R16386 Vbias Vbias.n404 0.252372
R16387 Vbias Vbias.n401 0.252372
R16388 Vbias Vbias.n398 0.252372
R16389 Vbias.n380 Vbias 0.252372
R16390 Vbias Vbias.n997 0.237067
R16391 Vbias.n339 Vbias.n327 0.175179
R16392 Vbias.n444 Vbias.n443 0.175179
R16393 Vbias.n446 Vbias.n445 0.175179
R16394 Vbias.n573 Vbias.n272 0.175179
R16395 Vbias.n581 Vbias.n580 0.175179
R16396 Vbias.n583 Vbias.n582 0.175179
R16397 Vbias.n193 Vbias.n146 0.175179
R16398 Vbias.n777 Vbias.n776 0.175179
R16399 Vbias.n775 Vbias.n774 0.175179
R16400 Vbias.n785 Vbias.n99 0.175179
R16401 Vbias.n905 Vbias.n904 0.175179
R16402 Vbias.n907 Vbias.n906 0.175179
R16403 Vbias.n93 Vbias.n50 0.175179
R16404 Vbias.n916 Vbias.n915 0.175179
R16405 Vbias.n342 Vbias.n322 0.175179
R16406 Vbias.n452 Vbias.n451 0.175179
R16407 Vbias.n450 Vbias.n449 0.175179
R16408 Vbias.n570 Vbias.n269 0.175179
R16409 Vbias.n589 Vbias.n588 0.175179
R16410 Vbias.n587 Vbias.n586 0.175179
R16411 Vbias.n196 Vbias.n149 0.175179
R16412 Vbias.n769 Vbias.n768 0.175179
R16413 Vbias.n771 Vbias.n770 0.175179
R16414 Vbias.n788 Vbias.n102 0.175179
R16415 Vbias.n899 Vbias.n898 0.175179
R16416 Vbias.n897 Vbias.n896 0.175179
R16417 Vbias.n90 Vbias.n47 0.175179
R16418 Vbias.n922 Vbias.n921 0.175179
R16419 Vbias.n345 Vbias.n319 0.175179
R16420 Vbias.n456 Vbias.n455 0.175179
R16421 Vbias.n458 Vbias.n457 0.175179
R16422 Vbias.n567 Vbias.n266 0.175179
R16423 Vbias.n593 Vbias.n592 0.175179
R16424 Vbias.n595 Vbias.n594 0.175179
R16425 Vbias.n199 Vbias.n152 0.175179
R16426 Vbias.n765 Vbias.n764 0.175179
R16427 Vbias.n763 Vbias.n762 0.175179
R16428 Vbias.n791 Vbias.n105 0.175179
R16429 Vbias.n891 Vbias.n890 0.175179
R16430 Vbias.n893 Vbias.n892 0.175179
R16431 Vbias.n87 Vbias.n44 0.175179
R16432 Vbias.n926 Vbias.n925 0.175179
R16433 Vbias.n348 Vbias.n316 0.175179
R16434 Vbias.n464 Vbias.n463 0.175179
R16435 Vbias.n462 Vbias.n461 0.175179
R16436 Vbias.n564 Vbias.n263 0.175179
R16437 Vbias.n601 Vbias.n600 0.175179
R16438 Vbias.n599 Vbias.n598 0.175179
R16439 Vbias.n202 Vbias.n155 0.175179
R16440 Vbias.n757 Vbias.n756 0.175179
R16441 Vbias.n759 Vbias.n758 0.175179
R16442 Vbias.n794 Vbias.n108 0.175179
R16443 Vbias.n887 Vbias.n886 0.175179
R16444 Vbias.n885 Vbias.n884 0.175179
R16445 Vbias.n84 Vbias.n41 0.175179
R16446 Vbias.n932 Vbias.n931 0.175179
R16447 Vbias.n351 Vbias.n313 0.175179
R16448 Vbias.n468 Vbias.n467 0.175179
R16449 Vbias.n470 Vbias.n469 0.175179
R16450 Vbias.n561 Vbias.n260 0.175179
R16451 Vbias.n605 Vbias.n604 0.175179
R16452 Vbias.n607 Vbias.n606 0.175179
R16453 Vbias.n205 Vbias.n158 0.175179
R16454 Vbias.n753 Vbias.n752 0.175179
R16455 Vbias.n751 Vbias.n750 0.175179
R16456 Vbias.n797 Vbias.n111 0.175179
R16457 Vbias.n879 Vbias.n878 0.175179
R16458 Vbias.n881 Vbias.n880 0.175179
R16459 Vbias.n81 Vbias.n38 0.175179
R16460 Vbias.n936 Vbias.n935 0.175179
R16461 Vbias.n354 Vbias.n310 0.175179
R16462 Vbias.n476 Vbias.n475 0.175179
R16463 Vbias.n474 Vbias.n473 0.175179
R16464 Vbias.n558 Vbias.n257 0.175179
R16465 Vbias.n613 Vbias.n612 0.175179
R16466 Vbias.n611 Vbias.n610 0.175179
R16467 Vbias.n208 Vbias.n161 0.175179
R16468 Vbias.n745 Vbias.n744 0.175179
R16469 Vbias.n747 Vbias.n746 0.175179
R16470 Vbias.n800 Vbias.n114 0.175179
R16471 Vbias.n875 Vbias.n874 0.175179
R16472 Vbias.n873 Vbias.n872 0.175179
R16473 Vbias.n78 Vbias.n35 0.175179
R16474 Vbias.n942 Vbias.n941 0.175179
R16475 Vbias.n357 Vbias.n307 0.175179
R16476 Vbias.n480 Vbias.n479 0.175179
R16477 Vbias.n482 Vbias.n481 0.175179
R16478 Vbias.n555 Vbias.n254 0.175179
R16479 Vbias.n617 Vbias.n616 0.175179
R16480 Vbias.n619 Vbias.n618 0.175179
R16481 Vbias.n211 Vbias.n164 0.175179
R16482 Vbias.n741 Vbias.n740 0.175179
R16483 Vbias.n739 Vbias.n738 0.175179
R16484 Vbias.n803 Vbias.n117 0.175179
R16485 Vbias.n867 Vbias.n866 0.175179
R16486 Vbias.n869 Vbias.n868 0.175179
R16487 Vbias.n75 Vbias.n32 0.175179
R16488 Vbias.n946 Vbias.n945 0.175179
R16489 Vbias.n360 Vbias.n304 0.175179
R16490 Vbias.n488 Vbias.n487 0.175179
R16491 Vbias.n486 Vbias.n485 0.175179
R16492 Vbias.n552 Vbias.n251 0.175179
R16493 Vbias.n625 Vbias.n624 0.175179
R16494 Vbias.n623 Vbias.n622 0.175179
R16495 Vbias.n214 Vbias.n167 0.175179
R16496 Vbias.n733 Vbias.n732 0.175179
R16497 Vbias.n735 Vbias.n734 0.175179
R16498 Vbias.n806 Vbias.n120 0.175179
R16499 Vbias.n863 Vbias.n862 0.175179
R16500 Vbias.n861 Vbias.n860 0.175179
R16501 Vbias.n72 Vbias.n29 0.175179
R16502 Vbias.n952 Vbias.n951 0.175179
R16503 Vbias.n363 Vbias.n301 0.175179
R16504 Vbias.n492 Vbias.n491 0.175179
R16505 Vbias.n494 Vbias.n493 0.175179
R16506 Vbias.n549 Vbias.n248 0.175179
R16507 Vbias.n629 Vbias.n628 0.175179
R16508 Vbias.n631 Vbias.n630 0.175179
R16509 Vbias.n217 Vbias.n170 0.175179
R16510 Vbias.n729 Vbias.n728 0.175179
R16511 Vbias.n727 Vbias.n726 0.175179
R16512 Vbias.n809 Vbias.n123 0.175179
R16513 Vbias.n855 Vbias.n854 0.175179
R16514 Vbias.n857 Vbias.n856 0.175179
R16515 Vbias.n69 Vbias.n26 0.175179
R16516 Vbias.n956 Vbias.n955 0.175179
R16517 Vbias.n366 Vbias.n298 0.175179
R16518 Vbias.n500 Vbias.n499 0.175179
R16519 Vbias.n498 Vbias.n497 0.175179
R16520 Vbias.n546 Vbias.n245 0.175179
R16521 Vbias.n637 Vbias.n636 0.175179
R16522 Vbias.n635 Vbias.n634 0.175179
R16523 Vbias.n220 Vbias.n173 0.175179
R16524 Vbias.n721 Vbias.n720 0.175179
R16525 Vbias.n723 Vbias.n722 0.175179
R16526 Vbias.n812 Vbias.n126 0.175179
R16527 Vbias.n851 Vbias.n850 0.175179
R16528 Vbias.n849 Vbias.n848 0.175179
R16529 Vbias.n66 Vbias.n23 0.175179
R16530 Vbias.n962 Vbias.n961 0.175179
R16531 Vbias.n369 Vbias.n295 0.175179
R16532 Vbias.n504 Vbias.n503 0.175179
R16533 Vbias.n506 Vbias.n505 0.175179
R16534 Vbias.n543 Vbias.n242 0.175179
R16535 Vbias.n641 Vbias.n640 0.175179
R16536 Vbias.n643 Vbias.n642 0.175179
R16537 Vbias.n223 Vbias.n176 0.175179
R16538 Vbias.n717 Vbias.n716 0.175179
R16539 Vbias.n715 Vbias.n714 0.175179
R16540 Vbias.n815 Vbias.n129 0.175179
R16541 Vbias.n843 Vbias.n842 0.175179
R16542 Vbias.n845 Vbias.n844 0.175179
R16543 Vbias.n63 Vbias.n20 0.175179
R16544 Vbias.n966 Vbias.n965 0.175179
R16545 Vbias.n372 Vbias.n292 0.175179
R16546 Vbias.n512 Vbias.n511 0.175179
R16547 Vbias.n510 Vbias.n509 0.175179
R16548 Vbias.n540 Vbias.n239 0.175179
R16549 Vbias.n649 Vbias.n648 0.175179
R16550 Vbias.n647 Vbias.n646 0.175179
R16551 Vbias.n226 Vbias.n179 0.175179
R16552 Vbias.n709 Vbias.n708 0.175179
R16553 Vbias.n711 Vbias.n710 0.175179
R16554 Vbias.n818 Vbias.n132 0.175179
R16555 Vbias.n839 Vbias.n838 0.175179
R16556 Vbias.n837 Vbias.n836 0.175179
R16557 Vbias.n60 Vbias.n17 0.175179
R16558 Vbias.n972 Vbias.n971 0.175179
R16559 Vbias.n375 Vbias.n289 0.175179
R16560 Vbias.n516 Vbias.n515 0.175179
R16561 Vbias.n518 Vbias.n517 0.175179
R16562 Vbias.n537 Vbias.n236 0.175179
R16563 Vbias.n653 Vbias.n652 0.175179
R16564 Vbias.n655 Vbias.n654 0.175179
R16565 Vbias.n229 Vbias.n182 0.175179
R16566 Vbias.n705 Vbias.n704 0.175179
R16567 Vbias.n703 Vbias.n702 0.175179
R16568 Vbias.n821 Vbias.n135 0.175179
R16569 Vbias.n831 Vbias.n830 0.175179
R16570 Vbias.n833 Vbias.n832 0.175179
R16571 Vbias.n57 Vbias.n12 0.175179
R16572 Vbias.n976 Vbias.n975 0.175179
R16573 Vbias.n396 Vbias.n335 0.175179
R16574 Vbias.n395 Vbias.n394 0.175179
R16575 Vbias.n521 Vbias.n281 0.175179
R16576 Vbias.n534 Vbias.n533 0.175179
R16577 Vbias.n532 Vbias.n531 0.175179
R16578 Vbias.n658 Vbias.n232 0.175179
R16579 Vbias.n689 Vbias.n688 0.175179
R16580 Vbias.n687 Vbias.n686 0.175179
R16581 Vbias.n699 Vbias.n138 0.175179
R16582 Vbias.n825 Vbias.n824 0.175179
R16583 Vbias.n827 Vbias.n826 0.175179
R16584 Vbias.n667 Vbias.n7 0.175179
R16585 Vbias.n983 Vbias.n982 0.175179
R16586 Vbias.n981 Vbias.n9 0.175179
R16587 Vbias.n913 Vbias.n912 0.175179
R16588 Vbias.n988 Vbias.n3 0.175179
R16589 Vbias.n987 Vbias.n986 0.175179
R16590 Vbias.n911 Vbias.n95 0.175179
R16591 Vbias.n910 Vbias.n909 0.175179
R16592 Vbias.n670 Vbias.n4 0.175179
R16593 Vbias.n675 Vbias.n674 0.175179
R16594 Vbias.n902 Vbias.n96 0.175179
R16595 Vbias.n783 Vbias.n782 0.175179
R16596 Vbias.n679 Vbias.n185 0.175179
R16597 Vbias.n696 Vbias.n695 0.175179
R16598 Vbias.n781 Vbias.n142 0.175179
R16599 Vbias.n780 Vbias.n779 0.175179
R16600 Vbias.n694 Vbias.n187 0.175179
R16601 Vbias.n693 Vbias.n692 0.175179
R16602 Vbias.n191 Vbias.n143 0.175179
R16603 Vbias.n277 Vbias.n276 0.175179
R16604 Vbias.n661 Vbias.n188 0.175179
R16605 Vbias.n528 Vbias.n527 0.175179
R16606 Vbias.n578 Vbias.n577 0.175179
R16607 Vbias.n576 Vbias.n575 0.175179
R16608 Vbias.n526 Vbias.n285 0.175179
R16609 Vbias.n525 Vbias.n524 0.175179
R16610 Vbias.n325 Vbias.n278 0.175179
R16611 Vbias.n441 Vbias.n440 0.175179
R16612 Vbias.n391 Vbias.n286 0.175179
R16613 Vbias.n383 Vbias.n382 0.175179
R16614 Vbias.n439 Vbias.n331 0.175179
R16615 Vbias.n392 Vbias 0.0972718
R16616 Vbias Vbias.n386 0.0972718
R16617 Vbias Vbias.n662 0.0972718
R16618 Vbias.n684 Vbias 0.0972718
R16619 Vbias Vbias.n680 0.0972718
R16620 Vbias Vbias.n671 0.0972718
R16621 Vbias.n14 Vbias 0.0972718
R16622 Vbias Vbias.n990 0.0972718
R16623 Vbias.n979 Vbias 0.0972718
R16624 Vbias Vbias.n978 0.0972718
R16625 Vbias.n969 Vbias 0.0972718
R16626 Vbias Vbias.n968 0.0972718
R16627 Vbias.n959 Vbias 0.0972718
R16628 Vbias Vbias.n958 0.0972718
R16629 Vbias.n949 Vbias 0.0972718
R16630 Vbias Vbias.n948 0.0972718
R16631 Vbias.n939 Vbias 0.0972718
R16632 Vbias Vbias.n938 0.0972718
R16633 Vbias.n929 Vbias 0.0972718
R16634 Vbias Vbias.n928 0.0972718
R16635 Vbias.n919 Vbias 0.0972718
R16636 Vbias Vbias.n918 0.0972718
R16637 Vbias.n914 Vbias 0.0972718
R16638 Vbias Vbias.n923 0.0972718
R16639 Vbias.n924 Vbias 0.0972718
R16640 Vbias Vbias.n933 0.0972718
R16641 Vbias.n934 Vbias 0.0972718
R16642 Vbias Vbias.n943 0.0972718
R16643 Vbias.n944 Vbias 0.0972718
R16644 Vbias Vbias.n953 0.0972718
R16645 Vbias.n954 Vbias 0.0972718
R16646 Vbias Vbias.n963 0.0972718
R16647 Vbias.n964 Vbias 0.0972718
R16648 Vbias Vbias.n973 0.0972718
R16649 Vbias.n974 Vbias 0.0972718
R16650 Vbias.n15 Vbias 0.0972718
R16651 Vbias.n985 Vbias 0.0972718
R16652 Vbias Vbias.n984 0.0972718
R16653 Vbias.n58 Vbias 0.0972718
R16654 Vbias.n61 Vbias 0.0972718
R16655 Vbias.n64 Vbias 0.0972718
R16656 Vbias.n67 Vbias 0.0972718
R16657 Vbias.n70 Vbias 0.0972718
R16658 Vbias.n73 Vbias 0.0972718
R16659 Vbias.n76 Vbias 0.0972718
R16660 Vbias.n79 Vbias 0.0972718
R16661 Vbias.n82 Vbias 0.0972718
R16662 Vbias.n85 Vbias 0.0972718
R16663 Vbias.n88 Vbias 0.0972718
R16664 Vbias.n91 Vbias 0.0972718
R16665 Vbias.n94 Vbias 0.0972718
R16666 Vbias.n908 Vbias 0.0972718
R16667 Vbias.n895 Vbias 0.0972718
R16668 Vbias.n894 Vbias 0.0972718
R16669 Vbias.n883 Vbias 0.0972718
R16670 Vbias.n882 Vbias 0.0972718
R16671 Vbias.n871 Vbias 0.0972718
R16672 Vbias.n870 Vbias 0.0972718
R16673 Vbias.n859 Vbias 0.0972718
R16674 Vbias.n858 Vbias 0.0972718
R16675 Vbias.n847 Vbias 0.0972718
R16676 Vbias.n846 Vbias 0.0972718
R16677 Vbias.n835 Vbias 0.0972718
R16678 Vbias.n834 Vbias 0.0972718
R16679 Vbias Vbias.n668 0.0972718
R16680 Vbias Vbias.n676 0.0972718
R16681 Vbias.n828 Vbias 0.0972718
R16682 Vbias.n829 Vbias 0.0972718
R16683 Vbias.n840 Vbias 0.0972718
R16684 Vbias.n841 Vbias 0.0972718
R16685 Vbias.n852 Vbias 0.0972718
R16686 Vbias.n853 Vbias 0.0972718
R16687 Vbias.n864 Vbias 0.0972718
R16688 Vbias.n865 Vbias 0.0972718
R16689 Vbias.n876 Vbias 0.0972718
R16690 Vbias.n877 Vbias 0.0972718
R16691 Vbias.n888 Vbias 0.0972718
R16692 Vbias.n889 Vbias 0.0972718
R16693 Vbias.n900 Vbias 0.0972718
R16694 Vbias.n903 Vbias 0.0972718
R16695 Vbias Vbias.n786 0.0972718
R16696 Vbias Vbias.n789 0.0972718
R16697 Vbias Vbias.n792 0.0972718
R16698 Vbias Vbias.n795 0.0972718
R16699 Vbias Vbias.n798 0.0972718
R16700 Vbias Vbias.n801 0.0972718
R16701 Vbias Vbias.n804 0.0972718
R16702 Vbias Vbias.n807 0.0972718
R16703 Vbias Vbias.n810 0.0972718
R16704 Vbias Vbias.n813 0.0972718
R16705 Vbias Vbias.n816 0.0972718
R16706 Vbias Vbias.n819 0.0972718
R16707 Vbias Vbias.n822 0.0972718
R16708 Vbias.n823 Vbias 0.0972718
R16709 Vbias.n697 Vbias 0.0972718
R16710 Vbias.n700 Vbias 0.0972718
R16711 Vbias.n701 Vbias 0.0972718
R16712 Vbias.n712 Vbias 0.0972718
R16713 Vbias.n713 Vbias 0.0972718
R16714 Vbias.n724 Vbias 0.0972718
R16715 Vbias.n725 Vbias 0.0972718
R16716 Vbias.n736 Vbias 0.0972718
R16717 Vbias.n737 Vbias 0.0972718
R16718 Vbias.n748 Vbias 0.0972718
R16719 Vbias.n749 Vbias 0.0972718
R16720 Vbias.n760 Vbias 0.0972718
R16721 Vbias.n761 Vbias 0.0972718
R16722 Vbias.n772 Vbias 0.0972718
R16723 Vbias.n773 Vbias 0.0972718
R16724 Vbias.n778 Vbias 0.0972718
R16725 Vbias.n767 Vbias 0.0972718
R16726 Vbias.n766 Vbias 0.0972718
R16727 Vbias.n755 Vbias 0.0972718
R16728 Vbias.n754 Vbias 0.0972718
R16729 Vbias.n743 Vbias 0.0972718
R16730 Vbias.n742 Vbias 0.0972718
R16731 Vbias.n731 Vbias 0.0972718
R16732 Vbias.n730 Vbias 0.0972718
R16733 Vbias.n719 Vbias 0.0972718
R16734 Vbias.n718 Vbias 0.0972718
R16735 Vbias.n707 Vbias 0.0972718
R16736 Vbias.n706 Vbias 0.0972718
R16737 Vbias.n685 Vbias 0.0972718
R16738 Vbias.n691 Vbias 0.0972718
R16739 Vbias Vbias.n690 0.0972718
R16740 Vbias Vbias.n230 0.0972718
R16741 Vbias Vbias.n227 0.0972718
R16742 Vbias Vbias.n224 0.0972718
R16743 Vbias Vbias.n221 0.0972718
R16744 Vbias Vbias.n218 0.0972718
R16745 Vbias Vbias.n215 0.0972718
R16746 Vbias Vbias.n212 0.0972718
R16747 Vbias Vbias.n209 0.0972718
R16748 Vbias Vbias.n206 0.0972718
R16749 Vbias Vbias.n203 0.0972718
R16750 Vbias Vbias.n200 0.0972718
R16751 Vbias Vbias.n197 0.0972718
R16752 Vbias Vbias.n194 0.0972718
R16753 Vbias Vbias.n584 0.0972718
R16754 Vbias.n585 Vbias 0.0972718
R16755 Vbias Vbias.n596 0.0972718
R16756 Vbias.n597 Vbias 0.0972718
R16757 Vbias Vbias.n608 0.0972718
R16758 Vbias.n609 Vbias 0.0972718
R16759 Vbias Vbias.n620 0.0972718
R16760 Vbias.n621 Vbias 0.0972718
R16761 Vbias Vbias.n632 0.0972718
R16762 Vbias.n633 Vbias 0.0972718
R16763 Vbias Vbias.n644 0.0972718
R16764 Vbias.n645 Vbias 0.0972718
R16765 Vbias Vbias.n656 0.0972718
R16766 Vbias Vbias.n659 0.0972718
R16767 Vbias.n529 Vbias 0.0972718
R16768 Vbias.n530 Vbias 0.0972718
R16769 Vbias.n651 Vbias 0.0972718
R16770 Vbias Vbias.n650 0.0972718
R16771 Vbias.n639 Vbias 0.0972718
R16772 Vbias Vbias.n638 0.0972718
R16773 Vbias.n627 Vbias 0.0972718
R16774 Vbias Vbias.n626 0.0972718
R16775 Vbias.n615 Vbias 0.0972718
R16776 Vbias Vbias.n614 0.0972718
R16777 Vbias.n603 Vbias 0.0972718
R16778 Vbias Vbias.n602 0.0972718
R16779 Vbias.n591 Vbias 0.0972718
R16780 Vbias Vbias.n590 0.0972718
R16781 Vbias.n579 Vbias 0.0972718
R16782 Vbias.n574 Vbias 0.0972718
R16783 Vbias.n571 Vbias 0.0972718
R16784 Vbias.n568 Vbias 0.0972718
R16785 Vbias.n565 Vbias 0.0972718
R16786 Vbias.n562 Vbias 0.0972718
R16787 Vbias.n559 Vbias 0.0972718
R16788 Vbias.n556 Vbias 0.0972718
R16789 Vbias.n553 Vbias 0.0972718
R16790 Vbias.n550 Vbias 0.0972718
R16791 Vbias.n547 Vbias 0.0972718
R16792 Vbias.n544 Vbias 0.0972718
R16793 Vbias.n541 Vbias 0.0972718
R16794 Vbias.n538 Vbias 0.0972718
R16795 Vbias.n535 Vbias 0.0972718
R16796 Vbias.n523 Vbias 0.0972718
R16797 Vbias Vbias.n522 0.0972718
R16798 Vbias Vbias.n519 0.0972718
R16799 Vbias.n508 Vbias 0.0972718
R16800 Vbias Vbias.n507 0.0972718
R16801 Vbias.n496 Vbias 0.0972718
R16802 Vbias Vbias.n495 0.0972718
R16803 Vbias.n484 Vbias 0.0972718
R16804 Vbias Vbias.n483 0.0972718
R16805 Vbias.n472 Vbias 0.0972718
R16806 Vbias Vbias.n471 0.0972718
R16807 Vbias.n460 Vbias 0.0972718
R16808 Vbias Vbias.n459 0.0972718
R16809 Vbias.n448 Vbias 0.0972718
R16810 Vbias Vbias.n447 0.0972718
R16811 Vbias.n442 Vbias 0.0972718
R16812 Vbias Vbias.n453 0.0972718
R16813 Vbias.n454 Vbias 0.0972718
R16814 Vbias Vbias.n465 0.0972718
R16815 Vbias.n466 Vbias 0.0972718
R16816 Vbias Vbias.n477 0.0972718
R16817 Vbias.n478 Vbias 0.0972718
R16818 Vbias Vbias.n489 0.0972718
R16819 Vbias.n490 Vbias 0.0972718
R16820 Vbias Vbias.n501 0.0972718
R16821 Vbias.n502 Vbias 0.0972718
R16822 Vbias Vbias.n513 0.0972718
R16823 Vbias.n514 Vbias 0.0972718
R16824 Vbias.n393 Vbias 0.0972718
R16825 Vbias Vbias.n384 0.0972718
R16826 Vbias Vbias.n377 0.0972718
R16827 Vbias Vbias.n376 0.0972718
R16828 Vbias Vbias.n373 0.0972718
R16829 Vbias Vbias.n370 0.0972718
R16830 Vbias Vbias.n367 0.0972718
R16831 Vbias Vbias.n364 0.0972718
R16832 Vbias Vbias.n361 0.0972718
R16833 Vbias Vbias.n358 0.0972718
R16834 Vbias Vbias.n355 0.0972718
R16835 Vbias Vbias.n352 0.0972718
R16836 Vbias Vbias.n349 0.0972718
R16837 Vbias Vbias.n346 0.0972718
R16838 Vbias Vbias.n343 0.0972718
R16839 Vbias Vbias.n340 0.0972718
R16840 Vbias.n437 Vbias 0.0972718
R16841 Vbias.n434 Vbias 0.0972718
R16842 Vbias.n431 Vbias 0.0972718
R16843 Vbias.n428 Vbias 0.0972718
R16844 Vbias.n425 Vbias 0.0972718
R16845 Vbias.n422 Vbias 0.0972718
R16846 Vbias.n419 Vbias 0.0972718
R16847 Vbias.n416 Vbias 0.0972718
R16848 Vbias.n413 Vbias 0.0972718
R16849 Vbias.n410 Vbias 0.0972718
R16850 Vbias.n407 Vbias 0.0972718
R16851 Vbias.n404 Vbias 0.0972718
R16852 Vbias.n401 Vbias 0.0972718
R16853 Vbias.n398 Vbias 0.0972718
R16854 Vbias.n380 Vbias 0.0972718
R16855 Vbias.n332 Vbias 0.0489375
R16856 Vbias.n378 Vbias 0.0489375
R16857 Vbias.n379 Vbias 0.0489375
R16858 Vbias.n329 Vbias 0.0489375
R16859 Vbias.n287 Vbias 0.0489375
R16860 Vbias.n279 Vbias 0.0489375
R16861 Vbias.n283 Vbias 0.0489375
R16862 Vbias.n275 Vbias 0.0489375
R16863 Vbias.n189 Vbias 0.0489375
R16864 Vbias.n144 Vbias 0.0489375
R16865 Vbias.n184 Vbias 0.0489375
R16866 Vbias.n140 Vbias 0.0489375
R16867 Vbias.n673 Vbias 0.0489375
R16868 Vbias.n97 Vbias 0.0489375
R16869 Vbias.n5 Vbias 0.0489375
R16870 Vbias.n52 Vbias 0.0489375
R16871 Vbias.n53 Vbias 0.0489375
R16872 Vbias.n49 Vbias 0.0489375
R16873 Vbias.n435 Vbias 0.0489375
R16874 Vbias.n338 Vbias 0.0489375
R16875 Vbias.n328 Vbias 0.0489375
R16876 Vbias.n326 Vbias 0.0489375
R16877 Vbias.n572 Vbias 0.0489375
R16878 Vbias.n273 Vbias 0.0489375
R16879 Vbias.n271 Vbias 0.0489375
R16880 Vbias.n192 Vbias 0.0489375
R16881 Vbias.n145 Vbias 0.0489375
R16882 Vbias.n147 Vbias 0.0489375
R16883 Vbias.n784 Vbias 0.0489375
R16884 Vbias.n100 Vbias 0.0489375
R16885 Vbias.n98 Vbias 0.0489375
R16886 Vbias.n92 Vbias 0.0489375
R16887 Vbias.n51 Vbias 0.0489375
R16888 Vbias.n48 Vbias 0.0489375
R16889 Vbias.n432 Vbias 0.0489375
R16890 Vbias.n341 Vbias 0.0489375
R16891 Vbias.n321 Vbias 0.0489375
R16892 Vbias.n323 Vbias 0.0489375
R16893 Vbias.n569 Vbias 0.0489375
R16894 Vbias.n268 Vbias 0.0489375
R16895 Vbias.n270 Vbias 0.0489375
R16896 Vbias.n195 Vbias 0.0489375
R16897 Vbias.n150 Vbias 0.0489375
R16898 Vbias.n148 Vbias 0.0489375
R16899 Vbias.n787 Vbias 0.0489375
R16900 Vbias.n101 Vbias 0.0489375
R16901 Vbias.n103 Vbias 0.0489375
R16902 Vbias.n89 Vbias 0.0489375
R16903 Vbias.n46 Vbias 0.0489375
R16904 Vbias.n43 Vbias 0.0489375
R16905 Vbias.n429 Vbias 0.0489375
R16906 Vbias.n344 Vbias 0.0489375
R16907 Vbias.n320 Vbias 0.0489375
R16908 Vbias.n318 Vbias 0.0489375
R16909 Vbias.n566 Vbias 0.0489375
R16910 Vbias.n267 Vbias 0.0489375
R16911 Vbias.n265 Vbias 0.0489375
R16912 Vbias.n198 Vbias 0.0489375
R16913 Vbias.n151 Vbias 0.0489375
R16914 Vbias.n153 Vbias 0.0489375
R16915 Vbias.n790 Vbias 0.0489375
R16916 Vbias.n106 Vbias 0.0489375
R16917 Vbias.n104 Vbias 0.0489375
R16918 Vbias.n86 Vbias 0.0489375
R16919 Vbias.n45 Vbias 0.0489375
R16920 Vbias.n42 Vbias 0.0489375
R16921 Vbias.n426 Vbias 0.0489375
R16922 Vbias.n347 Vbias 0.0489375
R16923 Vbias.n315 Vbias 0.0489375
R16924 Vbias.n317 Vbias 0.0489375
R16925 Vbias.n563 Vbias 0.0489375
R16926 Vbias.n262 Vbias 0.0489375
R16927 Vbias.n264 Vbias 0.0489375
R16928 Vbias.n201 Vbias 0.0489375
R16929 Vbias.n156 Vbias 0.0489375
R16930 Vbias.n154 Vbias 0.0489375
R16931 Vbias.n793 Vbias 0.0489375
R16932 Vbias.n107 Vbias 0.0489375
R16933 Vbias.n109 Vbias 0.0489375
R16934 Vbias.n83 Vbias 0.0489375
R16935 Vbias.n40 Vbias 0.0489375
R16936 Vbias.n37 Vbias 0.0489375
R16937 Vbias.n423 Vbias 0.0489375
R16938 Vbias.n350 Vbias 0.0489375
R16939 Vbias.n314 Vbias 0.0489375
R16940 Vbias.n312 Vbias 0.0489375
R16941 Vbias.n560 Vbias 0.0489375
R16942 Vbias.n261 Vbias 0.0489375
R16943 Vbias.n259 Vbias 0.0489375
R16944 Vbias.n204 Vbias 0.0489375
R16945 Vbias.n157 Vbias 0.0489375
R16946 Vbias.n159 Vbias 0.0489375
R16947 Vbias.n796 Vbias 0.0489375
R16948 Vbias.n112 Vbias 0.0489375
R16949 Vbias.n110 Vbias 0.0489375
R16950 Vbias.n80 Vbias 0.0489375
R16951 Vbias.n39 Vbias 0.0489375
R16952 Vbias.n36 Vbias 0.0489375
R16953 Vbias.n420 Vbias 0.0489375
R16954 Vbias.n353 Vbias 0.0489375
R16955 Vbias.n309 Vbias 0.0489375
R16956 Vbias.n311 Vbias 0.0489375
R16957 Vbias.n557 Vbias 0.0489375
R16958 Vbias.n256 Vbias 0.0489375
R16959 Vbias.n258 Vbias 0.0489375
R16960 Vbias.n207 Vbias 0.0489375
R16961 Vbias.n162 Vbias 0.0489375
R16962 Vbias.n160 Vbias 0.0489375
R16963 Vbias.n799 Vbias 0.0489375
R16964 Vbias.n113 Vbias 0.0489375
R16965 Vbias.n115 Vbias 0.0489375
R16966 Vbias.n77 Vbias 0.0489375
R16967 Vbias.n34 Vbias 0.0489375
R16968 Vbias.n31 Vbias 0.0489375
R16969 Vbias.n417 Vbias 0.0489375
R16970 Vbias.n356 Vbias 0.0489375
R16971 Vbias.n308 Vbias 0.0489375
R16972 Vbias.n306 Vbias 0.0489375
R16973 Vbias.n554 Vbias 0.0489375
R16974 Vbias.n255 Vbias 0.0489375
R16975 Vbias.n253 Vbias 0.0489375
R16976 Vbias.n210 Vbias 0.0489375
R16977 Vbias.n163 Vbias 0.0489375
R16978 Vbias.n165 Vbias 0.0489375
R16979 Vbias.n802 Vbias 0.0489375
R16980 Vbias.n118 Vbias 0.0489375
R16981 Vbias.n116 Vbias 0.0489375
R16982 Vbias.n74 Vbias 0.0489375
R16983 Vbias.n33 Vbias 0.0489375
R16984 Vbias.n30 Vbias 0.0489375
R16985 Vbias.n414 Vbias 0.0489375
R16986 Vbias.n359 Vbias 0.0489375
R16987 Vbias.n303 Vbias 0.0489375
R16988 Vbias.n305 Vbias 0.0489375
R16989 Vbias.n551 Vbias 0.0489375
R16990 Vbias.n250 Vbias 0.0489375
R16991 Vbias.n252 Vbias 0.0489375
R16992 Vbias.n213 Vbias 0.0489375
R16993 Vbias.n168 Vbias 0.0489375
R16994 Vbias.n166 Vbias 0.0489375
R16995 Vbias.n805 Vbias 0.0489375
R16996 Vbias.n119 Vbias 0.0489375
R16997 Vbias.n121 Vbias 0.0489375
R16998 Vbias.n71 Vbias 0.0489375
R16999 Vbias.n28 Vbias 0.0489375
R17000 Vbias.n25 Vbias 0.0489375
R17001 Vbias.n411 Vbias 0.0489375
R17002 Vbias.n362 Vbias 0.0489375
R17003 Vbias.n302 Vbias 0.0489375
R17004 Vbias.n300 Vbias 0.0489375
R17005 Vbias.n548 Vbias 0.0489375
R17006 Vbias.n249 Vbias 0.0489375
R17007 Vbias.n247 Vbias 0.0489375
R17008 Vbias.n216 Vbias 0.0489375
R17009 Vbias.n169 Vbias 0.0489375
R17010 Vbias.n171 Vbias 0.0489375
R17011 Vbias.n808 Vbias 0.0489375
R17012 Vbias.n124 Vbias 0.0489375
R17013 Vbias.n122 Vbias 0.0489375
R17014 Vbias.n68 Vbias 0.0489375
R17015 Vbias.n27 Vbias 0.0489375
R17016 Vbias.n24 Vbias 0.0489375
R17017 Vbias.n408 Vbias 0.0489375
R17018 Vbias.n365 Vbias 0.0489375
R17019 Vbias.n297 Vbias 0.0489375
R17020 Vbias.n299 Vbias 0.0489375
R17021 Vbias.n545 Vbias 0.0489375
R17022 Vbias.n244 Vbias 0.0489375
R17023 Vbias.n246 Vbias 0.0489375
R17024 Vbias.n219 Vbias 0.0489375
R17025 Vbias.n174 Vbias 0.0489375
R17026 Vbias.n172 Vbias 0.0489375
R17027 Vbias.n811 Vbias 0.0489375
R17028 Vbias.n125 Vbias 0.0489375
R17029 Vbias.n127 Vbias 0.0489375
R17030 Vbias.n65 Vbias 0.0489375
R17031 Vbias.n22 Vbias 0.0489375
R17032 Vbias.n19 Vbias 0.0489375
R17033 Vbias.n405 Vbias 0.0489375
R17034 Vbias.n368 Vbias 0.0489375
R17035 Vbias.n296 Vbias 0.0489375
R17036 Vbias.n294 Vbias 0.0489375
R17037 Vbias.n542 Vbias 0.0489375
R17038 Vbias.n243 Vbias 0.0489375
R17039 Vbias.n241 Vbias 0.0489375
R17040 Vbias.n222 Vbias 0.0489375
R17041 Vbias.n175 Vbias 0.0489375
R17042 Vbias.n177 Vbias 0.0489375
R17043 Vbias.n814 Vbias 0.0489375
R17044 Vbias.n130 Vbias 0.0489375
R17045 Vbias.n128 Vbias 0.0489375
R17046 Vbias.n62 Vbias 0.0489375
R17047 Vbias.n21 Vbias 0.0489375
R17048 Vbias.n18 Vbias 0.0489375
R17049 Vbias.n402 Vbias 0.0489375
R17050 Vbias.n371 Vbias 0.0489375
R17051 Vbias.n291 Vbias 0.0489375
R17052 Vbias.n293 Vbias 0.0489375
R17053 Vbias.n539 Vbias 0.0489375
R17054 Vbias.n238 Vbias 0.0489375
R17055 Vbias.n240 Vbias 0.0489375
R17056 Vbias.n225 Vbias 0.0489375
R17057 Vbias.n180 Vbias 0.0489375
R17058 Vbias.n178 Vbias 0.0489375
R17059 Vbias.n817 Vbias 0.0489375
R17060 Vbias.n131 Vbias 0.0489375
R17061 Vbias.n133 Vbias 0.0489375
R17062 Vbias.n59 Vbias 0.0489375
R17063 Vbias.n16 Vbias 0.0489375
R17064 Vbias.n11 Vbias 0.0489375
R17065 Vbias.n399 Vbias 0.0489375
R17066 Vbias.n374 Vbias 0.0489375
R17067 Vbias.n290 Vbias 0.0489375
R17068 Vbias.n288 Vbias 0.0489375
R17069 Vbias.n536 Vbias 0.0489375
R17070 Vbias.n237 Vbias 0.0489375
R17071 Vbias.n235 Vbias 0.0489375
R17072 Vbias.n228 Vbias 0.0489375
R17073 Vbias.n181 Vbias 0.0489375
R17074 Vbias.n183 Vbias 0.0489375
R17075 Vbias.n820 Vbias 0.0489375
R17076 Vbias.n136 Vbias 0.0489375
R17077 Vbias.n134 Vbias 0.0489375
R17078 Vbias.n56 Vbias 0.0489375
R17079 Vbias.n13 Vbias 0.0489375
R17080 Vbias.n10 Vbias 0.0489375
R17081 Vbias.n333 Vbias 0.0489375
R17082 Vbias.n334 Vbias 0.0489375
R17083 Vbias.n336 Vbias 0.0489375
R17084 Vbias.n520 Vbias 0.0489375
R17085 Vbias.n280 Vbias 0.0489375
R17086 Vbias.n282 Vbias 0.0489375
R17087 Vbias.n657 Vbias 0.0489375
R17088 Vbias.n231 Vbias 0.0489375
R17089 Vbias.n233 Vbias 0.0489375
R17090 Vbias.n698 Vbias 0.0489375
R17091 Vbias.n139 Vbias 0.0489375
R17092 Vbias.n137 Vbias 0.0489375
R17093 Vbias.n666 Vbias 0.0489375
R17094 Vbias.n6 Vbias 0.0489375
R17095 Vbias.n8 Vbias 0.0489375
R17096 Vbias.n1 Vbias 0.0489375
R17097 Vbias.n2 Vbias 0.0489375
R17098 Vbias.n55 Vbias 0.0489375
R17099 Vbias.n669 Vbias 0.0489375
R17100 Vbias.n901 Vbias 0.0489375
R17101 Vbias.n678 Vbias 0.0489375
R17102 Vbias.n141 Vbias 0.0489375
R17103 Vbias.n186 Vbias 0.0489375
R17104 Vbias.n190 Vbias 0.0489375
R17105 Vbias.n660 Vbias 0.0489375
R17106 Vbias.n274 Vbias 0.0489375
R17107 Vbias.n284 Vbias 0.0489375
R17108 Vbias.n324 Vbias 0.0489375
R17109 Vbias.n390 Vbias 0.0489375
R17110 Vbias.n330 Vbias 0.0489375
R17111 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R17112 XThR.Tn[12].n2 XThR.Tn[12].n1 243.679
R17113 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R17114 XThR.Tn[12].n2 XThR.Tn[12].n0 205.28
R17115 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R17116 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R17117 XThR.Tn[12] XThR.Tn[12].n78 161.363
R17118 XThR.Tn[12] XThR.Tn[12].n73 161.363
R17119 XThR.Tn[12] XThR.Tn[12].n68 161.363
R17120 XThR.Tn[12] XThR.Tn[12].n63 161.363
R17121 XThR.Tn[12] XThR.Tn[12].n58 161.363
R17122 XThR.Tn[12] XThR.Tn[12].n53 161.363
R17123 XThR.Tn[12] XThR.Tn[12].n48 161.363
R17124 XThR.Tn[12] XThR.Tn[12].n43 161.363
R17125 XThR.Tn[12] XThR.Tn[12].n38 161.363
R17126 XThR.Tn[12] XThR.Tn[12].n33 161.363
R17127 XThR.Tn[12] XThR.Tn[12].n28 161.363
R17128 XThR.Tn[12] XThR.Tn[12].n23 161.363
R17129 XThR.Tn[12] XThR.Tn[12].n18 161.363
R17130 XThR.Tn[12] XThR.Tn[12].n13 161.363
R17131 XThR.Tn[12] XThR.Tn[12].n8 161.363
R17132 XThR.Tn[12] XThR.Tn[12].n6 161.363
R17133 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R17134 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R17135 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R17136 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R17137 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R17138 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R17139 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R17140 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R17141 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R17142 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R17143 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R17144 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R17145 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R17146 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R17147 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R17148 XThR.Tn[12].n78 XThR.Tn[12].t18 161.106
R17149 XThR.Tn[12].n73 XThR.Tn[12].t24 161.106
R17150 XThR.Tn[12].n68 XThR.Tn[12].t67 161.106
R17151 XThR.Tn[12].n63 XThR.Tn[12].t52 161.106
R17152 XThR.Tn[12].n58 XThR.Tn[12].t16 161.106
R17153 XThR.Tn[12].n53 XThR.Tn[12].t40 161.106
R17154 XThR.Tn[12].n48 XThR.Tn[12].t22 161.106
R17155 XThR.Tn[12].n43 XThR.Tn[12].t65 161.106
R17156 XThR.Tn[12].n38 XThR.Tn[12].t51 161.106
R17157 XThR.Tn[12].n33 XThR.Tn[12].t56 161.106
R17158 XThR.Tn[12].n28 XThR.Tn[12].t39 161.106
R17159 XThR.Tn[12].n23 XThR.Tn[12].t66 161.106
R17160 XThR.Tn[12].n18 XThR.Tn[12].t38 161.106
R17161 XThR.Tn[12].n13 XThR.Tn[12].t20 161.106
R17162 XThR.Tn[12].n8 XThR.Tn[12].t43 161.106
R17163 XThR.Tn[12].n6 XThR.Tn[12].t28 161.106
R17164 XThR.Tn[12].n79 XThR.Tn[12].t58 159.978
R17165 XThR.Tn[12].n74 XThR.Tn[12].t62 159.978
R17166 XThR.Tn[12].n69 XThR.Tn[12].t47 159.978
R17167 XThR.Tn[12].n64 XThR.Tn[12].t31 159.978
R17168 XThR.Tn[12].n59 XThR.Tn[12].t55 159.978
R17169 XThR.Tn[12].n54 XThR.Tn[12].t19 159.978
R17170 XThR.Tn[12].n49 XThR.Tn[12].t61 159.978
R17171 XThR.Tn[12].n44 XThR.Tn[12].t44 159.978
R17172 XThR.Tn[12].n39 XThR.Tn[12].t29 159.978
R17173 XThR.Tn[12].n34 XThR.Tn[12].t37 159.978
R17174 XThR.Tn[12].n29 XThR.Tn[12].t17 159.978
R17175 XThR.Tn[12].n24 XThR.Tn[12].t46 159.978
R17176 XThR.Tn[12].n19 XThR.Tn[12].t15 159.978
R17177 XThR.Tn[12].n14 XThR.Tn[12].t60 159.978
R17178 XThR.Tn[12].n9 XThR.Tn[12].t21 159.978
R17179 XThR.Tn[12].n78 XThR.Tn[12].t69 145.038
R17180 XThR.Tn[12].n73 XThR.Tn[12].t32 145.038
R17181 XThR.Tn[12].n68 XThR.Tn[12].t73 145.038
R17182 XThR.Tn[12].n63 XThR.Tn[12].t57 145.038
R17183 XThR.Tn[12].n58 XThR.Tn[12].t25 145.038
R17184 XThR.Tn[12].n53 XThR.Tn[12].t68 145.038
R17185 XThR.Tn[12].n48 XThR.Tn[12].t12 145.038
R17186 XThR.Tn[12].n43 XThR.Tn[12].t59 145.038
R17187 XThR.Tn[12].n38 XThR.Tn[12].t54 145.038
R17188 XThR.Tn[12].n33 XThR.Tn[12].t23 145.038
R17189 XThR.Tn[12].n28 XThR.Tn[12].t48 145.038
R17190 XThR.Tn[12].n23 XThR.Tn[12].t70 145.038
R17191 XThR.Tn[12].n18 XThR.Tn[12].t45 145.038
R17192 XThR.Tn[12].n13 XThR.Tn[12].t30 145.038
R17193 XThR.Tn[12].n8 XThR.Tn[12].t53 145.038
R17194 XThR.Tn[12].n6 XThR.Tn[12].t36 145.038
R17195 XThR.Tn[12].n79 XThR.Tn[12].t27 143.911
R17196 XThR.Tn[12].n74 XThR.Tn[12].t50 143.911
R17197 XThR.Tn[12].n69 XThR.Tn[12].t34 143.911
R17198 XThR.Tn[12].n64 XThR.Tn[12].t13 143.911
R17199 XThR.Tn[12].n59 XThR.Tn[12].t42 143.911
R17200 XThR.Tn[12].n54 XThR.Tn[12].t26 143.911
R17201 XThR.Tn[12].n49 XThR.Tn[12].t35 143.911
R17202 XThR.Tn[12].n44 XThR.Tn[12].t14 143.911
R17203 XThR.Tn[12].n39 XThR.Tn[12].t72 143.911
R17204 XThR.Tn[12].n34 XThR.Tn[12].t41 143.911
R17205 XThR.Tn[12].n29 XThR.Tn[12].t64 143.911
R17206 XThR.Tn[12].n24 XThR.Tn[12].t33 143.911
R17207 XThR.Tn[12].n19 XThR.Tn[12].t63 143.911
R17208 XThR.Tn[12].n14 XThR.Tn[12].t49 143.911
R17209 XThR.Tn[12].n9 XThR.Tn[12].t71 143.911
R17210 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17211 XThR.Tn[12].n85 XThR.Tn[12].t6 26.5955
R17212 XThR.Tn[12].n85 XThR.Tn[12].t4 26.5955
R17213 XThR.Tn[12].n86 XThR.Tn[12].t7 26.5955
R17214 XThR.Tn[12].n86 XThR.Tn[12].t5 26.5955
R17215 XThR.Tn[12].n0 XThR.Tn[12].t0 26.5955
R17216 XThR.Tn[12].n0 XThR.Tn[12].t2 26.5955
R17217 XThR.Tn[12].n1 XThR.Tn[12].t3 26.5955
R17218 XThR.Tn[12].n1 XThR.Tn[12].t1 26.5955
R17219 XThR.Tn[12].n4 XThR.Tn[12].t10 24.9236
R17220 XThR.Tn[12].n4 XThR.Tn[12].t8 24.9236
R17221 XThR.Tn[12].n3 XThR.Tn[12].t11 24.9236
R17222 XThR.Tn[12].n3 XThR.Tn[12].t9 24.9236
R17223 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R17224 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R17225 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R17226 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R17227 XThR.Tn[12] XThR.Tn[12].n7 5.34038
R17228 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R17229 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R17230 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R17231 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R17232 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R17233 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R17234 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R17235 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R17236 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R17237 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R17238 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R17239 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R17240 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R17241 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R17242 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R17243 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R17244 XThR.Tn[12].n12 XThR.Tn[12] 2.52282
R17245 XThR.Tn[12].n17 XThR.Tn[12] 2.52282
R17246 XThR.Tn[12].n22 XThR.Tn[12] 2.52282
R17247 XThR.Tn[12].n27 XThR.Tn[12] 2.52282
R17248 XThR.Tn[12].n32 XThR.Tn[12] 2.52282
R17249 XThR.Tn[12].n37 XThR.Tn[12] 2.52282
R17250 XThR.Tn[12].n42 XThR.Tn[12] 2.52282
R17251 XThR.Tn[12].n47 XThR.Tn[12] 2.52282
R17252 XThR.Tn[12].n52 XThR.Tn[12] 2.52282
R17253 XThR.Tn[12].n57 XThR.Tn[12] 2.52282
R17254 XThR.Tn[12].n62 XThR.Tn[12] 2.52282
R17255 XThR.Tn[12].n67 XThR.Tn[12] 2.52282
R17256 XThR.Tn[12].n72 XThR.Tn[12] 2.52282
R17257 XThR.Tn[12].n77 XThR.Tn[12] 2.52282
R17258 XThR.Tn[12].n82 XThR.Tn[12] 2.52282
R17259 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R17260 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R17261 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R17262 XThR.Tn[12].n80 XThR.Tn[12] 1.08677
R17263 XThR.Tn[12].n75 XThR.Tn[12] 1.08677
R17264 XThR.Tn[12].n70 XThR.Tn[12] 1.08677
R17265 XThR.Tn[12].n65 XThR.Tn[12] 1.08677
R17266 XThR.Tn[12].n60 XThR.Tn[12] 1.08677
R17267 XThR.Tn[12].n55 XThR.Tn[12] 1.08677
R17268 XThR.Tn[12].n50 XThR.Tn[12] 1.08677
R17269 XThR.Tn[12].n45 XThR.Tn[12] 1.08677
R17270 XThR.Tn[12].n40 XThR.Tn[12] 1.08677
R17271 XThR.Tn[12].n35 XThR.Tn[12] 1.08677
R17272 XThR.Tn[12].n30 XThR.Tn[12] 1.08677
R17273 XThR.Tn[12].n25 XThR.Tn[12] 1.08677
R17274 XThR.Tn[12].n20 XThR.Tn[12] 1.08677
R17275 XThR.Tn[12].n15 XThR.Tn[12] 1.08677
R17276 XThR.Tn[12].n10 XThR.Tn[12] 1.08677
R17277 XThR.Tn[12] XThR.Tn[12].n12 0.839786
R17278 XThR.Tn[12] XThR.Tn[12].n17 0.839786
R17279 XThR.Tn[12] XThR.Tn[12].n22 0.839786
R17280 XThR.Tn[12] XThR.Tn[12].n27 0.839786
R17281 XThR.Tn[12] XThR.Tn[12].n32 0.839786
R17282 XThR.Tn[12] XThR.Tn[12].n37 0.839786
R17283 XThR.Tn[12] XThR.Tn[12].n42 0.839786
R17284 XThR.Tn[12] XThR.Tn[12].n47 0.839786
R17285 XThR.Tn[12] XThR.Tn[12].n52 0.839786
R17286 XThR.Tn[12] XThR.Tn[12].n57 0.839786
R17287 XThR.Tn[12] XThR.Tn[12].n62 0.839786
R17288 XThR.Tn[12] XThR.Tn[12].n67 0.839786
R17289 XThR.Tn[12] XThR.Tn[12].n72 0.839786
R17290 XThR.Tn[12] XThR.Tn[12].n77 0.839786
R17291 XThR.Tn[12] XThR.Tn[12].n82 0.839786
R17292 XThR.Tn[12].n7 XThR.Tn[12] 0.499542
R17293 XThR.Tn[12].n81 XThR.Tn[12] 0.063
R17294 XThR.Tn[12].n76 XThR.Tn[12] 0.063
R17295 XThR.Tn[12].n71 XThR.Tn[12] 0.063
R17296 XThR.Tn[12].n66 XThR.Tn[12] 0.063
R17297 XThR.Tn[12].n61 XThR.Tn[12] 0.063
R17298 XThR.Tn[12].n56 XThR.Tn[12] 0.063
R17299 XThR.Tn[12].n51 XThR.Tn[12] 0.063
R17300 XThR.Tn[12].n46 XThR.Tn[12] 0.063
R17301 XThR.Tn[12].n41 XThR.Tn[12] 0.063
R17302 XThR.Tn[12].n36 XThR.Tn[12] 0.063
R17303 XThR.Tn[12].n31 XThR.Tn[12] 0.063
R17304 XThR.Tn[12].n26 XThR.Tn[12] 0.063
R17305 XThR.Tn[12].n21 XThR.Tn[12] 0.063
R17306 XThR.Tn[12].n16 XThR.Tn[12] 0.063
R17307 XThR.Tn[12].n11 XThR.Tn[12] 0.063
R17308 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R17309 XThR.Tn[12] XThR.Tn[12].n83 0.038
R17310 XThR.Tn[12].n7 XThR.Tn[12] 0.0143889
R17311 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00771154
R17312 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00771154
R17313 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00771154
R17314 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00771154
R17315 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00771154
R17316 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00771154
R17317 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00771154
R17318 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00771154
R17319 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00771154
R17320 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00771154
R17321 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00771154
R17322 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00771154
R17323 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00771154
R17324 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00771154
R17325 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00771154
R17326 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R17327 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R17328 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R17329 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R17330 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R17331 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R17332 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R17333 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R17334 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R17335 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R17336 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R17337 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R17338 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R17339 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R17340 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R17341 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R17342 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R17343 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R17344 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R17345 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R17346 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R17347 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R17348 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R17349 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R17350 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R17351 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R17352 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R17353 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R17354 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R17355 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R17356 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R17357 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R17358 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R17359 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R17360 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R17361 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R17362 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R17363 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R17364 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R17365 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R17366 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R17367 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R17368 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R17369 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R17370 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R17371 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R17372 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R17373 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R17374 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R17375 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R17376 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R17377 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R17378 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R17379 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R17380 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R17381 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R17382 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R17383 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R17384 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R17385 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R17386 XThC.XTBN.Y.n192 XThC.XTBN.Y.n191 208.964
R17387 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R17388 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R17389 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R17390 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R17391 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R17392 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R17393 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R17394 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R17395 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R17396 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R17397 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R17398 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R17399 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R17400 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R17401 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R17402 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R17403 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R17404 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R17405 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R17406 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R17407 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R17408 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R17409 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R17410 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R17411 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R17412 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R17413 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R17414 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R17415 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R17416 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R17417 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R17418 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R17419 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R17420 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R17421 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R17422 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R17423 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R17424 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R17425 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R17426 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R17427 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R17428 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R17429 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R17430 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R17431 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R17432 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R17433 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R17434 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R17435 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R17436 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R17437 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R17438 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R17439 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R17440 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R17441 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R17442 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R17443 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R17444 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R17445 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R17446 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R17447 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R17448 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R17449 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R17450 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R17451 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R17452 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R17453 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R17454 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R17455 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R17456 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R17457 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R17458 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R17459 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R17460 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R17461 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R17462 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R17463 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R17464 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R17465 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R17466 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R17467 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R17468 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R17469 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R17470 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R17471 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R17472 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R17473 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R17474 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R17475 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R17476 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R17477 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R17478 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R17479 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R17480 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R17481 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R17482 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R17483 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R17484 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R17485 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R17486 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R17487 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R17488 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R17489 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R17490 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R17491 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R17492 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R17493 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R17494 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R17495 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R17496 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R17497 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R17498 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R17499 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R17500 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R17501 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R17502 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R17503 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R17504 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R17505 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R17506 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R17507 XThC.XTBN.Y XThC.XTBN.Y.n188 96.8352
R17508 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R17509 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R17510 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R17511 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R17512 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R17513 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R17514 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R17515 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R17516 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R17517 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R17518 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R17519 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R17520 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R17521 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R17522 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R17523 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R17524 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R17525 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R17526 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R17527 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R17528 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R17529 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R17530 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R17531 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R17532 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R17533 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R17534 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R17535 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R17536 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R17537 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R17538 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R17539 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R17540 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R17541 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R17542 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R17543 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R17544 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R17545 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R17546 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R17547 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R17548 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R17549 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R17550 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R17551 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R17552 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R17553 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R17554 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R17555 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R17556 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R17557 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R17558 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R17559 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R17560 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R17561 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R17562 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R17563 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R17564 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R17565 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R17566 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R17567 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R17568 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R17569 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R17570 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R17571 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R17572 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R17573 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R17574 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R17575 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R17576 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R17577 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R17578 XThC.XTBN.Y.n191 XThC.XTBN.Y.t0 26.5955
R17579 XThC.XTBN.Y.n191 XThC.XTBN.Y.t1 26.5955
R17580 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 24.9236
R17581 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 24.9236
R17582 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R17583 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R17584 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R17585 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R17586 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R17587 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R17588 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R17589 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R17590 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R17591 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R17592 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R17593 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R17594 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R17595 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R17596 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R17597 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R17598 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R17599 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R17600 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R17601 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R17602 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R17603 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R17604 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R17605 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R17606 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R17607 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R17608 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R17609 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R17610 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R17611 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R17612 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R17613 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R17614 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R17615 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R17616 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R17617 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R17618 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R17619 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R17620 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R17621 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R17622 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R17623 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R17624 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R17625 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R17626 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R17627 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R17628 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R17629 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R17630 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R17631 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R17632 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R17633 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R17634 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R17635 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R17636 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R17637 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R17638 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R17639 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R17640 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R17641 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R17642 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R17643 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R17644 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R17645 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R17646 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R17647 XThC.XTBN.Y XThC.XTBN.Y.n190 12.5445
R17648 XThC.XTBN.Y XThC.XTBN.Y.n189 11.2645
R17649 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R17650 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R17651 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R17652 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R17653 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R17654 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R17655 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R17656 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R17657 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R17658 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R17659 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R17660 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R17661 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R17662 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R17663 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R17664 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R17665 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R17666 XThC.XTBN.Y.n189 XThC.XTBN.Y 6.1445
R17667 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R17668 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R17669 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R17670 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R17671 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R17672 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R17673 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R17674 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R17675 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R17676 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R17677 XThC.XTBN.Y.n190 XThC.XTBN.Y 4.8645
R17678 XThC.XTBN.Y.n189 XThC.XTBN.Y 4.65505
R17679 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R17680 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R17681 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R17682 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R17683 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R17684 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R17685 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R17686 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R17687 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R17688 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R17689 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R17690 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R17691 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R17692 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R17693 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R17694 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R17695 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R17696 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R17697 XThC.XTBN.Y.n192 XThC.XTBN.Y 2.0485
R17698 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R17699 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R17700 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R17701 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R17702 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R17703 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R17704 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R17705 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R17706 XThC.XTBN.Y XThC.XTBN.Y.n192 1.55202
R17707 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R17708 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R17709 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R17710 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R17711 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R17712 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R17713 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R17714 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R17715 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R17716 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R17717 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R17718 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R17719 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R17720 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R17721 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R17722 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R17723 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R17724 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R17725 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R17726 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R17727 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R17728 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R17729 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R17730 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R17731 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R17732 XThC.Tn[6].n73 XThC.Tn[6].n71 332.332
R17733 XThC.Tn[6].n73 XThC.Tn[6].n72 296.493
R17734 XThC.Tn[6].n68 XThC.Tn[6].n66 161.365
R17735 XThC.Tn[6].n64 XThC.Tn[6].n62 161.365
R17736 XThC.Tn[6].n60 XThC.Tn[6].n58 161.365
R17737 XThC.Tn[6].n56 XThC.Tn[6].n54 161.365
R17738 XThC.Tn[6].n52 XThC.Tn[6].n50 161.365
R17739 XThC.Tn[6].n48 XThC.Tn[6].n46 161.365
R17740 XThC.Tn[6].n44 XThC.Tn[6].n42 161.365
R17741 XThC.Tn[6].n40 XThC.Tn[6].n38 161.365
R17742 XThC.Tn[6].n36 XThC.Tn[6].n34 161.365
R17743 XThC.Tn[6].n32 XThC.Tn[6].n30 161.365
R17744 XThC.Tn[6].n28 XThC.Tn[6].n26 161.365
R17745 XThC.Tn[6].n24 XThC.Tn[6].n22 161.365
R17746 XThC.Tn[6].n20 XThC.Tn[6].n18 161.365
R17747 XThC.Tn[6].n16 XThC.Tn[6].n14 161.365
R17748 XThC.Tn[6].n12 XThC.Tn[6].n10 161.365
R17749 XThC.Tn[6].n9 XThC.Tn[6].n7 161.365
R17750 XThC.Tn[6].n66 XThC.Tn[6].t34 161.202
R17751 XThC.Tn[6].n62 XThC.Tn[6].t24 161.202
R17752 XThC.Tn[6].n58 XThC.Tn[6].t43 161.202
R17753 XThC.Tn[6].n54 XThC.Tn[6].t41 161.202
R17754 XThC.Tn[6].n50 XThC.Tn[6].t32 161.202
R17755 XThC.Tn[6].n46 XThC.Tn[6].t21 161.202
R17756 XThC.Tn[6].n42 XThC.Tn[6].t19 161.202
R17757 XThC.Tn[6].n38 XThC.Tn[6].t31 161.202
R17758 XThC.Tn[6].n34 XThC.Tn[6].t29 161.202
R17759 XThC.Tn[6].n30 XThC.Tn[6].t22 161.202
R17760 XThC.Tn[6].n26 XThC.Tn[6].t38 161.202
R17761 XThC.Tn[6].n22 XThC.Tn[6].t37 161.202
R17762 XThC.Tn[6].n18 XThC.Tn[6].t18 161.202
R17763 XThC.Tn[6].n14 XThC.Tn[6].t17 161.202
R17764 XThC.Tn[6].n10 XThC.Tn[6].t13 161.202
R17765 XThC.Tn[6].n7 XThC.Tn[6].t26 161.202
R17766 XThC.Tn[6].n66 XThC.Tn[6].t30 145.137
R17767 XThC.Tn[6].n62 XThC.Tn[6].t20 145.137
R17768 XThC.Tn[6].n58 XThC.Tn[6].t39 145.137
R17769 XThC.Tn[6].n54 XThC.Tn[6].t36 145.137
R17770 XThC.Tn[6].n50 XThC.Tn[6].t28 145.137
R17771 XThC.Tn[6].n46 XThC.Tn[6].t15 145.137
R17772 XThC.Tn[6].n42 XThC.Tn[6].t14 145.137
R17773 XThC.Tn[6].n38 XThC.Tn[6].t27 145.137
R17774 XThC.Tn[6].n34 XThC.Tn[6].t25 145.137
R17775 XThC.Tn[6].n30 XThC.Tn[6].t16 145.137
R17776 XThC.Tn[6].n26 XThC.Tn[6].t35 145.137
R17777 XThC.Tn[6].n22 XThC.Tn[6].t33 145.137
R17778 XThC.Tn[6].n18 XThC.Tn[6].t12 145.137
R17779 XThC.Tn[6].n14 XThC.Tn[6].t42 145.137
R17780 XThC.Tn[6].n10 XThC.Tn[6].t40 145.137
R17781 XThC.Tn[6].n7 XThC.Tn[6].t23 145.137
R17782 XThC.Tn[6].n2 XThC.Tn[6].n0 135.248
R17783 XThC.Tn[6].n2 XThC.Tn[6].n1 98.982
R17784 XThC.Tn[6].n4 XThC.Tn[6].n3 98.982
R17785 XThC.Tn[6].n6 XThC.Tn[6].n5 98.982
R17786 XThC.Tn[6].n4 XThC.Tn[6].n2 36.2672
R17787 XThC.Tn[6].n6 XThC.Tn[6].n4 36.2672
R17788 XThC.Tn[6].n70 XThC.Tn[6].n6 32.6405
R17789 XThC.Tn[6].n71 XThC.Tn[6].t1 26.5955
R17790 XThC.Tn[6].n71 XThC.Tn[6].t0 26.5955
R17791 XThC.Tn[6].n72 XThC.Tn[6].t3 26.5955
R17792 XThC.Tn[6].n72 XThC.Tn[6].t2 26.5955
R17793 XThC.Tn[6].n0 XThC.Tn[6].t11 24.9236
R17794 XThC.Tn[6].n0 XThC.Tn[6].t10 24.9236
R17795 XThC.Tn[6].n1 XThC.Tn[6].t9 24.9236
R17796 XThC.Tn[6].n1 XThC.Tn[6].t8 24.9236
R17797 XThC.Tn[6].n3 XThC.Tn[6].t6 24.9236
R17798 XThC.Tn[6].n3 XThC.Tn[6].t5 24.9236
R17799 XThC.Tn[6].n5 XThC.Tn[6].t4 24.9236
R17800 XThC.Tn[6].n5 XThC.Tn[6].t7 24.9236
R17801 XThC.Tn[6].n74 XThC.Tn[6].n73 18.5605
R17802 XThC.Tn[6].n74 XThC.Tn[6].n70 11.5205
R17803 XThC.Tn[6] XThC.Tn[6].n9 8.0245
R17804 XThC.Tn[6].n69 XThC.Tn[6].n68 7.9105
R17805 XThC.Tn[6].n65 XThC.Tn[6].n64 7.9105
R17806 XThC.Tn[6].n61 XThC.Tn[6].n60 7.9105
R17807 XThC.Tn[6].n57 XThC.Tn[6].n56 7.9105
R17808 XThC.Tn[6].n53 XThC.Tn[6].n52 7.9105
R17809 XThC.Tn[6].n49 XThC.Tn[6].n48 7.9105
R17810 XThC.Tn[6].n45 XThC.Tn[6].n44 7.9105
R17811 XThC.Tn[6].n41 XThC.Tn[6].n40 7.9105
R17812 XThC.Tn[6].n37 XThC.Tn[6].n36 7.9105
R17813 XThC.Tn[6].n33 XThC.Tn[6].n32 7.9105
R17814 XThC.Tn[6].n29 XThC.Tn[6].n28 7.9105
R17815 XThC.Tn[6].n25 XThC.Tn[6].n24 7.9105
R17816 XThC.Tn[6].n21 XThC.Tn[6].n20 7.9105
R17817 XThC.Tn[6].n17 XThC.Tn[6].n16 7.9105
R17818 XThC.Tn[6].n13 XThC.Tn[6].n12 7.9105
R17819 XThC.Tn[6].n70 XThC.Tn[6] 5.42203
R17820 XThC.Tn[6] XThC.Tn[6].n74 0.6405
R17821 XThC.Tn[6].n13 XThC.Tn[6] 0.235138
R17822 XThC.Tn[6].n17 XThC.Tn[6] 0.235138
R17823 XThC.Tn[6].n21 XThC.Tn[6] 0.235138
R17824 XThC.Tn[6].n25 XThC.Tn[6] 0.235138
R17825 XThC.Tn[6].n29 XThC.Tn[6] 0.235138
R17826 XThC.Tn[6].n33 XThC.Tn[6] 0.235138
R17827 XThC.Tn[6].n37 XThC.Tn[6] 0.235138
R17828 XThC.Tn[6].n41 XThC.Tn[6] 0.235138
R17829 XThC.Tn[6].n45 XThC.Tn[6] 0.235138
R17830 XThC.Tn[6].n49 XThC.Tn[6] 0.235138
R17831 XThC.Tn[6].n53 XThC.Tn[6] 0.235138
R17832 XThC.Tn[6].n57 XThC.Tn[6] 0.235138
R17833 XThC.Tn[6].n61 XThC.Tn[6] 0.235138
R17834 XThC.Tn[6].n65 XThC.Tn[6] 0.235138
R17835 XThC.Tn[6].n69 XThC.Tn[6] 0.235138
R17836 XThC.Tn[6] XThC.Tn[6].n13 0.114505
R17837 XThC.Tn[6] XThC.Tn[6].n17 0.114505
R17838 XThC.Tn[6] XThC.Tn[6].n21 0.114505
R17839 XThC.Tn[6] XThC.Tn[6].n25 0.114505
R17840 XThC.Tn[6] XThC.Tn[6].n29 0.114505
R17841 XThC.Tn[6] XThC.Tn[6].n33 0.114505
R17842 XThC.Tn[6] XThC.Tn[6].n37 0.114505
R17843 XThC.Tn[6] XThC.Tn[6].n41 0.114505
R17844 XThC.Tn[6] XThC.Tn[6].n45 0.114505
R17845 XThC.Tn[6] XThC.Tn[6].n49 0.114505
R17846 XThC.Tn[6] XThC.Tn[6].n53 0.114505
R17847 XThC.Tn[6] XThC.Tn[6].n57 0.114505
R17848 XThC.Tn[6] XThC.Tn[6].n61 0.114505
R17849 XThC.Tn[6] XThC.Tn[6].n65 0.114505
R17850 XThC.Tn[6] XThC.Tn[6].n69 0.114505
R17851 XThC.Tn[6].n68 XThC.Tn[6].n67 0.0599512
R17852 XThC.Tn[6].n64 XThC.Tn[6].n63 0.0599512
R17853 XThC.Tn[6].n60 XThC.Tn[6].n59 0.0599512
R17854 XThC.Tn[6].n56 XThC.Tn[6].n55 0.0599512
R17855 XThC.Tn[6].n52 XThC.Tn[6].n51 0.0599512
R17856 XThC.Tn[6].n48 XThC.Tn[6].n47 0.0599512
R17857 XThC.Tn[6].n44 XThC.Tn[6].n43 0.0599512
R17858 XThC.Tn[6].n40 XThC.Tn[6].n39 0.0599512
R17859 XThC.Tn[6].n36 XThC.Tn[6].n35 0.0599512
R17860 XThC.Tn[6].n32 XThC.Tn[6].n31 0.0599512
R17861 XThC.Tn[6].n28 XThC.Tn[6].n27 0.0599512
R17862 XThC.Tn[6].n24 XThC.Tn[6].n23 0.0599512
R17863 XThC.Tn[6].n20 XThC.Tn[6].n19 0.0599512
R17864 XThC.Tn[6].n16 XThC.Tn[6].n15 0.0599512
R17865 XThC.Tn[6].n12 XThC.Tn[6].n11 0.0599512
R17866 XThC.Tn[6].n9 XThC.Tn[6].n8 0.0599512
R17867 XThC.Tn[6].n67 XThC.Tn[6] 0.0469286
R17868 XThC.Tn[6].n63 XThC.Tn[6] 0.0469286
R17869 XThC.Tn[6].n59 XThC.Tn[6] 0.0469286
R17870 XThC.Tn[6].n55 XThC.Tn[6] 0.0469286
R17871 XThC.Tn[6].n51 XThC.Tn[6] 0.0469286
R17872 XThC.Tn[6].n47 XThC.Tn[6] 0.0469286
R17873 XThC.Tn[6].n43 XThC.Tn[6] 0.0469286
R17874 XThC.Tn[6].n39 XThC.Tn[6] 0.0469286
R17875 XThC.Tn[6].n35 XThC.Tn[6] 0.0469286
R17876 XThC.Tn[6].n31 XThC.Tn[6] 0.0469286
R17877 XThC.Tn[6].n27 XThC.Tn[6] 0.0469286
R17878 XThC.Tn[6].n23 XThC.Tn[6] 0.0469286
R17879 XThC.Tn[6].n19 XThC.Tn[6] 0.0469286
R17880 XThC.Tn[6].n15 XThC.Tn[6] 0.0469286
R17881 XThC.Tn[6].n11 XThC.Tn[6] 0.0469286
R17882 XThC.Tn[6].n8 XThC.Tn[6] 0.0469286
R17883 XThC.Tn[6].n67 XThC.Tn[6] 0.0401341
R17884 XThC.Tn[6].n63 XThC.Tn[6] 0.0401341
R17885 XThC.Tn[6].n59 XThC.Tn[6] 0.0401341
R17886 XThC.Tn[6].n55 XThC.Tn[6] 0.0401341
R17887 XThC.Tn[6].n51 XThC.Tn[6] 0.0401341
R17888 XThC.Tn[6].n47 XThC.Tn[6] 0.0401341
R17889 XThC.Tn[6].n43 XThC.Tn[6] 0.0401341
R17890 XThC.Tn[6].n39 XThC.Tn[6] 0.0401341
R17891 XThC.Tn[6].n35 XThC.Tn[6] 0.0401341
R17892 XThC.Tn[6].n31 XThC.Tn[6] 0.0401341
R17893 XThC.Tn[6].n27 XThC.Tn[6] 0.0401341
R17894 XThC.Tn[6].n23 XThC.Tn[6] 0.0401341
R17895 XThC.Tn[6].n19 XThC.Tn[6] 0.0401341
R17896 XThC.Tn[6].n15 XThC.Tn[6] 0.0401341
R17897 XThC.Tn[6].n11 XThC.Tn[6] 0.0401341
R17898 XThC.Tn[6].n8 XThC.Tn[6] 0.0401341
R17899 XThR.Tn[9].n87 XThR.Tn[9].n86 256.104
R17900 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R17901 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R17902 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R17903 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R17904 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R17905 XThR.Tn[9] XThR.Tn[9].n78 161.363
R17906 XThR.Tn[9] XThR.Tn[9].n73 161.363
R17907 XThR.Tn[9] XThR.Tn[9].n68 161.363
R17908 XThR.Tn[9] XThR.Tn[9].n63 161.363
R17909 XThR.Tn[9] XThR.Tn[9].n58 161.363
R17910 XThR.Tn[9] XThR.Tn[9].n53 161.363
R17911 XThR.Tn[9] XThR.Tn[9].n48 161.363
R17912 XThR.Tn[9] XThR.Tn[9].n43 161.363
R17913 XThR.Tn[9] XThR.Tn[9].n38 161.363
R17914 XThR.Tn[9] XThR.Tn[9].n33 161.363
R17915 XThR.Tn[9] XThR.Tn[9].n28 161.363
R17916 XThR.Tn[9] XThR.Tn[9].n23 161.363
R17917 XThR.Tn[9] XThR.Tn[9].n18 161.363
R17918 XThR.Tn[9] XThR.Tn[9].n13 161.363
R17919 XThR.Tn[9] XThR.Tn[9].n8 161.363
R17920 XThR.Tn[9] XThR.Tn[9].n6 161.363
R17921 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R17922 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R17923 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R17924 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R17925 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R17926 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R17927 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R17928 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R17929 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R17930 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R17931 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R17932 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R17933 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R17934 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R17935 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R17936 XThR.Tn[9].n78 XThR.Tn[9].t63 161.106
R17937 XThR.Tn[9].n73 XThR.Tn[9].t69 161.106
R17938 XThR.Tn[9].n68 XThR.Tn[9].t47 161.106
R17939 XThR.Tn[9].n63 XThR.Tn[9].t34 161.106
R17940 XThR.Tn[9].n58 XThR.Tn[9].t62 161.106
R17941 XThR.Tn[9].n53 XThR.Tn[9].t24 161.106
R17942 XThR.Tn[9].n48 XThR.Tn[9].t66 161.106
R17943 XThR.Tn[9].n43 XThR.Tn[9].t45 161.106
R17944 XThR.Tn[9].n38 XThR.Tn[9].t32 161.106
R17945 XThR.Tn[9].n33 XThR.Tn[9].t37 161.106
R17946 XThR.Tn[9].n28 XThR.Tn[9].t23 161.106
R17947 XThR.Tn[9].n23 XThR.Tn[9].t46 161.106
R17948 XThR.Tn[9].n18 XThR.Tn[9].t21 161.106
R17949 XThR.Tn[9].n13 XThR.Tn[9].t64 161.106
R17950 XThR.Tn[9].n8 XThR.Tn[9].t28 161.106
R17951 XThR.Tn[9].n6 XThR.Tn[9].t71 161.106
R17952 XThR.Tn[9].n79 XThR.Tn[9].t54 159.978
R17953 XThR.Tn[9].n74 XThR.Tn[9].t61 159.978
R17954 XThR.Tn[9].n69 XThR.Tn[9].t43 159.978
R17955 XThR.Tn[9].n64 XThR.Tn[9].t27 159.978
R17956 XThR.Tn[9].n59 XThR.Tn[9].t52 159.978
R17957 XThR.Tn[9].n54 XThR.Tn[9].t18 159.978
R17958 XThR.Tn[9].n49 XThR.Tn[9].t60 159.978
R17959 XThR.Tn[9].n44 XThR.Tn[9].t40 159.978
R17960 XThR.Tn[9].n39 XThR.Tn[9].t25 159.978
R17961 XThR.Tn[9].n34 XThR.Tn[9].t33 159.978
R17962 XThR.Tn[9].n29 XThR.Tn[9].t16 159.978
R17963 XThR.Tn[9].n24 XThR.Tn[9].t42 159.978
R17964 XThR.Tn[9].n19 XThR.Tn[9].t15 159.978
R17965 XThR.Tn[9].n14 XThR.Tn[9].t59 159.978
R17966 XThR.Tn[9].n9 XThR.Tn[9].t19 159.978
R17967 XThR.Tn[9].n78 XThR.Tn[9].t49 145.038
R17968 XThR.Tn[9].n73 XThR.Tn[9].t14 145.038
R17969 XThR.Tn[9].n68 XThR.Tn[9].t57 145.038
R17970 XThR.Tn[9].n63 XThR.Tn[9].t38 145.038
R17971 XThR.Tn[9].n58 XThR.Tn[9].t70 145.038
R17972 XThR.Tn[9].n53 XThR.Tn[9].t48 145.038
R17973 XThR.Tn[9].n48 XThR.Tn[9].t58 145.038
R17974 XThR.Tn[9].n43 XThR.Tn[9].t39 145.038
R17975 XThR.Tn[9].n38 XThR.Tn[9].t36 145.038
R17976 XThR.Tn[9].n33 XThR.Tn[9].t67 145.038
R17977 XThR.Tn[9].n28 XThR.Tn[9].t31 145.038
R17978 XThR.Tn[9].n23 XThR.Tn[9].t56 145.038
R17979 XThR.Tn[9].n18 XThR.Tn[9].t29 145.038
R17980 XThR.Tn[9].n13 XThR.Tn[9].t72 145.038
R17981 XThR.Tn[9].n8 XThR.Tn[9].t35 145.038
R17982 XThR.Tn[9].n6 XThR.Tn[9].t17 145.038
R17983 XThR.Tn[9].n79 XThR.Tn[9].t68 143.911
R17984 XThR.Tn[9].n74 XThR.Tn[9].t30 143.911
R17985 XThR.Tn[9].n69 XThR.Tn[9].t12 143.911
R17986 XThR.Tn[9].n64 XThR.Tn[9].t53 143.911
R17987 XThR.Tn[9].n59 XThR.Tn[9].t22 143.911
R17988 XThR.Tn[9].n54 XThR.Tn[9].t65 143.911
R17989 XThR.Tn[9].n49 XThR.Tn[9].t13 143.911
R17990 XThR.Tn[9].n44 XThR.Tn[9].t55 143.911
R17991 XThR.Tn[9].n39 XThR.Tn[9].t51 143.911
R17992 XThR.Tn[9].n34 XThR.Tn[9].t20 143.911
R17993 XThR.Tn[9].n29 XThR.Tn[9].t44 143.911
R17994 XThR.Tn[9].n24 XThR.Tn[9].t73 143.911
R17995 XThR.Tn[9].n19 XThR.Tn[9].t41 143.911
R17996 XThR.Tn[9].n14 XThR.Tn[9].t26 143.911
R17997 XThR.Tn[9].n9 XThR.Tn[9].t50 143.911
R17998 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R17999 XThR.Tn[9].n0 XThR.Tn[9].t2 26.5955
R18000 XThR.Tn[9].n0 XThR.Tn[9].t0 26.5955
R18001 XThR.Tn[9].n85 XThR.Tn[9].t10 26.5955
R18002 XThR.Tn[9].n85 XThR.Tn[9].t8 26.5955
R18003 XThR.Tn[9].n86 XThR.Tn[9].t11 26.5955
R18004 XThR.Tn[9].n86 XThR.Tn[9].t9 26.5955
R18005 XThR.Tn[9].n1 XThR.Tn[9].t3 26.5955
R18006 XThR.Tn[9].n1 XThR.Tn[9].t1 26.5955
R18007 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R18008 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R18009 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R18010 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R18011 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R18012 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R18013 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R18014 XThR.Tn[9] XThR.Tn[9].n7 5.34038
R18015 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R18016 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R18017 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R18018 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R18019 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R18020 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R18021 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R18022 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R18023 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R18024 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R18025 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R18026 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R18027 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R18028 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R18029 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R18030 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R18031 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R18032 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R18033 XThR.Tn[9].n12 XThR.Tn[9] 2.52282
R18034 XThR.Tn[9].n17 XThR.Tn[9] 2.52282
R18035 XThR.Tn[9].n22 XThR.Tn[9] 2.52282
R18036 XThR.Tn[9].n27 XThR.Tn[9] 2.52282
R18037 XThR.Tn[9].n32 XThR.Tn[9] 2.52282
R18038 XThR.Tn[9].n37 XThR.Tn[9] 2.52282
R18039 XThR.Tn[9].n42 XThR.Tn[9] 2.52282
R18040 XThR.Tn[9].n47 XThR.Tn[9] 2.52282
R18041 XThR.Tn[9].n52 XThR.Tn[9] 2.52282
R18042 XThR.Tn[9].n57 XThR.Tn[9] 2.52282
R18043 XThR.Tn[9].n62 XThR.Tn[9] 2.52282
R18044 XThR.Tn[9].n67 XThR.Tn[9] 2.52282
R18045 XThR.Tn[9].n72 XThR.Tn[9] 2.52282
R18046 XThR.Tn[9].n77 XThR.Tn[9] 2.52282
R18047 XThR.Tn[9].n82 XThR.Tn[9] 2.52282
R18048 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R18049 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R18050 XThR.Tn[9].n80 XThR.Tn[9] 1.08677
R18051 XThR.Tn[9].n75 XThR.Tn[9] 1.08677
R18052 XThR.Tn[9].n70 XThR.Tn[9] 1.08677
R18053 XThR.Tn[9].n65 XThR.Tn[9] 1.08677
R18054 XThR.Tn[9].n60 XThR.Tn[9] 1.08677
R18055 XThR.Tn[9].n55 XThR.Tn[9] 1.08677
R18056 XThR.Tn[9].n50 XThR.Tn[9] 1.08677
R18057 XThR.Tn[9].n45 XThR.Tn[9] 1.08677
R18058 XThR.Tn[9].n40 XThR.Tn[9] 1.08677
R18059 XThR.Tn[9].n35 XThR.Tn[9] 1.08677
R18060 XThR.Tn[9].n30 XThR.Tn[9] 1.08677
R18061 XThR.Tn[9].n25 XThR.Tn[9] 1.08677
R18062 XThR.Tn[9].n20 XThR.Tn[9] 1.08677
R18063 XThR.Tn[9].n15 XThR.Tn[9] 1.08677
R18064 XThR.Tn[9].n10 XThR.Tn[9] 1.08677
R18065 XThR.Tn[9] XThR.Tn[9].n12 0.839786
R18066 XThR.Tn[9] XThR.Tn[9].n17 0.839786
R18067 XThR.Tn[9] XThR.Tn[9].n22 0.839786
R18068 XThR.Tn[9] XThR.Tn[9].n27 0.839786
R18069 XThR.Tn[9] XThR.Tn[9].n32 0.839786
R18070 XThR.Tn[9] XThR.Tn[9].n37 0.839786
R18071 XThR.Tn[9] XThR.Tn[9].n42 0.839786
R18072 XThR.Tn[9] XThR.Tn[9].n47 0.839786
R18073 XThR.Tn[9] XThR.Tn[9].n52 0.839786
R18074 XThR.Tn[9] XThR.Tn[9].n57 0.839786
R18075 XThR.Tn[9] XThR.Tn[9].n62 0.839786
R18076 XThR.Tn[9] XThR.Tn[9].n67 0.839786
R18077 XThR.Tn[9] XThR.Tn[9].n72 0.839786
R18078 XThR.Tn[9] XThR.Tn[9].n77 0.839786
R18079 XThR.Tn[9] XThR.Tn[9].n82 0.839786
R18080 XThR.Tn[9].n7 XThR.Tn[9] 0.499542
R18081 XThR.Tn[9].n81 XThR.Tn[9] 0.063
R18082 XThR.Tn[9].n76 XThR.Tn[9] 0.063
R18083 XThR.Tn[9].n71 XThR.Tn[9] 0.063
R18084 XThR.Tn[9].n66 XThR.Tn[9] 0.063
R18085 XThR.Tn[9].n61 XThR.Tn[9] 0.063
R18086 XThR.Tn[9].n56 XThR.Tn[9] 0.063
R18087 XThR.Tn[9].n51 XThR.Tn[9] 0.063
R18088 XThR.Tn[9].n46 XThR.Tn[9] 0.063
R18089 XThR.Tn[9].n41 XThR.Tn[9] 0.063
R18090 XThR.Tn[9].n36 XThR.Tn[9] 0.063
R18091 XThR.Tn[9].n31 XThR.Tn[9] 0.063
R18092 XThR.Tn[9].n26 XThR.Tn[9] 0.063
R18093 XThR.Tn[9].n21 XThR.Tn[9] 0.063
R18094 XThR.Tn[9].n16 XThR.Tn[9] 0.063
R18095 XThR.Tn[9].n11 XThR.Tn[9] 0.063
R18096 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R18097 XThR.Tn[9] XThR.Tn[9].n83 0.038
R18098 XThR.Tn[9].n7 XThR.Tn[9] 0.0143889
R18099 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00771154
R18100 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00771154
R18101 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00771154
R18102 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00771154
R18103 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00771154
R18104 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00771154
R18105 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00771154
R18106 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00771154
R18107 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00771154
R18108 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00771154
R18109 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00771154
R18110 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00771154
R18111 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00771154
R18112 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00771154
R18113 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00771154
R18114 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18115 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18116 XThC.Tn[5].n71 XThC.Tn[5].n69 161.365
R18117 XThC.Tn[5].n67 XThC.Tn[5].n65 161.365
R18118 XThC.Tn[5].n63 XThC.Tn[5].n61 161.365
R18119 XThC.Tn[5].n59 XThC.Tn[5].n57 161.365
R18120 XThC.Tn[5].n55 XThC.Tn[5].n53 161.365
R18121 XThC.Tn[5].n51 XThC.Tn[5].n49 161.365
R18122 XThC.Tn[5].n47 XThC.Tn[5].n45 161.365
R18123 XThC.Tn[5].n43 XThC.Tn[5].n41 161.365
R18124 XThC.Tn[5].n39 XThC.Tn[5].n37 161.365
R18125 XThC.Tn[5].n35 XThC.Tn[5].n33 161.365
R18126 XThC.Tn[5].n31 XThC.Tn[5].n29 161.365
R18127 XThC.Tn[5].n27 XThC.Tn[5].n25 161.365
R18128 XThC.Tn[5].n23 XThC.Tn[5].n21 161.365
R18129 XThC.Tn[5].n19 XThC.Tn[5].n17 161.365
R18130 XThC.Tn[5].n15 XThC.Tn[5].n13 161.365
R18131 XThC.Tn[5].n12 XThC.Tn[5].n10 161.365
R18132 XThC.Tn[5].n69 XThC.Tn[5].t41 161.202
R18133 XThC.Tn[5].n65 XThC.Tn[5].t30 161.202
R18134 XThC.Tn[5].n61 XThC.Tn[5].t18 161.202
R18135 XThC.Tn[5].n57 XThC.Tn[5].t16 161.202
R18136 XThC.Tn[5].n53 XThC.Tn[5].t39 161.202
R18137 XThC.Tn[5].n49 XThC.Tn[5].t26 161.202
R18138 XThC.Tn[5].n45 XThC.Tn[5].t25 161.202
R18139 XThC.Tn[5].n41 XThC.Tn[5].t37 161.202
R18140 XThC.Tn[5].n37 XThC.Tn[5].t35 161.202
R18141 XThC.Tn[5].n33 XThC.Tn[5].t27 161.202
R18142 XThC.Tn[5].n29 XThC.Tn[5].t14 161.202
R18143 XThC.Tn[5].n25 XThC.Tn[5].t13 161.202
R18144 XThC.Tn[5].n21 XThC.Tn[5].t24 161.202
R18145 XThC.Tn[5].n17 XThC.Tn[5].t23 161.202
R18146 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18147 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18148 XThC.Tn[5].n69 XThC.Tn[5].t22 145.137
R18149 XThC.Tn[5].n65 XThC.Tn[5].t12 145.137
R18150 XThC.Tn[5].n61 XThC.Tn[5].t32 145.137
R18151 XThC.Tn[5].n57 XThC.Tn[5].t31 145.137
R18152 XThC.Tn[5].n53 XThC.Tn[5].t21 145.137
R18153 XThC.Tn[5].n49 XThC.Tn[5].t42 145.137
R18154 XThC.Tn[5].n45 XThC.Tn[5].t40 145.137
R18155 XThC.Tn[5].n41 XThC.Tn[5].t20 145.137
R18156 XThC.Tn[5].n37 XThC.Tn[5].t17 145.137
R18157 XThC.Tn[5].n33 XThC.Tn[5].t43 145.137
R18158 XThC.Tn[5].n29 XThC.Tn[5].t29 145.137
R18159 XThC.Tn[5].n25 XThC.Tn[5].t28 145.137
R18160 XThC.Tn[5].n21 XThC.Tn[5].t38 145.137
R18161 XThC.Tn[5].n17 XThC.Tn[5].t36 145.137
R18162 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18163 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18164 XThC.Tn[5].n6 XThC.Tn[5].n4 135.249
R18165 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18166 XThC.Tn[5].n6 XThC.Tn[5].n5 98.981
R18167 XThC.Tn[5].n8 XThC.Tn[5].n7 98.981
R18168 XThC.Tn[5].n8 XThC.Tn[5].n6 36.2672
R18169 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18170 XThC.Tn[5].n73 XThC.Tn[5].n9 32.6405
R18171 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R18172 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R18173 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R18174 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R18175 XThC.Tn[5].n3 XThC.Tn[5].t1 24.9236
R18176 XThC.Tn[5].n3 XThC.Tn[5].t0 24.9236
R18177 XThC.Tn[5].n4 XThC.Tn[5].t8 24.9236
R18178 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R18179 XThC.Tn[5].n5 XThC.Tn[5].t10 24.9236
R18180 XThC.Tn[5].n5 XThC.Tn[5].t9 24.9236
R18181 XThC.Tn[5].n7 XThC.Tn[5].t3 24.9236
R18182 XThC.Tn[5].n7 XThC.Tn[5].t2 24.9236
R18183 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18184 XThC.Tn[5] XThC.Tn[5].n12 8.0245
R18185 XThC.Tn[5].n72 XThC.Tn[5].n71 7.9105
R18186 XThC.Tn[5].n68 XThC.Tn[5].n67 7.9105
R18187 XThC.Tn[5].n64 XThC.Tn[5].n63 7.9105
R18188 XThC.Tn[5].n60 XThC.Tn[5].n59 7.9105
R18189 XThC.Tn[5].n56 XThC.Tn[5].n55 7.9105
R18190 XThC.Tn[5].n52 XThC.Tn[5].n51 7.9105
R18191 XThC.Tn[5].n48 XThC.Tn[5].n47 7.9105
R18192 XThC.Tn[5].n44 XThC.Tn[5].n43 7.9105
R18193 XThC.Tn[5].n40 XThC.Tn[5].n39 7.9105
R18194 XThC.Tn[5].n36 XThC.Tn[5].n35 7.9105
R18195 XThC.Tn[5].n32 XThC.Tn[5].n31 7.9105
R18196 XThC.Tn[5].n28 XThC.Tn[5].n27 7.9105
R18197 XThC.Tn[5].n24 XThC.Tn[5].n23 7.9105
R18198 XThC.Tn[5].n20 XThC.Tn[5].n19 7.9105
R18199 XThC.Tn[5].n16 XThC.Tn[5].n15 7.9105
R18200 XThC.Tn[5] XThC.Tn[5].n73 6.7205
R18201 XThC.Tn[5].n73 XThC.Tn[5] 5.69842
R18202 XThC.Tn[5].n16 XThC.Tn[5] 0.235138
R18203 XThC.Tn[5].n20 XThC.Tn[5] 0.235138
R18204 XThC.Tn[5].n24 XThC.Tn[5] 0.235138
R18205 XThC.Tn[5].n28 XThC.Tn[5] 0.235138
R18206 XThC.Tn[5].n32 XThC.Tn[5] 0.235138
R18207 XThC.Tn[5].n36 XThC.Tn[5] 0.235138
R18208 XThC.Tn[5].n40 XThC.Tn[5] 0.235138
R18209 XThC.Tn[5].n44 XThC.Tn[5] 0.235138
R18210 XThC.Tn[5].n48 XThC.Tn[5] 0.235138
R18211 XThC.Tn[5].n52 XThC.Tn[5] 0.235138
R18212 XThC.Tn[5].n56 XThC.Tn[5] 0.235138
R18213 XThC.Tn[5].n60 XThC.Tn[5] 0.235138
R18214 XThC.Tn[5].n64 XThC.Tn[5] 0.235138
R18215 XThC.Tn[5].n68 XThC.Tn[5] 0.235138
R18216 XThC.Tn[5].n72 XThC.Tn[5] 0.235138
R18217 XThC.Tn[5] XThC.Tn[5].n16 0.114505
R18218 XThC.Tn[5] XThC.Tn[5].n20 0.114505
R18219 XThC.Tn[5] XThC.Tn[5].n24 0.114505
R18220 XThC.Tn[5] XThC.Tn[5].n28 0.114505
R18221 XThC.Tn[5] XThC.Tn[5].n32 0.114505
R18222 XThC.Tn[5] XThC.Tn[5].n36 0.114505
R18223 XThC.Tn[5] XThC.Tn[5].n40 0.114505
R18224 XThC.Tn[5] XThC.Tn[5].n44 0.114505
R18225 XThC.Tn[5] XThC.Tn[5].n48 0.114505
R18226 XThC.Tn[5] XThC.Tn[5].n52 0.114505
R18227 XThC.Tn[5] XThC.Tn[5].n56 0.114505
R18228 XThC.Tn[5] XThC.Tn[5].n60 0.114505
R18229 XThC.Tn[5] XThC.Tn[5].n64 0.114505
R18230 XThC.Tn[5] XThC.Tn[5].n68 0.114505
R18231 XThC.Tn[5] XThC.Tn[5].n72 0.114505
R18232 XThC.Tn[5].n71 XThC.Tn[5].n70 0.0599512
R18233 XThC.Tn[5].n67 XThC.Tn[5].n66 0.0599512
R18234 XThC.Tn[5].n63 XThC.Tn[5].n62 0.0599512
R18235 XThC.Tn[5].n59 XThC.Tn[5].n58 0.0599512
R18236 XThC.Tn[5].n55 XThC.Tn[5].n54 0.0599512
R18237 XThC.Tn[5].n51 XThC.Tn[5].n50 0.0599512
R18238 XThC.Tn[5].n47 XThC.Tn[5].n46 0.0599512
R18239 XThC.Tn[5].n43 XThC.Tn[5].n42 0.0599512
R18240 XThC.Tn[5].n39 XThC.Tn[5].n38 0.0599512
R18241 XThC.Tn[5].n35 XThC.Tn[5].n34 0.0599512
R18242 XThC.Tn[5].n31 XThC.Tn[5].n30 0.0599512
R18243 XThC.Tn[5].n27 XThC.Tn[5].n26 0.0599512
R18244 XThC.Tn[5].n23 XThC.Tn[5].n22 0.0599512
R18245 XThC.Tn[5].n19 XThC.Tn[5].n18 0.0599512
R18246 XThC.Tn[5].n15 XThC.Tn[5].n14 0.0599512
R18247 XThC.Tn[5].n12 XThC.Tn[5].n11 0.0599512
R18248 XThC.Tn[5].n70 XThC.Tn[5] 0.0469286
R18249 XThC.Tn[5].n66 XThC.Tn[5] 0.0469286
R18250 XThC.Tn[5].n62 XThC.Tn[5] 0.0469286
R18251 XThC.Tn[5].n58 XThC.Tn[5] 0.0469286
R18252 XThC.Tn[5].n54 XThC.Tn[5] 0.0469286
R18253 XThC.Tn[5].n50 XThC.Tn[5] 0.0469286
R18254 XThC.Tn[5].n46 XThC.Tn[5] 0.0469286
R18255 XThC.Tn[5].n42 XThC.Tn[5] 0.0469286
R18256 XThC.Tn[5].n38 XThC.Tn[5] 0.0469286
R18257 XThC.Tn[5].n34 XThC.Tn[5] 0.0469286
R18258 XThC.Tn[5].n30 XThC.Tn[5] 0.0469286
R18259 XThC.Tn[5].n26 XThC.Tn[5] 0.0469286
R18260 XThC.Tn[5].n22 XThC.Tn[5] 0.0469286
R18261 XThC.Tn[5].n18 XThC.Tn[5] 0.0469286
R18262 XThC.Tn[5].n14 XThC.Tn[5] 0.0469286
R18263 XThC.Tn[5].n11 XThC.Tn[5] 0.0469286
R18264 XThC.Tn[5].n70 XThC.Tn[5] 0.0401341
R18265 XThC.Tn[5].n66 XThC.Tn[5] 0.0401341
R18266 XThC.Tn[5].n62 XThC.Tn[5] 0.0401341
R18267 XThC.Tn[5].n58 XThC.Tn[5] 0.0401341
R18268 XThC.Tn[5].n54 XThC.Tn[5] 0.0401341
R18269 XThC.Tn[5].n50 XThC.Tn[5] 0.0401341
R18270 XThC.Tn[5].n46 XThC.Tn[5] 0.0401341
R18271 XThC.Tn[5].n42 XThC.Tn[5] 0.0401341
R18272 XThC.Tn[5].n38 XThC.Tn[5] 0.0401341
R18273 XThC.Tn[5].n34 XThC.Tn[5] 0.0401341
R18274 XThC.Tn[5].n30 XThC.Tn[5] 0.0401341
R18275 XThC.Tn[5].n26 XThC.Tn[5] 0.0401341
R18276 XThC.Tn[5].n22 XThC.Tn[5] 0.0401341
R18277 XThC.Tn[5].n18 XThC.Tn[5] 0.0401341
R18278 XThC.Tn[5].n14 XThC.Tn[5] 0.0401341
R18279 XThC.Tn[5].n11 XThC.Tn[5] 0.0401341
R18280 XThC.Tn[9].n70 XThC.Tn[9].n69 265.341
R18281 XThC.Tn[9].n74 XThC.Tn[9].n72 243.68
R18282 XThC.Tn[9].n2 XThC.Tn[9].n0 241.847
R18283 XThC.Tn[9].n74 XThC.Tn[9].n73 205.28
R18284 XThC.Tn[9].n70 XThC.Tn[9].n68 202.094
R18285 XThC.Tn[9].n2 XThC.Tn[9].n1 185
R18286 XThC.Tn[9].n64 XThC.Tn[9].n62 161.365
R18287 XThC.Tn[9].n60 XThC.Tn[9].n58 161.365
R18288 XThC.Tn[9].n56 XThC.Tn[9].n54 161.365
R18289 XThC.Tn[9].n52 XThC.Tn[9].n50 161.365
R18290 XThC.Tn[9].n48 XThC.Tn[9].n46 161.365
R18291 XThC.Tn[9].n44 XThC.Tn[9].n42 161.365
R18292 XThC.Tn[9].n40 XThC.Tn[9].n38 161.365
R18293 XThC.Tn[9].n36 XThC.Tn[9].n34 161.365
R18294 XThC.Tn[9].n32 XThC.Tn[9].n30 161.365
R18295 XThC.Tn[9].n28 XThC.Tn[9].n26 161.365
R18296 XThC.Tn[9].n24 XThC.Tn[9].n22 161.365
R18297 XThC.Tn[9].n20 XThC.Tn[9].n18 161.365
R18298 XThC.Tn[9].n16 XThC.Tn[9].n14 161.365
R18299 XThC.Tn[9].n12 XThC.Tn[9].n10 161.365
R18300 XThC.Tn[9].n8 XThC.Tn[9].n6 161.365
R18301 XThC.Tn[9].n5 XThC.Tn[9].n3 161.365
R18302 XThC.Tn[9].n62 XThC.Tn[9].t20 161.202
R18303 XThC.Tn[9].n58 XThC.Tn[9].t41 161.202
R18304 XThC.Tn[9].n54 XThC.Tn[9].t29 161.202
R18305 XThC.Tn[9].n50 XThC.Tn[9].t27 161.202
R18306 XThC.Tn[9].n46 XThC.Tn[9].t18 161.202
R18307 XThC.Tn[9].n42 XThC.Tn[9].t37 161.202
R18308 XThC.Tn[9].n38 XThC.Tn[9].t36 161.202
R18309 XThC.Tn[9].n34 XThC.Tn[9].t16 161.202
R18310 XThC.Tn[9].n30 XThC.Tn[9].t14 161.202
R18311 XThC.Tn[9].n26 XThC.Tn[9].t38 161.202
R18312 XThC.Tn[9].n22 XThC.Tn[9].t25 161.202
R18313 XThC.Tn[9].n18 XThC.Tn[9].t24 161.202
R18314 XThC.Tn[9].n14 XThC.Tn[9].t35 161.202
R18315 XThC.Tn[9].n10 XThC.Tn[9].t34 161.202
R18316 XThC.Tn[9].n6 XThC.Tn[9].t30 161.202
R18317 XThC.Tn[9].n3 XThC.Tn[9].t12 161.202
R18318 XThC.Tn[9].n62 XThC.Tn[9].t33 145.137
R18319 XThC.Tn[9].n58 XThC.Tn[9].t23 145.137
R18320 XThC.Tn[9].n54 XThC.Tn[9].t43 145.137
R18321 XThC.Tn[9].n50 XThC.Tn[9].t42 145.137
R18322 XThC.Tn[9].n46 XThC.Tn[9].t32 145.137
R18323 XThC.Tn[9].n42 XThC.Tn[9].t21 145.137
R18324 XThC.Tn[9].n38 XThC.Tn[9].t19 145.137
R18325 XThC.Tn[9].n34 XThC.Tn[9].t31 145.137
R18326 XThC.Tn[9].n30 XThC.Tn[9].t28 145.137
R18327 XThC.Tn[9].n26 XThC.Tn[9].t22 145.137
R18328 XThC.Tn[9].n22 XThC.Tn[9].t40 145.137
R18329 XThC.Tn[9].n18 XThC.Tn[9].t39 145.137
R18330 XThC.Tn[9].n14 XThC.Tn[9].t17 145.137
R18331 XThC.Tn[9].n10 XThC.Tn[9].t15 145.137
R18332 XThC.Tn[9].n6 XThC.Tn[9].t13 145.137
R18333 XThC.Tn[9].n3 XThC.Tn[9].t26 145.137
R18334 XThC.Tn[9].n72 XThC.Tn[9].t1 26.5955
R18335 XThC.Tn[9].n72 XThC.Tn[9].t0 26.5955
R18336 XThC.Tn[9].n69 XThC.Tn[9].t10 26.5955
R18337 XThC.Tn[9].n69 XThC.Tn[9].t9 26.5955
R18338 XThC.Tn[9].n68 XThC.Tn[9].t8 26.5955
R18339 XThC.Tn[9].n68 XThC.Tn[9].t11 26.5955
R18340 XThC.Tn[9].n73 XThC.Tn[9].t3 26.5955
R18341 XThC.Tn[9].n73 XThC.Tn[9].t2 26.5955
R18342 XThC.Tn[9].n1 XThC.Tn[9].t6 24.9236
R18343 XThC.Tn[9].n1 XThC.Tn[9].t7 24.9236
R18344 XThC.Tn[9].n0 XThC.Tn[9].t5 24.9236
R18345 XThC.Tn[9].n0 XThC.Tn[9].t4 24.9236
R18346 XThC.Tn[9] XThC.Tn[9].n74 22.9652
R18347 XThC.Tn[9] XThC.Tn[9].n2 18.8943
R18348 XThC.Tn[9].n71 XThC.Tn[9].n70 13.9299
R18349 XThC.Tn[9] XThC.Tn[9].n71 13.9299
R18350 XThC.Tn[9] XThC.Tn[9].n5 8.0245
R18351 XThC.Tn[9].n65 XThC.Tn[9].n64 7.9105
R18352 XThC.Tn[9].n61 XThC.Tn[9].n60 7.9105
R18353 XThC.Tn[9].n57 XThC.Tn[9].n56 7.9105
R18354 XThC.Tn[9].n53 XThC.Tn[9].n52 7.9105
R18355 XThC.Tn[9].n49 XThC.Tn[9].n48 7.9105
R18356 XThC.Tn[9].n45 XThC.Tn[9].n44 7.9105
R18357 XThC.Tn[9].n41 XThC.Tn[9].n40 7.9105
R18358 XThC.Tn[9].n37 XThC.Tn[9].n36 7.9105
R18359 XThC.Tn[9].n33 XThC.Tn[9].n32 7.9105
R18360 XThC.Tn[9].n29 XThC.Tn[9].n28 7.9105
R18361 XThC.Tn[9].n25 XThC.Tn[9].n24 7.9105
R18362 XThC.Tn[9].n21 XThC.Tn[9].n20 7.9105
R18363 XThC.Tn[9].n17 XThC.Tn[9].n16 7.9105
R18364 XThC.Tn[9].n13 XThC.Tn[9].n12 7.9105
R18365 XThC.Tn[9].n9 XThC.Tn[9].n8 7.9105
R18366 XThC.Tn[9].n67 XThC.Tn[9].n66 7.44831
R18367 XThC.Tn[9].n67 XThC.Tn[9] 6.34069
R18368 XThC.Tn[9].n66 XThC.Tn[9] 4.25199
R18369 XThC.Tn[9] XThC.Tn[9].n67 1.79489
R18370 XThC.Tn[9].n71 XThC.Tn[9] 1.19676
R18371 XThC.Tn[9].n66 XThC.Tn[9] 0.657022
R18372 XThC.Tn[9].n9 XThC.Tn[9] 0.235138
R18373 XThC.Tn[9].n13 XThC.Tn[9] 0.235138
R18374 XThC.Tn[9].n17 XThC.Tn[9] 0.235138
R18375 XThC.Tn[9].n21 XThC.Tn[9] 0.235138
R18376 XThC.Tn[9].n25 XThC.Tn[9] 0.235138
R18377 XThC.Tn[9].n29 XThC.Tn[9] 0.235138
R18378 XThC.Tn[9].n33 XThC.Tn[9] 0.235138
R18379 XThC.Tn[9].n37 XThC.Tn[9] 0.235138
R18380 XThC.Tn[9].n41 XThC.Tn[9] 0.235138
R18381 XThC.Tn[9].n45 XThC.Tn[9] 0.235138
R18382 XThC.Tn[9].n49 XThC.Tn[9] 0.235138
R18383 XThC.Tn[9].n53 XThC.Tn[9] 0.235138
R18384 XThC.Tn[9].n57 XThC.Tn[9] 0.235138
R18385 XThC.Tn[9].n61 XThC.Tn[9] 0.235138
R18386 XThC.Tn[9].n65 XThC.Tn[9] 0.235138
R18387 XThC.Tn[9] XThC.Tn[9].n9 0.114505
R18388 XThC.Tn[9] XThC.Tn[9].n13 0.114505
R18389 XThC.Tn[9] XThC.Tn[9].n17 0.114505
R18390 XThC.Tn[9] XThC.Tn[9].n21 0.114505
R18391 XThC.Tn[9] XThC.Tn[9].n25 0.114505
R18392 XThC.Tn[9] XThC.Tn[9].n29 0.114505
R18393 XThC.Tn[9] XThC.Tn[9].n33 0.114505
R18394 XThC.Tn[9] XThC.Tn[9].n37 0.114505
R18395 XThC.Tn[9] XThC.Tn[9].n41 0.114505
R18396 XThC.Tn[9] XThC.Tn[9].n45 0.114505
R18397 XThC.Tn[9] XThC.Tn[9].n49 0.114505
R18398 XThC.Tn[9] XThC.Tn[9].n53 0.114505
R18399 XThC.Tn[9] XThC.Tn[9].n57 0.114505
R18400 XThC.Tn[9] XThC.Tn[9].n61 0.114505
R18401 XThC.Tn[9] XThC.Tn[9].n65 0.114505
R18402 XThC.Tn[9].n64 XThC.Tn[9].n63 0.0599512
R18403 XThC.Tn[9].n60 XThC.Tn[9].n59 0.0599512
R18404 XThC.Tn[9].n56 XThC.Tn[9].n55 0.0599512
R18405 XThC.Tn[9].n52 XThC.Tn[9].n51 0.0599512
R18406 XThC.Tn[9].n48 XThC.Tn[9].n47 0.0599512
R18407 XThC.Tn[9].n44 XThC.Tn[9].n43 0.0599512
R18408 XThC.Tn[9].n40 XThC.Tn[9].n39 0.0599512
R18409 XThC.Tn[9].n36 XThC.Tn[9].n35 0.0599512
R18410 XThC.Tn[9].n32 XThC.Tn[9].n31 0.0599512
R18411 XThC.Tn[9].n28 XThC.Tn[9].n27 0.0599512
R18412 XThC.Tn[9].n24 XThC.Tn[9].n23 0.0599512
R18413 XThC.Tn[9].n20 XThC.Tn[9].n19 0.0599512
R18414 XThC.Tn[9].n16 XThC.Tn[9].n15 0.0599512
R18415 XThC.Tn[9].n12 XThC.Tn[9].n11 0.0599512
R18416 XThC.Tn[9].n8 XThC.Tn[9].n7 0.0599512
R18417 XThC.Tn[9].n5 XThC.Tn[9].n4 0.0599512
R18418 XThC.Tn[9].n63 XThC.Tn[9] 0.0469286
R18419 XThC.Tn[9].n59 XThC.Tn[9] 0.0469286
R18420 XThC.Tn[9].n55 XThC.Tn[9] 0.0469286
R18421 XThC.Tn[9].n51 XThC.Tn[9] 0.0469286
R18422 XThC.Tn[9].n47 XThC.Tn[9] 0.0469286
R18423 XThC.Tn[9].n43 XThC.Tn[9] 0.0469286
R18424 XThC.Tn[9].n39 XThC.Tn[9] 0.0469286
R18425 XThC.Tn[9].n35 XThC.Tn[9] 0.0469286
R18426 XThC.Tn[9].n31 XThC.Tn[9] 0.0469286
R18427 XThC.Tn[9].n27 XThC.Tn[9] 0.0469286
R18428 XThC.Tn[9].n23 XThC.Tn[9] 0.0469286
R18429 XThC.Tn[9].n19 XThC.Tn[9] 0.0469286
R18430 XThC.Tn[9].n15 XThC.Tn[9] 0.0469286
R18431 XThC.Tn[9].n11 XThC.Tn[9] 0.0469286
R18432 XThC.Tn[9].n7 XThC.Tn[9] 0.0469286
R18433 XThC.Tn[9].n4 XThC.Tn[9] 0.0469286
R18434 XThC.Tn[9].n63 XThC.Tn[9] 0.0401341
R18435 XThC.Tn[9].n59 XThC.Tn[9] 0.0401341
R18436 XThC.Tn[9].n55 XThC.Tn[9] 0.0401341
R18437 XThC.Tn[9].n51 XThC.Tn[9] 0.0401341
R18438 XThC.Tn[9].n47 XThC.Tn[9] 0.0401341
R18439 XThC.Tn[9].n43 XThC.Tn[9] 0.0401341
R18440 XThC.Tn[9].n39 XThC.Tn[9] 0.0401341
R18441 XThC.Tn[9].n35 XThC.Tn[9] 0.0401341
R18442 XThC.Tn[9].n31 XThC.Tn[9] 0.0401341
R18443 XThC.Tn[9].n27 XThC.Tn[9] 0.0401341
R18444 XThC.Tn[9].n23 XThC.Tn[9] 0.0401341
R18445 XThC.Tn[9].n19 XThC.Tn[9] 0.0401341
R18446 XThC.Tn[9].n15 XThC.Tn[9] 0.0401341
R18447 XThC.Tn[9].n11 XThC.Tn[9] 0.0401341
R18448 XThC.Tn[9].n7 XThC.Tn[9] 0.0401341
R18449 XThC.Tn[9].n4 XThC.Tn[9] 0.0401341
R18450 XThC.Tn[11].n70 XThC.Tn[11].n69 265.341
R18451 XThC.Tn[11].n74 XThC.Tn[11].n72 243.68
R18452 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R18453 XThC.Tn[11].n74 XThC.Tn[11].n73 205.28
R18454 XThC.Tn[11].n70 XThC.Tn[11].n68 202.094
R18455 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R18456 XThC.Tn[11].n64 XThC.Tn[11].n62 161.365
R18457 XThC.Tn[11].n60 XThC.Tn[11].n58 161.365
R18458 XThC.Tn[11].n56 XThC.Tn[11].n54 161.365
R18459 XThC.Tn[11].n52 XThC.Tn[11].n50 161.365
R18460 XThC.Tn[11].n48 XThC.Tn[11].n46 161.365
R18461 XThC.Tn[11].n44 XThC.Tn[11].n42 161.365
R18462 XThC.Tn[11].n40 XThC.Tn[11].n38 161.365
R18463 XThC.Tn[11].n36 XThC.Tn[11].n34 161.365
R18464 XThC.Tn[11].n32 XThC.Tn[11].n30 161.365
R18465 XThC.Tn[11].n28 XThC.Tn[11].n26 161.365
R18466 XThC.Tn[11].n24 XThC.Tn[11].n22 161.365
R18467 XThC.Tn[11].n20 XThC.Tn[11].n18 161.365
R18468 XThC.Tn[11].n16 XThC.Tn[11].n14 161.365
R18469 XThC.Tn[11].n12 XThC.Tn[11].n10 161.365
R18470 XThC.Tn[11].n8 XThC.Tn[11].n6 161.365
R18471 XThC.Tn[11].n5 XThC.Tn[11].n3 161.365
R18472 XThC.Tn[11].n62 XThC.Tn[11].t24 161.202
R18473 XThC.Tn[11].n58 XThC.Tn[11].t14 161.202
R18474 XThC.Tn[11].n54 XThC.Tn[11].t33 161.202
R18475 XThC.Tn[11].n50 XThC.Tn[11].t30 161.202
R18476 XThC.Tn[11].n46 XThC.Tn[11].t22 161.202
R18477 XThC.Tn[11].n42 XThC.Tn[11].t41 161.202
R18478 XThC.Tn[11].n38 XThC.Tn[11].t40 161.202
R18479 XThC.Tn[11].n34 XThC.Tn[11].t21 161.202
R18480 XThC.Tn[11].n30 XThC.Tn[11].t19 161.202
R18481 XThC.Tn[11].n26 XThC.Tn[11].t42 161.202
R18482 XThC.Tn[11].n22 XThC.Tn[11].t29 161.202
R18483 XThC.Tn[11].n18 XThC.Tn[11].t28 161.202
R18484 XThC.Tn[11].n14 XThC.Tn[11].t39 161.202
R18485 XThC.Tn[11].n10 XThC.Tn[11].t37 161.202
R18486 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R18487 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R18488 XThC.Tn[11].n62 XThC.Tn[11].t27 145.137
R18489 XThC.Tn[11].n58 XThC.Tn[11].t17 145.137
R18490 XThC.Tn[11].n54 XThC.Tn[11].t36 145.137
R18491 XThC.Tn[11].n50 XThC.Tn[11].t34 145.137
R18492 XThC.Tn[11].n46 XThC.Tn[11].t26 145.137
R18493 XThC.Tn[11].n42 XThC.Tn[11].t15 145.137
R18494 XThC.Tn[11].n38 XThC.Tn[11].t13 145.137
R18495 XThC.Tn[11].n34 XThC.Tn[11].t25 145.137
R18496 XThC.Tn[11].n30 XThC.Tn[11].t23 145.137
R18497 XThC.Tn[11].n26 XThC.Tn[11].t16 145.137
R18498 XThC.Tn[11].n22 XThC.Tn[11].t32 145.137
R18499 XThC.Tn[11].n18 XThC.Tn[11].t31 145.137
R18500 XThC.Tn[11].n14 XThC.Tn[11].t12 145.137
R18501 XThC.Tn[11].n10 XThC.Tn[11].t43 145.137
R18502 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R18503 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R18504 XThC.Tn[11].n69 XThC.Tn[11].t7 26.5955
R18505 XThC.Tn[11].n69 XThC.Tn[11].t9 26.5955
R18506 XThC.Tn[11].n72 XThC.Tn[11].t2 26.5955
R18507 XThC.Tn[11].n72 XThC.Tn[11].t5 26.5955
R18508 XThC.Tn[11].n73 XThC.Tn[11].t4 26.5955
R18509 XThC.Tn[11].n73 XThC.Tn[11].t3 26.5955
R18510 XThC.Tn[11].n68 XThC.Tn[11].t11 26.5955
R18511 XThC.Tn[11].n68 XThC.Tn[11].t0 26.5955
R18512 XThC.Tn[11].n1 XThC.Tn[11].t6 24.9236
R18513 XThC.Tn[11].n1 XThC.Tn[11].t10 24.9236
R18514 XThC.Tn[11].n0 XThC.Tn[11].t8 24.9236
R18515 XThC.Tn[11].n0 XThC.Tn[11].t1 24.9236
R18516 XThC.Tn[11] XThC.Tn[11].n74 22.9652
R18517 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R18518 XThC.Tn[11].n71 XThC.Tn[11].n70 13.9299
R18519 XThC.Tn[11] XThC.Tn[11].n71 13.9299
R18520 XThC.Tn[11] XThC.Tn[11].n5 8.0245
R18521 XThC.Tn[11].n65 XThC.Tn[11].n64 7.9105
R18522 XThC.Tn[11].n61 XThC.Tn[11].n60 7.9105
R18523 XThC.Tn[11].n57 XThC.Tn[11].n56 7.9105
R18524 XThC.Tn[11].n53 XThC.Tn[11].n52 7.9105
R18525 XThC.Tn[11].n49 XThC.Tn[11].n48 7.9105
R18526 XThC.Tn[11].n45 XThC.Tn[11].n44 7.9105
R18527 XThC.Tn[11].n41 XThC.Tn[11].n40 7.9105
R18528 XThC.Tn[11].n37 XThC.Tn[11].n36 7.9105
R18529 XThC.Tn[11].n33 XThC.Tn[11].n32 7.9105
R18530 XThC.Tn[11].n29 XThC.Tn[11].n28 7.9105
R18531 XThC.Tn[11].n25 XThC.Tn[11].n24 7.9105
R18532 XThC.Tn[11].n21 XThC.Tn[11].n20 7.9105
R18533 XThC.Tn[11].n17 XThC.Tn[11].n16 7.9105
R18534 XThC.Tn[11].n13 XThC.Tn[11].n12 7.9105
R18535 XThC.Tn[11].n9 XThC.Tn[11].n8 7.9105
R18536 XThC.Tn[11].n67 XThC.Tn[11].n66 7.44831
R18537 XThC.Tn[11].n67 XThC.Tn[11] 6.34069
R18538 XThC.Tn[11].n66 XThC.Tn[11] 4.37928
R18539 XThC.Tn[11] XThC.Tn[11].n67 1.79489
R18540 XThC.Tn[11].n71 XThC.Tn[11] 1.19676
R18541 XThC.Tn[11].n66 XThC.Tn[11] 1.0918
R18542 XThC.Tn[11].n9 XThC.Tn[11] 0.235138
R18543 XThC.Tn[11].n13 XThC.Tn[11] 0.235138
R18544 XThC.Tn[11].n17 XThC.Tn[11] 0.235138
R18545 XThC.Tn[11].n21 XThC.Tn[11] 0.235138
R18546 XThC.Tn[11].n25 XThC.Tn[11] 0.235138
R18547 XThC.Tn[11].n29 XThC.Tn[11] 0.235138
R18548 XThC.Tn[11].n33 XThC.Tn[11] 0.235138
R18549 XThC.Tn[11].n37 XThC.Tn[11] 0.235138
R18550 XThC.Tn[11].n41 XThC.Tn[11] 0.235138
R18551 XThC.Tn[11].n45 XThC.Tn[11] 0.235138
R18552 XThC.Tn[11].n49 XThC.Tn[11] 0.235138
R18553 XThC.Tn[11].n53 XThC.Tn[11] 0.235138
R18554 XThC.Tn[11].n57 XThC.Tn[11] 0.235138
R18555 XThC.Tn[11].n61 XThC.Tn[11] 0.235138
R18556 XThC.Tn[11].n65 XThC.Tn[11] 0.235138
R18557 XThC.Tn[11] XThC.Tn[11].n9 0.114505
R18558 XThC.Tn[11] XThC.Tn[11].n13 0.114505
R18559 XThC.Tn[11] XThC.Tn[11].n17 0.114505
R18560 XThC.Tn[11] XThC.Tn[11].n21 0.114505
R18561 XThC.Tn[11] XThC.Tn[11].n25 0.114505
R18562 XThC.Tn[11] XThC.Tn[11].n29 0.114505
R18563 XThC.Tn[11] XThC.Tn[11].n33 0.114505
R18564 XThC.Tn[11] XThC.Tn[11].n37 0.114505
R18565 XThC.Tn[11] XThC.Tn[11].n41 0.114505
R18566 XThC.Tn[11] XThC.Tn[11].n45 0.114505
R18567 XThC.Tn[11] XThC.Tn[11].n49 0.114505
R18568 XThC.Tn[11] XThC.Tn[11].n53 0.114505
R18569 XThC.Tn[11] XThC.Tn[11].n57 0.114505
R18570 XThC.Tn[11] XThC.Tn[11].n61 0.114505
R18571 XThC.Tn[11] XThC.Tn[11].n65 0.114505
R18572 XThC.Tn[11].n64 XThC.Tn[11].n63 0.0599512
R18573 XThC.Tn[11].n60 XThC.Tn[11].n59 0.0599512
R18574 XThC.Tn[11].n56 XThC.Tn[11].n55 0.0599512
R18575 XThC.Tn[11].n52 XThC.Tn[11].n51 0.0599512
R18576 XThC.Tn[11].n48 XThC.Tn[11].n47 0.0599512
R18577 XThC.Tn[11].n44 XThC.Tn[11].n43 0.0599512
R18578 XThC.Tn[11].n40 XThC.Tn[11].n39 0.0599512
R18579 XThC.Tn[11].n36 XThC.Tn[11].n35 0.0599512
R18580 XThC.Tn[11].n32 XThC.Tn[11].n31 0.0599512
R18581 XThC.Tn[11].n28 XThC.Tn[11].n27 0.0599512
R18582 XThC.Tn[11].n24 XThC.Tn[11].n23 0.0599512
R18583 XThC.Tn[11].n20 XThC.Tn[11].n19 0.0599512
R18584 XThC.Tn[11].n16 XThC.Tn[11].n15 0.0599512
R18585 XThC.Tn[11].n12 XThC.Tn[11].n11 0.0599512
R18586 XThC.Tn[11].n8 XThC.Tn[11].n7 0.0599512
R18587 XThC.Tn[11].n5 XThC.Tn[11].n4 0.0599512
R18588 XThC.Tn[11].n63 XThC.Tn[11] 0.0469286
R18589 XThC.Tn[11].n59 XThC.Tn[11] 0.0469286
R18590 XThC.Tn[11].n55 XThC.Tn[11] 0.0469286
R18591 XThC.Tn[11].n51 XThC.Tn[11] 0.0469286
R18592 XThC.Tn[11].n47 XThC.Tn[11] 0.0469286
R18593 XThC.Tn[11].n43 XThC.Tn[11] 0.0469286
R18594 XThC.Tn[11].n39 XThC.Tn[11] 0.0469286
R18595 XThC.Tn[11].n35 XThC.Tn[11] 0.0469286
R18596 XThC.Tn[11].n31 XThC.Tn[11] 0.0469286
R18597 XThC.Tn[11].n27 XThC.Tn[11] 0.0469286
R18598 XThC.Tn[11].n23 XThC.Tn[11] 0.0469286
R18599 XThC.Tn[11].n19 XThC.Tn[11] 0.0469286
R18600 XThC.Tn[11].n15 XThC.Tn[11] 0.0469286
R18601 XThC.Tn[11].n11 XThC.Tn[11] 0.0469286
R18602 XThC.Tn[11].n7 XThC.Tn[11] 0.0469286
R18603 XThC.Tn[11].n4 XThC.Tn[11] 0.0469286
R18604 XThC.Tn[11].n63 XThC.Tn[11] 0.0401341
R18605 XThC.Tn[11].n59 XThC.Tn[11] 0.0401341
R18606 XThC.Tn[11].n55 XThC.Tn[11] 0.0401341
R18607 XThC.Tn[11].n51 XThC.Tn[11] 0.0401341
R18608 XThC.Tn[11].n47 XThC.Tn[11] 0.0401341
R18609 XThC.Tn[11].n43 XThC.Tn[11] 0.0401341
R18610 XThC.Tn[11].n39 XThC.Tn[11] 0.0401341
R18611 XThC.Tn[11].n35 XThC.Tn[11] 0.0401341
R18612 XThC.Tn[11].n31 XThC.Tn[11] 0.0401341
R18613 XThC.Tn[11].n27 XThC.Tn[11] 0.0401341
R18614 XThC.Tn[11].n23 XThC.Tn[11] 0.0401341
R18615 XThC.Tn[11].n19 XThC.Tn[11] 0.0401341
R18616 XThC.Tn[11].n15 XThC.Tn[11] 0.0401341
R18617 XThC.Tn[11].n11 XThC.Tn[11] 0.0401341
R18618 XThC.Tn[11].n7 XThC.Tn[11] 0.0401341
R18619 XThC.Tn[11].n4 XThC.Tn[11] 0.0401341
R18620 XThC.Tn[12].n70 XThC.Tn[12].n69 256.104
R18621 XThC.Tn[12].n74 XThC.Tn[12].n72 243.68
R18622 XThC.Tn[12].n2 XThC.Tn[12].n0 241.847
R18623 XThC.Tn[12].n74 XThC.Tn[12].n73 205.28
R18624 XThC.Tn[12].n70 XThC.Tn[12].n68 202.095
R18625 XThC.Tn[12].n2 XThC.Tn[12].n1 185
R18626 XThC.Tn[12].n64 XThC.Tn[12].n62 161.365
R18627 XThC.Tn[12].n60 XThC.Tn[12].n58 161.365
R18628 XThC.Tn[12].n56 XThC.Tn[12].n54 161.365
R18629 XThC.Tn[12].n52 XThC.Tn[12].n50 161.365
R18630 XThC.Tn[12].n48 XThC.Tn[12].n46 161.365
R18631 XThC.Tn[12].n44 XThC.Tn[12].n42 161.365
R18632 XThC.Tn[12].n40 XThC.Tn[12].n38 161.365
R18633 XThC.Tn[12].n36 XThC.Tn[12].n34 161.365
R18634 XThC.Tn[12].n32 XThC.Tn[12].n30 161.365
R18635 XThC.Tn[12].n28 XThC.Tn[12].n26 161.365
R18636 XThC.Tn[12].n24 XThC.Tn[12].n22 161.365
R18637 XThC.Tn[12].n20 XThC.Tn[12].n18 161.365
R18638 XThC.Tn[12].n16 XThC.Tn[12].n14 161.365
R18639 XThC.Tn[12].n12 XThC.Tn[12].n10 161.365
R18640 XThC.Tn[12].n8 XThC.Tn[12].n6 161.365
R18641 XThC.Tn[12].n5 XThC.Tn[12].n3 161.365
R18642 XThC.Tn[12].n62 XThC.Tn[12].t41 161.202
R18643 XThC.Tn[12].n58 XThC.Tn[12].t31 161.202
R18644 XThC.Tn[12].n54 XThC.Tn[12].t18 161.202
R18645 XThC.Tn[12].n50 XThC.Tn[12].t15 161.202
R18646 XThC.Tn[12].n46 XThC.Tn[12].t39 161.202
R18647 XThC.Tn[12].n42 XThC.Tn[12].t26 161.202
R18648 XThC.Tn[12].n38 XThC.Tn[12].t25 161.202
R18649 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R18650 XThC.Tn[12].n30 XThC.Tn[12].t36 161.202
R18651 XThC.Tn[12].n26 XThC.Tn[12].t27 161.202
R18652 XThC.Tn[12].n22 XThC.Tn[12].t14 161.202
R18653 XThC.Tn[12].n18 XThC.Tn[12].t13 161.202
R18654 XThC.Tn[12].n14 XThC.Tn[12].t24 161.202
R18655 XThC.Tn[12].n10 XThC.Tn[12].t22 161.202
R18656 XThC.Tn[12].n6 XThC.Tn[12].t20 161.202
R18657 XThC.Tn[12].n3 XThC.Tn[12].t35 161.202
R18658 XThC.Tn[12].n62 XThC.Tn[12].t12 145.137
R18659 XThC.Tn[12].n58 XThC.Tn[12].t34 145.137
R18660 XThC.Tn[12].n54 XThC.Tn[12].t21 145.137
R18661 XThC.Tn[12].n50 XThC.Tn[12].t19 145.137
R18662 XThC.Tn[12].n46 XThC.Tn[12].t43 145.137
R18663 XThC.Tn[12].n42 XThC.Tn[12].t32 145.137
R18664 XThC.Tn[12].n38 XThC.Tn[12].t30 145.137
R18665 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R18666 XThC.Tn[12].n30 XThC.Tn[12].t40 145.137
R18667 XThC.Tn[12].n26 XThC.Tn[12].t33 145.137
R18668 XThC.Tn[12].n22 XThC.Tn[12].t17 145.137
R18669 XThC.Tn[12].n18 XThC.Tn[12].t16 145.137
R18670 XThC.Tn[12].n14 XThC.Tn[12].t29 145.137
R18671 XThC.Tn[12].n10 XThC.Tn[12].t28 145.137
R18672 XThC.Tn[12].n6 XThC.Tn[12].t23 145.137
R18673 XThC.Tn[12].n3 XThC.Tn[12].t37 145.137
R18674 XThC.Tn[12].n72 XThC.Tn[12].t1 26.5955
R18675 XThC.Tn[12].n72 XThC.Tn[12].t0 26.5955
R18676 XThC.Tn[12].n68 XThC.Tn[12].t5 26.5955
R18677 XThC.Tn[12].n68 XThC.Tn[12].t6 26.5955
R18678 XThC.Tn[12].n69 XThC.Tn[12].t4 26.5955
R18679 XThC.Tn[12].n69 XThC.Tn[12].t7 26.5955
R18680 XThC.Tn[12].n73 XThC.Tn[12].t3 26.5955
R18681 XThC.Tn[12].n73 XThC.Tn[12].t2 26.5955
R18682 XThC.Tn[12].n1 XThC.Tn[12].t9 24.9236
R18683 XThC.Tn[12].n1 XThC.Tn[12].t8 24.9236
R18684 XThC.Tn[12].n0 XThC.Tn[12].t11 24.9236
R18685 XThC.Tn[12].n0 XThC.Tn[12].t10 24.9236
R18686 XThC.Tn[12] XThC.Tn[12].n74 22.9652
R18687 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R18688 XThC.Tn[12].n71 XThC.Tn[12].n70 13.9299
R18689 XThC.Tn[12] XThC.Tn[12].n71 13.9299
R18690 XThC.Tn[12] XThC.Tn[12].n5 8.0245
R18691 XThC.Tn[12].n65 XThC.Tn[12].n64 7.9105
R18692 XThC.Tn[12].n61 XThC.Tn[12].n60 7.9105
R18693 XThC.Tn[12].n57 XThC.Tn[12].n56 7.9105
R18694 XThC.Tn[12].n53 XThC.Tn[12].n52 7.9105
R18695 XThC.Tn[12].n49 XThC.Tn[12].n48 7.9105
R18696 XThC.Tn[12].n45 XThC.Tn[12].n44 7.9105
R18697 XThC.Tn[12].n41 XThC.Tn[12].n40 7.9105
R18698 XThC.Tn[12].n37 XThC.Tn[12].n36 7.9105
R18699 XThC.Tn[12].n33 XThC.Tn[12].n32 7.9105
R18700 XThC.Tn[12].n29 XThC.Tn[12].n28 7.9105
R18701 XThC.Tn[12].n25 XThC.Tn[12].n24 7.9105
R18702 XThC.Tn[12].n21 XThC.Tn[12].n20 7.9105
R18703 XThC.Tn[12].n17 XThC.Tn[12].n16 7.9105
R18704 XThC.Tn[12].n13 XThC.Tn[12].n12 7.9105
R18705 XThC.Tn[12].n9 XThC.Tn[12].n8 7.9105
R18706 XThC.Tn[12].n67 XThC.Tn[12].n66 7.4309
R18707 XThC.Tn[12].n66 XThC.Tn[12] 4.71945
R18708 XThC.Tn[12].n71 XThC.Tn[12].n67 2.99115
R18709 XThC.Tn[12].n71 XThC.Tn[12] 2.87153
R18710 XThC.Tn[12].n67 XThC.Tn[12] 2.2734
R18711 XThC.Tn[12].n66 XThC.Tn[12] 0.88175
R18712 XThC.Tn[12].n9 XThC.Tn[12] 0.235138
R18713 XThC.Tn[12].n13 XThC.Tn[12] 0.235138
R18714 XThC.Tn[12].n17 XThC.Tn[12] 0.235138
R18715 XThC.Tn[12].n21 XThC.Tn[12] 0.235138
R18716 XThC.Tn[12].n25 XThC.Tn[12] 0.235138
R18717 XThC.Tn[12].n29 XThC.Tn[12] 0.235138
R18718 XThC.Tn[12].n33 XThC.Tn[12] 0.235138
R18719 XThC.Tn[12].n37 XThC.Tn[12] 0.235138
R18720 XThC.Tn[12].n41 XThC.Tn[12] 0.235138
R18721 XThC.Tn[12].n45 XThC.Tn[12] 0.235138
R18722 XThC.Tn[12].n49 XThC.Tn[12] 0.235138
R18723 XThC.Tn[12].n53 XThC.Tn[12] 0.235138
R18724 XThC.Tn[12].n57 XThC.Tn[12] 0.235138
R18725 XThC.Tn[12].n61 XThC.Tn[12] 0.235138
R18726 XThC.Tn[12].n65 XThC.Tn[12] 0.235138
R18727 XThC.Tn[12] XThC.Tn[12].n9 0.114505
R18728 XThC.Tn[12] XThC.Tn[12].n13 0.114505
R18729 XThC.Tn[12] XThC.Tn[12].n17 0.114505
R18730 XThC.Tn[12] XThC.Tn[12].n21 0.114505
R18731 XThC.Tn[12] XThC.Tn[12].n25 0.114505
R18732 XThC.Tn[12] XThC.Tn[12].n29 0.114505
R18733 XThC.Tn[12] XThC.Tn[12].n33 0.114505
R18734 XThC.Tn[12] XThC.Tn[12].n37 0.114505
R18735 XThC.Tn[12] XThC.Tn[12].n41 0.114505
R18736 XThC.Tn[12] XThC.Tn[12].n45 0.114505
R18737 XThC.Tn[12] XThC.Tn[12].n49 0.114505
R18738 XThC.Tn[12] XThC.Tn[12].n53 0.114505
R18739 XThC.Tn[12] XThC.Tn[12].n57 0.114505
R18740 XThC.Tn[12] XThC.Tn[12].n61 0.114505
R18741 XThC.Tn[12] XThC.Tn[12].n65 0.114505
R18742 XThC.Tn[12].n64 XThC.Tn[12].n63 0.0599512
R18743 XThC.Tn[12].n60 XThC.Tn[12].n59 0.0599512
R18744 XThC.Tn[12].n56 XThC.Tn[12].n55 0.0599512
R18745 XThC.Tn[12].n52 XThC.Tn[12].n51 0.0599512
R18746 XThC.Tn[12].n48 XThC.Tn[12].n47 0.0599512
R18747 XThC.Tn[12].n44 XThC.Tn[12].n43 0.0599512
R18748 XThC.Tn[12].n40 XThC.Tn[12].n39 0.0599512
R18749 XThC.Tn[12].n36 XThC.Tn[12].n35 0.0599512
R18750 XThC.Tn[12].n32 XThC.Tn[12].n31 0.0599512
R18751 XThC.Tn[12].n28 XThC.Tn[12].n27 0.0599512
R18752 XThC.Tn[12].n24 XThC.Tn[12].n23 0.0599512
R18753 XThC.Tn[12].n20 XThC.Tn[12].n19 0.0599512
R18754 XThC.Tn[12].n16 XThC.Tn[12].n15 0.0599512
R18755 XThC.Tn[12].n12 XThC.Tn[12].n11 0.0599512
R18756 XThC.Tn[12].n8 XThC.Tn[12].n7 0.0599512
R18757 XThC.Tn[12].n5 XThC.Tn[12].n4 0.0599512
R18758 XThC.Tn[12].n63 XThC.Tn[12] 0.0469286
R18759 XThC.Tn[12].n59 XThC.Tn[12] 0.0469286
R18760 XThC.Tn[12].n55 XThC.Tn[12] 0.0469286
R18761 XThC.Tn[12].n51 XThC.Tn[12] 0.0469286
R18762 XThC.Tn[12].n47 XThC.Tn[12] 0.0469286
R18763 XThC.Tn[12].n43 XThC.Tn[12] 0.0469286
R18764 XThC.Tn[12].n39 XThC.Tn[12] 0.0469286
R18765 XThC.Tn[12].n35 XThC.Tn[12] 0.0469286
R18766 XThC.Tn[12].n31 XThC.Tn[12] 0.0469286
R18767 XThC.Tn[12].n27 XThC.Tn[12] 0.0469286
R18768 XThC.Tn[12].n23 XThC.Tn[12] 0.0469286
R18769 XThC.Tn[12].n19 XThC.Tn[12] 0.0469286
R18770 XThC.Tn[12].n15 XThC.Tn[12] 0.0469286
R18771 XThC.Tn[12].n11 XThC.Tn[12] 0.0469286
R18772 XThC.Tn[12].n7 XThC.Tn[12] 0.0469286
R18773 XThC.Tn[12].n4 XThC.Tn[12] 0.0469286
R18774 XThC.Tn[12].n63 XThC.Tn[12] 0.0401341
R18775 XThC.Tn[12].n59 XThC.Tn[12] 0.0401341
R18776 XThC.Tn[12].n55 XThC.Tn[12] 0.0401341
R18777 XThC.Tn[12].n51 XThC.Tn[12] 0.0401341
R18778 XThC.Tn[12].n47 XThC.Tn[12] 0.0401341
R18779 XThC.Tn[12].n43 XThC.Tn[12] 0.0401341
R18780 XThC.Tn[12].n39 XThC.Tn[12] 0.0401341
R18781 XThC.Tn[12].n35 XThC.Tn[12] 0.0401341
R18782 XThC.Tn[12].n31 XThC.Tn[12] 0.0401341
R18783 XThC.Tn[12].n27 XThC.Tn[12] 0.0401341
R18784 XThC.Tn[12].n23 XThC.Tn[12] 0.0401341
R18785 XThC.Tn[12].n19 XThC.Tn[12] 0.0401341
R18786 XThC.Tn[12].n15 XThC.Tn[12] 0.0401341
R18787 XThC.Tn[12].n11 XThC.Tn[12] 0.0401341
R18788 XThC.Tn[12].n7 XThC.Tn[12] 0.0401341
R18789 XThC.Tn[12].n4 XThC.Tn[12] 0.0401341
R18790 XThC.Tn[13].n70 XThC.Tn[13].n69 265.341
R18791 XThC.Tn[13].n74 XThC.Tn[13].n72 243.68
R18792 XThC.Tn[13].n2 XThC.Tn[13].n0 241.847
R18793 XThC.Tn[13].n74 XThC.Tn[13].n73 205.28
R18794 XThC.Tn[13].n70 XThC.Tn[13].n68 202.094
R18795 XThC.Tn[13].n2 XThC.Tn[13].n1 185
R18796 XThC.Tn[13].n64 XThC.Tn[13].n62 161.365
R18797 XThC.Tn[13].n60 XThC.Tn[13].n58 161.365
R18798 XThC.Tn[13].n56 XThC.Tn[13].n54 161.365
R18799 XThC.Tn[13].n52 XThC.Tn[13].n50 161.365
R18800 XThC.Tn[13].n48 XThC.Tn[13].n46 161.365
R18801 XThC.Tn[13].n44 XThC.Tn[13].n42 161.365
R18802 XThC.Tn[13].n40 XThC.Tn[13].n38 161.365
R18803 XThC.Tn[13].n36 XThC.Tn[13].n34 161.365
R18804 XThC.Tn[13].n32 XThC.Tn[13].n30 161.365
R18805 XThC.Tn[13].n28 XThC.Tn[13].n26 161.365
R18806 XThC.Tn[13].n24 XThC.Tn[13].n22 161.365
R18807 XThC.Tn[13].n20 XThC.Tn[13].n18 161.365
R18808 XThC.Tn[13].n16 XThC.Tn[13].n14 161.365
R18809 XThC.Tn[13].n12 XThC.Tn[13].n10 161.365
R18810 XThC.Tn[13].n8 XThC.Tn[13].n6 161.365
R18811 XThC.Tn[13].n5 XThC.Tn[13].n3 161.365
R18812 XThC.Tn[13].n62 XThC.Tn[13].t33 161.202
R18813 XThC.Tn[13].n58 XThC.Tn[13].t23 161.202
R18814 XThC.Tn[13].n54 XThC.Tn[13].t42 161.202
R18815 XThC.Tn[13].n50 XThC.Tn[13].t39 161.202
R18816 XThC.Tn[13].n46 XThC.Tn[13].t31 161.202
R18817 XThC.Tn[13].n42 XThC.Tn[13].t18 161.202
R18818 XThC.Tn[13].n38 XThC.Tn[13].t17 161.202
R18819 XThC.Tn[13].n34 XThC.Tn[13].t30 161.202
R18820 XThC.Tn[13].n30 XThC.Tn[13].t28 161.202
R18821 XThC.Tn[13].n26 XThC.Tn[13].t19 161.202
R18822 XThC.Tn[13].n22 XThC.Tn[13].t38 161.202
R18823 XThC.Tn[13].n18 XThC.Tn[13].t37 161.202
R18824 XThC.Tn[13].n14 XThC.Tn[13].t16 161.202
R18825 XThC.Tn[13].n10 XThC.Tn[13].t14 161.202
R18826 XThC.Tn[13].n6 XThC.Tn[13].t12 161.202
R18827 XThC.Tn[13].n3 XThC.Tn[13].t27 161.202
R18828 XThC.Tn[13].n62 XThC.Tn[13].t36 145.137
R18829 XThC.Tn[13].n58 XThC.Tn[13].t26 145.137
R18830 XThC.Tn[13].n54 XThC.Tn[13].t13 145.137
R18831 XThC.Tn[13].n50 XThC.Tn[13].t43 145.137
R18832 XThC.Tn[13].n46 XThC.Tn[13].t35 145.137
R18833 XThC.Tn[13].n42 XThC.Tn[13].t24 145.137
R18834 XThC.Tn[13].n38 XThC.Tn[13].t22 145.137
R18835 XThC.Tn[13].n34 XThC.Tn[13].t34 145.137
R18836 XThC.Tn[13].n30 XThC.Tn[13].t32 145.137
R18837 XThC.Tn[13].n26 XThC.Tn[13].t25 145.137
R18838 XThC.Tn[13].n22 XThC.Tn[13].t41 145.137
R18839 XThC.Tn[13].n18 XThC.Tn[13].t40 145.137
R18840 XThC.Tn[13].n14 XThC.Tn[13].t21 145.137
R18841 XThC.Tn[13].n10 XThC.Tn[13].t20 145.137
R18842 XThC.Tn[13].n6 XThC.Tn[13].t15 145.137
R18843 XThC.Tn[13].n3 XThC.Tn[13].t29 145.137
R18844 XThC.Tn[13].n72 XThC.Tn[13].t1 26.5955
R18845 XThC.Tn[13].n72 XThC.Tn[13].t0 26.5955
R18846 XThC.Tn[13].n69 XThC.Tn[13].t4 26.5955
R18847 XThC.Tn[13].n69 XThC.Tn[13].t7 26.5955
R18848 XThC.Tn[13].n68 XThC.Tn[13].t6 26.5955
R18849 XThC.Tn[13].n68 XThC.Tn[13].t5 26.5955
R18850 XThC.Tn[13].n73 XThC.Tn[13].t3 26.5955
R18851 XThC.Tn[13].n73 XThC.Tn[13].t2 26.5955
R18852 XThC.Tn[13].n1 XThC.Tn[13].t8 24.9236
R18853 XThC.Tn[13].n1 XThC.Tn[13].t10 24.9236
R18854 XThC.Tn[13].n0 XThC.Tn[13].t11 24.9236
R18855 XThC.Tn[13].n0 XThC.Tn[13].t9 24.9236
R18856 XThC.Tn[13] XThC.Tn[13].n74 22.9652
R18857 XThC.Tn[13] XThC.Tn[13].n2 18.8943
R18858 XThC.Tn[13].n71 XThC.Tn[13].n70 13.9299
R18859 XThC.Tn[13] XThC.Tn[13].n71 13.9299
R18860 XThC.Tn[13] XThC.Tn[13].n5 8.0245
R18861 XThC.Tn[13].n65 XThC.Tn[13].n64 7.9105
R18862 XThC.Tn[13].n61 XThC.Tn[13].n60 7.9105
R18863 XThC.Tn[13].n57 XThC.Tn[13].n56 7.9105
R18864 XThC.Tn[13].n53 XThC.Tn[13].n52 7.9105
R18865 XThC.Tn[13].n49 XThC.Tn[13].n48 7.9105
R18866 XThC.Tn[13].n45 XThC.Tn[13].n44 7.9105
R18867 XThC.Tn[13].n41 XThC.Tn[13].n40 7.9105
R18868 XThC.Tn[13].n37 XThC.Tn[13].n36 7.9105
R18869 XThC.Tn[13].n33 XThC.Tn[13].n32 7.9105
R18870 XThC.Tn[13].n29 XThC.Tn[13].n28 7.9105
R18871 XThC.Tn[13].n25 XThC.Tn[13].n24 7.9105
R18872 XThC.Tn[13].n21 XThC.Tn[13].n20 7.9105
R18873 XThC.Tn[13].n17 XThC.Tn[13].n16 7.9105
R18874 XThC.Tn[13].n13 XThC.Tn[13].n12 7.9105
R18875 XThC.Tn[13].n9 XThC.Tn[13].n8 7.9105
R18876 XThC.Tn[13].n67 XThC.Tn[13].n66 7.46054
R18877 XThC.Tn[13].n67 XThC.Tn[13] 6.34069
R18878 XThC.Tn[13].n66 XThC.Tn[13] 4.78838
R18879 XThC.Tn[13] XThC.Tn[13].n67 1.79489
R18880 XThC.Tn[13].n66 XThC.Tn[13] 1.51436
R18881 XThC.Tn[13].n71 XThC.Tn[13] 1.19676
R18882 XThC.Tn[13].n9 XThC.Tn[13] 0.235138
R18883 XThC.Tn[13].n13 XThC.Tn[13] 0.235138
R18884 XThC.Tn[13].n17 XThC.Tn[13] 0.235138
R18885 XThC.Tn[13].n21 XThC.Tn[13] 0.235138
R18886 XThC.Tn[13].n25 XThC.Tn[13] 0.235138
R18887 XThC.Tn[13].n29 XThC.Tn[13] 0.235138
R18888 XThC.Tn[13].n33 XThC.Tn[13] 0.235138
R18889 XThC.Tn[13].n37 XThC.Tn[13] 0.235138
R18890 XThC.Tn[13].n41 XThC.Tn[13] 0.235138
R18891 XThC.Tn[13].n45 XThC.Tn[13] 0.235138
R18892 XThC.Tn[13].n49 XThC.Tn[13] 0.235138
R18893 XThC.Tn[13].n53 XThC.Tn[13] 0.235138
R18894 XThC.Tn[13].n57 XThC.Tn[13] 0.235138
R18895 XThC.Tn[13].n61 XThC.Tn[13] 0.235138
R18896 XThC.Tn[13].n65 XThC.Tn[13] 0.235138
R18897 XThC.Tn[13] XThC.Tn[13].n9 0.114505
R18898 XThC.Tn[13] XThC.Tn[13].n13 0.114505
R18899 XThC.Tn[13] XThC.Tn[13].n17 0.114505
R18900 XThC.Tn[13] XThC.Tn[13].n21 0.114505
R18901 XThC.Tn[13] XThC.Tn[13].n25 0.114505
R18902 XThC.Tn[13] XThC.Tn[13].n29 0.114505
R18903 XThC.Tn[13] XThC.Tn[13].n33 0.114505
R18904 XThC.Tn[13] XThC.Tn[13].n37 0.114505
R18905 XThC.Tn[13] XThC.Tn[13].n41 0.114505
R18906 XThC.Tn[13] XThC.Tn[13].n45 0.114505
R18907 XThC.Tn[13] XThC.Tn[13].n49 0.114505
R18908 XThC.Tn[13] XThC.Tn[13].n53 0.114505
R18909 XThC.Tn[13] XThC.Tn[13].n57 0.114505
R18910 XThC.Tn[13] XThC.Tn[13].n61 0.114505
R18911 XThC.Tn[13] XThC.Tn[13].n65 0.114505
R18912 XThC.Tn[13].n64 XThC.Tn[13].n63 0.0599512
R18913 XThC.Tn[13].n60 XThC.Tn[13].n59 0.0599512
R18914 XThC.Tn[13].n56 XThC.Tn[13].n55 0.0599512
R18915 XThC.Tn[13].n52 XThC.Tn[13].n51 0.0599512
R18916 XThC.Tn[13].n48 XThC.Tn[13].n47 0.0599512
R18917 XThC.Tn[13].n44 XThC.Tn[13].n43 0.0599512
R18918 XThC.Tn[13].n40 XThC.Tn[13].n39 0.0599512
R18919 XThC.Tn[13].n36 XThC.Tn[13].n35 0.0599512
R18920 XThC.Tn[13].n32 XThC.Tn[13].n31 0.0599512
R18921 XThC.Tn[13].n28 XThC.Tn[13].n27 0.0599512
R18922 XThC.Tn[13].n24 XThC.Tn[13].n23 0.0599512
R18923 XThC.Tn[13].n20 XThC.Tn[13].n19 0.0599512
R18924 XThC.Tn[13].n16 XThC.Tn[13].n15 0.0599512
R18925 XThC.Tn[13].n12 XThC.Tn[13].n11 0.0599512
R18926 XThC.Tn[13].n8 XThC.Tn[13].n7 0.0599512
R18927 XThC.Tn[13].n5 XThC.Tn[13].n4 0.0599512
R18928 XThC.Tn[13].n63 XThC.Tn[13] 0.0469286
R18929 XThC.Tn[13].n59 XThC.Tn[13] 0.0469286
R18930 XThC.Tn[13].n55 XThC.Tn[13] 0.0469286
R18931 XThC.Tn[13].n51 XThC.Tn[13] 0.0469286
R18932 XThC.Tn[13].n47 XThC.Tn[13] 0.0469286
R18933 XThC.Tn[13].n43 XThC.Tn[13] 0.0469286
R18934 XThC.Tn[13].n39 XThC.Tn[13] 0.0469286
R18935 XThC.Tn[13].n35 XThC.Tn[13] 0.0469286
R18936 XThC.Tn[13].n31 XThC.Tn[13] 0.0469286
R18937 XThC.Tn[13].n27 XThC.Tn[13] 0.0469286
R18938 XThC.Tn[13].n23 XThC.Tn[13] 0.0469286
R18939 XThC.Tn[13].n19 XThC.Tn[13] 0.0469286
R18940 XThC.Tn[13].n15 XThC.Tn[13] 0.0469286
R18941 XThC.Tn[13].n11 XThC.Tn[13] 0.0469286
R18942 XThC.Tn[13].n7 XThC.Tn[13] 0.0469286
R18943 XThC.Tn[13].n4 XThC.Tn[13] 0.0469286
R18944 XThC.Tn[13].n63 XThC.Tn[13] 0.0401341
R18945 XThC.Tn[13].n59 XThC.Tn[13] 0.0401341
R18946 XThC.Tn[13].n55 XThC.Tn[13] 0.0401341
R18947 XThC.Tn[13].n51 XThC.Tn[13] 0.0401341
R18948 XThC.Tn[13].n47 XThC.Tn[13] 0.0401341
R18949 XThC.Tn[13].n43 XThC.Tn[13] 0.0401341
R18950 XThC.Tn[13].n39 XThC.Tn[13] 0.0401341
R18951 XThC.Tn[13].n35 XThC.Tn[13] 0.0401341
R18952 XThC.Tn[13].n31 XThC.Tn[13] 0.0401341
R18953 XThC.Tn[13].n27 XThC.Tn[13] 0.0401341
R18954 XThC.Tn[13].n23 XThC.Tn[13] 0.0401341
R18955 XThC.Tn[13].n19 XThC.Tn[13] 0.0401341
R18956 XThC.Tn[13].n15 XThC.Tn[13] 0.0401341
R18957 XThC.Tn[13].n11 XThC.Tn[13] 0.0401341
R18958 XThC.Tn[13].n7 XThC.Tn[13] 0.0401341
R18959 XThC.Tn[13].n4 XThC.Tn[13] 0.0401341
R18960 XThC.Tn[0].n74 XThC.Tn[0].n73 332.332
R18961 XThC.Tn[0].n74 XThC.Tn[0].n72 296.493
R18962 XThC.Tn[0].n68 XThC.Tn[0].n66 161.365
R18963 XThC.Tn[0].n64 XThC.Tn[0].n62 161.365
R18964 XThC.Tn[0].n60 XThC.Tn[0].n58 161.365
R18965 XThC.Tn[0].n56 XThC.Tn[0].n54 161.365
R18966 XThC.Tn[0].n52 XThC.Tn[0].n50 161.365
R18967 XThC.Tn[0].n48 XThC.Tn[0].n46 161.365
R18968 XThC.Tn[0].n44 XThC.Tn[0].n42 161.365
R18969 XThC.Tn[0].n40 XThC.Tn[0].n38 161.365
R18970 XThC.Tn[0].n36 XThC.Tn[0].n34 161.365
R18971 XThC.Tn[0].n32 XThC.Tn[0].n30 161.365
R18972 XThC.Tn[0].n28 XThC.Tn[0].n26 161.365
R18973 XThC.Tn[0].n24 XThC.Tn[0].n22 161.365
R18974 XThC.Tn[0].n20 XThC.Tn[0].n18 161.365
R18975 XThC.Tn[0].n16 XThC.Tn[0].n14 161.365
R18976 XThC.Tn[0].n12 XThC.Tn[0].n10 161.365
R18977 XThC.Tn[0].n9 XThC.Tn[0].n7 161.365
R18978 XThC.Tn[0].n66 XThC.Tn[0].t29 161.202
R18979 XThC.Tn[0].n62 XThC.Tn[0].t19 161.202
R18980 XThC.Tn[0].n58 XThC.Tn[0].t38 161.202
R18981 XThC.Tn[0].n54 XThC.Tn[0].t36 161.202
R18982 XThC.Tn[0].n50 XThC.Tn[0].t27 161.202
R18983 XThC.Tn[0].n46 XThC.Tn[0].t16 161.202
R18984 XThC.Tn[0].n42 XThC.Tn[0].t15 161.202
R18985 XThC.Tn[0].n38 XThC.Tn[0].t26 161.202
R18986 XThC.Tn[0].n34 XThC.Tn[0].t25 161.202
R18987 XThC.Tn[0].n30 XThC.Tn[0].t17 161.202
R18988 XThC.Tn[0].n26 XThC.Tn[0].t34 161.202
R18989 XThC.Tn[0].n22 XThC.Tn[0].t32 161.202
R18990 XThC.Tn[0].n18 XThC.Tn[0].t13 161.202
R18991 XThC.Tn[0].n14 XThC.Tn[0].t12 161.202
R18992 XThC.Tn[0].n10 XThC.Tn[0].t41 161.202
R18993 XThC.Tn[0].n7 XThC.Tn[0].t22 161.202
R18994 XThC.Tn[0].n66 XThC.Tn[0].t24 145.137
R18995 XThC.Tn[0].n62 XThC.Tn[0].t14 145.137
R18996 XThC.Tn[0].n58 XThC.Tn[0].t33 145.137
R18997 XThC.Tn[0].n54 XThC.Tn[0].t31 145.137
R18998 XThC.Tn[0].n50 XThC.Tn[0].t23 145.137
R18999 XThC.Tn[0].n46 XThC.Tn[0].t42 145.137
R19000 XThC.Tn[0].n42 XThC.Tn[0].t40 145.137
R19001 XThC.Tn[0].n38 XThC.Tn[0].t21 145.137
R19002 XThC.Tn[0].n34 XThC.Tn[0].t20 145.137
R19003 XThC.Tn[0].n30 XThC.Tn[0].t43 145.137
R19004 XThC.Tn[0].n26 XThC.Tn[0].t30 145.137
R19005 XThC.Tn[0].n22 XThC.Tn[0].t28 145.137
R19006 XThC.Tn[0].n18 XThC.Tn[0].t39 145.137
R19007 XThC.Tn[0].n14 XThC.Tn[0].t37 145.137
R19008 XThC.Tn[0].n10 XThC.Tn[0].t35 145.137
R19009 XThC.Tn[0].n7 XThC.Tn[0].t18 145.137
R19010 XThC.Tn[0].n2 XThC.Tn[0].n0 135.248
R19011 XThC.Tn[0].n2 XThC.Tn[0].n1 98.982
R19012 XThC.Tn[0].n4 XThC.Tn[0].n3 98.982
R19013 XThC.Tn[0].n6 XThC.Tn[0].n5 98.982
R19014 XThC.Tn[0].n4 XThC.Tn[0].n2 36.2672
R19015 XThC.Tn[0].n6 XThC.Tn[0].n4 36.2672
R19016 XThC.Tn[0].n71 XThC.Tn[0].n6 32.6405
R19017 XThC.Tn[0].n72 XThC.Tn[0].t1 26.5955
R19018 XThC.Tn[0].n72 XThC.Tn[0].t0 26.5955
R19019 XThC.Tn[0].n73 XThC.Tn[0].t3 26.5955
R19020 XThC.Tn[0].n73 XThC.Tn[0].t2 26.5955
R19021 XThC.Tn[0].n0 XThC.Tn[0].t11 24.9236
R19022 XThC.Tn[0].n0 XThC.Tn[0].t10 24.9236
R19023 XThC.Tn[0].n1 XThC.Tn[0].t8 24.9236
R19024 XThC.Tn[0].n1 XThC.Tn[0].t9 24.9236
R19025 XThC.Tn[0].n3 XThC.Tn[0].t7 24.9236
R19026 XThC.Tn[0].n3 XThC.Tn[0].t6 24.9236
R19027 XThC.Tn[0].n5 XThC.Tn[0].t5 24.9236
R19028 XThC.Tn[0].n5 XThC.Tn[0].t4 24.9236
R19029 XThC.Tn[0].n75 XThC.Tn[0].n74 18.5605
R19030 XThC.Tn[0].n75 XThC.Tn[0].n71 11.5205
R19031 XThC.Tn[0] XThC.Tn[0].n9 8.0245
R19032 XThC.Tn[0].n69 XThC.Tn[0].n68 7.9105
R19033 XThC.Tn[0].n65 XThC.Tn[0].n64 7.9105
R19034 XThC.Tn[0].n61 XThC.Tn[0].n60 7.9105
R19035 XThC.Tn[0].n57 XThC.Tn[0].n56 7.9105
R19036 XThC.Tn[0].n53 XThC.Tn[0].n52 7.9105
R19037 XThC.Tn[0].n49 XThC.Tn[0].n48 7.9105
R19038 XThC.Tn[0].n45 XThC.Tn[0].n44 7.9105
R19039 XThC.Tn[0].n41 XThC.Tn[0].n40 7.9105
R19040 XThC.Tn[0].n37 XThC.Tn[0].n36 7.9105
R19041 XThC.Tn[0].n33 XThC.Tn[0].n32 7.9105
R19042 XThC.Tn[0].n29 XThC.Tn[0].n28 7.9105
R19043 XThC.Tn[0].n25 XThC.Tn[0].n24 7.9105
R19044 XThC.Tn[0].n21 XThC.Tn[0].n20 7.9105
R19045 XThC.Tn[0].n17 XThC.Tn[0].n16 7.9105
R19046 XThC.Tn[0].n13 XThC.Tn[0].n12 7.9105
R19047 XThC.Tn[0].n70 XThC.Tn[0] 5.90911
R19048 XThC.Tn[0].n71 XThC.Tn[0].n70 4.6005
R19049 XThC.Tn[0].n70 XThC.Tn[0] 1.89022
R19050 XThC.Tn[0] XThC.Tn[0].n75 0.6405
R19051 XThC.Tn[0].n13 XThC.Tn[0] 0.235138
R19052 XThC.Tn[0].n17 XThC.Tn[0] 0.235138
R19053 XThC.Tn[0].n21 XThC.Tn[0] 0.235138
R19054 XThC.Tn[0].n25 XThC.Tn[0] 0.235138
R19055 XThC.Tn[0].n29 XThC.Tn[0] 0.235138
R19056 XThC.Tn[0].n33 XThC.Tn[0] 0.235138
R19057 XThC.Tn[0].n37 XThC.Tn[0] 0.235138
R19058 XThC.Tn[0].n41 XThC.Tn[0] 0.235138
R19059 XThC.Tn[0].n45 XThC.Tn[0] 0.235138
R19060 XThC.Tn[0].n49 XThC.Tn[0] 0.235138
R19061 XThC.Tn[0].n53 XThC.Tn[0] 0.235138
R19062 XThC.Tn[0].n57 XThC.Tn[0] 0.235138
R19063 XThC.Tn[0].n61 XThC.Tn[0] 0.235138
R19064 XThC.Tn[0].n65 XThC.Tn[0] 0.235138
R19065 XThC.Tn[0].n69 XThC.Tn[0] 0.235138
R19066 XThC.Tn[0] XThC.Tn[0].n13 0.114505
R19067 XThC.Tn[0] XThC.Tn[0].n17 0.114505
R19068 XThC.Tn[0] XThC.Tn[0].n21 0.114505
R19069 XThC.Tn[0] XThC.Tn[0].n25 0.114505
R19070 XThC.Tn[0] XThC.Tn[0].n29 0.114505
R19071 XThC.Tn[0] XThC.Tn[0].n33 0.114505
R19072 XThC.Tn[0] XThC.Tn[0].n37 0.114505
R19073 XThC.Tn[0] XThC.Tn[0].n41 0.114505
R19074 XThC.Tn[0] XThC.Tn[0].n45 0.114505
R19075 XThC.Tn[0] XThC.Tn[0].n49 0.114505
R19076 XThC.Tn[0] XThC.Tn[0].n53 0.114505
R19077 XThC.Tn[0] XThC.Tn[0].n57 0.114505
R19078 XThC.Tn[0] XThC.Tn[0].n61 0.114505
R19079 XThC.Tn[0] XThC.Tn[0].n65 0.114505
R19080 XThC.Tn[0] XThC.Tn[0].n69 0.114505
R19081 XThC.Tn[0].n68 XThC.Tn[0].n67 0.0599512
R19082 XThC.Tn[0].n64 XThC.Tn[0].n63 0.0599512
R19083 XThC.Tn[0].n60 XThC.Tn[0].n59 0.0599512
R19084 XThC.Tn[0].n56 XThC.Tn[0].n55 0.0599512
R19085 XThC.Tn[0].n52 XThC.Tn[0].n51 0.0599512
R19086 XThC.Tn[0].n48 XThC.Tn[0].n47 0.0599512
R19087 XThC.Tn[0].n44 XThC.Tn[0].n43 0.0599512
R19088 XThC.Tn[0].n40 XThC.Tn[0].n39 0.0599512
R19089 XThC.Tn[0].n36 XThC.Tn[0].n35 0.0599512
R19090 XThC.Tn[0].n32 XThC.Tn[0].n31 0.0599512
R19091 XThC.Tn[0].n28 XThC.Tn[0].n27 0.0599512
R19092 XThC.Tn[0].n24 XThC.Tn[0].n23 0.0599512
R19093 XThC.Tn[0].n20 XThC.Tn[0].n19 0.0599512
R19094 XThC.Tn[0].n16 XThC.Tn[0].n15 0.0599512
R19095 XThC.Tn[0].n12 XThC.Tn[0].n11 0.0599512
R19096 XThC.Tn[0].n9 XThC.Tn[0].n8 0.0599512
R19097 XThC.Tn[0].n67 XThC.Tn[0] 0.0469286
R19098 XThC.Tn[0].n63 XThC.Tn[0] 0.0469286
R19099 XThC.Tn[0].n59 XThC.Tn[0] 0.0469286
R19100 XThC.Tn[0].n55 XThC.Tn[0] 0.0469286
R19101 XThC.Tn[0].n51 XThC.Tn[0] 0.0469286
R19102 XThC.Tn[0].n47 XThC.Tn[0] 0.0469286
R19103 XThC.Tn[0].n43 XThC.Tn[0] 0.0469286
R19104 XThC.Tn[0].n39 XThC.Tn[0] 0.0469286
R19105 XThC.Tn[0].n35 XThC.Tn[0] 0.0469286
R19106 XThC.Tn[0].n31 XThC.Tn[0] 0.0469286
R19107 XThC.Tn[0].n27 XThC.Tn[0] 0.0469286
R19108 XThC.Tn[0].n23 XThC.Tn[0] 0.0469286
R19109 XThC.Tn[0].n19 XThC.Tn[0] 0.0469286
R19110 XThC.Tn[0].n15 XThC.Tn[0] 0.0469286
R19111 XThC.Tn[0].n11 XThC.Tn[0] 0.0469286
R19112 XThC.Tn[0].n8 XThC.Tn[0] 0.0469286
R19113 XThC.Tn[0].n67 XThC.Tn[0] 0.0401341
R19114 XThC.Tn[0].n63 XThC.Tn[0] 0.0401341
R19115 XThC.Tn[0].n59 XThC.Tn[0] 0.0401341
R19116 XThC.Tn[0].n55 XThC.Tn[0] 0.0401341
R19117 XThC.Tn[0].n51 XThC.Tn[0] 0.0401341
R19118 XThC.Tn[0].n47 XThC.Tn[0] 0.0401341
R19119 XThC.Tn[0].n43 XThC.Tn[0] 0.0401341
R19120 XThC.Tn[0].n39 XThC.Tn[0] 0.0401341
R19121 XThC.Tn[0].n35 XThC.Tn[0] 0.0401341
R19122 XThC.Tn[0].n31 XThC.Tn[0] 0.0401341
R19123 XThC.Tn[0].n27 XThC.Tn[0] 0.0401341
R19124 XThC.Tn[0].n23 XThC.Tn[0] 0.0401341
R19125 XThC.Tn[0].n19 XThC.Tn[0] 0.0401341
R19126 XThC.Tn[0].n15 XThC.Tn[0] 0.0401341
R19127 XThC.Tn[0].n11 XThC.Tn[0] 0.0401341
R19128 XThC.Tn[0].n8 XThC.Tn[0] 0.0401341
R19129 XThC.XTB4.Y.n21 XThC.XTB4.Y.t0 235.56
R19130 XThC.XTB4.Y.n3 XThC.XTB4.Y.t3 212.081
R19131 XThC.XTB4.Y.n2 XThC.XTB4.Y.t2 212.081
R19132 XThC.XTB4.Y.n8 XThC.XTB4.Y.t17 212.081
R19133 XThC.XTB4.Y.n0 XThC.XTB4.Y.t13 212.081
R19134 XThC.XTB4.Y.n12 XThC.XTB4.Y.t8 212.081
R19135 XThC.XTB4.Y.n13 XThC.XTB4.Y.t12 212.081
R19136 XThC.XTB4.Y.n15 XThC.XTB4.Y.t6 212.081
R19137 XThC.XTB4.Y.n11 XThC.XTB4.Y.t16 212.081
R19138 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 173.761
R19139 XThC.XTB4.Y.n14 XThC.XTB4.Y 158.656
R19140 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 152
R19141 XThC.XTB4.Y.n5 XThC.XTB4.Y.n1 152
R19142 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 152
R19143 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 152
R19144 XThC.XTB4.Y.n3 XThC.XTB4.Y.t14 139.78
R19145 XThC.XTB4.Y.n2 XThC.XTB4.Y.t10 139.78
R19146 XThC.XTB4.Y.n8 XThC.XTB4.Y.t7 139.78
R19147 XThC.XTB4.Y.n0 XThC.XTB4.Y.t4 139.78
R19148 XThC.XTB4.Y.n12 XThC.XTB4.Y.t11 139.78
R19149 XThC.XTB4.Y.n13 XThC.XTB4.Y.t15 139.78
R19150 XThC.XTB4.Y.n15 XThC.XTB4.Y.t9 139.78
R19151 XThC.XTB4.Y.n11 XThC.XTB4.Y.t5 139.78
R19152 XThC.XTB4.Y.n20 XThC.XTB4.Y.t1 133.386
R19153 XThC.XTB4.Y.n19 XThC.XTB4.Y.n10 72.9296
R19154 XThC.XTB4.Y.n13 XThC.XTB4.Y.n12 61.346
R19155 XThC.XTB4.Y.n7 XThC.XTB4.Y.n1 49.6611
R19156 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 45.2793
R19157 XThC.XTB4.Y.n4 XThC.XTB4.Y.n2 42.3581
R19158 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 38.1854
R19159 XThC.XTB4.Y.n16 XThC.XTB4.Y.n11 30.6732
R19160 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R19161 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R19162 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 30.6732
R19163 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 21.7605
R19164 XThC.XTB4.Y XThC.XTB4.Y.n20 19.5051
R19165 XThC.XTB4.Y.n4 XThC.XTB4.Y.n3 18.9884
R19166 XThC.XTB4.Y.n9 XThC.XTB4.Y.n0 16.0672
R19167 XThC.XTB4.Y.n17 XThC.XTB4.Y 14.7905
R19168 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 11.994
R19169 XThC.XTB4.Y.n10 XThC.XTB4.Y 11.5205
R19170 XThC.XTB4.Y.n6 XThC.XTB4.Y 10.2405
R19171 XThC.XTB4.Y.n2 XThC.XTB4.Y.n1 7.30353
R19172 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 7.24578
R19173 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 4.38232
R19174 XThC.XTB4.Y.n21 XThC.XTB4.Y 2.22659
R19175 XThC.XTB4.Y XThC.XTB4.Y.n21 1.55202
R19176 XThC.XTB4.Y.n18 XThC.XTB4.Y 0.966538
R19177 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19178 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19179 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19180 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19181 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19182 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19183 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19184 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19185 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19186 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19187 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19188 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19189 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19190 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19191 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19192 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19193 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19194 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19195 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19196 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19197 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19198 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19199 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19200 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19201 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19202 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19203 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19204 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19205 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19206 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19207 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19208 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19209 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19210 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19211 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19212 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19213 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19214 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19215 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19216 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19217 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19218 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19219 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19220 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19221 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19222 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19223 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19224 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19225 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19226 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19227 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19228 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19229 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19230 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19231 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19232 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19233 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19234 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19235 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19236 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19237 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19238 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19239 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19240 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19241 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19242 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19243 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19244 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19245 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19246 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19247 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19248 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19249 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19250 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19251 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19252 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19253 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19254 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19255 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19256 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19257 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19258 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19259 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19260 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19261 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19262 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19263 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19264 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19265 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19266 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19267 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19268 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19269 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19270 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19271 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19272 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R19273 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19274 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19275 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R19276 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19277 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19278 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19279 XThR.Tn[3].n1 XThR.Tn[3].t3 26.5955
R19280 XThR.Tn[3].n1 XThR.Tn[3].t6 26.5955
R19281 XThR.Tn[3].n0 XThR.Tn[3].t4 26.5955
R19282 XThR.Tn[3].n0 XThR.Tn[3].t5 26.5955
R19283 XThR.Tn[3].n3 XThR.Tn[3].t10 24.9236
R19284 XThR.Tn[3].n3 XThR.Tn[3].t7 24.9236
R19285 XThR.Tn[3].n4 XThR.Tn[3].t9 24.9236
R19286 XThR.Tn[3].n4 XThR.Tn[3].t8 24.9236
R19287 XThR.Tn[3].n5 XThR.Tn[3].t11 24.9236
R19288 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19289 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19290 XThR.Tn[3].n6 XThR.Tn[3].t0 24.9236
R19291 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19292 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19293 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19294 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19295 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19296 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19297 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19298 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19299 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19300 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19301 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19302 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19303 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19304 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19305 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19306 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19307 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19308 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19309 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19310 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19311 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19312 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19313 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19314 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19315 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19316 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19317 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19318 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19319 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19320 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19321 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19322 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19323 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19324 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19325 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19326 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19327 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19328 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19329 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19330 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19331 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19332 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19333 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19334 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19335 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19336 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19337 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19338 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19339 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19340 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19341 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19342 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19343 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19344 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19345 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19346 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19347 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19348 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19349 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19350 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19351 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19352 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19353 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19354 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19355 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19356 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19357 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19358 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19359 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19360 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19361 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19362 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19363 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19364 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19365 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19366 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19367 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19368 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19369 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19370 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19371 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19372 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19373 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19374 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19375 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19376 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19377 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19378 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19379 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19380 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19381 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19382 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19383 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19384 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19385 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19386 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19387 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19388 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19389 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19390 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19391 XThR.Tn[5].n88 XThR.Tn[5].n87 332.332
R19392 XThR.Tn[5].n88 XThR.Tn[5].n86 296.493
R19393 XThR.Tn[5] XThR.Tn[5].n79 161.363
R19394 XThR.Tn[5] XThR.Tn[5].n74 161.363
R19395 XThR.Tn[5] XThR.Tn[5].n69 161.363
R19396 XThR.Tn[5] XThR.Tn[5].n64 161.363
R19397 XThR.Tn[5] XThR.Tn[5].n59 161.363
R19398 XThR.Tn[5] XThR.Tn[5].n54 161.363
R19399 XThR.Tn[5] XThR.Tn[5].n49 161.363
R19400 XThR.Tn[5] XThR.Tn[5].n44 161.363
R19401 XThR.Tn[5] XThR.Tn[5].n39 161.363
R19402 XThR.Tn[5] XThR.Tn[5].n34 161.363
R19403 XThR.Tn[5] XThR.Tn[5].n29 161.363
R19404 XThR.Tn[5] XThR.Tn[5].n24 161.363
R19405 XThR.Tn[5] XThR.Tn[5].n19 161.363
R19406 XThR.Tn[5] XThR.Tn[5].n14 161.363
R19407 XThR.Tn[5] XThR.Tn[5].n9 161.363
R19408 XThR.Tn[5] XThR.Tn[5].n7 161.363
R19409 XThR.Tn[5].n81 XThR.Tn[5].n80 161.3
R19410 XThR.Tn[5].n76 XThR.Tn[5].n75 161.3
R19411 XThR.Tn[5].n71 XThR.Tn[5].n70 161.3
R19412 XThR.Tn[5].n66 XThR.Tn[5].n65 161.3
R19413 XThR.Tn[5].n61 XThR.Tn[5].n60 161.3
R19414 XThR.Tn[5].n56 XThR.Tn[5].n55 161.3
R19415 XThR.Tn[5].n51 XThR.Tn[5].n50 161.3
R19416 XThR.Tn[5].n46 XThR.Tn[5].n45 161.3
R19417 XThR.Tn[5].n41 XThR.Tn[5].n40 161.3
R19418 XThR.Tn[5].n36 XThR.Tn[5].n35 161.3
R19419 XThR.Tn[5].n31 XThR.Tn[5].n30 161.3
R19420 XThR.Tn[5].n26 XThR.Tn[5].n25 161.3
R19421 XThR.Tn[5].n21 XThR.Tn[5].n20 161.3
R19422 XThR.Tn[5].n16 XThR.Tn[5].n15 161.3
R19423 XThR.Tn[5].n11 XThR.Tn[5].n10 161.3
R19424 XThR.Tn[5].n79 XThR.Tn[5].t62 161.106
R19425 XThR.Tn[5].n74 XThR.Tn[5].t70 161.106
R19426 XThR.Tn[5].n69 XThR.Tn[5].t52 161.106
R19427 XThR.Tn[5].n64 XThR.Tn[5].t35 161.106
R19428 XThR.Tn[5].n59 XThR.Tn[5].t60 161.106
R19429 XThR.Tn[5].n54 XThR.Tn[5].t24 161.106
R19430 XThR.Tn[5].n49 XThR.Tn[5].t68 161.106
R19431 XThR.Tn[5].n44 XThR.Tn[5].t49 161.106
R19432 XThR.Tn[5].n39 XThR.Tn[5].t32 161.106
R19433 XThR.Tn[5].n34 XThR.Tn[5].t40 161.106
R19434 XThR.Tn[5].n29 XThR.Tn[5].t22 161.106
R19435 XThR.Tn[5].n24 XThR.Tn[5].t51 161.106
R19436 XThR.Tn[5].n19 XThR.Tn[5].t21 161.106
R19437 XThR.Tn[5].n14 XThR.Tn[5].t66 161.106
R19438 XThR.Tn[5].n9 XThR.Tn[5].t26 161.106
R19439 XThR.Tn[5].n7 XThR.Tn[5].t72 161.106
R19440 XThR.Tn[5].n80 XThR.Tn[5].t59 159.978
R19441 XThR.Tn[5].n75 XThR.Tn[5].t64 159.978
R19442 XThR.Tn[5].n70 XThR.Tn[5].t47 159.978
R19443 XThR.Tn[5].n65 XThR.Tn[5].t31 159.978
R19444 XThR.Tn[5].n60 XThR.Tn[5].t57 159.978
R19445 XThR.Tn[5].n55 XThR.Tn[5].t20 159.978
R19446 XThR.Tn[5].n50 XThR.Tn[5].t63 159.978
R19447 XThR.Tn[5].n45 XThR.Tn[5].t45 159.978
R19448 XThR.Tn[5].n40 XThR.Tn[5].t29 159.978
R19449 XThR.Tn[5].n35 XThR.Tn[5].t37 159.978
R19450 XThR.Tn[5].n30 XThR.Tn[5].t19 159.978
R19451 XThR.Tn[5].n25 XThR.Tn[5].t46 159.978
R19452 XThR.Tn[5].n20 XThR.Tn[5].t18 159.978
R19453 XThR.Tn[5].n15 XThR.Tn[5].t61 159.978
R19454 XThR.Tn[5].n10 XThR.Tn[5].t23 159.978
R19455 XThR.Tn[5].n79 XThR.Tn[5].t54 145.038
R19456 XThR.Tn[5].n74 XThR.Tn[5].t12 145.038
R19457 XThR.Tn[5].n69 XThR.Tn[5].t56 145.038
R19458 XThR.Tn[5].n64 XThR.Tn[5].t41 145.038
R19459 XThR.Tn[5].n59 XThR.Tn[5].t71 145.038
R19460 XThR.Tn[5].n54 XThR.Tn[5].t53 145.038
R19461 XThR.Tn[5].n49 XThR.Tn[5].t58 145.038
R19462 XThR.Tn[5].n44 XThR.Tn[5].t42 145.038
R19463 XThR.Tn[5].n39 XThR.Tn[5].t38 145.038
R19464 XThR.Tn[5].n34 XThR.Tn[5].t69 145.038
R19465 XThR.Tn[5].n29 XThR.Tn[5].t30 145.038
R19466 XThR.Tn[5].n24 XThR.Tn[5].t55 145.038
R19467 XThR.Tn[5].n19 XThR.Tn[5].t28 145.038
R19468 XThR.Tn[5].n14 XThR.Tn[5].t73 145.038
R19469 XThR.Tn[5].n9 XThR.Tn[5].t39 145.038
R19470 XThR.Tn[5].n7 XThR.Tn[5].t17 145.038
R19471 XThR.Tn[5].n80 XThR.Tn[5].t27 143.911
R19472 XThR.Tn[5].n75 XThR.Tn[5].t50 143.911
R19473 XThR.Tn[5].n70 XThR.Tn[5].t34 143.911
R19474 XThR.Tn[5].n65 XThR.Tn[5].t15 143.911
R19475 XThR.Tn[5].n60 XThR.Tn[5].t44 143.911
R19476 XThR.Tn[5].n55 XThR.Tn[5].t25 143.911
R19477 XThR.Tn[5].n50 XThR.Tn[5].t36 143.911
R19478 XThR.Tn[5].n45 XThR.Tn[5].t16 143.911
R19479 XThR.Tn[5].n40 XThR.Tn[5].t14 143.911
R19480 XThR.Tn[5].n35 XThR.Tn[5].t43 143.911
R19481 XThR.Tn[5].n30 XThR.Tn[5].t67 143.911
R19482 XThR.Tn[5].n25 XThR.Tn[5].t33 143.911
R19483 XThR.Tn[5].n20 XThR.Tn[5].t65 143.911
R19484 XThR.Tn[5].n15 XThR.Tn[5].t48 143.911
R19485 XThR.Tn[5].n10 XThR.Tn[5].t13 143.911
R19486 XThR.Tn[5].n2 XThR.Tn[5].n0 135.249
R19487 XThR.Tn[5].n2 XThR.Tn[5].n1 98.981
R19488 XThR.Tn[5].n4 XThR.Tn[5].n3 98.981
R19489 XThR.Tn[5].n6 XThR.Tn[5].n5 98.981
R19490 XThR.Tn[5].n4 XThR.Tn[5].n2 36.2672
R19491 XThR.Tn[5].n6 XThR.Tn[5].n4 36.2672
R19492 XThR.Tn[5].n85 XThR.Tn[5].n6 32.6405
R19493 XThR.Tn[5].n87 XThR.Tn[5].t1 26.5955
R19494 XThR.Tn[5].n87 XThR.Tn[5].t0 26.5955
R19495 XThR.Tn[5].n86 XThR.Tn[5].t2 26.5955
R19496 XThR.Tn[5].n86 XThR.Tn[5].t3 26.5955
R19497 XThR.Tn[5].n0 XThR.Tn[5].t8 24.9236
R19498 XThR.Tn[5].n0 XThR.Tn[5].t9 24.9236
R19499 XThR.Tn[5].n1 XThR.Tn[5].t11 24.9236
R19500 XThR.Tn[5].n1 XThR.Tn[5].t10 24.9236
R19501 XThR.Tn[5].n3 XThR.Tn[5].t6 24.9236
R19502 XThR.Tn[5].n3 XThR.Tn[5].t5 24.9236
R19503 XThR.Tn[5].n5 XThR.Tn[5].t7 24.9236
R19504 XThR.Tn[5].n5 XThR.Tn[5].t4 24.9236
R19505 XThR.Tn[5].n89 XThR.Tn[5].n88 18.5605
R19506 XThR.Tn[5].n89 XThR.Tn[5].n85 11.5205
R19507 XThR.Tn[5].n85 XThR.Tn[5] 5.71508
R19508 XThR.Tn[5] XThR.Tn[5].n8 5.34038
R19509 XThR.Tn[5].n13 XThR.Tn[5].n12 4.5005
R19510 XThR.Tn[5].n18 XThR.Tn[5].n17 4.5005
R19511 XThR.Tn[5].n23 XThR.Tn[5].n22 4.5005
R19512 XThR.Tn[5].n28 XThR.Tn[5].n27 4.5005
R19513 XThR.Tn[5].n33 XThR.Tn[5].n32 4.5005
R19514 XThR.Tn[5].n38 XThR.Tn[5].n37 4.5005
R19515 XThR.Tn[5].n43 XThR.Tn[5].n42 4.5005
R19516 XThR.Tn[5].n48 XThR.Tn[5].n47 4.5005
R19517 XThR.Tn[5].n53 XThR.Tn[5].n52 4.5005
R19518 XThR.Tn[5].n58 XThR.Tn[5].n57 4.5005
R19519 XThR.Tn[5].n63 XThR.Tn[5].n62 4.5005
R19520 XThR.Tn[5].n68 XThR.Tn[5].n67 4.5005
R19521 XThR.Tn[5].n73 XThR.Tn[5].n72 4.5005
R19522 XThR.Tn[5].n78 XThR.Tn[5].n77 4.5005
R19523 XThR.Tn[5].n83 XThR.Tn[5].n82 4.5005
R19524 XThR.Tn[5].n84 XThR.Tn[5] 3.70586
R19525 XThR.Tn[5].n13 XThR.Tn[5] 2.52282
R19526 XThR.Tn[5].n18 XThR.Tn[5] 2.52282
R19527 XThR.Tn[5].n23 XThR.Tn[5] 2.52282
R19528 XThR.Tn[5].n28 XThR.Tn[5] 2.52282
R19529 XThR.Tn[5].n33 XThR.Tn[5] 2.52282
R19530 XThR.Tn[5].n38 XThR.Tn[5] 2.52282
R19531 XThR.Tn[5].n43 XThR.Tn[5] 2.52282
R19532 XThR.Tn[5].n48 XThR.Tn[5] 2.52282
R19533 XThR.Tn[5].n53 XThR.Tn[5] 2.52282
R19534 XThR.Tn[5].n58 XThR.Tn[5] 2.52282
R19535 XThR.Tn[5].n63 XThR.Tn[5] 2.52282
R19536 XThR.Tn[5].n68 XThR.Tn[5] 2.52282
R19537 XThR.Tn[5].n73 XThR.Tn[5] 2.52282
R19538 XThR.Tn[5].n78 XThR.Tn[5] 2.52282
R19539 XThR.Tn[5].n83 XThR.Tn[5] 2.52282
R19540 XThR.Tn[5].n81 XThR.Tn[5] 1.08677
R19541 XThR.Tn[5].n76 XThR.Tn[5] 1.08677
R19542 XThR.Tn[5].n71 XThR.Tn[5] 1.08677
R19543 XThR.Tn[5].n66 XThR.Tn[5] 1.08677
R19544 XThR.Tn[5].n61 XThR.Tn[5] 1.08677
R19545 XThR.Tn[5].n56 XThR.Tn[5] 1.08677
R19546 XThR.Tn[5].n51 XThR.Tn[5] 1.08677
R19547 XThR.Tn[5].n46 XThR.Tn[5] 1.08677
R19548 XThR.Tn[5].n41 XThR.Tn[5] 1.08677
R19549 XThR.Tn[5].n36 XThR.Tn[5] 1.08677
R19550 XThR.Tn[5].n31 XThR.Tn[5] 1.08677
R19551 XThR.Tn[5].n26 XThR.Tn[5] 1.08677
R19552 XThR.Tn[5].n21 XThR.Tn[5] 1.08677
R19553 XThR.Tn[5].n16 XThR.Tn[5] 1.08677
R19554 XThR.Tn[5].n11 XThR.Tn[5] 1.08677
R19555 XThR.Tn[5] XThR.Tn[5].n13 0.839786
R19556 XThR.Tn[5] XThR.Tn[5].n18 0.839786
R19557 XThR.Tn[5] XThR.Tn[5].n23 0.839786
R19558 XThR.Tn[5] XThR.Tn[5].n28 0.839786
R19559 XThR.Tn[5] XThR.Tn[5].n33 0.839786
R19560 XThR.Tn[5] XThR.Tn[5].n38 0.839786
R19561 XThR.Tn[5] XThR.Tn[5].n43 0.839786
R19562 XThR.Tn[5] XThR.Tn[5].n48 0.839786
R19563 XThR.Tn[5] XThR.Tn[5].n53 0.839786
R19564 XThR.Tn[5] XThR.Tn[5].n58 0.839786
R19565 XThR.Tn[5] XThR.Tn[5].n63 0.839786
R19566 XThR.Tn[5] XThR.Tn[5].n68 0.839786
R19567 XThR.Tn[5] XThR.Tn[5].n73 0.839786
R19568 XThR.Tn[5] XThR.Tn[5].n78 0.839786
R19569 XThR.Tn[5] XThR.Tn[5].n83 0.839786
R19570 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19571 XThR.Tn[5].n8 XThR.Tn[5] 0.499542
R19572 XThR.Tn[5].n82 XThR.Tn[5] 0.063
R19573 XThR.Tn[5].n77 XThR.Tn[5] 0.063
R19574 XThR.Tn[5].n72 XThR.Tn[5] 0.063
R19575 XThR.Tn[5].n67 XThR.Tn[5] 0.063
R19576 XThR.Tn[5].n62 XThR.Tn[5] 0.063
R19577 XThR.Tn[5].n57 XThR.Tn[5] 0.063
R19578 XThR.Tn[5].n52 XThR.Tn[5] 0.063
R19579 XThR.Tn[5].n47 XThR.Tn[5] 0.063
R19580 XThR.Tn[5].n42 XThR.Tn[5] 0.063
R19581 XThR.Tn[5].n37 XThR.Tn[5] 0.063
R19582 XThR.Tn[5].n32 XThR.Tn[5] 0.063
R19583 XThR.Tn[5].n27 XThR.Tn[5] 0.063
R19584 XThR.Tn[5].n22 XThR.Tn[5] 0.063
R19585 XThR.Tn[5].n17 XThR.Tn[5] 0.063
R19586 XThR.Tn[5].n12 XThR.Tn[5] 0.063
R19587 XThR.Tn[5].n84 XThR.Tn[5] 0.0540714
R19588 XThR.Tn[5] XThR.Tn[5].n84 0.038
R19589 XThR.Tn[5].n8 XThR.Tn[5] 0.0143889
R19590 XThR.Tn[5].n82 XThR.Tn[5].n81 0.00771154
R19591 XThR.Tn[5].n77 XThR.Tn[5].n76 0.00771154
R19592 XThR.Tn[5].n72 XThR.Tn[5].n71 0.00771154
R19593 XThR.Tn[5].n67 XThR.Tn[5].n66 0.00771154
R19594 XThR.Tn[5].n62 XThR.Tn[5].n61 0.00771154
R19595 XThR.Tn[5].n57 XThR.Tn[5].n56 0.00771154
R19596 XThR.Tn[5].n52 XThR.Tn[5].n51 0.00771154
R19597 XThR.Tn[5].n47 XThR.Tn[5].n46 0.00771154
R19598 XThR.Tn[5].n42 XThR.Tn[5].n41 0.00771154
R19599 XThR.Tn[5].n37 XThR.Tn[5].n36 0.00771154
R19600 XThR.Tn[5].n32 XThR.Tn[5].n31 0.00771154
R19601 XThR.Tn[5].n27 XThR.Tn[5].n26 0.00771154
R19602 XThR.Tn[5].n22 XThR.Tn[5].n21 0.00771154
R19603 XThR.Tn[5].n17 XThR.Tn[5].n16 0.00771154
R19604 XThR.Tn[5].n12 XThR.Tn[5].n11 0.00771154
R19605 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R19606 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R19607 XThC.Tn[4].n71 XThC.Tn[4].n69 161.365
R19608 XThC.Tn[4].n67 XThC.Tn[4].n65 161.365
R19609 XThC.Tn[4].n63 XThC.Tn[4].n61 161.365
R19610 XThC.Tn[4].n59 XThC.Tn[4].n57 161.365
R19611 XThC.Tn[4].n55 XThC.Tn[4].n53 161.365
R19612 XThC.Tn[4].n51 XThC.Tn[4].n49 161.365
R19613 XThC.Tn[4].n47 XThC.Tn[4].n45 161.365
R19614 XThC.Tn[4].n43 XThC.Tn[4].n41 161.365
R19615 XThC.Tn[4].n39 XThC.Tn[4].n37 161.365
R19616 XThC.Tn[4].n35 XThC.Tn[4].n33 161.365
R19617 XThC.Tn[4].n31 XThC.Tn[4].n29 161.365
R19618 XThC.Tn[4].n27 XThC.Tn[4].n25 161.365
R19619 XThC.Tn[4].n23 XThC.Tn[4].n21 161.365
R19620 XThC.Tn[4].n19 XThC.Tn[4].n17 161.365
R19621 XThC.Tn[4].n15 XThC.Tn[4].n13 161.365
R19622 XThC.Tn[4].n12 XThC.Tn[4].n10 161.365
R19623 XThC.Tn[4].n69 XThC.Tn[4].t32 161.202
R19624 XThC.Tn[4].n65 XThC.Tn[4].t22 161.202
R19625 XThC.Tn[4].n61 XThC.Tn[4].t41 161.202
R19626 XThC.Tn[4].n57 XThC.Tn[4].t38 161.202
R19627 XThC.Tn[4].n53 XThC.Tn[4].t30 161.202
R19628 XThC.Tn[4].n49 XThC.Tn[4].t17 161.202
R19629 XThC.Tn[4].n45 XThC.Tn[4].t16 161.202
R19630 XThC.Tn[4].n41 XThC.Tn[4].t29 161.202
R19631 XThC.Tn[4].n37 XThC.Tn[4].t27 161.202
R19632 XThC.Tn[4].n33 XThC.Tn[4].t18 161.202
R19633 XThC.Tn[4].n29 XThC.Tn[4].t37 161.202
R19634 XThC.Tn[4].n25 XThC.Tn[4].t36 161.202
R19635 XThC.Tn[4].n21 XThC.Tn[4].t15 161.202
R19636 XThC.Tn[4].n17 XThC.Tn[4].t13 161.202
R19637 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R19638 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R19639 XThC.Tn[4].n69 XThC.Tn[4].t35 145.137
R19640 XThC.Tn[4].n65 XThC.Tn[4].t25 145.137
R19641 XThC.Tn[4].n61 XThC.Tn[4].t12 145.137
R19642 XThC.Tn[4].n57 XThC.Tn[4].t42 145.137
R19643 XThC.Tn[4].n53 XThC.Tn[4].t34 145.137
R19644 XThC.Tn[4].n49 XThC.Tn[4].t23 145.137
R19645 XThC.Tn[4].n45 XThC.Tn[4].t21 145.137
R19646 XThC.Tn[4].n41 XThC.Tn[4].t33 145.137
R19647 XThC.Tn[4].n37 XThC.Tn[4].t31 145.137
R19648 XThC.Tn[4].n33 XThC.Tn[4].t24 145.137
R19649 XThC.Tn[4].n29 XThC.Tn[4].t40 145.137
R19650 XThC.Tn[4].n25 XThC.Tn[4].t39 145.137
R19651 XThC.Tn[4].n21 XThC.Tn[4].t20 145.137
R19652 XThC.Tn[4].n17 XThC.Tn[4].t19 145.137
R19653 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R19654 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R19655 XThC.Tn[4].n6 XThC.Tn[4].n4 135.248
R19656 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R19657 XThC.Tn[4].n6 XThC.Tn[4].n5 98.982
R19658 XThC.Tn[4].n8 XThC.Tn[4].n7 98.982
R19659 XThC.Tn[4].n8 XThC.Tn[4].n6 36.2672
R19660 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R19661 XThC.Tn[4].n73 XThC.Tn[4].n9 32.6405
R19662 XThC.Tn[4].n1 XThC.Tn[4].t7 26.5955
R19663 XThC.Tn[4].n1 XThC.Tn[4].t6 26.5955
R19664 XThC.Tn[4].n0 XThC.Tn[4].t5 26.5955
R19665 XThC.Tn[4].n0 XThC.Tn[4].t4 26.5955
R19666 XThC.Tn[4].n3 XThC.Tn[4].t1 24.9236
R19667 XThC.Tn[4].n3 XThC.Tn[4].t0 24.9236
R19668 XThC.Tn[4].n4 XThC.Tn[4].t8 24.9236
R19669 XThC.Tn[4].n4 XThC.Tn[4].t11 24.9236
R19670 XThC.Tn[4].n5 XThC.Tn[4].t10 24.9236
R19671 XThC.Tn[4].n5 XThC.Tn[4].t9 24.9236
R19672 XThC.Tn[4].n7 XThC.Tn[4].t3 24.9236
R19673 XThC.Tn[4].n7 XThC.Tn[4].t2 24.9236
R19674 XThC.Tn[4].n74 XThC.Tn[4].n2 18.5605
R19675 XThC.Tn[4].n74 XThC.Tn[4].n73 11.5205
R19676 XThC.Tn[4] XThC.Tn[4].n12 8.0245
R19677 XThC.Tn[4].n72 XThC.Tn[4].n71 7.9105
R19678 XThC.Tn[4].n68 XThC.Tn[4].n67 7.9105
R19679 XThC.Tn[4].n64 XThC.Tn[4].n63 7.9105
R19680 XThC.Tn[4].n60 XThC.Tn[4].n59 7.9105
R19681 XThC.Tn[4].n56 XThC.Tn[4].n55 7.9105
R19682 XThC.Tn[4].n52 XThC.Tn[4].n51 7.9105
R19683 XThC.Tn[4].n48 XThC.Tn[4].n47 7.9105
R19684 XThC.Tn[4].n44 XThC.Tn[4].n43 7.9105
R19685 XThC.Tn[4].n40 XThC.Tn[4].n39 7.9105
R19686 XThC.Tn[4].n36 XThC.Tn[4].n35 7.9105
R19687 XThC.Tn[4].n32 XThC.Tn[4].n31 7.9105
R19688 XThC.Tn[4].n28 XThC.Tn[4].n27 7.9105
R19689 XThC.Tn[4].n24 XThC.Tn[4].n23 7.9105
R19690 XThC.Tn[4].n20 XThC.Tn[4].n19 7.9105
R19691 XThC.Tn[4].n16 XThC.Tn[4].n15 7.9105
R19692 XThC.Tn[4].n73 XThC.Tn[4] 5.77342
R19693 XThC.Tn[4] XThC.Tn[4].n74 0.6405
R19694 XThC.Tn[4].n16 XThC.Tn[4] 0.235138
R19695 XThC.Tn[4].n20 XThC.Tn[4] 0.235138
R19696 XThC.Tn[4].n24 XThC.Tn[4] 0.235138
R19697 XThC.Tn[4].n28 XThC.Tn[4] 0.235138
R19698 XThC.Tn[4].n32 XThC.Tn[4] 0.235138
R19699 XThC.Tn[4].n36 XThC.Tn[4] 0.235138
R19700 XThC.Tn[4].n40 XThC.Tn[4] 0.235138
R19701 XThC.Tn[4].n44 XThC.Tn[4] 0.235138
R19702 XThC.Tn[4].n48 XThC.Tn[4] 0.235138
R19703 XThC.Tn[4].n52 XThC.Tn[4] 0.235138
R19704 XThC.Tn[4].n56 XThC.Tn[4] 0.235138
R19705 XThC.Tn[4].n60 XThC.Tn[4] 0.235138
R19706 XThC.Tn[4].n64 XThC.Tn[4] 0.235138
R19707 XThC.Tn[4].n68 XThC.Tn[4] 0.235138
R19708 XThC.Tn[4].n72 XThC.Tn[4] 0.235138
R19709 XThC.Tn[4] XThC.Tn[4].n16 0.114505
R19710 XThC.Tn[4] XThC.Tn[4].n20 0.114505
R19711 XThC.Tn[4] XThC.Tn[4].n24 0.114505
R19712 XThC.Tn[4] XThC.Tn[4].n28 0.114505
R19713 XThC.Tn[4] XThC.Tn[4].n32 0.114505
R19714 XThC.Tn[4] XThC.Tn[4].n36 0.114505
R19715 XThC.Tn[4] XThC.Tn[4].n40 0.114505
R19716 XThC.Tn[4] XThC.Tn[4].n44 0.114505
R19717 XThC.Tn[4] XThC.Tn[4].n48 0.114505
R19718 XThC.Tn[4] XThC.Tn[4].n52 0.114505
R19719 XThC.Tn[4] XThC.Tn[4].n56 0.114505
R19720 XThC.Tn[4] XThC.Tn[4].n60 0.114505
R19721 XThC.Tn[4] XThC.Tn[4].n64 0.114505
R19722 XThC.Tn[4] XThC.Tn[4].n68 0.114505
R19723 XThC.Tn[4] XThC.Tn[4].n72 0.114505
R19724 XThC.Tn[4].n71 XThC.Tn[4].n70 0.0599512
R19725 XThC.Tn[4].n67 XThC.Tn[4].n66 0.0599512
R19726 XThC.Tn[4].n63 XThC.Tn[4].n62 0.0599512
R19727 XThC.Tn[4].n59 XThC.Tn[4].n58 0.0599512
R19728 XThC.Tn[4].n55 XThC.Tn[4].n54 0.0599512
R19729 XThC.Tn[4].n51 XThC.Tn[4].n50 0.0599512
R19730 XThC.Tn[4].n47 XThC.Tn[4].n46 0.0599512
R19731 XThC.Tn[4].n43 XThC.Tn[4].n42 0.0599512
R19732 XThC.Tn[4].n39 XThC.Tn[4].n38 0.0599512
R19733 XThC.Tn[4].n35 XThC.Tn[4].n34 0.0599512
R19734 XThC.Tn[4].n31 XThC.Tn[4].n30 0.0599512
R19735 XThC.Tn[4].n27 XThC.Tn[4].n26 0.0599512
R19736 XThC.Tn[4].n23 XThC.Tn[4].n22 0.0599512
R19737 XThC.Tn[4].n19 XThC.Tn[4].n18 0.0599512
R19738 XThC.Tn[4].n15 XThC.Tn[4].n14 0.0599512
R19739 XThC.Tn[4].n12 XThC.Tn[4].n11 0.0599512
R19740 XThC.Tn[4].n70 XThC.Tn[4] 0.0469286
R19741 XThC.Tn[4].n66 XThC.Tn[4] 0.0469286
R19742 XThC.Tn[4].n62 XThC.Tn[4] 0.0469286
R19743 XThC.Tn[4].n58 XThC.Tn[4] 0.0469286
R19744 XThC.Tn[4].n54 XThC.Tn[4] 0.0469286
R19745 XThC.Tn[4].n50 XThC.Tn[4] 0.0469286
R19746 XThC.Tn[4].n46 XThC.Tn[4] 0.0469286
R19747 XThC.Tn[4].n42 XThC.Tn[4] 0.0469286
R19748 XThC.Tn[4].n38 XThC.Tn[4] 0.0469286
R19749 XThC.Tn[4].n34 XThC.Tn[4] 0.0469286
R19750 XThC.Tn[4].n30 XThC.Tn[4] 0.0469286
R19751 XThC.Tn[4].n26 XThC.Tn[4] 0.0469286
R19752 XThC.Tn[4].n22 XThC.Tn[4] 0.0469286
R19753 XThC.Tn[4].n18 XThC.Tn[4] 0.0469286
R19754 XThC.Tn[4].n14 XThC.Tn[4] 0.0469286
R19755 XThC.Tn[4].n11 XThC.Tn[4] 0.0469286
R19756 XThC.Tn[4].n70 XThC.Tn[4] 0.0401341
R19757 XThC.Tn[4].n66 XThC.Tn[4] 0.0401341
R19758 XThC.Tn[4].n62 XThC.Tn[4] 0.0401341
R19759 XThC.Tn[4].n58 XThC.Tn[4] 0.0401341
R19760 XThC.Tn[4].n54 XThC.Tn[4] 0.0401341
R19761 XThC.Tn[4].n50 XThC.Tn[4] 0.0401341
R19762 XThC.Tn[4].n46 XThC.Tn[4] 0.0401341
R19763 XThC.Tn[4].n42 XThC.Tn[4] 0.0401341
R19764 XThC.Tn[4].n38 XThC.Tn[4] 0.0401341
R19765 XThC.Tn[4].n34 XThC.Tn[4] 0.0401341
R19766 XThC.Tn[4].n30 XThC.Tn[4] 0.0401341
R19767 XThC.Tn[4].n26 XThC.Tn[4] 0.0401341
R19768 XThC.Tn[4].n22 XThC.Tn[4] 0.0401341
R19769 XThC.Tn[4].n18 XThC.Tn[4] 0.0401341
R19770 XThC.Tn[4].n14 XThC.Tn[4] 0.0401341
R19771 XThC.Tn[4].n11 XThC.Tn[4] 0.0401341
R19772 Iout.n1020 Iout.t148 239.927
R19773 Iout.n509 Iout.t20 239.927
R19774 Iout.n513 Iout.t65 239.927
R19775 Iout.n507 Iout.t112 239.927
R19776 Iout.n504 Iout.t241 239.927
R19777 Iout.n500 Iout.t197 239.927
R19778 Iout.n192 Iout.t157 239.927
R19779 Iout.n195 Iout.t253 239.927
R19780 Iout.n199 Iout.t140 239.927
R19781 Iout.n202 Iout.t231 239.927
R19782 Iout.n206 Iout.t194 239.927
R19783 Iout.n210 Iout.t83 239.927
R19784 Iout.n214 Iout.t90 239.927
R19785 Iout.n218 Iout.t33 239.927
R19786 Iout.n222 Iout.t206 239.927
R19787 Iout.n226 Iout.t208 239.927
R19788 Iout.n232 Iout.t159 239.927
R19789 Iout.n235 Iout.t114 239.927
R19790 Iout.n238 Iout.t143 239.927
R19791 Iout.n241 Iout.t18 239.927
R19792 Iout.n244 Iout.t131 239.927
R19793 Iout.n247 Iout.t215 239.927
R19794 Iout.n250 Iout.t173 239.927
R19795 Iout.n255 Iout.t47 239.927
R19796 Iout.n252 Iout.t29 239.927
R19797 Iout.n489 Iout.t38 239.927
R19798 Iout.n494 Iout.t34 239.927
R19799 Iout.n491 Iout.t55 239.927
R19800 Iout.n519 Iout.t2 239.927
R19801 Iout.n149 Iout.t228 239.927
R19802 Iout.n146 Iout.t227 239.927
R19803 Iout.n1010 Iout.t149 239.927
R19804 Iout.n1007 Iout.t191 239.927
R19805 Iout.n140 Iout.t86 239.927
R19806 Iout.n143 Iout.t239 239.927
R19807 Iout.n525 Iout.t130 239.927
R19808 Iout.n480 Iout.t58 239.927
R19809 Iout.n483 Iout.t243 239.927
R19810 Iout.n478 Iout.t167 239.927
R19811 Iout.n259 Iout.t134 239.927
R19812 Iout.n186 Iout.t19 239.927
R19813 Iout.n271 Iout.t45 239.927
R19814 Iout.n180 Iout.t43 239.927
R19815 Iout.n283 Iout.t101 239.927
R19816 Iout.n174 Iout.t4 239.927
R19817 Iout.n168 Iout.t203 239.927
R19818 Iout.n301 Iout.t153 239.927
R19819 Iout.n289 Iout.t74 239.927
R19820 Iout.n177 Iout.t78 239.927
R19821 Iout.n277 Iout.t195 239.927
R19822 Iout.n183 Iout.t174 239.927
R19823 Iout.n265 Iout.t117 239.927
R19824 Iout.n189 Iout.t255 239.927
R19825 Iout.n472 Iout.t201 239.927
R19826 Iout.n469 Iout.t166 239.927
R19827 Iout.n156 Iout.t220 239.927
R19828 Iout.n531 Iout.t59 239.927
R19829 Iout.n534 Iout.t146 239.927
R19830 Iout.n536 Iout.t75 239.927
R19831 Iout.n133 Iout.t113 239.927
R19832 Iout.n136 Iout.t91 239.927
R19833 Iout.n542 Iout.t119 239.927
R19834 Iout.n460 Iout.t186 239.927
R19835 Iout.n463 Iout.t158 239.927
R19836 Iout.n458 Iout.t27 239.927
R19837 Iout.n305 Iout.t181 239.927
R19838 Iout.n308 Iout.t237 239.927
R19839 Iout.n311 Iout.t154 239.927
R19840 Iout.n314 Iout.t10 239.927
R19841 Iout.n317 Iout.t250 239.927
R19842 Iout.n320 Iout.t7 239.927
R19843 Iout.n392 Iout.t152 239.927
R19844 Iout.n378 Iout.t12 239.927
R19845 Iout.n376 Iout.t121 239.927
R19846 Iout.n394 Iout.t165 239.927
R19847 Iout.n408 Iout.t61 239.927
R19848 Iout.n410 Iout.t199 239.927
R19849 Iout.n424 Iout.t190 239.927
R19850 Iout.n426 Iout.t88 239.927
R19851 Iout.n447 Iout.t232 239.927
R19852 Iout.n452 Iout.t129 239.927
R19853 Iout.n449 Iout.t252 239.927
R19854 Iout.n548 Iout.t122 239.927
R19855 Iout.n130 Iout.t87 239.927
R19856 Iout.n559 Iout.t14 239.927
R19857 Iout.n557 Iout.t178 239.927
R19858 Iout.n554 Iout.t171 239.927
R19859 Iout.n434 Iout.t155 239.927
R19860 Iout.n438 Iout.t6 239.927
R19861 Iout.n441 Iout.t214 239.927
R19862 Iout.n432 Iout.t106 239.927
R19863 Iout.n418 Iout.t198 239.927
R19864 Iout.n416 Iout.t51 239.927
R19865 Iout.n402 Iout.t172 239.927
R19866 Iout.n357 Iout.t107 239.927
R19867 Iout.n360 Iout.t147 239.927
R19868 Iout.n363 Iout.t31 239.927
R19869 Iout.n366 Iout.t226 239.927
R19870 Iout.n354 Iout.t209 239.927
R19871 Iout.n351 Iout.t13 239.927
R19872 Iout.n348 Iout.t213 239.927
R19873 Iout.n345 Iout.t210 239.927
R19874 Iout.n342 Iout.t205 239.927
R19875 Iout.n339 Iout.t230 239.927
R19876 Iout.n336 Iout.t17 239.927
R19877 Iout.n333 Iout.t234 239.927
R19878 Iout.n117 Iout.t124 239.927
R19879 Iout.n582 Iout.t222 239.927
R19880 Iout.n111 Iout.t105 239.927
R19881 Iout.n594 Iout.t175 239.927
R19882 Iout.n105 Iout.t251 239.927
R19883 Iout.n606 Iout.t39 239.927
R19884 Iout.n99 Iout.t246 239.927
R19885 Iout.n618 Iout.t132 239.927
R19886 Iout.n624 Iout.t202 239.927
R19887 Iout.n90 Iout.t254 239.927
R19888 Iout.n636 Iout.t64 239.927
R19889 Iout.n81 Iout.t110 239.927
R19890 Iout.n648 Iout.t71 239.927
R19891 Iout.n96 Iout.t1 239.927
R19892 Iout.n612 Iout.t62 239.927
R19893 Iout.n102 Iout.t240 239.927
R19894 Iout.n600 Iout.t22 239.927
R19895 Iout.n108 Iout.t9 239.927
R19896 Iout.n588 Iout.t179 239.927
R19897 Iout.n687 Iout.t170 239.927
R19898 Iout.n684 Iout.t116 239.927
R19899 Iout.n681 Iout.t247 239.927
R19900 Iout.n678 Iout.t40 239.927
R19901 Iout.n675 Iout.t94 239.927
R19902 Iout.n672 Iout.t185 239.927
R19903 Iout.n747 Iout.t53 239.927
R19904 Iout.n50 Iout.t56 239.927
R19905 Iout.n759 Iout.t126 239.927
R19906 Iout.n44 Iout.t100 239.927
R19907 Iout.n771 Iout.t69 239.927
R19908 Iout.n42 Iout.t30 239.927
R19909 Iout.n56 Iout.t32 239.927
R19910 Iout.n735 Iout.t200 239.927
R19911 Iout.n62 Iout.t68 239.927
R19912 Iout.n723 Iout.t109 239.927
R19913 Iout.n717 Iout.t125 239.927
R19914 Iout.n65 Iout.t82 239.927
R19915 Iout.n729 Iout.t169 239.927
R19916 Iout.n59 Iout.t5 239.927
R19917 Iout.n805 Iout.t123 239.927
R19918 Iout.n808 Iout.t80 239.927
R19919 Iout.n811 Iout.t70 239.927
R19920 Iout.n814 Iout.t8 239.927
R19921 Iout.n817 Iout.t211 239.927
R19922 Iout.n820 Iout.t36 239.927
R19923 Iout.n823 Iout.t156 239.927
R19924 Iout.n802 Iout.t238 239.927
R19925 Iout.n799 Iout.t23 239.927
R19926 Iout.n890 Iout.t76 239.927
R19927 Iout.n888 Iout.t192 239.927
R19928 Iout.n881 Iout.t103 239.927
R19929 Iout.n869 Iout.t49 239.927
R19930 Iout.n867 Iout.t37 239.927
R19931 Iout.n855 Iout.t72 239.927
R19932 Iout.n853 Iout.t150 239.927
R19933 Iout.n841 Iout.t41 239.927
R19934 Iout.n839 Iout.t46 239.927
R19935 Iout.n827 Iout.t176 239.927
R19936 Iout.n883 Iout.t162 239.927
R19937 Iout.n895 Iout.t219 239.927
R19938 Iout.n897 Iout.t44 239.927
R19939 Iout.n909 Iout.t16 239.927
R19940 Iout.n911 Iout.t95 239.927
R19941 Iout.n923 Iout.t135 239.927
R19942 Iout.n926 Iout.t108 239.927
R19943 Iout.n22 Iout.t224 239.927
R19944 Iout.n876 Iout.t104 239.927
R19945 Iout.n874 Iout.t182 239.927
R19946 Iout.n862 Iout.t188 239.927
R19947 Iout.n860 Iout.t164 239.927
R19948 Iout.n848 Iout.t236 239.927
R19949 Iout.n846 Iout.t151 239.927
R19950 Iout.n834 Iout.t25 239.927
R19951 Iout.n832 Iout.t52 239.927
R19952 Iout.n902 Iout.t137 239.927
R19953 Iout.n904 Iout.t248 239.927
R19954 Iout.n916 Iout.t249 239.927
R19955 Iout.n918 Iout.t184 239.927
R19956 Iout.n931 Iout.t67 239.927
R19957 Iout.n934 Iout.t73 239.927
R19958 Iout.n796 Iout.t77 239.927
R19959 Iout.n793 Iout.t111 239.927
R19960 Iout.n790 Iout.t144 239.927
R19961 Iout.n787 Iout.t28 239.927
R19962 Iout.n784 Iout.t221 239.927
R19963 Iout.n781 Iout.t235 239.927
R19964 Iout.n938 Iout.t244 239.927
R19965 Iout.n741 Iout.t63 239.927
R19966 Iout.n53 Iout.t145 239.927
R19967 Iout.n753 Iout.t98 239.927
R19968 Iout.n47 Iout.t168 239.927
R19969 Iout.n765 Iout.t127 239.927
R19970 Iout.n38 Iout.t92 239.927
R19971 Iout.n777 Iout.t81 239.927
R19972 Iout.n71 Iout.t136 239.927
R19973 Iout.n705 Iout.t11 239.927
R19974 Iout.n77 Iout.t128 239.927
R19975 Iout.n944 Iout.t216 239.927
R19976 Iout.n19 Iout.t85 239.927
R19977 Iout.n68 Iout.t242 239.927
R19978 Iout.n711 Iout.t233 239.927
R19979 Iout.n74 Iout.t223 239.927
R19980 Iout.n699 Iout.t26 239.927
R19981 Iout.n950 Iout.t187 239.927
R19982 Iout.n953 Iout.t204 239.927
R19983 Iout.n669 Iout.t141 239.927
R19984 Iout.n666 Iout.t163 239.927
R19985 Iout.n663 Iout.t3 239.927
R19986 Iout.n660 Iout.t35 239.927
R19987 Iout.n657 Iout.t245 239.927
R19988 Iout.n654 Iout.t180 239.927
R19989 Iout.n690 Iout.t97 239.927
R19990 Iout.n695 Iout.t54 239.927
R19991 Iout.n692 Iout.t225 239.927
R19992 Iout.n957 Iout.t89 239.927
R19993 Iout.n114 Iout.t133 239.927
R19994 Iout.n576 Iout.t177 239.927
R19995 Iout.n573 Iout.t161 239.927
R19996 Iout.n963 Iout.t48 239.927
R19997 Iout.n14 Iout.t142 239.927
R19998 Iout.n93 Iout.t42 239.927
R19999 Iout.n630 Iout.t84 239.927
R20000 Iout.n87 Iout.t138 239.927
R20001 Iout.n642 Iout.t120 239.927
R20002 Iout.n85 Iout.t60 239.927
R20003 Iout.n563 Iout.t15 239.927
R20004 Iout.n969 Iout.t189 239.927
R20005 Iout.n972 Iout.t118 239.927
R20006 Iout.n569 Iout.t79 239.927
R20007 Iout.n123 Iout.t96 239.927
R20008 Iout.n120 Iout.t21 239.927
R20009 Iout.n976 Iout.t207 239.927
R20010 Iout.n400 Iout.t50 239.927
R20011 Iout.n386 Iout.t99 239.927
R20012 Iout.n384 Iout.t24 239.927
R20013 Iout.n370 Iout.t139 239.927
R20014 Iout.n982 Iout.t115 239.927
R20015 Iout.n9 Iout.t0 239.927
R20016 Iout.n127 Iout.t160 239.927
R20017 Iout.n988 Iout.t102 239.927
R20018 Iout.n991 Iout.t196 239.927
R20019 Iout.n323 Iout.t212 239.927
R20020 Iout.n326 Iout.t229 239.927
R20021 Iout.n329 Iout.t193 239.927
R20022 Iout.n995 Iout.t57 239.927
R20023 Iout.n1001 Iout.t217 239.927
R20024 Iout.n4 Iout.t218 239.927
R20025 Iout.n295 Iout.t66 239.927
R20026 Iout.n172 Iout.t183 239.927
R20027 Iout.n1014 Iout.t93 239.927
R20028 Iout.n1021 Iout.n1020 7.9105
R20029 Iout.n510 Iout.n509 7.9105
R20030 Iout.n514 Iout.n513 7.9105
R20031 Iout.n508 Iout.n507 7.9105
R20032 Iout.n505 Iout.n504 7.9105
R20033 Iout.n501 Iout.n500 7.9105
R20034 Iout.n193 Iout.n192 7.9105
R20035 Iout.n196 Iout.n195 7.9105
R20036 Iout.n200 Iout.n199 7.9105
R20037 Iout.n203 Iout.n202 7.9105
R20038 Iout.n207 Iout.n206 7.9105
R20039 Iout.n211 Iout.n210 7.9105
R20040 Iout.n215 Iout.n214 7.9105
R20041 Iout.n219 Iout.n218 7.9105
R20042 Iout.n223 Iout.n222 7.9105
R20043 Iout.n227 Iout.n226 7.9105
R20044 Iout.n233 Iout.n232 7.9105
R20045 Iout.n236 Iout.n235 7.9105
R20046 Iout.n239 Iout.n238 7.9105
R20047 Iout.n242 Iout.n241 7.9105
R20048 Iout.n245 Iout.n244 7.9105
R20049 Iout.n248 Iout.n247 7.9105
R20050 Iout.n251 Iout.n250 7.9105
R20051 Iout.n256 Iout.n255 7.9105
R20052 Iout.n253 Iout.n252 7.9105
R20053 Iout.n490 Iout.n489 7.9105
R20054 Iout.n495 Iout.n494 7.9105
R20055 Iout.n492 Iout.n491 7.9105
R20056 Iout.n520 Iout.n519 7.9105
R20057 Iout.n150 Iout.n149 7.9105
R20058 Iout.n147 Iout.n146 7.9105
R20059 Iout.n1011 Iout.n1010 7.9105
R20060 Iout.n1008 Iout.n1007 7.9105
R20061 Iout.n141 Iout.n140 7.9105
R20062 Iout.n144 Iout.n143 7.9105
R20063 Iout.n526 Iout.n525 7.9105
R20064 Iout.n481 Iout.n480 7.9105
R20065 Iout.n484 Iout.n483 7.9105
R20066 Iout.n479 Iout.n478 7.9105
R20067 Iout.n260 Iout.n259 7.9105
R20068 Iout.n187 Iout.n186 7.9105
R20069 Iout.n272 Iout.n271 7.9105
R20070 Iout.n181 Iout.n180 7.9105
R20071 Iout.n284 Iout.n283 7.9105
R20072 Iout.n175 Iout.n174 7.9105
R20073 Iout.n169 Iout.n168 7.9105
R20074 Iout.n302 Iout.n301 7.9105
R20075 Iout.n290 Iout.n289 7.9105
R20076 Iout.n178 Iout.n177 7.9105
R20077 Iout.n278 Iout.n277 7.9105
R20078 Iout.n184 Iout.n183 7.9105
R20079 Iout.n266 Iout.n265 7.9105
R20080 Iout.n190 Iout.n189 7.9105
R20081 Iout.n473 Iout.n472 7.9105
R20082 Iout.n470 Iout.n469 7.9105
R20083 Iout.n157 Iout.n156 7.9105
R20084 Iout.n532 Iout.n531 7.9105
R20085 Iout.n535 Iout.n534 7.9105
R20086 Iout.n537 Iout.n536 7.9105
R20087 Iout.n134 Iout.n133 7.9105
R20088 Iout.n137 Iout.n136 7.9105
R20089 Iout.n543 Iout.n542 7.9105
R20090 Iout.n461 Iout.n460 7.9105
R20091 Iout.n464 Iout.n463 7.9105
R20092 Iout.n459 Iout.n458 7.9105
R20093 Iout.n306 Iout.n305 7.9105
R20094 Iout.n309 Iout.n308 7.9105
R20095 Iout.n312 Iout.n311 7.9105
R20096 Iout.n315 Iout.n314 7.9105
R20097 Iout.n318 Iout.n317 7.9105
R20098 Iout.n321 Iout.n320 7.9105
R20099 Iout.n393 Iout.n392 7.9105
R20100 Iout.n379 Iout.n378 7.9105
R20101 Iout.n377 Iout.n376 7.9105
R20102 Iout.n395 Iout.n394 7.9105
R20103 Iout.n409 Iout.n408 7.9105
R20104 Iout.n411 Iout.n410 7.9105
R20105 Iout.n425 Iout.n424 7.9105
R20106 Iout.n427 Iout.n426 7.9105
R20107 Iout.n448 Iout.n447 7.9105
R20108 Iout.n453 Iout.n452 7.9105
R20109 Iout.n450 Iout.n449 7.9105
R20110 Iout.n549 Iout.n548 7.9105
R20111 Iout.n131 Iout.n130 7.9105
R20112 Iout.n560 Iout.n559 7.9105
R20113 Iout.n558 Iout.n557 7.9105
R20114 Iout.n555 Iout.n554 7.9105
R20115 Iout.n435 Iout.n434 7.9105
R20116 Iout.n439 Iout.n438 7.9105
R20117 Iout.n442 Iout.n441 7.9105
R20118 Iout.n433 Iout.n432 7.9105
R20119 Iout.n419 Iout.n418 7.9105
R20120 Iout.n417 Iout.n416 7.9105
R20121 Iout.n403 Iout.n402 7.9105
R20122 Iout.n358 Iout.n357 7.9105
R20123 Iout.n361 Iout.n360 7.9105
R20124 Iout.n364 Iout.n363 7.9105
R20125 Iout.n367 Iout.n366 7.9105
R20126 Iout.n355 Iout.n354 7.9105
R20127 Iout.n352 Iout.n351 7.9105
R20128 Iout.n349 Iout.n348 7.9105
R20129 Iout.n346 Iout.n345 7.9105
R20130 Iout.n343 Iout.n342 7.9105
R20131 Iout.n340 Iout.n339 7.9105
R20132 Iout.n337 Iout.n336 7.9105
R20133 Iout.n334 Iout.n333 7.9105
R20134 Iout.n118 Iout.n117 7.9105
R20135 Iout.n583 Iout.n582 7.9105
R20136 Iout.n112 Iout.n111 7.9105
R20137 Iout.n595 Iout.n594 7.9105
R20138 Iout.n106 Iout.n105 7.9105
R20139 Iout.n607 Iout.n606 7.9105
R20140 Iout.n100 Iout.n99 7.9105
R20141 Iout.n619 Iout.n618 7.9105
R20142 Iout.n625 Iout.n624 7.9105
R20143 Iout.n91 Iout.n90 7.9105
R20144 Iout.n637 Iout.n636 7.9105
R20145 Iout.n82 Iout.n81 7.9105
R20146 Iout.n649 Iout.n648 7.9105
R20147 Iout.n97 Iout.n96 7.9105
R20148 Iout.n613 Iout.n612 7.9105
R20149 Iout.n103 Iout.n102 7.9105
R20150 Iout.n601 Iout.n600 7.9105
R20151 Iout.n109 Iout.n108 7.9105
R20152 Iout.n589 Iout.n588 7.9105
R20153 Iout.n688 Iout.n687 7.9105
R20154 Iout.n685 Iout.n684 7.9105
R20155 Iout.n682 Iout.n681 7.9105
R20156 Iout.n679 Iout.n678 7.9105
R20157 Iout.n676 Iout.n675 7.9105
R20158 Iout.n673 Iout.n672 7.9105
R20159 Iout.n748 Iout.n747 7.9105
R20160 Iout.n51 Iout.n50 7.9105
R20161 Iout.n760 Iout.n759 7.9105
R20162 Iout.n45 Iout.n44 7.9105
R20163 Iout.n772 Iout.n771 7.9105
R20164 Iout.n43 Iout.n42 7.9105
R20165 Iout.n57 Iout.n56 7.9105
R20166 Iout.n736 Iout.n735 7.9105
R20167 Iout.n63 Iout.n62 7.9105
R20168 Iout.n724 Iout.n723 7.9105
R20169 Iout.n718 Iout.n717 7.9105
R20170 Iout.n66 Iout.n65 7.9105
R20171 Iout.n730 Iout.n729 7.9105
R20172 Iout.n60 Iout.n59 7.9105
R20173 Iout.n806 Iout.n805 7.9105
R20174 Iout.n809 Iout.n808 7.9105
R20175 Iout.n812 Iout.n811 7.9105
R20176 Iout.n815 Iout.n814 7.9105
R20177 Iout.n818 Iout.n817 7.9105
R20178 Iout.n821 Iout.n820 7.9105
R20179 Iout.n824 Iout.n823 7.9105
R20180 Iout.n803 Iout.n802 7.9105
R20181 Iout.n800 Iout.n799 7.9105
R20182 Iout.n891 Iout.n890 7.9105
R20183 Iout.n889 Iout.n888 7.9105
R20184 Iout.n882 Iout.n881 7.9105
R20185 Iout.n870 Iout.n869 7.9105
R20186 Iout.n868 Iout.n867 7.9105
R20187 Iout.n856 Iout.n855 7.9105
R20188 Iout.n854 Iout.n853 7.9105
R20189 Iout.n842 Iout.n841 7.9105
R20190 Iout.n840 Iout.n839 7.9105
R20191 Iout.n828 Iout.n827 7.9105
R20192 Iout.n884 Iout.n883 7.9105
R20193 Iout.n896 Iout.n895 7.9105
R20194 Iout.n898 Iout.n897 7.9105
R20195 Iout.n910 Iout.n909 7.9105
R20196 Iout.n912 Iout.n911 7.9105
R20197 Iout.n924 Iout.n923 7.9105
R20198 Iout.n927 Iout.n926 7.9105
R20199 Iout.n23 Iout.n22 7.9105
R20200 Iout.n877 Iout.n876 7.9105
R20201 Iout.n875 Iout.n874 7.9105
R20202 Iout.n863 Iout.n862 7.9105
R20203 Iout.n861 Iout.n860 7.9105
R20204 Iout.n849 Iout.n848 7.9105
R20205 Iout.n847 Iout.n846 7.9105
R20206 Iout.n835 Iout.n834 7.9105
R20207 Iout.n833 Iout.n832 7.9105
R20208 Iout.n903 Iout.n902 7.9105
R20209 Iout.n905 Iout.n904 7.9105
R20210 Iout.n917 Iout.n916 7.9105
R20211 Iout.n919 Iout.n918 7.9105
R20212 Iout.n932 Iout.n931 7.9105
R20213 Iout.n935 Iout.n934 7.9105
R20214 Iout.n797 Iout.n796 7.9105
R20215 Iout.n794 Iout.n793 7.9105
R20216 Iout.n791 Iout.n790 7.9105
R20217 Iout.n788 Iout.n787 7.9105
R20218 Iout.n785 Iout.n784 7.9105
R20219 Iout.n782 Iout.n781 7.9105
R20220 Iout.n939 Iout.n938 7.9105
R20221 Iout.n742 Iout.n741 7.9105
R20222 Iout.n54 Iout.n53 7.9105
R20223 Iout.n754 Iout.n753 7.9105
R20224 Iout.n48 Iout.n47 7.9105
R20225 Iout.n766 Iout.n765 7.9105
R20226 Iout.n39 Iout.n38 7.9105
R20227 Iout.n778 Iout.n777 7.9105
R20228 Iout.n72 Iout.n71 7.9105
R20229 Iout.n706 Iout.n705 7.9105
R20230 Iout.n78 Iout.n77 7.9105
R20231 Iout.n945 Iout.n944 7.9105
R20232 Iout.n20 Iout.n19 7.9105
R20233 Iout.n69 Iout.n68 7.9105
R20234 Iout.n712 Iout.n711 7.9105
R20235 Iout.n75 Iout.n74 7.9105
R20236 Iout.n700 Iout.n699 7.9105
R20237 Iout.n951 Iout.n950 7.9105
R20238 Iout.n954 Iout.n953 7.9105
R20239 Iout.n670 Iout.n669 7.9105
R20240 Iout.n667 Iout.n666 7.9105
R20241 Iout.n664 Iout.n663 7.9105
R20242 Iout.n661 Iout.n660 7.9105
R20243 Iout.n658 Iout.n657 7.9105
R20244 Iout.n655 Iout.n654 7.9105
R20245 Iout.n691 Iout.n690 7.9105
R20246 Iout.n696 Iout.n695 7.9105
R20247 Iout.n693 Iout.n692 7.9105
R20248 Iout.n958 Iout.n957 7.9105
R20249 Iout.n115 Iout.n114 7.9105
R20250 Iout.n577 Iout.n576 7.9105
R20251 Iout.n574 Iout.n573 7.9105
R20252 Iout.n964 Iout.n963 7.9105
R20253 Iout.n15 Iout.n14 7.9105
R20254 Iout.n94 Iout.n93 7.9105
R20255 Iout.n631 Iout.n630 7.9105
R20256 Iout.n88 Iout.n87 7.9105
R20257 Iout.n643 Iout.n642 7.9105
R20258 Iout.n86 Iout.n85 7.9105
R20259 Iout.n564 Iout.n563 7.9105
R20260 Iout.n970 Iout.n969 7.9105
R20261 Iout.n973 Iout.n972 7.9105
R20262 Iout.n570 Iout.n569 7.9105
R20263 Iout.n124 Iout.n123 7.9105
R20264 Iout.n121 Iout.n120 7.9105
R20265 Iout.n977 Iout.n976 7.9105
R20266 Iout.n401 Iout.n400 7.9105
R20267 Iout.n387 Iout.n386 7.9105
R20268 Iout.n385 Iout.n384 7.9105
R20269 Iout.n371 Iout.n370 7.9105
R20270 Iout.n983 Iout.n982 7.9105
R20271 Iout.n10 Iout.n9 7.9105
R20272 Iout.n128 Iout.n127 7.9105
R20273 Iout.n989 Iout.n988 7.9105
R20274 Iout.n992 Iout.n991 7.9105
R20275 Iout.n324 Iout.n323 7.9105
R20276 Iout.n327 Iout.n326 7.9105
R20277 Iout.n330 Iout.n329 7.9105
R20278 Iout.n996 Iout.n995 7.9105
R20279 Iout.n1002 Iout.n1001 7.9105
R20280 Iout.n5 Iout.n4 7.9105
R20281 Iout.n296 Iout.n295 7.9105
R20282 Iout.n173 Iout.n172 7.9105
R20283 Iout.n1015 Iout.n1014 7.9105
R20284 Iout.n886 Iout.n885 3.86101
R20285 Iout.n880 Iout.n879 3.86101
R20286 Iout.n894 Iout.n893 3.86101
R20287 Iout.n872 Iout.n871 3.86101
R20288 Iout.n900 Iout.n899 3.86101
R20289 Iout.n866 Iout.n865 3.86101
R20290 Iout.n908 Iout.n907 3.86101
R20291 Iout.n858 Iout.n857 3.86101
R20292 Iout.n914 Iout.n913 3.86101
R20293 Iout.n852 Iout.n851 3.86101
R20294 Iout.n922 Iout.n921 3.86101
R20295 Iout.n844 Iout.n843 3.86101
R20296 Iout.n929 Iout.n928 3.86101
R20297 Iout.n838 Iout.n837 3.86101
R20298 Iout.n925 Iout.n21 3.86101
R20299 Iout.n830 Iout.n829 3.86101
R20300 Iout.n879 Iout.n878 3.4105
R20301 Iout.n887 Iout.n886 3.4105
R20302 Iout.n893 Iout.n892 3.4105
R20303 Iout.n798 Iout.n28 3.4105
R20304 Iout.n801 Iout.n29 3.4105
R20305 Iout.n804 Iout.n30 3.4105
R20306 Iout.n807 Iout.n31 3.4105
R20307 Iout.n873 Iout.n872 3.4105
R20308 Iout.n744 Iout.n743 3.4105
R20309 Iout.n740 Iout.n739 3.4105
R20310 Iout.n732 Iout.n731 3.4105
R20311 Iout.n728 Iout.n727 3.4105
R20312 Iout.n720 Iout.n719 3.4105
R20313 Iout.n795 Iout.n27 3.4105
R20314 Iout.n901 Iout.n900 3.4105
R20315 Iout.n722 Iout.n721 3.4105
R20316 Iout.n726 Iout.n725 3.4105
R20317 Iout.n734 Iout.n733 3.4105
R20318 Iout.n738 Iout.n737 3.4105
R20319 Iout.n746 Iout.n745 3.4105
R20320 Iout.n750 Iout.n749 3.4105
R20321 Iout.n752 Iout.n751 3.4105
R20322 Iout.n810 Iout.n32 3.4105
R20323 Iout.n865 Iout.n864 3.4105
R20324 Iout.n668 Iout.n55 3.4105
R20325 Iout.n671 Iout.n58 3.4105
R20326 Iout.n674 Iout.n61 3.4105
R20327 Iout.n677 Iout.n64 3.4105
R20328 Iout.n680 Iout.n67 3.4105
R20329 Iout.n683 Iout.n70 3.4105
R20330 Iout.n686 Iout.n73 3.4105
R20331 Iout.n714 Iout.n713 3.4105
R20332 Iout.n716 Iout.n715 3.4105
R20333 Iout.n792 Iout.n26 3.4105
R20334 Iout.n907 Iout.n906 3.4105
R20335 Iout.n587 Iout.n586 3.4105
R20336 Iout.n591 Iout.n590 3.4105
R20337 Iout.n599 Iout.n598 3.4105
R20338 Iout.n603 Iout.n602 3.4105
R20339 Iout.n611 Iout.n610 3.4105
R20340 Iout.n615 Iout.n614 3.4105
R20341 Iout.n623 Iout.n622 3.4105
R20342 Iout.n627 Iout.n626 3.4105
R20343 Iout.n665 Iout.n52 3.4105
R20344 Iout.n758 Iout.n757 3.4105
R20345 Iout.n756 Iout.n755 3.4105
R20346 Iout.n813 Iout.n33 3.4105
R20347 Iout.n859 Iout.n858 3.4105
R20348 Iout.n629 Iout.n628 3.4105
R20349 Iout.n621 Iout.n620 3.4105
R20350 Iout.n617 Iout.n616 3.4105
R20351 Iout.n609 Iout.n608 3.4105
R20352 Iout.n605 Iout.n604 3.4105
R20353 Iout.n597 Iout.n596 3.4105
R20354 Iout.n593 Iout.n592 3.4105
R20355 Iout.n585 Iout.n584 3.4105
R20356 Iout.n581 Iout.n580 3.4105
R20357 Iout.n579 Iout.n578 3.4105
R20358 Iout.n689 Iout.n76 3.4105
R20359 Iout.n710 Iout.n709 3.4105
R20360 Iout.n708 Iout.n707 3.4105
R20361 Iout.n789 Iout.n25 3.4105
R20362 Iout.n915 Iout.n914 3.4105
R20363 Iout.n572 Iout.n571 3.4105
R20364 Iout.n335 Iout.n116 3.4105
R20365 Iout.n338 Iout.n113 3.4105
R20366 Iout.n341 Iout.n110 3.4105
R20367 Iout.n344 Iout.n107 3.4105
R20368 Iout.n347 Iout.n104 3.4105
R20369 Iout.n350 Iout.n101 3.4105
R20370 Iout.n353 Iout.n98 3.4105
R20371 Iout.n356 Iout.n95 3.4105
R20372 Iout.n359 Iout.n92 3.4105
R20373 Iout.n633 Iout.n632 3.4105
R20374 Iout.n635 Iout.n634 3.4105
R20375 Iout.n662 Iout.n49 3.4105
R20376 Iout.n762 Iout.n761 3.4105
R20377 Iout.n764 Iout.n763 3.4105
R20378 Iout.n816 Iout.n34 3.4105
R20379 Iout.n851 Iout.n850 3.4105
R20380 Iout.n399 Iout.n398 3.4105
R20381 Iout.n405 Iout.n404 3.4105
R20382 Iout.n415 Iout.n414 3.4105
R20383 Iout.n421 Iout.n420 3.4105
R20384 Iout.n431 Iout.n430 3.4105
R20385 Iout.n444 Iout.n443 3.4105
R20386 Iout.n440 Iout.n159 3.4105
R20387 Iout.n437 Iout.n436 3.4105
R20388 Iout.n553 Iout.n552 3.4105
R20389 Iout.n556 Iout.n119 3.4105
R20390 Iout.n562 Iout.n561 3.4105
R20391 Iout.n568 Iout.n567 3.4105
R20392 Iout.n566 Iout.n565 3.4105
R20393 Iout.n575 Iout.n79 3.4105
R20394 Iout.n698 Iout.n697 3.4105
R20395 Iout.n702 Iout.n701 3.4105
R20396 Iout.n704 Iout.n703 3.4105
R20397 Iout.n786 Iout.n24 3.4105
R20398 Iout.n921 Iout.n920 3.4105
R20399 Iout.n129 Iout.n125 3.4105
R20400 Iout.n547 Iout.n546 3.4105
R20401 Iout.n551 Iout.n550 3.4105
R20402 Iout.n451 Iout.n158 3.4105
R20403 Iout.n455 Iout.n454 3.4105
R20404 Iout.n446 Iout.n445 3.4105
R20405 Iout.n429 Iout.n428 3.4105
R20406 Iout.n423 Iout.n422 3.4105
R20407 Iout.n413 Iout.n412 3.4105
R20408 Iout.n407 Iout.n406 3.4105
R20409 Iout.n397 Iout.n396 3.4105
R20410 Iout.n391 Iout.n390 3.4105
R20411 Iout.n389 Iout.n388 3.4105
R20412 Iout.n362 Iout.n89 3.4105
R20413 Iout.n641 Iout.n640 3.4105
R20414 Iout.n639 Iout.n638 3.4105
R20415 Iout.n659 Iout.n46 3.4105
R20416 Iout.n770 Iout.n769 3.4105
R20417 Iout.n768 Iout.n767 3.4105
R20418 Iout.n819 Iout.n35 3.4105
R20419 Iout.n845 Iout.n844 3.4105
R20420 Iout.n325 Iout.n165 3.4105
R20421 Iout.n322 Iout.n164 3.4105
R20422 Iout.n319 Iout.n163 3.4105
R20423 Iout.n316 Iout.n162 3.4105
R20424 Iout.n313 Iout.n161 3.4105
R20425 Iout.n310 Iout.n160 3.4105
R20426 Iout.n307 Iout.n155 3.4105
R20427 Iout.n457 Iout.n456 3.4105
R20428 Iout.n466 Iout.n465 3.4105
R20429 Iout.n462 Iout.n126 3.4105
R20430 Iout.n545 Iout.n544 3.4105
R20431 Iout.n541 Iout.n540 3.4105
R20432 Iout.n135 Iout.n3 3.4105
R20433 Iout.n987 Iout.n986 3.4105
R20434 Iout.n985 Iout.n984 3.4105
R20435 Iout.n122 Iout.n8 3.4105
R20436 Iout.n968 Iout.n967 3.4105
R20437 Iout.n966 Iout.n965 3.4105
R20438 Iout.n694 Iout.n13 3.4105
R20439 Iout.n949 Iout.n948 3.4105
R20440 Iout.n947 Iout.n946 3.4105
R20441 Iout.n783 Iout.n18 3.4105
R20442 Iout.n930 Iout.n929 3.4105
R20443 Iout.n1004 Iout.n1003 3.4105
R20444 Iout.n539 Iout.n538 3.4105
R20445 Iout.n533 Iout.n132 3.4105
R20446 Iout.n530 Iout.n529 3.4105
R20447 Iout.n468 Iout.n467 3.4105
R20448 Iout.n471 Iout.n153 3.4105
R20449 Iout.n475 Iout.n474 3.4105
R20450 Iout.n264 Iout.n263 3.4105
R20451 Iout.n268 Iout.n267 3.4105
R20452 Iout.n276 Iout.n275 3.4105
R20453 Iout.n280 Iout.n279 3.4105
R20454 Iout.n288 Iout.n287 3.4105
R20455 Iout.n292 Iout.n291 3.4105
R20456 Iout.n300 Iout.n299 3.4105
R20457 Iout.n328 Iout.n166 3.4105
R20458 Iout.n381 Iout.n380 3.4105
R20459 Iout.n383 Iout.n382 3.4105
R20460 Iout.n365 Iout.n83 3.4105
R20461 Iout.n645 Iout.n644 3.4105
R20462 Iout.n647 Iout.n646 3.4105
R20463 Iout.n656 Iout.n40 3.4105
R20464 Iout.n774 Iout.n773 3.4105
R20465 Iout.n776 Iout.n775 3.4105
R20466 Iout.n822 Iout.n36 3.4105
R20467 Iout.n837 Iout.n836 3.4105
R20468 Iout.n298 Iout.n297 3.4105
R20469 Iout.n294 Iout.n293 3.4105
R20470 Iout.n286 Iout.n285 3.4105
R20471 Iout.n282 Iout.n281 3.4105
R20472 Iout.n274 Iout.n273 3.4105
R20473 Iout.n270 Iout.n269 3.4105
R20474 Iout.n262 Iout.n261 3.4105
R20475 Iout.n477 Iout.n476 3.4105
R20476 Iout.n486 Iout.n485 3.4105
R20477 Iout.n482 Iout.n151 3.4105
R20478 Iout.n528 Iout.n527 3.4105
R20479 Iout.n524 Iout.n523 3.4105
R20480 Iout.n142 Iout.n138 3.4105
R20481 Iout.n1006 Iout.n1005 3.4105
R20482 Iout.n1009 Iout.n0 3.4105
R20483 Iout.n1000 Iout.n999 3.4105
R20484 Iout.n998 Iout.n997 3.4105
R20485 Iout.n990 Iout.n6 3.4105
R20486 Iout.n981 Iout.n980 3.4105
R20487 Iout.n979 Iout.n978 3.4105
R20488 Iout.n971 Iout.n11 3.4105
R20489 Iout.n962 Iout.n961 3.4105
R20490 Iout.n960 Iout.n959 3.4105
R20491 Iout.n952 Iout.n16 3.4105
R20492 Iout.n943 Iout.n942 3.4105
R20493 Iout.n941 Iout.n940 3.4105
R20494 Iout.n933 Iout.n21 3.4105
R20495 Iout.n1017 Iout.n1016 3.4105
R20496 Iout.n148 Iout.n2 3.4105
R20497 Iout.n518 Iout.n517 3.4105
R20498 Iout.n522 Iout.n521 3.4105
R20499 Iout.n493 Iout.n139 3.4105
R20500 Iout.n497 Iout.n496 3.4105
R20501 Iout.n488 Iout.n487 3.4105
R20502 Iout.n254 Iout.n154 3.4105
R20503 Iout.n258 Iout.n257 3.4105
R20504 Iout.n249 Iout.n188 3.4105
R20505 Iout.n246 Iout.n185 3.4105
R20506 Iout.n243 Iout.n182 3.4105
R20507 Iout.n240 Iout.n179 3.4105
R20508 Iout.n237 Iout.n176 3.4105
R20509 Iout.n234 Iout.n170 3.4105
R20510 Iout.n231 Iout.n230 3.4105
R20511 Iout.n171 Iout.n167 3.4105
R20512 Iout.n304 Iout.n303 3.4105
R20513 Iout.n332 Iout.n331 3.4105
R20514 Iout.n375 Iout.n374 3.4105
R20515 Iout.n373 Iout.n372 3.4105
R20516 Iout.n369 Iout.n368 3.4105
R20517 Iout.n84 Iout.n80 3.4105
R20518 Iout.n651 Iout.n650 3.4105
R20519 Iout.n653 Iout.n652 3.4105
R20520 Iout.n41 Iout.n37 3.4105
R20521 Iout.n780 Iout.n779 3.4105
R20522 Iout.n826 Iout.n825 3.4105
R20523 Iout.n831 Iout.n830 3.4105
R20524 Iout.n229 Iout.n228 3.4105
R20525 Iout.n225 Iout.n224 3.4105
R20526 Iout.n221 Iout.n220 3.4105
R20527 Iout.n217 Iout.n216 3.4105
R20528 Iout.n213 Iout.n212 3.4105
R20529 Iout.n209 Iout.n208 3.4105
R20530 Iout.n205 Iout.n204 3.4105
R20531 Iout.n201 Iout.n191 3.4105
R20532 Iout.n198 Iout.n197 3.4105
R20533 Iout.n194 Iout.n152 3.4105
R20534 Iout.n499 Iout.n498 3.4105
R20535 Iout.n503 Iout.n502 3.4105
R20536 Iout.n506 Iout.n145 3.4105
R20537 Iout.n516 Iout.n515 3.4105
R20538 Iout.n512 Iout.n511 3.4105
R20539 Iout.n1019 Iout.n1018 3.4105
R20540 Iout.n936 Iout.n23 1.43848
R20541 Iout.n936 Iout.n935 1.34612
R20542 Iout.n939 Iout.n937 1.34612
R20543 Iout.n20 Iout.n17 1.34612
R20544 Iout.n955 Iout.n954 1.34612
R20545 Iout.n958 Iout.n956 1.34612
R20546 Iout.n15 Iout.n12 1.34612
R20547 Iout.n974 Iout.n973 1.34612
R20548 Iout.n977 Iout.n975 1.34612
R20549 Iout.n10 Iout.n7 1.34612
R20550 Iout.n993 Iout.n992 1.34612
R20551 Iout.n996 Iout.n994 1.34612
R20552 Iout.n5 Iout.n1 1.34612
R20553 Iout.n1012 Iout.n1011 1.34612
R20554 Iout.n1015 Iout.n1013 1.34612
R20555 Iout.n1022 Iout.n1021 1.34612
R20556 Iout.n197 Iout.n154 0.451012
R20557 Iout.n476 Iout.n154 0.451012
R20558 Iout.n476 Iout.n475 0.451012
R20559 Iout.n475 Iout.n155 0.451012
R20560 Iout.n445 Iout.n155 0.451012
R20561 Iout.n445 Iout.n444 0.451012
R20562 Iout.n444 Iout.n107 0.451012
R20563 Iout.n604 Iout.n107 0.451012
R20564 Iout.n604 Iout.n603 0.451012
R20565 Iout.n603 Iout.n64 0.451012
R20566 Iout.n733 Iout.n64 0.451012
R20567 Iout.n733 Iout.n732 0.451012
R20568 Iout.n732 Iout.n29 0.451012
R20569 Iout.n886 Iout.n29 0.451012
R20570 Iout.n258 Iout.n191 0.451012
R20571 Iout.n262 Iout.n258 0.451012
R20572 Iout.n263 Iout.n262 0.451012
R20573 Iout.n263 Iout.n160 0.451012
R20574 Iout.n429 Iout.n160 0.451012
R20575 Iout.n430 Iout.n429 0.451012
R20576 Iout.n430 Iout.n104 0.451012
R20577 Iout.n609 Iout.n104 0.451012
R20578 Iout.n610 Iout.n609 0.451012
R20579 Iout.n610 Iout.n61 0.451012
R20580 Iout.n738 Iout.n61 0.451012
R20581 Iout.n739 Iout.n738 0.451012
R20582 Iout.n739 Iout.n30 0.451012
R20583 Iout.n879 Iout.n30 0.451012
R20584 Iout.n487 Iout.n152 0.451012
R20585 Iout.n487 Iout.n486 0.451012
R20586 Iout.n486 Iout.n153 0.451012
R20587 Iout.n456 Iout.n153 0.451012
R20588 Iout.n456 Iout.n455 0.451012
R20589 Iout.n455 Iout.n159 0.451012
R20590 Iout.n159 Iout.n110 0.451012
R20591 Iout.n597 Iout.n110 0.451012
R20592 Iout.n598 Iout.n597 0.451012
R20593 Iout.n598 Iout.n67 0.451012
R20594 Iout.n726 Iout.n67 0.451012
R20595 Iout.n727 Iout.n726 0.451012
R20596 Iout.n727 Iout.n28 0.451012
R20597 Iout.n893 Iout.n28 0.451012
R20598 Iout.n204 Iout.n188 0.451012
R20599 Iout.n269 Iout.n188 0.451012
R20600 Iout.n269 Iout.n268 0.451012
R20601 Iout.n268 Iout.n161 0.451012
R20602 Iout.n422 Iout.n161 0.451012
R20603 Iout.n422 Iout.n421 0.451012
R20604 Iout.n421 Iout.n101 0.451012
R20605 Iout.n616 Iout.n101 0.451012
R20606 Iout.n616 Iout.n615 0.451012
R20607 Iout.n615 Iout.n58 0.451012
R20608 Iout.n745 Iout.n58 0.451012
R20609 Iout.n745 Iout.n744 0.451012
R20610 Iout.n744 Iout.n31 0.451012
R20611 Iout.n872 Iout.n31 0.451012
R20612 Iout.n498 Iout.n497 0.451012
R20613 Iout.n497 Iout.n151 0.451012
R20614 Iout.n467 Iout.n151 0.451012
R20615 Iout.n467 Iout.n466 0.451012
R20616 Iout.n466 Iout.n158 0.451012
R20617 Iout.n436 Iout.n158 0.451012
R20618 Iout.n436 Iout.n113 0.451012
R20619 Iout.n592 Iout.n113 0.451012
R20620 Iout.n592 Iout.n591 0.451012
R20621 Iout.n591 Iout.n70 0.451012
R20622 Iout.n721 Iout.n70 0.451012
R20623 Iout.n721 Iout.n720 0.451012
R20624 Iout.n720 Iout.n27 0.451012
R20625 Iout.n900 Iout.n27 0.451012
R20626 Iout.n208 Iout.n185 0.451012
R20627 Iout.n274 Iout.n185 0.451012
R20628 Iout.n275 Iout.n274 0.451012
R20629 Iout.n275 Iout.n162 0.451012
R20630 Iout.n413 Iout.n162 0.451012
R20631 Iout.n414 Iout.n413 0.451012
R20632 Iout.n414 Iout.n98 0.451012
R20633 Iout.n621 Iout.n98 0.451012
R20634 Iout.n622 Iout.n621 0.451012
R20635 Iout.n622 Iout.n55 0.451012
R20636 Iout.n750 Iout.n55 0.451012
R20637 Iout.n751 Iout.n750 0.451012
R20638 Iout.n751 Iout.n32 0.451012
R20639 Iout.n865 Iout.n32 0.451012
R20640 Iout.n502 Iout.n139 0.451012
R20641 Iout.n528 Iout.n139 0.451012
R20642 Iout.n529 Iout.n528 0.451012
R20643 Iout.n529 Iout.n126 0.451012
R20644 Iout.n551 Iout.n126 0.451012
R20645 Iout.n552 Iout.n551 0.451012
R20646 Iout.n552 Iout.n116 0.451012
R20647 Iout.n585 Iout.n116 0.451012
R20648 Iout.n586 Iout.n585 0.451012
R20649 Iout.n586 Iout.n73 0.451012
R20650 Iout.n714 Iout.n73 0.451012
R20651 Iout.n715 Iout.n714 0.451012
R20652 Iout.n715 Iout.n26 0.451012
R20653 Iout.n907 Iout.n26 0.451012
R20654 Iout.n212 Iout.n182 0.451012
R20655 Iout.n281 Iout.n182 0.451012
R20656 Iout.n281 Iout.n280 0.451012
R20657 Iout.n280 Iout.n163 0.451012
R20658 Iout.n406 Iout.n163 0.451012
R20659 Iout.n406 Iout.n405 0.451012
R20660 Iout.n405 Iout.n95 0.451012
R20661 Iout.n628 Iout.n95 0.451012
R20662 Iout.n628 Iout.n627 0.451012
R20663 Iout.n627 Iout.n52 0.451012
R20664 Iout.n757 Iout.n52 0.451012
R20665 Iout.n757 Iout.n756 0.451012
R20666 Iout.n756 Iout.n33 0.451012
R20667 Iout.n858 Iout.n33 0.451012
R20668 Iout.n522 Iout.n145 0.451012
R20669 Iout.n523 Iout.n522 0.451012
R20670 Iout.n523 Iout.n132 0.451012
R20671 Iout.n545 Iout.n132 0.451012
R20672 Iout.n546 Iout.n545 0.451012
R20673 Iout.n546 Iout.n119 0.451012
R20674 Iout.n572 Iout.n119 0.451012
R20675 Iout.n580 Iout.n572 0.451012
R20676 Iout.n580 Iout.n579 0.451012
R20677 Iout.n579 Iout.n76 0.451012
R20678 Iout.n709 Iout.n76 0.451012
R20679 Iout.n709 Iout.n708 0.451012
R20680 Iout.n708 Iout.n25 0.451012
R20681 Iout.n914 Iout.n25 0.451012
R20682 Iout.n216 Iout.n179 0.451012
R20683 Iout.n286 Iout.n179 0.451012
R20684 Iout.n287 Iout.n286 0.451012
R20685 Iout.n287 Iout.n164 0.451012
R20686 Iout.n397 Iout.n164 0.451012
R20687 Iout.n398 Iout.n397 0.451012
R20688 Iout.n398 Iout.n92 0.451012
R20689 Iout.n633 Iout.n92 0.451012
R20690 Iout.n634 Iout.n633 0.451012
R20691 Iout.n634 Iout.n49 0.451012
R20692 Iout.n762 Iout.n49 0.451012
R20693 Iout.n763 Iout.n762 0.451012
R20694 Iout.n763 Iout.n34 0.451012
R20695 Iout.n851 Iout.n34 0.451012
R20696 Iout.n517 Iout.n516 0.451012
R20697 Iout.n517 Iout.n138 0.451012
R20698 Iout.n539 Iout.n138 0.451012
R20699 Iout.n540 Iout.n539 0.451012
R20700 Iout.n540 Iout.n125 0.451012
R20701 Iout.n562 Iout.n125 0.451012
R20702 Iout.n567 Iout.n562 0.451012
R20703 Iout.n567 Iout.n566 0.451012
R20704 Iout.n566 Iout.n79 0.451012
R20705 Iout.n698 Iout.n79 0.451012
R20706 Iout.n702 Iout.n698 0.451012
R20707 Iout.n703 Iout.n702 0.451012
R20708 Iout.n703 Iout.n24 0.451012
R20709 Iout.n921 Iout.n24 0.451012
R20710 Iout.n220 Iout.n176 0.451012
R20711 Iout.n293 Iout.n176 0.451012
R20712 Iout.n293 Iout.n292 0.451012
R20713 Iout.n292 Iout.n165 0.451012
R20714 Iout.n390 Iout.n165 0.451012
R20715 Iout.n390 Iout.n389 0.451012
R20716 Iout.n389 Iout.n89 0.451012
R20717 Iout.n640 Iout.n89 0.451012
R20718 Iout.n640 Iout.n639 0.451012
R20719 Iout.n639 Iout.n46 0.451012
R20720 Iout.n769 Iout.n46 0.451012
R20721 Iout.n769 Iout.n768 0.451012
R20722 Iout.n768 Iout.n35 0.451012
R20723 Iout.n844 Iout.n35 0.451012
R20724 Iout.n511 Iout.n2 0.451012
R20725 Iout.n1005 Iout.n2 0.451012
R20726 Iout.n1005 Iout.n1004 0.451012
R20727 Iout.n1004 Iout.n3 0.451012
R20728 Iout.n986 Iout.n3 0.451012
R20729 Iout.n986 Iout.n985 0.451012
R20730 Iout.n985 Iout.n8 0.451012
R20731 Iout.n967 Iout.n8 0.451012
R20732 Iout.n967 Iout.n966 0.451012
R20733 Iout.n966 Iout.n13 0.451012
R20734 Iout.n948 Iout.n13 0.451012
R20735 Iout.n948 Iout.n947 0.451012
R20736 Iout.n947 Iout.n18 0.451012
R20737 Iout.n929 Iout.n18 0.451012
R20738 Iout.n224 Iout.n170 0.451012
R20739 Iout.n298 Iout.n170 0.451012
R20740 Iout.n299 Iout.n298 0.451012
R20741 Iout.n299 Iout.n166 0.451012
R20742 Iout.n381 Iout.n166 0.451012
R20743 Iout.n382 Iout.n381 0.451012
R20744 Iout.n382 Iout.n83 0.451012
R20745 Iout.n645 Iout.n83 0.451012
R20746 Iout.n646 Iout.n645 0.451012
R20747 Iout.n646 Iout.n40 0.451012
R20748 Iout.n774 Iout.n40 0.451012
R20749 Iout.n775 Iout.n774 0.451012
R20750 Iout.n775 Iout.n36 0.451012
R20751 Iout.n837 Iout.n36 0.451012
R20752 Iout.n1018 Iout.n1017 0.451012
R20753 Iout.n1017 Iout.n0 0.451012
R20754 Iout.n999 Iout.n0 0.451012
R20755 Iout.n999 Iout.n998 0.451012
R20756 Iout.n998 Iout.n6 0.451012
R20757 Iout.n980 Iout.n6 0.451012
R20758 Iout.n980 Iout.n979 0.451012
R20759 Iout.n979 Iout.n11 0.451012
R20760 Iout.n961 Iout.n11 0.451012
R20761 Iout.n961 Iout.n960 0.451012
R20762 Iout.n960 Iout.n16 0.451012
R20763 Iout.n942 Iout.n16 0.451012
R20764 Iout.n942 Iout.n941 0.451012
R20765 Iout.n941 Iout.n21 0.451012
R20766 Iout.n230 Iout.n229 0.451012
R20767 Iout.n230 Iout.n167 0.451012
R20768 Iout.n304 Iout.n167 0.451012
R20769 Iout.n332 Iout.n304 0.451012
R20770 Iout.n374 Iout.n332 0.451012
R20771 Iout.n374 Iout.n373 0.451012
R20772 Iout.n373 Iout.n369 0.451012
R20773 Iout.n369 Iout.n80 0.451012
R20774 Iout.n651 Iout.n80 0.451012
R20775 Iout.n652 Iout.n651 0.451012
R20776 Iout.n652 Iout.n37 0.451012
R20777 Iout.n780 Iout.n37 0.451012
R20778 Iout.n826 Iout.n780 0.451012
R20779 Iout.n830 Iout.n826 0.451012
R20780 Iout.n231 Iout 0.2919
R20781 Iout.n303 Iout 0.2919
R20782 Iout Iout.n300 0.2919
R20783 Iout.n375 Iout 0.2919
R20784 Iout.n380 Iout 0.2919
R20785 Iout.n391 Iout 0.2919
R20786 Iout.n368 Iout 0.2919
R20787 Iout Iout.n365 0.2919
R20788 Iout Iout.n362 0.2919
R20789 Iout Iout.n359 0.2919
R20790 Iout.n650 Iout 0.2919
R20791 Iout Iout.n647 0.2919
R20792 Iout.n638 Iout 0.2919
R20793 Iout Iout.n635 0.2919
R20794 Iout.n626 Iout 0.2919
R20795 Iout.n41 Iout 0.2919
R20796 Iout.n773 Iout 0.2919
R20797 Iout Iout.n770 0.2919
R20798 Iout.n761 Iout 0.2919
R20799 Iout Iout.n758 0.2919
R20800 Iout.n749 Iout 0.2919
R20801 Iout.n825 Iout 0.2919
R20802 Iout Iout.n822 0.2919
R20803 Iout Iout.n819 0.2919
R20804 Iout Iout.n816 0.2919
R20805 Iout Iout.n813 0.2919
R20806 Iout Iout.n810 0.2919
R20807 Iout Iout.n807 0.2919
R20808 Iout.n829 Iout 0.2919
R20809 Iout.n838 Iout 0.2919
R20810 Iout.n843 Iout 0.2919
R20811 Iout.n852 Iout 0.2919
R20812 Iout.n857 Iout 0.2919
R20813 Iout.n866 Iout 0.2919
R20814 Iout.n871 Iout 0.2919
R20815 Iout.n880 Iout 0.2919
R20816 Iout Iout.n925 0.2919
R20817 Iout.n928 Iout 0.2919
R20818 Iout.n922 Iout 0.2919
R20819 Iout.n913 Iout 0.2919
R20820 Iout.n908 Iout 0.2919
R20821 Iout.n899 Iout 0.2919
R20822 Iout.n894 Iout 0.2919
R20823 Iout.n885 Iout 0.2919
R20824 Iout.n831 Iout 0.2919
R20825 Iout.n836 Iout 0.2919
R20826 Iout.n845 Iout 0.2919
R20827 Iout.n850 Iout 0.2919
R20828 Iout.n859 Iout 0.2919
R20829 Iout.n864 Iout 0.2919
R20830 Iout.n873 Iout 0.2919
R20831 Iout.n878 Iout 0.2919
R20832 Iout.n887 Iout 0.2919
R20833 Iout.n892 Iout 0.2919
R20834 Iout.n933 Iout 0.2919
R20835 Iout.n930 Iout 0.2919
R20836 Iout.n920 Iout 0.2919
R20837 Iout.n915 Iout 0.2919
R20838 Iout.n906 Iout 0.2919
R20839 Iout.n901 Iout 0.2919
R20840 Iout.n940 Iout 0.2919
R20841 Iout Iout.n783 0.2919
R20842 Iout Iout.n786 0.2919
R20843 Iout Iout.n789 0.2919
R20844 Iout Iout.n792 0.2919
R20845 Iout Iout.n795 0.2919
R20846 Iout Iout.n798 0.2919
R20847 Iout Iout.n801 0.2919
R20848 Iout Iout.n804 0.2919
R20849 Iout.n779 Iout 0.2919
R20850 Iout Iout.n776 0.2919
R20851 Iout.n767 Iout 0.2919
R20852 Iout Iout.n764 0.2919
R20853 Iout.n755 Iout 0.2919
R20854 Iout Iout.n752 0.2919
R20855 Iout.n743 Iout 0.2919
R20856 Iout Iout.n740 0.2919
R20857 Iout.n731 Iout 0.2919
R20858 Iout Iout.n728 0.2919
R20859 Iout.n719 Iout 0.2919
R20860 Iout Iout.n943 0.2919
R20861 Iout.n946 Iout 0.2919
R20862 Iout Iout.n704 0.2919
R20863 Iout.n707 Iout 0.2919
R20864 Iout Iout.n716 0.2919
R20865 Iout.n952 Iout 0.2919
R20866 Iout.n949 Iout 0.2919
R20867 Iout.n701 Iout 0.2919
R20868 Iout Iout.n710 0.2919
R20869 Iout.n713 Iout 0.2919
R20870 Iout Iout.n722 0.2919
R20871 Iout.n725 Iout 0.2919
R20872 Iout Iout.n734 0.2919
R20873 Iout.n737 Iout 0.2919
R20874 Iout Iout.n746 0.2919
R20875 Iout.n653 Iout 0.2919
R20876 Iout.n656 Iout 0.2919
R20877 Iout.n659 Iout 0.2919
R20878 Iout.n662 Iout 0.2919
R20879 Iout.n665 Iout 0.2919
R20880 Iout.n668 Iout 0.2919
R20881 Iout.n671 Iout 0.2919
R20882 Iout.n674 Iout 0.2919
R20883 Iout.n677 Iout 0.2919
R20884 Iout.n680 Iout 0.2919
R20885 Iout.n683 Iout 0.2919
R20886 Iout.n686 Iout 0.2919
R20887 Iout.n959 Iout 0.2919
R20888 Iout Iout.n694 0.2919
R20889 Iout.n697 Iout 0.2919
R20890 Iout.n689 Iout 0.2919
R20891 Iout Iout.n962 0.2919
R20892 Iout.n965 Iout 0.2919
R20893 Iout Iout.n575 0.2919
R20894 Iout.n578 Iout 0.2919
R20895 Iout Iout.n587 0.2919
R20896 Iout.n590 Iout 0.2919
R20897 Iout Iout.n599 0.2919
R20898 Iout.n602 Iout 0.2919
R20899 Iout Iout.n611 0.2919
R20900 Iout.n614 Iout 0.2919
R20901 Iout Iout.n623 0.2919
R20902 Iout.n84 Iout 0.2919
R20903 Iout.n644 Iout 0.2919
R20904 Iout Iout.n641 0.2919
R20905 Iout.n632 Iout 0.2919
R20906 Iout Iout.n629 0.2919
R20907 Iout.n620 Iout 0.2919
R20908 Iout Iout.n617 0.2919
R20909 Iout.n608 Iout 0.2919
R20910 Iout Iout.n605 0.2919
R20911 Iout.n596 Iout 0.2919
R20912 Iout Iout.n593 0.2919
R20913 Iout.n584 Iout 0.2919
R20914 Iout Iout.n581 0.2919
R20915 Iout.n971 Iout 0.2919
R20916 Iout.n968 Iout 0.2919
R20917 Iout.n565 Iout 0.2919
R20918 Iout.n978 Iout 0.2919
R20919 Iout Iout.n122 0.2919
R20920 Iout Iout.n568 0.2919
R20921 Iout.n571 Iout 0.2919
R20922 Iout Iout.n335 0.2919
R20923 Iout Iout.n338 0.2919
R20924 Iout Iout.n341 0.2919
R20925 Iout Iout.n344 0.2919
R20926 Iout Iout.n347 0.2919
R20927 Iout Iout.n350 0.2919
R20928 Iout Iout.n353 0.2919
R20929 Iout Iout.n356 0.2919
R20930 Iout.n372 Iout 0.2919
R20931 Iout.n383 Iout 0.2919
R20932 Iout.n388 Iout 0.2919
R20933 Iout.n399 Iout 0.2919
R20934 Iout.n404 Iout 0.2919
R20935 Iout.n415 Iout 0.2919
R20936 Iout.n420 Iout 0.2919
R20937 Iout.n431 Iout 0.2919
R20938 Iout.n443 Iout 0.2919
R20939 Iout Iout.n440 0.2919
R20940 Iout Iout.n437 0.2919
R20941 Iout.n553 Iout 0.2919
R20942 Iout.n556 Iout 0.2919
R20943 Iout.n561 Iout 0.2919
R20944 Iout Iout.n981 0.2919
R20945 Iout.n984 Iout 0.2919
R20946 Iout.n990 Iout 0.2919
R20947 Iout.n987 Iout 0.2919
R20948 Iout Iout.n129 0.2919
R20949 Iout Iout.n547 0.2919
R20950 Iout.n550 Iout 0.2919
R20951 Iout Iout.n451 0.2919
R20952 Iout.n454 Iout 0.2919
R20953 Iout.n446 Iout 0.2919
R20954 Iout.n428 Iout 0.2919
R20955 Iout.n423 Iout 0.2919
R20956 Iout.n412 Iout 0.2919
R20957 Iout.n407 Iout 0.2919
R20958 Iout.n396 Iout 0.2919
R20959 Iout.n331 Iout 0.2919
R20960 Iout Iout.n328 0.2919
R20961 Iout Iout.n325 0.2919
R20962 Iout Iout.n322 0.2919
R20963 Iout Iout.n319 0.2919
R20964 Iout Iout.n316 0.2919
R20965 Iout Iout.n313 0.2919
R20966 Iout Iout.n310 0.2919
R20967 Iout Iout.n307 0.2919
R20968 Iout.n457 Iout 0.2919
R20969 Iout.n465 Iout 0.2919
R20970 Iout Iout.n462 0.2919
R20971 Iout.n544 Iout 0.2919
R20972 Iout Iout.n541 0.2919
R20973 Iout Iout.n135 0.2919
R20974 Iout.n997 Iout 0.2919
R20975 Iout Iout.n1000 0.2919
R20976 Iout.n1003 Iout 0.2919
R20977 Iout.n538 Iout 0.2919
R20978 Iout.n533 Iout 0.2919
R20979 Iout.n530 Iout 0.2919
R20980 Iout Iout.n468 0.2919
R20981 Iout Iout.n471 0.2919
R20982 Iout.n474 Iout 0.2919
R20983 Iout Iout.n264 0.2919
R20984 Iout.n267 Iout 0.2919
R20985 Iout Iout.n276 0.2919
R20986 Iout.n279 Iout 0.2919
R20987 Iout Iout.n288 0.2919
R20988 Iout.n291 Iout 0.2919
R20989 Iout.n171 Iout 0.2919
R20990 Iout.n297 Iout 0.2919
R20991 Iout Iout.n294 0.2919
R20992 Iout.n285 Iout 0.2919
R20993 Iout Iout.n282 0.2919
R20994 Iout.n273 Iout 0.2919
R20995 Iout Iout.n270 0.2919
R20996 Iout.n261 Iout 0.2919
R20997 Iout.n477 Iout 0.2919
R20998 Iout.n485 Iout 0.2919
R20999 Iout Iout.n482 0.2919
R21000 Iout.n527 Iout 0.2919
R21001 Iout Iout.n524 0.2919
R21002 Iout Iout.n142 0.2919
R21003 Iout.n1006 Iout 0.2919
R21004 Iout.n1009 Iout 0.2919
R21005 Iout.n1016 Iout 0.2919
R21006 Iout Iout.n148 0.2919
R21007 Iout Iout.n518 0.2919
R21008 Iout.n521 Iout 0.2919
R21009 Iout Iout.n493 0.2919
R21010 Iout.n496 Iout 0.2919
R21011 Iout.n488 Iout 0.2919
R21012 Iout Iout.n254 0.2919
R21013 Iout.n257 Iout 0.2919
R21014 Iout.n249 Iout 0.2919
R21015 Iout.n246 Iout 0.2919
R21016 Iout.n243 Iout 0.2919
R21017 Iout.n240 Iout 0.2919
R21018 Iout.n237 Iout 0.2919
R21019 Iout.n234 Iout 0.2919
R21020 Iout.n228 Iout 0.2919
R21021 Iout Iout.n225 0.2919
R21022 Iout Iout.n221 0.2919
R21023 Iout Iout.n217 0.2919
R21024 Iout Iout.n213 0.2919
R21025 Iout Iout.n209 0.2919
R21026 Iout Iout.n205 0.2919
R21027 Iout Iout.n201 0.2919
R21028 Iout Iout.n198 0.2919
R21029 Iout Iout.n194 0.2919
R21030 Iout.n499 Iout 0.2919
R21031 Iout.n503 Iout 0.2919
R21032 Iout.n506 Iout 0.2919
R21033 Iout.n515 Iout 0.2919
R21034 Iout Iout.n512 0.2919
R21035 Iout.n1019 Iout 0.2919
R21036 Iout.n1013 Iout.n1012 0.092855
R21037 Iout.n1012 Iout.n1 0.092855
R21038 Iout.n994 Iout.n1 0.092855
R21039 Iout.n994 Iout.n993 0.092855
R21040 Iout.n993 Iout.n7 0.092855
R21041 Iout.n975 Iout.n7 0.092855
R21042 Iout.n975 Iout.n974 0.092855
R21043 Iout.n974 Iout.n12 0.092855
R21044 Iout.n956 Iout.n12 0.092855
R21045 Iout.n956 Iout.n955 0.092855
R21046 Iout.n955 Iout.n17 0.092855
R21047 Iout.n937 Iout.n17 0.092855
R21048 Iout.n937 Iout.n936 0.092855
R21049 Iout.n197 Iout 0.0818902
R21050 Iout.n191 Iout 0.0818902
R21051 Iout.n152 Iout 0.0818902
R21052 Iout.n204 Iout 0.0818902
R21053 Iout.n498 Iout 0.0818902
R21054 Iout.n208 Iout 0.0818902
R21055 Iout.n502 Iout 0.0818902
R21056 Iout.n212 Iout 0.0818902
R21057 Iout.n145 Iout 0.0818902
R21058 Iout.n216 Iout 0.0818902
R21059 Iout.n516 Iout 0.0818902
R21060 Iout.n220 Iout 0.0818902
R21061 Iout.n511 Iout 0.0818902
R21062 Iout.n224 Iout 0.0818902
R21063 Iout.n1018 Iout 0.0818902
R21064 Iout.n229 Iout 0.0818902
R21065 Iout.n1013 Iout 0.072645
R21066 Iout.n302 Iout 0.0532071
R21067 Iout Iout.n377 0.0532071
R21068 Iout.n379 Iout 0.0532071
R21069 Iout.n367 Iout 0.0532071
R21070 Iout.n364 Iout 0.0532071
R21071 Iout.n361 Iout 0.0532071
R21072 Iout.n649 Iout 0.0532071
R21073 Iout Iout.n82 0.0532071
R21074 Iout.n637 Iout 0.0532071
R21075 Iout Iout.n91 0.0532071
R21076 Iout Iout.n43 0.0532071
R21077 Iout.n772 Iout 0.0532071
R21078 Iout Iout.n45 0.0532071
R21079 Iout.n760 Iout 0.0532071
R21080 Iout Iout.n51 0.0532071
R21081 Iout.n824 Iout 0.0532071
R21082 Iout.n821 Iout 0.0532071
R21083 Iout.n818 Iout 0.0532071
R21084 Iout.n815 Iout 0.0532071
R21085 Iout.n812 Iout 0.0532071
R21086 Iout.n809 Iout 0.0532071
R21087 Iout.n828 Iout 0.0532071
R21088 Iout Iout.n840 0.0532071
R21089 Iout.n842 Iout 0.0532071
R21090 Iout Iout.n854 0.0532071
R21091 Iout.n856 Iout 0.0532071
R21092 Iout Iout.n868 0.0532071
R21093 Iout.n870 Iout 0.0532071
R21094 Iout.n927 Iout 0.0532071
R21095 Iout Iout.n924 0.0532071
R21096 Iout.n912 Iout 0.0532071
R21097 Iout Iout.n910 0.0532071
R21098 Iout.n898 Iout 0.0532071
R21099 Iout Iout.n896 0.0532071
R21100 Iout.n884 Iout 0.0532071
R21101 Iout Iout.n882 0.0532071
R21102 Iout Iout.n833 0.0532071
R21103 Iout.n835 Iout 0.0532071
R21104 Iout Iout.n847 0.0532071
R21105 Iout.n849 Iout 0.0532071
R21106 Iout Iout.n861 0.0532071
R21107 Iout.n863 Iout 0.0532071
R21108 Iout Iout.n875 0.0532071
R21109 Iout.n877 Iout 0.0532071
R21110 Iout Iout.n889 0.0532071
R21111 Iout Iout.n932 0.0532071
R21112 Iout.n919 Iout 0.0532071
R21113 Iout Iout.n917 0.0532071
R21114 Iout.n905 Iout 0.0532071
R21115 Iout Iout.n903 0.0532071
R21116 Iout.n891 Iout 0.0532071
R21117 Iout.n782 Iout 0.0532071
R21118 Iout.n785 Iout 0.0532071
R21119 Iout.n788 Iout 0.0532071
R21120 Iout.n791 Iout 0.0532071
R21121 Iout.n794 Iout 0.0532071
R21122 Iout.n797 Iout 0.0532071
R21123 Iout.n800 Iout 0.0532071
R21124 Iout.n803 Iout 0.0532071
R21125 Iout.n806 Iout 0.0532071
R21126 Iout.n778 Iout 0.0532071
R21127 Iout Iout.n39 0.0532071
R21128 Iout.n766 Iout 0.0532071
R21129 Iout Iout.n48 0.0532071
R21130 Iout.n754 Iout 0.0532071
R21131 Iout Iout.n54 0.0532071
R21132 Iout.n742 Iout 0.0532071
R21133 Iout Iout.n60 0.0532071
R21134 Iout.n730 Iout 0.0532071
R21135 Iout Iout.n66 0.0532071
R21136 Iout.n945 Iout 0.0532071
R21137 Iout.n78 Iout 0.0532071
R21138 Iout.n706 Iout 0.0532071
R21139 Iout Iout.n72 0.0532071
R21140 Iout.n718 Iout 0.0532071
R21141 Iout Iout.n951 0.0532071
R21142 Iout.n700 Iout 0.0532071
R21143 Iout Iout.n75 0.0532071
R21144 Iout.n712 Iout 0.0532071
R21145 Iout Iout.n69 0.0532071
R21146 Iout.n724 Iout 0.0532071
R21147 Iout Iout.n63 0.0532071
R21148 Iout.n736 Iout 0.0532071
R21149 Iout Iout.n57 0.0532071
R21150 Iout.n748 Iout 0.0532071
R21151 Iout Iout.n655 0.0532071
R21152 Iout Iout.n658 0.0532071
R21153 Iout Iout.n661 0.0532071
R21154 Iout Iout.n664 0.0532071
R21155 Iout Iout.n667 0.0532071
R21156 Iout Iout.n670 0.0532071
R21157 Iout Iout.n673 0.0532071
R21158 Iout Iout.n676 0.0532071
R21159 Iout Iout.n679 0.0532071
R21160 Iout Iout.n682 0.0532071
R21161 Iout Iout.n685 0.0532071
R21162 Iout.n693 Iout 0.0532071
R21163 Iout.n696 Iout 0.0532071
R21164 Iout Iout.n691 0.0532071
R21165 Iout Iout.n688 0.0532071
R21166 Iout.n964 Iout 0.0532071
R21167 Iout.n574 Iout 0.0532071
R21168 Iout.n577 Iout 0.0532071
R21169 Iout Iout.n115 0.0532071
R21170 Iout.n589 Iout 0.0532071
R21171 Iout Iout.n109 0.0532071
R21172 Iout.n601 Iout 0.0532071
R21173 Iout Iout.n103 0.0532071
R21174 Iout.n613 Iout 0.0532071
R21175 Iout Iout.n97 0.0532071
R21176 Iout.n625 Iout 0.0532071
R21177 Iout Iout.n86 0.0532071
R21178 Iout.n643 Iout 0.0532071
R21179 Iout Iout.n88 0.0532071
R21180 Iout.n631 Iout 0.0532071
R21181 Iout Iout.n94 0.0532071
R21182 Iout.n619 Iout 0.0532071
R21183 Iout Iout.n100 0.0532071
R21184 Iout.n607 Iout 0.0532071
R21185 Iout Iout.n106 0.0532071
R21186 Iout.n595 Iout 0.0532071
R21187 Iout Iout.n112 0.0532071
R21188 Iout.n583 Iout 0.0532071
R21189 Iout Iout.n970 0.0532071
R21190 Iout.n564 Iout 0.0532071
R21191 Iout Iout.n118 0.0532071
R21192 Iout.n121 Iout 0.0532071
R21193 Iout.n124 Iout 0.0532071
R21194 Iout.n570 Iout 0.0532071
R21195 Iout.n334 Iout 0.0532071
R21196 Iout.n337 Iout 0.0532071
R21197 Iout.n340 Iout 0.0532071
R21198 Iout.n343 Iout 0.0532071
R21199 Iout.n346 Iout 0.0532071
R21200 Iout.n349 Iout 0.0532071
R21201 Iout.n352 Iout 0.0532071
R21202 Iout.n355 Iout 0.0532071
R21203 Iout.n358 Iout 0.0532071
R21204 Iout.n371 Iout 0.0532071
R21205 Iout Iout.n385 0.0532071
R21206 Iout.n387 Iout 0.0532071
R21207 Iout Iout.n401 0.0532071
R21208 Iout.n403 Iout 0.0532071
R21209 Iout Iout.n417 0.0532071
R21210 Iout.n419 Iout 0.0532071
R21211 Iout Iout.n433 0.0532071
R21212 Iout.n442 Iout 0.0532071
R21213 Iout.n439 Iout 0.0532071
R21214 Iout.n435 Iout 0.0532071
R21215 Iout Iout.n555 0.0532071
R21216 Iout Iout.n558 0.0532071
R21217 Iout.n983 Iout 0.0532071
R21218 Iout.n560 Iout 0.0532071
R21219 Iout Iout.n989 0.0532071
R21220 Iout.n128 Iout 0.0532071
R21221 Iout.n131 Iout 0.0532071
R21222 Iout.n549 Iout 0.0532071
R21223 Iout.n450 Iout 0.0532071
R21224 Iout.n453 Iout 0.0532071
R21225 Iout Iout.n448 0.0532071
R21226 Iout.n427 Iout 0.0532071
R21227 Iout Iout.n425 0.0532071
R21228 Iout.n411 Iout 0.0532071
R21229 Iout Iout.n409 0.0532071
R21230 Iout.n395 Iout 0.0532071
R21231 Iout Iout.n393 0.0532071
R21232 Iout.n330 Iout 0.0532071
R21233 Iout.n327 Iout 0.0532071
R21234 Iout.n324 Iout 0.0532071
R21235 Iout.n321 Iout 0.0532071
R21236 Iout.n318 Iout 0.0532071
R21237 Iout.n315 Iout 0.0532071
R21238 Iout.n312 Iout 0.0532071
R21239 Iout.n309 Iout 0.0532071
R21240 Iout.n306 Iout 0.0532071
R21241 Iout Iout.n459 0.0532071
R21242 Iout.n464 Iout 0.0532071
R21243 Iout.n461 Iout 0.0532071
R21244 Iout.n543 Iout 0.0532071
R21245 Iout.n137 Iout 0.0532071
R21246 Iout.n134 Iout 0.0532071
R21247 Iout.n1002 Iout 0.0532071
R21248 Iout.n537 Iout 0.0532071
R21249 Iout Iout.n535 0.0532071
R21250 Iout Iout.n532 0.0532071
R21251 Iout.n157 Iout 0.0532071
R21252 Iout.n470 Iout 0.0532071
R21253 Iout.n473 Iout 0.0532071
R21254 Iout.n190 Iout 0.0532071
R21255 Iout.n266 Iout 0.0532071
R21256 Iout Iout.n184 0.0532071
R21257 Iout.n278 Iout 0.0532071
R21258 Iout Iout.n178 0.0532071
R21259 Iout.n290 Iout 0.0532071
R21260 Iout Iout.n169 0.0532071
R21261 Iout Iout.n173 0.0532071
R21262 Iout.n296 Iout 0.0532071
R21263 Iout Iout.n175 0.0532071
R21264 Iout.n284 Iout 0.0532071
R21265 Iout Iout.n181 0.0532071
R21266 Iout.n272 Iout 0.0532071
R21267 Iout Iout.n187 0.0532071
R21268 Iout.n260 Iout 0.0532071
R21269 Iout Iout.n479 0.0532071
R21270 Iout.n484 Iout 0.0532071
R21271 Iout.n481 Iout 0.0532071
R21272 Iout.n526 Iout 0.0532071
R21273 Iout.n144 Iout 0.0532071
R21274 Iout.n141 Iout 0.0532071
R21275 Iout Iout.n1008 0.0532071
R21276 Iout.n147 Iout 0.0532071
R21277 Iout.n150 Iout 0.0532071
R21278 Iout.n520 Iout 0.0532071
R21279 Iout.n492 Iout 0.0532071
R21280 Iout.n495 Iout 0.0532071
R21281 Iout Iout.n490 0.0532071
R21282 Iout.n253 Iout 0.0532071
R21283 Iout.n256 Iout 0.0532071
R21284 Iout Iout.n251 0.0532071
R21285 Iout Iout.n248 0.0532071
R21286 Iout Iout.n245 0.0532071
R21287 Iout Iout.n242 0.0532071
R21288 Iout Iout.n239 0.0532071
R21289 Iout Iout.n236 0.0532071
R21290 Iout Iout.n233 0.0532071
R21291 Iout.n227 Iout 0.0532071
R21292 Iout.n223 Iout 0.0532071
R21293 Iout.n219 Iout 0.0532071
R21294 Iout.n215 Iout 0.0532071
R21295 Iout.n211 Iout 0.0532071
R21296 Iout.n207 Iout 0.0532071
R21297 Iout.n203 Iout 0.0532071
R21298 Iout.n200 Iout 0.0532071
R21299 Iout.n196 Iout 0.0532071
R21300 Iout.n193 Iout 0.0532071
R21301 Iout Iout.n501 0.0532071
R21302 Iout Iout.n505 0.0532071
R21303 Iout Iout.n508 0.0532071
R21304 Iout.n514 Iout 0.0532071
R21305 Iout.n510 Iout 0.0532071
R21306 Iout.n1020 Iout 0.03925
R21307 Iout.n509 Iout 0.03925
R21308 Iout.n513 Iout 0.03925
R21309 Iout.n507 Iout 0.03925
R21310 Iout.n504 Iout 0.03925
R21311 Iout.n500 Iout 0.03925
R21312 Iout.n192 Iout 0.03925
R21313 Iout.n195 Iout 0.03925
R21314 Iout.n199 Iout 0.03925
R21315 Iout.n202 Iout 0.03925
R21316 Iout.n206 Iout 0.03925
R21317 Iout.n210 Iout 0.03925
R21318 Iout.n214 Iout 0.03925
R21319 Iout.n218 Iout 0.03925
R21320 Iout.n222 Iout 0.03925
R21321 Iout.n226 Iout 0.03925
R21322 Iout.n232 Iout 0.03925
R21323 Iout.n235 Iout 0.03925
R21324 Iout.n238 Iout 0.03925
R21325 Iout.n241 Iout 0.03925
R21326 Iout.n244 Iout 0.03925
R21327 Iout.n247 Iout 0.03925
R21328 Iout.n250 Iout 0.03925
R21329 Iout.n255 Iout 0.03925
R21330 Iout.n252 Iout 0.03925
R21331 Iout.n489 Iout 0.03925
R21332 Iout.n494 Iout 0.03925
R21333 Iout.n491 Iout 0.03925
R21334 Iout.n519 Iout 0.03925
R21335 Iout.n149 Iout 0.03925
R21336 Iout.n146 Iout 0.03925
R21337 Iout.n1010 Iout 0.03925
R21338 Iout.n1007 Iout 0.03925
R21339 Iout.n140 Iout 0.03925
R21340 Iout.n143 Iout 0.03925
R21341 Iout.n525 Iout 0.03925
R21342 Iout.n480 Iout 0.03925
R21343 Iout.n483 Iout 0.03925
R21344 Iout.n478 Iout 0.03925
R21345 Iout.n259 Iout 0.03925
R21346 Iout.n186 Iout 0.03925
R21347 Iout.n271 Iout 0.03925
R21348 Iout.n180 Iout 0.03925
R21349 Iout.n283 Iout 0.03925
R21350 Iout.n174 Iout 0.03925
R21351 Iout.n168 Iout 0.03925
R21352 Iout.n301 Iout 0.03925
R21353 Iout.n289 Iout 0.03925
R21354 Iout.n177 Iout 0.03925
R21355 Iout.n277 Iout 0.03925
R21356 Iout.n183 Iout 0.03925
R21357 Iout.n265 Iout 0.03925
R21358 Iout.n189 Iout 0.03925
R21359 Iout.n472 Iout 0.03925
R21360 Iout.n469 Iout 0.03925
R21361 Iout.n156 Iout 0.03925
R21362 Iout.n531 Iout 0.03925
R21363 Iout.n534 Iout 0.03925
R21364 Iout.n536 Iout 0.03925
R21365 Iout.n133 Iout 0.03925
R21366 Iout.n136 Iout 0.03925
R21367 Iout.n542 Iout 0.03925
R21368 Iout.n460 Iout 0.03925
R21369 Iout.n463 Iout 0.03925
R21370 Iout.n458 Iout 0.03925
R21371 Iout.n305 Iout 0.03925
R21372 Iout.n308 Iout 0.03925
R21373 Iout.n311 Iout 0.03925
R21374 Iout.n314 Iout 0.03925
R21375 Iout.n317 Iout 0.03925
R21376 Iout.n320 Iout 0.03925
R21377 Iout.n392 Iout 0.03925
R21378 Iout.n378 Iout 0.03925
R21379 Iout.n376 Iout 0.03925
R21380 Iout.n394 Iout 0.03925
R21381 Iout.n408 Iout 0.03925
R21382 Iout.n410 Iout 0.03925
R21383 Iout.n424 Iout 0.03925
R21384 Iout.n426 Iout 0.03925
R21385 Iout.n447 Iout 0.03925
R21386 Iout.n452 Iout 0.03925
R21387 Iout.n449 Iout 0.03925
R21388 Iout.n548 Iout 0.03925
R21389 Iout.n130 Iout 0.03925
R21390 Iout.n559 Iout 0.03925
R21391 Iout.n557 Iout 0.03925
R21392 Iout.n554 Iout 0.03925
R21393 Iout.n434 Iout 0.03925
R21394 Iout.n438 Iout 0.03925
R21395 Iout.n441 Iout 0.03925
R21396 Iout.n432 Iout 0.03925
R21397 Iout.n418 Iout 0.03925
R21398 Iout.n416 Iout 0.03925
R21399 Iout.n402 Iout 0.03925
R21400 Iout.n357 Iout 0.03925
R21401 Iout.n360 Iout 0.03925
R21402 Iout.n363 Iout 0.03925
R21403 Iout.n366 Iout 0.03925
R21404 Iout.n354 Iout 0.03925
R21405 Iout.n351 Iout 0.03925
R21406 Iout.n348 Iout 0.03925
R21407 Iout.n345 Iout 0.03925
R21408 Iout.n342 Iout 0.03925
R21409 Iout.n339 Iout 0.03925
R21410 Iout.n336 Iout 0.03925
R21411 Iout.n333 Iout 0.03925
R21412 Iout.n117 Iout 0.03925
R21413 Iout.n582 Iout 0.03925
R21414 Iout.n111 Iout 0.03925
R21415 Iout.n594 Iout 0.03925
R21416 Iout.n105 Iout 0.03925
R21417 Iout.n606 Iout 0.03925
R21418 Iout.n99 Iout 0.03925
R21419 Iout.n618 Iout 0.03925
R21420 Iout.n624 Iout 0.03925
R21421 Iout.n90 Iout 0.03925
R21422 Iout.n636 Iout 0.03925
R21423 Iout.n81 Iout 0.03925
R21424 Iout.n648 Iout 0.03925
R21425 Iout.n96 Iout 0.03925
R21426 Iout.n612 Iout 0.03925
R21427 Iout.n102 Iout 0.03925
R21428 Iout.n600 Iout 0.03925
R21429 Iout.n108 Iout 0.03925
R21430 Iout.n588 Iout 0.03925
R21431 Iout.n687 Iout 0.03925
R21432 Iout.n684 Iout 0.03925
R21433 Iout.n681 Iout 0.03925
R21434 Iout.n678 Iout 0.03925
R21435 Iout.n675 Iout 0.03925
R21436 Iout.n672 Iout 0.03925
R21437 Iout.n747 Iout 0.03925
R21438 Iout.n50 Iout 0.03925
R21439 Iout.n759 Iout 0.03925
R21440 Iout.n44 Iout 0.03925
R21441 Iout.n771 Iout 0.03925
R21442 Iout.n42 Iout 0.03925
R21443 Iout.n56 Iout 0.03925
R21444 Iout.n735 Iout 0.03925
R21445 Iout.n62 Iout 0.03925
R21446 Iout.n723 Iout 0.03925
R21447 Iout.n717 Iout 0.03925
R21448 Iout.n65 Iout 0.03925
R21449 Iout.n729 Iout 0.03925
R21450 Iout.n59 Iout 0.03925
R21451 Iout.n805 Iout 0.03925
R21452 Iout.n808 Iout 0.03925
R21453 Iout.n811 Iout 0.03925
R21454 Iout.n814 Iout 0.03925
R21455 Iout.n817 Iout 0.03925
R21456 Iout.n820 Iout 0.03925
R21457 Iout.n823 Iout 0.03925
R21458 Iout.n802 Iout 0.03925
R21459 Iout.n799 Iout 0.03925
R21460 Iout.n890 Iout 0.03925
R21461 Iout.n888 Iout 0.03925
R21462 Iout.n881 Iout 0.03925
R21463 Iout.n869 Iout 0.03925
R21464 Iout.n867 Iout 0.03925
R21465 Iout.n855 Iout 0.03925
R21466 Iout.n853 Iout 0.03925
R21467 Iout.n841 Iout 0.03925
R21468 Iout.n839 Iout 0.03925
R21469 Iout.n827 Iout 0.03925
R21470 Iout.n883 Iout 0.03925
R21471 Iout.n895 Iout 0.03925
R21472 Iout.n897 Iout 0.03925
R21473 Iout.n909 Iout 0.03925
R21474 Iout.n911 Iout 0.03925
R21475 Iout.n923 Iout 0.03925
R21476 Iout.n926 Iout 0.03925
R21477 Iout.n22 Iout 0.03925
R21478 Iout.n876 Iout 0.03925
R21479 Iout.n874 Iout 0.03925
R21480 Iout.n862 Iout 0.03925
R21481 Iout.n860 Iout 0.03925
R21482 Iout.n848 Iout 0.03925
R21483 Iout.n846 Iout 0.03925
R21484 Iout.n834 Iout 0.03925
R21485 Iout.n832 Iout 0.03925
R21486 Iout.n902 Iout 0.03925
R21487 Iout.n904 Iout 0.03925
R21488 Iout.n916 Iout 0.03925
R21489 Iout.n918 Iout 0.03925
R21490 Iout.n931 Iout 0.03925
R21491 Iout.n934 Iout 0.03925
R21492 Iout.n796 Iout 0.03925
R21493 Iout.n793 Iout 0.03925
R21494 Iout.n790 Iout 0.03925
R21495 Iout.n787 Iout 0.03925
R21496 Iout.n784 Iout 0.03925
R21497 Iout.n781 Iout 0.03925
R21498 Iout.n938 Iout 0.03925
R21499 Iout.n741 Iout 0.03925
R21500 Iout.n53 Iout 0.03925
R21501 Iout.n753 Iout 0.03925
R21502 Iout.n47 Iout 0.03925
R21503 Iout.n765 Iout 0.03925
R21504 Iout.n38 Iout 0.03925
R21505 Iout.n777 Iout 0.03925
R21506 Iout.n71 Iout 0.03925
R21507 Iout.n705 Iout 0.03925
R21508 Iout.n77 Iout 0.03925
R21509 Iout.n944 Iout 0.03925
R21510 Iout.n19 Iout 0.03925
R21511 Iout.n68 Iout 0.03925
R21512 Iout.n711 Iout 0.03925
R21513 Iout.n74 Iout 0.03925
R21514 Iout.n699 Iout 0.03925
R21515 Iout.n950 Iout 0.03925
R21516 Iout.n953 Iout 0.03925
R21517 Iout.n669 Iout 0.03925
R21518 Iout.n666 Iout 0.03925
R21519 Iout.n663 Iout 0.03925
R21520 Iout.n660 Iout 0.03925
R21521 Iout.n657 Iout 0.03925
R21522 Iout.n654 Iout 0.03925
R21523 Iout.n690 Iout 0.03925
R21524 Iout.n695 Iout 0.03925
R21525 Iout.n692 Iout 0.03925
R21526 Iout.n957 Iout 0.03925
R21527 Iout.n114 Iout 0.03925
R21528 Iout.n576 Iout 0.03925
R21529 Iout.n573 Iout 0.03925
R21530 Iout.n963 Iout 0.03925
R21531 Iout.n14 Iout 0.03925
R21532 Iout.n93 Iout 0.03925
R21533 Iout.n630 Iout 0.03925
R21534 Iout.n87 Iout 0.03925
R21535 Iout.n642 Iout 0.03925
R21536 Iout.n85 Iout 0.03925
R21537 Iout.n563 Iout 0.03925
R21538 Iout.n969 Iout 0.03925
R21539 Iout.n972 Iout 0.03925
R21540 Iout.n569 Iout 0.03925
R21541 Iout.n123 Iout 0.03925
R21542 Iout.n120 Iout 0.03925
R21543 Iout.n976 Iout 0.03925
R21544 Iout.n400 Iout 0.03925
R21545 Iout.n386 Iout 0.03925
R21546 Iout.n384 Iout 0.03925
R21547 Iout.n370 Iout 0.03925
R21548 Iout.n982 Iout 0.03925
R21549 Iout.n9 Iout 0.03925
R21550 Iout.n127 Iout 0.03925
R21551 Iout.n988 Iout 0.03925
R21552 Iout.n991 Iout 0.03925
R21553 Iout.n323 Iout 0.03925
R21554 Iout.n326 Iout 0.03925
R21555 Iout.n329 Iout 0.03925
R21556 Iout.n995 Iout 0.03925
R21557 Iout.n1001 Iout 0.03925
R21558 Iout.n4 Iout 0.03925
R21559 Iout.n295 Iout 0.03925
R21560 Iout.n172 Iout 0.03925
R21561 Iout.n1014 Iout 0.03925
R21562 Iout.n1022 Iout 0.02071
R21563 Iout Iout.n1022 0.00379
R21564 Iout.n303 Iout.n302 0.00105952
R21565 Iout.n377 Iout.n375 0.00105952
R21566 Iout.n380 Iout.n379 0.00105952
R21567 Iout.n368 Iout.n367 0.00105952
R21568 Iout.n365 Iout.n364 0.00105952
R21569 Iout.n362 Iout.n361 0.00105952
R21570 Iout.n650 Iout.n649 0.00105952
R21571 Iout.n647 Iout.n82 0.00105952
R21572 Iout.n638 Iout.n637 0.00105952
R21573 Iout.n635 Iout.n91 0.00105952
R21574 Iout.n43 Iout.n41 0.00105952
R21575 Iout.n773 Iout.n772 0.00105952
R21576 Iout.n770 Iout.n45 0.00105952
R21577 Iout.n761 Iout.n760 0.00105952
R21578 Iout.n758 Iout.n51 0.00105952
R21579 Iout.n825 Iout.n824 0.00105952
R21580 Iout.n822 Iout.n821 0.00105952
R21581 Iout.n819 Iout.n818 0.00105952
R21582 Iout.n816 Iout.n815 0.00105952
R21583 Iout.n813 Iout.n812 0.00105952
R21584 Iout.n810 Iout.n809 0.00105952
R21585 Iout.n829 Iout.n828 0.00105952
R21586 Iout.n840 Iout.n838 0.00105952
R21587 Iout.n843 Iout.n842 0.00105952
R21588 Iout.n854 Iout.n852 0.00105952
R21589 Iout.n857 Iout.n856 0.00105952
R21590 Iout.n868 Iout.n866 0.00105952
R21591 Iout.n871 Iout.n870 0.00105952
R21592 Iout.n925 Iout.n23 0.00105952
R21593 Iout.n928 Iout.n927 0.00105952
R21594 Iout.n924 Iout.n922 0.00105952
R21595 Iout.n913 Iout.n912 0.00105952
R21596 Iout.n910 Iout.n908 0.00105952
R21597 Iout.n899 Iout.n898 0.00105952
R21598 Iout.n896 Iout.n894 0.00105952
R21599 Iout.n885 Iout.n884 0.00105952
R21600 Iout.n882 Iout.n880 0.00105952
R21601 Iout.n833 Iout.n831 0.00105952
R21602 Iout.n836 Iout.n835 0.00105952
R21603 Iout.n847 Iout.n845 0.00105952
R21604 Iout.n850 Iout.n849 0.00105952
R21605 Iout.n861 Iout.n859 0.00105952
R21606 Iout.n864 Iout.n863 0.00105952
R21607 Iout.n875 Iout.n873 0.00105952
R21608 Iout.n878 Iout.n877 0.00105952
R21609 Iout.n889 Iout.n887 0.00105952
R21610 Iout.n935 Iout.n933 0.00105952
R21611 Iout.n932 Iout.n930 0.00105952
R21612 Iout.n920 Iout.n919 0.00105952
R21613 Iout.n917 Iout.n915 0.00105952
R21614 Iout.n906 Iout.n905 0.00105952
R21615 Iout.n903 Iout.n901 0.00105952
R21616 Iout.n892 Iout.n891 0.00105952
R21617 Iout.n940 Iout.n939 0.00105952
R21618 Iout.n783 Iout.n782 0.00105952
R21619 Iout.n786 Iout.n785 0.00105952
R21620 Iout.n789 Iout.n788 0.00105952
R21621 Iout.n792 Iout.n791 0.00105952
R21622 Iout.n795 Iout.n794 0.00105952
R21623 Iout.n798 Iout.n797 0.00105952
R21624 Iout.n801 Iout.n800 0.00105952
R21625 Iout.n804 Iout.n803 0.00105952
R21626 Iout.n807 Iout.n806 0.00105952
R21627 Iout.n779 Iout.n778 0.00105952
R21628 Iout.n776 Iout.n39 0.00105952
R21629 Iout.n767 Iout.n766 0.00105952
R21630 Iout.n764 Iout.n48 0.00105952
R21631 Iout.n755 Iout.n754 0.00105952
R21632 Iout.n752 Iout.n54 0.00105952
R21633 Iout.n743 Iout.n742 0.00105952
R21634 Iout.n740 Iout.n60 0.00105952
R21635 Iout.n731 Iout.n730 0.00105952
R21636 Iout.n728 Iout.n66 0.00105952
R21637 Iout.n943 Iout.n20 0.00105952
R21638 Iout.n946 Iout.n945 0.00105952
R21639 Iout.n704 Iout.n78 0.00105952
R21640 Iout.n707 Iout.n706 0.00105952
R21641 Iout.n716 Iout.n72 0.00105952
R21642 Iout.n719 Iout.n718 0.00105952
R21643 Iout.n954 Iout.n952 0.00105952
R21644 Iout.n951 Iout.n949 0.00105952
R21645 Iout.n701 Iout.n700 0.00105952
R21646 Iout.n710 Iout.n75 0.00105952
R21647 Iout.n713 Iout.n712 0.00105952
R21648 Iout.n722 Iout.n69 0.00105952
R21649 Iout.n725 Iout.n724 0.00105952
R21650 Iout.n734 Iout.n63 0.00105952
R21651 Iout.n737 Iout.n736 0.00105952
R21652 Iout.n746 Iout.n57 0.00105952
R21653 Iout.n749 Iout.n748 0.00105952
R21654 Iout.n655 Iout.n653 0.00105952
R21655 Iout.n658 Iout.n656 0.00105952
R21656 Iout.n661 Iout.n659 0.00105952
R21657 Iout.n664 Iout.n662 0.00105952
R21658 Iout.n667 Iout.n665 0.00105952
R21659 Iout.n670 Iout.n668 0.00105952
R21660 Iout.n673 Iout.n671 0.00105952
R21661 Iout.n676 Iout.n674 0.00105952
R21662 Iout.n679 Iout.n677 0.00105952
R21663 Iout.n682 Iout.n680 0.00105952
R21664 Iout.n685 Iout.n683 0.00105952
R21665 Iout.n959 Iout.n958 0.00105952
R21666 Iout.n694 Iout.n693 0.00105952
R21667 Iout.n697 Iout.n696 0.00105952
R21668 Iout.n691 Iout.n689 0.00105952
R21669 Iout.n688 Iout.n686 0.00105952
R21670 Iout.n962 Iout.n15 0.00105952
R21671 Iout.n965 Iout.n964 0.00105952
R21672 Iout.n575 Iout.n574 0.00105952
R21673 Iout.n578 Iout.n577 0.00105952
R21674 Iout.n587 Iout.n115 0.00105952
R21675 Iout.n590 Iout.n589 0.00105952
R21676 Iout.n599 Iout.n109 0.00105952
R21677 Iout.n602 Iout.n601 0.00105952
R21678 Iout.n611 Iout.n103 0.00105952
R21679 Iout.n614 Iout.n613 0.00105952
R21680 Iout.n623 Iout.n97 0.00105952
R21681 Iout.n626 Iout.n625 0.00105952
R21682 Iout.n86 Iout.n84 0.00105952
R21683 Iout.n644 Iout.n643 0.00105952
R21684 Iout.n641 Iout.n88 0.00105952
R21685 Iout.n632 Iout.n631 0.00105952
R21686 Iout.n629 Iout.n94 0.00105952
R21687 Iout.n620 Iout.n619 0.00105952
R21688 Iout.n617 Iout.n100 0.00105952
R21689 Iout.n608 Iout.n607 0.00105952
R21690 Iout.n605 Iout.n106 0.00105952
R21691 Iout.n596 Iout.n595 0.00105952
R21692 Iout.n593 Iout.n112 0.00105952
R21693 Iout.n584 Iout.n583 0.00105952
R21694 Iout.n973 Iout.n971 0.00105952
R21695 Iout.n970 Iout.n968 0.00105952
R21696 Iout.n565 Iout.n564 0.00105952
R21697 Iout.n581 Iout.n118 0.00105952
R21698 Iout.n978 Iout.n977 0.00105952
R21699 Iout.n122 Iout.n121 0.00105952
R21700 Iout.n568 Iout.n124 0.00105952
R21701 Iout.n571 Iout.n570 0.00105952
R21702 Iout.n335 Iout.n334 0.00105952
R21703 Iout.n338 Iout.n337 0.00105952
R21704 Iout.n341 Iout.n340 0.00105952
R21705 Iout.n344 Iout.n343 0.00105952
R21706 Iout.n347 Iout.n346 0.00105952
R21707 Iout.n350 Iout.n349 0.00105952
R21708 Iout.n353 Iout.n352 0.00105952
R21709 Iout.n356 Iout.n355 0.00105952
R21710 Iout.n359 Iout.n358 0.00105952
R21711 Iout.n372 Iout.n371 0.00105952
R21712 Iout.n385 Iout.n383 0.00105952
R21713 Iout.n388 Iout.n387 0.00105952
R21714 Iout.n401 Iout.n399 0.00105952
R21715 Iout.n404 Iout.n403 0.00105952
R21716 Iout.n417 Iout.n415 0.00105952
R21717 Iout.n420 Iout.n419 0.00105952
R21718 Iout.n433 Iout.n431 0.00105952
R21719 Iout.n443 Iout.n442 0.00105952
R21720 Iout.n440 Iout.n439 0.00105952
R21721 Iout.n437 Iout.n435 0.00105952
R21722 Iout.n555 Iout.n553 0.00105952
R21723 Iout.n558 Iout.n556 0.00105952
R21724 Iout.n981 Iout.n10 0.00105952
R21725 Iout.n984 Iout.n983 0.00105952
R21726 Iout.n561 Iout.n560 0.00105952
R21727 Iout.n992 Iout.n990 0.00105952
R21728 Iout.n989 Iout.n987 0.00105952
R21729 Iout.n129 Iout.n128 0.00105952
R21730 Iout.n547 Iout.n131 0.00105952
R21731 Iout.n550 Iout.n549 0.00105952
R21732 Iout.n451 Iout.n450 0.00105952
R21733 Iout.n454 Iout.n453 0.00105952
R21734 Iout.n448 Iout.n446 0.00105952
R21735 Iout.n428 Iout.n427 0.00105952
R21736 Iout.n425 Iout.n423 0.00105952
R21737 Iout.n412 Iout.n411 0.00105952
R21738 Iout.n409 Iout.n407 0.00105952
R21739 Iout.n396 Iout.n395 0.00105952
R21740 Iout.n393 Iout.n391 0.00105952
R21741 Iout.n331 Iout.n330 0.00105952
R21742 Iout.n328 Iout.n327 0.00105952
R21743 Iout.n325 Iout.n324 0.00105952
R21744 Iout.n322 Iout.n321 0.00105952
R21745 Iout.n319 Iout.n318 0.00105952
R21746 Iout.n316 Iout.n315 0.00105952
R21747 Iout.n313 Iout.n312 0.00105952
R21748 Iout.n310 Iout.n309 0.00105952
R21749 Iout.n307 Iout.n306 0.00105952
R21750 Iout.n459 Iout.n457 0.00105952
R21751 Iout.n465 Iout.n464 0.00105952
R21752 Iout.n462 Iout.n461 0.00105952
R21753 Iout.n544 Iout.n543 0.00105952
R21754 Iout.n541 Iout.n137 0.00105952
R21755 Iout.n997 Iout.n996 0.00105952
R21756 Iout.n135 Iout.n134 0.00105952
R21757 Iout.n1000 Iout.n5 0.00105952
R21758 Iout.n1003 Iout.n1002 0.00105952
R21759 Iout.n538 Iout.n537 0.00105952
R21760 Iout.n535 Iout.n533 0.00105952
R21761 Iout.n532 Iout.n530 0.00105952
R21762 Iout.n468 Iout.n157 0.00105952
R21763 Iout.n471 Iout.n470 0.00105952
R21764 Iout.n474 Iout.n473 0.00105952
R21765 Iout.n264 Iout.n190 0.00105952
R21766 Iout.n267 Iout.n266 0.00105952
R21767 Iout.n276 Iout.n184 0.00105952
R21768 Iout.n279 Iout.n278 0.00105952
R21769 Iout.n288 Iout.n178 0.00105952
R21770 Iout.n291 Iout.n290 0.00105952
R21771 Iout.n300 Iout.n169 0.00105952
R21772 Iout.n173 Iout.n171 0.00105952
R21773 Iout.n297 Iout.n296 0.00105952
R21774 Iout.n294 Iout.n175 0.00105952
R21775 Iout.n285 Iout.n284 0.00105952
R21776 Iout.n282 Iout.n181 0.00105952
R21777 Iout.n273 Iout.n272 0.00105952
R21778 Iout.n270 Iout.n187 0.00105952
R21779 Iout.n261 Iout.n260 0.00105952
R21780 Iout.n479 Iout.n477 0.00105952
R21781 Iout.n485 Iout.n484 0.00105952
R21782 Iout.n482 Iout.n481 0.00105952
R21783 Iout.n527 Iout.n526 0.00105952
R21784 Iout.n524 Iout.n144 0.00105952
R21785 Iout.n142 Iout.n141 0.00105952
R21786 Iout.n1008 Iout.n1006 0.00105952
R21787 Iout.n1011 Iout.n1009 0.00105952
R21788 Iout.n1016 Iout.n1015 0.00105952
R21789 Iout.n148 Iout.n147 0.00105952
R21790 Iout.n518 Iout.n150 0.00105952
R21791 Iout.n521 Iout.n520 0.00105952
R21792 Iout.n493 Iout.n492 0.00105952
R21793 Iout.n496 Iout.n495 0.00105952
R21794 Iout.n490 Iout.n488 0.00105952
R21795 Iout.n254 Iout.n253 0.00105952
R21796 Iout.n257 Iout.n256 0.00105952
R21797 Iout.n251 Iout.n249 0.00105952
R21798 Iout.n248 Iout.n246 0.00105952
R21799 Iout.n245 Iout.n243 0.00105952
R21800 Iout.n242 Iout.n240 0.00105952
R21801 Iout.n239 Iout.n237 0.00105952
R21802 Iout.n236 Iout.n234 0.00105952
R21803 Iout.n233 Iout.n231 0.00105952
R21804 Iout.n228 Iout.n227 0.00105952
R21805 Iout.n225 Iout.n223 0.00105952
R21806 Iout.n221 Iout.n219 0.00105952
R21807 Iout.n217 Iout.n215 0.00105952
R21808 Iout.n213 Iout.n211 0.00105952
R21809 Iout.n209 Iout.n207 0.00105952
R21810 Iout.n205 Iout.n203 0.00105952
R21811 Iout.n201 Iout.n200 0.00105952
R21812 Iout.n198 Iout.n196 0.00105952
R21813 Iout.n194 Iout.n193 0.00105952
R21814 Iout.n501 Iout.n499 0.00105952
R21815 Iout.n505 Iout.n503 0.00105952
R21816 Iout.n508 Iout.n506 0.00105952
R21817 Iout.n515 Iout.n514 0.00105952
R21818 Iout.n512 Iout.n510 0.00105952
R21819 Iout.n1021 Iout.n1019 0.00105952
R21820 XThC.Tn[2].n74 XThC.Tn[2].n72 332.332
R21821 XThC.Tn[2].n74 XThC.Tn[2].n73 296.493
R21822 XThC.Tn[2].n68 XThC.Tn[2].n66 161.365
R21823 XThC.Tn[2].n64 XThC.Tn[2].n62 161.365
R21824 XThC.Tn[2].n60 XThC.Tn[2].n58 161.365
R21825 XThC.Tn[2].n56 XThC.Tn[2].n54 161.365
R21826 XThC.Tn[2].n52 XThC.Tn[2].n50 161.365
R21827 XThC.Tn[2].n48 XThC.Tn[2].n46 161.365
R21828 XThC.Tn[2].n44 XThC.Tn[2].n42 161.365
R21829 XThC.Tn[2].n40 XThC.Tn[2].n38 161.365
R21830 XThC.Tn[2].n36 XThC.Tn[2].n34 161.365
R21831 XThC.Tn[2].n32 XThC.Tn[2].n30 161.365
R21832 XThC.Tn[2].n28 XThC.Tn[2].n26 161.365
R21833 XThC.Tn[2].n24 XThC.Tn[2].n22 161.365
R21834 XThC.Tn[2].n20 XThC.Tn[2].n18 161.365
R21835 XThC.Tn[2].n16 XThC.Tn[2].n14 161.365
R21836 XThC.Tn[2].n12 XThC.Tn[2].n10 161.365
R21837 XThC.Tn[2].n9 XThC.Tn[2].n7 161.365
R21838 XThC.Tn[2].n66 XThC.Tn[2].t24 161.202
R21839 XThC.Tn[2].n62 XThC.Tn[2].t14 161.202
R21840 XThC.Tn[2].n58 XThC.Tn[2].t33 161.202
R21841 XThC.Tn[2].n54 XThC.Tn[2].t30 161.202
R21842 XThC.Tn[2].n50 XThC.Tn[2].t22 161.202
R21843 XThC.Tn[2].n46 XThC.Tn[2].t41 161.202
R21844 XThC.Tn[2].n42 XThC.Tn[2].t40 161.202
R21845 XThC.Tn[2].n38 XThC.Tn[2].t21 161.202
R21846 XThC.Tn[2].n34 XThC.Tn[2].t19 161.202
R21847 XThC.Tn[2].n30 XThC.Tn[2].t42 161.202
R21848 XThC.Tn[2].n26 XThC.Tn[2].t29 161.202
R21849 XThC.Tn[2].n22 XThC.Tn[2].t28 161.202
R21850 XThC.Tn[2].n18 XThC.Tn[2].t39 161.202
R21851 XThC.Tn[2].n14 XThC.Tn[2].t37 161.202
R21852 XThC.Tn[2].n10 XThC.Tn[2].t35 161.202
R21853 XThC.Tn[2].n7 XThC.Tn[2].t18 161.202
R21854 XThC.Tn[2].n66 XThC.Tn[2].t27 145.137
R21855 XThC.Tn[2].n62 XThC.Tn[2].t17 145.137
R21856 XThC.Tn[2].n58 XThC.Tn[2].t36 145.137
R21857 XThC.Tn[2].n54 XThC.Tn[2].t34 145.137
R21858 XThC.Tn[2].n50 XThC.Tn[2].t26 145.137
R21859 XThC.Tn[2].n46 XThC.Tn[2].t15 145.137
R21860 XThC.Tn[2].n42 XThC.Tn[2].t13 145.137
R21861 XThC.Tn[2].n38 XThC.Tn[2].t25 145.137
R21862 XThC.Tn[2].n34 XThC.Tn[2].t23 145.137
R21863 XThC.Tn[2].n30 XThC.Tn[2].t16 145.137
R21864 XThC.Tn[2].n26 XThC.Tn[2].t32 145.137
R21865 XThC.Tn[2].n22 XThC.Tn[2].t31 145.137
R21866 XThC.Tn[2].n18 XThC.Tn[2].t12 145.137
R21867 XThC.Tn[2].n14 XThC.Tn[2].t43 145.137
R21868 XThC.Tn[2].n10 XThC.Tn[2].t38 145.137
R21869 XThC.Tn[2].n7 XThC.Tn[2].t20 145.137
R21870 XThC.Tn[2].n2 XThC.Tn[2].n0 135.248
R21871 XThC.Tn[2].n2 XThC.Tn[2].n1 98.982
R21872 XThC.Tn[2].n4 XThC.Tn[2].n3 98.982
R21873 XThC.Tn[2].n6 XThC.Tn[2].n5 98.982
R21874 XThC.Tn[2].n4 XThC.Tn[2].n2 36.2672
R21875 XThC.Tn[2].n6 XThC.Tn[2].n4 36.2672
R21876 XThC.Tn[2].n71 XThC.Tn[2].n6 32.6405
R21877 XThC.Tn[2].n72 XThC.Tn[2].t1 26.5955
R21878 XThC.Tn[2].n72 XThC.Tn[2].t0 26.5955
R21879 XThC.Tn[2].n73 XThC.Tn[2].t3 26.5955
R21880 XThC.Tn[2].n73 XThC.Tn[2].t2 26.5955
R21881 XThC.Tn[2].n0 XThC.Tn[2].t11 24.9236
R21882 XThC.Tn[2].n0 XThC.Tn[2].t8 24.9236
R21883 XThC.Tn[2].n1 XThC.Tn[2].t9 24.9236
R21884 XThC.Tn[2].n1 XThC.Tn[2].t10 24.9236
R21885 XThC.Tn[2].n3 XThC.Tn[2].t5 24.9236
R21886 XThC.Tn[2].n3 XThC.Tn[2].t4 24.9236
R21887 XThC.Tn[2].n5 XThC.Tn[2].t7 24.9236
R21888 XThC.Tn[2].n5 XThC.Tn[2].t6 24.9236
R21889 XThC.Tn[2].n75 XThC.Tn[2].n74 18.5605
R21890 XThC.Tn[2].n75 XThC.Tn[2].n71 11.5205
R21891 XThC.Tn[2] XThC.Tn[2].n9 8.0245
R21892 XThC.Tn[2].n69 XThC.Tn[2].n68 7.9105
R21893 XThC.Tn[2].n65 XThC.Tn[2].n64 7.9105
R21894 XThC.Tn[2].n61 XThC.Tn[2].n60 7.9105
R21895 XThC.Tn[2].n57 XThC.Tn[2].n56 7.9105
R21896 XThC.Tn[2].n53 XThC.Tn[2].n52 7.9105
R21897 XThC.Tn[2].n49 XThC.Tn[2].n48 7.9105
R21898 XThC.Tn[2].n45 XThC.Tn[2].n44 7.9105
R21899 XThC.Tn[2].n41 XThC.Tn[2].n40 7.9105
R21900 XThC.Tn[2].n37 XThC.Tn[2].n36 7.9105
R21901 XThC.Tn[2].n33 XThC.Tn[2].n32 7.9105
R21902 XThC.Tn[2].n29 XThC.Tn[2].n28 7.9105
R21903 XThC.Tn[2].n25 XThC.Tn[2].n24 7.9105
R21904 XThC.Tn[2].n21 XThC.Tn[2].n20 7.9105
R21905 XThC.Tn[2].n17 XThC.Tn[2].n16 7.9105
R21906 XThC.Tn[2].n13 XThC.Tn[2].n12 7.9105
R21907 XThC.Tn[2].n70 XThC.Tn[2] 5.58686
R21908 XThC.Tn[2].n71 XThC.Tn[2].n70 4.6005
R21909 XThC.Tn[2].n70 XThC.Tn[2] 1.83383
R21910 XThC.Tn[2] XThC.Tn[2].n75 0.6405
R21911 XThC.Tn[2].n13 XThC.Tn[2] 0.235138
R21912 XThC.Tn[2].n17 XThC.Tn[2] 0.235138
R21913 XThC.Tn[2].n21 XThC.Tn[2] 0.235138
R21914 XThC.Tn[2].n25 XThC.Tn[2] 0.235138
R21915 XThC.Tn[2].n29 XThC.Tn[2] 0.235138
R21916 XThC.Tn[2].n33 XThC.Tn[2] 0.235138
R21917 XThC.Tn[2].n37 XThC.Tn[2] 0.235138
R21918 XThC.Tn[2].n41 XThC.Tn[2] 0.235138
R21919 XThC.Tn[2].n45 XThC.Tn[2] 0.235138
R21920 XThC.Tn[2].n49 XThC.Tn[2] 0.235138
R21921 XThC.Tn[2].n53 XThC.Tn[2] 0.235138
R21922 XThC.Tn[2].n57 XThC.Tn[2] 0.235138
R21923 XThC.Tn[2].n61 XThC.Tn[2] 0.235138
R21924 XThC.Tn[2].n65 XThC.Tn[2] 0.235138
R21925 XThC.Tn[2].n69 XThC.Tn[2] 0.235138
R21926 XThC.Tn[2] XThC.Tn[2].n13 0.114505
R21927 XThC.Tn[2] XThC.Tn[2].n17 0.114505
R21928 XThC.Tn[2] XThC.Tn[2].n21 0.114505
R21929 XThC.Tn[2] XThC.Tn[2].n25 0.114505
R21930 XThC.Tn[2] XThC.Tn[2].n29 0.114505
R21931 XThC.Tn[2] XThC.Tn[2].n33 0.114505
R21932 XThC.Tn[2] XThC.Tn[2].n37 0.114505
R21933 XThC.Tn[2] XThC.Tn[2].n41 0.114505
R21934 XThC.Tn[2] XThC.Tn[2].n45 0.114505
R21935 XThC.Tn[2] XThC.Tn[2].n49 0.114505
R21936 XThC.Tn[2] XThC.Tn[2].n53 0.114505
R21937 XThC.Tn[2] XThC.Tn[2].n57 0.114505
R21938 XThC.Tn[2] XThC.Tn[2].n61 0.114505
R21939 XThC.Tn[2] XThC.Tn[2].n65 0.114505
R21940 XThC.Tn[2] XThC.Tn[2].n69 0.114505
R21941 XThC.Tn[2].n68 XThC.Tn[2].n67 0.0599512
R21942 XThC.Tn[2].n64 XThC.Tn[2].n63 0.0599512
R21943 XThC.Tn[2].n60 XThC.Tn[2].n59 0.0599512
R21944 XThC.Tn[2].n56 XThC.Tn[2].n55 0.0599512
R21945 XThC.Tn[2].n52 XThC.Tn[2].n51 0.0599512
R21946 XThC.Tn[2].n48 XThC.Tn[2].n47 0.0599512
R21947 XThC.Tn[2].n44 XThC.Tn[2].n43 0.0599512
R21948 XThC.Tn[2].n40 XThC.Tn[2].n39 0.0599512
R21949 XThC.Tn[2].n36 XThC.Tn[2].n35 0.0599512
R21950 XThC.Tn[2].n32 XThC.Tn[2].n31 0.0599512
R21951 XThC.Tn[2].n28 XThC.Tn[2].n27 0.0599512
R21952 XThC.Tn[2].n24 XThC.Tn[2].n23 0.0599512
R21953 XThC.Tn[2].n20 XThC.Tn[2].n19 0.0599512
R21954 XThC.Tn[2].n16 XThC.Tn[2].n15 0.0599512
R21955 XThC.Tn[2].n12 XThC.Tn[2].n11 0.0599512
R21956 XThC.Tn[2].n9 XThC.Tn[2].n8 0.0599512
R21957 XThC.Tn[2].n67 XThC.Tn[2] 0.0469286
R21958 XThC.Tn[2].n63 XThC.Tn[2] 0.0469286
R21959 XThC.Tn[2].n59 XThC.Tn[2] 0.0469286
R21960 XThC.Tn[2].n55 XThC.Tn[2] 0.0469286
R21961 XThC.Tn[2].n51 XThC.Tn[2] 0.0469286
R21962 XThC.Tn[2].n47 XThC.Tn[2] 0.0469286
R21963 XThC.Tn[2].n43 XThC.Tn[2] 0.0469286
R21964 XThC.Tn[2].n39 XThC.Tn[2] 0.0469286
R21965 XThC.Tn[2].n35 XThC.Tn[2] 0.0469286
R21966 XThC.Tn[2].n31 XThC.Tn[2] 0.0469286
R21967 XThC.Tn[2].n27 XThC.Tn[2] 0.0469286
R21968 XThC.Tn[2].n23 XThC.Tn[2] 0.0469286
R21969 XThC.Tn[2].n19 XThC.Tn[2] 0.0469286
R21970 XThC.Tn[2].n15 XThC.Tn[2] 0.0469286
R21971 XThC.Tn[2].n11 XThC.Tn[2] 0.0469286
R21972 XThC.Tn[2].n8 XThC.Tn[2] 0.0469286
R21973 XThC.Tn[2].n67 XThC.Tn[2] 0.0401341
R21974 XThC.Tn[2].n63 XThC.Tn[2] 0.0401341
R21975 XThC.Tn[2].n59 XThC.Tn[2] 0.0401341
R21976 XThC.Tn[2].n55 XThC.Tn[2] 0.0401341
R21977 XThC.Tn[2].n51 XThC.Tn[2] 0.0401341
R21978 XThC.Tn[2].n47 XThC.Tn[2] 0.0401341
R21979 XThC.Tn[2].n43 XThC.Tn[2] 0.0401341
R21980 XThC.Tn[2].n39 XThC.Tn[2] 0.0401341
R21981 XThC.Tn[2].n35 XThC.Tn[2] 0.0401341
R21982 XThC.Tn[2].n31 XThC.Tn[2] 0.0401341
R21983 XThC.Tn[2].n27 XThC.Tn[2] 0.0401341
R21984 XThC.Tn[2].n23 XThC.Tn[2] 0.0401341
R21985 XThC.Tn[2].n19 XThC.Tn[2] 0.0401341
R21986 XThC.Tn[2].n15 XThC.Tn[2] 0.0401341
R21987 XThC.Tn[2].n11 XThC.Tn[2] 0.0401341
R21988 XThC.Tn[2].n8 XThC.Tn[2] 0.0401341
R21989 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R21990 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R21991 XThC.Tn[1].n71 XThC.Tn[1].n69 161.365
R21992 XThC.Tn[1].n67 XThC.Tn[1].n65 161.365
R21993 XThC.Tn[1].n63 XThC.Tn[1].n61 161.365
R21994 XThC.Tn[1].n59 XThC.Tn[1].n57 161.365
R21995 XThC.Tn[1].n55 XThC.Tn[1].n53 161.365
R21996 XThC.Tn[1].n51 XThC.Tn[1].n49 161.365
R21997 XThC.Tn[1].n47 XThC.Tn[1].n45 161.365
R21998 XThC.Tn[1].n43 XThC.Tn[1].n41 161.365
R21999 XThC.Tn[1].n39 XThC.Tn[1].n37 161.365
R22000 XThC.Tn[1].n35 XThC.Tn[1].n33 161.365
R22001 XThC.Tn[1].n31 XThC.Tn[1].n29 161.365
R22002 XThC.Tn[1].n27 XThC.Tn[1].n25 161.365
R22003 XThC.Tn[1].n23 XThC.Tn[1].n21 161.365
R22004 XThC.Tn[1].n19 XThC.Tn[1].n17 161.365
R22005 XThC.Tn[1].n15 XThC.Tn[1].n13 161.365
R22006 XThC.Tn[1].n12 XThC.Tn[1].n10 161.365
R22007 XThC.Tn[1].n69 XThC.Tn[1].t35 161.202
R22008 XThC.Tn[1].n65 XThC.Tn[1].t25 161.202
R22009 XThC.Tn[1].n61 XThC.Tn[1].t12 161.202
R22010 XThC.Tn[1].n57 XThC.Tn[1].t41 161.202
R22011 XThC.Tn[1].n53 XThC.Tn[1].t33 161.202
R22012 XThC.Tn[1].n49 XThC.Tn[1].t20 161.202
R22013 XThC.Tn[1].n45 XThC.Tn[1].t19 161.202
R22014 XThC.Tn[1].n41 XThC.Tn[1].t32 161.202
R22015 XThC.Tn[1].n37 XThC.Tn[1].t30 161.202
R22016 XThC.Tn[1].n33 XThC.Tn[1].t21 161.202
R22017 XThC.Tn[1].n29 XThC.Tn[1].t40 161.202
R22018 XThC.Tn[1].n25 XThC.Tn[1].t39 161.202
R22019 XThC.Tn[1].n21 XThC.Tn[1].t18 161.202
R22020 XThC.Tn[1].n17 XThC.Tn[1].t16 161.202
R22021 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R22022 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R22023 XThC.Tn[1].n69 XThC.Tn[1].t38 145.137
R22024 XThC.Tn[1].n65 XThC.Tn[1].t28 145.137
R22025 XThC.Tn[1].n61 XThC.Tn[1].t15 145.137
R22026 XThC.Tn[1].n57 XThC.Tn[1].t13 145.137
R22027 XThC.Tn[1].n53 XThC.Tn[1].t37 145.137
R22028 XThC.Tn[1].n49 XThC.Tn[1].t26 145.137
R22029 XThC.Tn[1].n45 XThC.Tn[1].t24 145.137
R22030 XThC.Tn[1].n41 XThC.Tn[1].t36 145.137
R22031 XThC.Tn[1].n37 XThC.Tn[1].t34 145.137
R22032 XThC.Tn[1].n33 XThC.Tn[1].t27 145.137
R22033 XThC.Tn[1].n29 XThC.Tn[1].t43 145.137
R22034 XThC.Tn[1].n25 XThC.Tn[1].t42 145.137
R22035 XThC.Tn[1].n21 XThC.Tn[1].t23 145.137
R22036 XThC.Tn[1].n17 XThC.Tn[1].t22 145.137
R22037 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R22038 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R22039 XThC.Tn[1].n5 XThC.Tn[1].n3 135.249
R22040 XThC.Tn[1].n5 XThC.Tn[1].n4 98.981
R22041 XThC.Tn[1].n7 XThC.Tn[1].n6 98.981
R22042 XThC.Tn[1].n9 XThC.Tn[1].n8 98.981
R22043 XThC.Tn[1].n7 XThC.Tn[1].n5 36.2672
R22044 XThC.Tn[1].n9 XThC.Tn[1].n7 36.2672
R22045 XThC.Tn[1].n74 XThC.Tn[1].n9 32.6405
R22046 XThC.Tn[1].n1 XThC.Tn[1].t1 26.5955
R22047 XThC.Tn[1].n1 XThC.Tn[1].t0 26.5955
R22048 XThC.Tn[1].n0 XThC.Tn[1].t3 26.5955
R22049 XThC.Tn[1].n0 XThC.Tn[1].t2 26.5955
R22050 XThC.Tn[1].n3 XThC.Tn[1].t11 24.9236
R22051 XThC.Tn[1].n3 XThC.Tn[1].t10 24.9236
R22052 XThC.Tn[1].n4 XThC.Tn[1].t9 24.9236
R22053 XThC.Tn[1].n4 XThC.Tn[1].t8 24.9236
R22054 XThC.Tn[1].n6 XThC.Tn[1].t7 24.9236
R22055 XThC.Tn[1].n6 XThC.Tn[1].t6 24.9236
R22056 XThC.Tn[1].n8 XThC.Tn[1].t5 24.9236
R22057 XThC.Tn[1].n8 XThC.Tn[1].t4 24.9236
R22058 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R22059 XThC.Tn[1] XThC.Tn[1].n12 8.0245
R22060 XThC.Tn[1].n72 XThC.Tn[1].n71 7.9105
R22061 XThC.Tn[1].n68 XThC.Tn[1].n67 7.9105
R22062 XThC.Tn[1].n64 XThC.Tn[1].n63 7.9105
R22063 XThC.Tn[1].n60 XThC.Tn[1].n59 7.9105
R22064 XThC.Tn[1].n56 XThC.Tn[1].n55 7.9105
R22065 XThC.Tn[1].n52 XThC.Tn[1].n51 7.9105
R22066 XThC.Tn[1].n48 XThC.Tn[1].n47 7.9105
R22067 XThC.Tn[1].n44 XThC.Tn[1].n43 7.9105
R22068 XThC.Tn[1].n40 XThC.Tn[1].n39 7.9105
R22069 XThC.Tn[1].n36 XThC.Tn[1].n35 7.9105
R22070 XThC.Tn[1].n32 XThC.Tn[1].n31 7.9105
R22071 XThC.Tn[1].n28 XThC.Tn[1].n27 7.9105
R22072 XThC.Tn[1].n24 XThC.Tn[1].n23 7.9105
R22073 XThC.Tn[1].n20 XThC.Tn[1].n19 7.9105
R22074 XThC.Tn[1].n16 XThC.Tn[1].n15 7.9105
R22075 XThC.Tn[1] XThC.Tn[1].n74 6.7205
R22076 XThC.Tn[1].n73 XThC.Tn[1] 6.08068
R22077 XThC.Tn[1].n74 XThC.Tn[1].n73 4.65249
R22078 XThC.Tn[1].n73 XThC.Tn[1] 1.8942
R22079 XThC.Tn[1].n16 XThC.Tn[1] 0.235138
R22080 XThC.Tn[1].n20 XThC.Tn[1] 0.235138
R22081 XThC.Tn[1].n24 XThC.Tn[1] 0.235138
R22082 XThC.Tn[1].n28 XThC.Tn[1] 0.235138
R22083 XThC.Tn[1].n32 XThC.Tn[1] 0.235138
R22084 XThC.Tn[1].n36 XThC.Tn[1] 0.235138
R22085 XThC.Tn[1].n40 XThC.Tn[1] 0.235138
R22086 XThC.Tn[1].n44 XThC.Tn[1] 0.235138
R22087 XThC.Tn[1].n48 XThC.Tn[1] 0.235138
R22088 XThC.Tn[1].n52 XThC.Tn[1] 0.235138
R22089 XThC.Tn[1].n56 XThC.Tn[1] 0.235138
R22090 XThC.Tn[1].n60 XThC.Tn[1] 0.235138
R22091 XThC.Tn[1].n64 XThC.Tn[1] 0.235138
R22092 XThC.Tn[1].n68 XThC.Tn[1] 0.235138
R22093 XThC.Tn[1].n72 XThC.Tn[1] 0.235138
R22094 XThC.Tn[1] XThC.Tn[1].n16 0.114505
R22095 XThC.Tn[1] XThC.Tn[1].n20 0.114505
R22096 XThC.Tn[1] XThC.Tn[1].n24 0.114505
R22097 XThC.Tn[1] XThC.Tn[1].n28 0.114505
R22098 XThC.Tn[1] XThC.Tn[1].n32 0.114505
R22099 XThC.Tn[1] XThC.Tn[1].n36 0.114505
R22100 XThC.Tn[1] XThC.Tn[1].n40 0.114505
R22101 XThC.Tn[1] XThC.Tn[1].n44 0.114505
R22102 XThC.Tn[1] XThC.Tn[1].n48 0.114505
R22103 XThC.Tn[1] XThC.Tn[1].n52 0.114505
R22104 XThC.Tn[1] XThC.Tn[1].n56 0.114505
R22105 XThC.Tn[1] XThC.Tn[1].n60 0.114505
R22106 XThC.Tn[1] XThC.Tn[1].n64 0.114505
R22107 XThC.Tn[1] XThC.Tn[1].n68 0.114505
R22108 XThC.Tn[1] XThC.Tn[1].n72 0.114505
R22109 XThC.Tn[1].n71 XThC.Tn[1].n70 0.0599512
R22110 XThC.Tn[1].n67 XThC.Tn[1].n66 0.0599512
R22111 XThC.Tn[1].n63 XThC.Tn[1].n62 0.0599512
R22112 XThC.Tn[1].n59 XThC.Tn[1].n58 0.0599512
R22113 XThC.Tn[1].n55 XThC.Tn[1].n54 0.0599512
R22114 XThC.Tn[1].n51 XThC.Tn[1].n50 0.0599512
R22115 XThC.Tn[1].n47 XThC.Tn[1].n46 0.0599512
R22116 XThC.Tn[1].n43 XThC.Tn[1].n42 0.0599512
R22117 XThC.Tn[1].n39 XThC.Tn[1].n38 0.0599512
R22118 XThC.Tn[1].n35 XThC.Tn[1].n34 0.0599512
R22119 XThC.Tn[1].n31 XThC.Tn[1].n30 0.0599512
R22120 XThC.Tn[1].n27 XThC.Tn[1].n26 0.0599512
R22121 XThC.Tn[1].n23 XThC.Tn[1].n22 0.0599512
R22122 XThC.Tn[1].n19 XThC.Tn[1].n18 0.0599512
R22123 XThC.Tn[1].n15 XThC.Tn[1].n14 0.0599512
R22124 XThC.Tn[1].n12 XThC.Tn[1].n11 0.0599512
R22125 XThC.Tn[1].n70 XThC.Tn[1] 0.0469286
R22126 XThC.Tn[1].n66 XThC.Tn[1] 0.0469286
R22127 XThC.Tn[1].n62 XThC.Tn[1] 0.0469286
R22128 XThC.Tn[1].n58 XThC.Tn[1] 0.0469286
R22129 XThC.Tn[1].n54 XThC.Tn[1] 0.0469286
R22130 XThC.Tn[1].n50 XThC.Tn[1] 0.0469286
R22131 XThC.Tn[1].n46 XThC.Tn[1] 0.0469286
R22132 XThC.Tn[1].n42 XThC.Tn[1] 0.0469286
R22133 XThC.Tn[1].n38 XThC.Tn[1] 0.0469286
R22134 XThC.Tn[1].n34 XThC.Tn[1] 0.0469286
R22135 XThC.Tn[1].n30 XThC.Tn[1] 0.0469286
R22136 XThC.Tn[1].n26 XThC.Tn[1] 0.0469286
R22137 XThC.Tn[1].n22 XThC.Tn[1] 0.0469286
R22138 XThC.Tn[1].n18 XThC.Tn[1] 0.0469286
R22139 XThC.Tn[1].n14 XThC.Tn[1] 0.0469286
R22140 XThC.Tn[1].n11 XThC.Tn[1] 0.0469286
R22141 XThC.Tn[1].n70 XThC.Tn[1] 0.0401341
R22142 XThC.Tn[1].n66 XThC.Tn[1] 0.0401341
R22143 XThC.Tn[1].n62 XThC.Tn[1] 0.0401341
R22144 XThC.Tn[1].n58 XThC.Tn[1] 0.0401341
R22145 XThC.Tn[1].n54 XThC.Tn[1] 0.0401341
R22146 XThC.Tn[1].n50 XThC.Tn[1] 0.0401341
R22147 XThC.Tn[1].n46 XThC.Tn[1] 0.0401341
R22148 XThC.Tn[1].n42 XThC.Tn[1] 0.0401341
R22149 XThC.Tn[1].n38 XThC.Tn[1] 0.0401341
R22150 XThC.Tn[1].n34 XThC.Tn[1] 0.0401341
R22151 XThC.Tn[1].n30 XThC.Tn[1] 0.0401341
R22152 XThC.Tn[1].n26 XThC.Tn[1] 0.0401341
R22153 XThC.Tn[1].n22 XThC.Tn[1] 0.0401341
R22154 XThC.Tn[1].n18 XThC.Tn[1] 0.0401341
R22155 XThC.Tn[1].n14 XThC.Tn[1] 0.0401341
R22156 XThC.Tn[1].n11 XThC.Tn[1] 0.0401341
R22157 XThC.Tn[3].n2 XThC.Tn[3].n1 332.332
R22158 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R22159 XThC.Tn[3].n71 XThC.Tn[3].n69 161.365
R22160 XThC.Tn[3].n67 XThC.Tn[3].n65 161.365
R22161 XThC.Tn[3].n63 XThC.Tn[3].n61 161.365
R22162 XThC.Tn[3].n59 XThC.Tn[3].n57 161.365
R22163 XThC.Tn[3].n55 XThC.Tn[3].n53 161.365
R22164 XThC.Tn[3].n51 XThC.Tn[3].n49 161.365
R22165 XThC.Tn[3].n47 XThC.Tn[3].n45 161.365
R22166 XThC.Tn[3].n43 XThC.Tn[3].n41 161.365
R22167 XThC.Tn[3].n39 XThC.Tn[3].n37 161.365
R22168 XThC.Tn[3].n35 XThC.Tn[3].n33 161.365
R22169 XThC.Tn[3].n31 XThC.Tn[3].n29 161.365
R22170 XThC.Tn[3].n27 XThC.Tn[3].n25 161.365
R22171 XThC.Tn[3].n23 XThC.Tn[3].n21 161.365
R22172 XThC.Tn[3].n19 XThC.Tn[3].n17 161.365
R22173 XThC.Tn[3].n15 XThC.Tn[3].n13 161.365
R22174 XThC.Tn[3].n12 XThC.Tn[3].n10 161.365
R22175 XThC.Tn[3].n69 XThC.Tn[3].t16 161.202
R22176 XThC.Tn[3].n65 XThC.Tn[3].t38 161.202
R22177 XThC.Tn[3].n61 XThC.Tn[3].t25 161.202
R22178 XThC.Tn[3].n57 XThC.Tn[3].t22 161.202
R22179 XThC.Tn[3].n53 XThC.Tn[3].t14 161.202
R22180 XThC.Tn[3].n49 XThC.Tn[3].t33 161.202
R22181 XThC.Tn[3].n45 XThC.Tn[3].t32 161.202
R22182 XThC.Tn[3].n41 XThC.Tn[3].t13 161.202
R22183 XThC.Tn[3].n37 XThC.Tn[3].t43 161.202
R22184 XThC.Tn[3].n33 XThC.Tn[3].t34 161.202
R22185 XThC.Tn[3].n29 XThC.Tn[3].t21 161.202
R22186 XThC.Tn[3].n25 XThC.Tn[3].t20 161.202
R22187 XThC.Tn[3].n21 XThC.Tn[3].t31 161.202
R22188 XThC.Tn[3].n17 XThC.Tn[3].t29 161.202
R22189 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R22190 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R22191 XThC.Tn[3].n69 XThC.Tn[3].t19 145.137
R22192 XThC.Tn[3].n65 XThC.Tn[3].t41 145.137
R22193 XThC.Tn[3].n61 XThC.Tn[3].t28 145.137
R22194 XThC.Tn[3].n57 XThC.Tn[3].t26 145.137
R22195 XThC.Tn[3].n53 XThC.Tn[3].t18 145.137
R22196 XThC.Tn[3].n49 XThC.Tn[3].t39 145.137
R22197 XThC.Tn[3].n45 XThC.Tn[3].t37 145.137
R22198 XThC.Tn[3].n41 XThC.Tn[3].t17 145.137
R22199 XThC.Tn[3].n37 XThC.Tn[3].t15 145.137
R22200 XThC.Tn[3].n33 XThC.Tn[3].t40 145.137
R22201 XThC.Tn[3].n29 XThC.Tn[3].t24 145.137
R22202 XThC.Tn[3].n25 XThC.Tn[3].t23 145.137
R22203 XThC.Tn[3].n21 XThC.Tn[3].t36 145.137
R22204 XThC.Tn[3].n17 XThC.Tn[3].t35 145.137
R22205 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R22206 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R22207 XThC.Tn[3].n6 XThC.Tn[3].n4 135.249
R22208 XThC.Tn[3].n9 XThC.Tn[3].n3 98.981
R22209 XThC.Tn[3].n6 XThC.Tn[3].n5 98.981
R22210 XThC.Tn[3].n8 XThC.Tn[3].n7 98.981
R22211 XThC.Tn[3].n8 XThC.Tn[3].n6 36.2672
R22212 XThC.Tn[3].n9 XThC.Tn[3].n8 36.2672
R22213 XThC.Tn[3].n74 XThC.Tn[3].n9 32.6405
R22214 XThC.Tn[3].n1 XThC.Tn[3].t7 26.5955
R22215 XThC.Tn[3].n1 XThC.Tn[3].t6 26.5955
R22216 XThC.Tn[3].n0 XThC.Tn[3].t5 26.5955
R22217 XThC.Tn[3].n0 XThC.Tn[3].t4 26.5955
R22218 XThC.Tn[3].n3 XThC.Tn[3].t1 24.9236
R22219 XThC.Tn[3].n3 XThC.Tn[3].t0 24.9236
R22220 XThC.Tn[3].n4 XThC.Tn[3].t11 24.9236
R22221 XThC.Tn[3].n4 XThC.Tn[3].t10 24.9236
R22222 XThC.Tn[3].n5 XThC.Tn[3].t9 24.9236
R22223 XThC.Tn[3].n5 XThC.Tn[3].t8 24.9236
R22224 XThC.Tn[3].n7 XThC.Tn[3].t3 24.9236
R22225 XThC.Tn[3].n7 XThC.Tn[3].t2 24.9236
R22226 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R22227 XThC.Tn[3] XThC.Tn[3].n12 8.0245
R22228 XThC.Tn[3].n72 XThC.Tn[3].n71 7.9105
R22229 XThC.Tn[3].n68 XThC.Tn[3].n67 7.9105
R22230 XThC.Tn[3].n64 XThC.Tn[3].n63 7.9105
R22231 XThC.Tn[3].n60 XThC.Tn[3].n59 7.9105
R22232 XThC.Tn[3].n56 XThC.Tn[3].n55 7.9105
R22233 XThC.Tn[3].n52 XThC.Tn[3].n51 7.9105
R22234 XThC.Tn[3].n48 XThC.Tn[3].n47 7.9105
R22235 XThC.Tn[3].n44 XThC.Tn[3].n43 7.9105
R22236 XThC.Tn[3].n40 XThC.Tn[3].n39 7.9105
R22237 XThC.Tn[3].n36 XThC.Tn[3].n35 7.9105
R22238 XThC.Tn[3].n32 XThC.Tn[3].n31 7.9105
R22239 XThC.Tn[3].n28 XThC.Tn[3].n27 7.9105
R22240 XThC.Tn[3].n24 XThC.Tn[3].n23 7.9105
R22241 XThC.Tn[3].n20 XThC.Tn[3].n19 7.9105
R22242 XThC.Tn[3].n16 XThC.Tn[3].n15 7.9105
R22243 XThC.Tn[3].n73 XThC.Tn[3] 7.48718
R22244 XThC.Tn[3] XThC.Tn[3].n74 6.7205
R22245 XThC.Tn[3].n74 XThC.Tn[3].n73 5.06464
R22246 XThC.Tn[3].n73 XThC.Tn[3] 1.18175
R22247 XThC.Tn[3].n16 XThC.Tn[3] 0.235138
R22248 XThC.Tn[3].n20 XThC.Tn[3] 0.235138
R22249 XThC.Tn[3].n24 XThC.Tn[3] 0.235138
R22250 XThC.Tn[3].n28 XThC.Tn[3] 0.235138
R22251 XThC.Tn[3].n32 XThC.Tn[3] 0.235138
R22252 XThC.Tn[3].n36 XThC.Tn[3] 0.235138
R22253 XThC.Tn[3].n40 XThC.Tn[3] 0.235138
R22254 XThC.Tn[3].n44 XThC.Tn[3] 0.235138
R22255 XThC.Tn[3].n48 XThC.Tn[3] 0.235138
R22256 XThC.Tn[3].n52 XThC.Tn[3] 0.235138
R22257 XThC.Tn[3].n56 XThC.Tn[3] 0.235138
R22258 XThC.Tn[3].n60 XThC.Tn[3] 0.235138
R22259 XThC.Tn[3].n64 XThC.Tn[3] 0.235138
R22260 XThC.Tn[3].n68 XThC.Tn[3] 0.235138
R22261 XThC.Tn[3].n72 XThC.Tn[3] 0.235138
R22262 XThC.Tn[3] XThC.Tn[3].n16 0.114505
R22263 XThC.Tn[3] XThC.Tn[3].n20 0.114505
R22264 XThC.Tn[3] XThC.Tn[3].n24 0.114505
R22265 XThC.Tn[3] XThC.Tn[3].n28 0.114505
R22266 XThC.Tn[3] XThC.Tn[3].n32 0.114505
R22267 XThC.Tn[3] XThC.Tn[3].n36 0.114505
R22268 XThC.Tn[3] XThC.Tn[3].n40 0.114505
R22269 XThC.Tn[3] XThC.Tn[3].n44 0.114505
R22270 XThC.Tn[3] XThC.Tn[3].n48 0.114505
R22271 XThC.Tn[3] XThC.Tn[3].n52 0.114505
R22272 XThC.Tn[3] XThC.Tn[3].n56 0.114505
R22273 XThC.Tn[3] XThC.Tn[3].n60 0.114505
R22274 XThC.Tn[3] XThC.Tn[3].n64 0.114505
R22275 XThC.Tn[3] XThC.Tn[3].n68 0.114505
R22276 XThC.Tn[3] XThC.Tn[3].n72 0.114505
R22277 XThC.Tn[3].n71 XThC.Tn[3].n70 0.0599512
R22278 XThC.Tn[3].n67 XThC.Tn[3].n66 0.0599512
R22279 XThC.Tn[3].n63 XThC.Tn[3].n62 0.0599512
R22280 XThC.Tn[3].n59 XThC.Tn[3].n58 0.0599512
R22281 XThC.Tn[3].n55 XThC.Tn[3].n54 0.0599512
R22282 XThC.Tn[3].n51 XThC.Tn[3].n50 0.0599512
R22283 XThC.Tn[3].n47 XThC.Tn[3].n46 0.0599512
R22284 XThC.Tn[3].n43 XThC.Tn[3].n42 0.0599512
R22285 XThC.Tn[3].n39 XThC.Tn[3].n38 0.0599512
R22286 XThC.Tn[3].n35 XThC.Tn[3].n34 0.0599512
R22287 XThC.Tn[3].n31 XThC.Tn[3].n30 0.0599512
R22288 XThC.Tn[3].n27 XThC.Tn[3].n26 0.0599512
R22289 XThC.Tn[3].n23 XThC.Tn[3].n22 0.0599512
R22290 XThC.Tn[3].n19 XThC.Tn[3].n18 0.0599512
R22291 XThC.Tn[3].n15 XThC.Tn[3].n14 0.0599512
R22292 XThC.Tn[3].n12 XThC.Tn[3].n11 0.0599512
R22293 XThC.Tn[3].n70 XThC.Tn[3] 0.0469286
R22294 XThC.Tn[3].n66 XThC.Tn[3] 0.0469286
R22295 XThC.Tn[3].n62 XThC.Tn[3] 0.0469286
R22296 XThC.Tn[3].n58 XThC.Tn[3] 0.0469286
R22297 XThC.Tn[3].n54 XThC.Tn[3] 0.0469286
R22298 XThC.Tn[3].n50 XThC.Tn[3] 0.0469286
R22299 XThC.Tn[3].n46 XThC.Tn[3] 0.0469286
R22300 XThC.Tn[3].n42 XThC.Tn[3] 0.0469286
R22301 XThC.Tn[3].n38 XThC.Tn[3] 0.0469286
R22302 XThC.Tn[3].n34 XThC.Tn[3] 0.0469286
R22303 XThC.Tn[3].n30 XThC.Tn[3] 0.0469286
R22304 XThC.Tn[3].n26 XThC.Tn[3] 0.0469286
R22305 XThC.Tn[3].n22 XThC.Tn[3] 0.0469286
R22306 XThC.Tn[3].n18 XThC.Tn[3] 0.0469286
R22307 XThC.Tn[3].n14 XThC.Tn[3] 0.0469286
R22308 XThC.Tn[3].n11 XThC.Tn[3] 0.0469286
R22309 XThC.Tn[3].n70 XThC.Tn[3] 0.0401341
R22310 XThC.Tn[3].n66 XThC.Tn[3] 0.0401341
R22311 XThC.Tn[3].n62 XThC.Tn[3] 0.0401341
R22312 XThC.Tn[3].n58 XThC.Tn[3] 0.0401341
R22313 XThC.Tn[3].n54 XThC.Tn[3] 0.0401341
R22314 XThC.Tn[3].n50 XThC.Tn[3] 0.0401341
R22315 XThC.Tn[3].n46 XThC.Tn[3] 0.0401341
R22316 XThC.Tn[3].n42 XThC.Tn[3] 0.0401341
R22317 XThC.Tn[3].n38 XThC.Tn[3] 0.0401341
R22318 XThC.Tn[3].n34 XThC.Tn[3] 0.0401341
R22319 XThC.Tn[3].n30 XThC.Tn[3] 0.0401341
R22320 XThC.Tn[3].n26 XThC.Tn[3] 0.0401341
R22321 XThC.Tn[3].n22 XThC.Tn[3] 0.0401341
R22322 XThC.Tn[3].n18 XThC.Tn[3] 0.0401341
R22323 XThC.Tn[3].n14 XThC.Tn[3] 0.0401341
R22324 XThC.Tn[3].n11 XThC.Tn[3] 0.0401341
R22325 XThR.Tn[10].n5 XThR.Tn[10].n4 256.103
R22326 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R22327 XThR.Tn[10].n88 XThR.Tn[10].n86 241.847
R22328 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R22329 XThR.Tn[10].n5 XThR.Tn[10].n3 202.095
R22330 XThR.Tn[10].n88 XThR.Tn[10].n87 185
R22331 XThR.Tn[10] XThR.Tn[10].n79 161.363
R22332 XThR.Tn[10] XThR.Tn[10].n74 161.363
R22333 XThR.Tn[10] XThR.Tn[10].n69 161.363
R22334 XThR.Tn[10] XThR.Tn[10].n64 161.363
R22335 XThR.Tn[10] XThR.Tn[10].n59 161.363
R22336 XThR.Tn[10] XThR.Tn[10].n54 161.363
R22337 XThR.Tn[10] XThR.Tn[10].n49 161.363
R22338 XThR.Tn[10] XThR.Tn[10].n44 161.363
R22339 XThR.Tn[10] XThR.Tn[10].n39 161.363
R22340 XThR.Tn[10] XThR.Tn[10].n34 161.363
R22341 XThR.Tn[10] XThR.Tn[10].n29 161.363
R22342 XThR.Tn[10] XThR.Tn[10].n24 161.363
R22343 XThR.Tn[10] XThR.Tn[10].n19 161.363
R22344 XThR.Tn[10] XThR.Tn[10].n14 161.363
R22345 XThR.Tn[10] XThR.Tn[10].n9 161.363
R22346 XThR.Tn[10] XThR.Tn[10].n7 161.363
R22347 XThR.Tn[10].n81 XThR.Tn[10].n80 161.3
R22348 XThR.Tn[10].n76 XThR.Tn[10].n75 161.3
R22349 XThR.Tn[10].n71 XThR.Tn[10].n70 161.3
R22350 XThR.Tn[10].n66 XThR.Tn[10].n65 161.3
R22351 XThR.Tn[10].n61 XThR.Tn[10].n60 161.3
R22352 XThR.Tn[10].n56 XThR.Tn[10].n55 161.3
R22353 XThR.Tn[10].n51 XThR.Tn[10].n50 161.3
R22354 XThR.Tn[10].n46 XThR.Tn[10].n45 161.3
R22355 XThR.Tn[10].n41 XThR.Tn[10].n40 161.3
R22356 XThR.Tn[10].n36 XThR.Tn[10].n35 161.3
R22357 XThR.Tn[10].n31 XThR.Tn[10].n30 161.3
R22358 XThR.Tn[10].n26 XThR.Tn[10].n25 161.3
R22359 XThR.Tn[10].n21 XThR.Tn[10].n20 161.3
R22360 XThR.Tn[10].n16 XThR.Tn[10].n15 161.3
R22361 XThR.Tn[10].n11 XThR.Tn[10].n10 161.3
R22362 XThR.Tn[10].n79 XThR.Tn[10].t37 161.106
R22363 XThR.Tn[10].n74 XThR.Tn[10].t45 161.106
R22364 XThR.Tn[10].n69 XThR.Tn[10].t27 161.106
R22365 XThR.Tn[10].n64 XThR.Tn[10].t72 161.106
R22366 XThR.Tn[10].n59 XThR.Tn[10].t35 161.106
R22367 XThR.Tn[10].n54 XThR.Tn[10].t61 161.106
R22368 XThR.Tn[10].n49 XThR.Tn[10].t43 161.106
R22369 XThR.Tn[10].n44 XThR.Tn[10].t24 161.106
R22370 XThR.Tn[10].n39 XThR.Tn[10].t69 161.106
R22371 XThR.Tn[10].n34 XThR.Tn[10].t15 161.106
R22372 XThR.Tn[10].n29 XThR.Tn[10].t59 161.106
R22373 XThR.Tn[10].n24 XThR.Tn[10].t26 161.106
R22374 XThR.Tn[10].n19 XThR.Tn[10].t58 161.106
R22375 XThR.Tn[10].n14 XThR.Tn[10].t41 161.106
R22376 XThR.Tn[10].n9 XThR.Tn[10].t63 161.106
R22377 XThR.Tn[10].n7 XThR.Tn[10].t47 161.106
R22378 XThR.Tn[10].n80 XThR.Tn[10].t34 159.978
R22379 XThR.Tn[10].n75 XThR.Tn[10].t39 159.978
R22380 XThR.Tn[10].n70 XThR.Tn[10].t22 159.978
R22381 XThR.Tn[10].n65 XThR.Tn[10].t68 159.978
R22382 XThR.Tn[10].n60 XThR.Tn[10].t32 159.978
R22383 XThR.Tn[10].n55 XThR.Tn[10].t57 159.978
R22384 XThR.Tn[10].n50 XThR.Tn[10].t38 159.978
R22385 XThR.Tn[10].n45 XThR.Tn[10].t20 159.978
R22386 XThR.Tn[10].n40 XThR.Tn[10].t66 159.978
R22387 XThR.Tn[10].n35 XThR.Tn[10].t12 159.978
R22388 XThR.Tn[10].n30 XThR.Tn[10].t56 159.978
R22389 XThR.Tn[10].n25 XThR.Tn[10].t21 159.978
R22390 XThR.Tn[10].n20 XThR.Tn[10].t55 159.978
R22391 XThR.Tn[10].n15 XThR.Tn[10].t36 159.978
R22392 XThR.Tn[10].n10 XThR.Tn[10].t60 159.978
R22393 XThR.Tn[10].n79 XThR.Tn[10].t29 145.038
R22394 XThR.Tn[10].n74 XThR.Tn[10].t49 145.038
R22395 XThR.Tn[10].n69 XThR.Tn[10].t31 145.038
R22396 XThR.Tn[10].n64 XThR.Tn[10].t16 145.038
R22397 XThR.Tn[10].n59 XThR.Tn[10].t46 145.038
R22398 XThR.Tn[10].n54 XThR.Tn[10].t28 145.038
R22399 XThR.Tn[10].n49 XThR.Tn[10].t33 145.038
R22400 XThR.Tn[10].n44 XThR.Tn[10].t17 145.038
R22401 XThR.Tn[10].n39 XThR.Tn[10].t14 145.038
R22402 XThR.Tn[10].n34 XThR.Tn[10].t44 145.038
R22403 XThR.Tn[10].n29 XThR.Tn[10].t67 145.038
R22404 XThR.Tn[10].n24 XThR.Tn[10].t30 145.038
R22405 XThR.Tn[10].n19 XThR.Tn[10].t65 145.038
R22406 XThR.Tn[10].n14 XThR.Tn[10].t48 145.038
R22407 XThR.Tn[10].n9 XThR.Tn[10].t13 145.038
R22408 XThR.Tn[10].n7 XThR.Tn[10].t54 145.038
R22409 XThR.Tn[10].n80 XThR.Tn[10].t64 143.911
R22410 XThR.Tn[10].n75 XThR.Tn[10].t25 143.911
R22411 XThR.Tn[10].n70 XThR.Tn[10].t71 143.911
R22412 XThR.Tn[10].n65 XThR.Tn[10].t52 143.911
R22413 XThR.Tn[10].n60 XThR.Tn[10].t19 143.911
R22414 XThR.Tn[10].n55 XThR.Tn[10].t62 143.911
R22415 XThR.Tn[10].n50 XThR.Tn[10].t73 143.911
R22416 XThR.Tn[10].n45 XThR.Tn[10].t53 143.911
R22417 XThR.Tn[10].n40 XThR.Tn[10].t51 143.911
R22418 XThR.Tn[10].n35 XThR.Tn[10].t18 143.911
R22419 XThR.Tn[10].n30 XThR.Tn[10].t42 143.911
R22420 XThR.Tn[10].n25 XThR.Tn[10].t70 143.911
R22421 XThR.Tn[10].n20 XThR.Tn[10].t40 143.911
R22422 XThR.Tn[10].n15 XThR.Tn[10].t23 143.911
R22423 XThR.Tn[10].n10 XThR.Tn[10].t50 143.911
R22424 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R22425 XThR.Tn[10].n3 XThR.Tn[10].t3 26.5955
R22426 XThR.Tn[10].n3 XThR.Tn[10].t8 26.5955
R22427 XThR.Tn[10].n4 XThR.Tn[10].t10 26.5955
R22428 XThR.Tn[10].n4 XThR.Tn[10].t1 26.5955
R22429 XThR.Tn[10].n0 XThR.Tn[10].t6 26.5955
R22430 XThR.Tn[10].n0 XThR.Tn[10].t4 26.5955
R22431 XThR.Tn[10].n1 XThR.Tn[10].t7 26.5955
R22432 XThR.Tn[10].n1 XThR.Tn[10].t5 26.5955
R22433 XThR.Tn[10].n86 XThR.Tn[10].t2 24.9236
R22434 XThR.Tn[10].n86 XThR.Tn[10].t11 24.9236
R22435 XThR.Tn[10].n87 XThR.Tn[10].t9 24.9236
R22436 XThR.Tn[10].n87 XThR.Tn[10].t0 24.9236
R22437 XThR.Tn[10] XThR.Tn[10].n88 18.8943
R22438 XThR.Tn[10].n6 XThR.Tn[10].n5 13.5534
R22439 XThR.Tn[10].n85 XThR.Tn[10] 7.84567
R22440 XThR.Tn[10] XThR.Tn[10].n85 6.34069
R22441 XThR.Tn[10] XThR.Tn[10].n8 5.34038
R22442 XThR.Tn[10].n13 XThR.Tn[10].n12 4.5005
R22443 XThR.Tn[10].n18 XThR.Tn[10].n17 4.5005
R22444 XThR.Tn[10].n23 XThR.Tn[10].n22 4.5005
R22445 XThR.Tn[10].n28 XThR.Tn[10].n27 4.5005
R22446 XThR.Tn[10].n33 XThR.Tn[10].n32 4.5005
R22447 XThR.Tn[10].n38 XThR.Tn[10].n37 4.5005
R22448 XThR.Tn[10].n43 XThR.Tn[10].n42 4.5005
R22449 XThR.Tn[10].n48 XThR.Tn[10].n47 4.5005
R22450 XThR.Tn[10].n53 XThR.Tn[10].n52 4.5005
R22451 XThR.Tn[10].n58 XThR.Tn[10].n57 4.5005
R22452 XThR.Tn[10].n63 XThR.Tn[10].n62 4.5005
R22453 XThR.Tn[10].n68 XThR.Tn[10].n67 4.5005
R22454 XThR.Tn[10].n73 XThR.Tn[10].n72 4.5005
R22455 XThR.Tn[10].n78 XThR.Tn[10].n77 4.5005
R22456 XThR.Tn[10].n83 XThR.Tn[10].n82 4.5005
R22457 XThR.Tn[10].n84 XThR.Tn[10] 3.70586
R22458 XThR.Tn[10].n13 XThR.Tn[10] 2.52282
R22459 XThR.Tn[10].n18 XThR.Tn[10] 2.52282
R22460 XThR.Tn[10].n23 XThR.Tn[10] 2.52282
R22461 XThR.Tn[10].n28 XThR.Tn[10] 2.52282
R22462 XThR.Tn[10].n33 XThR.Tn[10] 2.52282
R22463 XThR.Tn[10].n38 XThR.Tn[10] 2.52282
R22464 XThR.Tn[10].n43 XThR.Tn[10] 2.52282
R22465 XThR.Tn[10].n48 XThR.Tn[10] 2.52282
R22466 XThR.Tn[10].n53 XThR.Tn[10] 2.52282
R22467 XThR.Tn[10].n58 XThR.Tn[10] 2.52282
R22468 XThR.Tn[10].n63 XThR.Tn[10] 2.52282
R22469 XThR.Tn[10].n68 XThR.Tn[10] 2.52282
R22470 XThR.Tn[10].n73 XThR.Tn[10] 2.52282
R22471 XThR.Tn[10].n78 XThR.Tn[10] 2.52282
R22472 XThR.Tn[10].n83 XThR.Tn[10] 2.52282
R22473 XThR.Tn[10].n85 XThR.Tn[10] 1.79489
R22474 XThR.Tn[10].n6 XThR.Tn[10] 1.50638
R22475 XThR.Tn[10] XThR.Tn[10].n6 1.19676
R22476 XThR.Tn[10].n81 XThR.Tn[10] 1.08677
R22477 XThR.Tn[10].n76 XThR.Tn[10] 1.08677
R22478 XThR.Tn[10].n71 XThR.Tn[10] 1.08677
R22479 XThR.Tn[10].n66 XThR.Tn[10] 1.08677
R22480 XThR.Tn[10].n61 XThR.Tn[10] 1.08677
R22481 XThR.Tn[10].n56 XThR.Tn[10] 1.08677
R22482 XThR.Tn[10].n51 XThR.Tn[10] 1.08677
R22483 XThR.Tn[10].n46 XThR.Tn[10] 1.08677
R22484 XThR.Tn[10].n41 XThR.Tn[10] 1.08677
R22485 XThR.Tn[10].n36 XThR.Tn[10] 1.08677
R22486 XThR.Tn[10].n31 XThR.Tn[10] 1.08677
R22487 XThR.Tn[10].n26 XThR.Tn[10] 1.08677
R22488 XThR.Tn[10].n21 XThR.Tn[10] 1.08677
R22489 XThR.Tn[10].n16 XThR.Tn[10] 1.08677
R22490 XThR.Tn[10].n11 XThR.Tn[10] 1.08677
R22491 XThR.Tn[10] XThR.Tn[10].n13 0.839786
R22492 XThR.Tn[10] XThR.Tn[10].n18 0.839786
R22493 XThR.Tn[10] XThR.Tn[10].n23 0.839786
R22494 XThR.Tn[10] XThR.Tn[10].n28 0.839786
R22495 XThR.Tn[10] XThR.Tn[10].n33 0.839786
R22496 XThR.Tn[10] XThR.Tn[10].n38 0.839786
R22497 XThR.Tn[10] XThR.Tn[10].n43 0.839786
R22498 XThR.Tn[10] XThR.Tn[10].n48 0.839786
R22499 XThR.Tn[10] XThR.Tn[10].n53 0.839786
R22500 XThR.Tn[10] XThR.Tn[10].n58 0.839786
R22501 XThR.Tn[10] XThR.Tn[10].n63 0.839786
R22502 XThR.Tn[10] XThR.Tn[10].n68 0.839786
R22503 XThR.Tn[10] XThR.Tn[10].n73 0.839786
R22504 XThR.Tn[10] XThR.Tn[10].n78 0.839786
R22505 XThR.Tn[10] XThR.Tn[10].n83 0.839786
R22506 XThR.Tn[10].n8 XThR.Tn[10] 0.499542
R22507 XThR.Tn[10].n82 XThR.Tn[10] 0.063
R22508 XThR.Tn[10].n77 XThR.Tn[10] 0.063
R22509 XThR.Tn[10].n72 XThR.Tn[10] 0.063
R22510 XThR.Tn[10].n67 XThR.Tn[10] 0.063
R22511 XThR.Tn[10].n62 XThR.Tn[10] 0.063
R22512 XThR.Tn[10].n57 XThR.Tn[10] 0.063
R22513 XThR.Tn[10].n52 XThR.Tn[10] 0.063
R22514 XThR.Tn[10].n47 XThR.Tn[10] 0.063
R22515 XThR.Tn[10].n42 XThR.Tn[10] 0.063
R22516 XThR.Tn[10].n37 XThR.Tn[10] 0.063
R22517 XThR.Tn[10].n32 XThR.Tn[10] 0.063
R22518 XThR.Tn[10].n27 XThR.Tn[10] 0.063
R22519 XThR.Tn[10].n22 XThR.Tn[10] 0.063
R22520 XThR.Tn[10].n17 XThR.Tn[10] 0.063
R22521 XThR.Tn[10].n12 XThR.Tn[10] 0.063
R22522 XThR.Tn[10].n84 XThR.Tn[10] 0.0540714
R22523 XThR.Tn[10] XThR.Tn[10].n84 0.038
R22524 XThR.Tn[10].n8 XThR.Tn[10] 0.0143889
R22525 XThR.Tn[10].n82 XThR.Tn[10].n81 0.00771154
R22526 XThR.Tn[10].n77 XThR.Tn[10].n76 0.00771154
R22527 XThR.Tn[10].n72 XThR.Tn[10].n71 0.00771154
R22528 XThR.Tn[10].n67 XThR.Tn[10].n66 0.00771154
R22529 XThR.Tn[10].n62 XThR.Tn[10].n61 0.00771154
R22530 XThR.Tn[10].n57 XThR.Tn[10].n56 0.00771154
R22531 XThR.Tn[10].n52 XThR.Tn[10].n51 0.00771154
R22532 XThR.Tn[10].n47 XThR.Tn[10].n46 0.00771154
R22533 XThR.Tn[10].n42 XThR.Tn[10].n41 0.00771154
R22534 XThR.Tn[10].n37 XThR.Tn[10].n36 0.00771154
R22535 XThR.Tn[10].n32 XThR.Tn[10].n31 0.00771154
R22536 XThR.Tn[10].n27 XThR.Tn[10].n26 0.00771154
R22537 XThR.Tn[10].n22 XThR.Tn[10].n21 0.00771154
R22538 XThR.Tn[10].n17 XThR.Tn[10].n16 0.00771154
R22539 XThR.Tn[10].n12 XThR.Tn[10].n11 0.00771154
R22540 XThC.Tn[14].n70 XThC.Tn[14].n69 256.104
R22541 XThC.Tn[14].n74 XThC.Tn[14].n73 243.679
R22542 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22543 XThC.Tn[14].n74 XThC.Tn[14].n72 205.28
R22544 XThC.Tn[14].n70 XThC.Tn[14].n68 202.095
R22545 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22546 XThC.Tn[14].n64 XThC.Tn[14].n62 161.365
R22547 XThC.Tn[14].n60 XThC.Tn[14].n58 161.365
R22548 XThC.Tn[14].n56 XThC.Tn[14].n54 161.365
R22549 XThC.Tn[14].n52 XThC.Tn[14].n50 161.365
R22550 XThC.Tn[14].n48 XThC.Tn[14].n46 161.365
R22551 XThC.Tn[14].n44 XThC.Tn[14].n42 161.365
R22552 XThC.Tn[14].n40 XThC.Tn[14].n38 161.365
R22553 XThC.Tn[14].n36 XThC.Tn[14].n34 161.365
R22554 XThC.Tn[14].n32 XThC.Tn[14].n30 161.365
R22555 XThC.Tn[14].n28 XThC.Tn[14].n26 161.365
R22556 XThC.Tn[14].n24 XThC.Tn[14].n22 161.365
R22557 XThC.Tn[14].n20 XThC.Tn[14].n18 161.365
R22558 XThC.Tn[14].n16 XThC.Tn[14].n14 161.365
R22559 XThC.Tn[14].n12 XThC.Tn[14].n10 161.365
R22560 XThC.Tn[14].n8 XThC.Tn[14].n6 161.365
R22561 XThC.Tn[14].n5 XThC.Tn[14].n3 161.365
R22562 XThC.Tn[14].n62 XThC.Tn[14].t12 161.202
R22563 XThC.Tn[14].n58 XThC.Tn[14].t33 161.202
R22564 XThC.Tn[14].n54 XThC.Tn[14].t21 161.202
R22565 XThC.Tn[14].n50 XThC.Tn[14].t19 161.202
R22566 XThC.Tn[14].n46 XThC.Tn[14].t42 161.202
R22567 XThC.Tn[14].n42 XThC.Tn[14].t30 161.202
R22568 XThC.Tn[14].n38 XThC.Tn[14].t27 161.202
R22569 XThC.Tn[14].n34 XThC.Tn[14].t41 161.202
R22570 XThC.Tn[14].n30 XThC.Tn[14].t39 161.202
R22571 XThC.Tn[14].n26 XThC.Tn[14].t31 161.202
R22572 XThC.Tn[14].n22 XThC.Tn[14].t17 161.202
R22573 XThC.Tn[14].n18 XThC.Tn[14].t14 161.202
R22574 XThC.Tn[14].n14 XThC.Tn[14].t26 161.202
R22575 XThC.Tn[14].n10 XThC.Tn[14].t25 161.202
R22576 XThC.Tn[14].n6 XThC.Tn[14].t22 161.202
R22577 XThC.Tn[14].n3 XThC.Tn[14].t38 161.202
R22578 XThC.Tn[14].n62 XThC.Tn[14].t18 145.137
R22579 XThC.Tn[14].n58 XThC.Tn[14].t40 145.137
R22580 XThC.Tn[14].n54 XThC.Tn[14].t28 145.137
R22581 XThC.Tn[14].n50 XThC.Tn[14].t24 145.137
R22582 XThC.Tn[14].n46 XThC.Tn[14].t16 145.137
R22583 XThC.Tn[14].n42 XThC.Tn[14].t36 145.137
R22584 XThC.Tn[14].n38 XThC.Tn[14].t35 145.137
R22585 XThC.Tn[14].n34 XThC.Tn[14].t15 145.137
R22586 XThC.Tn[14].n30 XThC.Tn[14].t13 145.137
R22587 XThC.Tn[14].n26 XThC.Tn[14].t37 145.137
R22588 XThC.Tn[14].n22 XThC.Tn[14].t23 145.137
R22589 XThC.Tn[14].n18 XThC.Tn[14].t20 145.137
R22590 XThC.Tn[14].n14 XThC.Tn[14].t34 145.137
R22591 XThC.Tn[14].n10 XThC.Tn[14].t32 145.137
R22592 XThC.Tn[14].n6 XThC.Tn[14].t29 145.137
R22593 XThC.Tn[14].n3 XThC.Tn[14].t43 145.137
R22594 XThC.Tn[14].n68 XThC.Tn[14].t8 26.5955
R22595 XThC.Tn[14].n68 XThC.Tn[14].t9 26.5955
R22596 XThC.Tn[14].n69 XThC.Tn[14].t11 26.5955
R22597 XThC.Tn[14].n69 XThC.Tn[14].t10 26.5955
R22598 XThC.Tn[14].n72 XThC.Tn[14].t1 26.5955
R22599 XThC.Tn[14].n72 XThC.Tn[14].t0 26.5955
R22600 XThC.Tn[14].n73 XThC.Tn[14].t3 26.5955
R22601 XThC.Tn[14].n73 XThC.Tn[14].t2 26.5955
R22602 XThC.Tn[14].n1 XThC.Tn[14].t5 24.9236
R22603 XThC.Tn[14].n1 XThC.Tn[14].t7 24.9236
R22604 XThC.Tn[14].n0 XThC.Tn[14].t4 24.9236
R22605 XThC.Tn[14].n0 XThC.Tn[14].t6 24.9236
R22606 XThC.Tn[14] XThC.Tn[14].n74 22.9652
R22607 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22608 XThC.Tn[14].n71 XThC.Tn[14].n70 13.9299
R22609 XThC.Tn[14] XThC.Tn[14].n71 13.9299
R22610 XThC.Tn[14] XThC.Tn[14].n5 8.0245
R22611 XThC.Tn[14].n65 XThC.Tn[14].n64 7.9105
R22612 XThC.Tn[14].n61 XThC.Tn[14].n60 7.9105
R22613 XThC.Tn[14].n57 XThC.Tn[14].n56 7.9105
R22614 XThC.Tn[14].n53 XThC.Tn[14].n52 7.9105
R22615 XThC.Tn[14].n49 XThC.Tn[14].n48 7.9105
R22616 XThC.Tn[14].n45 XThC.Tn[14].n44 7.9105
R22617 XThC.Tn[14].n41 XThC.Tn[14].n40 7.9105
R22618 XThC.Tn[14].n37 XThC.Tn[14].n36 7.9105
R22619 XThC.Tn[14].n33 XThC.Tn[14].n32 7.9105
R22620 XThC.Tn[14].n29 XThC.Tn[14].n28 7.9105
R22621 XThC.Tn[14].n25 XThC.Tn[14].n24 7.9105
R22622 XThC.Tn[14].n21 XThC.Tn[14].n20 7.9105
R22623 XThC.Tn[14].n17 XThC.Tn[14].n16 7.9105
R22624 XThC.Tn[14].n13 XThC.Tn[14].n12 7.9105
R22625 XThC.Tn[14].n9 XThC.Tn[14].n8 7.9105
R22626 XThC.Tn[14].n67 XThC.Tn[14].n66 7.51947
R22627 XThC.Tn[14].n66 XThC.Tn[14] 5.85107
R22628 XThC.Tn[14].n71 XThC.Tn[14].n67 2.99115
R22629 XThC.Tn[14].n71 XThC.Tn[14] 2.87153
R22630 XThC.Tn[14].n67 XThC.Tn[14] 2.2734
R22631 XThC.Tn[14].n66 XThC.Tn[14] 1.06164
R22632 XThC.Tn[14].n9 XThC.Tn[14] 0.235138
R22633 XThC.Tn[14].n13 XThC.Tn[14] 0.235138
R22634 XThC.Tn[14].n17 XThC.Tn[14] 0.235138
R22635 XThC.Tn[14].n21 XThC.Tn[14] 0.235138
R22636 XThC.Tn[14].n25 XThC.Tn[14] 0.235138
R22637 XThC.Tn[14].n29 XThC.Tn[14] 0.235138
R22638 XThC.Tn[14].n33 XThC.Tn[14] 0.235138
R22639 XThC.Tn[14].n37 XThC.Tn[14] 0.235138
R22640 XThC.Tn[14].n41 XThC.Tn[14] 0.235138
R22641 XThC.Tn[14].n45 XThC.Tn[14] 0.235138
R22642 XThC.Tn[14].n49 XThC.Tn[14] 0.235138
R22643 XThC.Tn[14].n53 XThC.Tn[14] 0.235138
R22644 XThC.Tn[14].n57 XThC.Tn[14] 0.235138
R22645 XThC.Tn[14].n61 XThC.Tn[14] 0.235138
R22646 XThC.Tn[14].n65 XThC.Tn[14] 0.235138
R22647 XThC.Tn[14] XThC.Tn[14].n9 0.114505
R22648 XThC.Tn[14] XThC.Tn[14].n13 0.114505
R22649 XThC.Tn[14] XThC.Tn[14].n17 0.114505
R22650 XThC.Tn[14] XThC.Tn[14].n21 0.114505
R22651 XThC.Tn[14] XThC.Tn[14].n25 0.114505
R22652 XThC.Tn[14] XThC.Tn[14].n29 0.114505
R22653 XThC.Tn[14] XThC.Tn[14].n33 0.114505
R22654 XThC.Tn[14] XThC.Tn[14].n37 0.114505
R22655 XThC.Tn[14] XThC.Tn[14].n41 0.114505
R22656 XThC.Tn[14] XThC.Tn[14].n45 0.114505
R22657 XThC.Tn[14] XThC.Tn[14].n49 0.114505
R22658 XThC.Tn[14] XThC.Tn[14].n53 0.114505
R22659 XThC.Tn[14] XThC.Tn[14].n57 0.114505
R22660 XThC.Tn[14] XThC.Tn[14].n61 0.114505
R22661 XThC.Tn[14] XThC.Tn[14].n65 0.114505
R22662 XThC.Tn[14].n64 XThC.Tn[14].n63 0.0599512
R22663 XThC.Tn[14].n60 XThC.Tn[14].n59 0.0599512
R22664 XThC.Tn[14].n56 XThC.Tn[14].n55 0.0599512
R22665 XThC.Tn[14].n52 XThC.Tn[14].n51 0.0599512
R22666 XThC.Tn[14].n48 XThC.Tn[14].n47 0.0599512
R22667 XThC.Tn[14].n44 XThC.Tn[14].n43 0.0599512
R22668 XThC.Tn[14].n40 XThC.Tn[14].n39 0.0599512
R22669 XThC.Tn[14].n36 XThC.Tn[14].n35 0.0599512
R22670 XThC.Tn[14].n32 XThC.Tn[14].n31 0.0599512
R22671 XThC.Tn[14].n28 XThC.Tn[14].n27 0.0599512
R22672 XThC.Tn[14].n24 XThC.Tn[14].n23 0.0599512
R22673 XThC.Tn[14].n20 XThC.Tn[14].n19 0.0599512
R22674 XThC.Tn[14].n16 XThC.Tn[14].n15 0.0599512
R22675 XThC.Tn[14].n12 XThC.Tn[14].n11 0.0599512
R22676 XThC.Tn[14].n8 XThC.Tn[14].n7 0.0599512
R22677 XThC.Tn[14].n5 XThC.Tn[14].n4 0.0599512
R22678 XThC.Tn[14].n63 XThC.Tn[14] 0.0469286
R22679 XThC.Tn[14].n59 XThC.Tn[14] 0.0469286
R22680 XThC.Tn[14].n55 XThC.Tn[14] 0.0469286
R22681 XThC.Tn[14].n51 XThC.Tn[14] 0.0469286
R22682 XThC.Tn[14].n47 XThC.Tn[14] 0.0469286
R22683 XThC.Tn[14].n43 XThC.Tn[14] 0.0469286
R22684 XThC.Tn[14].n39 XThC.Tn[14] 0.0469286
R22685 XThC.Tn[14].n35 XThC.Tn[14] 0.0469286
R22686 XThC.Tn[14].n31 XThC.Tn[14] 0.0469286
R22687 XThC.Tn[14].n27 XThC.Tn[14] 0.0469286
R22688 XThC.Tn[14].n23 XThC.Tn[14] 0.0469286
R22689 XThC.Tn[14].n19 XThC.Tn[14] 0.0469286
R22690 XThC.Tn[14].n15 XThC.Tn[14] 0.0469286
R22691 XThC.Tn[14].n11 XThC.Tn[14] 0.0469286
R22692 XThC.Tn[14].n7 XThC.Tn[14] 0.0469286
R22693 XThC.Tn[14].n4 XThC.Tn[14] 0.0469286
R22694 XThC.Tn[14].n63 XThC.Tn[14] 0.0401341
R22695 XThC.Tn[14].n59 XThC.Tn[14] 0.0401341
R22696 XThC.Tn[14].n55 XThC.Tn[14] 0.0401341
R22697 XThC.Tn[14].n51 XThC.Tn[14] 0.0401341
R22698 XThC.Tn[14].n47 XThC.Tn[14] 0.0401341
R22699 XThC.Tn[14].n43 XThC.Tn[14] 0.0401341
R22700 XThC.Tn[14].n39 XThC.Tn[14] 0.0401341
R22701 XThC.Tn[14].n35 XThC.Tn[14] 0.0401341
R22702 XThC.Tn[14].n31 XThC.Tn[14] 0.0401341
R22703 XThC.Tn[14].n27 XThC.Tn[14] 0.0401341
R22704 XThC.Tn[14].n23 XThC.Tn[14] 0.0401341
R22705 XThC.Tn[14].n19 XThC.Tn[14] 0.0401341
R22706 XThC.Tn[14].n15 XThC.Tn[14] 0.0401341
R22707 XThC.Tn[14].n11 XThC.Tn[14] 0.0401341
R22708 XThC.Tn[14].n7 XThC.Tn[14] 0.0401341
R22709 XThC.Tn[14].n4 XThC.Tn[14] 0.0401341
R22710 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R22711 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R22712 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R22713 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R22714 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R22715 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R22716 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R22717 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R22718 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R22719 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22720 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22721 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22722 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22723 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22724 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22725 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22726 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22727 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22728 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22729 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22730 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22731 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22732 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22733 XThC.XTB1.Y.n0 XThC.XTB1.Y.t2 132.067
R22734 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22735 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22736 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22737 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22738 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22739 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22740 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22741 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22742 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22743 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22744 XThC.XTB1.Y.n2 XThC.XTB1.Y.t1 26.5955
R22745 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22746 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22747 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22748 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22749 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22750 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22751 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22752 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22753 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22754 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22755 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22756 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22757 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22758 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22759 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22760 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22761 XThC.Tn[8].n71 XThC.Tn[8].n70 256.104
R22762 XThC.Tn[8].n75 XThC.Tn[8].n74 243.679
R22763 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22764 XThC.Tn[8].n75 XThC.Tn[8].n73 205.28
R22765 XThC.Tn[8].n71 XThC.Tn[8].n69 202.095
R22766 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22767 XThC.Tn[8].n65 XThC.Tn[8].n63 161.365
R22768 XThC.Tn[8].n61 XThC.Tn[8].n59 161.365
R22769 XThC.Tn[8].n57 XThC.Tn[8].n55 161.365
R22770 XThC.Tn[8].n53 XThC.Tn[8].n51 161.365
R22771 XThC.Tn[8].n49 XThC.Tn[8].n47 161.365
R22772 XThC.Tn[8].n45 XThC.Tn[8].n43 161.365
R22773 XThC.Tn[8].n41 XThC.Tn[8].n39 161.365
R22774 XThC.Tn[8].n37 XThC.Tn[8].n35 161.365
R22775 XThC.Tn[8].n33 XThC.Tn[8].n31 161.365
R22776 XThC.Tn[8].n29 XThC.Tn[8].n27 161.365
R22777 XThC.Tn[8].n25 XThC.Tn[8].n23 161.365
R22778 XThC.Tn[8].n21 XThC.Tn[8].n19 161.365
R22779 XThC.Tn[8].n17 XThC.Tn[8].n15 161.365
R22780 XThC.Tn[8].n13 XThC.Tn[8].n11 161.365
R22781 XThC.Tn[8].n9 XThC.Tn[8].n7 161.365
R22782 XThC.Tn[8].n6 XThC.Tn[8].n4 161.365
R22783 XThC.Tn[8].n63 XThC.Tn[8].t15 161.202
R22784 XThC.Tn[8].n59 XThC.Tn[8].t37 161.202
R22785 XThC.Tn[8].n55 XThC.Tn[8].t24 161.202
R22786 XThC.Tn[8].n51 XThC.Tn[8].t21 161.202
R22787 XThC.Tn[8].n47 XThC.Tn[8].t13 161.202
R22788 XThC.Tn[8].n43 XThC.Tn[8].t32 161.202
R22789 XThC.Tn[8].n39 XThC.Tn[8].t31 161.202
R22790 XThC.Tn[8].n35 XThC.Tn[8].t12 161.202
R22791 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R22792 XThC.Tn[8].n27 XThC.Tn[8].t33 161.202
R22793 XThC.Tn[8].n23 XThC.Tn[8].t20 161.202
R22794 XThC.Tn[8].n19 XThC.Tn[8].t19 161.202
R22795 XThC.Tn[8].n15 XThC.Tn[8].t30 161.202
R22796 XThC.Tn[8].n11 XThC.Tn[8].t28 161.202
R22797 XThC.Tn[8].n7 XThC.Tn[8].t26 161.202
R22798 XThC.Tn[8].n4 XThC.Tn[8].t41 161.202
R22799 XThC.Tn[8].n63 XThC.Tn[8].t18 145.137
R22800 XThC.Tn[8].n59 XThC.Tn[8].t40 145.137
R22801 XThC.Tn[8].n55 XThC.Tn[8].t27 145.137
R22802 XThC.Tn[8].n51 XThC.Tn[8].t25 145.137
R22803 XThC.Tn[8].n47 XThC.Tn[8].t17 145.137
R22804 XThC.Tn[8].n43 XThC.Tn[8].t38 145.137
R22805 XThC.Tn[8].n39 XThC.Tn[8].t36 145.137
R22806 XThC.Tn[8].n35 XThC.Tn[8].t16 145.137
R22807 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R22808 XThC.Tn[8].n27 XThC.Tn[8].t39 145.137
R22809 XThC.Tn[8].n23 XThC.Tn[8].t23 145.137
R22810 XThC.Tn[8].n19 XThC.Tn[8].t22 145.137
R22811 XThC.Tn[8].n15 XThC.Tn[8].t35 145.137
R22812 XThC.Tn[8].n11 XThC.Tn[8].t34 145.137
R22813 XThC.Tn[8].n7 XThC.Tn[8].t29 145.137
R22814 XThC.Tn[8].n4 XThC.Tn[8].t43 145.137
R22815 XThC.Tn[8].n69 XThC.Tn[8].t9 26.5955
R22816 XThC.Tn[8].n69 XThC.Tn[8].t10 26.5955
R22817 XThC.Tn[8].n70 XThC.Tn[8].t8 26.5955
R22818 XThC.Tn[8].n70 XThC.Tn[8].t11 26.5955
R22819 XThC.Tn[8].n73 XThC.Tn[8].t2 26.5955
R22820 XThC.Tn[8].n73 XThC.Tn[8].t1 26.5955
R22821 XThC.Tn[8].n74 XThC.Tn[8].t0 26.5955
R22822 XThC.Tn[8].n74 XThC.Tn[8].t3 26.5955
R22823 XThC.Tn[8].n1 XThC.Tn[8].t7 24.9236
R22824 XThC.Tn[8].n1 XThC.Tn[8].t6 24.9236
R22825 XThC.Tn[8].n0 XThC.Tn[8].t5 24.9236
R22826 XThC.Tn[8].n0 XThC.Tn[8].t4 24.9236
R22827 XThC.Tn[8] XThC.Tn[8].n75 22.9652
R22828 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22829 XThC.Tn[8].n72 XThC.Tn[8].n71 13.9299
R22830 XThC.Tn[8] XThC.Tn[8].n72 13.9299
R22831 XThC.Tn[8] XThC.Tn[8].n6 8.0245
R22832 XThC.Tn[8].n66 XThC.Tn[8].n65 7.9105
R22833 XThC.Tn[8].n62 XThC.Tn[8].n61 7.9105
R22834 XThC.Tn[8].n58 XThC.Tn[8].n57 7.9105
R22835 XThC.Tn[8].n54 XThC.Tn[8].n53 7.9105
R22836 XThC.Tn[8].n50 XThC.Tn[8].n49 7.9105
R22837 XThC.Tn[8].n46 XThC.Tn[8].n45 7.9105
R22838 XThC.Tn[8].n42 XThC.Tn[8].n41 7.9105
R22839 XThC.Tn[8].n38 XThC.Tn[8].n37 7.9105
R22840 XThC.Tn[8].n34 XThC.Tn[8].n33 7.9105
R22841 XThC.Tn[8].n30 XThC.Tn[8].n29 7.9105
R22842 XThC.Tn[8].n26 XThC.Tn[8].n25 7.9105
R22843 XThC.Tn[8].n22 XThC.Tn[8].n21 7.9105
R22844 XThC.Tn[8].n18 XThC.Tn[8].n17 7.9105
R22845 XThC.Tn[8].n14 XThC.Tn[8].n13 7.9105
R22846 XThC.Tn[8].n10 XThC.Tn[8].n9 7.9105
R22847 XThC.Tn[8].n68 XThC.Tn[8].n67 7.42331
R22848 XThC.Tn[8].n67 XThC.Tn[8] 4.24005
R22849 XThC.Tn[8].n72 XThC.Tn[8].n68 2.99115
R22850 XThC.Tn[8].n72 XThC.Tn[8] 2.87153
R22851 XThC.Tn[8].n68 XThC.Tn[8] 2.2734
R22852 XThC.Tn[8].n3 XThC.Tn[8] 0.672375
R22853 XThC.Tn[8].n10 XThC.Tn[8] 0.235138
R22854 XThC.Tn[8].n14 XThC.Tn[8] 0.235138
R22855 XThC.Tn[8].n18 XThC.Tn[8] 0.235138
R22856 XThC.Tn[8].n22 XThC.Tn[8] 0.235138
R22857 XThC.Tn[8].n26 XThC.Tn[8] 0.235138
R22858 XThC.Tn[8].n30 XThC.Tn[8] 0.235138
R22859 XThC.Tn[8].n34 XThC.Tn[8] 0.235138
R22860 XThC.Tn[8].n38 XThC.Tn[8] 0.235138
R22861 XThC.Tn[8].n42 XThC.Tn[8] 0.235138
R22862 XThC.Tn[8].n46 XThC.Tn[8] 0.235138
R22863 XThC.Tn[8].n50 XThC.Tn[8] 0.235138
R22864 XThC.Tn[8].n54 XThC.Tn[8] 0.235138
R22865 XThC.Tn[8].n58 XThC.Tn[8] 0.235138
R22866 XThC.Tn[8].n62 XThC.Tn[8] 0.235138
R22867 XThC.Tn[8].n66 XThC.Tn[8] 0.235138
R22868 XThC.Tn[8].n67 XThC.Tn[8].n3 0.220435
R22869 XThC.Tn[8].n3 XThC.Tn[8] 0.168469
R22870 XThC.Tn[8] XThC.Tn[8].n10 0.114505
R22871 XThC.Tn[8] XThC.Tn[8].n14 0.114505
R22872 XThC.Tn[8] XThC.Tn[8].n18 0.114505
R22873 XThC.Tn[8] XThC.Tn[8].n22 0.114505
R22874 XThC.Tn[8] XThC.Tn[8].n26 0.114505
R22875 XThC.Tn[8] XThC.Tn[8].n30 0.114505
R22876 XThC.Tn[8] XThC.Tn[8].n34 0.114505
R22877 XThC.Tn[8] XThC.Tn[8].n38 0.114505
R22878 XThC.Tn[8] XThC.Tn[8].n42 0.114505
R22879 XThC.Tn[8] XThC.Tn[8].n46 0.114505
R22880 XThC.Tn[8] XThC.Tn[8].n50 0.114505
R22881 XThC.Tn[8] XThC.Tn[8].n54 0.114505
R22882 XThC.Tn[8] XThC.Tn[8].n58 0.114505
R22883 XThC.Tn[8] XThC.Tn[8].n62 0.114505
R22884 XThC.Tn[8] XThC.Tn[8].n66 0.114505
R22885 XThC.Tn[8].n65 XThC.Tn[8].n64 0.0599512
R22886 XThC.Tn[8].n61 XThC.Tn[8].n60 0.0599512
R22887 XThC.Tn[8].n57 XThC.Tn[8].n56 0.0599512
R22888 XThC.Tn[8].n53 XThC.Tn[8].n52 0.0599512
R22889 XThC.Tn[8].n49 XThC.Tn[8].n48 0.0599512
R22890 XThC.Tn[8].n45 XThC.Tn[8].n44 0.0599512
R22891 XThC.Tn[8].n41 XThC.Tn[8].n40 0.0599512
R22892 XThC.Tn[8].n37 XThC.Tn[8].n36 0.0599512
R22893 XThC.Tn[8].n33 XThC.Tn[8].n32 0.0599512
R22894 XThC.Tn[8].n29 XThC.Tn[8].n28 0.0599512
R22895 XThC.Tn[8].n25 XThC.Tn[8].n24 0.0599512
R22896 XThC.Tn[8].n21 XThC.Tn[8].n20 0.0599512
R22897 XThC.Tn[8].n17 XThC.Tn[8].n16 0.0599512
R22898 XThC.Tn[8].n13 XThC.Tn[8].n12 0.0599512
R22899 XThC.Tn[8].n9 XThC.Tn[8].n8 0.0599512
R22900 XThC.Tn[8].n6 XThC.Tn[8].n5 0.0599512
R22901 XThC.Tn[8].n64 XThC.Tn[8] 0.0469286
R22902 XThC.Tn[8].n60 XThC.Tn[8] 0.0469286
R22903 XThC.Tn[8].n56 XThC.Tn[8] 0.0469286
R22904 XThC.Tn[8].n52 XThC.Tn[8] 0.0469286
R22905 XThC.Tn[8].n48 XThC.Tn[8] 0.0469286
R22906 XThC.Tn[8].n44 XThC.Tn[8] 0.0469286
R22907 XThC.Tn[8].n40 XThC.Tn[8] 0.0469286
R22908 XThC.Tn[8].n36 XThC.Tn[8] 0.0469286
R22909 XThC.Tn[8].n32 XThC.Tn[8] 0.0469286
R22910 XThC.Tn[8].n28 XThC.Tn[8] 0.0469286
R22911 XThC.Tn[8].n24 XThC.Tn[8] 0.0469286
R22912 XThC.Tn[8].n20 XThC.Tn[8] 0.0469286
R22913 XThC.Tn[8].n16 XThC.Tn[8] 0.0469286
R22914 XThC.Tn[8].n12 XThC.Tn[8] 0.0469286
R22915 XThC.Tn[8].n8 XThC.Tn[8] 0.0469286
R22916 XThC.Tn[8].n5 XThC.Tn[8] 0.0469286
R22917 XThC.Tn[8].n64 XThC.Tn[8] 0.0401341
R22918 XThC.Tn[8].n60 XThC.Tn[8] 0.0401341
R22919 XThC.Tn[8].n56 XThC.Tn[8] 0.0401341
R22920 XThC.Tn[8].n52 XThC.Tn[8] 0.0401341
R22921 XThC.Tn[8].n48 XThC.Tn[8] 0.0401341
R22922 XThC.Tn[8].n44 XThC.Tn[8] 0.0401341
R22923 XThC.Tn[8].n40 XThC.Tn[8] 0.0401341
R22924 XThC.Tn[8].n36 XThC.Tn[8] 0.0401341
R22925 XThC.Tn[8].n32 XThC.Tn[8] 0.0401341
R22926 XThC.Tn[8].n28 XThC.Tn[8] 0.0401341
R22927 XThC.Tn[8].n24 XThC.Tn[8] 0.0401341
R22928 XThC.Tn[8].n20 XThC.Tn[8] 0.0401341
R22929 XThC.Tn[8].n16 XThC.Tn[8] 0.0401341
R22930 XThC.Tn[8].n12 XThC.Tn[8] 0.0401341
R22931 XThC.Tn[8].n8 XThC.Tn[8] 0.0401341
R22932 XThC.Tn[8].n5 XThC.Tn[8] 0.0401341
R22933 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R22934 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R22935 XThR.Tn[1] XThR.Tn[1].n82 161.363
R22936 XThR.Tn[1] XThR.Tn[1].n77 161.363
R22937 XThR.Tn[1] XThR.Tn[1].n72 161.363
R22938 XThR.Tn[1] XThR.Tn[1].n67 161.363
R22939 XThR.Tn[1] XThR.Tn[1].n62 161.363
R22940 XThR.Tn[1] XThR.Tn[1].n57 161.363
R22941 XThR.Tn[1] XThR.Tn[1].n52 161.363
R22942 XThR.Tn[1] XThR.Tn[1].n47 161.363
R22943 XThR.Tn[1] XThR.Tn[1].n42 161.363
R22944 XThR.Tn[1] XThR.Tn[1].n37 161.363
R22945 XThR.Tn[1] XThR.Tn[1].n32 161.363
R22946 XThR.Tn[1] XThR.Tn[1].n27 161.363
R22947 XThR.Tn[1] XThR.Tn[1].n22 161.363
R22948 XThR.Tn[1] XThR.Tn[1].n17 161.363
R22949 XThR.Tn[1] XThR.Tn[1].n12 161.363
R22950 XThR.Tn[1] XThR.Tn[1].n10 161.363
R22951 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R22952 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R22953 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R22954 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R22955 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R22956 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R22957 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R22958 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R22959 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R22960 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R22961 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R22962 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R22963 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R22964 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R22965 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R22966 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R22967 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R22968 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R22969 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R22970 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R22971 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R22972 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R22973 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R22974 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R22975 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R22976 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R22977 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R22978 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R22979 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R22980 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R22981 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R22982 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R22983 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R22984 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R22985 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R22986 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R22987 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R22988 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R22989 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R22990 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R22991 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R22992 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R22993 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R22994 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R22995 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R22996 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R22997 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R22998 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R22999 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R23000 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R23001 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R23002 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R23003 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R23004 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R23005 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R23006 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R23007 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R23008 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R23009 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R23010 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R23011 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R23012 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R23013 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R23014 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R23015 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R23016 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R23017 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R23018 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R23019 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R23020 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R23021 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R23022 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R23023 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R23024 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R23025 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R23026 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R23027 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R23028 XThR.Tn[1].n5 XThR.Tn[1].n3 135.249
R23029 XThR.Tn[1].n5 XThR.Tn[1].n4 98.981
R23030 XThR.Tn[1].n7 XThR.Tn[1].n6 98.981
R23031 XThR.Tn[1].n9 XThR.Tn[1].n8 98.981
R23032 XThR.Tn[1].n7 XThR.Tn[1].n5 36.2672
R23033 XThR.Tn[1].n9 XThR.Tn[1].n7 36.2672
R23034 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R23035 XThR.Tn[1].n1 XThR.Tn[1].t7 26.5955
R23036 XThR.Tn[1].n1 XThR.Tn[1].t6 26.5955
R23037 XThR.Tn[1].n0 XThR.Tn[1].t4 26.5955
R23038 XThR.Tn[1].n0 XThR.Tn[1].t5 26.5955
R23039 XThR.Tn[1].n3 XThR.Tn[1].t11 24.9236
R23040 XThR.Tn[1].n3 XThR.Tn[1].t8 24.9236
R23041 XThR.Tn[1].n4 XThR.Tn[1].t10 24.9236
R23042 XThR.Tn[1].n4 XThR.Tn[1].t9 24.9236
R23043 XThR.Tn[1].n6 XThR.Tn[1].t2 24.9236
R23044 XThR.Tn[1].n6 XThR.Tn[1].t1 24.9236
R23045 XThR.Tn[1].n8 XThR.Tn[1].t3 24.9236
R23046 XThR.Tn[1].n8 XThR.Tn[1].t0 24.9236
R23047 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R23048 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R23049 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R23050 XThR.Tn[1] XThR.Tn[1].n11 5.34038
R23051 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R23052 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R23053 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R23054 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R23055 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R23056 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R23057 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R23058 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R23059 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R23060 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R23061 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R23062 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R23063 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R23064 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R23065 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R23066 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R23067 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R23068 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R23069 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R23070 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R23071 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R23072 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R23073 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R23074 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R23075 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R23076 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R23077 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R23078 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R23079 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R23080 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R23081 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R23082 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R23083 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R23084 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R23085 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R23086 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R23087 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R23088 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R23089 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R23090 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R23091 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R23092 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R23093 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R23094 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R23095 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R23096 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R23097 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R23098 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R23099 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R23100 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R23101 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R23102 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R23103 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R23104 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R23105 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R23106 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R23107 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R23108 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R23109 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R23110 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R23111 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R23112 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R23113 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R23114 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R23115 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R23116 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R23117 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R23118 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R23119 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R23120 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R23121 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R23122 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R23123 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R23124 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R23125 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R23126 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R23127 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R23128 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R23129 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R23130 XThR.Tn[1] XThR.Tn[1].n87 0.038
R23131 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R23132 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R23133 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R23134 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R23135 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R23136 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R23137 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R23138 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R23139 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R23140 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R23141 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R23142 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R23143 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R23144 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R23145 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R23146 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R23147 XThC.Tn[7].n5 XThC.Tn[7].n4 255.096
R23148 XThC.Tn[7].n2 XThC.Tn[7].n0 236.589
R23149 XThC.Tn[7].n5 XThC.Tn[7].n3 201.845
R23150 XThC.Tn[7].n2 XThC.Tn[7].n1 200.321
R23151 XThC.Tn[7].n67 XThC.Tn[7].n65 161.365
R23152 XThC.Tn[7].n63 XThC.Tn[7].n61 161.365
R23153 XThC.Tn[7].n59 XThC.Tn[7].n57 161.365
R23154 XThC.Tn[7].n55 XThC.Tn[7].n53 161.365
R23155 XThC.Tn[7].n51 XThC.Tn[7].n49 161.365
R23156 XThC.Tn[7].n47 XThC.Tn[7].n45 161.365
R23157 XThC.Tn[7].n43 XThC.Tn[7].n41 161.365
R23158 XThC.Tn[7].n39 XThC.Tn[7].n37 161.365
R23159 XThC.Tn[7].n35 XThC.Tn[7].n33 161.365
R23160 XThC.Tn[7].n31 XThC.Tn[7].n29 161.365
R23161 XThC.Tn[7].n27 XThC.Tn[7].n25 161.365
R23162 XThC.Tn[7].n23 XThC.Tn[7].n21 161.365
R23163 XThC.Tn[7].n19 XThC.Tn[7].n17 161.365
R23164 XThC.Tn[7].n15 XThC.Tn[7].n13 161.365
R23165 XThC.Tn[7].n11 XThC.Tn[7].n9 161.365
R23166 XThC.Tn[7].n8 XThC.Tn[7].n6 161.365
R23167 XThC.Tn[7].n65 XThC.Tn[7].t19 161.202
R23168 XThC.Tn[7].n61 XThC.Tn[7].t9 161.202
R23169 XThC.Tn[7].n57 XThC.Tn[7].t28 161.202
R23170 XThC.Tn[7].n53 XThC.Tn[7].t26 161.202
R23171 XThC.Tn[7].n49 XThC.Tn[7].t17 161.202
R23172 XThC.Tn[7].n45 XThC.Tn[7].t38 161.202
R23173 XThC.Tn[7].n41 XThC.Tn[7].t36 161.202
R23174 XThC.Tn[7].n37 XThC.Tn[7].t16 161.202
R23175 XThC.Tn[7].n33 XThC.Tn[7].t14 161.202
R23176 XThC.Tn[7].n29 XThC.Tn[7].t39 161.202
R23177 XThC.Tn[7].n25 XThC.Tn[7].t23 161.202
R23178 XThC.Tn[7].n21 XThC.Tn[7].t22 161.202
R23179 XThC.Tn[7].n17 XThC.Tn[7].t35 161.202
R23180 XThC.Tn[7].n13 XThC.Tn[7].t34 161.202
R23181 XThC.Tn[7].n9 XThC.Tn[7].t30 161.202
R23182 XThC.Tn[7].n6 XThC.Tn[7].t11 161.202
R23183 XThC.Tn[7].n65 XThC.Tn[7].t15 145.137
R23184 XThC.Tn[7].n61 XThC.Tn[7].t37 145.137
R23185 XThC.Tn[7].n57 XThC.Tn[7].t24 145.137
R23186 XThC.Tn[7].n53 XThC.Tn[7].t21 145.137
R23187 XThC.Tn[7].n49 XThC.Tn[7].t13 145.137
R23188 XThC.Tn[7].n45 XThC.Tn[7].t32 145.137
R23189 XThC.Tn[7].n41 XThC.Tn[7].t31 145.137
R23190 XThC.Tn[7].n37 XThC.Tn[7].t12 145.137
R23191 XThC.Tn[7].n33 XThC.Tn[7].t10 145.137
R23192 XThC.Tn[7].n29 XThC.Tn[7].t33 145.137
R23193 XThC.Tn[7].n25 XThC.Tn[7].t20 145.137
R23194 XThC.Tn[7].n21 XThC.Tn[7].t18 145.137
R23195 XThC.Tn[7].n17 XThC.Tn[7].t29 145.137
R23196 XThC.Tn[7].n13 XThC.Tn[7].t27 145.137
R23197 XThC.Tn[7].n9 XThC.Tn[7].t25 145.137
R23198 XThC.Tn[7].n6 XThC.Tn[7].t8 145.137
R23199 XThC.Tn[7].n4 XThC.Tn[7].t2 26.5955
R23200 XThC.Tn[7].n4 XThC.Tn[7].t1 26.5955
R23201 XThC.Tn[7].n3 XThC.Tn[7].t0 26.5955
R23202 XThC.Tn[7].n3 XThC.Tn[7].t3 26.5955
R23203 XThC.Tn[7] XThC.Tn[7].n5 26.4992
R23204 XThC.Tn[7].n0 XThC.Tn[7].t6 24.9236
R23205 XThC.Tn[7].n0 XThC.Tn[7].t5 24.9236
R23206 XThC.Tn[7].n1 XThC.Tn[7].t4 24.9236
R23207 XThC.Tn[7].n1 XThC.Tn[7].t7 24.9236
R23208 XThC.Tn[7].n70 XThC.Tn[7].n2 12.0894
R23209 XThC.Tn[7].n70 XThC.Tn[7] 9.64206
R23210 XThC.Tn[7].n69 XThC.Tn[7] 8.14595
R23211 XThC.Tn[7] XThC.Tn[7].n8 8.0245
R23212 XThC.Tn[7].n68 XThC.Tn[7].n67 7.9105
R23213 XThC.Tn[7].n64 XThC.Tn[7].n63 7.9105
R23214 XThC.Tn[7].n60 XThC.Tn[7].n59 7.9105
R23215 XThC.Tn[7].n56 XThC.Tn[7].n55 7.9105
R23216 XThC.Tn[7].n52 XThC.Tn[7].n51 7.9105
R23217 XThC.Tn[7].n48 XThC.Tn[7].n47 7.9105
R23218 XThC.Tn[7].n44 XThC.Tn[7].n43 7.9105
R23219 XThC.Tn[7].n40 XThC.Tn[7].n39 7.9105
R23220 XThC.Tn[7].n36 XThC.Tn[7].n35 7.9105
R23221 XThC.Tn[7].n32 XThC.Tn[7].n31 7.9105
R23222 XThC.Tn[7].n28 XThC.Tn[7].n27 7.9105
R23223 XThC.Tn[7].n24 XThC.Tn[7].n23 7.9105
R23224 XThC.Tn[7].n20 XThC.Tn[7].n19 7.9105
R23225 XThC.Tn[7].n16 XThC.Tn[7].n15 7.9105
R23226 XThC.Tn[7].n12 XThC.Tn[7].n11 7.9105
R23227 XThC.Tn[7].n69 XThC.Tn[7] 5.30358
R23228 XThC.Tn[7] XThC.Tn[7].n69 3.15894
R23229 XThC.Tn[7] XThC.Tn[7].n70 1.66284
R23230 XThC.Tn[7].n12 XThC.Tn[7] 0.235138
R23231 XThC.Tn[7].n16 XThC.Tn[7] 0.235138
R23232 XThC.Tn[7].n20 XThC.Tn[7] 0.235138
R23233 XThC.Tn[7].n24 XThC.Tn[7] 0.235138
R23234 XThC.Tn[7].n28 XThC.Tn[7] 0.235138
R23235 XThC.Tn[7].n32 XThC.Tn[7] 0.235138
R23236 XThC.Tn[7].n36 XThC.Tn[7] 0.235138
R23237 XThC.Tn[7].n40 XThC.Tn[7] 0.235138
R23238 XThC.Tn[7].n44 XThC.Tn[7] 0.235138
R23239 XThC.Tn[7].n48 XThC.Tn[7] 0.235138
R23240 XThC.Tn[7].n52 XThC.Tn[7] 0.235138
R23241 XThC.Tn[7].n56 XThC.Tn[7] 0.235138
R23242 XThC.Tn[7].n60 XThC.Tn[7] 0.235138
R23243 XThC.Tn[7].n64 XThC.Tn[7] 0.235138
R23244 XThC.Tn[7].n68 XThC.Tn[7] 0.235138
R23245 XThC.Tn[7] XThC.Tn[7].n12 0.114505
R23246 XThC.Tn[7] XThC.Tn[7].n16 0.114505
R23247 XThC.Tn[7] XThC.Tn[7].n20 0.114505
R23248 XThC.Tn[7] XThC.Tn[7].n24 0.114505
R23249 XThC.Tn[7] XThC.Tn[7].n28 0.114505
R23250 XThC.Tn[7] XThC.Tn[7].n32 0.114505
R23251 XThC.Tn[7] XThC.Tn[7].n36 0.114505
R23252 XThC.Tn[7] XThC.Tn[7].n40 0.114505
R23253 XThC.Tn[7] XThC.Tn[7].n44 0.114505
R23254 XThC.Tn[7] XThC.Tn[7].n48 0.114505
R23255 XThC.Tn[7] XThC.Tn[7].n52 0.114505
R23256 XThC.Tn[7] XThC.Tn[7].n56 0.114505
R23257 XThC.Tn[7] XThC.Tn[7].n60 0.114505
R23258 XThC.Tn[7] XThC.Tn[7].n64 0.114505
R23259 XThC.Tn[7] XThC.Tn[7].n68 0.114505
R23260 XThC.Tn[7].n67 XThC.Tn[7].n66 0.0599512
R23261 XThC.Tn[7].n63 XThC.Tn[7].n62 0.0599512
R23262 XThC.Tn[7].n59 XThC.Tn[7].n58 0.0599512
R23263 XThC.Tn[7].n55 XThC.Tn[7].n54 0.0599512
R23264 XThC.Tn[7].n51 XThC.Tn[7].n50 0.0599512
R23265 XThC.Tn[7].n47 XThC.Tn[7].n46 0.0599512
R23266 XThC.Tn[7].n43 XThC.Tn[7].n42 0.0599512
R23267 XThC.Tn[7].n39 XThC.Tn[7].n38 0.0599512
R23268 XThC.Tn[7].n35 XThC.Tn[7].n34 0.0599512
R23269 XThC.Tn[7].n31 XThC.Tn[7].n30 0.0599512
R23270 XThC.Tn[7].n27 XThC.Tn[7].n26 0.0599512
R23271 XThC.Tn[7].n23 XThC.Tn[7].n22 0.0599512
R23272 XThC.Tn[7].n19 XThC.Tn[7].n18 0.0599512
R23273 XThC.Tn[7].n15 XThC.Tn[7].n14 0.0599512
R23274 XThC.Tn[7].n11 XThC.Tn[7].n10 0.0599512
R23275 XThC.Tn[7].n8 XThC.Tn[7].n7 0.0599512
R23276 XThC.Tn[7].n66 XThC.Tn[7] 0.0469286
R23277 XThC.Tn[7].n62 XThC.Tn[7] 0.0469286
R23278 XThC.Tn[7].n58 XThC.Tn[7] 0.0469286
R23279 XThC.Tn[7].n54 XThC.Tn[7] 0.0469286
R23280 XThC.Tn[7].n50 XThC.Tn[7] 0.0469286
R23281 XThC.Tn[7].n46 XThC.Tn[7] 0.0469286
R23282 XThC.Tn[7].n42 XThC.Tn[7] 0.0469286
R23283 XThC.Tn[7].n38 XThC.Tn[7] 0.0469286
R23284 XThC.Tn[7].n34 XThC.Tn[7] 0.0469286
R23285 XThC.Tn[7].n30 XThC.Tn[7] 0.0469286
R23286 XThC.Tn[7].n26 XThC.Tn[7] 0.0469286
R23287 XThC.Tn[7].n22 XThC.Tn[7] 0.0469286
R23288 XThC.Tn[7].n18 XThC.Tn[7] 0.0469286
R23289 XThC.Tn[7].n14 XThC.Tn[7] 0.0469286
R23290 XThC.Tn[7].n10 XThC.Tn[7] 0.0469286
R23291 XThC.Tn[7].n7 XThC.Tn[7] 0.0469286
R23292 XThC.Tn[7].n66 XThC.Tn[7] 0.0401341
R23293 XThC.Tn[7].n62 XThC.Tn[7] 0.0401341
R23294 XThC.Tn[7].n58 XThC.Tn[7] 0.0401341
R23295 XThC.Tn[7].n54 XThC.Tn[7] 0.0401341
R23296 XThC.Tn[7].n50 XThC.Tn[7] 0.0401341
R23297 XThC.Tn[7].n46 XThC.Tn[7] 0.0401341
R23298 XThC.Tn[7].n42 XThC.Tn[7] 0.0401341
R23299 XThC.Tn[7].n38 XThC.Tn[7] 0.0401341
R23300 XThC.Tn[7].n34 XThC.Tn[7] 0.0401341
R23301 XThC.Tn[7].n30 XThC.Tn[7] 0.0401341
R23302 XThC.Tn[7].n26 XThC.Tn[7] 0.0401341
R23303 XThC.Tn[7].n22 XThC.Tn[7] 0.0401341
R23304 XThC.Tn[7].n18 XThC.Tn[7] 0.0401341
R23305 XThC.Tn[7].n14 XThC.Tn[7] 0.0401341
R23306 XThC.Tn[7].n10 XThC.Tn[7] 0.0401341
R23307 XThC.Tn[7].n7 XThC.Tn[7] 0.0401341
R23308 XThR.Tn[4].n2 XThR.Tn[4].n1 332.332
R23309 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R23310 XThR.Tn[4] XThR.Tn[4].n82 161.363
R23311 XThR.Tn[4] XThR.Tn[4].n77 161.363
R23312 XThR.Tn[4] XThR.Tn[4].n72 161.363
R23313 XThR.Tn[4] XThR.Tn[4].n67 161.363
R23314 XThR.Tn[4] XThR.Tn[4].n62 161.363
R23315 XThR.Tn[4] XThR.Tn[4].n57 161.363
R23316 XThR.Tn[4] XThR.Tn[4].n52 161.363
R23317 XThR.Tn[4] XThR.Tn[4].n47 161.363
R23318 XThR.Tn[4] XThR.Tn[4].n42 161.363
R23319 XThR.Tn[4] XThR.Tn[4].n37 161.363
R23320 XThR.Tn[4] XThR.Tn[4].n32 161.363
R23321 XThR.Tn[4] XThR.Tn[4].n27 161.363
R23322 XThR.Tn[4] XThR.Tn[4].n22 161.363
R23323 XThR.Tn[4] XThR.Tn[4].n17 161.363
R23324 XThR.Tn[4] XThR.Tn[4].n12 161.363
R23325 XThR.Tn[4] XThR.Tn[4].n10 161.363
R23326 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R23327 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R23328 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R23329 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R23330 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R23331 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R23332 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R23333 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R23334 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R23335 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R23336 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R23337 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R23338 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R23339 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R23340 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R23341 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R23342 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R23343 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R23344 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R23345 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R23346 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R23347 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R23348 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R23349 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R23350 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R23351 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R23352 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R23353 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R23354 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R23355 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R23356 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R23357 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R23358 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R23359 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R23360 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R23361 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R23362 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R23363 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R23364 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R23365 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R23366 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R23367 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R23368 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R23369 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R23370 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R23371 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R23372 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R23373 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R23374 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R23375 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R23376 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R23377 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R23378 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R23379 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R23380 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R23381 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R23382 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R23383 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R23384 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R23385 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R23386 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R23387 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R23388 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R23389 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R23390 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R23391 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R23392 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R23393 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R23394 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R23395 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R23396 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R23397 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R23398 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R23399 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R23400 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R23401 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R23402 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R23403 XThR.Tn[4].n5 XThR.Tn[4].n3 135.249
R23404 XThR.Tn[4].n5 XThR.Tn[4].n4 98.982
R23405 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R23406 XThR.Tn[4].n9 XThR.Tn[4].n8 98.982
R23407 XThR.Tn[4].n7 XThR.Tn[4].n5 36.2672
R23408 XThR.Tn[4].n9 XThR.Tn[4].n7 36.2672
R23409 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R23410 XThR.Tn[4].n1 XThR.Tn[4].t4 26.5955
R23411 XThR.Tn[4].n1 XThR.Tn[4].t7 26.5955
R23412 XThR.Tn[4].n0 XThR.Tn[4].t5 26.5955
R23413 XThR.Tn[4].n0 XThR.Tn[4].t6 26.5955
R23414 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R23415 XThR.Tn[4].n3 XThR.Tn[4].t9 24.9236
R23416 XThR.Tn[4].n4 XThR.Tn[4].t11 24.9236
R23417 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R23418 XThR.Tn[4].n6 XThR.Tn[4].t2 24.9236
R23419 XThR.Tn[4].n6 XThR.Tn[4].t1 24.9236
R23420 XThR.Tn[4].n8 XThR.Tn[4].t3 24.9236
R23421 XThR.Tn[4].n8 XThR.Tn[4].t0 24.9236
R23422 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R23423 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R23424 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R23425 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R23426 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R23427 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R23428 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R23429 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R23430 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R23431 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R23432 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R23433 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R23434 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R23435 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R23436 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R23437 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R23438 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R23439 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R23440 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R23441 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R23442 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R23443 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R23444 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R23445 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R23446 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R23447 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R23448 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R23449 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R23450 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R23451 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R23452 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R23453 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R23454 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R23455 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R23456 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R23457 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R23458 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R23459 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R23460 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R23461 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R23462 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R23463 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R23464 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R23465 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R23466 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R23467 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R23468 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R23469 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R23470 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R23471 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R23472 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R23473 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R23474 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R23475 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R23476 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R23477 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R23478 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R23479 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R23480 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R23481 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R23482 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R23483 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R23484 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R23485 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R23486 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R23487 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R23488 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R23489 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R23490 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R23491 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R23492 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R23493 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R23494 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R23495 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R23496 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R23497 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R23498 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R23499 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R23500 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R23501 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R23502 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R23503 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R23504 XThR.Tn[4] XThR.Tn[4].n87 0.038
R23505 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R23506 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R23507 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R23508 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R23509 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R23510 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R23511 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R23512 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R23513 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R23514 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R23515 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R23516 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R23517 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R23518 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R23519 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R23520 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R23521 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R23522 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R23523 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R23524 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R23525 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R23526 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R23527 XThR.Tn[11] XThR.Tn[11].n82 161.363
R23528 XThR.Tn[11] XThR.Tn[11].n77 161.363
R23529 XThR.Tn[11] XThR.Tn[11].n72 161.363
R23530 XThR.Tn[11] XThR.Tn[11].n67 161.363
R23531 XThR.Tn[11] XThR.Tn[11].n62 161.363
R23532 XThR.Tn[11] XThR.Tn[11].n57 161.363
R23533 XThR.Tn[11] XThR.Tn[11].n52 161.363
R23534 XThR.Tn[11] XThR.Tn[11].n47 161.363
R23535 XThR.Tn[11] XThR.Tn[11].n42 161.363
R23536 XThR.Tn[11] XThR.Tn[11].n37 161.363
R23537 XThR.Tn[11] XThR.Tn[11].n32 161.363
R23538 XThR.Tn[11] XThR.Tn[11].n27 161.363
R23539 XThR.Tn[11] XThR.Tn[11].n22 161.363
R23540 XThR.Tn[11] XThR.Tn[11].n17 161.363
R23541 XThR.Tn[11] XThR.Tn[11].n12 161.363
R23542 XThR.Tn[11] XThR.Tn[11].n10 161.363
R23543 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R23544 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R23545 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R23546 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R23547 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R23548 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R23549 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R23550 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R23551 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R23552 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R23553 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R23554 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R23555 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R23556 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R23557 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R23558 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R23559 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R23560 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R23561 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R23562 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R23563 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R23564 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R23565 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R23566 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R23567 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R23568 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R23569 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R23570 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R23571 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R23572 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R23573 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R23574 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R23575 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R23576 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R23577 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R23578 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R23579 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R23580 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R23581 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R23582 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R23583 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R23584 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R23585 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R23586 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R23587 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R23588 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R23589 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R23590 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R23591 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R23592 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R23593 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R23594 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R23595 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R23596 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R23597 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R23598 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R23599 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R23600 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R23601 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R23602 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R23603 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R23604 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R23605 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R23606 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R23607 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R23608 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R23609 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R23610 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R23611 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R23612 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R23613 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R23614 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R23615 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R23616 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R23617 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R23618 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R23619 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R23620 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R23621 XThR.Tn[11].n6 XThR.Tn[11].t11 26.5955
R23622 XThR.Tn[11].n6 XThR.Tn[11].t3 26.5955
R23623 XThR.Tn[11].n7 XThR.Tn[11].t9 26.5955
R23624 XThR.Tn[11].n7 XThR.Tn[11].t2 26.5955
R23625 XThR.Tn[11].n3 XThR.Tn[11].t4 26.5955
R23626 XThR.Tn[11].n3 XThR.Tn[11].t6 26.5955
R23627 XThR.Tn[11].n4 XThR.Tn[11].t5 26.5955
R23628 XThR.Tn[11].n4 XThR.Tn[11].t7 26.5955
R23629 XThR.Tn[11].n0 XThR.Tn[11].t1 24.9236
R23630 XThR.Tn[11].n0 XThR.Tn[11].t10 24.9236
R23631 XThR.Tn[11].n1 XThR.Tn[11].t0 24.9236
R23632 XThR.Tn[11].n1 XThR.Tn[11].t8 24.9236
R23633 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R23634 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R23635 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R23636 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R23637 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R23638 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R23639 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R23640 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R23641 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R23642 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R23643 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R23644 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R23645 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R23646 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R23647 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R23648 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R23649 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R23650 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R23651 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R23652 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R23653 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R23654 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R23655 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R23656 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R23657 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R23658 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R23659 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R23660 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R23661 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R23662 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R23663 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R23664 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R23665 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R23666 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R23667 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R23668 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R23669 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R23670 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R23671 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R23672 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R23673 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R23674 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R23675 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R23676 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R23677 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R23678 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R23679 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R23680 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R23681 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R23682 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R23683 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R23684 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R23685 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R23686 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R23687 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R23688 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R23689 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R23690 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R23691 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R23692 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R23693 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R23694 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R23695 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R23696 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R23697 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R23698 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R23699 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R23700 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R23701 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R23702 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R23703 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R23704 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R23705 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R23706 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R23707 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R23708 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R23709 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R23710 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R23711 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R23712 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R23713 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R23714 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R23715 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R23716 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R23717 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R23718 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R23719 XThR.Tn[11] XThR.Tn[11].n87 0.038
R23720 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R23721 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R23722 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R23723 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R23724 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R23725 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R23726 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R23727 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R23728 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R23729 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R23730 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R23731 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R23732 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R23733 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R23734 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R23735 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R23736 XThR.Tn[7].n5 XThR.Tn[7].n3 244.067
R23737 XThR.Tn[7].n2 XThR.Tn[7].n0 236.589
R23738 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23739 XThR.Tn[7].n2 XThR.Tn[7].n1 200.321
R23740 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23741 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23742 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23743 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23744 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23745 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23746 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23747 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23748 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23749 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23750 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23751 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23752 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23753 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23754 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23755 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23756 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23757 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23758 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23759 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23760 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23761 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23762 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23763 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23764 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23765 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23766 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23767 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23768 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23769 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23770 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23771 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23772 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23773 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23774 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23775 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23776 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23777 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23778 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23779 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23780 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23781 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23782 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23783 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23784 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23785 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23786 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23787 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23788 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23789 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23790 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23791 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23792 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23793 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23794 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23795 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23796 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23797 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23798 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23799 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23800 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23801 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23802 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23803 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23804 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23805 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23806 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23807 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23808 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23809 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23810 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23811 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23812 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23813 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23814 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23815 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23816 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23817 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23818 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23819 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23820 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23821 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23822 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23823 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23824 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23825 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23826 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23827 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23828 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23829 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23830 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23831 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23832 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23833 XThR.Tn[7].n4 XThR.Tn[7].t1 26.5955
R23834 XThR.Tn[7].n4 XThR.Tn[7].t0 26.5955
R23835 XThR.Tn[7].n3 XThR.Tn[7].t2 26.5955
R23836 XThR.Tn[7].n3 XThR.Tn[7].t3 26.5955
R23837 XThR.Tn[7].n0 XThR.Tn[7].t7 24.9236
R23838 XThR.Tn[7].n0 XThR.Tn[7].t4 24.9236
R23839 XThR.Tn[7].n1 XThR.Tn[7].t6 24.9236
R23840 XThR.Tn[7].n1 XThR.Tn[7].t5 24.9236
R23841 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23842 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23843 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23844 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23845 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R23846 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23847 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23848 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23849 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23850 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23851 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23852 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23853 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23854 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23855 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23856 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23857 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23858 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23859 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23860 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23861 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23862 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23863 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23864 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23865 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23866 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23867 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23868 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23869 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23870 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23871 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23872 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23873 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23874 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23875 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23876 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23877 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23878 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23879 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23880 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23881 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23882 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23883 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23884 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23885 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23886 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23887 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23888 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23889 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23890 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23891 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23892 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23893 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23894 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23895 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23896 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23897 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23898 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23899 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23900 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23901 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23902 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23903 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23904 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23905 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23906 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23907 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23908 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23909 XThR.Tn[7].n6 XThR.Tn[7] 0.830612
R23910 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23911 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23912 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23913 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23914 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23915 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23916 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23917 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23918 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23919 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23920 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23921 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23922 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23923 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23924 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23925 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23926 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R23927 XThR.Tn[7] XThR.Tn[7].n84 0.038
R23928 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R23929 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R23930 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R23931 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R23932 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R23933 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R23934 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R23935 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R23936 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R23937 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R23938 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R23939 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R23940 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R23941 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R23942 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R23943 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R23944 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23945 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23946 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23947 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23948 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23949 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23950 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23951 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23952 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23953 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23954 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23955 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23956 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23957 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23958 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23959 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23960 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23961 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23962 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23963 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23964 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23965 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23966 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23967 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23968 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23969 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23970 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23971 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23972 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23973 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23974 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23975 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23976 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23977 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23978 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23979 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23980 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23981 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23982 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23983 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23984 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23985 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23986 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23987 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23988 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23989 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23990 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23991 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23992 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23993 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23994 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23995 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23996 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23997 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23998 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23999 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R24000 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R24001 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R24002 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R24003 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R24004 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R24005 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R24006 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R24007 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R24008 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R24009 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R24010 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R24011 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R24012 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R24013 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R24014 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R24015 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R24016 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R24017 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R24018 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R24019 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R24020 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R24021 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R24022 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R24023 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R24024 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R24025 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R24026 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R24027 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R24028 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R24029 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R24030 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R24031 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R24032 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R24033 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R24034 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R24035 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R24036 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R24037 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R24038 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R24039 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R24040 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R24041 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R24042 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R24043 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R24044 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R24045 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R24046 XThR.Tn[0].n1 XThR.Tn[0].t3 26.5955
R24047 XThR.Tn[0].n1 XThR.Tn[0].t2 26.5955
R24048 XThR.Tn[0].n0 XThR.Tn[0].t4 26.5955
R24049 XThR.Tn[0].n0 XThR.Tn[0].t5 26.5955
R24050 XThR.Tn[0].n3 XThR.Tn[0].t7 24.9236
R24051 XThR.Tn[0].n3 XThR.Tn[0].t8 24.9236
R24052 XThR.Tn[0].n4 XThR.Tn[0].t6 24.9236
R24053 XThR.Tn[0].n4 XThR.Tn[0].t9 24.9236
R24054 XThR.Tn[0].n5 XThR.Tn[0].t11 24.9236
R24055 XThR.Tn[0].n5 XThR.Tn[0].t10 24.9236
R24056 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R24057 XThR.Tn[0].n6 XThR.Tn[0].t1 24.9236
R24058 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R24059 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R24060 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R24061 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R24062 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R24063 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R24064 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R24065 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R24066 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R24067 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R24068 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R24069 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R24070 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R24071 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R24072 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R24073 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R24074 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R24075 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R24076 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R24077 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R24078 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R24079 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R24080 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R24081 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R24082 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R24083 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R24084 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R24085 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R24086 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R24087 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R24088 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R24089 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R24090 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R24091 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R24092 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R24093 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R24094 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R24095 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R24096 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R24097 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R24098 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R24099 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R24100 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R24101 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R24102 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R24103 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R24104 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R24105 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R24106 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R24107 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R24108 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R24109 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R24110 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R24111 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R24112 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R24113 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R24114 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R24115 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R24116 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R24117 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R24118 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R24119 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R24120 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R24121 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R24122 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R24123 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R24124 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R24125 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R24126 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R24127 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R24128 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R24129 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R24130 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R24131 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R24132 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R24133 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R24134 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R24135 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R24136 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R24137 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R24138 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R24139 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R24140 XThR.Tn[0] XThR.Tn[0].n87 0.038
R24141 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R24142 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R24143 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R24144 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R24145 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R24146 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R24147 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R24148 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R24149 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R24150 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R24151 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R24152 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R24153 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R24154 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R24155 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R24156 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R24157 XThR.Tn[8].n5 XThR.Tn[8].n4 256.103
R24158 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R24159 XThR.Tn[8].n88 XThR.Tn[8].n87 241.847
R24160 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R24161 XThR.Tn[8].n5 XThR.Tn[8].n3 202.095
R24162 XThR.Tn[8].n88 XThR.Tn[8].n86 185
R24163 XThR.Tn[8] XThR.Tn[8].n79 161.363
R24164 XThR.Tn[8] XThR.Tn[8].n74 161.363
R24165 XThR.Tn[8] XThR.Tn[8].n69 161.363
R24166 XThR.Tn[8] XThR.Tn[8].n64 161.363
R24167 XThR.Tn[8] XThR.Tn[8].n59 161.363
R24168 XThR.Tn[8] XThR.Tn[8].n54 161.363
R24169 XThR.Tn[8] XThR.Tn[8].n49 161.363
R24170 XThR.Tn[8] XThR.Tn[8].n44 161.363
R24171 XThR.Tn[8] XThR.Tn[8].n39 161.363
R24172 XThR.Tn[8] XThR.Tn[8].n34 161.363
R24173 XThR.Tn[8] XThR.Tn[8].n29 161.363
R24174 XThR.Tn[8] XThR.Tn[8].n24 161.363
R24175 XThR.Tn[8] XThR.Tn[8].n19 161.363
R24176 XThR.Tn[8] XThR.Tn[8].n14 161.363
R24177 XThR.Tn[8] XThR.Tn[8].n9 161.363
R24178 XThR.Tn[8] XThR.Tn[8].n7 161.363
R24179 XThR.Tn[8].n81 XThR.Tn[8].n80 161.3
R24180 XThR.Tn[8].n76 XThR.Tn[8].n75 161.3
R24181 XThR.Tn[8].n71 XThR.Tn[8].n70 161.3
R24182 XThR.Tn[8].n66 XThR.Tn[8].n65 161.3
R24183 XThR.Tn[8].n61 XThR.Tn[8].n60 161.3
R24184 XThR.Tn[8].n56 XThR.Tn[8].n55 161.3
R24185 XThR.Tn[8].n51 XThR.Tn[8].n50 161.3
R24186 XThR.Tn[8].n46 XThR.Tn[8].n45 161.3
R24187 XThR.Tn[8].n41 XThR.Tn[8].n40 161.3
R24188 XThR.Tn[8].n36 XThR.Tn[8].n35 161.3
R24189 XThR.Tn[8].n31 XThR.Tn[8].n30 161.3
R24190 XThR.Tn[8].n26 XThR.Tn[8].n25 161.3
R24191 XThR.Tn[8].n21 XThR.Tn[8].n20 161.3
R24192 XThR.Tn[8].n16 XThR.Tn[8].n15 161.3
R24193 XThR.Tn[8].n11 XThR.Tn[8].n10 161.3
R24194 XThR.Tn[8].n79 XThR.Tn[8].t23 161.106
R24195 XThR.Tn[8].n74 XThR.Tn[8].t29 161.106
R24196 XThR.Tn[8].n69 XThR.Tn[8].t71 161.106
R24197 XThR.Tn[8].n64 XThR.Tn[8].t57 161.106
R24198 XThR.Tn[8].n59 XThR.Tn[8].t21 161.106
R24199 XThR.Tn[8].n54 XThR.Tn[8].t46 161.106
R24200 XThR.Tn[8].n49 XThR.Tn[8].t27 161.106
R24201 XThR.Tn[8].n44 XThR.Tn[8].t69 161.106
R24202 XThR.Tn[8].n39 XThR.Tn[8].t56 161.106
R24203 XThR.Tn[8].n34 XThR.Tn[8].t61 161.106
R24204 XThR.Tn[8].n29 XThR.Tn[8].t44 161.106
R24205 XThR.Tn[8].n24 XThR.Tn[8].t70 161.106
R24206 XThR.Tn[8].n19 XThR.Tn[8].t43 161.106
R24207 XThR.Tn[8].n14 XThR.Tn[8].t26 161.106
R24208 XThR.Tn[8].n9 XThR.Tn[8].t49 161.106
R24209 XThR.Tn[8].n7 XThR.Tn[8].t33 161.106
R24210 XThR.Tn[8].n80 XThR.Tn[8].t19 159.978
R24211 XThR.Tn[8].n75 XThR.Tn[8].t25 159.978
R24212 XThR.Tn[8].n70 XThR.Tn[8].t67 159.978
R24213 XThR.Tn[8].n65 XThR.Tn[8].t54 159.978
R24214 XThR.Tn[8].n60 XThR.Tn[8].t16 159.978
R24215 XThR.Tn[8].n55 XThR.Tn[8].t42 159.978
R24216 XThR.Tn[8].n50 XThR.Tn[8].t24 159.978
R24217 XThR.Tn[8].n45 XThR.Tn[8].t64 159.978
R24218 XThR.Tn[8].n40 XThR.Tn[8].t51 159.978
R24219 XThR.Tn[8].n35 XThR.Tn[8].t58 159.978
R24220 XThR.Tn[8].n30 XThR.Tn[8].t41 159.978
R24221 XThR.Tn[8].n25 XThR.Tn[8].t66 159.978
R24222 XThR.Tn[8].n20 XThR.Tn[8].t40 159.978
R24223 XThR.Tn[8].n15 XThR.Tn[8].t22 159.978
R24224 XThR.Tn[8].n10 XThR.Tn[8].t45 159.978
R24225 XThR.Tn[8].n79 XThR.Tn[8].t73 145.038
R24226 XThR.Tn[8].n74 XThR.Tn[8].t35 145.038
R24227 XThR.Tn[8].n69 XThR.Tn[8].t15 145.038
R24228 XThR.Tn[8].n64 XThR.Tn[8].t62 145.038
R24229 XThR.Tn[8].n59 XThR.Tn[8].t30 145.038
R24230 XThR.Tn[8].n54 XThR.Tn[8].t72 145.038
R24231 XThR.Tn[8].n49 XThR.Tn[8].t17 145.038
R24232 XThR.Tn[8].n44 XThR.Tn[8].t63 145.038
R24233 XThR.Tn[8].n39 XThR.Tn[8].t60 145.038
R24234 XThR.Tn[8].n34 XThR.Tn[8].t28 145.038
R24235 XThR.Tn[8].n29 XThR.Tn[8].t52 145.038
R24236 XThR.Tn[8].n24 XThR.Tn[8].t12 145.038
R24237 XThR.Tn[8].n19 XThR.Tn[8].t50 145.038
R24238 XThR.Tn[8].n14 XThR.Tn[8].t34 145.038
R24239 XThR.Tn[8].n9 XThR.Tn[8].t59 145.038
R24240 XThR.Tn[8].n7 XThR.Tn[8].t39 145.038
R24241 XThR.Tn[8].n80 XThR.Tn[8].t32 143.911
R24242 XThR.Tn[8].n75 XThR.Tn[8].t55 143.911
R24243 XThR.Tn[8].n70 XThR.Tn[8].t37 143.911
R24244 XThR.Tn[8].n65 XThR.Tn[8].t18 143.911
R24245 XThR.Tn[8].n60 XThR.Tn[8].t48 143.911
R24246 XThR.Tn[8].n55 XThR.Tn[8].t31 143.911
R24247 XThR.Tn[8].n50 XThR.Tn[8].t38 143.911
R24248 XThR.Tn[8].n45 XThR.Tn[8].t20 143.911
R24249 XThR.Tn[8].n40 XThR.Tn[8].t14 143.911
R24250 XThR.Tn[8].n35 XThR.Tn[8].t47 143.911
R24251 XThR.Tn[8].n30 XThR.Tn[8].t68 143.911
R24252 XThR.Tn[8].n25 XThR.Tn[8].t36 143.911
R24253 XThR.Tn[8].n20 XThR.Tn[8].t65 143.911
R24254 XThR.Tn[8].n15 XThR.Tn[8].t53 143.911
R24255 XThR.Tn[8].n10 XThR.Tn[8].t13 143.911
R24256 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R24257 XThR.Tn[8].n3 XThR.Tn[8].t9 26.5955
R24258 XThR.Tn[8].n3 XThR.Tn[8].t7 26.5955
R24259 XThR.Tn[8].n4 XThR.Tn[8].t11 26.5955
R24260 XThR.Tn[8].n4 XThR.Tn[8].t2 26.5955
R24261 XThR.Tn[8].n0 XThR.Tn[8].t5 26.5955
R24262 XThR.Tn[8].n0 XThR.Tn[8].t3 26.5955
R24263 XThR.Tn[8].n1 XThR.Tn[8].t6 26.5955
R24264 XThR.Tn[8].n1 XThR.Tn[8].t4 26.5955
R24265 XThR.Tn[8].n86 XThR.Tn[8].t1 24.9236
R24266 XThR.Tn[8].n86 XThR.Tn[8].t10 24.9236
R24267 XThR.Tn[8].n87 XThR.Tn[8].t0 24.9236
R24268 XThR.Tn[8].n87 XThR.Tn[8].t8 24.9236
R24269 XThR.Tn[8] XThR.Tn[8].n88 18.8943
R24270 XThR.Tn[8].n6 XThR.Tn[8].n5 13.5534
R24271 XThR.Tn[8].n85 XThR.Tn[8] 7.82692
R24272 XThR.Tn[8] XThR.Tn[8].n85 6.34069
R24273 XThR.Tn[8] XThR.Tn[8].n8 5.34038
R24274 XThR.Tn[8].n13 XThR.Tn[8].n12 4.5005
R24275 XThR.Tn[8].n18 XThR.Tn[8].n17 4.5005
R24276 XThR.Tn[8].n23 XThR.Tn[8].n22 4.5005
R24277 XThR.Tn[8].n28 XThR.Tn[8].n27 4.5005
R24278 XThR.Tn[8].n33 XThR.Tn[8].n32 4.5005
R24279 XThR.Tn[8].n38 XThR.Tn[8].n37 4.5005
R24280 XThR.Tn[8].n43 XThR.Tn[8].n42 4.5005
R24281 XThR.Tn[8].n48 XThR.Tn[8].n47 4.5005
R24282 XThR.Tn[8].n53 XThR.Tn[8].n52 4.5005
R24283 XThR.Tn[8].n58 XThR.Tn[8].n57 4.5005
R24284 XThR.Tn[8].n63 XThR.Tn[8].n62 4.5005
R24285 XThR.Tn[8].n68 XThR.Tn[8].n67 4.5005
R24286 XThR.Tn[8].n73 XThR.Tn[8].n72 4.5005
R24287 XThR.Tn[8].n78 XThR.Tn[8].n77 4.5005
R24288 XThR.Tn[8].n83 XThR.Tn[8].n82 4.5005
R24289 XThR.Tn[8].n84 XThR.Tn[8] 3.70586
R24290 XThR.Tn[8].n13 XThR.Tn[8] 2.52282
R24291 XThR.Tn[8].n18 XThR.Tn[8] 2.52282
R24292 XThR.Tn[8].n23 XThR.Tn[8] 2.52282
R24293 XThR.Tn[8].n28 XThR.Tn[8] 2.52282
R24294 XThR.Tn[8].n33 XThR.Tn[8] 2.52282
R24295 XThR.Tn[8].n38 XThR.Tn[8] 2.52282
R24296 XThR.Tn[8].n43 XThR.Tn[8] 2.52282
R24297 XThR.Tn[8].n48 XThR.Tn[8] 2.52282
R24298 XThR.Tn[8].n53 XThR.Tn[8] 2.52282
R24299 XThR.Tn[8].n58 XThR.Tn[8] 2.52282
R24300 XThR.Tn[8].n63 XThR.Tn[8] 2.52282
R24301 XThR.Tn[8].n68 XThR.Tn[8] 2.52282
R24302 XThR.Tn[8].n73 XThR.Tn[8] 2.52282
R24303 XThR.Tn[8].n78 XThR.Tn[8] 2.52282
R24304 XThR.Tn[8].n83 XThR.Tn[8] 2.52282
R24305 XThR.Tn[8].n85 XThR.Tn[8] 1.79489
R24306 XThR.Tn[8].n6 XThR.Tn[8] 1.50638
R24307 XThR.Tn[8] XThR.Tn[8].n6 1.19676
R24308 XThR.Tn[8].n81 XThR.Tn[8] 1.08677
R24309 XThR.Tn[8].n76 XThR.Tn[8] 1.08677
R24310 XThR.Tn[8].n71 XThR.Tn[8] 1.08677
R24311 XThR.Tn[8].n66 XThR.Tn[8] 1.08677
R24312 XThR.Tn[8].n61 XThR.Tn[8] 1.08677
R24313 XThR.Tn[8].n56 XThR.Tn[8] 1.08677
R24314 XThR.Tn[8].n51 XThR.Tn[8] 1.08677
R24315 XThR.Tn[8].n46 XThR.Tn[8] 1.08677
R24316 XThR.Tn[8].n41 XThR.Tn[8] 1.08677
R24317 XThR.Tn[8].n36 XThR.Tn[8] 1.08677
R24318 XThR.Tn[8].n31 XThR.Tn[8] 1.08677
R24319 XThR.Tn[8].n26 XThR.Tn[8] 1.08677
R24320 XThR.Tn[8].n21 XThR.Tn[8] 1.08677
R24321 XThR.Tn[8].n16 XThR.Tn[8] 1.08677
R24322 XThR.Tn[8].n11 XThR.Tn[8] 1.08677
R24323 XThR.Tn[8] XThR.Tn[8].n13 0.839786
R24324 XThR.Tn[8] XThR.Tn[8].n18 0.839786
R24325 XThR.Tn[8] XThR.Tn[8].n23 0.839786
R24326 XThR.Tn[8] XThR.Tn[8].n28 0.839786
R24327 XThR.Tn[8] XThR.Tn[8].n33 0.839786
R24328 XThR.Tn[8] XThR.Tn[8].n38 0.839786
R24329 XThR.Tn[8] XThR.Tn[8].n43 0.839786
R24330 XThR.Tn[8] XThR.Tn[8].n48 0.839786
R24331 XThR.Tn[8] XThR.Tn[8].n53 0.839786
R24332 XThR.Tn[8] XThR.Tn[8].n58 0.839786
R24333 XThR.Tn[8] XThR.Tn[8].n63 0.839786
R24334 XThR.Tn[8] XThR.Tn[8].n68 0.839786
R24335 XThR.Tn[8] XThR.Tn[8].n73 0.839786
R24336 XThR.Tn[8] XThR.Tn[8].n78 0.839786
R24337 XThR.Tn[8] XThR.Tn[8].n83 0.839786
R24338 XThR.Tn[8].n8 XThR.Tn[8] 0.499542
R24339 XThR.Tn[8].n82 XThR.Tn[8] 0.063
R24340 XThR.Tn[8].n77 XThR.Tn[8] 0.063
R24341 XThR.Tn[8].n72 XThR.Tn[8] 0.063
R24342 XThR.Tn[8].n67 XThR.Tn[8] 0.063
R24343 XThR.Tn[8].n62 XThR.Tn[8] 0.063
R24344 XThR.Tn[8].n57 XThR.Tn[8] 0.063
R24345 XThR.Tn[8].n52 XThR.Tn[8] 0.063
R24346 XThR.Tn[8].n47 XThR.Tn[8] 0.063
R24347 XThR.Tn[8].n42 XThR.Tn[8] 0.063
R24348 XThR.Tn[8].n37 XThR.Tn[8] 0.063
R24349 XThR.Tn[8].n32 XThR.Tn[8] 0.063
R24350 XThR.Tn[8].n27 XThR.Tn[8] 0.063
R24351 XThR.Tn[8].n22 XThR.Tn[8] 0.063
R24352 XThR.Tn[8].n17 XThR.Tn[8] 0.063
R24353 XThR.Tn[8].n12 XThR.Tn[8] 0.063
R24354 XThR.Tn[8].n84 XThR.Tn[8] 0.0540714
R24355 XThR.Tn[8] XThR.Tn[8].n84 0.038
R24356 XThR.Tn[8].n8 XThR.Tn[8] 0.0143889
R24357 XThR.Tn[8].n82 XThR.Tn[8].n81 0.00771154
R24358 XThR.Tn[8].n77 XThR.Tn[8].n76 0.00771154
R24359 XThR.Tn[8].n72 XThR.Tn[8].n71 0.00771154
R24360 XThR.Tn[8].n67 XThR.Tn[8].n66 0.00771154
R24361 XThR.Tn[8].n62 XThR.Tn[8].n61 0.00771154
R24362 XThR.Tn[8].n57 XThR.Tn[8].n56 0.00771154
R24363 XThR.Tn[8].n52 XThR.Tn[8].n51 0.00771154
R24364 XThR.Tn[8].n47 XThR.Tn[8].n46 0.00771154
R24365 XThR.Tn[8].n42 XThR.Tn[8].n41 0.00771154
R24366 XThR.Tn[8].n37 XThR.Tn[8].n36 0.00771154
R24367 XThR.Tn[8].n32 XThR.Tn[8].n31 0.00771154
R24368 XThR.Tn[8].n27 XThR.Tn[8].n26 0.00771154
R24369 XThR.Tn[8].n22 XThR.Tn[8].n21 0.00771154
R24370 XThR.Tn[8].n17 XThR.Tn[8].n16 0.00771154
R24371 XThR.Tn[8].n12 XThR.Tn[8].n11 0.00771154
R24372 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R24373 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R24374 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R24375 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R24376 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R24377 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R24378 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R24379 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R24380 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R24381 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R24382 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R24383 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R24384 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R24385 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R24386 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R24387 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R24388 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R24389 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R24390 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R24391 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R24392 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R24393 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R24394 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R24395 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R24396 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R24397 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R24398 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R24399 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R24400 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R24401 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R24402 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R24403 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R24404 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R24405 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R24406 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R24407 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R24408 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R24409 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R24410 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R24411 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R24412 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R24413 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R24414 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R24415 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R24416 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R24417 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R24418 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R24419 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R24420 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R24421 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R24422 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R24423 data[4].n3 data[4].t0 231.835
R24424 data[4].n0 data[4].t3 230.155
R24425 data[4].n0 data[4].t1 157.856
R24426 data[4].n3 data[4].t2 157.07
R24427 data[4].n1 data[4].n0 152
R24428 data[4].n4 data[4].n3 152
R24429 data[4].n2 data[4].n1 25.6681
R24430 data[4].n4 data[4].n2 10.7642
R24431 data[4].n2 data[4] 2.763
R24432 data[4].n1 data[4] 2.10199
R24433 data[4] data[4].n4 2.01193
R24434 XThR.Tn[13].n87 XThR.Tn[13].n86 256.104
R24435 XThR.Tn[13].n2 XThR.Tn[13].n1 243.68
R24436 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R24437 XThR.Tn[13].n2 XThR.Tn[13].n0 205.28
R24438 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R24439 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R24440 XThR.Tn[13] XThR.Tn[13].n78 161.363
R24441 XThR.Tn[13] XThR.Tn[13].n73 161.363
R24442 XThR.Tn[13] XThR.Tn[13].n68 161.363
R24443 XThR.Tn[13] XThR.Tn[13].n63 161.363
R24444 XThR.Tn[13] XThR.Tn[13].n58 161.363
R24445 XThR.Tn[13] XThR.Tn[13].n53 161.363
R24446 XThR.Tn[13] XThR.Tn[13].n48 161.363
R24447 XThR.Tn[13] XThR.Tn[13].n43 161.363
R24448 XThR.Tn[13] XThR.Tn[13].n38 161.363
R24449 XThR.Tn[13] XThR.Tn[13].n33 161.363
R24450 XThR.Tn[13] XThR.Tn[13].n28 161.363
R24451 XThR.Tn[13] XThR.Tn[13].n23 161.363
R24452 XThR.Tn[13] XThR.Tn[13].n18 161.363
R24453 XThR.Tn[13] XThR.Tn[13].n13 161.363
R24454 XThR.Tn[13] XThR.Tn[13].n8 161.363
R24455 XThR.Tn[13] XThR.Tn[13].n6 161.363
R24456 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R24457 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R24458 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R24459 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R24460 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R24461 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R24462 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R24463 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R24464 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R24465 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R24466 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R24467 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R24468 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R24469 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R24470 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R24471 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R24472 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R24473 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R24474 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R24475 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R24476 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R24477 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R24478 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R24479 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R24480 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R24481 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R24482 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R24483 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R24484 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R24485 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R24486 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R24487 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R24488 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R24489 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R24490 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R24491 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R24492 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R24493 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R24494 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R24495 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R24496 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R24497 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R24498 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R24499 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R24500 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R24501 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R24502 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R24503 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R24504 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R24505 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R24506 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R24507 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R24508 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R24509 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R24510 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R24511 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R24512 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R24513 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R24514 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R24515 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R24516 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R24517 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R24518 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R24519 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R24520 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R24521 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R24522 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R24523 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R24524 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R24525 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R24526 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R24527 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R24528 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R24529 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R24530 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R24531 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R24532 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R24533 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R24534 XThR.Tn[13].n85 XThR.Tn[13].t10 26.5955
R24535 XThR.Tn[13].n85 XThR.Tn[13].t8 26.5955
R24536 XThR.Tn[13].n86 XThR.Tn[13].t11 26.5955
R24537 XThR.Tn[13].n86 XThR.Tn[13].t9 26.5955
R24538 XThR.Tn[13].n0 XThR.Tn[13].t2 26.5955
R24539 XThR.Tn[13].n0 XThR.Tn[13].t0 26.5955
R24540 XThR.Tn[13].n1 XThR.Tn[13].t1 26.5955
R24541 XThR.Tn[13].n1 XThR.Tn[13].t3 26.5955
R24542 XThR.Tn[13].n4 XThR.Tn[13].t6 24.9236
R24543 XThR.Tn[13].n4 XThR.Tn[13].t4 24.9236
R24544 XThR.Tn[13].n3 XThR.Tn[13].t7 24.9236
R24545 XThR.Tn[13].n3 XThR.Tn[13].t5 24.9236
R24546 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R24547 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R24548 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R24549 XThR.Tn[13] XThR.Tn[13].n7 5.34038
R24550 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R24551 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R24552 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R24553 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R24554 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R24555 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R24556 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R24557 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R24558 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R24559 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R24560 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R24561 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R24562 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R24563 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R24564 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R24565 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R24566 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R24567 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R24568 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R24569 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R24570 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R24571 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R24572 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R24573 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R24574 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R24575 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R24576 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R24577 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R24578 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R24579 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R24580 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R24581 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R24582 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R24583 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R24584 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R24585 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R24586 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R24587 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R24588 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R24589 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R24590 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R24591 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R24592 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R24593 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R24594 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R24595 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R24596 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R24597 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R24598 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R24599 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R24600 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R24601 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R24602 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R24603 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R24604 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R24605 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R24606 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R24607 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R24608 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R24609 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R24610 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R24611 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R24612 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R24613 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R24614 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R24615 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R24616 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R24617 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R24618 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R24619 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R24620 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R24621 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R24622 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R24623 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R24624 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R24625 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R24626 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R24627 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R24628 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R24629 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R24630 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R24631 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R24632 XThR.Tn[13] XThR.Tn[13].n83 0.038
R24633 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R24634 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R24635 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R24636 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R24637 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R24638 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R24639 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R24640 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R24641 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R24642 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R24643 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R24644 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R24645 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R24646 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R24647 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R24648 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R24649 data[0].n1 data[0].t0 230.155
R24650 data[0].n0 data[0].t2 228.463
R24651 data[0].n1 data[0].t1 157.856
R24652 data[0].n0 data[0].t3 157.07
R24653 data[0].n2 data[0].n1 152.768
R24654 data[0].n4 data[0].n0 152.256
R24655 data[0].n3 data[0].n2 24.1398
R24656 data[0].n4 data[0].n3 9.48418
R24657 data[0] data[0].n4 6.1445
R24658 data[0].n2 data[0] 5.6325
R24659 data[0].n3 data[0] 2.638
R24660 XThR.XTB4.Y XThR.XTB4.Y.t0 230.518
R24661 XThR.XTB4.Y.n10 XThR.XTB4.Y.t12 212.081
R24662 XThR.XTB4.Y.n11 XThR.XTB4.Y.t2 212.081
R24663 XThR.XTB4.Y.n16 XThR.XTB4.Y.t7 212.081
R24664 XThR.XTB4.Y.n17 XThR.XTB4.Y.t6 212.081
R24665 XThR.XTB4.Y.n0 XThR.XTB4.Y.t17 212.081
R24666 XThR.XTB4.Y.n1 XThR.XTB4.Y.t5 212.081
R24667 XThR.XTB4.Y.n3 XThR.XTB4.Y.t15 212.081
R24668 XThR.XTB4.Y.n4 XThR.XTB4.Y.t4 212.081
R24669 XThR.XTB4.Y.n13 XThR.XTB4.Y.n12 173.761
R24670 XThR.XTB4.Y.n2 XThR.XTB4.Y 167.361
R24671 XThR.XTB4.Y.n19 XThR.XTB4.Y.n18 152
R24672 XThR.XTB4.Y.n15 XThR.XTB4.Y.n14 152
R24673 XThR.XTB4.Y.n13 XThR.XTB4.Y.n9 152
R24674 XThR.XTB4.Y.n6 XThR.XTB4.Y.n5 152
R24675 XThR.XTB4.Y.n10 XThR.XTB4.Y.t3 139.78
R24676 XThR.XTB4.Y.n11 XThR.XTB4.Y.t9 139.78
R24677 XThR.XTB4.Y.n16 XThR.XTB4.Y.t14 139.78
R24678 XThR.XTB4.Y.n17 XThR.XTB4.Y.t11 139.78
R24679 XThR.XTB4.Y.n0 XThR.XTB4.Y.t10 139.78
R24680 XThR.XTB4.Y.n1 XThR.XTB4.Y.t16 139.78
R24681 XThR.XTB4.Y.n3 XThR.XTB4.Y.t8 139.78
R24682 XThR.XTB4.Y.n4 XThR.XTB4.Y.t13 139.78
R24683 XThR.XTB4.Y.n21 XThR.XTB4.Y.t1 133.386
R24684 XThR.XTB4.Y.n20 XThR.XTB4.Y.n19 72.9296
R24685 XThR.XTB4.Y.n1 XThR.XTB4.Y.n0 61.346
R24686 XThR.XTB4.Y.n15 XThR.XTB4.Y.n9 49.6611
R24687 XThR.XTB4.Y.n18 XThR.XTB4.Y.n16 45.2793
R24688 XThR.XTB4.Y.n12 XThR.XTB4.Y.n11 42.3581
R24689 XThR.XTB4.Y.n20 XThR.XTB4.Y.n8 38.1854
R24690 XThR.XTB4.Y.n2 XThR.XTB4.Y.n1 30.6732
R24691 XThR.XTB4.Y.n3 XThR.XTB4.Y.n2 30.6732
R24692 XThR.XTB4.Y.n5 XThR.XTB4.Y.n3 30.6732
R24693 XThR.XTB4.Y.n5 XThR.XTB4.Y.n4 30.6732
R24694 XThR.XTB4.Y XThR.XTB4.Y.n21 28.966
R24695 XThR.XTB4.Y.n14 XThR.XTB4.Y.n13 21.7605
R24696 XThR.XTB4.Y.n14 XThR.XTB4.Y 21.1205
R24697 XThR.XTB4.Y.n12 XThR.XTB4.Y.n10 18.9884
R24698 XThR.XTB4.Y.n18 XThR.XTB4.Y.n17 16.0672
R24699 XThR.XTB4.Y.n21 XThR.XTB4.Y.n20 11.994
R24700 XThR.XTB4.Y.n22 XThR.XTB4.Y 11.6875
R24701 XThR.XTB4.Y.n8 XThR.XTB4.Y.n7 8.21182
R24702 XThR.XTB4.Y.n11 XThR.XTB4.Y.n9 7.30353
R24703 XThR.XTB4.Y.n8 XThR.XTB4.Y.n6 7.24578
R24704 XThR.XTB4.Y.n22 XThR.XTB4.Y 7.23528
R24705 XThR.XTB4.Y.n6 XThR.XTB4.Y 6.08654
R24706 XThR.XTB4.Y XThR.XTB4.Y.n22 5.04292
R24707 XThR.XTB4.Y.n16 XThR.XTB4.Y.n15 4.38232
R24708 XThR.XTB4.Y.n7 XThR.XTB4.Y 1.79489
R24709 XThR.XTB4.Y.n7 XThR.XTB4.Y 0.966538
R24710 XThR.XTB4.Y.n19 XThR.XTB4.Y 0.6405
R24711 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R24712 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R24713 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R24714 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R24715 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R24716 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R24717 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R24718 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R24719 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24720 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24721 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24722 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24723 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24724 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24725 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24726 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24727 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24728 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24729 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24730 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24731 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24732 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24733 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24734 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24735 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24736 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24737 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24738 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24739 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24740 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24741 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24742 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24743 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24744 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24745 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24746 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24747 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24748 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24749 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24750 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24751 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24752 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24753 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24754 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24755 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24756 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24757 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24758 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24759 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24760 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24761 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24762 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24763 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R24764 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R24765 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R24766 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R24767 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R24768 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R24769 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R24770 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R24771 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R24772 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R24773 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R24774 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R24775 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R24776 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R24777 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R24778 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R24779 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R24780 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R24781 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R24782 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R24783 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R24784 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R24785 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R24786 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R24787 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R24788 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R24789 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R24790 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R24791 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R24792 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R24793 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R24794 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R24795 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R24796 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R24797 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R24798 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R24799 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R24800 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R24801 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R24802 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R24803 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R24804 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R24805 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R24806 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R24807 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R24808 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R24809 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R24810 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R24811 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R24812 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R24813 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R24814 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R24815 data[6].n0 data[6].t0 230.576
R24816 data[6].n0 data[6].t1 158.275
R24817 data[6].n1 data[6].n0 152
R24818 data[6].n1 data[6] 11.9995
R24819 data[6] data[6].n1 6.66717
R24820 data[1].n4 data[1].t2 230.576
R24821 data[1].n1 data[1].t0 230.363
R24822 data[1].n0 data[1].t4 229.369
R24823 data[1].n4 data[1].t5 158.275
R24824 data[1].n1 data[1].t3 158.064
R24825 data[1].n0 data[1].t1 157.07
R24826 data[1].n2 data[1].n1 153.28
R24827 data[1].n7 data[1].n0 153.147
R24828 data[1].n5 data[1].n4 152
R24829 data[1].n7 data[1].n6 16.3874
R24830 data[1].n6 data[1].n5 14.9641
R24831 data[1].n3 data[1].n2 9.3005
R24832 data[1].n6 data[1].n3 6.49639
R24833 data[1] data[1].n7 3.24826
R24834 data[1].n2 data[1] 2.92621
R24835 data[1].n3 data[1] 2.15819
R24836 data[1].n5 data[1] 2.13383
R24837 data[2].n0 data[2].t0 230.576
R24838 data[2].n0 data[2].t1 158.275
R24839 data[2].n1 data[2].n0 152
R24840 data[2].n1 data[2] 12.7714
R24841 data[2] data[2].n1 2.13383
R24842 data[5].n4 data[5].t2 230.576
R24843 data[5].n1 data[5].t0 230.363
R24844 data[5].n0 data[5].t1 229.369
R24845 data[5].n4 data[5].t5 158.275
R24846 data[5].n1 data[5].t3 158.064
R24847 data[5].n0 data[5].t4 157.07
R24848 data[5].n2 data[5].n1 152.256
R24849 data[5].n7 data[5].n0 152.238
R24850 data[5].n5 data[5].n4 152
R24851 data[5].n7 data[5].n6 16.3874
R24852 data[5].n6 data[5].n5 14.6005
R24853 data[5].n3 data[5].n2 9.3005
R24854 data[5].n5 data[5] 6.66717
R24855 data[5].n6 data[5].n3 6.49639
R24856 data[5].n2 data[5] 6.1445
R24857 data[5] data[5].n7 5.68939
R24858 data[5].n3 data[5] 2.28319
R24859 bias[0] bias[0].t0 12.1467
R24860 bias[2].n0 bias[2].t0 56.8043
R24861 bias[2].n0 bias[2] 6.35112
R24862 bias[2] bias[2].n0 0.828709
R24863 data[3].n0 data[3].t1 230.576
R24864 data[3].n0 data[3].t0 158.275
R24865 data[3].n1 data[3].n0 153.553
R24866 data[3].n1 data[3] 11.6078
R24867 data[3] data[3].n1 2.90959
R24868 data[7].n0 data[7].t0 230.576
R24869 data[7].n0 data[7].t1 158.275
R24870 data[7].n1 data[7].n0 152
R24871 data[7].n1 data[7] 11.9995
R24872 data[7] data[7].n1 6.66717
R24873 bias[1] bias[1].t0 23.8076
C0 XA.XIR[9].XIC[6].icell.SM Iout 0.00388f
C1 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00214f
C2 XThR.XTBN.A a_n997_1803# 0.09118f
C3 XThR.XTB3.Y data[4] 0.03253f
C4 XThC.Tn[9] XThR.Tn[4] 0.28739f
C5 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.SM 0.00168f
C6 XThC.XTBN.Y XThC.Tn[12] 0.56523f
C7 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C8 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C9 XA.XIR[0].XIC[3].icell.SM VPWR 0.00158f
C10 XThC.XTB6.A a_6243_10571# 0.00295f
C11 XA.XIR[8].XIC_dummy_left.icell.Ien Vbias 0.00329f
C12 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04031f
C13 XThR.Tn[10] XA.XIR[11].XIC[12].icell.Ien 0.00338f
C14 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02762f
C15 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04031f
C16 XA.XIR[8].XIC[14].icell.SM Vbias 0.00701f
C17 XA.XIR[3].XIC[13].icell.Ien VPWR 0.1903f
C18 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00584f
C19 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10] 0.00341f
C20 XA.XIR[15].XIC[13].icell.PDM Iout 0.00117f
C21 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00256f
C22 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PUM 0.00465f
C23 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00584f
C24 XA.XIR[3].XIC[9].icell.Ien Iout 0.06417f
C25 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C26 XA.XIR[1].XIC[11].icell.PDM Iout 0.00117f
C27 XThC.Tn[0] XA.XIR[8].XIC_dummy_left.icell.Iout 0.00109f
C28 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[7].icell.Ien 0.00214f
C29 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PUM 0.00465f
C30 XThC.Tn[13] XThR.Tn[10] 0.2874f
C31 XThC.Tn[3] XThR.Tn[0] 0.28743f
C32 XA.XIR[7].XIC[6].icell.SM VPWR 0.00158f
C33 XA.XIR[2].XIC[6].icell.Ien VPWR 0.1903f
C34 XThC.Tn[5] XThR.Tn[5] 0.28739f
C35 a_n997_715# VPWR 0.02818f
C36 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C37 XA.XIR[2].XIC[2].icell.Ien Iout 0.06417f
C38 XA.XIR[1].XIC[8].icell.Ien VPWR 0.1903f
C39 XA.XIR[4].XIC[11].icell.PDM Iout 0.00117f
C40 XA.XIR[7].XIC[2].icell.SM Iout 0.00388f
C41 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.15202f
C42 XThC.Tn[6] XA.XIR[0].XIC[7].icell.Ien 0.002f
C43 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C44 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00214f
C45 XThR.Tn[13] XA.XIR[14].XIC[12].icell.SM 0.00121f
C46 XThC.Tn[10] XThC.Tn[12] 0.00453f
C47 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.SM 0.0039f
C48 a_3773_9615# Vbias 0.00846f
C49 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.0404f
C50 XA.XIR[13].XIC[14].icell.SM Iout 0.00388f
C51 XA.XIR[1].XIC[4].icell.Ien Iout 0.06417f
C52 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13] 0.00341f
C53 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00214f
C54 XThR.Tn[7] XA.XIR[8].XIC[3].icell.SM 0.00121f
C55 XA.XIR[12].XIC_dummy_right.icell.SM VPWR 0.00123f
C56 XThR.Tn[6] XA.XIR[7].XIC[14].icell.SM 0.00121f
C57 XA.XIR[5].XIC[4].icell.PDM Vbias 0.04261f
C58 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00584f
C59 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02762f
C60 XA.XIR[8].XIC[12].icell.Ien Iout 0.06417f
C61 XThC.XTB7.B data[2] 0.07481f
C62 XThR.Tn[8] XA.XIR[9].XIC[12].icell.Ien 0.00338f
C63 XThR.XTBN.A XThR.Tn[13] 0.00106f
C64 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C65 XA.XIR[15].XIC[0].icell.PUM VPWR 0.00937f
C66 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.SM 0.00168f
C67 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.15202f
C68 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00214f
C69 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PUM 0.00465f
C70 XThR.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.00341f
C71 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02762f
C72 XA.XIR[12].XIC[3].icell.PDM Vbias 0.04261f
C73 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Ien 0.00584f
C74 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C75 XThR.Tn[10] XA.XIR[11].XIC[4].icell.SM 0.00121f
C76 XThR.Tn[3] XA.XIR[3].XIC[5].icell.PDM 0.00341f
C77 a_5949_9615# VPWR 0.7053f
C78 XThR.Tn[1] XA.XIR[2].XIC[5].icell.Ien 0.00338f
C79 XA.XIR[11].XIC[9].icell.PDM Vbias 0.04261f
C80 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.03425f
C81 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.03425f
C82 XA.XIR[6].XIC[1].icell.PDM VPWR 0.00799f
C83 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C84 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04031f
C85 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PUM 0.00186f
C86 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.03554f
C87 XThR.XTB3.Y a_n997_2667# 0.002f
C88 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C89 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.15202f
C90 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.15202f
C91 XA.XIR[0].XIC[14].icell.Ien Iout 0.06389f
C92 XA.XIR[5].XIC[8].icell.PDM VPWR 0.00799f
C93 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C94 XThC.Tn[2] XThR.Tn[2] 0.28739f
C95 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C96 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.SM 0.0039f
C97 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.SM 0.0039f
C98 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.SM 0.0039f
C99 XA.XIR[3].XIC[3].icell.PUM Vbias 0.0031f
C100 XThR.Tn[13] XA.XIR[14].XIC[9].icell.Ien 0.00338f
C101 XThR.XTB6.A a_n1335_4229# 0.00304f
C102 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C103 XA.XIR[13].XIC[2].icell.PDM VPWR 0.00799f
C104 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00214f
C105 XThC.Tn[11] XThR.Tn[14] 0.28739f
C106 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.03425f
C107 XA.XIR[13].XIC[11].icell.Ien Iout 0.06417f
C108 XThC.XTB5.A VPWR 0.82807f
C109 XThR.Tn[3] VPWR 6.64542f
C110 XA.XIR[6].XIC[6].icell.SM Vbias 0.00701f
C111 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00584f
C112 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C113 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C114 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PUM 0.00465f
C115 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PUM 0.00465f
C116 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C117 XA.XIR[15].XIC[9].icell.PUM Vbias 0.0031f
C118 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00189f
C119 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C120 XA.XIR[12].XIC[7].icell.PDM VPWR 0.00799f
C121 XA.XIR[5].XIC[9].icell.Ien Vbias 0.21098f
C122 XThR.Tn[0] XA.XIR[1].XIC[12].icell.Ien 0.00338f
C123 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C124 XA.XIR[15].XIC[0].icell.SM Iout 0.00388f
C125 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.SM 0.0039f
C126 XThR.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.00338f
C127 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C128 XA.XIR[4].XIC[12].icell.PUM Vbias 0.0031f
C129 XA.XIR[8].XIC[1].icell.PDM Vbias 0.04261f
C130 XThR.XTB7.Y VPWR 1.14768f
C131 VPWR data[4] 0.5303f
C132 XA.XIR[11].XIC[1].icell.PDM Iout 0.00117f
C133 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.SM 0.00168f
C134 XA.XIR[2].XIC[5].icell.PDM Vbias 0.04261f
C135 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Iout 0.00347f
C136 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.03425f
C137 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11107f
C138 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C139 XA.XIR[13].XIC[2].icell.SM Vbias 0.00701f
C140 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.SM 0.00168f
C141 XThR.Tn[5] XA.XIR[6].XIC[14].icell.Ien 0.00338f
C142 XA.XIR[10].XIC[5].icell.PDM Iout 0.00117f
C143 XA.XIR[8].XIC[6].icell.PUM Vbias 0.0031f
C144 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C145 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.SM 0.0039f
C146 XA.XIR[15].XIC_15.icell.Ien VPWR 0.36724f
C147 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04031f
C148 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C149 XA.XIR[3].XIC[3].icell.SM VPWR 0.00158f
C150 XA.XIR[10].XIC[12].icell.SM VPWR 0.00158f
C151 XThR.XTB6.Y a_n997_1803# 0.00871f
C152 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.SM 0.0039f
C153 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.SM 0.00168f
C154 XA.XIR[12].XIC[4].icell.Ien Vbias 0.21098f
C155 XA.XIR[6].XIC[8].icell.Ien VPWR 0.1903f
C156 XThR.Tn[13] XA.XIR[14].XIC[10].icell.SM 0.00121f
C157 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.03425f
C158 XA.XIR[11].XIC[5].icell.SM Vbias 0.00701f
C159 XThC.XTBN.A XThC.Tn[9] 0.12399f
C160 XA.XIR[6].XIC[4].icell.Ien Iout 0.06417f
C161 XA.XIR[5].XIC[11].icell.PUM VPWR 0.00937f
C162 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.SM 0.0039f
C163 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7] 0.00341f
C164 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.03425f
C165 XThC.Tn[7] XThR.Tn[6] 0.28739f
C166 XThC.XTBN.Y a_10915_9569# 0.21503f
C167 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.SM 0.0039f
C168 XThR.Tn[10] XA.XIR[11].XIC[0].icell.Ien 0.00338f
C169 XA.XIR[15].XIC[5].icell.SM Iout 0.00388f
C170 XA.XIR[9].XIC_15.icell.PUM Vbias 0.0031f
C171 XThC.Tn[0] XThR.Tn[11] 0.28744f
C172 XA.XIR[10].XIC[7].icell.SM Vbias 0.00701f
C173 XA.XIR[4].XIC[12].icell.SM VPWR 0.00158f
C174 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00584f
C175 XThR.XTBN.Y XA.XIR[13].XIC_dummy_left.icell.Iout 0.00446f
C176 XA.XIR[3].XIC[3].icell.PDM VPWR 0.00799f
C177 XA.XIR[12].XIC[11].icell.PDM Iout 0.00117f
C178 XA.XIR[8].XIC[5].icell.PDM VPWR 0.00799f
C179 XA.XIR[14].XIC[2].icell.Ien VPWR 0.19084f
C180 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C181 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00584f
C182 XA.XIR[4].XIC[8].icell.SM Iout 0.00388f
C183 XA.XIR[0].XIC[8].icell.PUM Vbias 0.0031f
C184 XA.XIR[2].XIC[9].icell.PDM VPWR 0.00799f
C185 XThC.XTB7.A XThC.XTB7.B 0.35844f
C186 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C187 XA.XIR[13].XIC[4].icell.Ien VPWR 0.1903f
C188 XA.XIR[8].XIC[6].icell.SM VPWR 0.00158f
C189 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.SM 0.00168f
C190 XA.XIR[15].XIC[12].icell.PDM Iout 0.00117f
C191 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00584f
C192 XA.XIR[12].XIC[6].icell.PUM VPWR 0.00937f
C193 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12] 0.00341f
C194 XA.XIR[8].XIC[2].icell.SM Iout 0.00388f
C195 XThR.Tn[8] XA.XIR[9].XIC[2].icell.SM 0.00121f
C196 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02762f
C197 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.03425f
C198 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C199 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01577f
C200 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C201 XA.XIR[5].XIC_dummy_left.icell.Ien Vbias 0.00329f
C202 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.SM 0.0039f
C203 XA.XIR[2].XIC[9].icell.SM Vbias 0.00701f
C204 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04031f
C205 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C206 XA.XIR[11].XIC[7].icell.Ien VPWR 0.1903f
C207 XA.XIR[7].XIC[11].icell.PUM Vbias 0.0031f
C208 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C209 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PUM 0.00465f
C210 XA.XIR[5].XIC_15.icell.SM VPWR 0.00275f
C211 XThR.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.00338f
C212 XThC.XTB6.Y XThC.Tn[5] 0.20189f
C213 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C214 XA.XIR[11].XIC[3].icell.Ien Iout 0.06417f
C215 XA.XIR[1].XIC[11].icell.SM Vbias 0.00704f
C216 XA.XIR[10].XIC[9].icell.Ien VPWR 0.1903f
C217 XThC.Tn[13] XThR.Tn[13] 0.2874f
C218 XThR.Tn[3] XA.XIR[4].XIC[4].icell.Ien 0.00338f
C219 XA.XIR[9].XIC[11].icell.SM Iout 0.00388f
C220 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13] 0.00341f
C221 XA.XIR[10].XIC[5].icell.Ien Iout 0.06417f
C222 XThC.Tn[3] XThR.Tn[1] 0.28739f
C223 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.SM 0.00168f
C224 XThR.Tn[9] XA.XIR[10].XIC[5].icell.Ien 0.00338f
C225 XA.XIR[0].XIC[8].icell.SM VPWR 0.00158f
C226 a_n997_2667# VPWR 0.01642f
C227 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.03425f
C228 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.SM 0.0039f
C229 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C230 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C231 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C232 XA.XIR[0].XIC[4].icell.SM Iout 0.00367f
C233 XA.XIR[8].XIC[1].icell.PUM Vbias 0.0031f
C234 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04031f
C235 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.SM 0.00168f
C236 XThC.Tn[3] XThR.Tn[12] 0.28739f
C237 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.03425f
C238 XA.XIR[3].XIC[14].icell.Ien Iout 0.06417f
C239 XThC.Tn[12] XThR.Tn[8] 0.28739f
C240 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04031f
C241 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38708f
C242 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8] 0.00341f
C243 XA.XIR[2].XIC[11].icell.Ien VPWR 0.1903f
C244 XThR.Tn[7] Vbias 3.74624f
C245 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.SM 0.0039f
C246 XA.XIR[7].XIC[11].icell.SM VPWR 0.00158f
C247 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PUM 0.00465f
C248 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.03425f
C249 XA.XIR[7].XIC_15.icell.SM Vbias 0.00701f
C250 XThC.XTBN.Y XThC.Tn[1] 0.7252f
C251 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.SM 0.0039f
C252 XA.XIR[2].XIC[7].icell.Ien Iout 0.06417f
C253 XA.XIR[7].XIC[7].icell.SM Iout 0.00388f
C254 XA.XIR[7].XIC[5].icell.PDM Vbias 0.04261f
C255 XA.XIR[10].XIC_15.icell.SM Iout 0.0047f
C256 XThR.Tn[0] XA.XIR[1].XIC[2].icell.SM 0.00121f
C257 XA.XIR[1].XIC[13].icell.Ien VPWR 0.1903f
C258 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04031f
C259 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.15202f
C260 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.SM 0.00168f
C261 XThR.Tn[12] XA.XIR[13].XIC[3].icell.Ien 0.00338f
C262 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PUM 0.00465f
C263 XThC.Tn[7] XThR.Tn[4] 0.28739f
C264 XA.XIR[1].XIC[9].icell.Ien Iout 0.06417f
C265 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C266 a_n1049_7493# XA.XIR[1].XIC_dummy_left.icell.Iout 0.0013f
C267 XA.XIR[15].XIC[3].icell.PDM Vbias 0.04261f
C268 XA.XIR[4].XIC[2].icell.Ien Vbias 0.21098f
C269 XA.XIR[6].XIC[12].icell.PDM Vbias 0.04261f
C270 XA.XIR[10].XIC[10].icell.SM VPWR 0.00158f
C271 XThR.Tn[13] XA.XIR[14].XIC[14].icell.Ien 0.00338f
C272 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.04432f
C273 XThR.Tn[7] XA.XIR[8].XIC[8].icell.SM 0.00121f
C274 VPWR bias[1] 1.33312f
C275 XA.XIR[3].XIC[0].icell.SM VPWR 0.00158f
C276 XThC.XTB7.B a_5949_9615# 0.00927f
C277 XA.XIR[14].XIC[9].icell.PDM Vbias 0.04261f
C278 XThC.XTB4.Y XThC.Tn[5] 0.00814f
C279 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C280 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.SM 0.0039f
C281 XThC.Tn[2] XThR.Tn[10] 0.28739f
C282 XThR.Tn[5] XA.XIR[6].XIC[4].icell.SM 0.00121f
C283 XA.XIR[12].XIC[0].icell.Ien VPWR 0.1903f
C284 XThR.Tn[11] XA.XIR[12].XIC[6].icell.Ien 0.00338f
C285 XThC.XTB3.Y XThC.Tn[9] 0.00285f
C286 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.SM 0.00168f
C287 XThC.XTB6.Y a_10051_9569# 0.07626f
C288 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PDM 0.00172f
C289 XThR.Tn[10] XA.XIR[11].XIC_15.icell.Ien 0.00117f
C290 XThR.Tn[11] VPWR 7.58404f
C291 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.15202f
C292 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.SM 0.0039f
C293 XA.XIR[9].XIC[1].icell.PDM Vbias 0.04261f
C294 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04031f
C295 XA.XIR[7].XIC[9].icell.PDM VPWR 0.00799f
C296 XA.XIR[9].XIC[2].icell.PUM VPWR 0.00937f
C297 XThC.XTB5.A XThC.XTB7.B 0.30355f
C298 XA.XIR[12].XIC[12].icell.SM Vbias 0.00701f
C299 XThR.XTB6.A a_n1319_5611# 0.00467f
C300 XA.XIR[9].XIC[5].icell.Ien Vbias 0.21098f
C301 XThR.Tn[1] XA.XIR[2].XIC[10].icell.Ien 0.00338f
C302 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C303 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.SM 0.0039f
C304 XA.XIR[15].XIC[7].icell.PDM VPWR 0.0114f
C305 XA.XIR[4].XIC[4].icell.PUM VPWR 0.00937f
C306 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.SM 0.0039f
C307 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00214f
C308 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.15202f
C309 XA.XIR[6].XIC[4].icell.PDM Iout 0.00117f
C310 XA.XIR[10].XIC[13].icell.PUM VPWR 0.00937f
C311 XA.XIR[3].XIC[8].icell.PUM Vbias 0.0031f
C312 XA.XIR[5].XIC[11].icell.PDM Iout 0.00117f
C313 XA.XIR[14].XIC[1].icell.PDM Iout 0.00117f
C314 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00584f
C315 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C316 XA.XIR[1].XIC[6].icell.PDM Vbias 0.04261f
C317 XA.XIR[6].XIC[11].icell.SM Vbias 0.00701f
C318 a_8739_9569# VPWR 0.00583f
C319 XA.XIR[9].XIC[5].icell.PDM VPWR 0.00799f
C320 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00584f
C321 XThR.XTB7.A a_n1331_2891# 0.00995f
C322 XA.XIR[13].XIC[5].icell.PDM Iout 0.00117f
C323 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C324 XA.XIR[13].XIC[12].icell.SM VPWR 0.00158f
C325 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00584f
C326 XA.XIR[4].XIC[6].icell.PDM Vbias 0.04261f
C327 XA.XIR[5].XIC[14].icell.Ien Vbias 0.21098f
C328 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.SM 0.00168f
C329 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.SM 0.00168f
C330 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.03425f
C331 XA.XIR[12].XIC[10].icell.PDM Iout 0.00117f
C332 XA.XIR[9].XIC[7].icell.PUM VPWR 0.00937f
C333 XA.XIR[1].XIC[3].icell.PUM Vbias 0.0031f
C334 XA.XIR[3].XIC[14].icell.PDM Vbias 0.04261f
C335 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.SM 0.00168f
C336 XA.XIR[14].XIC[5].icell.SM Vbias 0.00701f
C337 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.SM 0.0039f
C338 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.SM 0.0039f
C339 XThR.XTBN.A a_n997_3979# 0.02087f
C340 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00584f
C341 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C342 XA.XIR[12].XIC_15.icell.PUM Vbias 0.0031f
C343 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.03425f
C344 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C345 XA.XIR[13].XIC[7].icell.SM Vbias 0.00701f
C346 XThC.Tn[0] XThR.Tn[14] 0.28742f
C347 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C348 XA.XIR[15].XIC[11].icell.PDM Iout 0.00117f
C349 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04031f
C350 XA.XIR[8].XIC[11].icell.PUM Vbias 0.0031f
C351 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02762f
C352 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.SM 0.0039f
C353 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C354 XThR.Tn[11] XA.XIR[12].XIC[0].icell.SM 0.00127f
C355 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.03425f
C356 XA.XIR[3].XIC[8].icell.SM VPWR 0.00158f
C357 XA.XIR[1].XIC[10].icell.PDM VPWR 0.00799f
C358 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.SM 0.00168f
C359 XA.XIR[12].XIC[9].icell.Ien Vbias 0.21098f
C360 XA.XIR[6].XIC[13].icell.Ien VPWR 0.1903f
C361 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PUM 0.00429f
C362 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00214f
C363 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14] 0.00341f
C364 XA.XIR[15].XIC_dummy_right.icell.SM VPWR 0.00123f
C365 XA.XIR[10].XIC[14].icell.Ien VPWR 0.19036f
C366 XA.XIR[3].XIC[4].icell.SM Iout 0.00388f
C367 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.SM 0.00168f
C368 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.SM 0.00168f
C369 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[4].icell.SM 0.0039f
C370 XA.XIR[4].XIC[10].icell.PDM VPWR 0.00799f
C371 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C372 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02762f
C373 XA.XIR[2].XIC[1].icell.SM VPWR 0.00158f
C374 XA.XIR[6].XIC[9].icell.Ien Iout 0.06417f
C375 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7] 0.00341f
C376 XA.XIR[7].XIC[3].icell.PUM VPWR 0.00937f
C377 XThR.XTB6.A XThR.Tn[5] 0.00361f
C378 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04031f
C379 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02762f
C380 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.SM 0.00168f
C381 XThR.Tn[13] XA.XIR[14].XIC[12].icell.Ien 0.00338f
C382 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02762f
C383 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00214f
C384 XA.XIR[1].XIC[3].icell.SM VPWR 0.00158f
C385 XA.XIR[9].XIC[0].icell.Ien Vbias 0.20951f
C386 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01577f
C387 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13] 0.00341f
C388 XA.XIR[14].XIC[7].icell.Ien VPWR 0.19084f
C389 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.SM 0.00168f
C390 XA.XIR[4].XIC[13].icell.SM Iout 0.00388f
C391 XA.XIR[3].XIC[6].icell.PDM Iout 0.00117f
C392 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C393 XA.XIR[14].XIC[3].icell.Ien Iout 0.06417f
C394 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.SM 0.00168f
C395 XA.XIR[0].XIC[13].icell.PUM Vbias 0.0031f
C396 XA.XIR[8].XIC[8].icell.PDM Iout 0.00117f
C397 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04031f
C398 XA.XIR[13].XIC[9].icell.Ien VPWR 0.1903f
C399 XA.XIR[8].XIC[11].icell.SM VPWR 0.00158f
C400 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.03023f
C401 XThC.Tn[11] VPWR 6.86576f
C402 XA.XIR[2].XIC[12].icell.PDM Iout 0.00117f
C403 XA.XIR[8].XIC_15.icell.SM Vbias 0.00701f
C404 XA.XIR[13].XIC[5].icell.Ien Iout 0.06417f
C405 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C406 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00584f
C407 XA.XIR[8].XIC[7].icell.SM Iout 0.00388f
C408 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.Ien 0.00584f
C409 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C410 XThR.Tn[8] XA.XIR[9].XIC[7].icell.SM 0.00121f
C411 XThR.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.00338f
C412 XThC.XTBN.A XThC.Tn[7] 0.01439f
C413 XThR.Tn[0] XA.XIR[0].XIC[9].icell.PDM 0.00341f
C414 XA.XIR[7].XIC_dummy_right.icell.PUM Vbias 0.00223f
C415 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.0404f
C416 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.15202f
C417 XA.XIR[2].XIC[14].icell.SM Vbias 0.00701f
C418 XA.XIR[12].XIC[10].icell.SM Vbias 0.00701f
C419 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.SM 0.0039f
C420 XThR.Tn[4] XA.XIR[5].XIC[9].icell.Ien 0.00338f
C421 XThR.Tn[1] XA.XIR[1].XIC[7].icell.PDM 0.00341f
C422 XA.XIR[5].XIC[1].icell.PUM Vbias 0.0031f
C423 XA.XIR[11].XIC[8].icell.Ien Iout 0.06417f
C424 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00214f
C425 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PUM 0.00465f
C426 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04031f
C427 XThR.XTBN.A XThR.Tn[7] 0.01439f
C428 XThR.Tn[3] XA.XIR[4].XIC[9].icell.Ien 0.00338f
C429 XThC.Tn[0] XA.XIR[2].XIC_dummy_left.icell.Iout 0.00109f
C430 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00584f
C431 XThR.XTBN.A a_n997_2891# 0.01719f
C432 XA.XIR[10].XIC[11].icell.PUM VPWR 0.00937f
C433 XA.XIR[0].XIC[13].icell.SM VPWR 0.00158f
C434 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5] 0.00341f
C435 XA.XIR[13].XIC_15.icell.SM Iout 0.0047f
C436 XThR.Tn[6] XThR.Tn[7] 0.06617f
C437 XA.XIR[10].XIC[0].icell.PDM Vbias 0.04207f
C438 XA.XIR[0].XIC[9].icell.SM Iout 0.00367f
C439 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00584f
C440 XA.XIR[12].XIC_dummy_left.icell.SM VPWR 0.00269f
C441 XThR.Tn[2] XA.XIR[2].XIC[4].icell.PDM 0.00341f
C442 XA.XIR[13].XIC[10].icell.SM VPWR 0.00158f
C443 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.03425f
C444 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04052f
C445 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PUM 0.00465f
C446 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04031f
C447 XThR.Tn[13] XA.XIR[14].XIC[4].icell.SM 0.00121f
C448 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[12].icell.Ien 0.00214f
C449 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C450 data[6] data[7] 0.04128f
C451 XA.XIR[6].XIC[3].icell.PUM Vbias 0.0031f
C452 XThC.Tn[2] XThR.Tn[13] 0.28739f
C453 XA.XIR[15].XIC[1].icell.PUM VPWR 0.00937f
C454 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6] 0.00341f
C455 XA.XIR[5].XIC[1].icell.Ien VPWR 0.1903f
C456 XA.XIR[2].XIC[12].icell.Ien Iout 0.06417f
C457 XA.XIR[15].XIC[4].icell.Ien Vbias 0.17899f
C458 XA.XIR[7].XIC[12].icell.SM Iout 0.00388f
C459 XThR.Tn[0] XA.XIR[1].XIC[7].icell.SM 0.00121f
C460 XA.XIR[5].XIC[4].icell.SM Vbias 0.00701f
C461 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.15202f
C462 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.SM 0.00168f
C463 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00214f
C464 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.SM 0.00168f
C465 XThR.Tn[14] VPWR 7.78627f
C466 XA.XIR[12].XIC[13].icell.PUM Vbias 0.0031f
C467 XThR.Tn[12] XA.XIR[13].XIC[8].icell.Ien 0.00338f
C468 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.03425f
C469 XA.XIR[11].XIC[0].icell.PDM VPWR 0.00799f
C470 XA.XIR[1].XIC[14].icell.Ien Iout 0.06417f
C471 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PUM 0.00102f
C472 XThC.Tn[5] Iout 0.83957f
C473 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.SM 0.0039f
C474 XA.XIR[4].XIC[7].icell.Ien Vbias 0.21098f
C475 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.SM 0.00168f
C476 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00584f
C477 XThC.Tn[5] XThR.Tn[9] 0.28739f
C478 XThC.Tn[1] XThR.Tn[8] 0.28739f
C479 XThR.Tn[7] XA.XIR[8].XIC[13].icell.SM 0.00121f
C480 XA.XIR[10].XIC[4].icell.PDM VPWR 0.00799f
C481 XA.XIR[10].XIC[12].icell.Ien VPWR 0.1903f
C482 XThR.XTB2.Y a_n1335_8107# 0.01006f
C483 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.SM 0.00168f
C484 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C485 XThR.Tn[5] XA.XIR[6].XIC[9].icell.SM 0.00121f
C486 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.0353f
C487 XThR.XTB6.Y a_n997_3979# 0.0046f
C488 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02762f
C489 bias[1] bias[0] 0.56718f
C490 XA.XIR[12].XIC[1].icell.Ien Iout 0.06417f
C491 XA.XIR[6].XIC[3].icell.SM VPWR 0.00158f
C492 XThR.Tn[13] XA.XIR[14].XIC[10].icell.Ien 0.00338f
C493 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.03425f
C494 VPWR data[1] 0.44103f
C495 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Ien 0.00232f
C496 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00214f
C497 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C498 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.15202f
C499 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C500 XA.XIR[13].XIC[13].icell.PUM VPWR 0.00937f
C501 XA.XIR[7].XIC[1].icell.Ien Vbias 0.21098f
C502 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.SM 0.00168f
C503 XA.XIR[15].XIC[6].icell.PUM VPWR 0.00937f
C504 XA.XIR[0].XIC[8].icell.PDM Vbias 0.04282f
C505 XA.XIR[5].XIC[6].icell.Ien VPWR 0.1903f
C506 XThC.XTB5.Y Vbias 0.01575f
C507 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PUM 0.00465f
C508 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.SM 0.00168f
C509 XThC.XTB7.B a_8739_9569# 0.0168f
C510 XThR.Tn[1] XA.XIR[2].XIC_15.icell.Ien 0.00117f
C511 XA.XIR[9].XIC[10].icell.Ien Vbias 0.21098f
C512 XA.XIR[5].XIC[2].icell.Ien Iout 0.06417f
C513 XA.XIR[10].XIC[4].icell.PUM Vbias 0.0031f
C514 XA.XIR[7].XIC[12].icell.PDM Iout 0.00117f
C515 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PUM 0.00465f
C516 XA.XIR[4].XIC[9].icell.PUM VPWR 0.00937f
C517 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.03425f
C518 XA.XIR[12].XIC[14].icell.Ien Vbias 0.21098f
C519 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00214f
C520 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.03425f
C521 XA.XIR[15].XIC[10].icell.PDM Iout 0.00117f
C522 XA.XIR[0].XIC[3].icell.Ien Vbias 0.21128f
C523 XThC.XTB3.Y XThC.Tn[7] 0.00819f
C524 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00214f
C525 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.SM 0.0039f
C526 XA.XIR[8].XIC[3].icell.PUM VPWR 0.00937f
C527 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.15202f
C528 XA.XIR[3].XIC[13].icell.PUM Vbias 0.0031f
C529 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C530 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00584f
C531 XThC.Tn[4] XThC.Tn[5] 0.4169f
C532 XThR.XTB2.Y a_n1049_7787# 0.2342f
C533 XA.XIR[0].XIC[12].icell.PDM VPWR 0.011f
C534 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02762f
C535 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.1106f
C536 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.SM 0.00168f
C537 XA.XIR[11].XIC[2].icell.SM VPWR 0.00158f
C538 XA.XIR[2].XIC[6].icell.PUM Vbias 0.0031f
C539 XA.XIR[7].XIC[6].icell.Ien Vbias 0.21098f
C540 XA.XIR[9].XIC[8].icell.PDM Iout 0.00117f
C541 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9] 0.00341f
C542 XA.XIR[13].XIC[14].icell.Ien VPWR 0.19036f
C543 XA.XIR[9].XIC[12].icell.PUM VPWR 0.00937f
C544 XThC.XTBN.Y Vbias 0.16321f
C545 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.SM 0.0039f
C546 XA.XIR[10].XIC[4].icell.SM VPWR 0.00158f
C547 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11] 0.00341f
C548 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00584f
C549 XA.XIR[1].XIC[8].icell.PUM Vbias 0.0031f
C550 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.03023f
C551 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02762f
C552 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.15202f
C553 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C554 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C555 XA.XIR[0].XIC[5].icell.PUM VPWR 0.00877f
C556 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04031f
C557 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Ien 0.00232f
C558 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C559 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C560 XThR.XTB6.Y a_n997_2891# 0.00466f
C561 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.SM 0.0039f
C562 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04031f
C563 XA.XIR[8].XIC_dummy_right.icell.PUM Vbias 0.00223f
C564 XA.XIR[3].XIC[13].icell.SM VPWR 0.00158f
C565 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C566 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C567 XThC.Tn[13] XThR.Tn[7] 0.2874f
C568 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.03425f
C569 XA.XIR[3].XIC[9].icell.SM Iout 0.00388f
C570 XA.XIR[1].XIC[13].icell.PDM Iout 0.00117f
C571 XThC.XTB7.B XThC.Tn[11] 0.03903f
C572 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.03425f
C573 XA.XIR[12].XIC[11].icell.PUM Vbias 0.0031f
C574 XA.XIR[6].XIC[14].icell.Ien Iout 0.06417f
C575 XA.XIR[2].XIC[6].icell.SM VPWR 0.00158f
C576 XA.XIR[7].XIC[8].icell.PUM VPWR 0.00937f
C577 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.SM 0.00168f
C578 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.SM 0.00168f
C579 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C580 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.SM 0.0039f
C581 XThC.Tn[10] Vbias 2.36503f
C582 XA.XIR[4].XIC[13].icell.PDM Iout 0.00117f
C583 XA.XIR[2].XIC[2].icell.SM Iout 0.00388f
C584 XA.XIR[1].XIC[8].icell.SM VPWR 0.00158f
C585 XA.XIR[10].XIC[10].icell.Ien VPWR 0.1903f
C586 XThR.Tn[1] XA.XIR[2].XIC[0].icell.SM 0.00121f
C587 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.SM 0.00168f
C588 a_4861_9615# Vbias 0.00548f
C589 XA.XIR[1].XIC[4].icell.SM Iout 0.00388f
C590 XA.XIR[14].XIC[8].icell.Ien Iout 0.06417f
C591 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C592 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00584f
C593 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PUM 0.00465f
C594 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.SM 0.00168f
C595 XA.XIR[15].XIC[12].icell.SM Vbias 0.00701f
C596 XThC.XTB3.Y a_3773_9615# 0.00124f
C597 XThR.XTBN.A a_n997_1579# 0.00199f
C598 XA.XIR[5].XIC[6].icell.PDM Vbias 0.04261f
C599 XA.XIR[13].XIC[11].icell.PUM VPWR 0.00937f
C600 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00584f
C601 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.15202f
C602 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.04036f
C603 XThR.Tn[11] XA.XIR[12].XIC[1].icell.SM 0.00121f
C604 XA.XIR[8].XIC[12].icell.SM Iout 0.00388f
C605 XThR.Tn[8] XA.XIR[9].XIC[12].icell.SM 0.00121f
C606 a_3773_9615# XThC.Tn[2] 0.01175f
C607 XThR.Tn[2] XA.XIR[3].XIC[7].icell.Ien 0.00338f
C608 XA.XIR[13].XIC[0].icell.PDM Vbias 0.04207f
C609 XThR.XTB3.Y VPWR 1.07975f
C610 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C611 XThR.Tn[4] XA.XIR[5].XIC[14].icell.Ien 0.00338f
C612 XThR.Tn[4] XA.XIR[4].XIC[6].icell.PDM 0.00341f
C613 XA.XIR[12].XIC[5].icell.PDM Vbias 0.04261f
C614 XA.XIR[12].XIC[12].icell.Ien Vbias 0.21098f
C615 XThC.Tn[12] XThR.Tn[3] 0.28739f
C616 XThR.XTB5.A XThR.XTB6.A 1.80461f
C617 XThR.Tn[3] XA.XIR[3].XIC[7].icell.PDM 0.00341f
C618 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C619 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Ien 0.00728f
C620 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PUM 0.00465f
C621 XThR.Tn[3] XA.XIR[4].XIC[14].icell.Ien 0.00338f
C622 XThC.XTB1.Y XThC.Tn[7] 0.0045f
C623 XThC.Tn[0] VPWR 5.9657f
C624 XThR.Tn[1] XA.XIR[2].XIC[5].icell.SM 0.00121f
C625 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.SM 0.00168f
C626 XA.XIR[6].XIC[3].icell.PDM VPWR 0.00799f
C627 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.04036f
C628 XThR.Tn[13] XA.XIR[14].XIC_15.icell.PDM 0.00172f
C629 XThR.Tn[13] XA.XIR[14].XIC_15.icell.Ien 0.00117f
C630 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.SM 0.0039f
C631 XA.XIR[0].XIC[14].icell.SM Iout 0.00367f
C632 XA.XIR[8].XIC[1].icell.Ien Vbias 0.21098f
C633 XA.XIR[14].XIC[0].icell.PDM VPWR 0.00799f
C634 XA.XIR[5].XIC[10].icell.PDM VPWR 0.00799f
C635 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PUM 0.00465f
C636 XThC.Tn[8] XThR.Tn[5] 0.28739f
C637 XA.XIR[3].XIC[3].icell.Ien Vbias 0.21098f
C638 XA.XIR[15].XIC_15.icell.PUM Vbias 0.0031f
C639 XA.XIR[13].XIC[4].icell.PDM VPWR 0.00799f
C640 XA.XIR[6].XIC[8].icell.PUM Vbias 0.0031f
C641 XA.XIR[13].XIC[12].icell.Ien VPWR 0.1903f
C642 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02762f
C643 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.03425f
C644 XThC.XTB7.Y a_7875_9569# 0.00476f
C645 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.SM 0.00168f
C646 XA.XIR[12].XIC[9].icell.PDM VPWR 0.00799f
C647 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C648 XA.XIR[15].XIC[9].icell.Ien Vbias 0.17899f
C649 XA.XIR[5].XIC[9].icell.SM Vbias 0.00701f
C650 XThR.Tn[0] XA.XIR[1].XIC[12].icell.SM 0.00121f
C651 XThC.XTB7.B data[1] 0.00593f
C652 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C653 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C654 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.03425f
C655 XA.XIR[9].XIC[2].icell.Ien VPWR 0.1903f
C656 XA.XIR[8].XIC[3].icell.PDM Vbias 0.04261f
C657 XA.XIR[3].XIC[1].icell.PDM Vbias 0.04261f
C658 XA.XIR[4].XIC[12].icell.Ien Vbias 0.21098f
C659 XA.XIR[11].XIC[3].icell.PDM Iout 0.00117f
C660 XThR.Tn[5] a_n1049_5317# 0.00158f
C661 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C662 a_6243_9615# XThC.Tn[5] 0.00158f
C663 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00214f
C664 XA.XIR[2].XIC[7].icell.PDM Vbias 0.04261f
C665 XThR.XTB6.A data[5] 0.37233f
C666 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.SM 0.0039f
C667 XA.XIR[13].XIC[4].icell.PUM Vbias 0.0031f
C668 XThR.Tn[5] XA.XIR[6].XIC[14].icell.SM 0.00121f
C669 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PUM 0.00102f
C670 XA.XIR[8].XIC[6].icell.Ien Vbias 0.21098f
C671 XThR.Tn[6] XA.XIR[7].XIC[1].icell.Ien 0.00338f
C672 XA.XIR[10].XIC[7].icell.PDM Iout 0.00117f
C673 XA.XIR[3].XIC[5].icell.PUM VPWR 0.00937f
C674 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04031f
C675 XA.XIR[12].XIC[4].icell.SM Vbias 0.00701f
C676 XA.XIR[6].XIC[8].icell.SM VPWR 0.00158f
C677 XA.XIR[6].XIC[4].icell.SM Iout 0.00388f
C678 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00584f
C679 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7] 0.00341f
C680 XA.XIR[5].XIC[11].icell.Ien VPWR 0.1903f
C681 XA.XIR[11].XIC[7].icell.PUM Vbias 0.0031f
C682 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PUM 0.00465f
C683 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.SM 0.0039f
C684 XA.XIR[9].XIC_15.icell.Ien Vbias 0.21234f
C685 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PUM 0.00441f
C686 XA.XIR[5].XIC[7].icell.Ien Iout 0.06417f
C687 XA.XIR[15].XIC[10].icell.SM Vbias 0.00701f
C688 XA.XIR[3].XIC[5].icell.PDM VPWR 0.00799f
C689 XA.XIR[8].XIC[7].icell.PDM VPWR 0.00799f
C690 XA.XIR[10].XIC[9].icell.PUM Vbias 0.0031f
C691 XA.XIR[4].XIC[14].icell.PUM VPWR 0.00937f
C692 XThR.Tn[14] XA.XIR[15].XIC[1].icell.Ien 0.00338f
C693 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.SM 0.00168f
C694 XA.XIR[14].XIC[2].icell.SM VPWR 0.00158f
C695 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C696 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00214f
C697 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC_15.icell.Ien 0.00214f
C698 XA.XIR[2].XIC[11].icell.PDM VPWR 0.00799f
C699 XA.XIR[0].XIC[8].icell.Ien Vbias 0.2113f
C700 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C701 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04031f
C702 XThC.Tn[14] XThR.Tn[2] 0.28745f
C703 XA.XIR[13].XIC[4].icell.SM VPWR 0.00158f
C704 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PUM 0.00465f
C705 XA.XIR[8].XIC[8].icell.PUM VPWR 0.00937f
C706 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C707 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00584f
C708 XThR.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.00338f
C709 XA.XIR[12].XIC[6].icell.Ien VPWR 0.1903f
C710 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00214f
C711 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12] 0.00341f
C712 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.03425f
C713 XA.XIR[12].XIC[10].icell.Ien Vbias 0.21098f
C714 XA.XIR[10].XIC_15.icell.Ien VPWR 0.25566f
C715 XA.XIR[11].XIC[7].icell.SM VPWR 0.00158f
C716 XThR.XTB6.Y a_n997_1579# 0.07626f
C717 XA.XIR[12].XIC[2].icell.Ien Iout 0.06417f
C718 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.SM 0.00168f
C719 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00214f
C720 XA.XIR[2].XIC[11].icell.PUM Vbias 0.0031f
C721 XA.XIR[7].XIC[11].icell.Ien Vbias 0.21098f
C722 XThR.Tn[4] XA.XIR[5].XIC[4].icell.SM 0.00121f
C723 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.03425f
C724 XA.XIR[11].XIC[3].icell.SM Iout 0.00388f
C725 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C726 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.SM 0.00168f
C727 XA.XIR[1].XIC[13].icell.PUM Vbias 0.0031f
C728 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C729 XThR.Tn[3] XA.XIR[4].XIC[4].icell.SM 0.00121f
C730 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.15202f
C731 XThR.Tn[14] XA.XIR[15].XIC[6].icell.Ien 0.00338f
C732 XA.XIR[0].XIC[10].icell.PUM VPWR 0.00877f
C733 XA.XIR[10].XIC[5].icell.SM Iout 0.00388f
C734 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C735 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00214f
C736 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.SM 0.00168f
C737 XThR.Tn[9] XA.XIR[10].XIC[5].icell.SM 0.00121f
C738 XA.XIR[15].XIC[13].icell.PUM Vbias 0.0031f
C739 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5] 0.00346f
C740 XThR.Tn[8] Vbias 3.74624f
C741 XA.XIR[13].XIC[10].icell.Ien VPWR 0.1903f
C742 XA.XIR[3].XIC[0].icell.Ien Vbias 0.20951f
C743 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04031f
C744 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04031f
C745 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C746 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C747 XThC.Tn[10] XThR.Tn[6] 0.28739f
C748 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PUM 0.00465f
C749 XA.XIR[3].XIC[14].icell.SM Iout 0.00388f
C750 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8] 0.00341f
C751 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04031f
C752 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00584f
C753 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[9].icell.SM 0.0039f
C754 XA.XIR[7].XIC[13].icell.PUM VPWR 0.00937f
C755 XA.XIR[2].XIC[11].icell.SM VPWR 0.00158f
C756 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PUM 0.00465f
C757 XA.XIR[11].XIC[1].icell.Ien Vbias 0.21098f
C758 XA.XIR[2].XIC_15.icell.SM Vbias 0.00701f
C759 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C760 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C761 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00214f
C762 XA.XIR[1].XIC[13].icell.SM VPWR 0.00158f
C763 XA.XIR[2].XIC[7].icell.SM Iout 0.00388f
C764 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PUM 0.00179f
C765 XThC.Tn[12] XThR.Tn[11] 0.28739f
C766 XA.XIR[7].XIC[7].icell.PDM Vbias 0.04261f
C767 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.04036f
C768 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C769 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.SM 0.0039f
C770 XA.XIR[9].XIC[0].icell.SM Vbias 0.00675f
C771 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PUM 0.00465f
C772 XThR.Tn[12] XA.XIR[13].XIC[3].icell.SM 0.00121f
C773 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.SM 0.00168f
C774 XA.XIR[1].XIC[9].icell.SM Iout 0.00388f
C775 XThC.Tn[2] XThR.Tn[7] 0.28739f
C776 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04052f
C777 XThR.XTB6.A XThR.Tn[9] 0.00838f
C778 XA.XIR[4].XIC[2].icell.SM Vbias 0.00701f
C779 XA.XIR[6].XIC[14].icell.PDM Vbias 0.04261f
C780 XA.XIR[15].XIC[5].icell.PDM Vbias 0.04261f
C781 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.15202f
C782 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.SM 0.00168f
C783 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C784 XA.XIR[3].XIC[2].icell.PUM VPWR 0.00937f
C785 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00214f
C786 XThC.XTB7.B XThC.Tn[0] 0.00139f
C787 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C788 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.15202f
C789 XA.XIR[12].XIC[0].icell.SM VPWR 0.00158f
C790 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.SM 0.00168f
C791 XThR.Tn[11] XA.XIR[12].XIC[6].icell.SM 0.00121f
C792 XA.XIR[15].XIC[14].icell.Ien Vbias 0.17899f
C793 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C794 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00584f
C795 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00584f
C796 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C797 XThC.XTB6.Y XThC.Tn[8] 0.02461f
C798 XThC.XTB5.Y XThC.Tn[13] 0.00145f
C799 XThR.Tn[2] XA.XIR[3].XIC[12].icell.Ien 0.00338f
C800 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.03425f
C801 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.SM 0.0039f
C802 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04052f
C803 XA.XIR[9].XIC[3].icell.PDM Vbias 0.04261f
C804 a_7651_9569# Vbias 0.00376f
C805 XThR.XTB7.A data[6] 0.00197f
C806 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C807 XThR.Tn[0] Iout 1.16239f
C808 XA.XIR[5].XIC[1].icell.SM VPWR 0.00158f
C809 XThR.XTB7.Y a_n1319_5317# 0.01283f
C810 XA.XIR[7].XIC[11].icell.PDM VPWR 0.00799f
C811 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.15202f
C812 XThC.XTB6.A a_7875_9569# 0.00149f
C813 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PUM 0.00465f
C814 XA.XIR[9].XIC[5].icell.SM Vbias 0.00701f
C815 XThR.Tn[1] XA.XIR[2].XIC[10].icell.SM 0.00121f
C816 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02762f
C817 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C818 a_n1049_6699# XThR.Tn[4] 0.00158f
C819 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00214f
C820 XA.XIR[15].XIC[9].icell.PDM VPWR 0.0114f
C821 XA.XIR[4].XIC[4].icell.Ien VPWR 0.1903f
C822 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02762f
C823 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PUM 0.00465f
C824 XA.XIR[6].XIC[6].icell.PDM Iout 0.00117f
C825 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Ien 0.00553f
C826 XA.XIR[3].XIC[8].icell.Ien Vbias 0.21098f
C827 XA.XIR[5].XIC[13].icell.PDM Iout 0.00117f
C828 XA.XIR[14].XIC[3].icell.PDM Iout 0.00117f
C829 XA.XIR[1].XIC[8].icell.PDM Vbias 0.04261f
C830 XA.XIR[6].XIC[13].icell.PUM Vbias 0.0031f
C831 XThC.Tn[1] XThR.Tn[3] 0.28739f
C832 a_9827_9569# VPWR 0.0017f
C833 XA.XIR[9].XIC[7].icell.PDM VPWR 0.00799f
C834 XA.XIR[13].XIC[7].icell.PDM Iout 0.00117f
C835 XThC.XTBN.Y XThC.Tn[13] 0.62331f
C836 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.SM 0.00168f
C837 XThC.Tn[10] XThR.Tn[4] 0.28739f
C838 XA.XIR[7].XIC[1].icell.SM Vbias 0.00701f
C839 XA.XIR[4].XIC[8].icell.PDM Vbias 0.04261f
C840 XA.XIR[5].XIC[14].icell.SM Vbias 0.00701f
C841 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C842 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C843 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00214f
C844 XA.XIR[15].XIC[11].icell.PUM Vbias 0.0031f
C845 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00584f
C846 XA.XIR[9].XIC[7].icell.Ien VPWR 0.1903f
C847 XA.XIR[1].XIC[3].icell.Ien Vbias 0.21104f
C848 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C849 XThC.XTB4.Y XThC.Tn[8] 0.01306f
C850 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00584f
C851 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C852 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C853 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00584f
C854 XA.XIR[14].XIC[7].icell.PUM Vbias 0.0031f
C855 XThC.Tn[0] XA.XIR[5].XIC_dummy_left.icell.Iout 0.00109f
C856 XA.XIR[9].XIC[3].icell.Ien Iout 0.06417f
C857 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.15202f
C858 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.SM 0.00168f
C859 XA.XIR[12].XIC_15.icell.Ien Vbias 0.21234f
C860 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C861 XThC.Tn[14] XThR.Tn[10] 0.28745f
C862 XThC.Tn[4] XThR.Tn[0] 0.28741f
C863 XA.XIR[13].XIC[9].icell.PUM Vbias 0.0031f
C864 XThC.Tn[6] XThR.Tn[5] 0.28739f
C865 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04031f
C866 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02762f
C867 XA.XIR[8].XIC[11].icell.Ien Vbias 0.21098f
C868 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00214f
C869 XA.XIR[3].XIC[10].icell.PUM VPWR 0.00937f
C870 XA.XIR[1].XIC[12].icell.PDM VPWR 0.008f
C871 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C872 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C873 XA.XIR[6].XIC[13].icell.SM VPWR 0.00158f
C874 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.03504f
C875 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14] 0.00341f
C876 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C877 XThC.Tn[11] XThC.Tn[12] 0.22144f
C878 XA.XIR[1].XIC[0].icell.PDM Iout 0.00117f
C879 XA.XIR[6].XIC[9].icell.SM Iout 0.00388f
C880 XA.XIR[2].XIC[3].icell.PUM VPWR 0.00937f
C881 XA.XIR[4].XIC[12].icell.PDM VPWR 0.00799f
C882 XA.XIR[7].XIC[3].icell.Ien VPWR 0.1903f
C883 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04031f
C884 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C885 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C886 XA.XIR[1].XIC[5].icell.PUM VPWR 0.00937f
C887 XA.XIR[5].XIC[12].icell.Ien Iout 0.06417f
C888 XA.XIR[4].XIC[0].icell.PDM Iout 0.00117f
C889 XThC.XTB7.B VPWR 1.32988f
C890 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C891 XA.XIR[13].XIC_15.icell.Ien VPWR 0.25566f
C892 XA.XIR[14].XIC[7].icell.SM VPWR 0.00158f
C893 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C894 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Iout 0.00347f
C895 XA.XIR[8].XIC[10].icell.PDM Iout 0.00117f
C896 XA.XIR[15].XIC[12].icell.Ien Vbias 0.17899f
C897 XA.XIR[3].XIC[8].icell.PDM Iout 0.00117f
C898 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C899 XA.XIR[14].XIC[3].icell.SM Iout 0.00388f
C900 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04031f
C901 XA.XIR[0].XIC[13].icell.Ien Vbias 0.2113f
C902 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00584f
C903 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[9].icell.Ien 0.00214f
C904 XThC.XTB5.Y data[3] 0.00931f
C905 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04031f
C906 XA.XIR[8].XIC[13].icell.PUM VPWR 0.00937f
C907 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C908 XThR.Tn[6] XA.XIR[7].XIC[11].icell.Ien 0.00338f
C909 XA.XIR[2].XIC[14].icell.PDM Iout 0.00117f
C910 XA.XIR[13].XIC[5].icell.SM Iout 0.00388f
C911 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.SM 0.00168f
C912 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.SM 0.0039f
C913 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.03592f
C914 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00584f
C915 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C916 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.15202f
C917 XThR.Tn[0] XA.XIR[0].XIC[11].icell.PDM 0.00341f
C918 XThR.Tn[2] XA.XIR[3].XIC[2].icell.SM 0.00121f
C919 XA.XIR[12].XIC[7].icell.Ien Iout 0.06417f
C920 XThR.XTBN.A XThR.Tn[8] 0.1369f
C921 XA.XIR[2].XIC_dummy_right.icell.PUM Vbias 0.00223f
C922 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02762f
C923 XThR.Tn[4] XA.XIR[5].XIC[9].icell.SM 0.00121f
C924 XA.XIR[10].XIC_dummy_right.icell.SM VPWR 0.00123f
C925 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.SM 0.00168f
C926 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.SM 0.00168f
C927 XThR.Tn[1] XA.XIR[1].XIC[9].icell.PDM 0.00341f
C928 XA.XIR[11].XIC[8].icell.SM Iout 0.00388f
C929 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00584f
C930 VPWR bias[0] 2.10172f
C931 XThC.Tn[3] XThR.Tn[2] 0.28739f
C932 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04031f
C933 XThR.Tn[3] XA.XIR[4].XIC[9].icell.SM 0.00121f
C934 XA.XIR[14].XIC[1].icell.Ien Vbias 0.21098f
C935 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.04036f
C936 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.15202f
C937 XThC.XTB7.Y a_6243_9615# 0.27822f
C938 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01499f
C939 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PUM 0.00465f
C940 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C941 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.15202f
C942 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5] 0.00341f
C943 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.04036f
C944 XThC.Tn[12] XThR.Tn[14] 0.28739f
C945 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.15202f
C946 XA.XIR[10].XIC[2].icell.PDM Vbias 0.04261f
C947 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02762f
C948 XThR.Tn[2] XA.XIR[2].XIC[6].icell.PDM 0.00341f
C949 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C950 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00214f
C951 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04031f
C952 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.03425f
C953 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.SM 0.00168f
C954 XThR.XTB7.B data[6] 0.07481f
C955 XA.XIR[6].XIC[3].icell.Ien Vbias 0.21098f
C956 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.15202f
C957 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Ien 0.00584f
C958 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C959 XThC.XTB2.Y XThC.Tn[8] 0.00167f
C960 XA.XIR[15].XIC[1].icell.Ien VPWR 0.32895f
C961 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00214f
C962 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PUM 0.00465f
C963 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11117f
C964 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6] 0.00341f
C965 XA.XIR[2].XIC[12].icell.SM Iout 0.00388f
C966 XA.XIR[15].XIC[4].icell.SM Vbias 0.00701f
C967 XA.XIR[5].XIC[6].icell.PUM Vbias 0.0031f
C968 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C969 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.03425f
C970 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12] 0.00341f
C971 XA.XIR[1].XIC[0].icell.Ien Iout 0.06411f
C972 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C973 XThR.Tn[12] XA.XIR[13].XIC[8].icell.SM 0.00121f
C974 XA.XIR[11].XIC[2].icell.PDM VPWR 0.00799f
C975 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Iout 0.00347f
C976 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.SM 0.0039f
C977 XA.XIR[1].XIC[14].icell.SM Iout 0.00388f
C978 XA.XIR[4].XIC[7].icell.SM Vbias 0.00701f
C979 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00584f
C980 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C981 XA.XIR[4].XIC[0].icell.Ien Iout 0.06411f
C982 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PUM 0.00186f
C983 XA.XIR[10].XIC[6].icell.PDM VPWR 0.00799f
C984 XThR.Tn[1] Iout 1.16236f
C985 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PUM 0.00429f
C986 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PUM 0.00179f
C987 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00584f
C988 XThC.XTBN.A XThC.Tn[10] 0.12148f
C989 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C990 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02762f
C991 XA.XIR[0].XIC_15.icell.SM Iout 0.00367f
C992 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C993 XA.XIR[8].XIC[1].icell.SM Vbias 0.00701f
C994 XThC.Tn[1] XThR.Tn[11] 0.28739f
C995 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02762f
C996 XThR.Tn[12] Iout 1.16233f
C997 XA.XIR[6].XIC[5].icell.PUM VPWR 0.00937f
C998 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C999 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C1000 XA.XIR[2].XIC[1].icell.Ien Vbias 0.21098f
C1001 XA.XIR[0].XIC[10].icell.PDM Vbias 0.04282f
C1002 XA.XIR[15].XIC[6].icell.Ien VPWR 0.32895f
C1003 XA.XIR[11].XIC[2].icell.Ien Vbias 0.21098f
C1004 XA.XIR[5].XIC[6].icell.SM VPWR 0.00158f
C1005 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.03425f
C1006 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Ien 0.00232f
C1007 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.15202f
C1008 XThC.XTB7.B a_9827_9569# 0.00228f
C1009 XA.XIR[15].XIC[10].icell.Ien Vbias 0.17899f
C1010 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00214f
C1011 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00584f
C1012 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.02762f
C1013 XA.XIR[9].XIC[10].icell.SM Vbias 0.00701f
C1014 XA.XIR[15].XIC[2].icell.Ien Iout 0.06807f
C1015 XThC.XTB7.A Vbias 0.0149f
C1016 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C1017 XA.XIR[7].XIC[14].icell.PDM Iout 0.00117f
C1018 XA.XIR[10].XIC[4].icell.Ien Vbias 0.21098f
C1019 XA.XIR[5].XIC[2].icell.SM Iout 0.00388f
C1020 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C1021 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.03425f
C1022 XA.XIR[4].XIC[9].icell.Ien VPWR 0.1903f
C1023 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18966f
C1024 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.SM 0.0039f
C1025 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PUM 0.00465f
C1026 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C1027 XA.XIR[4].XIC[5].icell.Ien Iout 0.06417f
C1028 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.03425f
C1029 XA.XIR[0].XIC[3].icell.SM Vbias 0.00716f
C1030 XA.XIR[8].XIC[3].icell.Ien VPWR 0.1903f
C1031 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C1032 XThC.XTB6.Y XThC.Tn[6] 0.00689f
C1033 XThR.Tn[6] XA.XIR[7].XIC[1].icell.SM 0.00121f
C1034 XA.XIR[3].XIC[13].icell.Ien Vbias 0.21098f
C1035 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C1036 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02762f
C1037 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C1038 XA.XIR[12].XIC[1].icell.SM VPWR 0.00158f
C1039 XThC.Tn[14] XThR.Tn[13] 0.28745f
C1040 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02762f
C1041 XA.XIR[0].XIC[14].icell.PDM VPWR 0.00783f
C1042 XThC.Tn[4] XThR.Tn[1] 0.2874f
C1043 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C1044 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PUM 0.0047f
C1045 XA.XIR[11].XIC[4].icell.PUM VPWR 0.00937f
C1046 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00214f
C1047 XThC.Tn[8] Iout 0.8379f
C1048 XA.XIR[9].XIC[10].icell.PDM Iout 0.00117f
C1049 XA.XIR[2].XIC[6].icell.Ien Vbias 0.21098f
C1050 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.SM 0.0039f
C1051 XA.XIR[7].XIC[6].icell.SM Vbias 0.00701f
C1052 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9] 0.00341f
C1053 XThC.Tn[8] XThR.Tn[9] 0.28739f
C1054 XA.XIR[9].XIC[12].icell.Ien VPWR 0.1903f
C1055 XA.XIR[10].XIC[6].icell.PUM VPWR 0.00937f
C1056 XA.XIR[9].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1057 XA.XIR[1].XIC[8].icell.Ien Vbias 0.21104f
C1058 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11] 0.00341f
C1059 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PUM 0.00465f
C1060 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C1061 XThR.Tn[14] XA.XIR[15].XIC[1].icell.SM 0.00121f
C1062 XThC.Tn[4] XThR.Tn[12] 0.28739f
C1063 XA.XIR[9].XIC[8].icell.Ien Iout 0.06417f
C1064 XThC.Tn[13] XThR.Tn[8] 0.2874f
C1065 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.15202f
C1066 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.SM 0.00168f
C1067 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18987f
C1068 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C1069 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[8].icell.Ien 0.00214f
C1070 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.SM 0.0039f
C1071 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04031f
C1072 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C1073 XThR.XTBN.A a_n997_3755# 0.01939f
C1074 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01577f
C1075 XThC.XTBN.Y XThC.Tn[2] 0.64352f
C1076 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Ien 0.00246f
C1077 XA.XIR[11].XIC[13].icell.SM Iout 0.00388f
C1078 XThR.XTB7.A XThR.Tn[5] 0.02751f
C1079 XA.XIR[1].XIC_15.icell.PDM Iout 0.00133f
C1080 XA.XIR[2].XIC[8].icell.PUM VPWR 0.00937f
C1081 XA.XIR[6].XIC[14].icell.SM Iout 0.00388f
C1082 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Ien 0.00214f
C1083 XA.XIR[7].XIC[8].icell.Ien VPWR 0.1903f
C1084 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C1085 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1086 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C1087 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C1088 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00584f
C1089 XThC.Tn[0] XA.XIR[12].XIC_dummy_left.icell.Iout 0.00109f
C1090 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[4].icell.Ien 0.00214f
C1091 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.Ien 0.00584f
C1092 XA.XIR[4].XIC_15.icell.PDM Iout 0.00133f
C1093 XA.XIR[0].XIC[0].icell.PUM VPWR 0.00877f
C1094 XA.XIR[1].XIC[10].icell.PUM VPWR 0.00937f
C1095 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.SM 0.0039f
C1096 XThC.XTB4.Y XThC.Tn[6] 0.00608f
C1097 XA.XIR[7].XIC[4].icell.Ien Iout 0.06417f
C1098 XThC.Tn[3] XThR.Tn[10] 0.28739f
C1099 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.04036f
C1100 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04031f
C1101 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02762f
C1102 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02762f
C1103 XThC.XTB3.Y XThC.Tn[10] 0.29462f
C1104 XA.XIR[13].XIC_dummy_right.icell.SM VPWR 0.00123f
C1105 a_5949_9615# Vbias 0.00634f
C1106 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.PDM 0.00591f
C1107 XA.XIR[14].XIC[8].icell.SM Iout 0.00388f
C1108 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.03425f
C1109 XA.XIR[6].XIC[1].icell.PDM Vbias 0.04261f
C1110 XThR.Tn[7] XA.XIR[8].XIC[5].icell.Ien 0.00338f
C1111 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.SM 0.0039f
C1112 XThC.XTB3.Y a_4861_9615# 0.0093f
C1113 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00584f
C1114 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00214f
C1115 XA.XIR[5].XIC[8].icell.PDM Vbias 0.04261f
C1116 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PUM 0.00465f
C1117 a_n1049_5611# XThR.Tn[6] 0.00158f
C1118 XThR.Tn[2] XA.XIR[3].XIC[7].icell.SM 0.00121f
C1119 XA.XIR[3].XIC_15.icell.SM Iout 0.0047f
C1120 XThR.Tn[12] XA.XIR[13].XIC[13].icell.SM 0.00121f
C1121 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00584f
C1122 XA.XIR[13].XIC[2].icell.PDM Vbias 0.04261f
C1123 a_n1049_8581# VPWR 0.71705f
C1124 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.SM 0.0039f
C1125 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00214f
C1126 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C1127 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.SM 0.00168f
C1128 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04031f
C1129 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.15202f
C1130 XThC.XTB5.A Vbias 0.00557f
C1131 XThR.Tn[3] Vbias 3.74868f
C1132 XThR.Tn[4] XA.XIR[4].XIC[8].icell.PDM 0.00341f
C1133 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C1134 XThR.Tn[4] XA.XIR[5].XIC[14].icell.SM 0.00121f
C1135 XA.XIR[12].XIC[7].icell.PDM Vbias 0.04261f
C1136 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12] 0.00341f
C1137 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.03425f
C1138 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C1139 XA.XIR[10].XIC[0].icell.Ien VPWR 0.1903f
C1140 XThR.Tn[3] XA.XIR[4].XIC[14].icell.SM 0.00121f
C1141 XThR.Tn[3] XA.XIR[3].XIC[9].icell.PDM 0.00341f
C1142 XThR.Tn[10] XA.XIR[11].XIC[6].icell.Ien 0.00338f
C1143 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C1144 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C1145 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.03425f
C1146 XA.XIR[6].XIC[5].icell.PDM VPWR 0.00799f
C1147 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00214f
C1148 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C1149 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.15202f
C1150 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PDM 0.00172f
C1151 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.03425f
C1152 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.15202f
C1153 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.SM 0.00168f
C1154 XA.XIR[14].XIC[2].icell.PDM VPWR 0.00799f
C1155 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.SM 0.00168f
C1156 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.15202f
C1157 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C1158 XA.XIR[5].XIC[12].icell.PDM VPWR 0.00799f
C1159 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00584f
C1160 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PUM 0.00465f
C1161 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C1162 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.03425f
C1163 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PUM 0.00465f
C1164 XThR.XTB4.Y data[6] 0.0086f
C1165 XA.XIR[10].XIC[12].icell.SM Vbias 0.00701f
C1166 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C1167 XA.XIR[13].XIC[6].icell.PDM VPWR 0.00799f
C1168 XA.XIR[15].XIC_15.icell.Ien Vbias 0.17891f
C1169 XA.XIR[5].XIC[0].icell.PDM Iout 0.00117f
C1170 XA.XIR[3].XIC[3].icell.SM Vbias 0.00701f
C1171 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC[14].icell.SM 0.0039f
C1172 XA.XIR[6].XIC[8].icell.Ien Vbias 0.21098f
C1173 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.15202f
C1174 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.Ien 0.00584f
C1175 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PUM 0.00465f
C1176 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00214f
C1177 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.03425f
C1178 XThC.XTB7.Y a_8963_9569# 0.00474f
C1179 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C1180 XA.XIR[5].XIC[11].icell.PUM Vbias 0.0031f
C1181 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02762f
C1182 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.SM 0.0039f
C1183 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C1184 XThC.Tn[1] XThR.Tn[14] 0.28739f
C1185 XA.XIR[9].XIC[2].icell.SM VPWR 0.00158f
C1186 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01432f
C1187 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C1188 XA.XIR[0].XIC_dummy_left.icell.SM VPWR 0.00269f
C1189 XA.XIR[8].XIC[5].icell.PDM Vbias 0.04261f
C1190 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02893f
C1191 XA.XIR[4].XIC[12].icell.SM Vbias 0.00701f
C1192 XA.XIR[3].XIC[3].icell.PDM Vbias 0.04261f
C1193 XThR.XTB2.Y a_n1049_7493# 0.02133f
C1194 XA.XIR[14].XIC[2].icell.Ien Vbias 0.21098f
C1195 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00214f
C1196 XThR.Tn[7] XA.XIR[8].XIC[0].icell.Ien 0.00338f
C1197 XA.XIR[11].XIC[5].icell.PDM Iout 0.00117f
C1198 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.SM 0.00168f
C1199 XA.XIR[11].XIC[11].icell.SM Iout 0.00388f
C1200 XA.XIR[2].XIC[9].icell.PDM Vbias 0.04261f
C1201 XA.XIR[13].XIC[4].icell.Ien Vbias 0.21098f
C1202 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C1203 XA.XIR[8].XIC[6].icell.SM Vbias 0.00701f
C1204 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C1205 XA.XIR[10].XIC[9].icell.PDM Iout 0.00117f
C1206 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04031f
C1207 XA.XIR[3].XIC[5].icell.Ien VPWR 0.1903f
C1208 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00584f
C1209 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.11103f
C1210 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.SM 0.00168f
C1211 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.03425f
C1212 XA.XIR[6].XIC[10].icell.PUM VPWR 0.00937f
C1213 XA.XIR[12].XIC[6].icell.PUM Vbias 0.0031f
C1214 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C1215 XThR.XTB6.Y a_n997_3755# 0.0046f
C1216 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00584f
C1217 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00214f
C1218 XA.XIR[10].XIC_15.icell.PUM Vbias 0.0031f
C1219 XA.XIR[11].XIC[7].icell.Ien Vbias 0.21098f
C1220 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.03425f
C1221 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[3].icell.Ien 0.00214f
C1222 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02762f
C1223 XA.XIR[5].XIC[11].icell.SM VPWR 0.00158f
C1224 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7] 0.00341f
C1225 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C1226 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C1227 XA.XIR[5].XIC_15.icell.SM Vbias 0.00701f
C1228 XThR.Tn[10] XA.XIR[11].XIC[0].icell.SM 0.00121f
C1229 XThC.Tn[12] VPWR 6.85795f
C1230 XA.XIR[15].XIC[7].icell.Ien Iout 0.06807f
C1231 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C1232 XA.XIR[10].XIC[9].icell.Ien Vbias 0.21098f
C1233 XA.XIR[4].XIC[14].icell.Ien VPWR 0.19036f
C1234 XA.XIR[5].XIC[7].icell.SM Iout 0.00388f
C1235 XA.XIR[3].XIC[7].icell.PDM VPWR 0.00799f
C1236 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.03549f
C1237 XA.XIR[8].XIC[9].icell.PDM VPWR 0.00799f
C1238 XA.XIR[14].XIC[4].icell.PUM VPWR 0.00937f
C1239 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C1240 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00584f
C1241 XA.XIR[4].XIC[10].icell.Ien Iout 0.06417f
C1242 XA.XIR[0].XIC[8].icell.SM Vbias 0.00716f
C1243 XA.XIR[2].XIC[13].icell.PDM VPWR 0.00799f
C1244 XThC.XTBN.A a_7651_9569# 0.02087f
C1245 XA.XIR[13].XIC[6].icell.PUM VPWR 0.00937f
C1246 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.SM 0.0039f
C1247 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04031f
C1248 XA.XIR[0].XIC[1].icell.Ien Iout 0.06389f
C1249 XThR.Tn[12] XA.XIR[13].XIC[11].icell.SM 0.00121f
C1250 XA.XIR[8].XIC[8].icell.Ien VPWR 0.1903f
C1251 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.03426f
C1252 XA.XIR[12].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1253 XThR.Tn[6] XA.XIR[7].XIC[6].icell.SM 0.00121f
C1254 XA.XIR[2].XIC[1].icell.PDM Iout 0.00117f
C1255 XA.XIR[12].XIC[6].icell.SM VPWR 0.00158f
C1256 a_n1049_7787# XThR.XTB3.Y 0.00124f
C1257 XA.XIR[8].XIC[4].icell.Ien Iout 0.06417f
C1258 XThR.XTB7.B XThR.Tn[5] 0.00705f
C1259 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12] 0.00341f
C1260 XThR.XTB6.Y a_n1049_5611# 0.26831f
C1261 XThR.Tn[8] XA.XIR[9].XIC[4].icell.Ien 0.00338f
C1262 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C1263 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07214f
C1264 XA.XIR[15].XIC_dummy_left.icell.Ien Vbias 0.00329f
C1265 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C1266 XA.XIR[12].XIC[2].icell.SM Iout 0.00388f
C1267 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C1268 XA.XIR[11].XIC[9].icell.PUM VPWR 0.00937f
C1269 XA.XIR[2].XIC[11].icell.Ien Vbias 0.21098f
C1270 XA.XIR[7].XIC[11].icell.SM Vbias 0.00701f
C1271 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00214f
C1272 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.39105f
C1273 XA.XIR[14].XIC[13].icell.SM Iout 0.00388f
C1274 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04031f
C1275 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.PDM 0.00586f
C1276 XA.XIR[1].XIC[13].icell.Ien Vbias 0.21104f
C1277 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00584f
C1278 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1279 XThR.Tn[14] XA.XIR[15].XIC[6].icell.SM 0.00121f
C1280 XA.XIR[9].XIC[13].icell.Ien Iout 0.06417f
C1281 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00584f
C1282 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.15202f
C1283 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18966f
C1284 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5] 0.00341f
C1285 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C1286 XA.XIR[10].XIC[10].icell.SM Vbias 0.00701f
C1287 XThC.Tn[3] XThR.Tn[13] 0.28739f
C1288 XA.XIR[3].XIC[0].icell.SM Vbias 0.00675f
C1289 bias[1] Vbias 0.05009f
C1290 XA.XIR[0].XIC[6].icell.Ien Iout 0.06389f
C1291 XThR.Tn[5] XA.XIR[6].XIC[1].icell.Ien 0.00338f
C1292 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04031f
C1293 XA.XIR[12].XIC[0].icell.Ien Vbias 0.20951f
C1294 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.SM 0.0039f
C1295 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.03425f
C1296 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04031f
C1297 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8] 0.00341f
C1298 XThC.Tn[6] Iout 0.83892f
C1299 XA.XIR[2].XIC[13].icell.PUM VPWR 0.00937f
C1300 XA.XIR[7].XIC[13].icell.Ien VPWR 0.1903f
C1301 XThC.Tn[6] XThR.Tn[9] 0.28739f
C1302 XThR.Tn[11] Vbias 3.74874f
C1303 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12] 0.00341f
C1304 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02762f
C1305 XThC.Tn[2] XThR.Tn[8] 0.28739f
C1306 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.15202f
C1307 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6] 0.00341f
C1308 XA.XIR[10].XIC_dummy_left.icell.SM VPWR 0.00269f
C1309 XA.XIR[7].XIC[9].icell.Ien Iout 0.06417f
C1310 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.SM 0.0039f
C1311 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01577f
C1312 XThR.Tn[0] XA.XIR[1].XIC[4].icell.Ien 0.00338f
C1313 XThR.Tn[7] XA.XIR[8].XIC_15.icell.PDM 0.00172f
C1314 XA.XIR[7].XIC[9].icell.PDM Vbias 0.04261f
C1315 XA.XIR[9].XIC[2].icell.PUM Vbias 0.0031f
C1316 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.SM 0.00168f
C1317 XA.XIR[11].XIC[9].icell.SM Iout 0.00388f
C1318 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.03425f
C1319 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C1320 XA.XIR[4].XIC[4].icell.PUM Vbias 0.0031f
C1321 XA.XIR[15].XIC[7].icell.PDM Vbias 0.04261f
C1322 XA.XIR[13].XIC[0].icell.Ien VPWR 0.1903f
C1323 XThR.Tn[7] XA.XIR[8].XIC[10].icell.Ien 0.00338f
C1324 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C1325 XThC.XTBN.Y a_2979_9615# 0.0607f
C1326 XA.XIR[10].XIC[13].icell.PUM Vbias 0.0031f
C1327 XA.XIR[12].XIC[2].icell.PUM VPWR 0.00937f
C1328 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C1329 XThR.Tn[5] XA.XIR[6].XIC[6].icell.Ien 0.00338f
C1330 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.SM 0.00168f
C1331 XThR.XTBN.A data[4] 0.02581f
C1332 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00584f
C1333 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C1334 XThR.Tn[2] XA.XIR[3].XIC[12].icell.SM 0.00121f
C1335 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Iout 0.00347f
C1336 a_8739_9569# Vbias 0.00278f
C1337 XA.XIR[2].XIC[0].icell.Ien Iout 0.06411f
C1338 XA.XIR[9].XIC[5].icell.PDM Vbias 0.04261f
C1339 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.15202f
C1340 data[2] data[3] 0.04128f
C1341 XThR.XTB5.A XThR.XTB7.A 0.07862f
C1342 XA.XIR[15].XIC[1].icell.SM VPWR 0.00158f
C1343 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00214f
C1344 XA.XIR[5].XIC[3].icell.PUM VPWR 0.00937f
C1345 XA.XIR[13].XIC[12].icell.SM Vbias 0.00701f
C1346 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00584f
C1347 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C1348 a_9827_9569# XThC.Tn[12] 0.19481f
C1349 XA.XIR[7].XIC[13].icell.PDM VPWR 0.00799f
C1350 XThC.XTB3.Y a_7651_9569# 0.00604f
C1351 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.03425f
C1352 XThC.XTB6.A data[0] 0.48493f
C1353 XThC.Tn[0] XThC.Tn[1] 1.17084f
C1354 XA.XIR[9].XIC[7].icell.PUM Vbias 0.0031f
C1355 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.SM 0.00168f
C1356 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PUM 0.00465f
C1357 XA.XIR[4].XIC[4].icell.SM VPWR 0.00158f
C1358 XThR.Tn[12] XA.XIR[13].XIC[9].icell.SM 0.00121f
C1359 XA.XIR[10].XIC[1].icell.Ien Iout 0.06417f
C1360 XA.XIR[7].XIC[1].icell.PDM Iout 0.00117f
C1361 XThR.Tn[9] XA.XIR[10].XIC[1].icell.Ien 0.00338f
C1362 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.15202f
C1363 XThC.Tn[4] XThC.Tn[6] 0.00202f
C1364 XA.XIR[1].XIC_15.icell.SM Iout 0.0047f
C1365 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.03425f
C1366 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.15202f
C1367 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PUM 0.00429f
C1368 XA.XIR[6].XIC[8].icell.PDM Iout 0.00117f
C1369 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Ien 0.00232f
C1370 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PUM 0.00465f
C1371 a_n1049_7787# VPWR 0.72173f
C1372 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[12].icell.Ien 0.00214f
C1373 XA.XIR[3].XIC[8].icell.SM Vbias 0.00701f
C1374 XA.XIR[5].XIC_15.icell.PDM Iout 0.00133f
C1375 XA.XIR[1].XIC[10].icell.PDM Vbias 0.04261f
C1376 XA.XIR[14].XIC[5].icell.PDM Iout 0.00117f
C1377 XA.XIR[14].XIC[11].icell.SM Iout 0.00388f
C1378 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.SM 0.00168f
C1379 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C1380 XA.XIR[6].XIC[13].icell.Ien Vbias 0.21098f
C1381 XA.XIR[9].XIC[9].icell.PDM VPWR 0.00799f
C1382 a_10915_9569# VPWR 0.00307f
C1383 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PUM 0.00465f
C1384 XA.XIR[10].XIC[14].icell.Ien Vbias 0.21098f
C1385 XA.XIR[0].XIC[1].icell.PDM VPWR 0.00774f
C1386 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.SM 0.0039f
C1387 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02762f
C1388 XA.XIR[13].XIC[9].icell.PDM Iout 0.00117f
C1389 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00584f
C1390 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C1391 XA.XIR[2].XIC[1].icell.SM Vbias 0.00701f
C1392 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.SM 0.00168f
C1393 XA.XIR[7].XIC[3].icell.PUM Vbias 0.0031f
C1394 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.SM 0.0039f
C1395 XA.XIR[4].XIC[10].icell.PDM Vbias 0.04261f
C1396 XA.XIR[5].XIC_dummy_right.icell.PUM Vbias 0.00223f
C1397 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C1398 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.SM 0.00168f
C1399 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.03425f
C1400 XA.XIR[9].XIC[7].icell.SM VPWR 0.00158f
C1401 XThC.Tn[14] XThR.Tn[7] 0.28745f
C1402 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02762f
C1403 XA.XIR[1].XIC[3].icell.SM Vbias 0.00704f
C1404 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.SM 0.00168f
C1405 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00256f
C1406 XA.XIR[13].XIC_15.icell.PUM Vbias 0.0031f
C1407 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C1408 XThC.XTB5.A a_7331_10587# 0.01243f
C1409 XThC.Tn[0] XA.XIR[15].XIC_dummy_left.icell.Iout 0.00109f
C1410 XA.XIR[14].XIC[7].icell.Ien Vbias 0.21098f
C1411 XA.XIR[9].XIC[3].icell.SM Iout 0.00388f
C1412 XThR.XTB7.A data[5] 0.06538f
C1413 XThC.XTB7.B XThC.Tn[12] 0.00772f
C1414 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.SM 0.0039f
C1415 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C1416 XA.XIR[13].XIC[9].icell.Ien Vbias 0.21098f
C1417 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PUM 0.00465f
C1418 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04031f
C1419 XA.XIR[8].XIC[11].icell.SM Vbias 0.00701f
C1420 XThR.XTBN.Y XThR.Tn[5] 0.59912f
C1421 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00214f
C1422 a_n1319_5317# VPWR 0.00672f
C1423 XA.XIR[11].XIC[13].icell.Ien Iout 0.06417f
C1424 XA.XIR[3].XIC[10].icell.Ien VPWR 0.1903f
C1425 XThC.Tn[11] Vbias 2.46509f
C1426 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10] 0.00341f
C1427 XA.XIR[1].XIC[14].icell.PDM VPWR 0.00809f
C1428 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01577f
C1429 XA.XIR[10].XIC[14].icell.PDM VPWR 0.00809f
C1430 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C1431 XThR.XTBN.A a_n997_2667# 0.01679f
C1432 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14] 0.00341f
C1433 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.SM 0.00168f
C1434 XA.XIR[1].XIC[2].icell.PDM Iout 0.00117f
C1435 XThR.Tn[3] XThR.Tn[4] 0.06967f
C1436 XA.XIR[3].XIC[6].icell.Ien Iout 0.06417f
C1437 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02762f
C1438 XA.XIR[2].XIC[3].icell.Ien VPWR 0.1903f
C1439 XA.XIR[4].XIC[14].icell.PDM VPWR 0.00809f
C1440 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01493f
C1441 XA.XIR[7].XIC[3].icell.SM VPWR 0.00158f
C1442 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00214f
C1443 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04031f
C1444 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07214f
C1445 XA.XIR[5].XIC[12].icell.SM Iout 0.00388f
C1446 XA.XIR[4].XIC[2].icell.PDM Iout 0.00117f
C1447 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00256f
C1448 XA.XIR[1].XIC[5].icell.Ien VPWR 0.1903f
C1449 XA.XIR[14].XIC[9].icell.PUM VPWR 0.00937f
C1450 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.SM 0.00168f
C1451 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.SM 0.0039f
C1452 XA.XIR[10].XIC[11].icell.PUM Vbias 0.0031f
C1453 XA.XIR[4].XIC_15.icell.Ien Iout 0.0642f
C1454 XA.XIR[0].XIC[13].icell.SM Vbias 0.00716f
C1455 XA.XIR[3].XIC[10].icell.PDM Iout 0.00117f
C1456 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.SM 0.00168f
C1457 XA.XIR[8].XIC[12].icell.PDM Iout 0.00117f
C1458 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Ien 0.00584f
C1459 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.04036f
C1460 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Ien 0.00214f
C1461 XA.XIR[8].XIC[13].icell.Ien VPWR 0.1903f
C1462 XThR.XTB4.Y XThR.Tn[5] 0.00751f
C1463 XThR.Tn[6] XA.XIR[7].XIC[11].icell.SM 0.00121f
C1464 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.SM 0.0039f
C1465 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C1466 XThC.Tn[13] XThR.Tn[3] 0.2874f
C1467 XThR.Tn[12] XA.XIR[13].XIC[13].icell.Ien 0.00338f
C1468 XA.XIR[13].XIC[10].icell.SM Vbias 0.00701f
C1469 XA.XIR[8].XIC[9].icell.Ien Iout 0.06417f
C1470 XThR.Tn[8] XA.XIR[9].XIC[9].icell.Ien 0.00338f
C1471 XThC.XTB7.A XThC.XTBN.A 0.197f
C1472 XA.XIR[11].XIC[14].icell.SM Iout 0.00388f
C1473 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02762f
C1474 XThC.Tn[1] VPWR 5.91915f
C1475 XThC.XTB1.Y a_7651_9569# 0.06353f
C1476 XThR.Tn[0] XA.XIR[0].XIC[13].icell.PDM 0.00341f
C1477 XA.XIR[12].XIC[7].icell.SM Iout 0.00388f
C1478 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.SM 0.00168f
C1479 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12] 0.00341f
C1480 XA.XIR[1].XIC[0].icell.PUM VPWR 0.00937f
C1481 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.SM 0.0039f
C1482 XA.XIR[6].XIC_15.icell.SM Iout 0.0047f
C1483 XA.XIR[15].XIC[1].icell.PUM Vbias 0.0031f
C1484 XA.XIR[5].XIC[1].icell.Ien Vbias 0.21098f
C1485 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C1486 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02762f
C1487 XThR.Tn[1] XA.XIR[1].XIC[11].icell.PDM 0.00341f
C1488 XA.XIR[4].XIC[0].icell.PUM VPWR 0.00937f
C1489 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04031f
C1490 XThR.Tn[10] XA.XIR[11].XIC[1].icell.SM 0.00121f
C1491 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C1492 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02762f
C1493 XThR.XTBN.A XThR.Tn[11] 0.11968f
C1494 XThR.Tn[14] Vbias 3.74893f
C1495 XA.XIR[11].XIC[0].icell.PDM Vbias 0.04207f
C1496 XThC.Tn[9] XThR.Tn[5] 0.28739f
C1497 XThR.Tn[1] XA.XIR[2].XIC[2].icell.Ien 0.00338f
C1498 XA.XIR[13].XIC_dummy_left.icell.SM VPWR 0.00269f
C1499 XA.XIR[0].XIC_15.icell.Ien VPWR 0.2554f
C1500 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.03425f
C1501 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.SM 0.0039f
C1502 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04031f
C1503 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02834f
C1504 XA.XIR[14].XIC[9].icell.SM Iout 0.00388f
C1505 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[3].icell.Ien 0.00214f
C1506 XA.XIR[0].XIC[11].icell.Ien Iout 0.06389f
C1507 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.15202f
C1508 XA.XIR[10].XIC[4].icell.PDM Vbias 0.04261f
C1509 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.15202f
C1510 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.15202f
C1511 XA.XIR[10].XIC[12].icell.Ien Vbias 0.21098f
C1512 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02762f
C1513 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C1514 XThR.Tn[2] XA.XIR[2].XIC[8].icell.PDM 0.00341f
C1515 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C1516 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00584f
C1517 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C1518 XA.XIR[6].XIC[0].icell.Ien VPWR 0.1903f
C1519 XThR.Tn[13] XA.XIR[14].XIC[6].icell.Ien 0.00338f
C1520 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04031f
C1521 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PUM 0.00465f
C1522 XThR.XTB5.A XThR.XTB7.B 0.30355f
C1523 XThC.Tn[8] data[0] 0.01643f
C1524 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C1525 data[1] Vbias 0.00255f
C1526 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.SM 0.0039f
C1527 a_n1319_6405# VPWR 0.00676f
C1528 XA.XIR[6].XIC[3].icell.SM Vbias 0.00701f
C1529 XA.XIR[13].XIC[13].icell.PUM Vbias 0.0031f
C1530 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00584f
C1531 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.25759f
C1532 XThR.Tn[12] XA.XIR[13].XIC[14].icell.SM 0.00121f
C1533 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02762f
C1534 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.15202f
C1535 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.SM 0.00168f
C1536 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[9].icell.Ien 0.00214f
C1537 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.Ien 0.00584f
C1538 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.03425f
C1539 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PUM 0.00465f
C1540 a_6243_9615# XThC.Tn[6] 0.26142f
C1541 XA.XIR[15].XIC[6].icell.PUM Vbias 0.0031f
C1542 XA.XIR[7].XIC[14].icell.Ien Iout 0.06417f
C1543 XThR.Tn[0] XA.XIR[1].XIC[9].icell.Ien 0.00338f
C1544 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.SM 0.00168f
C1545 XA.XIR[5].XIC[6].icell.Ien Vbias 0.21098f
C1546 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.SM 0.00168f
C1547 XA.XIR[11].XIC[4].icell.PDM VPWR 0.00799f
C1548 XA.XIR[11].XIC[11].icell.Ien Iout 0.06417f
C1549 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.SM 0.00168f
C1550 XA.XIR[4].XIC[9].icell.PUM Vbias 0.0031f
C1551 XA.XIR[4].XIC[0].icell.SM Iout 0.00388f
C1552 XThR.Tn[7] XA.XIR[8].XIC_15.icell.Ien 0.00117f
C1553 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.SM 0.0039f
C1554 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00584f
C1555 XA.XIR[10].XIC[8].icell.PDM VPWR 0.00799f
C1556 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00214f
C1557 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C1558 XA.XIR[13].XIC[1].icell.Ien Iout 0.06417f
C1559 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C1560 XThR.Tn[5] XA.XIR[6].XIC[11].icell.Ien 0.00338f
C1561 XA.XIR[8].XIC[3].icell.PUM Vbias 0.0031f
C1562 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C1563 XA.XIR[6].XIC[5].icell.Ien VPWR 0.1903f
C1564 XA.XIR[15].XIC_dummy_right.icell.Ien Vbias 0.00288f
C1565 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00214f
C1566 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00584f
C1567 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.SM 0.00168f
C1568 XA.XIR[15].XIC[6].icell.SM VPWR 0.00158f
C1569 XA.XIR[0].XIC[12].icell.PDM Vbias 0.04282f
C1570 XA.XIR[11].XIC[2].icell.SM Vbias 0.00701f
C1571 XA.XIR[5].XIC[8].icell.PUM VPWR 0.00937f
C1572 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02762f
C1573 XA.XIR[13].XIC[14].icell.Ien Vbias 0.21098f
C1574 XThR.XTB6.Y a_n997_2667# 0.00468f
C1575 XA.XIR[9].XIC[12].icell.PUM Vbias 0.0031f
C1576 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PUM 0.00465f
C1577 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02762f
C1578 XA.XIR[15].XIC[2].icell.SM Iout 0.00388f
C1579 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00214f
C1580 XThR.XTB7.B data[5] 0.00593f
C1581 XA.XIR[4].XIC[9].icell.SM VPWR 0.00158f
C1582 XA.XIR[10].XIC[4].icell.SM Vbias 0.00701f
C1583 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.03425f
C1584 XA.XIR[0].XIC[0].icell.SM VPWR 0.00158f
C1585 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02762f
C1586 XThR.Tn[12] XA.XIR[13].XIC[11].icell.Ien 0.00338f
C1587 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.03425f
C1588 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.SM 0.0039f
C1589 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02762f
C1590 XThC.XTB5.A XThC.XTBN.A 0.06305f
C1591 XA.XIR[4].XIC[5].icell.SM Iout 0.00388f
C1592 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.15202f
C1593 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C1594 XA.XIR[2].XIC[0].icell.PDM VPWR 0.00799f
C1595 XA.XIR[0].XIC[5].icell.PUM Vbias 0.0031f
C1596 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC[0].icell.Ien 0.00214f
C1597 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02762f
C1598 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00584f
C1599 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C1600 XA.XIR[8].XIC[3].icell.SM VPWR 0.00158f
C1601 XA.XIR[3].XIC[13].icell.SM Vbias 0.00701f
C1602 XA.XIR[10].XIC[13].icell.PDM VPWR 0.00799f
C1603 XThC.XTB7.A XThC.Tn[2] 0.12602f
C1604 XThR.Tn[13] XA.XIR[14].XIC[0].icell.SM 0.00127f
C1605 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Iout 0.00401f
C1606 XA.XIR[12].XIC[3].icell.PUM VPWR 0.00937f
C1607 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00584f
C1608 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C1609 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.Ien 0.00584f
C1610 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.SM 0.00168f
C1611 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.SM 0.00168f
C1612 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C1613 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.03425f
C1614 XA.XIR[14].XIC[13].icell.Ien Iout 0.06417f
C1615 XA.XIR[11].XIC[4].icell.Ien VPWR 0.1903f
C1616 XA.XIR[2].XIC[6].icell.SM Vbias 0.00701f
C1617 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04037f
C1618 XA.XIR[7].XIC[8].icell.PUM Vbias 0.0031f
C1619 XA.XIR[9].XIC[12].icell.PDM Iout 0.00117f
C1620 XA.XIR[13].XIC[14].icell.PDM VPWR 0.00809f
C1621 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02762f
C1622 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9] 0.00341f
C1623 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.SM 0.0039f
C1624 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.SM 0.0039f
C1625 XA.XIR[9].XIC[12].icell.SM VPWR 0.00158f
C1626 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00214f
C1627 XA.XIR[1].XIC[8].icell.SM Vbias 0.00704f
C1628 XA.XIR[10].XIC[6].icell.Ien VPWR 0.1903f
C1629 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11] 0.00341f
C1630 XA.XIR[1].XIC[1].icell.Ien Iout 0.06417f
C1631 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.15202f
C1632 XThC.Tn[11] XThR.Tn[6] 0.28739f
C1633 XA.XIR[10].XIC[10].icell.Ien Vbias 0.21098f
C1634 XA.XIR[9].XIC[8].icell.SM Iout 0.00388f
C1635 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00214f
C1636 XA.XIR[10].XIC[2].icell.Ien Iout 0.06417f
C1637 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C1638 XThR.Tn[9] XA.XIR[10].XIC[2].icell.Ien 0.00338f
C1639 XA.XIR[0].XIC[5].icell.SM VPWR 0.00158f
C1640 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00584f
C1641 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C1642 XThR.Tn[7] XA.XIR[8].XIC[0].icell.SM 0.00121f
C1643 XA.XIR[3].XIC_15.icell.Ien VPWR 0.25566f
C1644 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00584f
C1645 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C1646 XA.XIR[0].XIC[1].icell.SM Iout 0.00367f
C1647 XA.XIR[13].XIC[11].icell.PUM Vbias 0.0031f
C1648 XThC.Tn[13] XThR.Tn[11] 0.2874f
C1649 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PUM 0.00465f
C1650 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C1651 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00584f
C1652 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12] 0.00341f
C1653 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39036f
C1654 XA.XIR[3].XIC[11].icell.Ien Iout 0.06417f
C1655 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8] 0.00341f
C1656 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[8].icell.Ien 0.00214f
C1657 XA.XIR[2].XIC[8].icell.Ien VPWR 0.1903f
C1658 XThC.Tn[3] XThR.Tn[7] 0.28739f
C1659 XA.XIR[7].XIC[8].icell.SM VPWR 0.00158f
C1660 XThC.XTB7.B XThC.Tn[1] 0.0014f
C1661 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.3891f
C1662 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C1663 XA.XIR[2].XIC[4].icell.Ien Iout 0.06417f
C1664 XA.XIR[1].XIC[10].icell.Ien VPWR 0.1903f
C1665 XA.XIR[14].XIC[14].icell.SM Iout 0.00388f
C1666 XA.XIR[7].XIC[4].icell.SM Iout 0.00388f
C1667 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04031f
C1668 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.15202f
C1669 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[5].icell.Ien 0.00214f
C1670 XA.XIR[1].XIC[6].icell.Ien Iout 0.06417f
C1671 XThC.Tn[0] Vbias 1.72566f
C1672 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C1673 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C1674 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02762f
C1675 XA.XIR[6].XIC[3].icell.PDM Vbias 0.04261f
C1676 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PUM 0.00465f
C1677 XThR.Tn[7] XA.XIR[8].XIC[5].icell.SM 0.00121f
C1678 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C1679 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00214f
C1680 XThC.XTB3.Y a_5949_9615# 0.009f
C1681 XA.XIR[14].XIC[0].icell.PDM Vbias 0.04207f
C1682 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02809f
C1683 XA.XIR[5].XIC[10].icell.PDM Vbias 0.04261f
C1684 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.03425f
C1685 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.SM 0.0039f
C1686 XThR.XTB5.A XThR.XTBN.Y 0.00282f
C1687 XThR.Tn[5] XA.XIR[6].XIC[1].icell.SM 0.00121f
C1688 XA.XIR[6].XIC_dummy_left.icell.SM VPWR 0.00269f
C1689 XA.XIR[8].XIC[14].icell.Ien Iout 0.06417f
C1690 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PUM 0.00465f
C1691 XThR.Tn[8] XA.XIR[9].XIC[14].icell.Ien 0.00338f
C1692 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.03425f
C1693 XThR.Tn[11] XA.XIR[12].XIC[3].icell.Ien 0.00338f
C1694 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02762f
C1695 XA.XIR[13].XIC[4].icell.PDM Vbias 0.04261f
C1696 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1697 XA.XIR[13].XIC[12].icell.Ien Vbias 0.21098f
C1698 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.15202f
C1699 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C1700 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04031f
C1701 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00214f
C1702 XThR.Tn[4] XA.XIR[4].XIC[10].icell.PDM 0.00341f
C1703 XA.XIR[12].XIC[9].icell.PDM Vbias 0.04261f
C1704 XThR.XTB7.B XThR.Tn[9] 0.0565f
C1705 XA.XIR[7].XIC[0].icell.PDM VPWR 0.00799f
C1706 XThR.Tn[10] XA.XIR[11].XIC[6].icell.SM 0.00121f
C1707 XA.XIR[10].XIC[0].icell.SM VPWR 0.00158f
C1708 XThR.Tn[3] XA.XIR[3].XIC[11].icell.PDM 0.00341f
C1709 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00584f
C1710 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C1711 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C1712 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.SM 0.0039f
C1713 XA.XIR[9].XIC[2].icell.Ien Vbias 0.21098f
C1714 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02762f
C1715 XThR.Tn[1] XA.XIR[2].XIC[7].icell.Ien 0.00338f
C1716 XA.XIR[6].XIC[7].icell.PDM VPWR 0.00799f
C1717 XThC.Tn[2] XThR.Tn[3] 0.28739f
C1718 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.SM 0.00168f
C1719 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.15202f
C1720 XA.XIR[0].XIC_dummy_right.icell.SM VPWR 0.00123f
C1721 XA.XIR[14].XIC[4].icell.PDM VPWR 0.00799f
C1722 XThC.XTBN.Y XThC.Tn[14] 0.50214f
C1723 XA.XIR[5].XIC[14].icell.PDM VPWR 0.00809f
C1724 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.15202f
C1725 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.03425f
C1726 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.03425f
C1727 XThC.Tn[11] XThR.Tn[4] 0.28739f
C1728 XA.XIR[14].XIC[11].icell.Ien Iout 0.06417f
C1729 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.SM 0.0039f
C1730 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C1731 XA.XIR[3].XIC[5].icell.PUM Vbias 0.0031f
C1732 XA.XIR[13].XIC[8].icell.PDM VPWR 0.00799f
C1733 XA.XIR[5].XIC[2].icell.PDM Iout 0.00117f
C1734 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C1735 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C1736 XA.XIR[6].XIC[8].icell.SM Vbias 0.00701f
C1737 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.03023f
C1738 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PUM 0.00429f
C1739 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00584f
C1740 XThC.XTB7.Y a_10051_9569# 0.013f
C1741 XA.XIR[6].XIC[1].icell.Ien Iout 0.06417f
C1742 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.SM 0.00168f
C1743 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.15202f
C1744 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.SM 0.00168f
C1745 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PUM 0.00465f
C1746 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C1747 XThR.Tn[0] XA.XIR[1].XIC[14].icell.Ien 0.00338f
C1748 XA.XIR[5].XIC[11].icell.Ien Vbias 0.21098f
C1749 XThC.Tn[5] XThR.Tn[0] 0.28744f
C1750 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.15202f
C1751 XThC.Tn[7] XThR.Tn[5] 0.28739f
C1752 XA.XIR[12].XIC[1].icell.PDM Iout 0.00117f
C1753 XA.XIR[9].XIC[4].icell.PUM VPWR 0.00937f
C1754 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PUM 0.00465f
C1755 XThR.Tn[2] Iout 1.16236f
C1756 XA.XIR[3].XIC[5].icell.PDM Vbias 0.04261f
C1757 XA.XIR[4].XIC[14].icell.PUM Vbias 0.0031f
C1758 XA.XIR[14].XIC[2].icell.SM Vbias 0.00701f
C1759 XA.XIR[8].XIC[7].icell.PDM Vbias 0.04261f
C1760 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.SM 0.00168f
C1761 XA.XIR[11].XIC[7].icell.PDM Iout 0.00117f
C1762 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1763 XThC.Tn[11] XThC.Tn[13] 0.00226f
C1764 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.SM 0.00168f
C1765 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C1766 XA.XIR[11].XIC[12].icell.SM VPWR 0.00158f
C1767 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.SM 0.0039f
C1768 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02762f
C1769 XA.XIR[2].XIC[11].icell.PDM Vbias 0.04261f
C1770 XA.XIR[13].XIC[4].icell.SM Vbias 0.00701f
C1771 XA.XIR[8].XIC[8].icell.PUM Vbias 0.0031f
C1772 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00584f
C1773 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.SM 0.0039f
C1774 XA.XIR[10].XIC[12].icell.PDM VPWR 0.00799f
C1775 XA.XIR[3].XIC[5].icell.SM VPWR 0.00158f
C1776 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02762f
C1777 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C1778 XA.XIR[1].XIC[1].icell.PDM VPWR 0.00799f
C1779 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.03425f
C1780 XA.XIR[6].XIC[10].icell.Ien VPWR 0.1903f
C1781 XA.XIR[12].XIC[6].icell.Ien Vbias 0.21098f
C1782 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.15202f
C1783 XA.XIR[3].XIC[1].icell.SM Iout 0.00388f
C1784 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PDM 0.0059f
C1785 XA.XIR[10].XIC_15.icell.Ien Vbias 0.21234f
C1786 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PUM 0.00465f
C1787 XA.XIR[5].XIC[13].icell.PUM VPWR 0.00937f
C1788 VPWR Vbias 0.2165p
C1789 XA.XIR[11].XIC[7].icell.SM Vbias 0.00701f
C1790 XThR.Tn[4] XA.XIR[5].XIC[1].icell.Ien 0.00338f
C1791 XA.XIR[13].XIC[13].icell.PDM VPWR 0.00799f
C1792 XA.XIR[4].XIC[1].icell.PDM VPWR 0.00799f
C1793 XA.XIR[6].XIC[6].icell.Ien Iout 0.06417f
C1794 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7] 0.00341f
C1795 XThR.XTBN.Y XA.XIR[14].XIC_dummy_left.icell.Iout 0.00116f
C1796 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.SM 0.0039f
C1797 XA.XIR[15].XIC[7].icell.SM Iout 0.00388f
C1798 XA.XIR[3].XIC[9].icell.PDM VPWR 0.00799f
C1799 XA.XIR[4].XIC[14].icell.SM VPWR 0.00207f
C1800 XThR.Tn[3] XA.XIR[4].XIC[1].icell.Ien 0.00338f
C1801 XA.XIR[14].XIC[4].icell.Ien VPWR 0.19084f
C1802 XA.XIR[8].XIC[11].icell.PDM VPWR 0.00799f
C1803 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C1804 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13] 0.00341f
C1805 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00584f
C1806 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PUM 0.00465f
C1807 XA.XIR[4].XIC[10].icell.SM Iout 0.00388f
C1808 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07214f
C1809 XThC.XTBN.A a_8739_9569# 0.01719f
C1810 XA.XIR[0].XIC[10].icell.PUM Vbias 0.0031f
C1811 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C1812 XA.XIR[13].XIC[6].icell.Ien VPWR 0.1903f
C1813 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.04036f
C1814 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.0353f
C1815 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04031f
C1816 XA.XIR[8].XIC[8].icell.SM VPWR 0.00158f
C1817 XA.XIR[13].XIC[10].icell.Ien Vbias 0.21098f
C1818 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C1819 XA.XIR[2].XIC[3].icell.PDM Iout 0.00117f
C1820 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01577f
C1821 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00584f
C1822 XA.XIR[13].XIC[2].icell.Ien Iout 0.06417f
C1823 XA.XIR[12].XIC[8].icell.PUM VPWR 0.00937f
C1824 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1825 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12] 0.00341f
C1826 XA.XIR[8].XIC[4].icell.SM Iout 0.00388f
C1827 XThC.Tn[4] XThR.Tn[2] 0.28739f
C1828 XThR.Tn[8] XA.XIR[9].XIC[4].icell.SM 0.00121f
C1829 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C1830 XThR.XTB6.Y XThR.Tn[14] 0.00128f
C1831 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00584f
C1832 XThR.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.00353f
C1833 XA.XIR[2].XIC[11].icell.SM Vbias 0.00701f
C1834 XA.XIR[11].XIC[9].icell.Ien VPWR 0.1903f
C1835 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.SM 0.00168f
C1836 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.SM 0.0039f
C1837 XA.XIR[7].XIC[13].icell.PUM Vbias 0.0031f
C1838 XThR.Tn[4] XA.XIR[5].XIC[6].icell.Ien 0.00338f
C1839 XThC.Tn[13] XThR.Tn[14] 0.2874f
C1840 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1841 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.SM 0.00168f
C1842 XA.XIR[11].XIC[5].icell.Ien Iout 0.06417f
C1843 XA.XIR[1].XIC[13].icell.SM Vbias 0.00704f
C1844 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC[0].icell.Ien 0.00214f
C1845 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C1846 XThR.Tn[3] XA.XIR[4].XIC[6].icell.Ien 0.00338f
C1847 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C1848 XA.XIR[9].XIC[13].icell.SM Iout 0.00388f
C1849 XA.XIR[10].XIC[7].icell.Ien Iout 0.06417f
C1850 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C1851 XThR.Tn[9] XA.XIR[10].XIC[7].icell.Ien 0.00338f
C1852 a_7875_9569# XThC.Tn[9] 0.19329f
C1853 XA.XIR[0].XIC[10].icell.SM VPWR 0.00158f
C1854 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.SM 0.00168f
C1855 XThC.XTB6.A XThC.Tn[5] 0.00363f
C1856 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5] 0.00341f
C1857 XA.XIR[3].XIC[2].icell.PUM Vbias 0.0031f
C1858 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.SM 0.0039f
C1859 XThC.XTB2.Y XThC.Tn[9] 0.292f
C1860 XA.XIR[0].XIC[6].icell.SM Iout 0.00367f
C1861 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C1862 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.04036f
C1863 XA.XIR[2].XIC[0].icell.PUM VPWR 0.00937f
C1864 XThR.XTB3.Y XThR.Tn[6] 0.00298f
C1865 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C1866 XA.XIR[12].XIC[0].icell.SM Vbias 0.00675f
C1867 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PUM 0.00465f
C1868 XA.XIR[3].XIC_dummy_right.icell.SM VPWR 0.00123f
C1869 XThR.Tn[13] XA.XIR[14].XIC[1].icell.SM 0.00121f
C1870 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04031f
C1871 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8] 0.00341f
C1872 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C1873 XA.XIR[2].XIC[13].icell.Ien VPWR 0.1903f
C1874 XA.XIR[7].XIC[13].icell.SM VPWR 0.00158f
C1875 XA.XIR[11].XIC_15.icell.SM Iout 0.0047f
C1876 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PUM 0.00465f
C1877 XThR.XTB1.Y XThR.Tn[1] 0.0099f
C1878 XThR.XTBN.Y XThR.Tn[9] 0.48048f
C1879 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02762f
C1880 XThC.Tn[0] XThR.Tn[6] 0.28741f
C1881 XA.XIR[1].XIC[1].icell.PUM VPWR 0.00937f
C1882 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.SM 0.00168f
C1883 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6] 0.00341f
C1884 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1885 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PUM 0.00465f
C1886 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C1887 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.SM 0.0039f
C1888 XA.XIR[2].XIC[9].icell.Ien Iout 0.06417f
C1889 XThR.Tn[0] XA.XIR[1].XIC[4].icell.SM 0.00121f
C1890 XA.XIR[7].XIC[9].icell.SM Iout 0.00388f
C1891 XA.XIR[1].XIC_15.icell.Ien VPWR 0.25566f
C1892 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.15202f
C1893 XA.XIR[7].XIC[11].icell.PDM Vbias 0.04261f
C1894 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.15202f
C1895 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C1896 XThC.XTBN.A XThC.Tn[11] 0.12129f
C1897 XA.XIR[5].XIC[1].icell.SM Vbias 0.00701f
C1898 XA.XIR[11].XIC[10].icell.SM VPWR 0.00158f
C1899 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PUM 0.00465f
C1900 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02774f
C1901 XThR.XTB5.Y a_n1049_5317# 0.00907f
C1902 XA.XIR[4].XIC[1].icell.PUM VPWR 0.00937f
C1903 XThR.Tn[12] XA.XIR[13].XIC[5].icell.Ien 0.00338f
C1904 XA.XIR[1].XIC[11].icell.Ien Iout 0.06417f
C1905 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.SM 0.00168f
C1906 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C1907 XA.XIR[4].XIC[4].icell.Ien Vbias 0.21098f
C1908 XA.XIR[15].XIC[9].icell.PDM Vbias 0.04261f
C1909 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Ien 0.00584f
C1910 XThC.Tn[2] XThR.Tn[11] 0.28739f
C1911 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PUM 0.00465f
C1912 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C1913 XA.XIR[13].XIC[0].icell.SM VPWR 0.00158f
C1914 XThR.Tn[7] XA.XIR[8].XIC[10].icell.SM 0.00121f
C1915 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C1916 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02762f
C1917 XThC.XTBN.Y a_4067_9615# 0.08456f
C1918 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11] 0.00341f
C1919 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C1920 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.SM 0.0039f
C1921 XThR.Tn[5] XA.XIR[6].XIC[6].icell.SM 0.00121f
C1922 XThR.Tn[11] XA.XIR[12].XIC[8].icell.Ien 0.00338f
C1923 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PUM 0.00465f
C1924 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C1925 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[0].icell.SM 0.0039f
C1926 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Iout 0.00347f
C1927 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.SM 0.0039f
C1928 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.15202f
C1929 XA.XIR[9].XIC[7].icell.PDM Vbias 0.04261f
C1930 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C1931 a_9827_9569# Vbias 0.00417f
C1932 XA.XIR[15].XIC[3].icell.PUM VPWR 0.00937f
C1933 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07214f
C1934 XA.XIR[5].XIC[3].icell.Ien VPWR 0.1903f
C1935 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C1936 XThC.XTB3.Y a_8739_9569# 0.07285f
C1937 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C1938 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02762f
C1939 XA.XIR[9].XIC[7].icell.Ien Vbias 0.21098f
C1940 XThC.XTB6.Y XThC.Tn[7] 0.01462f
C1941 XThR.Tn[1] XA.XIR[2].XIC[12].icell.Ien 0.00338f
C1942 XThR.Tn[10] Iout 1.16231f
C1943 XA.XIR[4].XIC[6].icell.PUM VPWR 0.00937f
C1944 XA.XIR[7].XIC[3].icell.PDM Iout 0.00117f
C1945 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.SM 0.0039f
C1946 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.SM 0.0039f
C1947 XThR.Tn[9] XThR.Tn[10] 0.07779f
C1948 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1949 XA.XIR[11].XIC[13].icell.PUM VPWR 0.00937f
C1950 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[8].icell.Ien 0.00214f
C1951 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.15202f
C1952 XA.XIR[15].XIC[1].icell.PDM Iout 0.00117f
C1953 XA.XIR[6].XIC[10].icell.PDM Iout 0.00117f
C1954 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.03535f
C1955 XThC.Tn[5] XThR.Tn[1] 0.2874f
C1956 XA.XIR[10].XIC[11].icell.PDM VPWR 0.00799f
C1957 XThR.XTB5.Y data[7] 0.00931f
C1958 XThC.Tn[9] Iout 0.83793f
C1959 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00584f
C1960 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.SM 0.00168f
C1961 XThC.Tn[9] XThR.Tn[9] 0.28739f
C1962 XA.XIR[14].XIC[7].icell.PDM Iout 0.00117f
C1963 XA.XIR[3].XIC[10].icell.PUM Vbias 0.0031f
C1964 XA.XIR[14].XIC[12].icell.SM VPWR 0.00158f
C1965 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00584f
C1966 XA.XIR[1].XIC[12].icell.PDM Vbias 0.04261f
C1967 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00256f
C1968 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C1969 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00584f
C1970 XA.XIR[6].XIC[13].icell.SM Vbias 0.00701f
C1971 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.03425f
C1972 XThC.Tn[5] XThR.Tn[12] 0.28739f
C1973 XA.XIR[9].XIC[11].icell.PDM VPWR 0.00799f
C1974 XThC.Tn[14] XThR.Tn[8] 0.28745f
C1975 XA.XIR[13].XIC[12].icell.PDM VPWR 0.00799f
C1976 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PUM 0.00465f
C1977 XThR.XTB3.Y XThR.Tn[4] 0.00382f
C1978 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.SM 0.00168f
C1979 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.Ien 0.00584f
C1980 XA.XIR[0].XIC[3].icell.PDM VPWR 0.00774f
C1981 XA.XIR[4].XIC[12].icell.PDM Vbias 0.04261f
C1982 XA.XIR[2].XIC[3].icell.PUM Vbias 0.0031f
C1983 XA.XIR[7].XIC[3].icell.Ien Vbias 0.21098f
C1984 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C1985 XThC.XTB6.Y a_5949_10571# 0.01283f
C1986 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00584f
C1987 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C1988 XA.XIR[1].XIC[0].icell.SM VPWR 0.00158f
C1989 XThR.XTB3.Y a_n1049_7493# 0.23056f
C1990 XA.XIR[9].XIC[9].icell.PUM VPWR 0.00937f
C1991 XThC.XTB7.B Vbias 0.09241f
C1992 XThC.Tn[0] XThR.Tn[4] 0.28743f
C1993 XA.XIR[13].XIC_15.icell.Ien Vbias 0.21234f
C1994 XA.XIR[1].XIC[5].icell.PUM Vbias 0.0031f
C1995 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C1996 XThC.XTBN.Y XThC.Tn[3] 0.62681f
C1997 XA.XIR[10].XIC[1].icell.SM VPWR 0.00158f
C1998 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C1999 XA.XIR[14].XIC[7].icell.SM Vbias 0.00701f
C2000 XThR.XTBN.A VPWR 0.90694f
C2001 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C2002 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C2003 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02762f
C2004 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02762f
C2005 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.15202f
C2006 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.SM 0.0039f
C2007 XThC.XTBN.A data[1] 0.01444f
C2008 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.PDM 0.0059f
C2009 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00584f
C2010 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C2011 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00214f
C2012 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.03425f
C2013 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.SM 0.00168f
C2014 XThR.XTB5.Y a_n1049_6405# 0.24821f
C2015 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04031f
C2016 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.SM 0.00168f
C2017 XA.XIR[8].XIC[13].icell.PUM Vbias 0.0031f
C2018 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04038f
C2019 XA.XIR[11].XIC[14].icell.Ien VPWR 0.19036f
C2020 XThR.Tn[6] VPWR 6.58002f
C2021 XA.XIR[3].XIC[10].icell.SM VPWR 0.00158f
C2022 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2023 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C2024 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10] 0.00341f
C2025 XA.XIR[6].XIC_15.icell.Ien VPWR 0.25566f
C2026 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C2027 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01721f
C2028 XThC.XTB4.Y XThC.Tn[7] 0.01797f
C2029 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02762f
C2030 XThC.Tn[4] XThR.Tn[10] 0.28739f
C2031 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14] 0.00341f
C2032 XA.XIR[3].XIC[6].icell.SM Iout 0.00388f
C2033 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02762f
C2034 XA.XIR[1].XIC[4].icell.PDM Iout 0.00117f
C2035 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C2036 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.15202f
C2037 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[5].icell.SM 0.0039f
C2038 XA.XIR[2].XIC[3].icell.SM VPWR 0.00158f
C2039 XA.XIR[6].XIC[11].icell.Ien Iout 0.06417f
C2040 XA.XIR[7].XIC[5].icell.PUM VPWR 0.00937f
C2041 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01577f
C2042 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2043 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.03023f
C2044 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C2045 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PUM 0.00465f
C2046 XA.XIR[4].XIC[4].icell.PDM Iout 0.00117f
C2047 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.SM 0.0039f
C2048 XA.XIR[1].XIC[5].icell.SM VPWR 0.00158f
C2049 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00214f
C2050 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.SM 0.0039f
C2051 Vbias bias[0] 0.21039f
C2052 bias[1] bias[2] 0.16429f
C2053 XA.XIR[14].XIC[9].icell.Ien VPWR 0.19084f
C2054 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C2055 XA.XIR[1].XIC[1].icell.SM Iout 0.00388f
C2056 XA.XIR[3].XIC[12].icell.PDM Iout 0.00117f
C2057 a_4861_9615# XThC.Tn[3] 0.27012f
C2058 XA.XIR[0].XIC_15.icell.PUM Vbias 0.0031f
C2059 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C2060 XA.XIR[14].XIC[5].icell.Ien Iout 0.06417f
C2061 XA.XIR[8].XIC[14].icell.PDM Iout 0.00117f
C2062 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PDM 0.00172f
C2063 XA.XIR[8].XIC[13].icell.SM VPWR 0.00158f
C2064 XThC.Tn[0] XA.XIR[10].XIC_dummy_left.icell.Iout 0.00109f
C2065 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.389f
C2066 XA.XIR[13].XIC[7].icell.Ien Iout 0.06417f
C2067 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.15202f
C2068 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2069 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.SM 0.00168f
C2070 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.Ien 0.00256f
C2071 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C2072 XA.XIR[8].XIC[9].icell.SM Iout 0.00388f
C2073 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C2074 XThR.Tn[8] XA.XIR[9].XIC[9].icell.SM 0.00121f
C2075 XThR.Tn[0] XA.XIR[0].XIC_15.icell.PDM 0.00341f
C2076 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C2077 XThR.Tn[2] XA.XIR[3].XIC[4].icell.Ien 0.00338f
C2078 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2079 XThR.Tn[4] XA.XIR[5].XIC[11].icell.Ien 0.00338f
C2080 XA.XIR[15].XIC[1].icell.Ien Vbias 0.17899f
C2081 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.SM 0.0039f
C2082 XThR.Tn[1] XA.XIR[1].XIC[13].icell.PDM 0.00341f
C2083 XA.XIR[11].XIC[11].icell.PUM VPWR 0.00937f
C2084 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04031f
C2085 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C2086 XA.XIR[14].XIC_15.icell.SM Iout 0.0047f
C2087 XThR.Tn[3] XA.XIR[4].XIC[11].icell.Ien 0.00338f
C2088 a_7331_10587# VPWR 0.0063f
C2089 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00584f
C2090 XThR.Tn[1] XA.XIR[2].XIC[2].icell.SM 0.00121f
C2091 XA.XIR[11].XIC[2].icell.PDM Vbias 0.04261f
C2092 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02762f
C2093 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04031f
C2094 XA.XIR[14].XIC[10].icell.SM VPWR 0.00158f
C2095 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C2096 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11] 0.00341f
C2097 XA.XIR[10].XIC[6].icell.PDM Vbias 0.04261f
C2098 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00584f
C2099 XA.XIR[0].XIC[11].icell.SM Iout 0.00367f
C2100 XA.XIR[5].XIC[1].icell.PDM VPWR 0.00799f
C2101 XThR.Tn[2] XA.XIR[2].XIC[10].icell.PDM 0.00341f
C2102 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02762f
C2103 XThC.Tn[2] XThR.Tn[14] 0.28739f
C2104 XA.XIR[6].XIC[0].icell.SM VPWR 0.00158f
C2105 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.03425f
C2106 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04031f
C2107 XThR.Tn[13] XA.XIR[14].XIC[6].icell.SM 0.00121f
C2108 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.SM 0.00168f
C2109 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[13].icell.Ien 0.00214f
C2110 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00584f
C2111 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02762f
C2112 XA.XIR[6].XIC[5].icell.PUM Vbias 0.0031f
C2113 XThR.Tn[4] VPWR 6.61651f
C2114 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C2115 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.03425f
C2116 XA.XIR[2].XIC[14].icell.Ien Iout 0.06417f
C2117 XA.XIR[15].XIC[6].icell.Ien Vbias 0.17899f
C2118 XA.XIR[12].XIC[0].icell.PDM VPWR 0.00799f
C2119 XA.XIR[5].XIC[6].icell.SM Vbias 0.00701f
C2120 XThR.Tn[0] XA.XIR[1].XIC[9].icell.SM 0.00121f
C2121 XA.XIR[7].XIC[14].icell.SM Iout 0.00388f
C2122 a_n1049_7493# VPWR 0.72084f
C2123 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[10].icell.Ien 0.00214f
C2124 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C2125 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PUM 0.00465f
C2126 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C2127 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C2128 XA.XIR[11].XIC[6].icell.PDM VPWR 0.00799f
C2129 XA.XIR[1].XIC_dummy_right.icell.SM VPWR 0.00123f
C2130 XA.XIR[11].XIC[12].icell.Ien VPWR 0.1903f
C2131 XA.XIR[4].XIC[9].icell.Ien Vbias 0.21098f
C2132 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C2133 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00584f
C2134 XA.XIR[14].XIC[0].icell.Ien Iout 0.06411f
C2135 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C2136 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02762f
C2137 XA.XIR[0].XIC[0].icell.Ien Vbias 0.20991f
C2138 XA.XIR[10].XIC[10].icell.PDM VPWR 0.00799f
C2139 XThR.Tn[13] Iout 1.16236f
C2140 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.15202f
C2141 XThR.XTB6.Y VPWR 1.05512f
C2142 XThR.Tn[5] XA.XIR[6].XIC[11].icell.SM 0.00121f
C2143 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C2144 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PUM 0.00465f
C2145 XA.XIR[14].XIC[13].icell.PUM VPWR 0.00937f
C2146 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[14].icell.Ien 0.00214f
C2147 XA.XIR[8].XIC[3].icell.Ien Vbias 0.21098f
C2148 XThC.Tn[13] VPWR 6.87751f
C2149 XA.XIR[12].XIC[1].icell.SM Vbias 0.00701f
C2150 XA.XIR[6].XIC[5].icell.SM VPWR 0.00158f
C2151 XA.XIR[13].XIC[11].icell.PDM VPWR 0.00799f
C2152 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.15202f
C2153 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C2154 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C2155 XA.XIR[15].XIC[8].icell.PUM VPWR 0.00937f
C2156 XA.XIR[0].XIC[14].icell.PDM Vbias 0.04282f
C2157 XA.XIR[11].XIC[4].icell.PUM Vbias 0.0031f
C2158 XA.XIR[6].XIC[1].icell.SM Iout 0.00388f
C2159 XA.XIR[5].XIC[8].icell.Ien VPWR 0.1903f
C2160 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PUM 0.00102f
C2161 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11267f
C2162 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C2163 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.03425f
C2164 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C2165 XA.XIR[9].XIC[12].icell.Ien Vbias 0.21098f
C2166 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00584f
C2167 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.03425f
C2168 XA.XIR[5].XIC[4].icell.Ien Iout 0.06417f
C2169 XA.XIR[4].XIC[11].icell.PUM VPWR 0.00937f
C2170 XA.XIR[10].XIC[6].icell.PUM Vbias 0.0031f
C2171 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C2172 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00584f
C2173 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.SM 0.0039f
C2174 XA.XIR[0].XIC[2].icell.PUM VPWR 0.00877f
C2175 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C2176 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02762f
C2177 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C2178 XA.XIR[0].XIC[5].icell.Ien Vbias 0.2113f
C2179 XA.XIR[2].XIC[2].icell.PDM VPWR 0.00799f
C2180 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.PDM 0.00598f
C2181 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[5].icell.Ien 0.00214f
C2182 XA.XIR[13].XIC[1].icell.SM VPWR 0.00158f
C2183 XA.XIR[8].XIC[5].icell.PUM VPWR 0.00937f
C2184 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.SM 0.0039f
C2185 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02762f
C2186 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02762f
C2187 XThR.Tn[6] XA.XIR[7].XIC[3].icell.Ien 0.00338f
C2188 XA.XIR[3].XIC_15.icell.PUM Vbias 0.0031f
C2189 XThR.Tn[2] XA.XIR[3].XIC[1].icell.Ien 0.00338f
C2190 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C2191 XA.XIR[12].XIC[3].icell.Ien VPWR 0.1903f
C2192 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.SM 0.00168f
C2193 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PUM 0.00465f
C2194 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.SM 0.00168f
C2195 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00584f
C2196 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02812f
C2197 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1909f
C2198 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.SM 0.0039f
C2199 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C2200 XA.XIR[2].XIC[8].icell.PUM Vbias 0.0031f
C2201 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04031f
C2202 XA.XIR[11].XIC[4].icell.SM VPWR 0.00158f
C2203 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02762f
C2204 XA.XIR[10].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2205 XA.XIR[7].XIC[8].icell.Ien Vbias 0.21098f
C2206 XA.XIR[9].XIC[14].icell.PDM Iout 0.00117f
C2207 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02762f
C2208 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9] 0.00341f
C2209 XThR.Tn[4] XA.XIR[5].XIC[1].icell.SM 0.00121f
C2210 XThC.Tn[4] XThR.Tn[13] 0.28739f
C2211 XA.XIR[9].XIC[14].icell.PUM VPWR 0.00937f
C2212 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11] 0.00341f
C2213 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00584f
C2214 XA.XIR[1].XIC[10].icell.PUM Vbias 0.0031f
C2215 XA.XIR[10].XIC[6].icell.SM VPWR 0.00158f
C2216 XA.XIR[4].XIC_15.icell.SM VPWR 0.00275f
C2217 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.15202f
C2218 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.SM 0.0039f
C2219 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C2220 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.0353f
C2221 XThR.Tn[14] XA.XIR[15].XIC[3].icell.Ien 0.00338f
C2222 XThR.Tn[3] XA.XIR[4].XIC[1].icell.SM 0.00121f
C2223 XA.XIR[10].XIC[2].icell.SM Iout 0.00388f
C2224 XThC.XTB2.Y a_3773_9615# 0.2342f
C2225 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.SM 0.00168f
C2226 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00584f
C2227 XA.XIR[0].XIC[7].icell.PUM VPWR 0.00877f
C2228 XThR.Tn[9] XA.XIR[10].XIC[2].icell.SM 0.00121f
C2229 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Iout 0.00347f
C2230 XThC.Tn[7] Iout 0.84037f
C2231 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00584f
C2232 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C2233 XThC.Tn[7] XThR.Tn[9] 0.28739f
C2234 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.SM 0.0039f
C2235 XThC.Tn[3] XThR.Tn[8] 0.28739f
C2236 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PUM 0.00465f
C2237 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.04036f
C2238 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.03425f
C2239 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[3].icell.Ien 0.00214f
C2240 XThC.Tn[0] XA.XIR[13].XIC_dummy_left.icell.Iout 0.00109f
C2241 XA.XIR[3].XIC[11].icell.SM Iout 0.00388f
C2242 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C2243 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8] 0.00341f
C2244 XA.XIR[6].XIC_dummy_right.icell.SM VPWR 0.00123f
C2245 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.15202f
C2246 XA.XIR[7].XIC[10].icell.PUM VPWR 0.00937f
C2247 XA.XIR[2].XIC[8].icell.SM VPWR 0.00158f
C2248 a_n1049_8581# Vbias 0.00113f
C2249 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Ien 0.00584f
C2250 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C2251 XA.XIR[11].XIC[10].icell.Ien VPWR 0.1903f
C2252 XA.XIR[2].XIC[4].icell.SM Iout 0.00388f
C2253 XA.XIR[1].XIC[10].icell.SM VPWR 0.00158f
C2254 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04031f
C2255 XA.XIR[10].XIC[0].icell.Ien Vbias 0.20951f
C2256 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PUM 0.00465f
C2257 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00584f
C2258 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[13].icell.Ien 0.00214f
C2259 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PUM 0.00465f
C2260 XA.XIR[1].XIC[6].icell.SM Iout 0.00388f
C2261 XA.XIR[14].XIC[11].icell.PUM VPWR 0.00937f
C2262 XA.XIR[6].XIC[5].icell.PDM Vbias 0.04261f
C2263 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11] 0.00341f
C2264 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00584f
C2265 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.SM 0.00168f
C2266 VPWR data[3] 0.20846f
C2267 XThC.XTBN.A VPWR 0.88811f
C2268 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.15202f
C2269 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Ien 0.00232f
C2270 XA.XIR[5].XIC[12].icell.PDM Vbias 0.04261f
C2271 XA.XIR[14].XIC[2].icell.PDM Vbias 0.04261f
C2272 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00584f
C2273 XThC.Tn[5] XA.XIR[0].XIC[6].icell.Ien 0.0016f
C2274 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.15202f
C2275 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C2276 XThR.Tn[11] XA.XIR[12].XIC[3].icell.SM 0.00121f
C2277 XA.XIR[8].XIC[14].icell.SM Iout 0.00388f
C2278 a_9827_9569# XThC.Tn[13] 0.00173f
C2279 XA.XIR[2].XIC[1].icell.PUM VPWR 0.00937f
C2280 XThR.Tn[8] XA.XIR[9].XIC[14].icell.SM 0.00121f
C2281 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PUM 0.00465f
C2282 XThC.Tn[0] XThC.Tn[2] 0.1179f
C2283 XA.XIR[13].XIC[6].icell.PDM Vbias 0.04261f
C2284 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C2285 XThR.Tn[2] XA.XIR[3].XIC[9].icell.Ien 0.00338f
C2286 XA.XIR[11].XIC[0].icell.Ien VPWR 0.1903f
C2287 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.SM 0.00168f
C2288 XThC.Tn[5] XThC.Tn[6] 0.30991f
C2289 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04031f
C2290 XThR.Tn[4] XA.XIR[4].XIC[12].icell.PDM 0.00341f
C2291 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Ien 0.00584f
C2292 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2293 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02762f
C2294 XA.XIR[7].XIC[2].icell.PDM VPWR 0.00799f
C2295 XA.XIR[10].XIC[2].icell.PUM VPWR 0.00937f
C2296 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C2297 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.15202f
C2298 XThR.Tn[3] XA.XIR[3].XIC[13].icell.PDM 0.00341f
C2299 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14] 0.00341f
C2300 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2301 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C2302 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C2303 XA.XIR[9].XIC[2].icell.SM Vbias 0.00701f
C2304 XThR.Tn[1] XA.XIR[2].XIC[7].icell.SM 0.00121f
C2305 XA.XIR[6].XIC[9].icell.PDM VPWR 0.00799f
C2306 XA.XIR[15].XIC[0].icell.PDM VPWR 0.0114f
C2307 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C2308 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.SM 0.0039f
C2309 XThR.XTB6.A XThR.Tn[1] 0.00411f
C2310 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C2311 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2312 XA.XIR[14].XIC[6].icell.PDM VPWR 0.00799f
C2313 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C2314 XA.XIR[14].XIC[12].icell.Ien VPWR 0.19084f
C2315 XA.XIR[5].XIC[4].icell.PDM Iout 0.00117f
C2316 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.03425f
C2317 XA.XIR[3].XIC[5].icell.Ien Vbias 0.21098f
C2318 XA.XIR[13].XIC[10].icell.PDM VPWR 0.00799f
C2319 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C2320 XA.XIR[6].XIC[10].icell.PUM Vbias 0.0031f
C2321 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02762f
C2322 XThR.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.00338f
C2323 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.03574f
C2324 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.0353f
C2325 XThC.XTB7.Y XThC.Tn[8] 0.07806f
C2326 XThR.XTBN.Y XA.XIR[9].XIC_dummy_left.icell.Iout 0.00395f
C2327 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Ien 0.00595f
C2328 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C2329 XThC.XTB7.B XThC.Tn[13] 0.00276f
C2330 XThR.Tn[0] XA.XIR[1].XIC[14].icell.SM 0.00121f
C2331 XA.XIR[5].XIC[11].icell.SM Vbias 0.00701f
C2332 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.SM 0.00168f
C2333 XA.XIR[9].XIC[4].icell.Ien VPWR 0.1903f
C2334 XA.XIR[12].XIC[3].icell.PDM Iout 0.00117f
C2335 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.Ien 0.00584f
C2336 XThC.Tn[12] Vbias 2.48601f
C2337 XThR.Tn[0] XThR.Tn[1] 0.22353f
C2338 XA.XIR[3].XIC[7].icell.PDM Vbias 0.04261f
C2339 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.03425f
C2340 XA.XIR[4].XIC[14].icell.Ien Vbias 0.21098f
C2341 XA.XIR[14].XIC[4].icell.PUM Vbias 0.0031f
C2342 XA.XIR[8].XIC[9].icell.PDM Vbias 0.04261f
C2343 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PUM 0.00465f
C2344 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C2345 XA.XIR[11].XIC[9].icell.PDM Iout 0.00117f
C2346 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11153f
C2347 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.SM 0.00168f
C2348 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[4].icell.Ien 0.00214f
C2349 XA.XIR[2].XIC[13].icell.PDM Vbias 0.04261f
C2350 XA.XIR[13].XIC[6].icell.PUM Vbias 0.0031f
C2351 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.SM 0.0039f
C2352 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.15202f
C2353 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C2354 XA.XIR[8].XIC[8].icell.Ien Vbias 0.21098f
C2355 XA.XIR[3].XIC[7].icell.PUM VPWR 0.00937f
C2356 XA.XIR[1].XIC[3].icell.PDM VPWR 0.00799f
C2357 XA.XIR[6].XIC[10].icell.SM VPWR 0.00158f
C2358 XA.XIR[12].XIC[6].icell.SM Vbias 0.00701f
C2359 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02762f
C2360 XA.XIR[10].XIC_15.icell.PDM Vbias 0.04401f
C2361 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.03425f
C2362 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C2363 XA.XIR[5].XIC[13].icell.Ien VPWR 0.1903f
C2364 XA.XIR[11].XIC[9].icell.PUM Vbias 0.0031f
C2365 XA.XIR[6].XIC[6].icell.SM Iout 0.00388f
C2366 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7] 0.00341f
C2367 XA.XIR[4].XIC[3].icell.PDM VPWR 0.00799f
C2368 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[12].icell.Ien 0.00214f
C2369 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00584f
C2370 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C2371 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Iout 0.00347f
C2372 XA.XIR[0].XIC_dummy_left.icell.Ien Vbias 0.00487f
C2373 XThC.XTB3.Y VPWR 1.07065f
C2374 XA.XIR[5].XIC[9].icell.Ien Iout 0.06417f
C2375 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.SM 0.0039f
C2376 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2377 XThC.XTB1.Y XThC.Tn[0] 0.19116f
C2378 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02762f
C2379 XA.XIR[3].XIC[11].icell.PDM VPWR 0.00799f
C2380 XA.XIR[8].XIC[13].icell.PDM VPWR 0.00799f
C2381 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C2382 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13] 0.00341f
C2383 XA.XIR[14].XIC[4].icell.SM VPWR 0.00158f
C2384 XThC.Tn[14] XThR.Tn[3] 0.28745f
C2385 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PUM 0.00465f
C2386 XA.XIR[13].XIC_dummy_right.icell.Ien Vbias 0.00288f
C2387 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[13].icell.Ien 0.00214f
C2388 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.03425f
C2389 XThC.XTB7.A a_6243_10571# 0.0017f
C2390 XThC.Tn[2] VPWR 5.93664f
C2391 XA.XIR[8].XIC[1].icell.PDM Iout 0.00117f
C2392 XA.XIR[0].XIC[10].icell.Ien Vbias 0.2113f
C2393 XThC.XTBN.A a_9827_9569# 0.09118f
C2394 XA.XIR[13].XIC[6].icell.SM VPWR 0.00158f
C2395 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04031f
C2396 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04031f
C2397 XA.XIR[8].XIC[10].icell.PUM VPWR 0.00937f
C2398 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.PDM 0.00591f
C2399 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C2400 XA.XIR[2].XIC[5].icell.PDM Iout 0.00117f
C2401 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00256f
C2402 XThR.Tn[6] XA.XIR[7].XIC[8].icell.Ien 0.00338f
C2403 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07214f
C2404 XA.XIR[13].XIC[2].icell.SM Iout 0.00388f
C2405 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00584f
C2406 XA.XIR[11].XIC_15.icell.Ien VPWR 0.25566f
C2407 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00214f
C2408 XA.XIR[12].XIC[8].icell.Ien VPWR 0.1903f
C2409 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C2410 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2411 XThC.Tn[8] XThR.Tn[0] 0.28773f
C2412 XThC.Tn[10] XThR.Tn[5] 0.28739f
C2413 XThR.Tn[0] XA.XIR[0].XIC[2].icell.PDM 0.00341f
C2414 XA.XIR[12].XIC[4].icell.Ien Iout 0.06417f
C2415 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C2416 XA.XIR[2].XIC[13].icell.PUM Vbias 0.0031f
C2417 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C2418 XA.XIR[7].XIC[13].icell.Ien Vbias 0.21098f
C2419 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00214f
C2420 XThR.Tn[4] XA.XIR[5].XIC[6].icell.SM 0.00121f
C2421 XThR.Tn[1] XA.XIR[1].XIC[0].icell.PDM 0.00347f
C2422 XA.XIR[11].XIC[5].icell.SM Iout 0.00388f
C2423 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C2424 XA.XIR[1].XIC_15.icell.PUM Vbias 0.0031f
C2425 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C2426 XThR.Tn[3] XA.XIR[4].XIC[6].icell.SM 0.00121f
C2427 XThR.Tn[14] XA.XIR[15].XIC[8].icell.Ien 0.00338f
C2428 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.15202f
C2429 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.03425f
C2430 XA.XIR[14].XIC[10].icell.Ien VPWR 0.19084f
C2431 XA.XIR[10].XIC[7].icell.SM Iout 0.00388f
C2432 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C2433 XThC.XTB5.Y a_5155_9615# 0.24821f
C2434 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11] 0.00341f
C2435 XA.XIR[0].XIC[12].icell.PUM VPWR 0.00878f
C2436 XThR.Tn[9] XA.XIR[10].XIC[7].icell.SM 0.00121f
C2437 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C2438 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00214f
C2439 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5] 0.00341f
C2440 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PUM 0.00465f
C2441 XA.XIR[13].XIC[0].icell.Ien Vbias 0.20951f
C2442 XThC.XTB7.A a_4067_9615# 0.0127f
C2443 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PDM 0.00172f
C2444 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C2445 XThC.XTBN.A XThC.XTB7.B 0.35142f
C2446 XA.XIR[12].XIC[2].icell.PUM Vbias 0.0031f
C2447 XA.XIR[11].XIC_dummy_left.icell.SM VPWR 0.00269f
C2448 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04052f
C2449 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[10].icell.SM 0.0039f
C2450 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.03425f
C2451 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.15202f
C2452 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2453 XA.XIR[2].XIC[13].icell.SM VPWR 0.00158f
C2454 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01577f
C2455 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00584f
C2456 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PUM 0.00465f
C2457 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6] 0.00341f
C2458 XA.XIR[2].XIC[9].icell.SM Iout 0.00388f
C2459 XA.XIR[15].XIC[1].icell.SM Vbias 0.00701f
C2460 XA.XIR[7].XIC[13].icell.PDM Vbias 0.04261f
C2461 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14] 0.00341f
C2462 XA.XIR[5].XIC[3].icell.PUM Vbias 0.0031f
C2463 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.03425f
C2464 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.SM 0.00168f
C2465 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.SM 0.0039f
C2466 XThR.Tn[12] XA.XIR[13].XIC[5].icell.SM 0.00121f
C2467 XA.XIR[4].XIC[1].icell.Ien VPWR 0.1903f
C2468 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C2469 XA.XIR[1].XIC[11].icell.SM Iout 0.00388f
C2470 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C2471 XA.XIR[4].XIC[4].icell.SM Vbias 0.00701f
C2472 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.03425f
C2473 XA.XIR[13].XIC[2].icell.PUM VPWR 0.00937f
C2474 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.15202f
C2475 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00214f
C2476 XThC.XTBN.Y a_5155_9615# 0.07602f
C2477 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.15202f
C2478 XThR.Tn[11] XA.XIR[12].XIC[8].icell.SM 0.00121f
C2479 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[11].icell.Ien 0.00214f
C2480 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.SM 0.00168f
C2481 XThR.Tn[2] XA.XIR[3].XIC[14].icell.Ien 0.00338f
C2482 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.SM 0.0039f
C2483 XThC.XTB1.Y VPWR 1.1176f
C2484 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PUM 0.00176f
C2485 XA.XIR[9].XIC[9].icell.PDM Vbias 0.04261f
C2486 a_10915_9569# Vbias 0.00873f
C2487 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C2488 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02762f
C2489 XThR.Tn[7] Iout 1.16233f
C2490 XA.XIR[15].XIC[3].icell.Ien VPWR 0.32895f
C2491 XA.XIR[0].XIC[1].icell.PDM Vbias 0.04282f
C2492 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C2493 XA.XIR[5].XIC[3].icell.SM VPWR 0.00158f
C2494 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.SM 0.0039f
C2495 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.15202f
C2496 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02762f
C2497 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02762f
C2498 XA.XIR[7].XIC_15.icell.SM Iout 0.0047f
C2499 XThC.XTB7.A XThC.Tn[3] 0.03065f
C2500 XThR.Tn[1] XA.XIR[2].XIC[12].icell.SM 0.00121f
C2501 XA.XIR[9].XIC[7].icell.SM Vbias 0.00701f
C2502 XA.XIR[7].XIC[5].icell.PDM Iout 0.00117f
C2503 XA.XIR[4].XIC[6].icell.Ien VPWR 0.1903f
C2504 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.15235f
C2505 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01432f
C2506 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00214f
C2507 XA.XIR[15].XIC[3].icell.PDM Iout 0.00117f
C2508 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PUM 0.00465f
C2509 XA.XIR[4].XIC[2].icell.Ien Iout 0.06417f
C2510 XA.XIR[6].XIC[12].icell.PDM Iout 0.00117f
C2511 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C2512 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.SM 0.0039f
C2513 VPWR bias[2] 1.20331f
C2514 a_2979_9615# XThC.Tn[0] 0.28426f
C2515 XA.XIR[3].XIC[10].icell.Ien Vbias 0.21098f
C2516 XA.XIR[14].XIC[9].icell.PDM Iout 0.00117f
C2517 XA.XIR[1].XIC[14].icell.PDM Vbias 0.04261f
C2518 XA.XIR[6].XIC_15.icell.PUM Vbias 0.0031f
C2519 XA.XIR[9].XIC[13].icell.PDM VPWR 0.00799f
C2520 XA.XIR[10].XIC[14].icell.PDM Vbias 0.04261f
C2521 XThC.Tn[12] XThR.Tn[6] 0.28739f
C2522 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.SM 0.0039f
C2523 XA.XIR[0].XIC[5].icell.PDM VPWR 0.00908f
C2524 XA.XIR[7].XIC[0].icell.Ien VPWR 0.1903f
C2525 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.SM 0.0039f
C2526 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C2527 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C2528 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.03425f
C2529 XA.XIR[7].XIC[3].icell.SM Vbias 0.00701f
C2530 XA.XIR[2].XIC[3].icell.Ien Vbias 0.21098f
C2531 XA.XIR[4].XIC[14].icell.PDM Vbias 0.04261f
C2532 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.SM 0.00168f
C2533 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC_15.icell.Ien 0.00214f
C2534 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C2535 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C2536 XA.XIR[9].XIC[1].icell.PDM Iout 0.00117f
C2537 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9] 0.00341f
C2538 XA.XIR[1].XIC[2].icell.PUM VPWR 0.00937f
C2539 XA.XIR[9].XIC[9].icell.Ien VPWR 0.1903f
C2540 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00584f
C2541 XA.XIR[13].XIC_15.icell.PDM Vbias 0.04401f
C2542 XA.XIR[10].XIC[3].icell.PUM VPWR 0.00937f
C2543 XA.XIR[1].XIC[5].icell.Ien Vbias 0.21104f
C2544 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00584f
C2545 XThC.Tn[14] XThR.Tn[11] 0.28745f
C2546 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.SM 0.00168f
C2547 XA.XIR[14].XIC[9].icell.PUM Vbias 0.0031f
C2548 XA.XIR[12].XIC[12].icell.SM Iout 0.00388f
C2549 XA.XIR[9].XIC[5].icell.Ien Iout 0.06417f
C2550 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18966f
C2551 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C2552 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C2553 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.15202f
C2554 XThC.Tn[4] XThR.Tn[7] 0.28739f
C2555 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C2556 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04031f
C2557 XA.XIR[11].XIC[14].icell.PDM VPWR 0.00809f
C2558 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04031f
C2559 XA.XIR[8].XIC[13].icell.Ien Vbias 0.21098f
C2560 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04031f
C2561 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02771f
C2562 XThC.XTB7.B XThC.Tn[2] 0.00273f
C2563 XA.XIR[3].XIC[12].icell.PUM VPWR 0.00937f
C2564 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.SM 0.00168f
C2565 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10] 0.00341f
C2566 XThC.XTB7.Y XThC.Tn[6] 0.2144f
C2567 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14] 0.00341f
C2568 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.SM 0.00168f
C2569 XThC.Tn[1] Vbias 2.40549f
C2570 XA.XIR[1].XIC[6].icell.PDM Iout 0.00117f
C2571 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02762f
C2572 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C2573 XThC.XTB6.Y XThC.Tn[10] 0.02461f
C2574 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07214f
C2575 XA.XIR[6].XIC[11].icell.SM Iout 0.00388f
C2576 XA.XIR[2].XIC[5].icell.PUM VPWR 0.00937f
C2577 XA.XIR[14].XIC_15.icell.Ien VPWR 0.25598f
C2578 XA.XIR[7].XIC[5].icell.Ien VPWR 0.1903f
C2579 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PUM 0.00465f
C2580 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.03425f
C2581 XA.XIR[4].XIC[6].icell.PDM Iout 0.00117f
C2582 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Iout 0.00347f
C2583 XA.XIR[5].XIC[14].icell.Ien Iout 0.06417f
C2584 XA.XIR[1].XIC[7].icell.PUM VPWR 0.00937f
C2585 XThC.Tn[8] XThR.Tn[1] 0.28739f
C2586 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.SM 0.00168f
C2587 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PUM 0.00429f
C2588 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11] 0.00341f
C2589 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.15202f
C2590 XA.XIR[3].XIC[14].icell.PDM Iout 0.00117f
C2591 XA.XIR[0].XIC_15.icell.Ien Vbias 0.21265f
C2592 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.SM 0.0039f
C2593 XA.XIR[14].XIC[5].icell.SM Iout 0.00388f
C2594 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.SM 0.00168f
C2595 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.15202f
C2596 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01577f
C2597 XThR.Tn[7] XA.XIR[8].XIC[2].icell.Ien 0.00338f
C2598 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C2599 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C2600 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02762f
C2601 XThC.Tn[8] XThR.Tn[12] 0.28739f
C2602 XThR.Tn[6] XA.XIR[7].XIC[13].icell.Ien 0.00338f
C2603 XA.XIR[13].XIC[7].icell.SM Iout 0.00388f
C2604 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C2605 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00584f
C2606 XA.XIR[11].XIC_dummy_right.icell.SM VPWR 0.00123f
C2607 XA.XIR[6].XIC[0].icell.Ien Vbias 0.20951f
C2608 XA.XIR[12].XIC[9].icell.Ien Iout 0.06417f
C2609 XThR.Tn[2] XA.XIR[3].XIC[4].icell.SM 0.00121f
C2610 XThC.Tn[3] XThR.Tn[3] 0.28739f
C2611 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.SM 0.0039f
C2612 XThR.Tn[4] XA.XIR[5].XIC[11].icell.SM 0.00121f
C2613 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C2614 XThR.Tn[1] XA.XIR[1].XIC_15.icell.PDM 0.00341f
C2615 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14] 0.00341f
C2616 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00584f
C2617 XA.XIR[14].XIC[0].icell.PUM VPWR 0.00937f
C2618 XThC.Tn[12] XThR.Tn[4] 0.28739f
C2619 XThR.Tn[10] XA.XIR[11].XIC[3].icell.Ien 0.00338f
C2620 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04052f
C2621 XThR.Tn[3] XA.XIR[3].XIC[0].icell.PDM 0.00347f
C2622 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2623 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.15202f
C2624 XThR.Tn[3] XA.XIR[4].XIC[11].icell.SM 0.00121f
C2625 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.03425f
C2626 a_2979_9615# VPWR 0.70527f
C2627 XA.XIR[11].XIC[4].icell.PDM Vbias 0.04261f
C2628 XA.XIR[9].XIC[0].icell.Ien Iout 0.06411f
C2629 XThR.Tn[11] XA.XIR[12].XIC[13].icell.SM 0.00121f
C2630 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.15202f
C2631 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.15202f
C2632 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.15202f
C2633 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04031f
C2634 XThC.XTB4.Y XThC.Tn[10] 0.01391f
C2635 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.SM 0.00168f
C2636 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.03425f
C2637 XA.XIR[10].XIC[8].icell.PDM Vbias 0.04261f
C2638 XA.XIR[5].XIC[3].icell.PDM VPWR 0.00799f
C2639 XThR.Tn[2] XA.XIR[2].XIC[12].icell.PDM 0.00341f
C2640 XThC.XTB4.Y a_4861_9615# 0.23756f
C2641 XThC.Tn[6] XThR.Tn[0] 0.28748f
C2642 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[8].icell.Ien 0.00214f
C2643 XA.XIR[8].XIC_15.icell.SM Iout 0.0047f
C2644 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.04036f
C2645 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02762f
C2646 XA.XIR[6].XIC[2].icell.PUM VPWR 0.00937f
C2647 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C2648 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.15202f
C2649 XA.XIR[6].XIC[5].icell.Ien Vbias 0.21098f
C2650 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00214f
C2651 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PUM 0.00465f
C2652 XThC.XTB5.Y a_7875_9569# 0.00418f
C2653 XA.XIR[12].XIC[2].icell.PDM VPWR 0.00799f
C2654 XThC.Tn[12] XThC.Tn[13] 0.23689f
C2655 XA.XIR[2].XIC[14].icell.SM Iout 0.00388f
C2656 XA.XIR[15].XIC[6].icell.SM Vbias 0.00701f
C2657 XA.XIR[12].XIC[10].icell.SM Iout 0.00388f
C2658 XA.XIR[5].XIC[8].icell.PUM Vbias 0.0031f
C2659 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C2660 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.SM 0.00168f
C2661 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02762f
C2662 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.03425f
C2663 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C2664 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.SM 0.00168f
C2665 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PUM 0.00465f
C2666 XA.XIR[11].XIC[8].icell.PDM VPWR 0.00799f
C2667 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02762f
C2668 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02762f
C2669 XA.XIR[4].XIC[9].icell.SM Vbias 0.00701f
C2670 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C2671 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00584f
C2672 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.SM 0.00168f
C2673 XA.XIR[0].XIC[0].icell.SM Vbias 0.00691f
C2674 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00256f
C2675 XA.XIR[2].XIC[0].icell.PDM Vbias 0.04207f
C2676 XA.XIR[8].XIC[3].icell.SM Vbias 0.00701f
C2677 XA.XIR[10].XIC[0].icell.PDM Iout 0.00117f
C2678 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.03425f
C2679 XA.XIR[3].XIC[2].icell.Ien VPWR 0.1903f
C2680 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04037f
C2681 XA.XIR[10].XIC[13].icell.PDM Vbias 0.04261f
C2682 XA.XIR[6].XIC[7].icell.PUM VPWR 0.00937f
C2683 XA.XIR[12].XIC[3].icell.PUM Vbias 0.0031f
C2684 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.03425f
C2685 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Ien 0.00214f
C2686 XA.XIR[7].XIC_dummy_left.icell.SM VPWR 0.00269f
C2687 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.SM 0.00168f
C2688 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C2689 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00214f
C2690 XA.XIR[15].XIC[8].icell.Ien VPWR 0.32895f
C2691 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02762f
C2692 XA.XIR[11].XIC[4].icell.Ien Vbias 0.21098f
C2693 XA.XIR[5].XIC[8].icell.SM VPWR 0.00158f
C2694 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00214f
C2695 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.15202f
C2696 XThC.XTBN.Y a_7875_9569# 0.229f
C2697 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00584f
C2698 XA.XIR[13].XIC[14].icell.PDM Vbias 0.04261f
C2699 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[1].icell.Ien 0.00214f
C2700 XA.XIR[15].XIC[4].icell.Ien Iout 0.06807f
C2701 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.15202f
C2702 XA.XIR[5].XIC[4].icell.SM Iout 0.00388f
C2703 XA.XIR[9].XIC[12].icell.SM Vbias 0.00701f
C2704 XA.XIR[10].XIC[6].icell.Ien Vbias 0.21098f
C2705 XA.XIR[4].XIC[11].icell.Ien VPWR 0.1903f
C2706 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C2707 XA.XIR[8].XIC[0].icell.PDM VPWR 0.00799f
C2708 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C2709 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C2710 XThC.Tn[5] XThR.Tn[2] 0.28739f
C2711 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.SM 0.0039f
C2712 XA.XIR[11].XIC[13].icell.PDM VPWR 0.00799f
C2713 XA.XIR[4].XIC[7].icell.Ien Iout 0.06417f
C2714 XA.XIR[2].XIC[4].icell.PDM VPWR 0.00799f
C2715 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PUM 0.00465f
C2716 XA.XIR[0].XIC[5].icell.SM Vbias 0.00716f
C2717 XA.XIR[13].XIC[3].icell.PUM VPWR 0.00937f
C2718 XThC.Tn[14] XThR.Tn[14] 0.28745f
C2719 XA.XIR[8].XIC[5].icell.Ien VPWR 0.1903f
C2720 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.SM 0.00168f
C2721 XThR.Tn[6] XA.XIR[7].XIC[3].icell.SM 0.00121f
C2722 XA.XIR[3].XIC_15.icell.Ien Vbias 0.21234f
C2723 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C2724 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.03425f
C2725 XA.XIR[12].XIC[3].icell.SM VPWR 0.00158f
C2726 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PUM 0.00465f
C2727 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C2728 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C2729 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C2730 XA.XIR[14].XIC[14].icell.PDM VPWR 0.00809f
C2731 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.SM 0.00168f
C2732 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00584f
C2733 XA.XIR[1].XIC_dummy_left.icell.Ien Vbias 0.00393f
C2734 XA.XIR[11].XIC[6].icell.PUM VPWR 0.00937f
C2735 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Ien 0.00584f
C2736 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.SM 0.0039f
C2737 XA.XIR[2].XIC[8].icell.Ien Vbias 0.21098f
C2738 a_n1335_4229# data[4] 0.00451f
C2739 XA.XIR[7].XIC[8].icell.SM Vbias 0.00701f
C2740 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00214f
C2741 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04031f
C2742 XThR.Tn[11] XA.XIR[12].XIC[11].icell.SM 0.00121f
C2743 XA.XIR[7].XIC[1].icell.Ien Iout 0.06417f
C2744 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C2745 XA.XIR[9].XIC[14].icell.Ien VPWR 0.19036f
C2746 XThC.XTB2.Y XThC.Tn[10] 0.00106f
C2747 XA.XIR[10].XIC[8].icell.PUM VPWR 0.00937f
C2748 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C2749 XA.XIR[4].XIC_dummy_left.icell.Ien Vbias 0.00329f
C2750 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.SM 0.00168f
C2751 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11] 0.00341f
C2752 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02762f
C2753 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00256f
C2754 XA.XIR[1].XIC[10].icell.Ien Vbias 0.21104f
C2755 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[14].icell.Ien 0.00214f
C2756 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Iout 0.00347f
C2757 XThR.Tn[14] XA.XIR[15].XIC[3].icell.SM 0.00121f
C2758 XA.XIR[9].XIC[10].icell.Ien Iout 0.06417f
C2759 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C2760 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C2761 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18965f
C2762 XThC.XTB2.Y a_4861_9615# 0.00851f
C2763 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.15202f
C2764 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.SM 0.0039f
C2765 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[9].icell.Ien 0.00214f
C2766 XThC.Tn[1] XThR.Tn[6] 0.28739f
C2767 XA.XIR[12].XIC[14].icell.Ien Iout 0.06417f
C2768 XA.XIR[0].XIC[3].icell.Ien Iout 0.06389f
C2769 XThC.Tn[12] data[3] 0.00161f
C2770 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04031f
C2771 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.03023f
C2772 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2773 XThC.XTBN.A XThC.Tn[12] 0.22686f
C2774 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.Ien 0.00584f
C2775 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C2776 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.SM 0.00168f
C2777 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04031f
C2778 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8] 0.00341f
C2779 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02762f
C2780 XThR.Tn[5] a_n1049_5611# 0.27042f
C2781 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14] 0.00341f
C2782 XA.XIR[7].XIC[10].icell.Ien VPWR 0.1903f
C2783 XA.XIR[2].XIC[10].icell.PUM VPWR 0.00937f
C2784 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00584f
C2785 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C2786 XThC.Tn[3] XThR.Tn[11] 0.28739f
C2787 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.389f
C2788 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.SM 0.0039f
C2789 XA.XIR[1].XIC[12].icell.PUM VPWR 0.00937f
C2790 XA.XIR[7].XIC[6].icell.Ien Iout 0.06417f
C2791 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[5].icell.Ien 0.00214f
C2792 XA.XIR[14].XIC_dummy_right.icell.SM VPWR 0.00123f
C2793 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.Ien 0.00584f
C2794 XA.XIR[10].XIC[0].icell.SM Vbias 0.00675f
C2795 XA.XIR[7].XIC[0].icell.PDM Vbias 0.04207f
C2796 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04031f
C2797 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.SM 0.00168f
C2798 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.03425f
C2799 XThC.XTBN.Y Iout 0.00167f
C2800 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.03425f
C2801 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C2802 XA.XIR[6].XIC[7].icell.PDM Vbias 0.04261f
C2803 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C2804 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.SM 0.0039f
C2805 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C2806 XThR.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.00338f
C2807 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.15202f
C2808 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.SM 0.0039f
C2809 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.03425f
C2810 XA.XIR[8].XIC[0].icell.Ien VPWR 0.1903f
C2811 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00584f
C2812 XA.XIR[5].XIC[14].icell.PDM Vbias 0.04261f
C2813 XA.XIR[14].XIC[4].icell.PDM Vbias 0.04261f
C2814 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00214f
C2815 XThC.XTB5.Y XThC.Tn[4] 0.19958f
C2816 a_10915_9569# XThC.Tn[13] 0.01061f
C2817 XThR.Tn[5] XA.XIR[6].XIC[3].icell.Ien 0.00338f
C2818 XThC.XTB6.Y a_7651_9569# 0.0046f
C2819 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.03425f
C2820 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.SM 0.0039f
C2821 XA.XIR[13].XIC[8].icell.PDM Vbias 0.04261f
C2822 XThR.Tn[2] XA.XIR[3].XIC[9].icell.SM 0.00121f
C2823 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Ien 0.00584f
C2824 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00214f
C2825 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C2826 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PUM 0.00465f
C2827 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00584f
C2828 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04031f
C2829 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.15202f
C2830 XThR.Tn[4] XA.XIR[4].XIC[14].icell.PDM 0.00341f
C2831 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02762f
C2832 XA.XIR[7].XIC[4].icell.PDM VPWR 0.00799f
C2833 XThC.Tn[6] XThR.Tn[1] 0.2874f
C2834 XThR.Tn[3] XA.XIR[3].XIC_15.icell.PDM 0.00341f
C2835 XThR.Tn[10] XA.XIR[11].XIC[8].icell.Ien 0.00338f
C2836 XThR.XTB6.A XThR.XTB7.A 0.44014f
C2837 XThC.Tn[10] Iout 0.83837f
C2838 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C2839 XThC.Tn[10] XThR.Tn[9] 0.28739f
C2840 XA.XIR[9].XIC[4].icell.PUM Vbias 0.0031f
C2841 XA.XIR[6].XIC[11].icell.PDM VPWR 0.00799f
C2842 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.15202f
C2843 XA.XIR[4].XIC[1].icell.SM VPWR 0.00158f
C2844 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00214f
C2845 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.SM 0.00168f
C2846 XA.XIR[15].XIC[2].icell.PDM VPWR 0.0114f
C2847 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PUM 0.00465f
C2848 XThR.XTB5.A XThR.Tn[8] 0.00204f
C2849 XThC.Tn[6] XThR.Tn[12] 0.28739f
C2850 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.15202f
C2851 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02762f
C2852 XA.XIR[11].XIC[12].icell.SM Vbias 0.00701f
C2853 XA.XIR[14].XIC[8].icell.PDM VPWR 0.00799f
C2854 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C2855 XThR.XTB5.Y a_n997_1803# 0.06458f
C2856 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.PDM 0.0059f
C2857 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C2858 XA.XIR[15].XIC[12].icell.SM Iout 0.00388f
C2859 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Iout 0.00347f
C2860 XA.XIR[10].XIC[12].icell.PDM Vbias 0.04261f
C2861 XA.XIR[5].XIC[6].icell.PDM Iout 0.00117f
C2862 XThR.Tn[11] XA.XIR[12].XIC[9].icell.SM 0.00121f
C2863 XA.XIR[3].XIC[5].icell.SM Vbias 0.00701f
C2864 XThC.XTBN.Y XThC.Tn[4] 0.61061f
C2865 XA.XIR[1].XIC[1].icell.PDM Vbias 0.04261f
C2866 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00584f
C2867 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.Ien 0.00584f
C2868 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.15202f
C2869 XThC.Tn[1] XThR.Tn[4] 0.28739f
C2870 XA.XIR[6].XIC[10].icell.Ien Vbias 0.21098f
C2871 XA.XIR[9].XIC[0].icell.PDM VPWR 0.00799f
C2872 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[13].icell.Ien 0.00214f
C2873 XA.XIR[13].XIC[0].icell.PDM Iout 0.00117f
C2874 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.SM 0.00168f
C2875 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PUM 0.00465f
C2876 XA.XIR[4].XIC[1].icell.PDM Vbias 0.04261f
C2877 XA.XIR[5].XIC[13].icell.PUM Vbias 0.0031f
C2878 XA.XIR[13].XIC[13].icell.PDM Vbias 0.04261f
C2879 XThR.Tn[1] XA.XIR[2].XIC[0].icell.Ien 0.00338f
C2880 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.SM 0.0039f
C2881 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2882 XA.XIR[9].XIC[4].icell.SM VPWR 0.00158f
C2883 XA.XIR[12].XIC[5].icell.PDM Iout 0.00117f
C2884 XA.XIR[12].XIC[12].icell.Ien Iout 0.06417f
C2885 XThC.XTB4.Y a_7651_9569# 0.00497f
C2886 XA.XIR[4].XIC[14].icell.SM Vbias 0.00701f
C2887 XA.XIR[3].XIC[9].icell.PDM Vbias 0.04261f
C2888 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02762f
C2889 XA.XIR[8].XIC[11].icell.PDM Vbias 0.04261f
C2890 XA.XIR[14].XIC[4].icell.Ien Vbias 0.21098f
C2891 XThC.Tn[5] XThR.Tn[10] 0.28739f
C2892 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.03425f
C2893 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.03425f
C2894 XA.XIR[11].XIC[12].icell.PDM VPWR 0.00799f
C2895 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00214f
C2896 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C2897 XA.XIR[2].XIC_15.icell.PDM Vbias 0.04401f
C2898 XA.XIR[13].XIC[6].icell.Ien Vbias 0.21098f
C2899 XA.XIR[8].XIC[8].icell.SM Vbias 0.00701f
C2900 XThC.Tn[0] XA.XIR[4].XIC_dummy_left.icell.Iout 0.00109f
C2901 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.SM 0.0039f
C2902 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00584f
C2903 XA.XIR[1].XIC[5].icell.PDM VPWR 0.00799f
C2904 XA.XIR[8].XIC[1].icell.Ien Iout 0.06417f
C2905 XA.XIR[3].XIC[7].icell.Ien VPWR 0.1903f
C2906 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C2907 XThR.Tn[8] XA.XIR[9].XIC[1].icell.Ien 0.00338f
C2908 XA.XIR[11].XIC_15.icell.PUM Vbias 0.0031f
C2909 XA.XIR[12].XIC[8].icell.PUM Vbias 0.0031f
C2910 XA.XIR[14].XIC[13].icell.PDM VPWR 0.00799f
C2911 XA.XIR[6].XIC[12].icell.PUM VPWR 0.00937f
C2912 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00584f
C2913 XA.XIR[3].XIC[3].icell.Ien Iout 0.06417f
C2914 a_4861_9615# XThC.Tn[4] 0.00198f
C2915 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[4].icell.Ien 0.00214f
C2916 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7] 0.00341f
C2917 XA.XIR[11].XIC[9].icell.Ien Vbias 0.21098f
C2918 XA.XIR[4].XIC[5].icell.PDM VPWR 0.00799f
C2919 XA.XIR[5].XIC[13].icell.SM VPWR 0.00158f
C2920 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.SM 0.0039f
C2921 XThR.XTB5.Y XThR.Tn[13] 0.00145f
C2922 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04031f
C2923 XThC.XTBN.Y XA.XIR[0].XIC[11].icell.PDM 0.00104f
C2924 XA.XIR[15].XIC[9].icell.Ien Iout 0.06807f
C2925 XA.XIR[5].XIC[9].icell.SM Iout 0.00388f
C2926 XA.XIR[1].XIC[2].icell.Ien VPWR 0.1903f
C2927 XA.XIR[3].XIC[13].icell.PDM VPWR 0.00799f
C2928 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07214f
C2929 XA.XIR[14].XIC[6].icell.PUM VPWR 0.00937f
C2930 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13] 0.00341f
C2931 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.03426f
C2932 XA.XIR[8].XIC[3].icell.PDM Iout 0.00117f
C2933 XA.XIR[3].XIC[1].icell.PDM Iout 0.00117f
C2934 XA.XIR[4].XIC[12].icell.Ien Iout 0.06417f
C2935 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PUM 0.00465f
C2936 XA.XIR[13].XIC[8].icell.PUM VPWR 0.00937f
C2937 XA.XIR[0].XIC[10].icell.SM Vbias 0.00716f
C2938 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04031f
C2939 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04031f
C2940 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.SM 0.0039f
C2941 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C2942 XA.XIR[8].XIC[10].icell.Ien VPWR 0.1903f
C2943 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PUM 0.00444f
C2944 XA.XIR[2].XIC[7].icell.PDM Iout 0.00117f
C2945 XThR.Tn[6] XA.XIR[7].XIC[8].icell.SM 0.00121f
C2946 XA.XIR[12].XIC[8].icell.SM VPWR 0.00158f
C2947 XA.XIR[8].XIC[6].icell.Ien Iout 0.06417f
C2948 XThR.Tn[8] XA.XIR[9].XIC[6].icell.Ien 0.00338f
C2949 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14] 0.00341f
C2950 XA.XIR[12].XIC[4].icell.SM Iout 0.00388f
C2951 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.SM 0.00168f
C2952 XThR.Tn[0] XA.XIR[0].XIC[4].icell.PDM 0.00341f
C2953 XA.XIR[2].XIC[13].icell.Ien Vbias 0.21098f
C2954 XA.XIR[7].XIC[13].icell.SM Vbias 0.00701f
C2955 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.SM 0.0039f
C2956 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00214f
C2957 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PUM 0.00465f
C2958 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2959 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2960 XA.XIR[1].XIC[1].icell.PUM Vbias 0.0031f
C2961 XThR.Tn[1] XA.XIR[1].XIC[2].icell.PDM 0.00341f
C2962 XThR.Tn[0] XA.XIR[1].XIC[1].icell.Ien 0.00338f
C2963 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C2964 XA.XIR[1].XIC_15.icell.Ien Vbias 0.2124f
C2965 XThR.Tn[11] XA.XIR[12].XIC[13].icell.Ien 0.00338f
C2966 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C2967 XA.XIR[11].XIC[10].icell.SM Vbias 0.00701f
C2968 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04031f
C2969 XThR.Tn[14] XA.XIR[15].XIC[8].icell.SM 0.00121f
C2970 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02762f
C2971 XThC.Tn[3] XThR.Tn[14] 0.28739f
C2972 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.SM 0.00168f
C2973 XA.XIR[9].XIC_15.icell.Ien Iout 0.0642f
C2974 XA.XIR[4].XIC[1].icell.PUM Vbias 0.0031f
C2975 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C2976 XThC.XTB5.Y a_6243_9615# 0.00907f
C2977 XA.XIR[15].XIC[10].icell.SM Iout 0.00388f
C2978 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00214f
C2979 XA.XIR[0].XIC[12].icell.Ien VPWR 0.19211f
C2980 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.SM 0.00168f
C2981 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5] 0.00341f
C2982 XA.XIR[8].XIC_dummy_left.icell.SM VPWR 0.00269f
C2983 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Ien 0.00584f
C2984 XA.XIR[13].XIC[0].icell.SM Vbias 0.00675f
C2985 XA.XIR[0].XIC_dummy_right.icell.Ien Vbias 0.00307f
C2986 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.03425f
C2987 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.SM 0.0039f
C2988 XThC.XTB7.A a_5155_9615# 0.02287f
C2989 XA.XIR[0].XIC[8].icell.Ien Iout 0.06389f
C2990 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C2991 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PUM 0.00465f
C2992 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[12].icell.Ien 0.00214f
C2993 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C2994 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.SM 0.0039f
C2995 XThR.Tn[13] XA.XIR[14].XIC[3].icell.Ien 0.00338f
C2996 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04035f
C2997 XThC.XTB4.Y data[2] 0.0086f
C2998 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01577f
C2999 XA.XIR[7].XIC_15.icell.Ien VPWR 0.25566f
C3000 XA.XIR[12].XIC[10].icell.Ien Iout 0.06417f
C3001 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.SM 0.00168f
C3002 XThC.XTB2.Y a_7651_9569# 0.00191f
C3003 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.15202f
C3004 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6] 0.00341f
C3005 XA.XIR[5].XIC[0].icell.Ien VPWR 0.1903f
C3006 XA.XIR[15].XIC[3].icell.PUM Vbias 0.0031f
C3007 XA.XIR[7].XIC[11].icell.Ien Iout 0.06417f
C3008 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C3009 XA.XIR[5].XIC[3].icell.Ien Vbias 0.21098f
C3010 XA.XIR[7].XIC_15.icell.PDM Vbias 0.04401f
C3011 XThR.Tn[0] XA.XIR[1].XIC[6].icell.Ien 0.00338f
C3012 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C3013 XThR.XTB7.B XThR.XTB6.A 1.47641f
C3014 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C3015 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PUM 0.00465f
C3016 XA.XIR[14].XIC[1].icell.PUM VPWR 0.00937f
C3017 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PUM 0.00465f
C3018 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C3019 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00214f
C3020 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.1106f
C3021 XThC.Tn[14] VPWR 6.85545f
C3022 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.SM 0.00168f
C3023 XA.XIR[4].XIC[6].icell.PUM Vbias 0.0031f
C3024 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PUM 0.00465f
C3025 XThR.Tn[11] XA.XIR[12].XIC[14].icell.SM 0.00121f
C3026 XThR.Tn[7] XA.XIR[8].XIC[12].icell.Ien 0.00338f
C3027 XA.XIR[11].XIC[13].icell.PUM Vbias 0.0031f
C3028 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.SM 0.00168f
C3029 XThC.XTBN.Y a_6243_9615# 0.07731f
C3030 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C3031 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02762f
C3032 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C3033 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C3034 XA.XIR[10].XIC[11].icell.PDM Vbias 0.04261f
C3035 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PUM 0.00465f
C3036 XA.XIR[3].XIC[0].icell.Ien Iout 0.06411f
C3037 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PUM 0.00465f
C3038 XThR.Tn[8] Iout 1.16233f
C3039 XThR.Tn[5] XA.XIR[6].XIC[8].icell.Ien 0.00338f
C3040 XThR.Tn[8] XThR.Tn[9] 0.05786f
C3041 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C3042 XA.XIR[14].XIC[12].icell.SM Vbias 0.00701f
C3043 XThR.Tn[2] XA.XIR[3].XIC[14].icell.SM 0.00121f
C3044 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3045 XA.XIR[6].XIC[2].icell.Ien VPWR 0.1903f
C3046 XA.XIR[9].XIC[11].icell.PDM Vbias 0.04261f
C3047 XA.XIR[0].XIC[3].icell.PDM Vbias 0.04278f
C3048 XA.XIR[13].XIC[12].icell.PDM Vbias 0.04261f
C3049 XA.XIR[15].XIC[3].icell.SM VPWR 0.00158f
C3050 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01734f
C3051 XA.XIR[5].XIC[5].icell.PUM VPWR 0.00937f
C3052 XA.XIR[11].XIC[1].icell.Ien Iout 0.06417f
C3053 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00584f
C3054 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C3055 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3056 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.SM 0.0039f
C3057 XA.XIR[2].XIC_15.icell.SM Iout 0.0047f
C3058 XA.XIR[1].XIC[0].icell.SM Vbias 0.00679f
C3059 XA.XIR[9].XIC[9].icell.PUM Vbias 0.0031f
C3060 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01432f
C3061 XA.XIR[10].XIC[1].icell.SM Vbias 0.00701f
C3062 XA.XIR[7].XIC[7].icell.PDM Iout 0.00117f
C3063 XA.XIR[11].XIC[11].icell.PDM VPWR 0.00799f
C3064 XA.XIR[9].XIC[0].icell.SM Iout 0.00388f
C3065 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01785f
C3066 XA.XIR[4].XIC[6].icell.SM VPWR 0.00158f
C3067 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00584f
C3068 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.15202f
C3069 XA.XIR[4].XIC[2].icell.SM Iout 0.00388f
C3070 XA.XIR[6].XIC[14].icell.PDM Iout 0.00117f
C3071 XA.XIR[15].XIC[5].icell.PDM Iout 0.00117f
C3072 XThR.XTB2.Y data[5] 0.017f
C3073 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C3074 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.SM 0.0039f
C3075 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PUM 0.00465f
C3076 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[13].icell.Ien 0.00214f
C3077 XThC.Tn[5] XThR.Tn[13] 0.28739f
C3078 XThR.Tn[6] Vbias 3.74624f
C3079 XA.XIR[14].XIC[12].icell.PDM VPWR 0.00799f
C3080 XA.XIR[11].XIC[14].icell.Ien Vbias 0.21098f
C3081 XA.XIR[3].XIC[10].icell.SM Vbias 0.00701f
C3082 XA.XIR[6].XIC_15.icell.Ien Vbias 0.21234f
C3083 XA.XIR[15].XIC[14].icell.Ien Iout 0.06807f
C3084 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07214f
C3085 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PUM 0.00465f
C3086 XThR.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.00338f
C3087 XA.XIR[7].XIC[0].icell.SM VPWR 0.00158f
C3088 XA.XIR[0].XIC[7].icell.PDM VPWR 0.00773f
C3089 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.SM 0.00168f
C3090 XA.XIR[2].XIC[3].icell.SM Vbias 0.00701f
C3091 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.SM 0.0039f
C3092 XA.XIR[9].XIC[3].icell.PDM Iout 0.00117f
C3093 XA.XIR[14].XIC_15.icell.PUM Vbias 0.0031f
C3094 XA.XIR[7].XIC[5].icell.PUM Vbias 0.0031f
C3095 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9] 0.00341f
C3096 XThR.Tn[0] XThR.Tn[2] 0.00536f
C3097 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C3098 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C3099 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PUM 0.00465f
C3100 XA.XIR[9].XIC[9].icell.SM VPWR 0.00158f
C3101 XThC.Tn[4] XThR.Tn[8] 0.28739f
C3102 XThR.Tn[12] XA.XIR[13].XIC[1].icell.Ien 0.00338f
C3103 XA.XIR[10].XIC[3].icell.Ien VPWR 0.1903f
C3104 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.SM 0.00168f
C3105 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C3106 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C3107 XA.XIR[1].XIC[5].icell.SM Vbias 0.00704f
C3108 XA.XIR[14].XIC[9].icell.Ien Vbias 0.21098f
C3109 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C3110 XA.XIR[12].XIC[13].icell.SM VPWR 0.00158f
C3111 XA.XIR[9].XIC[5].icell.SM Iout 0.00388f
C3112 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[11].icell.Ien 0.00214f
C3113 XA.XIR[0].XIC[2].icell.SM VPWR 0.00158f
C3114 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04031f
C3115 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.SM 0.0039f
C3116 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.SM 0.00168f
C3117 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04052f
C3118 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00214f
C3119 XA.XIR[8].XIC[13].icell.SM Vbias 0.00701f
C3120 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04031f
C3121 XA.XIR[3].XIC[12].icell.Ien VPWR 0.1903f
C3122 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C3123 XA.XIR[2].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3124 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10] 0.00341f
C3125 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C3126 XA.XIR[3].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3127 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14] 0.00341f
C3128 XA.XIR[3].XIC[8].icell.Ien Iout 0.06417f
C3129 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C3130 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C3131 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Iout 0.00347f
C3132 XA.XIR[1].XIC[8].icell.PDM Iout 0.00117f
C3133 XThR.Tn[14] XA.XIR[15].XIC[13].icell.SM 0.00121f
C3134 XA.XIR[2].XIC[5].icell.Ien VPWR 0.1903f
C3135 XA.XIR[7].XIC[5].icell.SM VPWR 0.00158f
C3136 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00214f
C3137 XA.XIR[9].XIC[0].icell.PUM VPWR 0.00937f
C3138 XA.XIR[11].XIC[11].icell.PUM Vbias 0.0031f
C3139 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.SM 0.0039f
C3140 XThC.Tn[5] XA.XIR[0].XIC[6].icell.PDM 0.00343f
C3141 XA.XIR[4].XIC[8].icell.PDM Iout 0.00117f
C3142 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C3143 XA.XIR[1].XIC[7].icell.Ien VPWR 0.1903f
C3144 a_6243_10571# VPWR 0.00653f
C3145 XA.XIR[7].XIC[1].icell.SM Iout 0.00388f
C3146 XA.XIR[5].XIC[14].icell.SM Iout 0.00388f
C3147 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.15202f
C3148 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00214f
C3149 XThC.XTB6.Y a_5949_9615# 0.26831f
C3150 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.03511f
C3151 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C3152 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.04494f
C3153 XThC.Tn[1] XThC.Tn[2] 0.72045f
C3154 XThC.Tn[0] XThC.Tn[3] 0.12427f
C3155 XA.XIR[1].XIC[3].icell.Ien Iout 0.06417f
C3156 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C3157 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02762f
C3158 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.15202f
C3159 XThR.Tn[7] XA.XIR[8].XIC[2].icell.SM 0.00121f
C3160 XA.XIR[14].XIC[10].icell.SM Vbias 0.00701f
C3161 XA.XIR[8].XIC_15.icell.Ien VPWR 0.25566f
C3162 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02762f
C3163 XA.XIR[12].XIC_15.icell.Ien Iout 0.0642f
C3164 XThR.Tn[6] XA.XIR[7].XIC[13].icell.SM 0.00121f
C3165 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02762f
C3166 XThR.XTB7.A a_n1049_5317# 0.02018f
C3167 XA.XIR[5].XIC[1].icell.PDM Vbias 0.04261f
C3168 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.SM 0.0039f
C3169 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.SM 0.00168f
C3170 XA.XIR[8].XIC[11].icell.Ien Iout 0.06417f
C3171 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.PDM 0.00578f
C3172 XThR.Tn[8] XA.XIR[9].XIC[11].icell.Ien 0.00338f
C3173 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C3174 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00584f
C3175 XA.XIR[6].XIC[0].icell.SM Vbias 0.00675f
C3176 XThC.XTB5.A XThC.XTB6.Y 0.00193f
C3177 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.SM 0.0039f
C3178 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.SM 0.0039f
C3179 XThR.Tn[4] XA.XIR[4].XIC[1].icell.PDM 0.00341f
C3180 XThR.Tn[4] Vbias 3.74761f
C3181 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C3182 XA.XIR[5].XIC_dummy_left.icell.SM VPWR 0.00269f
C3183 XA.XIR[12].XIC[0].icell.PDM Vbias 0.04207f
C3184 XThR.Tn[10] XA.XIR[11].XIC[3].icell.SM 0.00121f
C3185 XThR.Tn[3] XA.XIR[3].XIC[2].icell.PDM 0.00341f
C3186 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C3187 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PUM 0.00465f
C3188 a_4067_9615# VPWR 0.70648f
C3189 XA.XIR[11].XIC[6].icell.PDM Vbias 0.04261f
C3190 a_n997_3755# XThR.Tn[9] 0.19352f
C3191 XThR.XTB2.Y XThR.Tn[9] 0.292f
C3192 XA.XIR[11].XIC[12].icell.Ien Vbias 0.21098f
C3193 XThR.Tn[1] XA.XIR[2].XIC[4].icell.Ien 0.00338f
C3194 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.SM 0.0039f
C3195 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04031f
C3196 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[4].icell.Ien 0.00214f
C3197 XA.XIR[10].XIC[10].icell.PDM Vbias 0.04261f
C3198 XA.XIR[15].XIC[12].icell.Ien Iout 0.06807f
C3199 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C3200 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.SM 0.0039f
C3201 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.15202f
C3202 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.15202f
C3203 XA.XIR[0].XIC[13].icell.Ien Iout 0.06389f
C3204 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.03425f
C3205 XA.XIR[5].XIC[5].icell.PDM VPWR 0.00799f
C3206 XThR.XTB5.Y a_n997_3979# 0.00418f
C3207 XThR.Tn[2] XA.XIR[2].XIC[14].icell.PDM 0.00341f
C3208 XThC.XTB4.Y a_5949_9615# 0.00465f
C3209 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C3210 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3211 XA.XIR[14].XIC[13].icell.PUM Vbias 0.0031f
C3212 XThR.Tn[13] XA.XIR[14].XIC[8].icell.Ien 0.00338f
C3213 XThC.Tn[13] Vbias 2.40092f
C3214 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PDM 0.00172f
C3215 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PUM 0.00465f
C3216 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.SM 0.00168f
C3217 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C3218 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02762f
C3219 XA.XIR[6].XIC[5].icell.SM Vbias 0.00701f
C3220 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00584f
C3221 XA.XIR[13].XIC[11].icell.PDM Vbias 0.04261f
C3222 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C3223 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C3224 XThC.XTB5.Y a_8963_9569# 0.00427f
C3225 XA.XIR[12].XIC[4].icell.PDM VPWR 0.00799f
C3226 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.Ien 0.00584f
C3227 XA.XIR[7].XIC_dummy_right.icell.SM VPWR 0.00123f
C3228 XA.XIR[12].XIC[11].icell.SM VPWR 0.00158f
C3229 XA.XIR[15].XIC[8].icell.PUM Vbias 0.0031f
C3230 XThR.Tn[0] XA.XIR[1].XIC[11].icell.Ien 0.00338f
C3231 XA.XIR[5].XIC[8].icell.Ien Vbias 0.21098f
C3232 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C3233 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C3234 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.03425f
C3235 XA.XIR[11].XIC[10].icell.PDM VPWR 0.00799f
C3236 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Iout 0.00347f
C3237 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C3238 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C3239 XA.XIR[4].XIC[11].icell.PUM Vbias 0.0031f
C3240 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C3241 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C3242 XA.XIR[14].XIC[1].icell.Ien Iout 0.06417f
C3243 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.SM 0.0039f
C3244 XA.XIR[0].XIC[2].icell.PUM Vbias 0.0031f
C3245 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PUM 0.00465f
C3246 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00584f
C3247 XA.XIR[8].XIC[0].icell.SM VPWR 0.00158f
C3248 XA.XIR[2].XIC[2].icell.PDM Vbias 0.04261f
C3249 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00214f
C3250 XA.XIR[14].XIC[11].icell.PDM VPWR 0.00799f
C3251 XA.XIR[13].XIC[1].icell.SM Vbias 0.00701f
C3252 XThR.Tn[14] XA.XIR[15].XIC[11].icell.SM 0.00121f
C3253 XThR.Tn[5] XA.XIR[6].XIC[13].icell.Ien 0.00338f
C3254 XThR.XTB7.B XThR.Tn[12] 0.00772f
C3255 XA.XIR[8].XIC[5].icell.PUM Vbias 0.0031f
C3256 XA.XIR[10].XIC[2].icell.PDM Iout 0.00117f
C3257 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04031f
C3258 XA.XIR[3].XIC[2].icell.SM VPWR 0.00158f
C3259 XA.XIR[12].XIC[3].icell.Ien Vbias 0.21098f
C3260 XThC.XTB1.Y XThC.Tn[1] 0.01447f
C3261 XA.XIR[6].XIC[7].icell.Ien VPWR 0.1903f
C3262 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.SM 0.00168f
C3263 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C3264 XA.XIR[14].XIC[14].icell.Ien Vbias 0.21098f
C3265 XThR.XTB7.A a_n1049_6405# 0.02287f
C3266 XA.XIR[15].XIC[8].icell.SM VPWR 0.00158f
C3267 XThC.Tn[3] VPWR 5.90764f
C3268 XA.XIR[6].XIC[3].icell.Ien Iout 0.06417f
C3269 XA.XIR[11].XIC[4].icell.SM Vbias 0.00701f
C3270 XThR.Tn[6] XThR.XTBN.A 0.00131f
C3271 XA.XIR[5].XIC[10].icell.PUM VPWR 0.00937f
C3272 XThC.XTBN.Y a_8963_9569# 0.22784f
C3273 XA.XIR[15].XIC[4].icell.SM Iout 0.00388f
C3274 XA.XIR[9].XIC[14].icell.PUM Vbias 0.0031f
C3275 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02762f
C3276 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C3277 XA.XIR[3].XIC[0].icell.PDM VPWR 0.00799f
C3278 XA.XIR[10].XIC[6].icell.SM Vbias 0.00701f
C3279 XA.XIR[4].XIC[11].icell.SM VPWR 0.00158f
C3280 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[7].icell.Ien 0.00214f
C3281 XA.XIR[12].XIC[14].icell.PUM VPWR 0.00937f
C3282 XA.XIR[8].XIC[2].icell.PDM VPWR 0.00799f
C3283 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C3284 XThR.XTB5.A XThR.XTB7.Y 0.00179f
C3285 XThR.XTB5.A data[4] 0.14415f
C3286 XA.XIR[4].XIC_15.icell.SM Vbias 0.00701f
C3287 XThC.Tn[9] XThR.Tn[0] 0.28777f
C3288 XA.XIR[2].XIC[6].icell.PDM VPWR 0.00799f
C3289 XThC.Tn[11] XThR.Tn[5] 0.28739f
C3290 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C3291 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C3292 XA.XIR[4].XIC[7].icell.SM Iout 0.00388f
C3293 XA.XIR[0].XIC[7].icell.PUM Vbias 0.0031f
C3294 XThR.XTB5.Y XThR.Tn[7] 0.00912f
C3295 XThR.Tn[1] XThR.Tn[2] 0.10497f
C3296 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.03425f
C3297 XA.XIR[13].XIC[3].icell.Ien VPWR 0.1903f
C3298 XThR.XTB5.Y a_n997_2891# 0.00424f
C3299 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.SM 0.0039f
C3300 XA.XIR[8].XIC[5].icell.SM VPWR 0.00158f
C3301 XThR.XTB1.Y a_n997_3979# 0.06353f
C3302 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C3303 XA.XIR[12].XIC[5].icell.PUM VPWR 0.00937f
C3304 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.03425f
C3305 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00584f
C3306 XA.XIR[8].XIC[1].icell.SM Iout 0.00388f
C3307 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.SM 0.00168f
C3308 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12] 0.00341f
C3309 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.Ien 0.00584f
C3310 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PUM 0.00465f
C3311 XThR.Tn[8] XA.XIR[9].XIC[1].icell.SM 0.00121f
C3312 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C3313 XA.XIR[11].XIC[6].icell.Ien VPWR 0.1903f
C3314 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04031f
C3315 XA.XIR[7].XIC[10].icell.PUM Vbias 0.0031f
C3316 XA.XIR[2].XIC[8].icell.SM Vbias 0.00701f
C3317 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38912f
C3318 XThR.Tn[4] XA.XIR[5].XIC[3].icell.Ien 0.00338f
C3319 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.SM 0.0039f
C3320 XA.XIR[11].XIC[10].icell.Ien Vbias 0.21098f
C3321 XA.XIR[2].XIC[1].icell.Ien Iout 0.06417f
C3322 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.0353f
C3323 XA.XIR[9].XIC[14].icell.SM VPWR 0.00207f
C3324 XA.XIR[11].XIC[2].icell.Ien Iout 0.06417f
C3325 XA.XIR[10].XIC[8].icell.Ien VPWR 0.1903f
C3326 XA.XIR[1].XIC[10].icell.SM Vbias 0.00704f
C3327 XA.XIR[15].XIC[10].icell.Ien Iout 0.06807f
C3328 XThR.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.00338f
C3329 XA.XIR[9].XIC[10].icell.SM Iout 0.00388f
C3330 XA.XIR[10].XIC[4].icell.Ien Iout 0.06417f
C3331 XThC.XTB2.Y a_5949_9615# 0.00844f
C3332 XThC.XTB7.B a_6243_10571# 0.00108f
C3333 XA.XIR[0].XIC[7].icell.SM VPWR 0.00158f
C3334 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.SM 0.00168f
C3335 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PUM 0.00471f
C3336 XThR.Tn[9] XA.XIR[10].XIC[4].icell.Ien 0.00338f
C3337 XA.XIR[14].XIC[11].icell.PUM Vbias 0.0031f
C3338 XThC.XTBN.A Vbias 0.01661f
C3339 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00584f
C3340 XThR.XTB7.B a_n1049_5317# 0.01743f
C3341 XA.XIR[0].XIC[3].icell.SM Iout 0.00367f
C3342 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Iout 0.00347f
C3343 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04031f
C3344 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C3345 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02762f
C3346 data[5] data[4] 0.64735f
C3347 XA.XIR[12].XIC[9].icell.SM VPWR 0.00158f
C3348 XA.XIR[2].XIC[1].icell.PUM Vbias 0.0031f
C3349 XThR.Tn[1] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00122f
C3350 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00584f
C3351 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C3352 XA.XIR[3].XIC[13].icell.Ien Iout 0.06417f
C3353 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8] 0.00341f
C3354 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04031f
C3355 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.15202f
C3356 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[9].icell.Ien 0.00214f
C3357 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.0404f
C3358 VPWR data[6] 0.21221f
C3359 XA.XIR[2].XIC[10].icell.Ien VPWR 0.1903f
C3360 XA.XIR[11].XIC[0].icell.Ien Vbias 0.20951f
C3361 XA.XIR[7].XIC[10].icell.SM VPWR 0.00158f
C3362 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C3363 XThC.Tn[8] XThR.Tn[2] 0.28739f
C3364 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[10].icell.Ien 0.00214f
C3365 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C3366 XA.XIR[1].XIC[12].icell.Ien VPWR 0.1903f
C3367 XA.XIR[2].XIC[6].icell.Ien Iout 0.06417f
C3368 XA.XIR[7].XIC[6].icell.SM Iout 0.00388f
C3369 XThR.Tn[0] XA.XIR[1].XIC[1].icell.SM 0.00121f
C3370 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04031f
C3371 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C3372 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.15202f
C3373 XA.XIR[10].XIC[2].icell.PUM Vbias 0.0031f
C3374 XA.XIR[7].XIC[2].icell.PDM Vbias 0.04261f
C3375 XA.XIR[1].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3376 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PUM 0.00465f
C3377 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[6].icell.Ien 0.00214f
C3378 XThR.Tn[12] XA.XIR[13].XIC[2].icell.Ien 0.00338f
C3379 XThR.Tn[14] XA.XIR[15].XIC[9].icell.SM 0.00121f
C3380 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C3381 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02762f
C3382 XA.XIR[1].XIC[8].icell.Ien Iout 0.06417f
C3383 XA.XIR[6].XIC[9].icell.PDM Vbias 0.04261f
C3384 XA.XIR[15].XIC[0].icell.PDM Vbias 0.04207f
C3385 XThR.XTBN.Y XA.XIR[6].XIC_dummy_left.icell.Ien 0.00159f
C3386 XThR.Tn[7] XA.XIR[8].XIC[7].icell.SM 0.00121f
C3387 XThR.XTB1.Y XThR.Tn[7] 0.00426f
C3388 a_n1335_4229# VPWR 0.00633f
C3389 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PUM 0.00465f
C3390 XA.XIR[14].XIC[6].icell.PDM Vbias 0.04261f
C3391 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C3392 XA.XIR[14].XIC[12].icell.Ien Vbias 0.21098f
C3393 XA.XIR[8].XIC_dummy_right.icell.SM VPWR 0.00123f
C3394 XThR.Tn[11] XA.XIR[12].XIC[5].icell.Ien 0.00338f
C3395 XThR.Tn[5] XA.XIR[6].XIC[3].icell.SM 0.00121f
C3396 XThC.XTB6.A XThC.Tn[9] 0.00838f
C3397 XThC.XTB6.Y a_8739_9569# 0.00466f
C3398 XA.XIR[13].XIC[10].icell.PDM Vbias 0.04261f
C3399 XThC.XTB7.A XThC.Tn[4] 0.0274f
C3400 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02762f
C3401 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C3402 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.03425f
C3403 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.15202f
C3404 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.SM 0.00168f
C3405 XA.XIR[11].XIC[0].icell.SM VPWR 0.00158f
C3406 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04031f
C3407 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00214f
C3408 XA.XIR[12].XIC[12].icell.PUM VPWR 0.00937f
C3409 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3410 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C3411 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.SM 0.00168f
C3412 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C3413 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PUM 0.00465f
C3414 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C3415 XA.XIR[7].XIC[6].icell.PDM VPWR 0.00799f
C3416 XThR.Tn[10] XA.XIR[11].XIC[8].icell.SM 0.00121f
C3417 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.SM 0.0039f
C3418 XA.XIR[9].XIC[4].icell.Ien Vbias 0.21098f
C3419 XThR.Tn[1] XA.XIR[2].XIC[9].icell.Ien 0.00338f
C3420 XA.XIR[15].XIC[4].icell.PDM VPWR 0.0114f
C3421 XA.XIR[4].XIC[3].icell.PUM VPWR 0.00937f
C3422 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C3423 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C3424 XThR.XTB6.Y XThR.Tn[6] 0.00639f
C3425 XA.XIR[6].XIC[13].icell.PDM VPWR 0.00799f
C3426 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PUM 0.00465f
C3427 XThC.Tn[13] XThR.Tn[6] 0.2874f
C3428 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.03425f
C3429 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C3430 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C3431 XA.XIR[6].XIC[1].icell.PDM Iout 0.00117f
C3432 XA.XIR[14].XIC[10].icell.PDM VPWR 0.00799f
C3433 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.15202f
C3434 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C3435 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02762f
C3436 XA.XIR[15].XIC[13].icell.SM VPWR 0.00158f
C3437 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.Ien 0.00584f
C3438 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.SM 0.0039f
C3439 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.SM 0.0039f
C3440 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C3441 XA.XIR[1].XIC[3].icell.PDM Vbias 0.04261f
C3442 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C3443 XA.XIR[5].XIC[8].icell.PDM Iout 0.00117f
C3444 XA.XIR[3].XIC[7].icell.PUM Vbias 0.0031f
C3445 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PUM 0.00465f
C3446 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01432f
C3447 XA.XIR[6].XIC[10].icell.SM Vbias 0.00701f
C3448 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00584f
C3449 XThR.XTB7.B a_n1049_6405# 0.00268f
C3450 XA.XIR[9].XIC[2].icell.PDM VPWR 0.00799f
C3451 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[1].icell.SM 0.0039f
C3452 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C3453 XA.XIR[13].XIC[2].icell.PDM Iout 0.00117f
C3454 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PUM 0.00465f
C3455 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Iout 0.00347f
C3456 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PUM 0.00465f
C3457 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00214f
C3458 XA.XIR[4].XIC[3].icell.PDM Vbias 0.04261f
C3459 XA.XIR[5].XIC[13].icell.Ien Vbias 0.21098f
C3460 XThR.Tn[3] Iout 1.16236f
C3461 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.03425f
C3462 XThC.Tn[5] XThR.Tn[7] 0.28739f
C3463 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C3464 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3465 XA.XIR[12].XIC[13].icell.Ien VPWR 0.1903f
C3466 XA.XIR[12].XIC[7].icell.PDM Iout 0.00117f
C3467 XA.XIR[9].XIC[6].icell.PUM VPWR 0.00937f
C3468 XThC.XTB3.Y Vbias 0.01225f
C3469 XThC.XTB7.B XThC.Tn[3] 0.00532f
C3470 XA.XIR[3].XIC[11].icell.PDM Vbias 0.04261f
C3471 XThC.XTB4.Y a_8739_9569# 0.00813f
C3472 XA.XIR[8].XIC[13].icell.PDM Vbias 0.04261f
C3473 XA.XIR[4].XIC_dummy_right.icell.PUM Vbias 0.00223f
C3474 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02762f
C3475 XA.XIR[14].XIC[4].icell.SM Vbias 0.00701f
C3476 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00214f
C3477 XThC.XTB7.Y XThC.Tn[7] 0.0835f
C3478 XThC.Tn[2] Vbias 2.61718f
C3479 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.SM 0.00168f
C3480 XThR.XTB4.Y XThR.Tn[12] 0.00209f
C3481 XA.XIR[13].XIC[6].icell.SM Vbias 0.00701f
C3482 XThC.XTB6.Y XThC.Tn[11] 0.02513f
C3483 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04031f
C3484 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C3485 XA.XIR[8].XIC[10].icell.PUM Vbias 0.0031f
C3486 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.SM 0.0039f
C3487 XA.XIR[11].XIC_15.icell.PDM Vbias 0.04401f
C3488 XA.XIR[3].XIC[7].icell.SM VPWR 0.00158f
C3489 XA.XIR[11].XIC_15.icell.Ien Vbias 0.21234f
C3490 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.0353f
C3491 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Ien 0.00584f
C3492 XA.XIR[1].XIC[7].icell.PDM VPWR 0.00799f
C3493 XA.XIR[12].XIC[8].icell.Ien Vbias 0.21098f
C3494 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C3495 XThR.Tn[14] XA.XIR[15].XIC[13].icell.Ien 0.00338f
C3496 XA.XIR[6].XIC[12].icell.Ien VPWR 0.1903f
C3497 XThC.Tn[9] XThR.Tn[1] 0.28739f
C3498 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.SM 0.00168f
C3499 XThR.XTB5.Y a_n997_1579# 0.00133f
C3500 XA.XIR[10].XIC[12].icell.SM Iout 0.00388f
C3501 XThR.Tn[10] XThR.Tn[12] 0.00142f
C3502 XA.XIR[15].XIC_15.icell.Ien Iout 0.0681f
C3503 XA.XIR[6].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3504 XA.XIR[3].XIC[3].icell.SM Iout 0.00388f
C3505 XThR.Tn[9] XA.XIR[10].XIC[12].icell.SM 0.00121f
C3506 XA.XIR[6].XIC[8].icell.Ien Iout 0.06417f
C3507 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01577f
C3508 XA.XIR[4].XIC[7].icell.PDM VPWR 0.00799f
C3509 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C3510 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7] 0.00341f
C3511 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.SM 0.00168f
C3512 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.SM 0.0039f
C3513 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04031f
C3514 XThC.Tn[9] XThR.Tn[12] 0.28739f
C3515 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.SM 0.0039f
C3516 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07214f
C3517 XA.XIR[1].XIC[2].icell.SM VPWR 0.00158f
C3518 XA.XIR[14].XIC[6].icell.Ien VPWR 0.19084f
C3519 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00584f
C3520 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13] 0.00341f
C3521 XA.XIR[14].XIC[10].icell.Ien Vbias 0.21098f
C3522 XA.XIR[12].XIC[14].icell.SM VPWR 0.00207f
C3523 XA.XIR[8].XIC[5].icell.PDM Iout 0.00117f
C3524 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.03425f
C3525 XA.XIR[4].XIC[12].icell.SM Iout 0.00388f
C3526 XA.XIR[0].XIC[12].icell.PUM Vbias 0.0031f
C3527 XA.XIR[3].XIC[3].icell.PDM Iout 0.00117f
C3528 XThR.XTBN.Y a_n1049_5317# 0.07731f
C3529 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04031f
C3530 XA.XIR[13].XIC[8].icell.Ien VPWR 0.1903f
C3531 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00584f
C3532 XA.XIR[14].XIC[2].icell.Ien Iout 0.06417f
C3533 XThC.Tn[4] XThR.Tn[3] 0.28739f
C3534 XA.XIR[8].XIC[10].icell.SM VPWR 0.00158f
C3535 XThR.Tn[4] XThR.XTB6.Y 0.00264f
C3536 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.03546f
C3537 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C3538 XA.XIR[2].XIC[9].icell.PDM Iout 0.00117f
C3539 XA.XIR[12].XIC[10].icell.PUM VPWR 0.00937f
C3540 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00584f
C3541 XA.XIR[13].XIC[4].icell.Ien Iout 0.06417f
C3542 XThC.Tn[13] XThR.Tn[4] 0.2874f
C3543 XA.XIR[8].XIC[6].icell.SM Iout 0.00388f
C3544 XThR.Tn[8] XA.XIR[9].XIC[6].icell.SM 0.00121f
C3545 XThR.XTB3.Y XThR.Tn[5] 0.00381f
C3546 XThR.Tn[0] XA.XIR[0].XIC[6].icell.PDM 0.00341f
C3547 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.03023f
C3548 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C3549 XA.XIR[2].XIC[13].icell.SM Vbias 0.00701f
C3550 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C3551 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.03425f
C3552 XA.XIR[7].XIC_15.icell.PUM Vbias 0.0031f
C3553 XThR.Tn[14] XA.XIR[15].XIC[14].icell.SM 0.00121f
C3554 XThC.XTB4.Y XThC.Tn[11] 0.30582f
C3555 XThR.Tn[4] XA.XIR[5].XIC[8].icell.Ien 0.00338f
C3556 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.SM 0.00168f
C3557 XThC.Tn[8] XThR.Tn[10] 0.28739f
C3558 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PUM 0.00186f
C3559 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C3560 XA.XIR[11].XIC[7].icell.Ien Iout 0.06417f
C3561 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C3562 XThR.Tn[1] XA.XIR[1].XIC[4].icell.PDM 0.00341f
C3563 XA.XIR[9].XIC[1].icell.PUM VPWR 0.00937f
C3564 XThC.Tn[0] XThR.Tn[5] 0.28743f
C3565 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C3566 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04031f
C3567 XThC.Tn[7] XThR.Tn[0] 0.2882f
C3568 XA.XIR[5].XIC_15.icell.SM Iout 0.0047f
C3569 XThR.Tn[3] XA.XIR[4].XIC[8].icell.Ien 0.00338f
C3570 XA.XIR[10].XIC[9].icell.Ien Iout 0.06417f
C3571 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C3572 XA.XIR[4].XIC[1].icell.Ien Vbias 0.21098f
C3573 XA.XIR[15].XIC[11].icell.SM VPWR 0.00158f
C3574 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00584f
C3575 XThC.Tn[8] XThC.Tn[9] 0.05322f
C3576 XA.XIR[0].XIC[12].icell.SM VPWR 0.00158f
C3577 XThR.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.00338f
C3578 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5] 0.00341f
C3579 XThR.XTB4.Y a_n1049_5317# 0.00463f
C3580 XA.XIR[3].XIC[0].icell.PUM VPWR 0.00937f
C3581 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00214f
C3582 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.SM 0.0039f
C3583 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C3584 XA.XIR[13].XIC[2].icell.PUM Vbias 0.0031f
C3585 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PUM 0.00465f
C3586 XThC.XTB7.A a_6243_9615# 0.02018f
C3587 XA.XIR[0].XIC[8].icell.SM Iout 0.00367f
C3588 XThC.Tn[12] XThC.Tn[14] 0.03994f
C3589 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3590 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.03425f
C3591 XThR.Tn[2] XA.XIR[2].XIC[1].icell.PDM 0.00341f
C3592 XThR.Tn[10] XA.XIR[11].XIC[13].icell.SM 0.00121f
C3593 XThR.Tn[13] XA.XIR[14].XIC[3].icell.SM 0.00121f
C3594 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04031f
C3595 XA.XIR[2].XIC_15.icell.Ien VPWR 0.25566f
C3596 XA.XIR[12].XIC[11].icell.Ien VPWR 0.1903f
C3597 XThC.XTB1.Y Vbias 0.01234f
C3598 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Iout 0.00347f
C3599 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C3600 a_n1319_5611# VPWR 0.00674f
C3601 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.SM 0.0039f
C3602 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6] 0.00341f
C3603 XA.XIR[2].XIC[11].icell.Ien Iout 0.06417f
C3604 XA.XIR[15].XIC[3].icell.Ien Vbias 0.17899f
C3605 XA.XIR[7].XIC[11].icell.SM Iout 0.00388f
C3606 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.03425f
C3607 XA.XIR[5].XIC[3].icell.SM Vbias 0.00701f
C3608 XThR.Tn[0] XA.XIR[1].XIC[6].icell.SM 0.00121f
C3609 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.15202f
C3610 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02762f
C3611 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.SM 0.00168f
C3612 XA.XIR[14].XIC[0].icell.SM VPWR 0.00158f
C3613 XThR.Tn[12] XA.XIR[13].XIC[7].icell.Ien 0.00338f
C3614 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C3615 XA.XIR[1].XIC[13].icell.Ien Iout 0.06417f
C3616 XA.XIR[4].XIC[6].icell.Ien Vbias 0.21098f
C3617 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PDM 0.00172f
C3618 XThR.Tn[7] XA.XIR[8].XIC[12].icell.SM 0.00121f
C3619 XThR.Tn[14] XA.XIR[15].XIC[11].icell.Ien 0.00338f
C3620 XA.XIR[10].XIC[1].icell.PDM VPWR 0.00799f
C3621 XA.XIR[10].XIC[10].icell.SM Iout 0.00388f
C3622 XA.XIR[15].XIC[14].icell.PUM VPWR 0.00937f
C3623 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.SM 0.0039f
C3624 XThR.Tn[9] XA.XIR[10].XIC[10].icell.SM 0.00121f
C3625 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.SM 0.0039f
C3626 XThR.Tn[5] XA.XIR[6].XIC[8].icell.SM 0.00121f
C3627 Vbias bias[2] 0.06133f
C3628 XA.XIR[3].XIC[0].icell.SM Iout 0.00388f
C3629 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.03425f
C3630 XThR.Tn[12] a_n997_1803# 0.18719f
C3631 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.PUM 0.00121f
C3632 XThR.XTBN.Y a_n1049_6405# 0.07602f
C3633 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.SM 0.00168f
C3634 XA.XIR[6].XIC[2].icell.SM VPWR 0.00158f
C3635 XA.XIR[12].XIC[0].icell.Ien Iout 0.06411f
C3636 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.SM 0.0039f
C3637 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC[0].icell.Ien 0.00214f
C3638 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.15202f
C3639 XThC.Tn[6] XThR.Tn[2] 0.28739f
C3640 XA.XIR[9].XIC[13].icell.PDM Vbias 0.04261f
C3641 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02762f
C3642 a_n1049_6699# XThR.XTB5.Y 0.0021f
C3643 XA.XIR[7].XIC[0].icell.Ien Vbias 0.20951f
C3644 XA.XIR[0].XIC[5].icell.PDM Vbias 0.04275f
C3645 XA.XIR[15].XIC[5].icell.PUM VPWR 0.00937f
C3646 XA.XIR[5].XIC[5].icell.Ien VPWR 0.1903f
C3647 XThR.Tn[11] Iout 1.16235f
C3648 XThR.Tn[9] XThR.Tn[11] 0.00252f
C3649 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3650 XA.XIR[1].XIC[2].icell.PUM Vbias 0.0031f
C3651 XA.XIR[9].XIC[9].icell.Ien Vbias 0.21098f
C3652 XA.XIR[10].XIC[3].icell.PUM Vbias 0.0031f
C3653 XA.XIR[4].XIC[8].icell.PUM VPWR 0.00937f
C3654 XA.XIR[7].XIC[9].icell.PDM Iout 0.00117f
C3655 XThR.Tn[1] XA.XIR[2].XIC[14].icell.Ien 0.00338f
C3656 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.SM 0.0039f
C3657 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[9].icell.Ien 0.00214f
C3658 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C3659 XA.XIR[15].XIC[7].icell.PDM Iout 0.00117f
C3660 XA.XIR[0].XIC[2].icell.Ien Vbias 0.2113f
C3661 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PUM 0.00102f
C3662 XA.XIR[11].XIC[14].icell.PDM Vbias 0.04261f
C3663 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.03425f
C3664 XA.XIR[3].XIC[12].icell.PUM Vbias 0.0031f
C3665 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02762f
C3666 XThR.XTB4.Y a_n1049_6405# 0.01546f
C3667 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00584f
C3668 XThR.Tn[5] VPWR 6.61445f
C3669 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00584f
C3670 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.03425f
C3671 XA.XIR[2].XIC[0].icell.SM VPWR 0.00158f
C3672 XA.XIR[14].XIC_15.icell.PDM Vbias 0.04401f
C3673 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01093f
C3674 XA.XIR[7].XIC[2].icell.PUM VPWR 0.00937f
C3675 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.15235f
C3676 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.Ien 0.00584f
C3677 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C3678 XA.XIR[11].XIC[1].icell.SM VPWR 0.00158f
C3679 XA.XIR[2].XIC[5].icell.PUM Vbias 0.0031f
C3680 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C3681 XA.XIR[15].XIC[9].icell.SM VPWR 0.00158f
C3682 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C3683 XA.XIR[9].XIC[5].icell.PDM Iout 0.00117f
C3684 XA.XIR[7].XIC[5].icell.Ien Vbias 0.21098f
C3685 XA.XIR[14].XIC_15.icell.Ien Vbias 0.21234f
C3686 XThR.XTBN.Y XA.XIR[7].XIC_dummy_left.icell.Ien 0.00158f
C3687 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.SM 0.00168f
C3688 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.03425f
C3689 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02762f
C3690 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9] 0.00341f
C3691 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.SM 0.0039f
C3692 XThC.Tn[2] XThR.Tn[6] 0.28739f
C3693 XThR.Tn[12] XThR.Tn[13] 0.06297f
C3694 XA.XIR[13].XIC[12].icell.SM Iout 0.00388f
C3695 XA.XIR[9].XIC[11].icell.PUM VPWR 0.00937f
C3696 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C3697 XA.XIR[1].XIC[7].icell.PUM Vbias 0.0031f
C3698 XA.XIR[10].XIC[3].icell.SM VPWR 0.00158f
C3699 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC_15.icell.Ien 0.00214f
C3700 XA.XIR[9].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.SM 0.0039f
C3701 XThC.XTB6.A a_5949_10571# 0.00467f
C3702 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04031f
C3703 XA.XIR[0].XIC[4].icell.PUM VPWR 0.00882f
C3704 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[4].icell.Ien 0.00214f
C3705 XThR.Tn[10] XA.XIR[11].XIC[11].icell.SM 0.00121f
C3706 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C3707 XThC.Tn[4] XThR.Tn[11] 0.28739f
C3708 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.SM 0.0039f
C3709 XA.XIR[8].XIC_15.icell.PUM Vbias 0.0031f
C3710 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04031f
C3711 XA.XIR[3].XIC[12].icell.SM VPWR 0.00158f
C3712 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00214f
C3713 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10] 0.00341f
C3714 XA.XIR[3].XIC[8].icell.SM Iout 0.00388f
C3715 XA.XIR[1].XIC[10].icell.PDM Iout 0.00117f
C3716 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.SM 0.00168f
C3717 XA.XIR[0].XIC[6].icell.Ien XA.XIR[0].XIC[6].icell.SM 0.0039f
C3718 XA.XIR[6].XIC[13].icell.Ien Iout 0.06417f
C3719 XA.XIR[2].XIC[5].icell.SM VPWR 0.00158f
C3720 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PUM 0.00465f
C3721 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02762f
C3722 XA.XIR[10].XIC[14].icell.Ien Iout 0.06417f
C3723 XA.XIR[7].XIC[7].icell.PUM VPWR 0.00937f
C3724 XThR.Tn[9] XA.XIR[10].XIC[14].icell.Ien 0.00338f
C3725 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[12].icell.Ien 0.00214f
C3726 XA.XIR[4].XIC[10].icell.PDM Iout 0.00117f
C3727 XA.XIR[1].XIC[7].icell.SM VPWR 0.00158f
C3728 XA.XIR[2].XIC[1].icell.SM Iout 0.00388f
C3729 XA.XIR[9].XIC_15.icell.SM VPWR 0.00275f
C3730 XA.XIR[5].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.SM 0.0039f
C3731 XThC.XTB5.Y XThC.Tn[5] 0.01095f
C3732 XA.XIR[15].XIC[12].icell.PUM VPWR 0.00937f
C3733 XThC.Tn[0] XA.XIR[11].XIC_dummy_left.icell.Iout 0.00109f
C3734 a_10915_9569# XThC.Tn[14] 0.20278f
C3735 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.SM 0.00168f
C3736 XThC.Tn[8] XThR.Tn[13] 0.28739f
C3737 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38996f
C3738 a_2979_9615# Vbias 0.00736f
C3739 XA.XIR[1].XIC[3].icell.SM Iout 0.00388f
C3740 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.SM 0.00168f
C3741 XA.XIR[14].XIC[7].icell.Ien Iout 0.06417f
C3742 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0404f
C3743 XA.XIR[10].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.SM 0.0039f
C3744 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.Ien 0.00584f
C3745 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.04498f
C3746 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[10].icell.Ien 0.00214f
C3747 XThR.Tn[6] XA.XIR[7].XIC_15.icell.PUM 0.00186f
C3748 XThC.Tn[7] XThR.Tn[1] 0.2877f
C3749 XA.XIR[13].XIC[9].icell.Ien Iout 0.06417f
C3750 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C3751 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.15202f
C3752 XA.XIR[5].XIC[3].icell.PDM Vbias 0.04261f
C3753 XA.XIR[8].XIC[11].icell.SM Iout 0.00388f
C3754 XThC.Tn[11] Iout 0.84142f
C3755 XThR.Tn[8] XA.XIR[9].XIC[11].icell.SM 0.00121f
C3756 XThC.Tn[11] XThR.Tn[9] 0.28739f
C3757 XA.XIR[6].XIC[2].icell.PUM Vbias 0.0031f
C3758 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C3759 XThR.Tn[2] XA.XIR[3].XIC[6].icell.Ien 0.00338f
C3760 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Iout 0.00347f
C3761 XThR.Tn[4] XA.XIR[4].XIC[3].icell.PDM 0.00341f
C3762 XThC.XTB2.Y data[1] 0.017f
C3763 XThR.Tn[4] XA.XIR[5].XIC[13].icell.Ien 0.00338f
C3764 XA.XIR[7].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.SM 0.0039f
C3765 XThC.Tn[7] XThR.Tn[12] 0.28739f
C3766 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02762f
C3767 XA.XIR[12].XIC[2].icell.PDM Vbias 0.04261f
C3768 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02762f
C3769 XThR.Tn[3] XA.XIR[3].XIC[4].icell.PDM 0.00341f
C3770 XThR.Tn[3] XA.XIR[4].XIC[13].icell.Ien 0.00338f
C3771 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04052f
C3772 a_5155_9615# VPWR 0.7051f
C3773 XA.XIR[11].XIC[8].icell.PDM Vbias 0.04261f
C3774 XThR.Tn[1] XA.XIR[2].XIC[4].icell.SM 0.00121f
C3775 XA.XIR[6].XIC[0].icell.PDM VPWR 0.00799f
C3776 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02762f
C3777 XThC.Tn[2] XThR.Tn[4] 0.28739f
C3778 XThC.XTBN.Y XThC.Tn[5] 0.60785f
C3779 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.SM 0.00168f
C3780 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04031f
C3781 XA.XIR[15].XIC[13].icell.Ien VPWR 0.32895f
C3782 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00584f
C3783 XA.XIR[0].XIC[13].icell.SM Iout 0.00367f
C3784 XA.XIR[5].XIC[7].icell.PDM VPWR 0.00799f
C3785 XA.XIR[3].XIC[2].icell.Ien Vbias 0.21098f
C3786 XThR.Tn[13] XA.XIR[14].XIC[8].icell.SM 0.00121f
C3787 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[14].icell.Ien 0.00214f
C3788 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.SM 0.0039f
C3789 XA.XIR[13].XIC[1].icell.PDM VPWR 0.00799f
C3790 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.03425f
C3791 XA.XIR[14].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.SM 0.0039f
C3792 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C3793 XA.XIR[13].XIC[10].icell.SM Iout 0.00388f
C3794 XA.XIR[6].XIC[7].icell.PUM Vbias 0.0031f
C3795 a_8963_9569# XA.XIR[0].XIC[10].icell.PDM 0.0029f
C3796 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C3797 XThC.Tn[6] XThR.Tn[10] 0.28739f
C3798 XThR.XTB7.B XThR.XTB7.A 0.35833f
C3799 XThC.XTB5.Y a_10051_9569# 0.00133f
C3800 XA.XIR[15].XIC[8].icell.Ien Vbias 0.17899f
C3801 XThC.XTBN.A data[3] 0.07741f
C3802 XA.XIR[12].XIC[6].icell.PDM VPWR 0.00799f
C3803 XA.XIR[2].XIC_dummy_right.icell.SM VPWR 0.00123f
C3804 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02762f
C3805 XThR.Tn[0] XA.XIR[1].XIC[11].icell.SM 0.00121f
C3806 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[11].icell.Ien 0.00214f
C3807 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.SM 0.00168f
C3808 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PUM 0.00465f
C3809 XA.XIR[5].XIC[8].icell.SM Vbias 0.00701f
C3810 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.SM 0.00168f
C3811 XA.XIR[5].XIC[1].icell.Ien Iout 0.06417f
C3812 XThR.Tn[10] XA.XIR[11].XIC[9].icell.SM 0.00121f
C3813 XThC.XTB7.A data[0] 0.86893f
C3814 XThC.Tn[7] XThC.Tn[8] 0.07597f
C3815 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC[0].icell.Ien 0.00214f
C3816 XA.XIR[4].XIC[11].icell.Ien Vbias 0.21098f
C3817 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.SM 0.00168f
C3818 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00584f
C3819 XA.XIR[8].XIC[0].icell.PDM Vbias 0.04207f
C3820 XThR.Tn[14] Iout 1.16234f
C3821 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PUM 0.00465f
C3822 XA.XIR[11].XIC[0].icell.PDM Iout 0.00117f
C3823 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Ien 0.00549f
C3824 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.03425f
C3825 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C3826 XA.XIR[11].XIC[13].icell.PDM Vbias 0.04261f
C3827 XA.XIR[2].XIC[4].icell.PDM Vbias 0.04261f
C3828 a_4861_9615# XThC.Tn[5] 0.00208f
C3829 XA.XIR[8].XIC[2].icell.PUM VPWR 0.00937f
C3830 XA.XIR[13].XIC[3].icell.PUM Vbias 0.0031f
C3831 XThR.Tn[5] XA.XIR[6].XIC[13].icell.SM 0.00121f
C3832 XThR.Tn[6] XA.XIR[7].XIC[0].icell.Ien 0.00338f
C3833 XA.XIR[8].XIC[5].icell.Ien Vbias 0.21098f
C3834 XA.XIR[10].XIC[4].icell.PDM Iout 0.00117f
C3835 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04031f
C3836 XA.XIR[15].XIC[14].icell.SM VPWR 0.00207f
C3837 XA.XIR[3].XIC[4].icell.PUM VPWR 0.00937f
C3838 XA.XIR[10].XIC[12].icell.Ien Iout 0.06417f
C3839 XThR.Tn[9] XA.XIR[10].XIC[12].icell.Ien 0.00338f
C3840 XA.XIR[6].XIC[7].icell.SM VPWR 0.00158f
C3841 XA.XIR[12].XIC[3].icell.SM Vbias 0.00701f
C3842 XThC.XTB6.Y VPWR 1.03148f
C3843 XA.XIR[14].XIC[14].icell.PDM Vbias 0.04261f
C3844 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00584f
C3845 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C3846 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PUM 0.00429f
C3847 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.SM 0.00168f
C3848 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C3849 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.1106f
C3850 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00214f
C3851 XA.XIR[15].XIC[10].icell.PUM VPWR 0.00937f
C3852 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02762f
C3853 XA.XIR[5].XIC[10].icell.Ien VPWR 0.1903f
C3854 XA.XIR[11].XIC[6].icell.PUM Vbias 0.0031f
C3855 XA.XIR[6].XIC[3].icell.SM Iout 0.00388f
C3856 XThC.XTBN.Y a_10051_9569# 0.23006f
C3857 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C3858 XThR.XTB7.A XThR.Tn[2] 0.12549f
C3859 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C3860 XA.XIR[9].XIC[14].icell.Ien Vbias 0.21098f
C3861 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.15202f
C3862 XA.XIR[4].XIC[13].icell.PUM VPWR 0.00937f
C3863 XThR.Tn[14] XA.XIR[15].XIC[0].icell.Ien 0.00377f
C3864 XA.XIR[10].XIC[8].icell.PUM Vbias 0.0031f
C3865 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02762f
C3866 XA.XIR[5].XIC[6].icell.Ien Iout 0.06417f
C3867 XA.XIR[3].XIC[2].icell.PDM VPWR 0.00799f
C3868 XA.XIR[8].XIC[4].icell.PDM VPWR 0.00799f
C3869 XA.XIR[14].XIC[1].icell.SM VPWR 0.00158f
C3870 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.15202f
C3871 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02762f
C3872 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.15202f
C3873 XA.XIR[2].XIC[8].icell.PDM VPWR 0.00799f
C3874 XA.XIR[0].XIC[7].icell.Ien Vbias 0.21134f
C3875 XA.XIR[13].XIC[3].icell.SM VPWR 0.00158f
C3876 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[6].icell.Ien 0.00214f
C3877 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00214f
C3878 XA.XIR[8].XIC[7].icell.PUM VPWR 0.00937f
C3879 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.02762f
C3880 XThR.Tn[6] XA.XIR[7].XIC[5].icell.Ien 0.00338f
C3881 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C3882 XA.XIR[12].XIC[5].icell.Ien VPWR 0.1903f
C3883 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12] 0.00341f
C3884 XA.XIR[11].XIC_dummy_right.icell.Ien Vbias 0.00288f
C3885 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.Ien 0.00584f
C3886 XThC.Tn[4] XThR.Tn[14] 0.28739f
C3887 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.03425f
C3888 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C3889 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.SM 0.00168f
C3890 XA.XIR[2].XIC[10].icell.PUM Vbias 0.0031f
C3891 XA.XIR[11].XIC[6].icell.SM VPWR 0.00158f
C3892 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04031f
C3893 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.SM 0.00168f
C3894 XA.XIR[7].XIC[10].icell.Ien Vbias 0.21098f
C3895 XThR.Tn[4] XA.XIR[5].XIC[3].icell.SM 0.00121f
C3896 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.0353f
C3897 XA.XIR[14].XIC_dummy_left.icell.Ien Vbias 0.00329f
C3898 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02762f
C3899 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3900 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Iout 0.00347f
C3901 XA.XIR[11].XIC[2].icell.SM Iout 0.00388f
C3902 XA.XIR[15].XIC[11].icell.Ien VPWR 0.32895f
C3903 XA.XIR[1].XIC[12].icell.PUM Vbias 0.0031f
C3904 XA.XIR[10].XIC[8].icell.SM VPWR 0.00158f
C3905 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.Ien 0.00584f
C3906 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.15202f
C3907 XThR.Tn[14] XA.XIR[15].XIC[5].icell.Ien 0.00338f
C3908 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02762f
C3909 XA.XIR[13].XIC[14].icell.Ien Iout 0.06417f
C3910 XThR.Tn[3] XA.XIR[4].XIC[3].icell.SM 0.00121f
C3911 XThC.XTB4.Y VPWR 0.91479f
C3912 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C3913 XA.XIR[10].XIC[4].icell.SM Iout 0.00388f
C3914 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.03431f
C3915 XThR.Tn[9] XA.XIR[10].XIC[4].icell.SM 0.00121f
C3916 XThC.XTB2.Y XThC.Tn[0] 0.00125f
C3917 XA.XIR[0].XIC[9].icell.PUM VPWR 0.00877f
C3918 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00214f
C3919 XA.XIR[12].XIC_15.icell.SM VPWR 0.00275f
C3920 XThC.Tn[0] XA.XIR[14].XIC_dummy_left.icell.Iout 0.00109f
C3921 XA.XIR[8].XIC[0].icell.Ien Vbias 0.20951f
C3922 XThR.Tn[10] XA.XIR[11].XIC[13].icell.Ien 0.00338f
C3923 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04031f
C3924 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[4].icell.Ien 0.00214f
C3925 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C3926 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C3927 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C3928 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04031f
C3929 XA.XIR[3].XIC[13].icell.SM Iout 0.00388f
C3930 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.SM 0.0039f
C3931 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8] 0.00341f
C3932 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.04591f
C3933 XA.XIR[7].XIC[12].icell.PUM VPWR 0.00937f
C3934 XThC.XTB5.A data[0] 0.14415f
C3935 XThR.XTB5.A VPWR 0.83125f
C3936 XA.XIR[2].XIC[10].icell.SM VPWR 0.00158f
C3937 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[2].icell.Ien 0.00214f
C3938 XA.XIR[2].XIC[6].icell.SM Iout 0.00388f
C3939 XA.XIR[1].XIC[12].icell.SM VPWR 0.00158f
C3940 XA.XIR[7].XIC[4].icell.PDM Vbias 0.04261f
C3941 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C3942 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.04036f
C3943 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04031f
C3944 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.SM 0.00168f
C3945 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PUM 0.00465f
C3946 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PUM 0.00465f
C3947 XThR.Tn[12] XA.XIR[13].XIC[2].icell.SM 0.00121f
C3948 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3949 XA.XIR[1].XIC[8].icell.SM Iout 0.00388f
C3950 XA.XIR[15].XIC[2].icell.PDM Vbias 0.04261f
C3951 XA.XIR[4].XIC[1].icell.SM Vbias 0.00701f
C3952 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00584f
C3953 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.SM 0.00168f
C3954 XA.XIR[6].XIC[11].icell.PDM Vbias 0.04261f
C3955 XThR.Tn[13] XA.XIR[14].XIC[13].icell.SM 0.00121f
C3956 XA.XIR[10].XIC[10].icell.Ien Iout 0.06417f
C3957 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C3958 XThR.Tn[9] XA.XIR[10].XIC[10].icell.Ien 0.00338f
C3959 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02762f
C3960 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.15202f
C3961 XA.XIR[3].XIC[1].icell.PUM VPWR 0.00937f
C3962 XThC.XTB7.B a_5155_9615# 0.00268f
C3963 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00584f
C3964 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Ien 0.00584f
C3965 XA.XIR[14].XIC[8].icell.PDM Vbias 0.04261f
C3966 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02762f
C3967 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PUM 0.00465f
C3968 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.15202f
C3969 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02762f
C3970 XThR.Tn[11] XA.XIR[12].XIC[5].icell.SM 0.00121f
C3971 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C3972 XThC.XTB6.Y a_9827_9569# 0.00871f
C3973 XThR.Tn[10] XA.XIR[11].XIC[14].icell.SM 0.00121f
C3974 XThR.Tn[2] XA.XIR[3].XIC[11].icell.Ien 0.00338f
C3975 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C3976 XA.XIR[11].XIC[2].icell.PUM VPWR 0.00937f
C3977 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.SM 0.00168f
C3978 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3979 XA.XIR[9].XIC[0].icell.PDM Vbias 0.04207f
C3980 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04031f
C3981 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PDM 0.00172f
C3982 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.03425f
C3983 XA.XIR[7].XIC[8].icell.PDM VPWR 0.00799f
C3984 XThR.XTB3.Y XThR.Tn[9] 0.00285f
C3985 XA.XIR[9].XIC[1].icell.Ien VPWR 0.1903f
C3986 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.15202f
C3987 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.SM 0.0039f
C3988 a_4067_9615# XThC.Tn[1] 0.00584f
C3989 XThC.Tn[6] XThR.Tn[13] 0.28739f
C3990 XA.XIR[9].XIC[4].icell.SM Vbias 0.00701f
C3991 XThR.Tn[1] XA.XIR[2].XIC[9].icell.SM 0.00121f
C3992 XA.XIR[15].XIC[6].icell.PDM VPWR 0.0114f
C3993 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07214f
C3994 XA.XIR[4].XIC[3].icell.Ien VPWR 0.1903f
C3995 VPWR data[5] 0.4402f
C3996 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.SM 0.00168f
C3997 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.03023f
C3998 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.PUM 0.00179f
C3999 XA.XIR[11].XIC[12].icell.PDM Vbias 0.04261f
C4000 XA.XIR[3].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.SM 0.0039f
C4001 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C4002 XThC.Tn[0] Iout 0.82545f
C4003 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C4004 XThC.Tn[0] XThR.Tn[9] 0.28741f
C4005 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C4006 XA.XIR[6].XIC[3].icell.PDM Iout 0.00117f
C4007 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.SM 0.00168f
C4008 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[14].icell.Ien 0.00214f
C4009 XA.XIR[3].XIC[7].icell.Ien Vbias 0.21098f
C4010 XA.XIR[14].XIC[0].icell.PDM Iout 0.00117f
C4011 XThR.XTB5.Y a_n997_3755# 0.00418f
C4012 XA.XIR[5].XIC[10].icell.PDM Iout 0.00117f
C4013 XA.XIR[1].XIC[5].icell.PDM Vbias 0.04261f
C4014 XThC.Tn[5] XThR.Tn[8] 0.28739f
C4015 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C4016 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C4017 XA.XIR[14].XIC[13].icell.PDM Vbias 0.04261f
C4018 XA.XIR[6].XIC[12].icell.PUM Vbias 0.0031f
C4019 XA.XIR[9].XIC[4].icell.PDM VPWR 0.00799f
C4020 a_7875_9569# VPWR 0.00639f
C4021 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PUM 0.00465f
C4022 XA.XIR[13].XIC[4].icell.PDM Iout 0.00117f
C4023 XA.XIR[13].XIC[12].icell.Ien Iout 0.06417f
C4024 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.SM 0.00168f
C4025 XA.XIR[5].XIC[13].icell.SM Vbias 0.00701f
C4026 XA.XIR[4].XIC[5].icell.PDM Vbias 0.04261f
C4027 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PUM 0.00102f
C4028 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.03425f
C4029 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00214f
C4030 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.03425f
C4031 XThC.XTB2.Y VPWR 0.97668f
C4032 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C4033 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C4034 XA.XIR[12].XIC[9].icell.PDM Iout 0.00117f
C4035 XThR.XTB7.A XThR.Tn[10] 0.00404f
C4036 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.1106f
C4037 XA.XIR[9].XIC[6].icell.Ien VPWR 0.1903f
C4038 XA.XIR[3].XIC[13].icell.PDM Vbias 0.04261f
C4039 XA.XIR[1].XIC[2].icell.Ien Vbias 0.21104f
C4040 XA.XIR[14].XIC[6].icell.PUM Vbias 0.0031f
C4041 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.03023f
C4042 XA.XIR[8].XIC_15.icell.PDM Vbias 0.04401f
C4043 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PUM 0.00429f
C4044 XThR.Tn[10] XA.XIR[11].XIC[11].icell.Ien 0.00338f
C4045 XA.XIR[9].XIC[2].icell.Ien Iout 0.06417f
C4046 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C4047 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.15202f
C4048 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C4049 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[5].icell.Ien 0.00214f
C4050 XA.XIR[13].XIC[8].icell.PUM Vbias 0.0031f
C4051 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02762f
C4052 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04031f
C4053 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PUM 0.00465f
C4054 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00584f
C4055 XA.XIR[8].XIC[10].icell.Ien Vbias 0.21098f
C4056 XThR.XTB5.Y a_n1049_5611# 0.0093f
C4057 XA.XIR[3].XIC[9].icell.PUM VPWR 0.00937f
C4058 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Ien 0.00584f
C4059 XA.XIR[1].XIC[9].icell.PDM VPWR 0.00799f
C4060 XThC.XTB3.Y XThC.Tn[2] 0.1864f
C4061 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02852f
C4062 XA.XIR[12].XIC[8].icell.SM Vbias 0.00701f
C4063 XA.XIR[6].XIC[12].icell.SM VPWR 0.00158f
C4064 XA.XIR[10].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.SM 0.0039f
C4065 XA.XIR[10].XIC[13].icell.SM VPWR 0.00158f
C4066 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C4067 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC_15.icell.Ien 0.00214f
C4068 XThC.Tn[1] XThC.Tn[3] 0.10977f
C4069 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7] 0.00341f
C4070 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02762f
C4071 XA.XIR[7].XIC[2].icell.Ien VPWR 0.1903f
C4072 XA.XIR[5].XIC_15.icell.Ien VPWR 0.25566f
C4073 XA.XIR[6].XIC[8].icell.SM Iout 0.00388f
C4074 XA.XIR[4].XIC[9].icell.PDM VPWR 0.00799f
C4075 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04031f
C4076 XA.XIR[14].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4077 XThR.Tn[13] XA.XIR[14].XIC[11].icell.SM 0.00121f
C4078 XThC.Tn[6] XThC.Tn[7] 0.1602f
C4079 XA.XIR[5].XIC[11].icell.Ien Iout 0.06417f
C4080 XA.XIR[8].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.SM 0.0039f
C4081 XA.XIR[1].XIC[4].icell.PUM VPWR 0.00937f
C4082 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C4083 XA.XIR[14].XIC[6].icell.SM VPWR 0.00158f
C4084 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13] 0.00341f
C4085 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[14].icell.Ien 0.00214f
C4086 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PUM 0.00465f
C4087 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C4088 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07214f
C4089 XA.XIR[3].XIC[5].icell.PDM Iout 0.00117f
C4090 XA.XIR[0].XIC[12].icell.Ien Vbias 0.2113f
C4091 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4092 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02762f
C4093 XA.XIR[14].XIC[2].icell.SM Iout 0.00388f
C4094 XA.XIR[8].XIC[7].icell.PDM Iout 0.00117f
C4095 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04031f
C4096 XA.XIR[13].XIC[8].icell.SM VPWR 0.00158f
C4097 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C4098 XA.XIR[8].XIC[12].icell.PUM VPWR 0.00937f
C4099 XThR.Tn[6] XA.XIR[7].XIC[10].icell.Ien 0.00338f
C4100 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C4101 XA.XIR[2].XIC[11].icell.PDM Iout 0.00117f
C4102 XA.XIR[13].XIC[4].icell.SM Iout 0.00388f
C4103 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00584f
C4104 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00214f
C4105 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.SM 0.0039f
C4106 XThC.Tn[8] XThR.Tn[7] 0.28739f
C4107 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C4108 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PUM 0.00465f
C4109 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.SM 0.00168f
C4110 XThR.Tn[0] XA.XIR[0].XIC[8].icell.PDM 0.00341f
C4111 XA.XIR[12].XIC[6].icell.Ien Iout 0.06417f
C4112 XA.XIR[2].XIC_15.icell.PUM Vbias 0.0031f
C4113 XThR.Tn[2] XA.XIR[3].XIC[1].icell.SM 0.00121f
C4114 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00214f
C4115 XA.XIR[7].XIC_15.icell.Ien Vbias 0.21234f
C4116 XThR.Tn[4] XA.XIR[5].XIC[8].icell.SM 0.00121f
C4117 XA.XIR[5].XIC[0].icell.Ien Vbias 0.20951f
C4118 XThR.Tn[1] XA.XIR[1].XIC[6].icell.PDM 0.00341f
C4119 XA.XIR[10].XIC_15.icell.Ien Iout 0.0642f
C4120 XA.XIR[13].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.SM 0.0039f
C4121 VPWR Iout 54.1536f
C4122 XA.XIR[11].XIC[7].icell.SM Iout 0.00388f
C4123 XThR.Tn[9] VPWR 7.55029f
C4124 XThC.XTB7.Y XThC.Tn[10] 0.07406f
C4125 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04031f
C4126 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.SM 0.00168f
C4127 XThR.Tn[9] XA.XIR[10].XIC_15.icell.Ien 0.00117f
C4128 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C4129 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04031f
C4130 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C4131 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C4132 XThR.Tn[3] XA.XIR[4].XIC[8].icell.SM 0.00121f
C4133 XA.XIR[14].XIC[1].icell.PUM Vbias 0.0031f
C4134 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.15202f
C4135 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[13].icell.Ien 0.00214f
C4136 XA.XIR[0].XIC[14].icell.PUM VPWR 0.00877f
C4137 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[9].icell.Ien 0.00214f
C4138 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.15202f
C4139 XThC.Tn[14] Vbias 2.45788f
C4140 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.SM 0.00168f
C4141 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5] 0.00341f
C4142 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.15202f
C4143 XThR.XTBN.Y XA.XIR[11].XIC_dummy_left.icell.Ien 0.0016f
C4144 XA.XIR[12].XIC[0].icell.PUM VPWR 0.00937f
C4145 XThR.Tn[2] XA.XIR[2].XIC[3].icell.PDM 0.00341f
C4146 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C4147 XA.XIR[13].XIC[10].icell.Ien Iout 0.06417f
C4148 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04031f
C4149 XA.XIR[0].XIC[11].icell.Ien XA.XIR[0].XIC[11].icell.SM 0.0039f
C4150 XA.XIR[6].XIC[2].icell.Ien Vbias 0.21098f
C4151 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.15202f
C4152 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04052f
C4153 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.Ien 0.00584f
C4154 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PUM 0.00465f
C4155 XA.XIR[15].XIC[0].icell.Ien VPWR 0.32895f
C4156 XA.XIR[5].XIC[0].icell.SM VPWR 0.00158f
C4157 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6] 0.00341f
C4158 XA.XIR[15].XIC[3].icell.SM Vbias 0.00701f
C4159 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C4160 XA.XIR[2].XIC[11].icell.SM Iout 0.00388f
C4161 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.03425f
C4162 XA.XIR[5].XIC[5].icell.PUM Vbias 0.0031f
C4163 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C4164 XA.XIR[5].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.SM 0.0039f
C4165 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C4166 XA.XIR[14].XIC[2].icell.PUM VPWR 0.00937f
C4167 XThR.Tn[12] XA.XIR[13].XIC[7].icell.SM 0.00121f
C4168 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.SM 0.00168f
C4169 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C4170 XA.XIR[1].XIC[13].icell.SM Iout 0.00388f
C4171 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02762f
C4172 XA.XIR[4].XIC[6].icell.SM Vbias 0.00701f
C4173 XA.XIR[11].XIC[11].icell.PDM Vbias 0.04261f
C4174 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.15202f
C4175 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00214f
C4176 XA.XIR[10].XIC[3].icell.PDM VPWR 0.00799f
C4177 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C4178 XThC.Tn[4] VPWR 5.88871f
C4179 XA.XIR[10].XIC[11].icell.SM VPWR 0.00158f
C4180 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PUM 0.00465f
C4181 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.15202f
C4182 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C4183 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C4184 XA.XIR[14].XIC[12].icell.PDM Vbias 0.04261f
C4185 XA.XIR[6].XIC[4].icell.PUM VPWR 0.00937f
C4186 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PUM 0.00465f
C4187 XA.XIR[12].XIC[0].icell.SM Iout 0.00388f
C4188 XThR.Tn[13] XA.XIR[14].XIC[9].icell.SM 0.00121f
C4189 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C4190 XA.XIR[9].XIC_15.icell.PDM Vbias 0.04401f
C4191 XA.XIR[7].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.SM 0.0039f
C4192 XThC.Tn[10] XThR.Tn[0] 0.28747f
C4193 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Ien 0.00309f
C4194 XThC.Tn[12] XThR.Tn[5] 0.28739f
C4195 XA.XIR[7].XIC[0].icell.SM Vbias 0.00675f
C4196 XA.XIR[0].XIC[7].icell.PDM Vbias 0.04278f
C4197 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Iout 0.00347f
C4198 XA.XIR[15].XIC[5].icell.Ien VPWR 0.32895f
C4199 XA.XIR[5].XIC[5].icell.SM VPWR 0.00158f
C4200 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.15202f
C4201 XThR.XTB7.B XThR.Tn[10] 0.06102f
C4202 XThC.XTB7.B a_7875_9569# 0.01174f
C4203 XThR.Tn[1] XA.XIR[2].XIC[14].icell.SM 0.00121f
C4204 XA.XIR[9].XIC[9].icell.SM Vbias 0.00701f
C4205 XA.XIR[7].XIC[11].icell.PDM Iout 0.00117f
C4206 XA.XIR[10].XIC[3].icell.Ien Vbias 0.21098f
C4207 XA.XIR[4].XIC[8].icell.Ien VPWR 0.1903f
C4208 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C4209 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C4210 XA.XIR[5].XIC[1].icell.SM Iout 0.00388f
C4211 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.SM 0.00168f
C4212 XA.XIR[1].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.SM 0.0039f
C4213 XA.XIR[12].XIC[13].icell.SM Vbias 0.00701f
C4214 XA.XIR[4].XIC[4].icell.Ien Iout 0.06417f
C4215 XA.XIR[15].XIC[9].icell.PDM Iout 0.00117f
C4216 XA.XIR[0].XIC[2].icell.SM Vbias 0.00716f
C4217 a_8963_9569# XThC.Tn[11] 0.19413f
C4218 XA.XIR[12].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.SM 0.0039f
C4219 XA.XIR[8].XIC[2].icell.Ien VPWR 0.1903f
C4220 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PUM 0.00465f
C4221 XA.XIR[3].XIC[12].icell.Ien Vbias 0.21098f
C4222 XA.XIR[10].XIC[14].icell.PUM VPWR 0.00937f
C4223 XA.XIR[15].XIC_15.icell.SM VPWR 0.00275f
C4224 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C4225 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PUM 0.00465f
C4226 XThR.Tn[2] XThR.XTB4.Y 0.0021f
C4227 XA.XIR[2].XIC[2].icell.PUM VPWR 0.00937f
C4228 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.15202f
C4229 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.SM 0.00168f
C4230 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.03591f
C4231 XA.XIR[0].XIC[11].icell.PDM VPWR 0.00774f
C4232 XA.XIR[11].XIC[3].icell.PUM VPWR 0.00937f
C4233 XA.XIR[2].XIC[5].icell.Ien Vbias 0.21098f
C4234 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[12].icell.Ien 0.00214f
C4235 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[3].icell.Ien 0.00214f
C4236 XA.XIR[9].XIC[7].icell.PDM Iout 0.00117f
C4237 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C4238 XA.XIR[7].XIC[5].icell.SM Vbias 0.00701f
C4239 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9] 0.00341f
C4240 XA.XIR[13].XIC[13].icell.SM VPWR 0.00158f
C4241 XA.XIR[9].XIC[11].icell.Ien VPWR 0.1903f
C4242 XThR.XTBN.Y XA.XIR[0].XIC_dummy_left.icell.Iout 0.00137f
C4243 XA.XIR[1].XIC[7].icell.Ien Vbias 0.21104f
C4244 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11] 0.00341f
C4245 XA.XIR[10].XIC[5].icell.PUM VPWR 0.00937f
C4246 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.Ien 0.00584f
C4247 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C4248 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C4249 XA.XIR[12].XIC[14].icell.PDM VPWR 0.00809f
C4250 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02762f
C4251 XA.XIR[9].XIC[7].icell.Ien Iout 0.06417f
C4252 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PUM 0.00465f
C4253 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C4254 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.15202f
C4255 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04031f
C4256 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18982f
C4257 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.SM 0.00168f
C4258 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PUM 0.00465f
C4259 XA.XIR[8].XIC_15.icell.Ien Vbias 0.21234f
C4260 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04031f
C4261 XThC.Tn[9] XThR.Tn[2] 0.28739f
C4262 XA.XIR[3].XIC[14].icell.PUM VPWR 0.00937f
C4263 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02762f
C4264 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C4265 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07555f
C4266 XA.XIR[1].XIC[12].icell.PDM Iout 0.00117f
C4267 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C4268 XA.XIR[2].XIC[7].icell.PUM VPWR 0.00937f
C4269 XA.XIR[6].XIC[13].icell.SM Iout 0.00388f
C4270 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.03425f
C4271 XA.XIR[7].XIC[7].icell.Ien VPWR 0.1903f
C4272 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04031f
C4273 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C4274 XA.XIR[5].XIC_dummy_right.icell.SM VPWR 0.00123f
C4275 XA.XIR[4].XIC[12].icell.PDM Iout 0.00117f
C4276 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C4277 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01444f
C4278 XA.XIR[7].XIC[3].icell.Ien Iout 0.06417f
C4279 XA.XIR[1].XIC[9].icell.PUM VPWR 0.00937f
C4280 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C4281 XThR.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.00338f
C4282 XA.XIR[10].XIC[9].icell.SM VPWR 0.00158f
C4283 XThC.XTB7.B Iout 0.00967f
C4284 XA.XIR[13].XIC_15.icell.Ien Iout 0.0642f
C4285 a_4067_9615# Vbias 0.00573f
C4286 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02762f
C4287 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C4288 XA.XIR[14].XIC[7].icell.SM Iout 0.00388f
C4289 XThC.XTB7.A XThC.Tn[5] 0.02758f
C4290 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PUM 0.00465f
C4291 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38919f
C4292 XThR.Tn[7] XA.XIR[8].XIC[4].icell.Ien 0.00338f
C4293 XThR.Tn[6] XA.XIR[7].XIC_15.icell.Ien 0.00117f
C4294 XA.XIR[5].XIC[5].icell.PDM Vbias 0.04261f
C4295 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.SM 0.00168f
C4296 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.Ien 0.00256f
C4297 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C4298 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C4299 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.04036f
C4300 data[1] data[0] 0.64735f
C4301 XThR.Tn[2] XA.XIR[3].XIC[6].icell.SM 0.00121f
C4302 XA.XIR[15].XIC_dummy_left.icell.SM VPWR 0.00269f
C4303 XThR.XTB7.B a_n997_1803# 0.00228f
C4304 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.15202f
C4305 XThR.Tn[4] XA.XIR[5].XIC[13].icell.SM 0.00121f
C4306 XThR.Tn[4] XA.XIR[4].XIC[5].icell.PDM 0.00341f
C4307 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.03425f
C4308 XThC.Tn[14] XThR.Tn[6] 0.28745f
C4309 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.15202f
C4310 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PUM 0.00465f
C4311 XA.XIR[12].XIC[4].icell.PDM Vbias 0.04261f
C4312 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.Ien 0.00584f
C4313 XA.XIR[12].XIC[11].icell.SM Vbias 0.00701f
C4314 XThR.Tn[10] XA.XIR[11].XIC[5].icell.Ien 0.00338f
C4315 XThR.Tn[3] XA.XIR[4].XIC[13].icell.SM 0.00121f
C4316 XThR.Tn[3] XA.XIR[3].XIC[6].icell.PDM 0.00341f
C4317 a_6243_9615# VPWR 0.70553f
C4318 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PUM 0.00465f
C4319 XA.XIR[11].XIC[10].icell.PDM Vbias 0.04261f
C4320 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.15202f
C4321 XA.XIR[6].XIC[2].icell.PDM VPWR 0.00799f
C4322 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.03425f
C4323 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04031f
C4324 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.15202f
C4325 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C4326 XA.XIR[10].XIC[12].icell.PUM VPWR 0.00937f
C4327 XThR.Tn[13] XA.XIR[14].XIC[14].icell.SM 0.00121f
C4328 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C4329 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.15202f
C4330 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02762f
C4331 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.SM 0.00168f
C4332 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C4333 XA.XIR[5].XIC[9].icell.PDM VPWR 0.00799f
C4334 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C4335 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02762f
C4336 XA.XIR[8].XIC[0].icell.SM Vbias 0.00675f
C4337 XA.XIR[6].XIC[8].icell.Ien XA.XIR[6].XIC[9].icell.Ien 0.00214f
C4338 XA.XIR[14].XIC[11].icell.PDM Vbias 0.04261f
C4339 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C4340 XThC.Tn[6] XThR.Tn[7] 0.28739f
C4341 XA.XIR[10].XIC[10].icell.Ien XA.XIR[10].XIC[11].icell.Ien 0.00214f
C4342 XA.XIR[3].XIC[2].icell.SM Vbias 0.00701f
C4343 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Iout 0.00347f
C4344 XA.XIR[13].XIC[3].icell.PDM VPWR 0.00799f
C4345 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.SM 0.00168f
C4346 XThC.XTB7.B XThC.Tn[4] 0.00356f
C4347 XA.XIR[6].XIC[7].icell.Ien Vbias 0.21098f
C4348 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.15202f
C4349 XA.XIR[13].XIC[11].icell.SM VPWR 0.00158f
C4350 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PUM 0.00268f
C4351 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.0284f
C4352 a_9827_9569# XA.XIR[0].XIC[11].icell.PDM 0.00136f
C4353 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C4354 XThC.XTB5.Y XThC.Tn[8] 0.01728f
C4355 XThC.XTB7.Y a_7651_9569# 0.00477f
C4356 XA.XIR[12].XIC[8].icell.PDM VPWR 0.00799f
C4357 XA.XIR[15].XIC[8].icell.SM Vbias 0.00701f
C4358 XThR.XTB1.Y data[4] 0.06453f
C4359 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02762f
C4360 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C4361 XThR.XTB5.Y a_n997_2667# 0.00427f
C4362 XThC.Tn[3] Vbias 2.45762f
C4363 XA.XIR[5].XIC[10].icell.PUM Vbias 0.0031f
C4364 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C4365 XThC.XTB6.A a_5155_10571# 0.00306f
C4366 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C4367 XA.XIR[15].XIC[1].icell.Ien Iout 0.06807f
C4368 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C4369 XThC.XTB6.Y XThC.Tn[12] 0.02863f
C4370 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.0353f
C4371 XA.XIR[9].XIC[1].icell.SM VPWR 0.00158f
C4372 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.03425f
C4373 XA.XIR[13].XIC[13].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00214f
C4374 XA.XIR[3].XIC[0].icell.PDM Vbias 0.04207f
C4375 XA.XIR[4].XIC[11].icell.SM Vbias 0.00701f
C4376 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00584f
C4377 XA.XIR[12].XIC[14].icell.PUM Vbias 0.0031f
C4378 XA.XIR[8].XIC[2].icell.PDM Vbias 0.04261f
C4379 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C4380 XThR.XTB7.B XThR.Tn[13] 0.00276f
C4381 XThC.Tn[10] XThR.Tn[1] 0.28739f
C4382 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.03425f
C4383 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02762f
C4384 XA.XIR[11].XIC[2].icell.PDM Iout 0.00117f
C4385 a_5949_9615# XThC.Tn[5] 0.27124f
C4386 XA.XIR[10].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.SM 0.0039f
C4387 XA.XIR[2].XIC[6].icell.PDM Vbias 0.04261f
C4388 XA.XIR[13].XIC[3].icell.Ien Vbias 0.21098f
C4389 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PUM 0.00186f
C4390 XThR.Tn[6] XA.XIR[7].XIC[0].icell.SM 0.00121f
C4391 XA.XIR[14].XIC[2].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00214f
C4392 XA.XIR[10].XIC[6].icell.PDM Iout 0.00117f
C4393 XA.XIR[8].XIC[5].icell.SM Vbias 0.00701f
C4394 XA.XIR[10].XIC[13].icell.Ien VPWR 0.1903f
C4395 XA.XIR[3].XIC[4].icell.Ien VPWR 0.1903f
C4396 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04031f
C4397 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C4398 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02762f
C4399 XThC.Tn[10] XThR.Tn[12] 0.28739f
C4400 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C4401 XA.XIR[12].XIC[5].icell.PUM Vbias 0.0031f
C4402 XA.XIR[6].XIC[9].icell.PUM VPWR 0.00937f
C4403 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C4404 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C4405 XThR.Tn[13] XA.XIR[14].XIC[11].icell.Ien 0.00338f
C4406 XA.XIR[11].XIC[6].icell.Ien Vbias 0.21098f
C4407 XA.XIR[15].XIC[0].icell.Ien XA.XIR[15].XIC[1].icell.Ien 0.00214f
C4408 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7] 0.00341f
C4409 XThR.Tn[4] XA.XIR[5].XIC[0].icell.Ien 0.00338f
C4410 XA.XIR[5].XIC[10].icell.SM VPWR 0.00158f
C4411 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.15202f
C4412 XA.XIR[9].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4413 XA.XIR[13].XIC[14].icell.PUM VPWR 0.00937f
C4414 XThC.XTBN.Y XThC.Tn[8] 0.50311f
C4415 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PUM 0.00465f
C4416 XThC.Tn[5] XThR.Tn[3] 0.28739f
C4417 XA.XIR[13].XIC[4].icell.Ien XA.XIR[13].XIC[5].icell.Ien 0.00214f
C4418 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C4419 XA.XIR[15].XIC[6].icell.Ien Iout 0.06807f
C4420 XA.XIR[5].XIC[6].icell.SM Iout 0.00388f
C4421 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C4422 XA.XIR[9].XIC[14].icell.SM Vbias 0.00701f
C4423 XA.XIR[3].XIC[4].icell.PDM VPWR 0.00799f
C4424 XThR.Tn[14] XA.XIR[15].XIC[0].icell.SM 0.00128f
C4425 XThC.XTB1.Y a_2979_9615# 0.21263f
C4426 XA.XIR[4].XIC[13].icell.Ien VPWR 0.1903f
C4427 XA.XIR[8].XIC[6].icell.PDM VPWR 0.00799f
C4428 XA.XIR[12].XIC[13].icell.PDM VPWR 0.00799f
C4429 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.04563f
C4430 XA.XIR[10].XIC[8].icell.Ien Vbias 0.21098f
C4431 XThC.Tn[14] XThR.Tn[4] 0.28745f
C4432 XA.XIR[14].XIC[3].icell.PUM VPWR 0.00937f
C4433 XA.XIR[3].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.SM 0.0039f
C4434 XA.XIR[4].XIC[9].icell.Ien Iout 0.06417f
C4435 XA.XIR[13].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.SM 0.0039f
C4436 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.04498f
C4437 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C4438 XA.XIR[0].XIC[7].icell.SM Vbias 0.00716f
C4439 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.SM 0.00168f
C4440 XA.XIR[2].XIC[10].icell.PDM VPWR 0.00799f
C4441 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04037f
C4442 XA.XIR[13].XIC[5].icell.PUM VPWR 0.00937f
C4443 XThC.Tn[0] XA.XIR[9].XIC_dummy_left.icell.Iout 0.00109f
C4444 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02762f
C4445 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C4446 XA.XIR[8].XIC[7].icell.Ien VPWR 0.1903f
C4447 XA.XIR[0].XIC[0].icell.Ien Iout 0.06382f
C4448 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01149f
C4449 XThC.XTB4.Y XThC.Tn[12] 0.00209f
C4450 XThR.Tn[6] XA.XIR[7].XIC[5].icell.SM 0.00121f
C4451 XThC.Tn[9] XThR.Tn[10] 0.28739f
C4452 XThC.Tn[1] XThR.Tn[5] 0.28739f
C4453 XA.XIR[6].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.SM 0.0039f
C4454 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C4455 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.SM 0.00168f
C4456 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12] 0.00341f
C4457 XA.XIR[12].XIC[5].icell.SM VPWR 0.00158f
C4458 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.15202f
C4459 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02762f
C4460 XA.XIR[8].XIC[3].icell.Ien Iout 0.06417f
C4461 XThR.Tn[8] XA.XIR[9].XIC[3].icell.Ien 0.00338f
C4462 XA.XIR[12].XIC[9].icell.SM Vbias 0.00701f
C4463 XA.XIR[10].XIC[14].icell.SM VPWR 0.00207f
C4464 XA.XIR[12].XIC[1].icell.SM Iout 0.00388f
C4465 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C4466 XA.XIR[11].XIC[8].icell.PUM VPWR 0.00937f
C4467 XA.XIR[2].XIC[10].icell.Ien Vbias 0.21098f
C4468 XThC.Tn[8] XThC.Tn[10] 0.00465f
C4469 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C4470 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04031f
C4471 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02762f
C4472 XA.XIR[7].XIC[10].icell.SM Vbias 0.00701f
C4473 XA.XIR[11].XIC[7].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00214f
C4474 XA.XIR[2].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.SM 0.0039f
C4475 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C4476 XA.XIR[10].XIC[10].icell.PUM VPWR 0.00937f
C4477 XThC.Tn[13] XThC.Tn[14] 0.38789f
C4478 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PUM 0.00465f
C4479 XA.XIR[1].XIC[12].icell.Ien Vbias 0.21104f
C4480 XThR.Tn[14] XA.XIR[15].XIC[5].icell.SM 0.00121f
C4481 XA.XIR[9].XIC[12].icell.Ien Iout 0.06417f
C4482 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.SM 0.00168f
C4483 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.15202f
C4484 XA.XIR[0].XIC[9].icell.Ien VPWR 0.19115f
C4485 XA.XIR[1].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.SM 0.0039f
C4486 XA.XIR[11].XIC_15.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Ien 0.00214f
C4487 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C4488 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02762f
C4489 XA.XIR[13].XIC[9].icell.SM VPWR 0.00158f
C4490 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C4491 XA.XIR[0].XIC[5].icell.Ien Iout 0.06389f
C4492 XThR.Tn[5] XA.XIR[6].XIC[0].icell.Ien 0.00338f
C4493 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04031f
C4494 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04031f
C4495 XThR.XTBN.Y a_n997_1803# 0.22873f
C4496 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04031f
C4497 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8] 0.00341f
C4498 XA.XIR[2].XIC[12].icell.PUM VPWR 0.00937f
C4499 XA.XIR[13].XIC[12].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00214f
C4500 XA.XIR[7].XIC[12].icell.Ien VPWR 0.1903f
C4501 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00584f
C4502 XA.XIR[11].XIC[0].icell.SM Vbias 0.00675f
C4503 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C4504 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.15202f
C4505 XA.XIR[7].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4506 XA.XIR[12].XIC[12].icell.PUM Vbias 0.0031f
C4507 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.Ien 0.00584f
C4508 XA.XIR[15].XIC[5].icell.Ien XA.XIR[15].XIC[6].icell.Ien 0.00214f
C4509 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PUM 0.00465f
C4510 XThR.Tn[0] XA.XIR[1].XIC[3].icell.Ien 0.00338f
C4511 XA.XIR[1].XIC[14].icell.PUM VPWR 0.00937f
C4512 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04031f
C4513 XA.XIR[8].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.SM 0.0039f
C4514 XA.XIR[7].XIC[6].icell.PDM Vbias 0.04261f
C4515 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.03425f
C4516 XA.XIR[7].XIC[8].icell.Ien Iout 0.06417f
C4517 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C4518 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.03425f
C4519 XA.XIR[6].XIC[13].icell.PDM Vbias 0.04261f
C4520 XA.XIR[10].XIC[11].icell.Ien VPWR 0.1903f
C4521 XA.XIR[15].XIC[4].icell.PDM Vbias 0.04261f
C4522 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C4523 XThR.XTB6.A a_n997_3755# 0.00149f
C4524 XA.XIR[4].XIC[3].icell.PUM Vbias 0.0031f
C4525 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C4526 XThR.Tn[7] XA.XIR[8].XIC[9].icell.Ien 0.00338f
C4527 XA.XIR[3].XIC[1].icell.Ien VPWR 0.1903f
C4528 XThC.XTB7.B a_6243_9615# 0.01743f
C4529 XA.XIR[9].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.SM 0.0039f
C4530 XThC.Tn[7] XThR.Tn[2] 0.28746f
C4531 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PUM 0.00465f
C4532 XA.XIR[14].XIC[10].icell.PDM Vbias 0.04261f
C4533 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00256f
C4534 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02762f
C4535 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PUM 0.00465f
C4536 XA.XIR[4].XIC[8].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00214f
C4537 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C4538 XA.XIR[15].XIC[13].icell.SM Vbias 0.00701f
C4539 XThR.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.00338f
C4540 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C4541 XA.XIR[12].XIC[1].icell.PUM VPWR 0.00937f
C4542 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PUM 0.00465f
C4543 XA.XIR[13].XIC[12].icell.PUM VPWR 0.00937f
C4544 XThR.Tn[2] XA.XIR[3].XIC[11].icell.SM 0.00121f
C4545 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02762f
C4546 XA.XIR[2].XIC[11].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00214f
C4547 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.SM 0.00168f
C4548 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.15202f
C4549 XA.XIR[9].XIC[2].icell.PDM Vbias 0.04261f
C4550 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.04036f
C4551 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02799f
C4552 XA.XIR[7].XIC[10].icell.PDM VPWR 0.00799f
C4553 XThR.Tn[0] XThR.XTB2.Y 0.00125f
C4554 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C4555 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.1106f
C4556 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02762f
C4557 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C4558 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PUM 0.00465f
C4559 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C4560 XA.XIR[9].XIC[6].icell.PUM Vbias 0.0031f
C4561 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C4562 XA.XIR[12].XIC[13].icell.Ien Vbias 0.21098f
C4563 XA.XIR[8].XIC[2].icell.Ien XA.XIR[8].XIC[3].icell.Ien 0.00214f
C4564 XA.XIR[10].XIC[0].icell.Ien Iout 0.06411f
C4565 XA.XIR[4].XIC[3].icell.SM VPWR 0.00158f
C4566 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.15202f
C4567 XA.XIR[1].XIC[13].icell.Ien XA.XIR[1].XIC[14].icell.Ien 0.00214f
C4568 XA.XIR[15].XIC[8].icell.PDM VPWR 0.0114f
C4569 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C4570 XThR.Tn[9] XA.XIR[10].XIC[0].icell.Ien 0.0037f
C4571 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C4572 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.SM 0.00168f
C4573 XA.XIR[6].XIC[5].icell.PDM Iout 0.00117f
C4574 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.15202f
C4575 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.15202f
C4576 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C4577 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C4578 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C4579 XThC.Tn[3] XThR.Tn[6] 0.28739f
C4580 XA.XIR[3].XIC[7].icell.SM Vbias 0.00701f
C4581 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02762f
C4582 XA.XIR[5].XIC[12].icell.PDM Iout 0.00117f
C4583 XA.XIR[14].XIC[2].icell.PDM Iout 0.00117f
C4584 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C4585 XA.XIR[1].XIC[7].icell.PDM Vbias 0.04261f
C4586 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.15202f
C4587 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.Ien 0.00584f
C4588 XA.XIR[6].XIC[12].icell.Ien Vbias 0.21098f
C4589 a_8963_9569# VPWR 0.0033f
C4590 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00584f
C4591 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.Ien 0.00584f
C4592 XA.XIR[9].XIC[6].icell.PDM VPWR 0.00799f
C4593 XThR.XTB7.A XThR.Tn[7] 0.00182f
C4594 VPWR data[0] 0.52929f
C4595 XThR.XTB7.A a_n997_2891# 0.00342f
C4596 XA.XIR[13].XIC[6].icell.PDM Iout 0.00117f
C4597 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.SM 0.00168f
C4598 XA.XIR[13].XIC[13].icell.Ien VPWR 0.1903f
C4599 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C4600 XA.XIR[4].XIC[7].icell.PDM Vbias 0.04261f
C4601 XA.XIR[5].XIC_15.icell.PUM Vbias 0.0031f
C4602 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02762f
C4603 XA.XIR[5].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.SM 0.0039f
C4604 XThC.Tn[5] XThR.Tn[11] 0.28739f
C4605 XA.XIR[12].XIC[12].icell.PDM VPWR 0.00799f
C4606 XA.XIR[9].XIC[6].icell.SM VPWR 0.00158f
C4607 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C4608 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C4609 XA.XIR[1].XIC[2].icell.SM Vbias 0.00704f
C4610 XA.XIR[3].XIC_15.icell.PDM Vbias 0.04401f
C4611 XA.XIR[14].XIC[6].icell.Ien Vbias 0.21098f
C4612 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.03579f
C4613 XA.XIR[12].XIC[0].icell.Ien XA.XIR[12].XIC[1].icell.Ien 0.00214f
C4614 XA.XIR[9].XIC[2].icell.SM Iout 0.00388f
C4615 XA.XIR[9].XIC[11].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00214f
C4616 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.PDM 0.00587f
C4617 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.SM 0.00168f
C4618 XA.XIR[12].XIC[14].icell.SM Vbias 0.00701f
C4619 XA.XIR[15].XIC[13].icell.PDM VPWR 0.0114f
C4620 XA.XIR[13].XIC[8].icell.Ien Vbias 0.21098f
C4621 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04031f
C4622 XA.XIR[13].XIC[11].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00214f
C4623 XA.XIR[8].XIC[10].icell.SM Vbias 0.00701f
C4624 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.03425f
C4625 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00584f
C4626 XThR.Tn[11] XA.XIR[12].XIC[1].icell.Ien 0.00338f
C4627 XA.XIR[3].XIC[9].icell.Ien VPWR 0.1903f
C4628 XA.XIR[4].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.SM 0.0039f
C4629 XA.XIR[1].XIC[11].icell.PDM VPWR 0.00799f
C4630 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.03433f
C4631 XA.XIR[12].XIC[10].icell.PUM Vbias 0.0031f
C4632 XA.XIR[6].XIC[14].icell.PUM VPWR 0.00937f
C4633 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PUM 0.00465f
C4634 XThC.XTB5.Y XThC.Tn[6] 0.00352f
C4635 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14] 0.00341f
C4636 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.0353f
C4637 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.Ien 0.00584f
C4638 XA.XIR[3].XIC[5].icell.Ien Iout 0.06417f
C4639 XA.XIR[0].XIC[4].icell.Ien XA.XIR[0].XIC[5].icell.Ien 0.00214f
C4640 XThC.Tn[9] XThR.Tn[13] 0.28739f
C4641 XA.XIR[2].XIC[2].icell.Ien VPWR 0.1903f
C4642 XA.XIR[7].XIC[2].icell.SM VPWR 0.00158f
C4643 XA.XIR[4].XIC[11].icell.PDM VPWR 0.00799f
C4644 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C4645 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04031f
C4646 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C4647 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02762f
C4648 XA.XIR[9].XIC[1].icell.PUM Vbias 0.0031f
C4649 XA.XIR[5].XIC[11].icell.SM Iout 0.00388f
C4650 XA.XIR[13].XIC[14].icell.SM VPWR 0.00207f
C4651 XA.XIR[1].XIC[4].icell.Ien VPWR 0.1903f
C4652 XA.XIR[14].XIC[8].icell.PUM VPWR 0.00937f
C4653 XThC.Tn[12] Iout 0.84307f
C4654 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.03425f
C4655 XA.XIR[15].XIC[11].icell.SM Vbias 0.00701f
C4656 XThC.Tn[12] XThR.Tn[9] 0.28739f
C4657 XA.XIR[4].XIC[14].icell.Ien Iout 0.06417f
C4658 XA.XIR[3].XIC[7].icell.PDM Iout 0.00117f
C4659 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04031f
C4660 XThC.Tn[8] XThR.Tn[8] 0.28739f
C4661 XA.XIR[8].XIC[9].icell.PDM Iout 0.00117f
C4662 XA.XIR[0].XIC[12].icell.SM Vbias 0.00716f
C4663 XA.XIR[12].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.SM 0.0039f
C4664 XA.XIR[13].XIC[10].icell.PUM VPWR 0.00937f
C4665 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.Ien 0.00584f
C4666 XA.XIR[8].XIC[12].icell.Ien VPWR 0.1903f
C4667 XA.XIR[8].XIC_dummy_right.icell.Ien Vbias 0.00288f
C4668 XA.XIR[2].XIC[13].icell.PDM Iout 0.00117f
C4669 XThR.Tn[6] XA.XIR[7].XIC[10].icell.SM 0.00121f
C4670 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04031f
C4671 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.03425f
C4672 XA.XIR[8].XIC[8].icell.Ien Iout 0.06417f
C4673 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PUM 0.00465f
C4674 XThR.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.00338f
C4675 XA.XIR[12].XIC[6].icell.SM Iout 0.00388f
C4676 XThR.Tn[0] XA.XIR[0].XIC[10].icell.PDM 0.00341f
C4677 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C4678 XA.XIR[2].XIC_15.icell.Ien Vbias 0.21234f
C4679 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C4680 XThC.XTBN.Y XThC.Tn[6] 0.61358f
C4681 XA.XIR[12].XIC[11].icell.Ien Vbias 0.21098f
C4682 XA.XIR[7].XIC[7].icell.Ien XA.XIR[7].XIC[8].icell.Ien 0.00214f
C4683 XThR.XTB7.B a_n997_3979# 0.01152f
C4684 XThC.Tn[3] XThR.Tn[4] 0.28739f
C4685 XA.XIR[10].XIC_15.icell.PDM Iout 0.00133f
C4686 XThR.Tn[1] XA.XIR[1].XIC[8].icell.PDM 0.00341f
C4687 XThR.Tn[9] XA.XIR[10].XIC_15.icell.PDM 0.00172f
C4688 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C4689 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04031f
C4690 XThR.XTBN.Y XA.XIR[8].XIC_dummy_left.icell.Ien 0.00243f
C4691 XA.XIR[14].XIC[0].icell.SM Vbias 0.00675f
C4692 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18971f
C4693 XThC.XTB7.Y a_5949_9615# 0.00153f
C4694 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C4695 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C4696 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5] 0.00341f
C4697 XThC.Tn[7] XThR.Tn[10] 0.28739f
C4698 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.15202f
C4699 XA.XIR[10].XIC[1].icell.PDM Vbias 0.04261f
C4700 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.15202f
C4701 XA.XIR[0].XIC[10].icell.Ien Iout 0.06389f
C4702 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Ien 0.00584f
C4703 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.SM 0.0039f
C4704 XA.XIR[15].XIC[14].icell.PUM Vbias 0.0031f
C4705 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C4706 XThR.Tn[2] XA.XIR[2].XIC[5].icell.PDM 0.00341f
C4707 XA.XIR[13].XIC[11].icell.Ien VPWR 0.1903f
C4708 XA.XIR[6].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.SM 0.0039f
C4709 XThR.Tn[13] XA.XIR[14].XIC[5].icell.Ien 0.00338f
C4710 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04031f
C4711 a_7651_9569# XThC.Tn[8] 0.1927f
C4712 XA.XIR[6].XIC[2].icell.SM Vbias 0.00701f
C4713 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02762f
C4714 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PUM 0.00465f
C4715 XThC.XTB5.A XThC.XTB7.Y 0.00179f
C4716 XA.XIR[15].XIC[0].icell.SM VPWR 0.00158f
C4717 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.15202f
C4718 XA.XIR[5].XIC[2].icell.PUM VPWR 0.00937f
C4719 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6] 0.00341f
C4720 XA.XIR[7].XIC[13].icell.Ien Iout 0.06417f
C4721 XA.XIR[15].XIC[5].icell.PUM Vbias 0.0031f
C4722 XThR.Tn[0] XA.XIR[1].XIC[8].icell.Ien 0.00338f
C4723 XA.XIR[5].XIC[5].icell.Ien Vbias 0.21098f
C4724 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C4725 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.SM 0.00168f
C4726 XA.XIR[11].XIC[1].icell.PDM VPWR 0.00799f
C4727 XA.XIR[13].XIC[10].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00214f
C4728 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C4729 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.03425f
C4730 XA.XIR[4].XIC[8].icell.PUM Vbias 0.0031f
C4731 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Iout 0.00347f
C4732 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02762f
C4733 XThR.Tn[7] XA.XIR[8].XIC[14].icell.Ien 0.00338f
C4734 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PUM 0.00465f
C4735 XThR.Tn[13] a_n997_1803# 0.0021f
C4736 XA.XIR[10].XIC[5].icell.PDM VPWR 0.00799f
C4737 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C4738 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.03425f
C4739 XA.XIR[13].XIC[0].icell.Ien Iout 0.06411f
C4740 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02771f
C4741 XThR.Tn[5] XA.XIR[6].XIC[10].icell.Ien 0.00338f
C4742 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.SM 0.00168f
C4743 XThR.XTB7.B XThR.Tn[7] 0.07415f
C4744 XThR.Tn[5] Vbias 3.74761f
C4745 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.03425f
C4746 XA.XIR[6].XIC[4].icell.Ien VPWR 0.1903f
C4747 XThR.XTB7.B a_n997_2891# 0.0168f
C4748 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02762f
C4749 XA.XIR[7].XIC[2].icell.PUM Vbias 0.0031f
C4750 XA.XIR[2].XIC[0].icell.SM Vbias 0.00675f
C4751 XA.XIR[15].XIC[5].icell.SM VPWR 0.00158f
C4752 XA.XIR[0].XIC[9].icell.PDM Vbias 0.04282f
C4753 XA.XIR[5].XIC[7].icell.PUM VPWR 0.00937f
C4754 XA.XIR[12].XIC[11].icell.PDM VPWR 0.00799f
C4755 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.03425f
C4756 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.Ien 0.00256f
C4757 XA.XIR[11].XIC[1].icell.SM Vbias 0.00701f
C4758 XA.XIR[13].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.SM 0.0039f
C4759 XA.XIR[15].XIC[9].icell.SM Vbias 0.00701f
C4760 XThC.XTB7.B a_8963_9569# 0.02071f
C4761 XThC.XTB7.B data[0] 0.0138f
C4762 XA.XIR[9].XIC[11].icell.PUM Vbias 0.0031f
C4763 XThC.Tn[12] XA.XIR[0].XIC[11].icell.PDM 0.00106f
C4764 XA.XIR[15].XIC[1].icell.SM Iout 0.00388f
C4765 XA.XIR[7].XIC[13].icell.PDM Iout 0.00117f
C4766 XA.XIR[10].XIC[3].icell.SM Vbias 0.00701f
C4767 XA.XIR[4].XIC[8].icell.SM VPWR 0.00158f
C4768 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C4769 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.Ien 0.00584f
C4770 XThC.Tn[5] XThR.Tn[14] 0.28739f
C4771 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.15202f
C4772 XThC.XTB6.A XThC.XTB7.A 0.44014f
C4773 XA.XIR[15].XIC[12].icell.PDM VPWR 0.0114f
C4774 XA.XIR[4].XIC[4].icell.SM Iout 0.00388f
C4775 XA.XIR[0].XIC[4].icell.PUM Vbias 0.0031f
C4776 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C4777 XA.XIR[8].XIC[2].icell.SM VPWR 0.00158f
C4778 XThR.XTB6.A data[4] 0.48493f
C4779 XA.XIR[6].XIC[13].icell.Ien XA.XIR[6].XIC[14].icell.Ien 0.00214f
C4780 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C4781 XThR.Tn[13] XA.XIR[14].XIC[0].icell.Ien 0.0037f
C4782 XA.XIR[3].XIC[12].icell.SM Vbias 0.00701f
C4783 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.Ien 0.00584f
C4784 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C4785 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.03425f
C4786 XA.XIR[0].XIC[13].icell.PDM VPWR 0.00774f
C4787 XThC.XTB2.Y XThC.Tn[1] 0.17879f
C4788 XA.XIR[11].XIC[3].icell.Ien VPWR 0.1903f
C4789 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C4790 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C4791 XA.XIR[7].XIC[7].icell.PUM Vbias 0.0031f
C4792 XA.XIR[11].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.SM 0.0039f
C4793 XA.XIR[2].XIC[5].icell.SM Vbias 0.00701f
C4794 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.SM 0.00168f
C4795 XA.XIR[9].XIC[9].icell.PDM Iout 0.00117f
C4796 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9] 0.00341f
C4797 XA.XIR[9].XIC[11].icell.SM VPWR 0.00158f
C4798 XA.XIR[10].XIC[5].icell.Ien VPWR 0.1903f
C4799 XA.XIR[5].XIC[1].icell.Ien XA.XIR[5].XIC[2].icell.Ien 0.00214f
C4800 XA.XIR[1].XIC[7].icell.SM Vbias 0.00704f
C4801 XA.XIR[9].XIC_15.icell.SM Vbias 0.00701f
C4802 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11] 0.00341f
C4803 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C4804 XA.XIR[15].XIC[12].icell.PUM Vbias 0.0031f
C4805 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.03425f
C4806 XA.XIR[9].XIC[7].icell.SM Iout 0.00388f
C4807 XA.XIR[0].XIC[4].icell.SM VPWR 0.00158f
C4808 XA.XIR[3].XIC_dummy_left.icell.Ien Vbias 0.00329f
C4809 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04031f
C4810 XA.XIR[10].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.SM 0.0039f
C4811 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C4812 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04031f
C4813 XA.XIR[14].XIC[7].icell.Ien XA.XIR[14].XIC[8].icell.Ien 0.00214f
C4814 XA.XIR[3].XIC[14].icell.Ien VPWR 0.19036f
C4815 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02762f
C4816 XThR.XTB2.Y a_n1049_5317# 0.00844f
C4817 XThR.XTBN.Y a_n997_3979# 0.23021f
C4818 XA.XIR[3].XIC[10].icell.Ien Iout 0.06417f
C4819 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.SM 0.00168f
C4820 XA.XIR[1].XIC[14].icell.PDM Iout 0.00117f
C4821 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C4822 XA.XIR[10].XIC_15.icell.SM VPWR 0.00275f
C4823 XA.XIR[2].XIC[7].icell.Ien VPWR 0.1903f
C4824 XA.XIR[10].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.SM 0.0039f
C4825 XA.XIR[10].XIC[14].icell.PDM Iout 0.00117f
C4826 XA.XIR[7].XIC[7].icell.SM VPWR 0.00158f
C4827 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04052f
C4828 XA.XIR[14].XIC_15.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Ien 0.00214f
C4829 XA.XIR[1].XIC[9].icell.Ien VPWR 0.1903f
C4830 XA.XIR[7].XIC[3].icell.SM Iout 0.00388f
C4831 XA.XIR[2].XIC[3].icell.Ien Iout 0.06417f
C4832 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C4833 XA.XIR[15].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.SM 0.0039f
C4834 XA.XIR[4].XIC[14].icell.PDM Iout 0.00117f
C4835 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02762f
C4836 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.15202f
C4837 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.SM 0.00168f
C4838 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C4839 XThR.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.00338f
C4840 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02762f
C4841 a_5155_9615# Vbias 0.00695f
C4842 XA.XIR[13].XIC_15.icell.PDM Iout 0.00133f
C4843 XA.XIR[1].XIC[5].icell.Ien Iout 0.06417f
C4844 XA.XIR[6].XIC[0].icell.PDM Vbias 0.04207f
C4845 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.SM 0.00168f
C4846 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C4847 XThR.Tn[7] XA.XIR[8].XIC[4].icell.SM 0.00121f
C4848 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PUM 0.00465f
C4849 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C4850 XThC.XTB3.Y a_4067_9615# 0.23056f
C4851 XA.XIR[15].XIC[13].icell.Ien Vbias 0.17899f
C4852 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.03425f
C4853 XA.XIR[5].XIC[7].icell.PDM Vbias 0.04261f
C4854 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C4855 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PUM 0.00429f
C4856 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C4857 XA.XIR[4].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.SM 0.0039f
C4858 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PUM 0.00465f
C4859 XThR.Tn[8] XA.XIR[9].XIC[13].icell.Ien 0.00338f
C4860 XThR.Tn[11] XA.XIR[12].XIC[2].icell.Ien 0.00338f
C4861 XA.XIR[8].XIC[13].icell.Ien Iout 0.06417f
C4862 a_4067_9615# XThC.Tn[2] 0.27699f
C4863 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.SM 0.00168f
C4864 XThC.Tn[7] XThR.Tn[13] 0.28739f
C4865 XThR.XTB4.Y a_n997_3979# 0.00497f
C4866 XA.XIR[13].XIC[1].icell.PDM Vbias 0.04261f
C4867 XA.XIR[2].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.SM 0.0039f
C4868 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.04036f
C4869 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02762f
C4870 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.15202f
C4871 XThR.Tn[4] XA.XIR[4].XIC[7].icell.PDM 0.00341f
C4872 XThC.Tn[1] Iout 0.84229f
C4873 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PUM 0.00186f
C4874 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.03425f
C4875 XThC.Tn[1] XThR.Tn[9] 0.28739f
C4876 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PUM 0.00465f
C4877 XA.XIR[12].XIC[6].icell.PDM Vbias 0.04261f
C4878 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PUM 0.00186f
C4879 XThR.Tn[3] XA.XIR[3].XIC[8].icell.PDM 0.00341f
C4880 XThC.XTB5.A XThC.XTB6.A 1.80461f
C4881 XThR.Tn[10] XA.XIR[11].XIC[5].icell.SM 0.00121f
C4882 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C4883 XThR.Tn[1] XA.XIR[2].XIC[6].icell.Ien 0.00338f
C4884 XThC.Tn[6] XThR.Tn[8] 0.28739f
C4885 XA.XIR[1].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.SM 0.0039f
C4886 XA.XIR[6].XIC[4].icell.PDM VPWR 0.00799f
C4887 XThR.XTB7.A a_n1049_6699# 0.02294f
C4888 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04052f
C4889 XA.XIR[3].XIC[4].icell.Ien XA.XIR[3].XIC[5].icell.Ien 0.00214f
C4890 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.15202f
C4891 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.15202f
C4892 XA.XIR[0].XIC_15.icell.Ien Iout 0.06388f
C4893 XThR.XTB5.Y VPWR 1.0269f
C4894 XA.XIR[14].XIC[1].icell.PDM VPWR 0.00799f
C4895 XA.XIR[8].XIC[2].icell.PUM Vbias 0.0031f
C4896 XA.XIR[5].XIC[11].icell.PDM VPWR 0.00799f
C4897 XThR.XTBN.Y XThR.Tn[7] 0.8998f
C4898 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PUM 0.00465f
C4899 XThR.XTBN.Y a_n997_2891# 0.22804f
C4900 XA.XIR[13].XIC[5].icell.PDM VPWR 0.00799f
C4901 XA.XIR[15].XIC[14].icell.SM Vbias 0.00701f
C4902 XA.XIR[3].XIC[4].icell.PUM Vbias 0.0031f
C4903 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02762f
C4904 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C4905 XA.XIR[6].XIC[7].icell.SM Vbias 0.00701f
C4906 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00584f
C4907 XThC.XTB6.Y Vbias 0.01503f
C4908 XA.XIR[7].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.SM 0.0039f
C4909 XA.XIR[6].XIC[0].icell.Ien Iout 0.06411f
C4910 XThC.XTB7.Y a_8739_9569# 0.00474f
C4911 XA.XIR[12].XIC[10].icell.PDM VPWR 0.00799f
C4912 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.Ien 0.00584f
C4913 XA.XIR[15].XIC[10].icell.PUM Vbias 0.0031f
C4914 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02762f
C4915 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.SM 0.00168f
C4916 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.SM 0.00168f
C4917 XThR.Tn[0] XA.XIR[1].XIC[13].icell.Ien 0.00338f
C4918 XA.XIR[5].XIC[10].icell.Ien Vbias 0.21098f
C4919 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.SM 0.00168f
C4920 XThR.XTB2.Y a_n1049_6405# 0.00847f
C4921 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.0353f
C4922 XThR.XTB7.B a_n997_1579# 0.00209f
C4923 XA.XIR[9].XIC[3].icell.PUM VPWR 0.00937f
C4924 XThC.XTB3.Y XThC.Tn[3] 0.01287f
C4925 XA.XIR[8].XIC[4].icell.PDM Vbias 0.04261f
C4926 XA.XIR[3].XIC[2].icell.PDM Vbias 0.04261f
C4927 XA.XIR[4].XIC[13].icell.PUM Vbias 0.0031f
C4928 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.Ien 0.00584f
C4929 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.SM 0.00168f
C4930 XA.XIR[14].XIC[1].icell.SM Vbias 0.00701f
C4931 XA.XIR[15].XIC[11].icell.PDM VPWR 0.0114f
C4932 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PUM 0.00465f
C4933 XA.XIR[11].XIC[4].icell.PDM Iout 0.00117f
C4934 XA.XIR[9].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.SM 0.0039f
C4935 XThR.Tn[5] XThR.Tn[6] 0.06649f
C4936 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00584f
C4937 XThC.Tn[2] XThC.Tn[3] 0.33669f
C4938 XA.XIR[2].XIC[8].icell.PDM Vbias 0.04261f
C4939 XA.XIR[13].XIC[3].icell.SM Vbias 0.00701f
C4940 XA.XIR[4].XIC[13].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00214f
C4941 XThR.Tn[5] XA.XIR[6].XIC_15.icell.Ien 0.00117f
C4942 XA.XIR[8].XIC[7].icell.PUM Vbias 0.0031f
C4943 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.SM 0.00168f
C4944 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C4945 XA.XIR[10].XIC[8].icell.PDM Iout 0.00117f
C4946 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04031f
C4947 XThR.XTB4.Y a_n997_2891# 0.00813f
C4948 XA.XIR[3].XIC[4].icell.SM VPWR 0.00158f
C4949 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C4950 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02762f
C4951 XA.XIR[6].XIC[9].icell.Ien VPWR 0.1903f
C4952 XA.XIR[12].XIC[5].icell.Ien Vbias 0.21098f
C4953 XThC.Tn[0] XA.XIR[3].XIC_dummy_left.icell.Iout 0.00109f
C4954 XA.XIR[11].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.SM 0.0039f
C4955 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.SM 0.00168f
C4956 XA.XIR[0].XIC[2].icell.Ien XA.XIR[0].XIC[2].icell.SM 0.0039f
C4957 XA.XIR[6].XIC[5].icell.Ien Iout 0.06417f
C4958 XA.XIR[5].XIC[12].icell.PUM VPWR 0.00937f
C4959 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7] 0.00341f
C4960 XA.XIR[11].XIC[6].icell.SM Vbias 0.00701f
C4961 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.Ien 0.00584f
C4962 XThR.Tn[10] a_n997_2891# 0.1927f
C4963 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.03425f
C4964 XA.XIR[9].XIC_dummy_right.icell.PUM Vbias 0.00223f
C4965 XA.XIR[15].XIC[6].icell.SM Iout 0.00388f
C4966 XA.XIR[3].XIC[6].icell.PDM VPWR 0.00799f
C4967 XA.XIR[10].XIC[8].icell.SM Vbias 0.00701f
C4968 XThR.Tn[3] XA.XIR[4].XIC[0].icell.Ien 0.00338f
C4969 XA.XIR[8].XIC[7].icell.Ien XA.XIR[8].XIC[8].icell.Ien 0.00214f
C4970 XA.XIR[8].XIC[8].icell.PDM VPWR 0.00799f
C4971 XA.XIR[4].XIC[13].icell.SM VPWR 0.00158f
C4972 XA.XIR[15].XIC[11].icell.Ien Vbias 0.17899f
C4973 XA.XIR[14].XIC[3].icell.Ien VPWR 0.19084f
C4974 XThC.Tn[9] XThR.Tn[7] 0.28739f
C4975 XThC.XTB4.Y Vbias 0.01548f
C4976 XA.XIR[2].XIC[12].icell.PDM VPWR 0.00799f
C4977 XA.XIR[4].XIC[9].icell.SM Iout 0.00388f
C4978 XA.XIR[13].XIC[5].icell.Ien VPWR 0.1903f
C4979 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C4980 XA.XIR[0].XIC[9].icell.PUM Vbias 0.0031f
C4981 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04031f
C4982 XA.XIR[8].XIC[7].icell.SM VPWR 0.00158f
C4983 XThR.XTB1.Y VPWR 1.13148f
C4984 XA.XIR[12].XIC_15.icell.SM Vbias 0.00701f
C4985 XA.XIR[0].XIC[0].icell.SM Iout 0.00367f
C4986 XThC.XTB2.Y a_3523_10575# 0.01006f
C4987 XA.XIR[2].XIC[0].icell.PDM Iout 0.00117f
C4988 XThC.XTB7.Y XThC.Tn[11] 0.07471f
C4989 XA.XIR[12].XIC[7].icell.PUM VPWR 0.00937f
C4990 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.Ien 0.00584f
C4991 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12] 0.00341f
C4992 XA.XIR[8].XIC[3].icell.SM Iout 0.00388f
C4993 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00584f
C4994 XThR.XTB6.Y a_n1319_5611# 0.01283f
C4995 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C4996 XThR.Tn[8] XA.XIR[9].XIC[3].icell.SM 0.00121f
C4997 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C4998 XA.XIR[10].XIC[13].icell.PDM Iout 0.00117f
C4999 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.04036f
C5000 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5001 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PUM 0.00465f
C5002 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02762f
C5003 XA.XIR[11].XIC[8].icell.Ien VPWR 0.1903f
C5004 XA.XIR[2].XIC[10].icell.SM Vbias 0.00701f
C5005 XA.XIR[7].XIC[12].icell.PUM Vbias 0.0031f
C5006 XA.XIR[7].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.SM 0.0039f
C5007 XThR.Tn[4] XA.XIR[5].XIC[5].icell.Ien 0.00338f
C5008 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02762f
C5009 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C5010 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.03425f
C5011 XA.XIR[11].XIC[4].icell.Ien Iout 0.06417f
C5012 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PUM 0.00465f
C5013 XA.XIR[1].XIC[12].icell.SM Vbias 0.00704f
C5014 XThR.Tn[3] XA.XIR[4].XIC[5].icell.Ien 0.00338f
C5015 XA.XIR[13].XIC_15.icell.SM VPWR 0.00275f
C5016 XA.XIR[13].XIC[14].icell.PDM Iout 0.00117f
C5017 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02832f
C5018 XA.XIR[9].XIC[12].icell.SM Iout 0.00388f
C5019 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C5020 XA.XIR[10].XIC[6].icell.Ien Iout 0.06417f
C5021 XA.XIR[0].XIC[9].icell.SM VPWR 0.00158f
C5022 XThR.Tn[9] XA.XIR[10].XIC[6].icell.Ien 0.00338f
C5023 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5] 0.00341f
C5024 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02762f
C5025 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02762f
C5026 XA.XIR[3].XIC[1].icell.PUM Vbias 0.0031f
C5027 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.Ien 0.00584f
C5028 XA.XIR[0].XIC[5].icell.SM Iout 0.00367f
C5029 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04031f
C5030 XThR.Tn[5] XA.XIR[6].XIC[0].icell.SM 0.00121f
C5031 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.Ien 0.00584f
C5032 XA.XIR[3].XIC_15.icell.Ien Iout 0.0642f
C5033 XThR.Tn[4] XThR.Tn[5] 0.07388f
C5034 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8] 0.00341f
C5035 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04031f
C5036 XThC.XTB5.A XThC.Tn[8] 0.00205f
C5037 XThC.Tn[8] XThR.Tn[3] 0.28739f
C5038 XA.XIR[2].XIC[12].icell.Ien VPWR 0.1903f
C5039 XA.XIR[0].XIC[9].icell.Ien XA.XIR[0].XIC[10].icell.Ien 0.00214f
C5040 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.PDM 0.00591f
C5041 XA.XIR[7].XIC[12].icell.SM VPWR 0.00158f
C5042 XA.XIR[11].XIC[2].icell.PUM Vbias 0.0031f
C5043 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PUM 0.00465f
C5044 XA.XIR[2].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5045 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Ien 0.00584f
C5046 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6] 0.00341f
C5047 XA.XIR[10].XIC[0].icell.PUM VPWR 0.00937f
C5048 XA.XIR[2].XIC[8].icell.Ien Iout 0.06417f
C5049 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.03023f
C5050 XA.XIR[7].XIC[8].icell.SM Iout 0.00388f
C5051 XA.XIR[1].XIC[14].icell.Ien VPWR 0.19036f
C5052 XThC.Tn[5] VPWR 5.90052f
C5053 XA.XIR[7].XIC[8].icell.PDM Vbias 0.04261f
C5054 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.SM 0.00168f
C5055 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.15202f
C5056 XThR.Tn[0] XA.XIR[1].XIC[3].icell.SM 0.00121f
C5057 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04052f
C5058 XA.XIR[5].XIC[6].icell.Ien XA.XIR[5].XIC[7].icell.Ien 0.00214f
C5059 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.SM 0.00168f
C5060 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.SM 0.0039f
C5061 XA.XIR[9].XIC[1].icell.Ien Vbias 0.21098f
C5062 XThR.Tn[12] XA.XIR[13].XIC[4].icell.Ien 0.00338f
C5063 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02762f
C5064 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PUM 0.00465f
C5065 XA.XIR[1].XIC[10].icell.Ien Iout 0.06417f
C5066 XThR.XTB7.B a_n1049_6699# 0.0036f
C5067 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.SM 0.00168f
C5068 XA.XIR[15].XIC[6].icell.PDM Vbias 0.04261f
C5069 XA.XIR[6].XIC_15.icell.PDM Vbias 0.04401f
C5070 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00584f
C5071 XA.XIR[4].XIC[3].icell.Ien Vbias 0.21098f
C5072 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C5073 XThR.Tn[7] XA.XIR[8].XIC[9].icell.SM 0.00121f
C5074 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11336f
C5075 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C5076 XThC.Tn[11] XThR.Tn[0] 0.28749f
C5077 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.03425f
C5078 XThC.Tn[13] XThR.Tn[5] 0.2874f
C5079 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.03425f
C5080 XA.XIR[12].XIC[1].icell.Ien VPWR 0.1903f
C5081 XThR.Tn[5] XA.XIR[6].XIC[5].icell.SM 0.00121f
C5082 XThR.Tn[11] XA.XIR[12].XIC[7].icell.Ien 0.00338f
C5083 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.03425f
C5084 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C5085 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00584f
C5086 XA.XIR[7].XIC[12].icell.Ien XA.XIR[7].XIC[13].icell.Ien 0.00214f
C5087 XA.XIR[9].XIC[4].icell.PDM Vbias 0.04261f
C5088 XThR.Tn[3] XA.XIR[4].XIC_15.icell.PDM 0.00172f
C5089 a_7875_9569# Vbias 0.00315f
C5090 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.15202f
C5091 XThR.XTBN.Y a_n997_1579# 0.23006f
C5092 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C5093 XA.XIR[7].XIC[12].icell.PDM VPWR 0.00799f
C5094 XThC.XTB2.Y Vbias 0.0123f
C5095 XThR.XTB7.Y a_n1049_5317# 0.27822f
C5096 XA.XIR[5].XIC[2].icell.Ien VPWR 0.1903f
C5097 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C5098 XA.XIR[9].XIC[6].icell.Ien Vbias 0.21098f
C5099 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.03425f
C5100 XA.XIR[7].XIC[0].icell.PDM Iout 0.00117f
C5101 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C5102 XThR.Tn[1] XA.XIR[2].XIC[11].icell.Ien 0.00338f
C5103 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PUM 0.00465f
C5104 XThR.Tn[9] XA.XIR[10].XIC[0].icell.SM 0.00127f
C5105 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.SM 0.00168f
C5106 XA.XIR[15].XIC[10].icell.PDM VPWR 0.0114f
C5107 XA.XIR[4].XIC[5].icell.PUM VPWR 0.00937f
C5108 XA.XIR[10].XIC[0].icell.SM Iout 0.00388f
C5109 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02762f
C5110 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02762f
C5111 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C5112 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.15202f
C5113 XA.XIR[6].XIC[7].icell.PDM Iout 0.00117f
C5114 XA.XIR[6].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.SM 0.0039f
C5115 XA.XIR[3].XIC[9].icell.PUM Vbias 0.0031f
C5116 XA.XIR[14].XIC[4].icell.PDM Iout 0.00117f
C5117 XA.XIR[1].XIC[9].icell.PDM Vbias 0.04261f
C5118 XA.XIR[5].XIC[14].icell.PDM Iout 0.00117f
C5119 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PUM 0.00465f
C5120 XA.XIR[6].XIC[12].icell.SM Vbias 0.00701f
C5121 XA.XIR[9].XIC[8].icell.PDM VPWR 0.00799f
C5122 a_10051_9569# VPWR 0.00319f
C5123 XA.XIR[10].XIC[13].icell.SM Vbias 0.00701f
C5124 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.Ien 0.00584f
C5125 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PUM 0.00465f
C5126 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Iout 0.00347f
C5127 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C5128 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.SM 0.00168f
C5129 XA.XIR[0].XIC[0].icell.PDM VPWR 0.00774f
C5130 XA.XIR[13].XIC[8].icell.PDM Iout 0.00117f
C5131 XA.XIR[4].XIC[9].icell.PDM Vbias 0.04261f
C5132 XA.XIR[7].XIC[2].icell.Ien Vbias 0.21098f
C5133 XA.XIR[5].XIC_15.icell.Ien Vbias 0.21234f
C5134 XA.XIR[9].XIC[8].icell.PUM VPWR 0.00937f
C5135 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.SM 0.00168f
C5136 XThC.Tn[10] XThR.Tn[2] 0.28739f
C5137 XA.XIR[1].XIC[4].icell.PUM Vbias 0.0031f
C5138 XA.XIR[14].XIC[6].icell.SM Vbias 0.00701f
C5139 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.15202f
C5140 XA.XIR[12].XIC_15.icell.PDM Vbias 0.04401f
C5141 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C5142 XA.XIR[12].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5143 XA.XIR[13].XIC[8].icell.SM Vbias 0.00701f
C5144 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04031f
C5145 XA.XIR[8].XIC[12].icell.PUM Vbias 0.0031f
C5146 XA.XIR[14].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.SM 0.0039f
C5147 XA.XIR[3].XIC[9].icell.SM VPWR 0.00158f
C5148 XThR.Tn[11] XThR.Tn[12] 0.11452f
C5149 XA.XIR[11].XIC[12].icell.SM Iout 0.00388f
C5150 XA.XIR[1].XIC[13].icell.PDM VPWR 0.00799f
C5151 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10] 0.00341f
C5152 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.SM 0.00168f
C5153 XA.XIR[6].XIC[14].icell.Ien VPWR 0.19036f
C5154 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.03425f
C5155 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.SM 0.00168f
C5156 XA.XIR[10].XIC[12].icell.PDM Iout 0.00117f
C5157 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14] 0.00341f
C5158 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04031f
C5159 XThR.Tn[3] a_n1049_6405# 0.00542f
C5160 XA.XIR[3].XIC[5].icell.SM Iout 0.00388f
C5161 XA.XIR[1].XIC[1].icell.PDM Iout 0.00117f
C5162 XA.XIR[4].XIC[13].icell.PDM VPWR 0.00799f
C5163 XA.XIR[2].XIC[2].icell.SM VPWR 0.00158f
C5164 XA.XIR[6].XIC[10].icell.Ien Iout 0.06417f
C5165 XA.XIR[7].XIC[4].icell.PUM VPWR 0.00937f
C5166 XThC.XTB7.A XThC.Tn[6] 0.10589f
C5167 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04031f
C5168 XA.XIR[13].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.SM 0.0039f
C5169 Vbias Iout 83.1596f
C5170 XA.XIR[1].XIC[4].icell.SM VPWR 0.00158f
C5171 XA.XIR[4].XIC[1].icell.PDM Iout 0.00117f
C5172 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5173 XA.XIR[13].XIC[13].icell.PDM Iout 0.00117f
C5174 XThR.Tn[9] Vbias 3.74874f
C5175 XA.XIR[14].XIC[8].icell.Ien VPWR 0.19084f
C5176 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02762f
C5177 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.Ien 0.00584f
C5178 XThR.XTB5.A XThR.XTBN.A 0.06303f
C5179 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.03023f
C5180 XA.XIR[4].XIC[14].icell.SM Iout 0.00388f
C5181 XA.XIR[3].XIC[9].icell.PDM Iout 0.00117f
C5182 XA.XIR[8].XIC[11].icell.PDM Iout 0.00117f
C5183 XA.XIR[0].XIC[14].icell.PUM Vbias 0.0031f
C5184 XA.XIR[14].XIC[4].icell.Ien Iout 0.06417f
C5185 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04031f
C5186 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00584f
C5187 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C5188 XA.XIR[13].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.SM 0.0039f
C5189 XA.XIR[8].XIC[12].icell.SM VPWR 0.00158f
C5190 XA.XIR[2].XIC_15.icell.PDM Iout 0.00133f
C5191 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.Ien 0.00584f
C5192 XA.XIR[13].XIC[6].icell.Ien Iout 0.06417f
C5193 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02762f
C5194 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C5195 XA.XIR[2].XIC[0].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00214f
C5196 XA.XIR[8].XIC[8].icell.SM Iout 0.00388f
C5197 XThR.Tn[12] XA.XIR[13].XIC[12].icell.SM 0.00121f
C5198 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.03425f
C5199 XThR.Tn[8] XA.XIR[9].XIC[8].icell.SM 0.00121f
C5200 XThC.Tn[8] XThR.Tn[11] 0.28739f
C5201 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PUM 0.00465f
C5202 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.SM 0.00168f
C5203 XThR.Tn[0] XA.XIR[0].XIC[12].icell.PDM 0.00341f
C5204 XThR.Tn[2] XA.XIR[3].XIC[3].icell.Ien 0.00338f
C5205 XThR.Tn[4] XA.XIR[5].XIC[10].icell.Ien 0.00338f
C5206 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39003f
C5207 XA.XIR[15].XIC[0].icell.Ien Vbias 0.17752f
C5208 XThR.Tn[1] XA.XIR[1].XIC[10].icell.PDM 0.00341f
C5209 XA.XIR[5].XIC[0].icell.SM Vbias 0.00675f
C5210 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PUM 0.00444f
C5211 XA.XIR[11].XIC[9].icell.Ien Iout 0.06417f
C5212 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C5213 XThR.XTBN.Y a_n1049_6699# 0.07601f
C5214 XThC.Tn[7] XThR.Tn[7] 0.28739f
C5215 XThR.Tn[3] XA.XIR[4].XIC[10].icell.Ien 0.00338f
C5216 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04031f
C5217 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C5218 XA.XIR[14].XIC[2].icell.PUM Vbias 0.0031f
C5219 XA.XIR[0].XIC[14].icell.SM VPWR 0.00207f
C5220 XA.XIR[13].XIC[0].icell.PUM VPWR 0.00937f
C5221 XThR.Tn[1] XA.XIR[2].XIC[1].icell.SM 0.00121f
C5222 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.SM 0.00168f
C5223 XThC.XTB7.B XThC.Tn[5] 0.00714f
C5224 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PUM 0.00465f
C5225 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04031f
C5226 XA.XIR[3].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.SM 0.0039f
C5227 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C5228 XA.XIR[10].XIC[3].icell.PDM Vbias 0.04261f
C5229 XA.XIR[0].XIC[10].icell.SM Iout 0.00367f
C5230 XA.XIR[10].XIC[11].icell.SM Vbias 0.00701f
C5231 XThC.Tn[4] Vbias 2.48532f
C5232 XThR.Tn[2] XA.XIR[2].XIC[7].icell.PDM 0.00341f
C5233 XThC.XTB6.Y XThC.Tn[13] 0.32552f
C5234 XThR.XTBN.A data[5] 0.0148f
C5235 XThR.Tn[13] XA.XIR[14].XIC[5].icell.SM 0.00121f
C5236 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04031f
C5237 XA.XIR[6].XIC[4].icell.PUM Vbias 0.0031f
C5238 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.SM 0.00168f
C5239 XA.XIR[15].XIC[2].icell.PUM VPWR 0.00937f
C5240 XThC.Tn[11] XThR.Tn[1] 0.28739f
C5241 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PUM 0.00186f
C5242 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.03425f
C5243 XA.XIR[15].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.SM 0.0039f
C5244 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.SM 0.00168f
C5245 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6] 0.00341f
C5246 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C5247 XA.XIR[15].XIC[5].icell.Ien Vbias 0.17899f
C5248 a_5949_9615# XThC.Tn[6] 0.0018f
C5249 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PUM 0.00465f
C5250 XA.XIR[2].XIC[13].icell.Ien Iout 0.06417f
C5251 XA.XIR[7].XIC[13].icell.SM Iout 0.00388f
C5252 XThR.Tn[0] XA.XIR[1].XIC[8].icell.SM 0.00121f
C5253 XA.XIR[5].XIC[5].icell.SM Vbias 0.00701f
C5254 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.15202f
C5255 XThC.XTB6.A data[1] 0.37233f
C5256 XThR.XTB4.Y a_n1049_6699# 0.23756f
C5257 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C5258 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C5259 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C5260 XThR.Tn[12] XA.XIR[13].XIC[9].icell.Ien 0.00338f
C5261 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C5262 XA.XIR[11].XIC[3].icell.PDM VPWR 0.00799f
C5263 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.SM 0.00168f
C5264 XA.XIR[1].XIC_15.icell.Ien Iout 0.0642f
C5265 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Ien 0.00232f
C5266 XA.XIR[11].XIC[10].icell.SM Iout 0.00388f
C5267 XA.XIR[4].XIC[8].icell.Ien Vbias 0.21098f
C5268 XThC.Tn[11] XThR.Tn[12] 0.28739f
C5269 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.03425f
C5270 XThR.Tn[7] XA.XIR[8].XIC[14].icell.SM 0.00121f
C5271 XA.XIR[10].XIC[7].icell.PDM VPWR 0.00799f
C5272 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C5273 XThR.XTB7.B XThR.Tn[8] 0.05091f
C5274 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C5275 XThR.XTB1.Y a_n1335_8331# 0.0097f
C5276 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PUM 0.00465f
C5277 XA.XIR[4].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.SM 0.0039f
C5278 XA.XIR[13].XIC[0].icell.SM Iout 0.00388f
C5279 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PUM 0.00465f
C5280 XThR.Tn[5] XA.XIR[6].XIC[10].icell.SM 0.00121f
C5281 XThC.XTBN.Y XThC.Tn[9] 0.49745f
C5282 XA.XIR[8].XIC[2].icell.Ien Vbias 0.21098f
C5283 XThC.Tn[6] XThR.Tn[3] 0.28739f
C5284 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C5285 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02762f
C5286 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Ien 0.00584f
C5287 XA.XIR[10].XIC[14].icell.PUM Vbias 0.0031f
C5288 XA.XIR[15].XIC_15.icell.SM Vbias 0.00701f
C5289 XA.XIR[6].XIC[4].icell.SM VPWR 0.00158f
C5290 XA.XIR[2].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.SM 0.0039f
C5291 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.15202f
C5292 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08547f
C5293 XA.XIR[2].XIC[2].icell.PUM Vbias 0.0031f
C5294 XA.XIR[15].XIC[7].icell.PUM VPWR 0.00937f
C5295 XA.XIR[0].XIC[11].icell.PDM Vbias 0.04282f
C5296 XA.XIR[11].XIC[3].icell.PUM Vbias 0.0031f
C5297 XA.XIR[5].XIC[7].icell.Ien VPWR 0.1903f
C5298 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PUM 0.00465f
C5299 XThR.XTB7.A a_n1049_5611# 0.01824f
C5300 XThC.XTB7.B a_10051_9569# 0.00209f
C5301 XThC.Tn[10] XThR.Tn[10] 0.28739f
C5302 XA.XIR[13].XIC[13].icell.SM Vbias 0.00701f
C5303 XThC.Tn[0] XThR.Tn[0] 0.28842f
C5304 XA.XIR[9].XIC[11].icell.Ien Vbias 0.21098f
C5305 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.SM 0.00168f
C5306 XA.XIR[5].XIC[3].icell.Ien Iout 0.06417f
C5307 XA.XIR[4].XIC[10].icell.PUM VPWR 0.00937f
C5308 XA.XIR[7].XIC_15.icell.PDM Iout 0.00133f
C5309 XA.XIR[8].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.SM 0.0039f
C5310 XA.XIR[10].XIC[5].icell.PUM Vbias 0.0031f
C5311 XThC.Tn[2] XThR.Tn[5] 0.28739f
C5312 XA.XIR[12].XIC[14].icell.PDM Vbias 0.04261f
C5313 XA.XIR[3].XIC[9].icell.Ien XA.XIR[3].XIC[10].icell.Ien 0.00214f
C5314 XA.XIR[0].XIC[1].icell.PUM VPWR 0.00877f
C5315 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02762f
C5316 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PUM 0.00465f
C5317 XThR.Tn[12] XA.XIR[13].XIC[10].icell.SM 0.00121f
C5318 XA.XIR[0].XIC[4].icell.Ien Vbias 0.21127f
C5319 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C5320 XThC.Tn[9] XThC.Tn[10] 0.07959f
C5321 XA.XIR[8].XIC[4].icell.PUM VPWR 0.00937f
C5322 XThR.XTB5.A XThR.XTB6.Y 0.00193f
C5323 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00584f
C5324 XThR.Tn[13] a_n997_1579# 0.19413f
C5325 XThR.Tn[2] XA.XIR[3].XIC[0].icell.Ien 0.00338f
C5326 XA.XIR[3].XIC[14].icell.PUM Vbias 0.0031f
C5327 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00584f
C5328 XThR.Tn[6] XA.XIR[7].XIC[2].icell.Ien 0.00338f
C5329 XA.XIR[10].XIC[11].icell.PDM Iout 0.00117f
C5330 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04031f
C5331 XA.XIR[12].XIC[2].icell.Ien VPWR 0.1903f
C5332 XA.XIR[15].XIC_15.icell.PDM Vbias 0.04401f
C5333 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00256f
C5334 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.Ien 0.00584f
C5335 XA.XIR[14].XIC[12].icell.SM Iout 0.00388f
C5336 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07079f
C5337 XA.XIR[11].XIC[3].icell.SM VPWR 0.00158f
C5338 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.SM 0.00168f
C5339 XA.XIR[7].XIC[7].icell.Ien Vbias 0.21098f
C5340 XA.XIR[9].XIC[11].icell.PDM Iout 0.00117f
C5341 XThC.XTB7.Y VPWR 1.07717f
C5342 XA.XIR[2].XIC[2].icell.Ien XA.XIR[2].XIC[3].icell.Ien 0.00214f
C5343 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C5344 XA.XIR[2].XIC[7].icell.PUM Vbias 0.0031f
C5345 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9] 0.00341f
C5346 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PUM 0.00465f
C5347 XA.XIR[13].XIC[12].icell.PDM Iout 0.00117f
C5348 XA.XIR[9].XIC[13].icell.PUM VPWR 0.00937f
C5349 XA.XIR[8].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.SM 0.0039f
C5350 XA.XIR[10].XIC[5].icell.SM VPWR 0.00158f
C5351 XA.XIR[1].XIC[9].icell.PUM Vbias 0.0031f
C5352 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C5353 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11] 0.00341f
C5354 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C5355 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.15202f
C5356 XA.XIR[10].XIC[9].icell.SM Vbias 0.00701f
C5357 XThR.Tn[14] XA.XIR[15].XIC[2].icell.Ien 0.00338f
C5358 XA.XIR[9].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.SM 0.0039f
C5359 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PUM 0.00465f
C5360 XA.XIR[1].XIC[0].icell.SM Iout 0.00388f
C5361 XA.XIR[10].XIC[1].icell.SM Iout 0.00388f
C5362 XThR.Tn[9] XA.XIR[10].XIC[1].icell.SM 0.00121f
C5363 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C5364 XA.XIR[0].XIC[6].icell.PUM VPWR 0.00877f
C5365 XA.XIR[1].XIC[4].icell.Ien XA.XIR[1].XIC[5].icell.Ien 0.00214f
C5366 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.SM 0.00168f
C5367 XThR.XTBN.A XThR.Tn[9] 0.12398f
C5368 XA.XIR[12].XIC_dummy_left.icell.Ien Vbias 0.00329f
C5369 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PUM 0.00465f
C5370 XA.XIR[3].XIC[14].icell.SM VPWR 0.00207f
C5371 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C5372 XA.XIR[11].XIC[14].icell.Ien Iout 0.06417f
C5373 XThR.Tn[6] Iout 1.1623f
C5374 XA.XIR[3].XIC[10].icell.SM Iout 0.00388f
C5375 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C5376 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.SM 0.00168f
C5377 XA.XIR[0].XIC[7].icell.Ien XA.XIR[0].XIC[7].icell.SM 0.0039f
C5378 XA.XIR[6].XIC_15.icell.Ien Iout 0.0642f
C5379 XA.XIR[2].XIC[7].icell.SM VPWR 0.00158f
C5380 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5381 XA.XIR[7].XIC[9].icell.PUM VPWR 0.00937f
C5382 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0279f
C5383 XA.XIR[1].XIC[9].icell.SM VPWR 0.00158f
C5384 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C5385 XA.XIR[8].XIC[12].icell.Ien XA.XIR[8].XIC[13].icell.Ien 0.00214f
C5386 XA.XIR[2].XIC[3].icell.SM Iout 0.00388f
C5387 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.SM 0.00168f
C5388 XThR.XTB6.A VPWR 0.68638f
C5389 XThC.Tn[8] XThR.Tn[14] 0.28739f
C5390 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04031f
C5391 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C5392 XA.XIR[5].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.SM 0.0039f
C5393 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C5394 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39f
C5395 a_6243_9615# Vbias 0.01019f
C5396 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C5397 XA.XIR[1].XIC[5].icell.SM Iout 0.00388f
C5398 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02762f
C5399 XA.XIR[14].XIC[9].icell.Ien Iout 0.06417f
C5400 XA.XIR[6].XIC[2].icell.PDM Vbias 0.04261f
C5401 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.03023f
C5402 XA.XIR[9].XIC[2].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00214f
C5403 XThR.XTB1.Y a_n1049_8581# 0.21263f
C5404 XA.XIR[10].XIC[12].icell.PUM Vbias 0.0031f
C5405 XA.XIR[12].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.SM 0.0039f
C5406 XThC.XTB3.Y a_5155_9615# 0.00913f
C5407 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.SM 0.00168f
C5408 XA.XIR[5].XIC[9].icell.PDM Vbias 0.04261f
C5409 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.0352f
C5410 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.15202f
C5411 XA.XIR[8].XIC[13].icell.SM Iout 0.00388f
C5412 XA.XIR[6].XIC[0].icell.PUM VPWR 0.00937f
C5413 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C5414 XThR.Tn[11] XA.XIR[12].XIC[2].icell.SM 0.00121f
C5415 XThR.Tn[8] XA.XIR[9].XIC[13].icell.SM 0.00121f
C5416 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C5417 XA.XIR[13].XIC[3].icell.PDM Vbias 0.04261f
C5418 XThR.Tn[2] XA.XIR[3].XIC[8].icell.Ien 0.00338f
C5419 XThR.Tn[12] XA.XIR[13].XIC[14].icell.Ien 0.00338f
C5420 XThR.Tn[0] VPWR 6.67008f
C5421 XA.XIR[13].XIC[11].icell.SM Vbias 0.00701f
C5422 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C5423 XThR.Tn[4] XA.XIR[5].XIC_15.icell.Ien 0.00117f
C5424 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04031f
C5425 XThR.Tn[4] XA.XIR[4].XIC[9].icell.PDM 0.00341f
C5426 XA.XIR[7].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.SM 0.0039f
C5427 XA.XIR[12].XIC[8].icell.PDM Vbias 0.04261f
C5428 XThR.XTB7.B a_n997_3755# 0.01174f
C5429 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C5430 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C5431 XA.XIR[10].XIC[1].icell.PUM VPWR 0.00937f
C5432 XThR.Tn[3] XA.XIR[4].XIC_15.icell.Ien 0.00117f
C5433 XThR.Tn[3] XA.XIR[3].XIC[10].icell.PDM 0.00341f
C5434 XThC.Tn[4] XThR.Tn[6] 0.28739f
C5435 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C5436 XA.XIR[9].XIC[1].icell.SM Vbias 0.00701f
C5437 XThR.Tn[1] XA.XIR[2].XIC[6].icell.SM 0.00121f
C5438 XA.XIR[6].XIC[6].icell.PDM VPWR 0.00799f
C5439 XThR.XTBN.Y XThR.Tn[8] 0.47811f
C5440 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C5441 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.Ien 0.00256f
C5442 XA.XIR[5].XIC[13].icell.PDM VPWR 0.00799f
C5443 XA.XIR[14].XIC[3].icell.PDM VPWR 0.00799f
C5444 XA.XIR[14].XIC[10].icell.SM Iout 0.00388f
C5445 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PUM 0.00465f
C5446 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.SM 0.00168f
C5447 XThC.Tn[6] XThR.Tn[11] 0.28739f
C5448 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.03425f
C5449 XA.XIR[10].XIC[13].icell.Ien Vbias 0.21098f
C5450 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C5451 XA.XIR[5].XIC[1].icell.PDM Iout 0.00117f
C5452 XA.XIR[13].XIC[7].icell.PDM VPWR 0.00799f
C5453 XA.XIR[3].XIC[4].icell.Ien Vbias 0.21098f
C5454 XA.XIR[15].XIC_dummy_right.icell.PUM Vbias 0.00223f
C5455 XA.XIR[0].XIC[14].icell.Ien XA.XIR[0].XIC_15.icell.Ien 0.00214f
C5456 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.SM 0.00168f
C5457 XA.XIR[6].XIC[9].icell.PUM Vbias 0.0031f
C5458 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C5459 XA.XIR[6].XIC[0].icell.SM Iout 0.00388f
C5460 XThC.XTB7.Y a_9827_9569# 0.00571f
C5461 XThR.XTB7.B a_n1049_5611# 0.00927f
C5462 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PUM 0.00465f
C5463 XA.XIR[5].XIC[10].icell.SM Vbias 0.00701f
C5464 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C5465 XThR.Tn[0] XA.XIR[1].XIC[13].icell.SM 0.00121f
C5466 XThR.Tn[4] Iout 1.16233f
C5467 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.Ien 0.00584f
C5468 XA.XIR[13].XIC[14].icell.PUM Vbias 0.0031f
C5469 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C5470 XA.XIR[5].XIC[11].icell.Ien XA.XIR[5].XIC[12].icell.Ien 0.00214f
C5471 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C5472 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02762f
C5473 XA.XIR[12].XIC[0].icell.PDM Iout 0.00117f
C5474 XA.XIR[9].XIC[3].icell.Ien VPWR 0.1903f
C5475 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00584f
C5476 XA.XIR[12].XIC[13].icell.PDM Vbias 0.04261f
C5477 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PUM 0.00465f
C5478 XA.XIR[3].XIC[4].icell.PDM Vbias 0.04261f
C5479 XA.XIR[8].XIC[6].icell.PDM Vbias 0.04261f
C5480 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C5481 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00584f
C5482 XA.XIR[4].XIC[13].icell.Ien Vbias 0.21098f
C5483 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C5484 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.03451f
C5485 XA.XIR[14].XIC[3].icell.PUM Vbias 0.0031f
C5486 XThR.XTB2.Y XThR.Tn[2] 0.00271f
C5487 XThC.XTB5.Y XThC.Tn[7] 0.00912f
C5488 XA.XIR[11].XIC[6].icell.PDM Iout 0.00117f
C5489 XA.XIR[11].XIC[12].icell.Ien Iout 0.06417f
C5490 XA.XIR[2].XIC[10].icell.PDM Vbias 0.04261f
C5491 XThC.Tn[10] XThR.Tn[13] 0.28739f
C5492 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.SM 0.00168f
C5493 XA.XIR[13].XIC[5].icell.PUM Vbias 0.0031f
C5494 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02762f
C5495 XThC.Tn[0] XThR.Tn[1] 0.28753f
C5496 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.03425f
C5497 XA.XIR[8].XIC[7].icell.Ien Vbias 0.21098f
C5498 XA.XIR[10].XIC[10].icell.PDM Iout 0.00117f
C5499 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04031f
C5500 XA.XIR[15].XIC[14].icell.PDM Vbias 0.04261f
C5501 XA.XIR[3].XIC[6].icell.PUM VPWR 0.00937f
C5502 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02762f
C5503 XA.XIR[1].XIC[0].icell.PDM VPWR 0.00799f
C5504 XThR.Tn[8] XThR.Tn[10] 0.00255f
C5505 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02762f
C5506 XA.XIR[12].XIC[5].icell.SM Vbias 0.00701f
C5507 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C5508 XA.XIR[6].XIC[9].icell.SM VPWR 0.00158f
C5509 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C5510 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PUM 0.00465f
C5511 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C5512 XThC.Tn[13] Iout 0.84238f
C5513 XThR.XTB7.A XThR.Tn[3] 0.0306f
C5514 XThC.Tn[13] XThR.Tn[9] 0.2874f
C5515 XA.XIR[10].XIC[14].icell.SM Vbias 0.00701f
C5516 XA.XIR[4].XIC[0].icell.PDM VPWR 0.00799f
C5517 XA.XIR[11].XIC[8].icell.PUM Vbias 0.0031f
C5518 XThR.Tn[4] XA.XIR[5].XIC[0].icell.SM 0.00121f
C5519 XThC.Tn[0] XThR.Tn[12] 0.28741f
C5520 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C5521 XA.XIR[5].XIC[12].icell.Ien VPWR 0.1903f
C5522 XA.XIR[6].XIC[5].icell.SM Iout 0.00388f
C5523 XThC.Tn[9] XThR.Tn[8] 0.28739f
C5524 XA.XIR[13].XIC[11].icell.PDM Iout 0.00117f
C5525 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7] 0.00341f
C5526 XThR.Tn[10] XA.XIR[11].XIC[1].icell.Ien 0.00338f
C5527 XA.XIR[5].XIC_dummy_right.icell.Ien Vbias 0.00288f
C5528 XA.XIR[3].XIC[8].icell.PDM VPWR 0.00799f
C5529 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00584f
C5530 XThR.Tn[3] XA.XIR[4].XIC[0].icell.SM 0.00121f
C5531 XThC.XTB6.A VPWR 0.68179f
C5532 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01577f
C5533 XA.XIR[5].XIC[8].icell.Ien Iout 0.06417f
C5534 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C5535 XA.XIR[10].XIC[10].icell.PUM Vbias 0.0031f
C5536 XA.XIR[14].XIC[3].icell.SM VPWR 0.00158f
C5537 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C5538 XA.XIR[8].XIC[10].icell.PDM VPWR 0.00799f
C5539 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.0353f
C5540 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13] 0.00341f
C5541 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.SM 0.00168f
C5542 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C5543 XA.XIR[0].XIC[9].icell.Ien Vbias 0.2113f
C5544 XThC.XTBN.A a_7875_9569# 0.01939f
C5545 XA.XIR[2].XIC[14].icell.PDM VPWR 0.00809f
C5546 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C5547 XThR.XTB7.A data[4] 0.8689f
C5548 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C5549 XA.XIR[13].XIC[5].icell.SM VPWR 0.00158f
C5550 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04031f
C5551 XThC.XTBN.Y XThC.Tn[7] 0.91493f
C5552 XA.XIR[12].XIC[6].icell.Ien XA.XIR[12].XIC[7].icell.Ien 0.00214f
C5553 XA.XIR[8].XIC[9].icell.PUM VPWR 0.00937f
C5554 XThC.Tn[4] XThR.Tn[4] 0.28739f
C5555 XThR.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.00338f
C5556 XA.XIR[13].XIC[9].icell.SM Vbias 0.00701f
C5557 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C5558 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C5559 XA.XIR[2].XIC[2].icell.PDM Iout 0.00117f
C5560 XThR.Tn[6] XA.XIR[7].XIC[7].icell.Ien 0.00338f
C5561 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C5562 XA.XIR[13].XIC[1].icell.SM Iout 0.00388f
C5563 XA.XIR[12].XIC[7].icell.Ien VPWR 0.1903f
C5564 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.SM 0.00168f
C5565 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12] 0.00341f
C5566 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.Ien 0.00584f
C5567 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Iout 0.00347f
C5568 XThC.XTB4.Y XThC.Tn[2] 0.0021f
C5569 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5570 XA.XIR[2].XIC[12].icell.PUM Vbias 0.0031f
C5571 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.03425f
C5572 XA.XIR[12].XIC[3].icell.Ien Iout 0.06417f
C5573 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C5574 XA.XIR[11].XIC[8].icell.SM VPWR 0.00158f
C5575 XA.XIR[7].XIC[12].icell.Ien Vbias 0.21098f
C5576 XThR.Tn[4] XA.XIR[5].XIC[5].icell.SM 0.00121f
C5577 XA.XIR[14].XIC[14].icell.Ien Iout 0.06417f
C5578 XA.XIR[11].XIC[4].icell.SM Iout 0.00388f
C5579 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.03425f
C5580 XA.XIR[1].XIC[14].icell.PUM Vbias 0.0031f
C5581 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.Ien 0.00584f
C5582 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C5583 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.15202f
C5584 XThR.Tn[14] XA.XIR[15].XIC[7].icell.Ien 0.00338f
C5585 XThR.Tn[3] XA.XIR[4].XIC[5].icell.SM 0.00121f
C5586 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PUM 0.00465f
C5587 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Iout 0.00347f
C5588 XA.XIR[10].XIC[6].icell.SM Iout 0.00388f
C5589 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.SM 0.00168f
C5590 XA.XIR[0].XIC[11].icell.PUM VPWR 0.00878f
C5591 XThR.Tn[9] XA.XIR[10].XIC[6].icell.SM 0.00121f
C5592 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5] 0.00341f
C5593 XA.XIR[10].XIC[11].icell.Ien Vbias 0.21098f
C5594 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.15202f
C5595 XA.XIR[4].XIC_15.icell.SM Iout 0.0047f
C5596 XA.XIR[3].XIC[1].icell.Ien Vbias 0.21098f
C5597 XThC.XTB7.A a_8739_10571# 0.00995f
C5598 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C5599 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38993f
C5600 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04031f
C5601 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PUM 0.00465f
C5602 XThR.XTB3.Y a_n1049_5317# 0.00899f
C5603 XA.XIR[12].XIC[1].icell.PUM Vbias 0.0031f
C5604 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PUM 0.00465f
C5605 XA.XIR[6].XIC[4].icell.Ien XA.XIR[6].XIC[5].icell.Ien 0.00214f
C5606 XA.XIR[13].XIC[12].icell.PUM Vbias 0.0031f
C5607 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PUM 0.00471f
C5608 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8] 0.00341f
C5609 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04031f
C5610 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C5611 XA.XIR[2].XIC[12].icell.SM VPWR 0.00158f
C5612 XA.XIR[7].XIC[14].icell.PUM VPWR 0.00937f
C5613 XThR.XTBN.Y a_n997_3755# 0.229f
C5614 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C5615 XA.XIR[1].XIC[0].icell.Ien VPWR 0.1903f
C5616 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C5617 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6] 0.00341f
C5618 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.15202f
C5619 XA.XIR[1].XIC[14].icell.SM VPWR 0.00207f
C5620 XA.XIR[2].XIC[8].icell.SM Iout 0.00388f
C5621 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C5622 XA.XIR[11].XIC[10].icell.Ien Iout 0.06417f
C5623 XA.XIR[7].XIC[10].icell.PDM Vbias 0.04261f
C5624 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C5625 XThR.Tn[12] XA.XIR[13].XIC[4].icell.SM 0.00121f
C5626 XA.XIR[4].XIC[0].icell.Ien VPWR 0.1903f
C5627 XA.XIR[1].XIC[10].icell.SM Iout 0.00388f
C5628 XThR.Tn[1] VPWR 6.67356f
C5629 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02762f
C5630 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PUM 0.00465f
C5631 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00584f
C5632 XA.XIR[15].XIC[8].icell.PDM Vbias 0.04261f
C5633 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C5634 XA.XIR[4].XIC[3].icell.SM Vbias 0.00701f
C5635 XA.XIR[0].XIC_15.icell.SM VPWR 0.00257f
C5636 XA.XIR[13].XIC[1].icell.PUM VPWR 0.00937f
C5637 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.15202f
C5638 XThC.XTBN.Y a_3773_9615# 0.08456f
C5639 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.15202f
C5640 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.Ien 0.00584f
C5641 XThR.XTB3.Y a_n1335_7243# 0.00941f
C5642 XThR.Tn[12] VPWR 7.57625f
C5643 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C5644 XThR.Tn[11] XA.XIR[12].XIC[7].icell.SM 0.00121f
C5645 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C5646 XThR.XTBN.Y a_n1049_5611# 0.0768f
C5647 XThR.Tn[2] XA.XIR[3].XIC[13].icell.Ien 0.00338f
C5648 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C5649 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.SM 0.00168f
C5650 a_8963_9569# Vbias 0.00243f
C5651 XA.XIR[9].XIC[6].icell.PDM Vbias 0.04261f
C5652 XThR.XTB4.Y a_n997_3755# 0.00497f
C5653 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C5654 data[0] Vbias 0.00282f
C5655 XA.XIR[15].XIC[2].icell.Ien VPWR 0.32895f
C5656 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PUM 0.00465f
C5657 XA.XIR[13].XIC[13].icell.Ien Vbias 0.21098f
C5658 XThC.Tn[6] XThR.Tn[14] 0.28739f
C5659 XA.XIR[11].XIC[0].icell.Ien Iout 0.06411f
C5660 XA.XIR[7].XIC[14].icell.PDM VPWR 0.00809f
C5661 XA.XIR[5].XIC[2].icell.SM VPWR 0.00158f
C5662 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C5663 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C5664 a_10051_9569# XThC.Tn[12] 0.00623f
C5665 XThC.XTB3.Y a_7875_9569# 0.0061f
C5666 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.15202f
C5667 XA.XIR[12].XIC[12].icell.PDM Vbias 0.04261f
C5668 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00214f
C5669 XA.XIR[9].XIC[6].icell.SM Vbias 0.00701f
C5670 XA.XIR[4].XIC[5].icell.Ien VPWR 0.1903f
C5671 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.03425f
C5672 XThR.Tn[1] XA.XIR[2].XIC[11].icell.SM 0.00121f
C5673 XA.XIR[7].XIC[2].icell.PDM Iout 0.00117f
C5674 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C5675 XThR.Tn[12] XA.XIR[13].XIC[10].icell.Ien 0.00338f
C5676 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C5677 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C5678 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C5679 XThR.XTB2.Y XThR.Tn[10] 0.00106f
C5680 XA.XIR[3].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.SM 0.0039f
C5681 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02762f
C5682 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C5683 XA.XIR[6].XIC[9].icell.PDM Iout 0.00117f
C5684 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PUM 0.00465f
C5685 XA.XIR[15].XIC[0].icell.PDM Iout 0.00117f
C5686 XThC.XTB2.Y XThC.Tn[2] 0.01113f
C5687 XA.XIR[15].XIC[13].icell.PDM Vbias 0.04261f
C5688 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5689 XA.XIR[3].XIC[9].icell.Ien Vbias 0.21098f
C5690 XA.XIR[1].XIC[11].icell.PDM Vbias 0.04261f
C5691 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C5692 XA.XIR[14].XIC[6].icell.PDM Iout 0.00117f
C5693 XA.XIR[14].XIC[12].icell.Ien Iout 0.06417f
C5694 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PUM 0.00465f
C5695 XA.XIR[6].XIC[14].icell.PUM Vbias 0.0031f
C5696 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02762f
C5697 XThR.XTB4.Y a_n1049_5611# 0.00465f
C5698 XThC.Tn[8] VPWR 6.8418f
C5699 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.03425f
C5700 XA.XIR[9].XIC[10].icell.PDM VPWR 0.00799f
C5701 XThR.XTB7.B XThR.Tn[3] 0.00532f
C5702 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5703 XA.XIR[13].XIC[10].icell.PDM Iout 0.00117f
C5704 XA.XIR[7].XIC_15.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Ien 0.00214f
C5705 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C5706 XA.XIR[0].XIC[2].icell.PDM VPWR 0.00774f
C5707 XThR.XTB3.Y a_n1049_6405# 0.00913f
C5708 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02762f
C5709 XA.XIR[4].XIC[11].icell.PDM Vbias 0.04261f
C5710 XA.XIR[11].XIC[3].icell.Ien XA.XIR[11].XIC[4].icell.Ien 0.00214f
C5711 XA.XIR[2].XIC[2].icell.Ien Vbias 0.21098f
C5712 XA.XIR[7].XIC[2].icell.SM Vbias 0.00701f
C5713 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.15202f
C5714 XA.XIR[9].XIC[8].icell.Ien VPWR 0.1903f
C5715 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C5716 XA.XIR[13].XIC[14].icell.SM Vbias 0.00701f
C5717 XA.XIR[1].XIC[4].icell.Ien Vbias 0.21104f
C5718 XA.XIR[7].XIC[0].icell.PUM VPWR 0.00937f
C5719 XA.XIR[14].XIC[8].icell.PUM Vbias 0.0031f
C5720 XThR.XTB7.B data[4] 0.01382f
C5721 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PUM 0.00465f
C5722 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C5723 XA.XIR[9].XIC[4].icell.Ien Iout 0.06417f
C5724 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C5725 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.SM 0.00168f
C5726 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.15202f
C5727 XThC.XTB6.A XThC.XTB7.B 1.47641f
C5728 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PUM 0.00465f
C5729 XA.XIR[10].XIC[5].icell.Ien XA.XIR[10].XIC[6].icell.Ien 0.00214f
C5730 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.03425f
C5731 XA.XIR[1].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.SM 0.0039f
C5732 XA.XIR[13].XIC[10].icell.PUM Vbias 0.0031f
C5733 XThR.XTB5.Y a_n1319_6405# 0.01188f
C5734 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04031f
C5735 a_n1049_5317# VPWR 0.72036f
C5736 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C5737 XA.XIR[11].XIC[13].icell.SM VPWR 0.00158f
C5738 XA.XIR[8].XIC[12].icell.Ien Vbias 0.21098f
C5739 XThR.XTB5.A bias[2] 0.00213f
C5740 XA.XIR[3].XIC[11].icell.PUM VPWR 0.00937f
C5741 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.0353f
C5742 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07214f
C5743 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10] 0.00341f
C5744 XA.XIR[6].XIC[14].icell.SM VPWR 0.00207f
C5745 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14] 0.00341f
C5746 XA.XIR[1].XIC[3].icell.PDM Iout 0.00117f
C5747 XA.XIR[6].XIC[10].icell.SM Iout 0.00388f
C5748 XA.XIR[7].XIC[4].icell.Ien VPWR 0.1903f
C5749 XA.XIR[2].XIC[4].icell.PUM VPWR 0.00937f
C5750 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07214f
C5751 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C5752 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C5753 XThR.Tn[2] XThR.Tn[3] 0.10553f
C5754 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C5755 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C5756 XA.XIR[1].XIC[6].icell.PUM VPWR 0.00937f
C5757 XA.XIR[4].XIC[3].icell.PDM Iout 0.00117f
C5758 XA.XIR[5].XIC[13].icell.Ien Iout 0.06417f
C5759 XA.XIR[8].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.SM 0.0039f
C5760 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C5761 XA.XIR[14].XIC[8].icell.SM VPWR 0.00158f
C5762 XA.XIR[3].XIC[14].icell.Ien XA.XIR[3].XIC_15.icell.Ien 0.00214f
C5763 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.15235f
C5764 XA.XIR[8].XIC[13].icell.PDM Iout 0.00117f
C5765 XA.XIR[3].XIC[11].icell.PDM Iout 0.00117f
C5766 XA.XIR[0].XIC[14].icell.Ien Vbias 0.2113f
C5767 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04052f
C5768 XA.XIR[14].XIC[4].icell.SM Iout 0.00388f
C5769 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.SM 0.00168f
C5770 XA.XIR[8].XIC[14].icell.PUM VPWR 0.00937f
C5771 XThC.Tn[2] Iout 0.84806f
C5772 XThC.Tn[2] XThR.Tn[9] 0.28739f
C5773 XThR.Tn[6] XA.XIR[7].XIC[12].icell.Ien 0.00338f
C5774 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00584f
C5775 XA.XIR[13].XIC[6].icell.SM Iout 0.00388f
C5776 XA.XIR[3].XIC_15.icell.SM VPWR 0.00275f
C5777 XA.XIR[4].XIC[4].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00214f
C5778 XA.XIR[13].XIC[11].icell.Ien Vbias 0.21098f
C5779 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.SM 0.00168f
C5780 XA.XIR[11].XIC_15.icell.PDM Iout 0.00133f
C5781 XThR.XTBN.Y a_n997_715# 0.21503f
C5782 XA.XIR[11].XIC_15.icell.Ien Iout 0.0642f
C5783 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.15202f
C5784 XA.XIR[12].XIC[8].icell.Ien Iout 0.06417f
C5785 XThR.Tn[0] XA.XIR[0].XIC[14].icell.PDM 0.00341f
C5786 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.03425f
C5787 XThR.Tn[2] XA.XIR[3].XIC[3].icell.SM 0.00121f
C5788 XA.XIR[1].XIC_dummy_left.icell.SM VPWR 0.00269f
C5789 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C5790 VPWR data[7] 0.212f
C5791 XThC.Tn[7] XThR.Tn[8] 0.28739f
C5792 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C5793 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.SM 0.00168f
C5794 XA.XIR[2].XIC[7].icell.Ien XA.XIR[2].XIC[8].icell.Ien 0.00214f
C5795 XThR.Tn[4] XA.XIR[5].XIC[10].icell.SM 0.00121f
C5796 XA.XIR[15].XIC[0].icell.SM Vbias 0.00675f
C5797 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.03547f
C5798 XThR.Tn[1] XA.XIR[1].XIC[12].icell.PDM 0.00341f
C5799 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C5800 XA.XIR[5].XIC[2].icell.PUM Vbias 0.0031f
C5801 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04031f
C5802 XThR.Tn[10] XA.XIR[11].XIC[2].icell.Ien 0.00338f
C5803 XA.XIR[4].XIC_dummy_left.icell.SM VPWR 0.00269f
C5804 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.15202f
C5805 XThR.Tn[3] XA.XIR[4].XIC[10].icell.SM 0.00121f
C5806 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.SM 0.00168f
C5807 XA.XIR[11].XIC[1].icell.PDM Vbias 0.04261f
C5808 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C5809 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.15202f
C5810 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.15202f
C5811 XA.XIR[1].XIC[9].icell.Ien XA.XIR[1].XIC[10].icell.Ien 0.00214f
C5812 XThR.XTB7.B a_n997_2667# 0.02071f
C5813 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C5814 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.03425f
C5815 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04031f
C5816 XA.XIR[14].XIC[10].icell.Ien Iout 0.06417f
C5817 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02762f
C5818 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.03425f
C5819 XA.XIR[10].XIC[5].icell.PDM Vbias 0.04261f
C5820 XA.XIR[5].XIC[0].icell.PDM VPWR 0.00799f
C5821 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C5822 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PUM 0.00465f
C5823 XThR.Tn[2] XA.XIR[2].XIC[9].icell.PDM 0.00341f
C5824 XA.XIR[6].XIC[1].icell.PUM VPWR 0.00937f
C5825 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04031f
C5826 XA.XIR[0].XIC[12].icell.Ien XA.XIR[0].XIC[12].icell.SM 0.0039f
C5827 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.03425f
C5828 XThC.XTB3.Y XThC.Tn[4] 0.00382f
C5829 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.15202f
C5830 XA.XIR[6].XIC[4].icell.Ien Vbias 0.21098f
C5831 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C5832 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.Ien 0.00584f
C5833 a_n1049_6405# VPWR 0.72095f
C5834 XThR.Tn[12] XA.XIR[13].XIC_15.icell.Ien 0.00117f
C5835 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.01438f
C5836 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C5837 XA.XIR[15].XIC[5].icell.SM Vbias 0.00701f
C5838 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C5839 XA.XIR[2].XIC[13].icell.SM Iout 0.00388f
C5840 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02762f
C5841 XThC.Tn[2] XThC.Tn[4] 0.02725f
C5842 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.03425f
C5843 XA.XIR[12].XIC[11].icell.PDM Vbias 0.04261f
C5844 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.SM 0.0039f
C5845 XA.XIR[5].XIC[7].icell.PUM Vbias 0.0031f
C5846 XA.XIR[5].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.SM 0.0039f
C5847 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C5848 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C5849 XA.XIR[11].XIC[5].icell.PDM VPWR 0.00799f
C5850 XA.XIR[4].XIC[8].icell.SM Vbias 0.00701f
C5851 XA.XIR[11].XIC[11].icell.SM VPWR 0.00158f
C5852 XA.XIR[9].XIC[7].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00214f
C5853 XA.XIR[4].XIC[1].icell.Ien Iout 0.06417f
C5854 XA.XIR[10].XIC[9].icell.PDM VPWR 0.00799f
C5855 XA.XIR[15].XIC[12].icell.PDM Vbias 0.04261f
C5856 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.03425f
C5857 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C5858 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.03425f
C5859 XThR.XTBN.Y XThR.Tn[3] 0.62502f
C5860 XA.XIR[12].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.SM 0.0039f
C5861 XA.XIR[8].XIC[2].icell.SM Vbias 0.00701f
C5862 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C5863 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01432f
C5864 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.SM 0.00168f
C5865 XA.XIR[6].XIC[6].icell.PUM VPWR 0.00937f
C5866 a_n1049_8581# XThR.Tn[0] 0.2685f
C5867 XThR.XTB7.B XThR.Tn[11] 0.03888f
C5868 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00584f
C5869 XThC.Tn[10] XThR.Tn[7] 0.28739f
C5870 XA.XIR[15].XIC[7].icell.Ien VPWR 0.32895f
C5871 XA.XIR[0].XIC[13].icell.PDM Vbias 0.04282f
C5872 XA.XIR[5].XIC[7].icell.SM VPWR 0.00158f
C5873 XA.XIR[11].XIC[3].icell.Ien Vbias 0.21098f
C5874 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C5875 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.03425f
C5876 XThC.XTB7.B XThC.Tn[8] 0.09736f
C5877 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.03425f
C5878 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.15202f
C5879 XA.XIR[9].XIC[11].icell.SM Vbias 0.00701f
C5880 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C5881 XA.XIR[15].XIC[3].icell.Ien Iout 0.06807f
C5882 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.389f
C5883 XA.XIR[5].XIC[3].icell.SM Iout 0.00388f
C5884 XA.XIR[10].XIC[5].icell.Ien Vbias 0.21098f
C5885 XThC.XTB7.Y XThC.Tn[12] 0.07222f
C5886 XA.XIR[4].XIC[10].icell.Ien VPWR 0.1903f
C5887 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18966f
C5888 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PUM 0.00465f
C5889 XA.XIR[4].XIC[6].icell.Ien Iout 0.06417f
C5890 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Iout 0.00347f
C5891 XA.XIR[14].XIC[0].icell.Ien XA.XIR[14].XIC[1].icell.Ien 0.00214f
C5892 XA.XIR[2].XIC[1].icell.PDM VPWR 0.00799f
C5893 XA.XIR[0].XIC[4].icell.SM Vbias 0.00716f
C5894 XA.XIR[11].XIC[14].icell.PUM VPWR 0.00937f
C5895 XA.XIR[12].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.SM 0.0039f
C5896 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C5897 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PUM 0.00465f
C5898 XA.XIR[8].XIC[4].icell.Ien VPWR 0.1903f
C5899 XA.XIR[3].XIC[14].icell.Ien Vbias 0.21098f
C5900 XThR.Tn[13] XA.XIR[14].XIC[1].icell.Ien 0.00338f
C5901 XThR.Tn[2] XA.XIR[3].XIC[0].icell.SM 0.00121f
C5902 XThR.Tn[6] XA.XIR[7].XIC[2].icell.SM 0.00121f
C5903 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C5904 XA.XIR[12].XIC[2].icell.SM VPWR 0.00158f
C5905 XA.XIR[14].XIC[13].icell.SM VPWR 0.00158f
C5906 XThC.Tn[2] XA.XIR[0].XIC[4].icell.Ien 0.00191f
C5907 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C5908 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C5909 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PUM 0.00465f
C5910 XA.XIR[11].XIC[5].icell.PUM VPWR 0.00937f
C5911 XA.XIR[2].XIC[7].icell.Ien Vbias 0.21098f
C5912 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04031f
C5913 XA.XIR[7].XIC[7].icell.SM Vbias 0.00701f
C5914 XA.XIR[9].XIC[13].icell.PDM Iout 0.00117f
C5915 XA.XIR[10].XIC_15.icell.SM Vbias 0.00701f
C5916 XA.XIR[7].XIC[3].icell.Ien XA.XIR[7].XIC[4].icell.Ien 0.00214f
C5917 XA.XIR[15].XIC[1].icell.Ien XA.XIR[15].XIC[2].icell.Ien 0.00214f
C5918 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9] 0.00341f
C5919 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.03425f
C5920 XA.XIR[7].XIC[0].icell.Ien Iout 0.06411f
C5921 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.SM 0.0039f
C5922 XA.XIR[9].XIC[13].icell.Ien VPWR 0.1903f
C5923 XA.XIR[10].XIC[7].icell.PUM VPWR 0.00937f
C5924 XA.XIR[1].XIC[9].icell.Ien Vbias 0.21104f
C5925 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C5926 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11] 0.00341f
C5927 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.Ien 0.00584f
C5928 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.03425f
C5929 XThR.Tn[14] XA.XIR[15].XIC[2].icell.SM 0.00121f
C5930 a_7331_10587# data[0] 0.00451f
C5931 XA.XIR[9].XIC[9].icell.Ien Iout 0.06417f
C5932 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.15202f
C5933 XThC.Tn[9] XThR.Tn[3] 0.28739f
C5934 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00584f
C5935 XA.XIR[0].XIC[6].icell.Ien VPWR 0.18973f
C5936 XThR.Tn[7] XA.XIR[8].XIC[1].icell.Ien 0.00338f
C5937 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C5938 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C5939 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.03425f
C5940 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C5941 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C5942 XA.XIR[0].XIC[2].icell.Ien Iout 0.06389f
C5943 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Iout 0.00347f
C5944 XA.XIR[11].XIC[14].icell.PDM Iout 0.00117f
C5945 XA.XIR[6].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.SM 0.0039f
C5946 XThC.Tn[6] VPWR 5.90436f
C5947 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.15222f
C5948 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8] 0.00341f
C5949 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C5950 XA.XIR[2].XIC[9].icell.PUM VPWR 0.00937f
C5951 XA.XIR[7].XIC[9].icell.Ien VPWR 0.1903f
C5952 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.15202f
C5953 XA.XIR[11].XIC[9].icell.SM VPWR 0.00158f
C5954 XA.XIR[14].XIC_15.icell.PDM Iout 0.00133f
C5955 XThC.Tn[12] XThR.Tn[0] 0.28786f
C5956 XA.XIR[1].XIC[11].icell.PUM VPWR 0.00937f
C5957 XA.XIR[7].XIC[5].icell.Ien Iout 0.06417f
C5958 XA.XIR[14].XIC_15.icell.Ien Iout 0.0642f
C5959 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04031f
C5960 XThC.Tn[14] XThR.Tn[5] 0.28745f
C5961 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.SM 0.00168f
C5962 XThR.XTBN.Y a_n997_2667# 0.22784f
C5963 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C5964 XA.XIR[12].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.SM 0.0039f
C5965 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PUM 0.00465f
C5966 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.SM 0.00168f
C5967 XA.XIR[6].XIC[4].icell.PDM Vbias 0.04261f
C5968 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C5969 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C5970 XThR.Tn[7] XA.XIR[8].XIC[6].icell.Ien 0.00338f
C5971 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C5972 XThC.XTB3.Y a_6243_9615# 0.00899f
C5973 XA.XIR[5].XIC[11].icell.PDM Vbias 0.04261f
C5974 XThR.Tn[8] a_n997_3979# 0.1927f
C5975 XA.XIR[14].XIC[1].icell.PDM Vbias 0.04261f
C5976 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C5977 XThR.Tn[5] XA.XIR[6].XIC[2].icell.Ien 0.00338f
C5978 XThR.Tn[8] XA.XIR[9].XIC_15.icell.PUM 0.00186f
C5979 XA.XIR[2].XIC[0].icell.Ien VPWR 0.1903f
C5980 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.03425f
C5981 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.SM 0.00168f
C5982 XA.XIR[13].XIC[5].icell.PDM Vbias 0.04261f
C5983 XThR.Tn[2] XA.XIR[3].XIC[8].icell.SM 0.00121f
C5984 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02762f
C5985 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.15202f
C5986 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02762f
C5987 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04031f
C5988 XThR.Tn[4] XA.XIR[4].XIC[11].icell.PDM 0.00341f
C5989 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01746f
C5990 XA.XIR[12].XIC[10].icell.PDM Vbias 0.04261f
C5991 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.03425f
C5992 XA.XIR[7].XIC[1].icell.PDM VPWR 0.00799f
C5993 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.Ien 0.00584f
C5994 XA.XIR[10].XIC[1].icell.Ien VPWR 0.1903f
C5995 XThR.Tn[10] XA.XIR[11].XIC[7].icell.Ien 0.00338f
C5996 XA.XIR[1].XIC_15.icell.SM VPWR 0.00275f
C5997 XThR.Tn[3] XA.XIR[3].XIC[12].icell.PDM 0.00341f
C5998 XA.XIR[8].XIC_15.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00214f
C5999 XA.XIR[11].XIC[12].icell.PUM VPWR 0.00937f
C6000 XThR.XTB4.Y a_n997_2667# 0.07199f
C6001 XA.XIR[9].XIC[3].icell.PUM Vbias 0.0031f
C6002 XA.XIR[6].XIC[8].icell.PDM VPWR 0.00799f
C6003 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.15202f
C6004 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02762f
C6005 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.15202f
C6006 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C6007 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.SM 0.00168f
C6008 XA.XIR[15].XIC[11].icell.PDM Vbias 0.04261f
C6009 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.15202f
C6010 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07214f
C6011 XA.XIR[14].XIC[5].icell.PDM VPWR 0.00799f
C6012 XA.XIR[14].XIC[11].icell.SM VPWR 0.00158f
C6013 XA.XIR[6].XIC[9].icell.Ien XA.XIR[6].XIC[10].icell.Ien 0.00214f
C6014 XThR.XTBN.Y XThR.Tn[11] 0.52266f
C6015 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C6016 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.03425f
C6017 XA.XIR[3].XIC[4].icell.SM Vbias 0.00701f
C6018 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C6019 XThC.Tn[11] XThR.Tn[2] 0.28739f
C6020 XA.XIR[13].XIC[9].icell.PDM VPWR 0.00799f
C6021 XA.XIR[5].XIC[3].icell.PDM Iout 0.00117f
C6022 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC[0].icell.Ien 0.00214f
C6023 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.15202f
C6024 XA.XIR[6].XIC[9].icell.Ien Vbias 0.21098f
C6025 XThC.XTB7.Y a_10915_9569# 0.06874f
C6026 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C6027 XThR.Tn[0] XA.XIR[1].XIC_15.icell.PUM 0.00186f
C6028 XA.XIR[5].XIC[12].icell.PUM Vbias 0.0031f
C6029 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.SM 0.00168f
C6030 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.SM 0.00168f
C6031 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C6032 XA.XIR[12].XIC[2].icell.PDM Iout 0.00117f
C6033 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PUM 0.00465f
C6034 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.SM 0.00168f
C6035 XA.XIR[9].XIC[3].icell.SM VPWR 0.00158f
C6036 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.03425f
C6037 XA.XIR[4].XIC[13].icell.SM Vbias 0.00701f
C6038 XA.XIR[3].XIC[6].icell.PDM Vbias 0.04261f
C6039 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.SM 0.00168f
C6040 XA.XIR[14].XIC[3].icell.Ien Vbias 0.21098f
C6041 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00584f
C6042 XA.XIR[8].XIC[8].icell.PDM Vbias 0.04261f
C6043 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C6044 XA.XIR[11].XIC[8].icell.PDM Iout 0.00117f
C6045 XThR.XTB7.Y a_n997_1803# 0.00571f
C6046 XA.XIR[11].XIC[13].icell.Ien VPWR 0.1903f
C6047 XThR.Tn[7] XThR.Tn[8] 0.07425f
C6048 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C6049 XA.XIR[10].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.SM 0.0039f
C6050 XA.XIR[2].XIC[12].icell.PDM Vbias 0.04261f
C6051 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C6052 XA.XIR[13].XIC[5].icell.Ien Vbias 0.21098f
C6053 XThC.XTB7.A XThC.Tn[7] 0.00184f
C6054 XA.XIR[8].XIC[7].icell.SM Vbias 0.00701f
C6055 XA.XIR[14].XIC[3].icell.Ien XA.XIR[14].XIC[4].icell.Ien 0.00214f
C6056 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C6057 XA.XIR[3].XIC[6].icell.Ien VPWR 0.1903f
C6058 XA.XIR[1].XIC[2].icell.PDM VPWR 0.00799f
C6059 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.15202f
C6060 XA.XIR[6].XIC[11].icell.PUM VPWR 0.00937f
C6061 XA.XIR[12].XIC[7].icell.PUM Vbias 0.0031f
C6062 XA.XIR[14].XIC[14].icell.PUM VPWR 0.00937f
C6063 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PUM 0.00465f
C6064 XA.XIR[3].XIC[2].icell.Ien Iout 0.06417f
C6065 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00584f
C6066 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.03425f
C6067 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.SM 0.00168f
C6068 XA.XIR[10].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6069 XA.XIR[4].XIC[2].icell.PDM VPWR 0.00799f
C6070 XA.XIR[11].XIC[8].icell.Ien Vbias 0.21098f
C6071 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7] 0.00341f
C6072 XA.XIR[5].XIC[12].icell.SM VPWR 0.00158f
C6073 XA.XIR[12].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.SM 0.0039f
C6074 XThR.Tn[10] XThR.Tn[11] 0.05908f
C6075 XA.XIR[13].XIC[5].icell.Ien XA.XIR[13].XIC[6].icell.Ien 0.00214f
C6076 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.SM 0.00168f
C6077 XA.XIR[15].XIC[8].icell.Ien Iout 0.06807f
C6078 XA.XIR[3].XIC[10].icell.PDM VPWR 0.00799f
C6079 XA.XIR[8].XIC[12].icell.PDM VPWR 0.00799f
C6080 XA.XIR[5].XIC[8].icell.SM Iout 0.00388f
C6081 XA.XIR[4].XIC_15.icell.Ien VPWR 0.25566f
C6082 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C6083 XA.XIR[14].XIC[5].icell.PUM VPWR 0.00937f
C6084 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.SM 0.00168f
C6085 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PUM 0.00429f
C6086 XA.XIR[13].XIC_15.icell.SM Vbias 0.00701f
C6087 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13] 0.00341f
C6088 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C6089 XA.XIR[3].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.SM 0.0039f
C6090 XThC.Tn[9] XThR.Tn[11] 0.28739f
C6091 XA.XIR[0].XIC[9].icell.SM Vbias 0.00716f
C6092 XThC.XTBN.A a_8963_9569# 0.01679f
C6093 XA.XIR[4].XIC[11].icell.Ien Iout 0.06417f
C6094 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6095 XA.XIR[8].XIC[0].icell.PDM Iout 0.00117f
C6096 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04031f
C6097 XThC.XTBN.A data[0] 0.02545f
C6098 XA.XIR[13].XIC[7].icell.PUM VPWR 0.00937f
C6099 XA.XIR[8].XIC[9].icell.Ien VPWR 0.1903f
C6100 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04031f
C6101 XA.XIR[2].XIC[4].icell.PDM Iout 0.00117f
C6102 XThR.Tn[6] XA.XIR[7].XIC[7].icell.SM 0.00121f
C6103 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02762f
C6104 XA.XIR[11].XIC[13].icell.PDM Iout 0.00117f
C6105 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C6106 XA.XIR[11].XIC[14].icell.SM VPWR 0.00207f
C6107 XA.XIR[4].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.SM 0.0039f
C6108 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C6109 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C6110 XA.XIR[12].XIC[7].icell.SM VPWR 0.00158f
C6111 XA.XIR[8].XIC[5].icell.Ien Iout 0.06417f
C6112 XA.XIR[6].XIC_15.icell.SM VPWR 0.00275f
C6113 XThR.Tn[8] XA.XIR[9].XIC[5].icell.Ien 0.00338f
C6114 XThR.XTB6.A a_n1319_5317# 0.00295f
C6115 XThR.Tn[0] XA.XIR[0].XIC[1].icell.PDM 0.00341f
C6116 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C6117 XA.XIR[12].XIC[3].icell.SM Iout 0.00388f
C6118 XA.XIR[11].XIC[8].icell.Ien XA.XIR[11].XIC[9].icell.Ien 0.00214f
C6119 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Ien 0.00584f
C6120 XA.XIR[2].XIC[12].icell.Ien Vbias 0.21098f
C6121 XA.XIR[11].XIC[10].icell.PUM VPWR 0.00937f
C6122 XA.XIR[7].XIC[12].icell.SM Vbias 0.00701f
C6123 XA.XIR[2].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.SM 0.0039f
C6124 XThC.XTB7.B XThC.Tn[6] 0.05039f
C6125 XA.XIR[14].XIC[14].icell.PDM Iout 0.00117f
C6126 XThC.XTB5.Y XThC.Tn[10] 0.01742f
C6127 XA.XIR[1].XIC[14].icell.Ien Vbias 0.21104f
C6128 XThC.Tn[5] Vbias 2.31635f
C6129 XThR.XTB2.Y a_n997_3979# 0.00191f
C6130 XThC.XTB6.Y XThC.Tn[14] 0.00128f
C6131 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.03425f
C6132 XThR.Tn[14] XA.XIR[15].XIC[7].icell.SM 0.00121f
C6133 XA.XIR[9].XIC[14].icell.Ien Iout 0.06417f
C6134 XA.XIR[14].XIC[9].icell.SM VPWR 0.00158f
C6135 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C6136 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.15202f
C6137 XA.XIR[0].XIC[11].icell.Ien VPWR 0.19072f
C6138 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.0404f
C6139 XA.XIR[1].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.SM 0.0039f
C6140 XThC.XTB5.Y a_4861_9615# 0.0021f
C6141 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C6142 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5] 0.00341f
C6143 XA.XIR[12].XIC[9].icell.Ien XA.XIR[12].XIC[10].icell.Ien 0.00214f
C6144 XThC.Tn[12] XThR.Tn[1] 0.28739f
C6145 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.SM 0.00168f
C6146 XA.XIR[0].XIC[7].icell.Ien Iout 0.06389f
C6147 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04052f
C6148 XA.XIR[2].XIC_dummy_left.icell.SM VPWR 0.00269f
C6149 XA.XIR[12].XIC[1].icell.Ien Vbias 0.21098f
C6150 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C6151 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.04036f
C6152 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.03431f
C6153 XThR.Tn[13] XA.XIR[14].XIC[2].icell.Ien 0.00338f
C6154 XA.XIR[11].XIC[0].icell.PUM VPWR 0.00937f
C6155 XA.XIR[7].XIC[14].icell.Ien VPWR 0.19036f
C6156 XThC.Tn[12] XThR.Tn[12] 0.28739f
C6157 XA.XIR[2].XIC[14].icell.PUM VPWR 0.00937f
C6158 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C6159 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00584f
C6160 XThR.XTB7.A VPWR 0.88595f
C6161 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.15202f
C6162 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6] 0.00341f
C6163 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.15202f
C6164 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.Ien 0.00584f
C6165 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.04497f
C6166 XA.XIR[15].XIC[6].icell.Ien XA.XIR[15].XIC[7].icell.Ien 0.00214f
C6167 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6168 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02762f
C6169 XThR.Tn[0] XA.XIR[1].XIC[5].icell.Ien 0.00338f
C6170 XA.XIR[5].XIC[2].icell.Ien Vbias 0.21098f
C6171 XA.XIR[7].XIC[10].icell.Ien Iout 0.06417f
C6172 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.SM 0.00168f
C6173 XA.XIR[11].XIC[11].icell.Ien VPWR 0.1903f
C6174 XA.XIR[7].XIC[12].icell.PDM Vbias 0.04261f
C6175 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.SM 0.00168f
C6176 XThC.Tn[7] XThR.Tn[3] 0.28739f
C6177 XA.XIR[4].XIC[0].icell.SM VPWR 0.00158f
C6178 XThC.XTBN.Y XThC.Tn[10] 0.51405f
C6179 XThR.XTB5.Y XThR.Tn[6] 0.00349f
C6180 XA.XIR[4].XIC[5].icell.PUM Vbias 0.0031f
C6181 XA.XIR[15].XIC[10].icell.PDM Vbias 0.04261f
C6182 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.SM 0.00168f
C6183 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02762f
C6184 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C6185 XA.XIR[13].XIC[1].icell.Ien VPWR 0.1903f
C6186 XThR.Tn[7] XA.XIR[8].XIC[11].icell.Ien 0.00338f
C6187 XA.XIR[9].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.SM 0.0039f
C6188 XA.XIR[14].XIC[12].icell.PUM VPWR 0.00937f
C6189 XThC.XTBN.Y a_4861_9615# 0.07601f
C6190 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.Ien 0.00584f
C6191 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.Ien 0.00584f
C6192 XA.XIR[4].XIC[9].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00214f
C6193 XThR.Tn[5] XA.XIR[6].XIC[7].icell.Ien 0.00338f
C6194 XA.XIR[8].XIC[0].icell.Ien Iout 0.06411f
C6195 XThR.Tn[8] XA.XIR[9].XIC[0].icell.Ien 0.00338f
C6196 XA.XIR[12].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.SM 0.0039f
C6197 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.02762f
C6198 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.SM 0.0039f
C6199 XThC.Tn[11] XThR.Tn[10] 0.28739f
C6200 XThC.Tn[1] XThR.Tn[0] 0.28784f
C6201 XThC.Tn[3] XThR.Tn[5] 0.28739f
C6202 XA.XIR[0].XIC[0].icell.Ien XA.XIR[0].XIC[1].icell.Ien 0.00214f
C6203 XThR.Tn[2] XA.XIR[3].XIC[13].icell.SM 0.00121f
C6204 XA.XIR[2].XIC[12].icell.Ien XA.XIR[2].XIC[13].icell.Ien 0.00214f
C6205 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C6206 XThC.XTB5.Y a_5155_10571# 0.01188f
C6207 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C6208 a_10051_9569# Vbias 0.00678f
C6209 XA.XIR[9].XIC[8].icell.PDM Vbias 0.04261f
C6210 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C6211 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.SM 0.00168f
C6212 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.03425f
C6213 XA.XIR[0].XIC[0].icell.PDM Vbias 0.04227f
C6214 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C6215 XA.XIR[15].XIC[2].icell.SM VPWR 0.00158f
C6216 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6217 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PUM 0.00465f
C6218 XA.XIR[5].XIC[4].icell.PUM VPWR 0.00937f
C6219 XThC.Tn[9] XThC.Tn[11] 0.00252f
C6220 XThR.XTB6.A a_n1319_6405# 0.00306f
C6221 XThC.XTB3.Y a_8963_9569# 0.002f
C6222 XThC.XTB3.Y data[0] 0.03253f
C6223 XA.XIR[9].XIC[8].icell.PUM Vbias 0.0031f
C6224 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02762f
C6225 XA.XIR[1].XIC[14].icell.Ien XA.XIR[1].XIC_15.icell.Ien 0.00214f
C6226 XA.XIR[4].XIC[5].icell.SM VPWR 0.00158f
C6227 XA.XIR[8].XIC[3].icell.Ien XA.XIR[8].XIC[4].icell.Ien 0.00214f
C6228 XA.XIR[7].XIC[4].icell.PDM Iout 0.00117f
C6229 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C6230 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.SM 0.0039f
C6231 XA.XIR[9].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.SM 0.0039f
C6232 XA.XIR[4].XIC[1].icell.SM Iout 0.00388f
C6233 XA.XIR[15].XIC[2].icell.PDM Iout 0.00117f
C6234 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.15202f
C6235 XA.XIR[6].XIC[11].icell.PDM Iout 0.00117f
C6236 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.03425f
C6237 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Ien 0.00584f
C6238 XA.XIR[3].XIC[9].icell.SM Vbias 0.00701f
C6239 XA.XIR[14].XIC[8].icell.PDM Iout 0.00117f
C6240 XA.XIR[1].XIC[13].icell.PDM Vbias 0.04261f
C6241 XA.XIR[14].XIC[13].icell.Ien VPWR 0.19084f
C6242 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C6243 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00584f
C6244 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.03023f
C6245 XA.XIR[6].XIC[14].icell.Ien Vbias 0.21098f
C6246 XA.XIR[9].XIC[12].icell.PDM VPWR 0.00799f
C6247 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00584f
C6248 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.Ien 0.00584f
C6249 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C6250 XA.XIR[0].XIC[4].icell.PDM VPWR 0.00777f
C6251 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.SM 0.00168f
C6252 XA.XIR[4].XIC[13].icell.PDM Vbias 0.04261f
C6253 XA.XIR[2].XIC[2].icell.SM Vbias 0.00701f
C6254 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C6255 XA.XIR[9].XIC[0].icell.PDM Iout 0.00117f
C6256 XA.XIR[5].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.SM 0.0039f
C6257 XA.XIR[7].XIC[4].icell.PUM Vbias 0.0031f
C6258 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9] 0.00341f
C6259 XA.XIR[1].XIC[1].icell.Ien VPWR 0.1903f
C6260 XThR.Tn[12] XA.XIR[13].XIC[0].icell.Ien 0.00368f
C6261 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C6262 XA.XIR[9].XIC[8].icell.SM VPWR 0.00158f
C6263 XA.XIR[13].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6264 XA.XIR[1].XIC[4].icell.SM Vbias 0.00704f
C6265 XA.XIR[10].XIC[2].icell.Ien VPWR 0.1903f
C6266 XA.XIR[14].XIC[8].icell.Ien Vbias 0.21098f
C6267 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.03425f
C6268 XA.XIR[9].XIC[12].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00214f
C6269 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.SM 0.00168f
C6270 XA.XIR[9].XIC[4].icell.SM Iout 0.00388f
C6271 XThR.Tn[11] XThR.Tn[13] 0.00153f
C6272 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C6273 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.03425f
C6274 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.03425f
C6275 XA.XIR[0].XIC[1].icell.SM VPWR 0.00158f
C6276 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04031f
C6277 XThC.Tn[0] XThR.Tn[2] 0.28748f
C6278 XA.XIR[11].XIC[12].icell.PDM Iout 0.00117f
C6279 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04031f
C6280 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C6281 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04031f
C6282 XA.XIR[8].XIC[12].icell.SM Vbias 0.00701f
C6283 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.Ien 0.00584f
C6284 XA.XIR[3].XIC[11].icell.Ien VPWR 0.1903f
C6285 XThC.Tn[9] XThR.Tn[14] 0.28739f
C6286 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10] 0.00341f
C6287 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02762f
C6288 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.15202f
C6289 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6290 XA.XIR[3].XIC[7].icell.Ien Iout 0.06417f
C6291 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14] 0.00341f
C6292 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.Ien 0.00584f
C6293 XA.XIR[1].XIC[5].icell.PDM Iout 0.00117f
C6294 XA.XIR[0].XIC[5].icell.Ien XA.XIR[0].XIC[6].icell.Ien 0.00214f
C6295 XA.XIR[14].XIC[13].icell.PDM Iout 0.00117f
C6296 XA.XIR[14].XIC[14].icell.SM VPWR 0.00207f
C6297 XA.XIR[7].XIC[4].icell.SM VPWR 0.00158f
C6298 XA.XIR[2].XIC[4].icell.Ien VPWR 0.1903f
C6299 XThR.Tn[1] a_n1049_7787# 0.26879f
C6300 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PUM 0.00465f
C6301 XA.XIR[10].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6302 XThC.XTB6.A XThC.Tn[1] 0.00411f
C6303 XA.XIR[4].XIC[5].icell.PDM Iout 0.00117f
C6304 XA.XIR[5].XIC[13].icell.SM Iout 0.00388f
C6305 XA.XIR[1].XIC[6].icell.Ien VPWR 0.1903f
C6306 XA.XIR[14].XIC[10].icell.PUM VPWR 0.00937f
C6307 XA.XIR[5].XIC[2].icell.Ien XA.XIR[5].XIC[3].icell.Ien 0.00214f
C6308 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C6309 XA.XIR[3].XIC[13].icell.PDM Iout 0.00117f
C6310 XA.XIR[1].XIC[2].icell.Ien Iout 0.06417f
C6311 a_5155_9615# XThC.Tn[3] 0.00508f
C6312 XA.XIR[4].XIC_dummy_right.icell.SM VPWR 0.00123f
C6313 XA.XIR[0].XIC[14].icell.SM Vbias 0.00716f
C6314 XA.XIR[8].XIC_15.icell.PDM Iout 0.00133f
C6315 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C6316 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C6317 XA.XIR[8].XIC[14].icell.Ien VPWR 0.19036f
C6318 XThR.Tn[7] XA.XIR[8].XIC[1].icell.SM 0.00121f
C6319 XThR.Tn[6] XA.XIR[7].XIC[12].icell.SM 0.00121f
C6320 XA.XIR[8].XIC[10].icell.Ien Iout 0.06417f
C6321 XThC.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.00109f
C6322 XThR.Tn[8] XA.XIR[9].XIC[10].icell.Ien 0.00338f
C6323 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PUM 0.00465f
C6324 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38912f
C6325 XThC.Tn[5] XThR.Tn[6] 0.28739f
C6326 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04675f
C6327 XThC.XTB1.Y data[0] 0.06453f
C6328 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.SM 0.00168f
C6329 XA.XIR[12].XIC[8].icell.SM Iout 0.00388f
C6330 XThR.XTB7.B VPWR 1.67447f
C6331 XA.XIR[7].XIC[8].icell.Ien XA.XIR[7].XIC[9].icell.Ien 0.00214f
C6332 XA.XIR[15].XIC[2].icell.PUM Vbias 0.0031f
C6333 XThR.Tn[1] XA.XIR[1].XIC[14].icell.PDM 0.00341f
C6334 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C6335 XThR.Tn[10] XA.XIR[11].XIC[2].icell.SM 0.00121f
C6336 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C6337 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.04036f
C6338 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PUM 0.00465f
C6339 XThC.Tn[7] XThR.Tn[11] 0.28739f
C6340 XA.XIR[11].XIC[3].icell.PDM Vbias 0.04261f
C6341 XThR.Tn[1] XA.XIR[2].XIC[3].icell.Ien 0.00338f
C6342 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.SM 0.00168f
C6343 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04031f
C6344 XA.XIR[14].XIC[11].icell.Ien VPWR 0.19084f
C6345 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PUM 0.00465f
C6346 XA.XIR[0].XIC[12].icell.Ien Iout 0.06389f
C6347 XA.XIR[10].XIC[7].icell.PDM Vbias 0.04261f
C6348 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.15202f
C6349 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.15202f
C6350 XA.XIR[5].XIC[2].icell.PDM VPWR 0.00799f
C6351 XThR.Tn[2] XA.XIR[2].XIC[11].icell.PDM 0.00341f
C6352 XA.XIR[6].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.SM 0.0039f
C6353 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02762f
C6354 XA.XIR[6].XIC[1].icell.Ien VPWR 0.1903f
C6355 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C6356 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Ien 0.00232f
C6357 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04031f
C6358 XThR.Tn[13] XA.XIR[14].XIC[7].icell.Ien 0.00338f
C6359 XThR.Tn[12] XA.XIR[13].XIC_15.icell.PDM 0.00172f
C6360 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.03425f
C6361 XA.XIR[6].XIC[4].icell.SM Vbias 0.00701f
C6362 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.Ien 0.00584f
C6363 XA.XIR[0].XIC_dummy_left.icell.PDM Vbias 0.00131f
C6364 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.15202f
C6365 XThC.XTB5.Y a_7651_9569# 0.00418f
C6366 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.SM 0.00168f
C6367 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C6368 XA.XIR[12].XIC[1].icell.PDM VPWR 0.00799f
C6369 XA.XIR[15].XIC[7].icell.PUM Vbias 0.0031f
C6370 XA.XIR[7].XIC_15.icell.Ien Iout 0.0642f
C6371 XThR.Tn[0] XA.XIR[1].XIC[10].icell.Ien 0.00338f
C6372 XThC.Tn[11] XThR.Tn[13] 0.28739f
C6373 XA.XIR[5].XIC[7].icell.Ien Vbias 0.21098f
C6374 XThR.Tn[2] VPWR 6.62952f
C6375 XA.XIR[5].XIC[0].icell.Ien Iout 0.06411f
C6376 XA.XIR[11].XIC[7].icell.PDM VPWR 0.00799f
C6377 XThC.Tn[1] XThR.Tn[1] 0.28739f
C6378 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C6379 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.SM 0.00168f
C6380 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C6381 XThR.Tn[13] XA.XIR[15].XIC_dummy_left.icell.PUM 0.00107f
C6382 XA.XIR[4].XIC[10].icell.PUM Vbias 0.0031f
C6383 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PUM 0.00465f
C6384 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.0353f
C6385 XA.XIR[0].XIC[1].icell.PUM Vbias 0.0031f
C6386 XThR.XTB7.Y a_n997_3979# 0.00477f
C6387 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.15202f
C6388 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C6389 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC[0].icell.Ien 0.00214f
C6390 XThC.Tn[14] Iout 0.84284f
C6391 XThC.Tn[14] XThR.Tn[9] 0.28745f
C6392 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PUM 0.00465f
C6393 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02762f
C6394 XThC.Tn[1] XThR.Tn[12] 0.28739f
C6395 XThR.Tn[5] XA.XIR[6].XIC[12].icell.Ien 0.00338f
C6396 XThC.Tn[10] XThR.Tn[8] 0.28739f
C6397 XA.XIR[8].XIC[4].icell.PUM Vbias 0.0031f
C6398 XA.XIR[3].XIC[1].icell.SM VPWR 0.00158f
C6399 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C6400 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PUM 0.00442f
C6401 XA.XIR[6].XIC[6].icell.Ien VPWR 0.1903f
C6402 XA.XIR[12].XIC[2].icell.Ien Vbias 0.21098f
C6403 XA.XIR[0].XIC_15.icell.Ien XA.XIR[0].XIC_15.icell.SM 0.0039f
C6404 XA.XIR[15].XIC[7].icell.SM VPWR 0.00158f
C6405 XA.XIR[7].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.SM 0.0039f
C6406 XA.XIR[0].XIC_15.icell.PDM Vbias 0.04422f
C6407 XA.XIR[5].XIC[9].icell.PUM VPWR 0.00937f
C6408 XA.XIR[11].XIC[3].icell.SM Vbias 0.00701f
C6409 XA.XIR[6].XIC[2].icell.Ien Iout 0.06417f
C6410 XThC.XTB7.Y Vbias 0.01727f
C6411 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C6412 XA.XIR[5].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.SM 0.0039f
C6413 XThC.XTBN.Y a_7651_9569# 0.23021f
C6414 XA.XIR[13].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.SM 0.0039f
C6415 XThC.Tn[5] XThR.Tn[4] 0.28739f
C6416 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C6417 XA.XIR[15].XIC[3].icell.SM Iout 0.00388f
C6418 XA.XIR[9].XIC[13].icell.PUM Vbias 0.0031f
C6419 XA.XIR[10].XIC[5].icell.SM Vbias 0.00701f
C6420 XA.XIR[4].XIC[10].icell.SM VPWR 0.00158f
C6421 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C6422 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.Ien 0.00584f
C6423 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.11857f
C6424 XA.XIR[10].XIC[0].icell.Ien XA.XIR[10].XIC[1].icell.Ien 0.00214f
C6425 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.PDM 0.00555f
C6426 XThC.XTB4.Y XThC.Tn[3] 0.18952f
C6427 XA.XIR[4].XIC[6].icell.SM Iout 0.00388f
C6428 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.15202f
C6429 XA.XIR[0].XIC[6].icell.PUM Vbias 0.0031f
C6430 XThC.Tn[0] XThR.Tn[10] 0.28736f
C6431 XA.XIR[2].XIC[3].icell.PDM VPWR 0.00799f
C6432 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.15202f
C6433 XA.XIR[11].XIC[11].icell.PDM Iout 0.00117f
C6434 XA.XIR[13].XIC[2].icell.Ien VPWR 0.1903f
C6435 XA.XIR[8].XIC[4].icell.SM VPWR 0.00158f
C6436 XA.XIR[6].XIC[14].icell.Ien XA.XIR[6].XIC_15.icell.Ien 0.00214f
C6437 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.03425f
C6438 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C6439 XA.XIR[3].XIC[14].icell.SM Vbias 0.00701f
C6440 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.Ien 0.00584f
C6441 XThR.Tn[13] XThR.Tn[14] 0.1554f
C6442 XA.XIR[12].XIC[4].icell.PUM VPWR 0.00937f
C6443 XA.XIR[14].XIC[12].icell.PDM Iout 0.00117f
C6444 XA.XIR[12].XIC[14].icell.Ien XA.XIR[12].XIC_15.icell.Ien 0.00214f
C6445 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.SM 0.00168f
C6446 XA.XIR[2].XIC[7].icell.SM Vbias 0.00701f
C6447 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04031f
C6448 XA.XIR[11].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.SM 0.0039f
C6449 XA.XIR[11].XIC[5].icell.Ien VPWR 0.1903f
C6450 XA.XIR[7].XIC[9].icell.PUM Vbias 0.0031f
C6451 XA.XIR[9].XIC_15.icell.PDM Iout 0.00133f
C6452 XThR.Tn[4] XA.XIR[5].XIC[2].icell.Ien 0.00338f
C6453 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9] 0.00341f
C6454 XA.XIR[9].XIC[13].icell.SM VPWR 0.00158f
C6455 XA.XIR[7].XIC[0].icell.SM Iout 0.00388f
C6456 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.15202f
C6457 XA.XIR[10].XIC[7].icell.Ien VPWR 0.1903f
C6458 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.SM 0.00168f
C6459 XA.XIR[15].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.SM 0.0039f
C6460 XA.XIR[1].XIC[9].icell.SM Vbias 0.00704f
C6461 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11] 0.00341f
C6462 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C6463 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C6464 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C6465 XA.XIR[3].XIC[1].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00214f
C6466 XThR.Tn[3] XA.XIR[4].XIC[2].icell.Ien 0.00338f
C6467 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C6468 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PUM 0.00465f
C6469 XA.XIR[13].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6470 XA.XIR[9].XIC[9].icell.SM Iout 0.00388f
C6471 XA.XIR[10].XIC[3].icell.Ien Iout 0.06417f
C6472 XA.XIR[0].XIC[6].icell.SM VPWR 0.00158f
C6473 XThR.XTB7.Y a_n997_2891# 0.00474f
C6474 XThC.XTB2.Y a_4067_9615# 0.02133f
C6475 XThR.Tn[9] XA.XIR[10].XIC[3].icell.Ien 0.00338f
C6476 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.SM 0.00168f
C6477 XA.XIR[10].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.SM 0.0039f
C6478 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C6479 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C6480 XA.XIR[12].XIC[13].icell.SM Iout 0.00388f
C6481 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02762f
C6482 XA.XIR[14].XIC[8].icell.Ien XA.XIR[14].XIC[9].icell.Ien 0.00214f
C6483 XA.XIR[0].XIC[2].icell.SM Iout 0.00367f
C6484 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C6485 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C6486 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04031f
C6487 XThR.XTBN.Y VPWR 4.54348f
C6488 XA.XIR[11].XIC_15.icell.SM VPWR 0.00275f
C6489 XA.XIR[3].XIC[12].icell.Ien Iout 0.06417f
C6490 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8] 0.00341f
C6491 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PUM 0.00465f
C6492 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.04036f
C6493 XA.XIR[2].XIC[9].icell.Ien VPWR 0.1903f
C6494 XThR.Tn[0] Vbias 3.76149f
C6495 XA.XIR[7].XIC[9].icell.SM VPWR 0.00158f
C6496 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C6497 XA.XIR[2].XIC[5].icell.Ien Iout 0.06417f
C6498 XA.XIR[15].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.SM 0.0039f
C6499 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PUM 0.00465f
C6500 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.15202f
C6501 XA.XIR[1].XIC[11].icell.Ien VPWR 0.1903f
C6502 XA.XIR[7].XIC[5].icell.SM Iout 0.00388f
C6503 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04031f
C6504 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C6505 XA.XIR[10].XIC[1].icell.PUM Vbias 0.0031f
C6506 XA.XIR[1].XIC[7].icell.Ien Iout 0.06417f
C6507 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.03425f
C6508 XA.XIR[6].XIC[6].icell.PDM Vbias 0.04261f
C6509 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C6510 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02762f
C6511 XThR.Tn[7] XA.XIR[8].XIC[6].icell.SM 0.00121f
C6512 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PUM 0.00465f
C6513 XThR.XTB2.Y a_n1049_6699# 0.00851f
C6514 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C6515 XThC.Tn[7] XThR.Tn[14] 0.28739f
C6516 XA.XIR[14].XIC[3].icell.PDM Vbias 0.04261f
C6517 XA.XIR[5].XIC[13].icell.PDM Vbias 0.04261f
C6518 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.15202f
C6519 XA.XIR[4].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.SM 0.0039f
C6520 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.SM 0.00168f
C6521 XA.XIR[8].XIC_15.icell.Ien Iout 0.0642f
C6522 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02762f
C6523 XThR.Tn[5] XA.XIR[6].XIC[2].icell.SM 0.00121f
C6524 a_10051_9569# XThC.Tn[13] 0.19413f
C6525 XThR.Tn[11] XA.XIR[12].XIC[4].icell.Ien 0.00338f
C6526 XThR.Tn[8] XA.XIR[9].XIC_15.icell.Ien 0.00117f
C6527 XThR.XTB4.Y VPWR 0.92827f
C6528 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C6529 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04052f
C6530 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C6531 XA.XIR[13].XIC[7].icell.PDM Vbias 0.04261f
C6532 XA.XIR[11].XIC[1].icell.PUM VPWR 0.00937f
C6533 XA.XIR[2].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.SM 0.0039f
C6534 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC[0].icell.Ien 0.00214f
C6535 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.15202f
C6536 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PUM 0.00465f
C6537 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04031f
C6538 XThR.Tn[4] XA.XIR[4].XIC[13].icell.PDM 0.00341f
C6539 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PUM 0.00465f
C6540 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C6541 XA.XIR[7].XIC[3].icell.PDM VPWR 0.00799f
C6542 XThR.Tn[10] VPWR 7.53208f
C6543 XThR.Tn[10] XA.XIR[11].XIC[7].icell.SM 0.00121f
C6544 XThR.Tn[3] XA.XIR[3].XIC[14].icell.PDM 0.00341f
C6545 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01745f
C6546 XA.XIR[9].XIC[3].icell.Ien Vbias 0.21098f
C6547 XThR.Tn[1] XA.XIR[2].XIC[8].icell.Ien 0.00338f
C6548 XA.XIR[15].XIC[1].icell.PDM VPWR 0.0114f
C6549 XA.XIR[6].XIC[10].icell.PDM VPWR 0.00799f
C6550 XA.XIR[1].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.SM 0.0039f
C6551 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C6552 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.SM 0.0039f
C6553 XThC.Tn[9] VPWR 6.83084f
C6554 XA.XIR[3].XIC[5].icell.Ien XA.XIR[3].XIC[6].icell.Ien 0.00214f
C6555 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC[0].icell.Ien 0.00214f
C6556 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.15202f
C6557 XThR.XTB5.A a_n1335_4229# 0.01243f
C6558 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02762f
C6559 XA.XIR[14].XIC[7].icell.PDM VPWR 0.00799f
C6560 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PUM 0.00465f
C6561 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.Ien 0.00584f
C6562 XA.XIR[5].XIC[5].icell.PDM Iout 0.00117f
C6563 XA.XIR[3].XIC[6].icell.PUM Vbias 0.0031f
C6564 XA.XIR[1].XIC[0].icell.PDM Vbias 0.04207f
C6565 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PUM 0.00465f
C6566 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02762f
C6567 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.SM 0.00168f
C6568 XA.XIR[6].XIC[9].icell.SM Vbias 0.00701f
C6569 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00584f
C6570 XA.XIR[15].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.SM 0.0039f
C6571 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C6572 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.Ien 0.00584f
C6573 XThR.Tn[0] XA.XIR[1].XIC_15.icell.Ien 0.00117f
C6574 XA.XIR[5].XIC[12].icell.Ien Vbias 0.21098f
C6575 XA.XIR[4].XIC[0].icell.PDM Vbias 0.04207f
C6576 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C6577 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C6578 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C6579 XA.XIR[12].XIC[4].icell.PDM Iout 0.00117f
C6580 XA.XIR[9].XIC[5].icell.PUM VPWR 0.00937f
C6581 XA.XIR[12].XIC[11].icell.SM Iout 0.00388f
C6582 XThC.XTB6.A Vbias 0.00648f
C6583 XA.XIR[4].XIC_15.icell.PUM Vbias 0.0031f
C6584 XA.XIR[8].XIC[10].icell.PDM Vbias 0.04261f
C6585 data[5] data[6] 0.01513f
C6586 XA.XIR[3].XIC[8].icell.PDM Vbias 0.04261f
C6587 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C6588 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C6589 XA.XIR[14].XIC[3].icell.SM Vbias 0.00701f
C6590 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C6591 XA.XIR[9].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.SM 0.0039f
C6592 XA.XIR[11].XIC[10].icell.PDM Iout 0.00117f
C6593 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00584f
C6594 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.SM 0.00168f
C6595 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02762f
C6596 XA.XIR[2].XIC[14].icell.PDM Vbias 0.04261f
C6597 XA.XIR[4].XIC[14].icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00214f
C6598 XA.XIR[13].XIC[5].icell.SM Vbias 0.00701f
C6599 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C6600 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.03425f
C6601 XA.XIR[8].XIC[9].icell.PUM Vbias 0.0031f
C6602 XA.XIR[3].XIC[6].icell.SM VPWR 0.00158f
C6603 XA.XIR[1].XIC[4].icell.PDM VPWR 0.00799f
C6604 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C6605 XA.XIR[8].XIC[0].icell.SM Iout 0.00388f
C6606 XA.XIR[6].XIC[11].icell.Ien VPWR 0.1903f
C6607 XThR.Tn[8] XA.XIR[9].XIC[0].icell.SM 0.00121f
C6608 XA.XIR[14].XIC[11].icell.PDM Iout 0.00117f
C6609 XThC.Tn[0] XThR.Tn[13] 0.28746f
C6610 XA.XIR[12].XIC[7].icell.Ien Vbias 0.21098f
C6611 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C6612 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.03425f
C6613 XA.XIR[3].XIC[2].icell.SM Iout 0.00388f
C6614 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C6615 a_4067_9615# XThC.Tn[4] 0.00141f
C6616 XA.XIR[6].XIC[7].icell.Ien Iout 0.06417f
C6617 XA.XIR[0].XIC[3].icell.Ien XA.XIR[0].XIC[3].icell.SM 0.0039f
C6618 XA.XIR[4].XIC[4].icell.PDM VPWR 0.00799f
C6619 XA.XIR[11].XIC[8].icell.SM Vbias 0.00701f
C6620 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7] 0.00341f
C6621 XA.XIR[5].XIC[14].icell.PUM VPWR 0.00937f
C6622 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04037f
C6623 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C6624 XA.XIR[15].XIC[8].icell.SM Iout 0.00388f
C6625 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C6626 XA.XIR[1].XIC[1].icell.SM VPWR 0.00158f
C6627 XA.XIR[8].XIC[8].icell.Ien XA.XIR[8].XIC[9].icell.Ien 0.00214f
C6628 XThC.Tn[3] Iout 0.8384f
C6629 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C6630 XThC.Tn[3] XThR.Tn[9] 0.28739f
C6631 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C6632 XA.XIR[3].XIC[12].icell.PDM VPWR 0.00799f
C6633 XA.XIR[8].XIC[14].icell.PDM VPWR 0.00809f
C6634 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C6635 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13] 0.00341f
C6636 XA.XIR[14].XIC[5].icell.Ien VPWR 0.19084f
C6637 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.03589f
C6638 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.15202f
C6639 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C6640 XA.XIR[3].XIC[0].icell.PDM Iout 0.00117f
C6641 XA.XIR[4].XIC[11].icell.SM Iout 0.00388f
C6642 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02762f
C6643 XThC.XTBN.A a_10051_9569# 0.00199f
C6644 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04031f
C6645 XA.XIR[8].XIC[2].icell.PDM Iout 0.00117f
C6646 XA.XIR[0].XIC[11].icell.PUM Vbias 0.0031f
C6647 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04031f
C6648 XA.XIR[13].XIC[7].icell.Ien VPWR 0.1903f
C6649 XThR.XTB6.A XThR.XTBN.A 0.0512f
C6650 XA.XIR[8].XIC[9].icell.SM VPWR 0.00158f
C6651 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6652 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6653 XA.XIR[2].XIC[6].icell.PDM Iout 0.00117f
C6654 XA.XIR[13].XIC[3].icell.Ien Iout 0.06417f
C6655 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C6656 XA.XIR[6].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6657 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02762f
C6658 XThR.XTB7.Y a_n997_1579# 0.013f
C6659 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.SM 0.00168f
C6660 XA.XIR[12].XIC[9].icell.PUM VPWR 0.00937f
C6661 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00584f
C6662 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.PDM 0.00591f
C6663 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.Ien 0.00584f
C6664 XA.XIR[8].XIC[5].icell.SM Iout 0.00388f
C6665 XThR.Tn[8] XA.XIR[9].XIC[5].icell.SM 0.00121f
C6666 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02762f
C6667 XThR.Tn[0] XA.XIR[0].XIC[3].icell.PDM 0.00341f
C6668 XA.XIR[2].XIC[12].icell.SM Vbias 0.00701f
C6669 XA.XIR[7].XIC[14].icell.PUM Vbias 0.0031f
C6670 a_n997_1803# VPWR 0.01991f
C6671 XA.XIR[7].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.SM 0.0039f
C6672 XThR.Tn[4] XA.XIR[5].XIC[7].icell.Ien 0.00338f
C6673 XA.XIR[14].XIC_15.icell.SM VPWR 0.00275f
C6674 XA.XIR[1].XIC[0].icell.Ien Vbias 0.20957f
C6675 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02762f
C6676 XThR.Tn[0] XA.XIR[1].XIC[0].icell.SM 0.00121f
C6677 XThR.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.00341f
C6678 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.03023f
C6679 XA.XIR[11].XIC[6].icell.Ien Iout 0.06417f
C6680 XThR.Tn[11] XA.XIR[12].XIC[12].icell.SM 0.00121f
C6681 XA.XIR[1].XIC[14].icell.SM Vbias 0.00704f
C6682 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Iout 0.00347f
C6683 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01432f
C6684 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.04036f
C6685 XThR.Tn[3] XA.XIR[4].XIC[7].icell.Ien 0.00338f
C6686 XThC.XTB7.A XThC.Tn[10] 0.00406f
C6687 XA.XIR[4].XIC[0].icell.Ien Vbias 0.20951f
C6688 XA.XIR[9].XIC[14].icell.SM Iout 0.00388f
C6689 XThR.Tn[1] Vbias 3.74893f
C6690 XA.XIR[0].XIC[11].icell.SM VPWR 0.00158f
C6691 XThC.XTB5.Y a_5949_9615# 0.0093f
C6692 XA.XIR[10].XIC[8].icell.Ien Iout 0.06417f
C6693 XThR.Tn[9] XA.XIR[10].XIC[8].icell.Ien 0.00338f
C6694 XA.XIR[3].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.SM 0.0039f
C6695 XThC.XTB3.Y XThC.Tn[5] 0.00384f
C6696 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PUM 0.00465f
C6697 XA.XIR[8].XIC[0].icell.PUM VPWR 0.00937f
C6698 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5] 0.00341f
C6699 XThC.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.00109f
C6700 XA.XIR[13].XIC[1].icell.PUM Vbias 0.0031f
C6701 XA.XIR[0].XIC_15.icell.SM Vbias 0.00716f
C6702 XThC.XTB7.A a_4861_9615# 0.02294f
C6703 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.Ien 0.00584f
C6704 XA.XIR[0].XIC[7].icell.SM Iout 0.00367f
C6705 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PUM 0.00465f
C6706 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02762f
C6707 XA.XIR[15].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.SM 0.0039f
C6708 XThC.Tn[3] XThC.Tn[4] 0.49877f
C6709 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.04036f
C6710 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02762f
C6711 XThR.Tn[12] Vbias 3.74784f
C6712 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PUM 0.00465f
C6713 XThR.Tn[13] XA.XIR[14].XIC[2].icell.SM 0.00121f
C6714 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PDM 0.00172f
C6715 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.SM 0.0039f
C6716 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.SM 0.00168f
C6717 XA.XIR[0].XIC[10].icell.Ien XA.XIR[0].XIC[11].icell.Ien 0.00214f
C6718 XA.XIR[7].XIC[14].icell.SM VPWR 0.00207f
C6719 XA.XIR[2].XIC[14].icell.Ien VPWR 0.19036f
C6720 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C6721 XA.XIR[12].XIC[9].icell.SM Iout 0.00388f
C6722 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C6723 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02762f
C6724 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6] 0.00341f
C6725 XA.XIR[2].XIC[10].icell.Ien Iout 0.06417f
C6726 XA.XIR[15].XIC[2].icell.Ien Vbias 0.17899f
C6727 XA.XIR[7].XIC[10].icell.SM Iout 0.00388f
C6728 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.15202f
C6729 XA.XIR[7].XIC[14].icell.PDM Vbias 0.04261f
C6730 XThR.Tn[0] XA.XIR[1].XIC[5].icell.SM 0.00121f
C6731 XA.XIR[5].XIC[2].icell.SM Vbias 0.00701f
C6732 XA.XIR[5].XIC[7].icell.Ien XA.XIR[5].XIC[8].icell.Ien 0.00214f
C6733 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C6734 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C6735 XA.XIR[14].XIC[0].icell.Ien VPWR 0.19084f
C6736 XA.XIR[8].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.SM 0.0039f
C6737 XThR.Tn[12] XA.XIR[13].XIC[6].icell.Ien 0.00338f
C6738 XA.XIR[4].XIC[2].icell.PUM VPWR 0.00937f
C6739 XA.XIR[1].XIC[12].icell.Ien Iout 0.06417f
C6740 XA.XIR[4].XIC[5].icell.Ien Vbias 0.21098f
C6741 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C6742 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00584f
C6743 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.SM 0.0039f
C6744 XThR.Tn[11] XA.XIR[12].XIC_15.icell.PUM 0.00186f
C6745 XThR.Tn[7] XA.XIR[8].XIC[11].icell.SM 0.00121f
C6746 XThR.Tn[13] VPWR 7.61336f
C6747 XThC.XTBN.Y a_5949_9615# 0.0768f
C6748 XThC.Tn[11] XThR.Tn[7] 0.28739f
C6749 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.03425f
C6750 XThR.Tn[11] XA.XIR[12].XIC[9].icell.Ien 0.00338f
C6751 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C6752 XThR.Tn[5] XA.XIR[6].XIC[7].icell.SM 0.00121f
C6753 XThC.XTB7.B XThC.Tn[9] 0.09571f
C6754 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Iout 0.00347f
C6755 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C6756 XThR.XTB2.Y XThR.Tn[8] 0.00167f
C6757 XThC.XTB7.Y XThC.Tn[13] 0.11626f
C6758 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C6759 XThR.Tn[2] XA.XIR[3].XIC_15.icell.PUM 0.00186f
C6760 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.SM 0.00168f
C6761 XA.XIR[6].XIC[1].icell.SM VPWR 0.00158f
C6762 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.15202f
C6763 XThC.Tn[8] Vbias 2.30271f
C6764 XA.XIR[7].XIC[13].icell.Ien XA.XIR[7].XIC[14].icell.Ien 0.00214f
C6765 XA.XIR[9].XIC[10].icell.PDM Vbias 0.04261f
C6766 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C6767 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.SM 0.00168f
C6768 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PUM 0.00465f
C6769 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.03425f
C6770 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.15202f
C6771 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02762f
C6772 XA.XIR[15].XIC[4].icell.PUM VPWR 0.00937f
C6773 XA.XIR[0].XIC[2].icell.PDM Vbias 0.04282f
C6774 XA.XIR[5].XIC[4].icell.Ien VPWR 0.1903f
C6775 XA.XIR[11].XIC[0].icell.SM Iout 0.00388f
C6776 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C6777 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PUM 0.00465f
C6778 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02762f
C6779 XA.XIR[15].XIC[9].icell.Ien XA.XIR[15].XIC[10].icell.Ien 0.00214f
C6780 XThC.XTB5.A XThC.XTBN.Y 0.00282f
C6781 XA.XIR[9].XIC[8].icell.Ien Vbias 0.21098f
C6782 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C6783 XThR.Tn[1] XA.XIR[2].XIC[13].icell.Ien 0.00338f
C6784 XA.XIR[7].XIC[6].icell.PDM Iout 0.00117f
C6785 XThR.XTB1.Y bias[2] 0.00393f
C6786 XThR.Tn[3] a_n1049_6699# 0.27008f
C6787 XA.XIR[4].XIC[7].icell.PUM VPWR 0.00937f
C6788 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PUM 0.00465f
C6789 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C6790 XA.XIR[6].XIC[13].icell.PDM Iout 0.00117f
C6791 XA.XIR[15].XIC[4].icell.PDM Iout 0.00117f
C6792 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C6793 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PUM 0.00471f
C6794 XA.XIR[12].XIC[2].icell.Ien XA.XIR[12].XIC[3].icell.Ien 0.00214f
C6795 XA.XIR[6].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.SM 0.0039f
C6796 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02762f
C6797 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PUM 0.00465f
C6798 XA.XIR[11].XIC[13].icell.SM Vbias 0.00701f
C6799 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.SM 0.00168f
C6800 XA.XIR[14].XIC[10].icell.PDM Iout 0.00117f
C6801 XA.XIR[3].XIC[11].icell.PUM Vbias 0.0031f
C6802 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C6803 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C6804 XA.XIR[1].XIC_15.icell.PDM Vbias 0.04401f
C6805 XA.XIR[15].XIC[13].icell.SM Iout 0.00388f
C6806 XA.XIR[6].XIC[14].icell.SM Vbias 0.00701f
C6807 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C6808 XA.XIR[9].XIC[14].icell.PDM VPWR 0.00809f
C6809 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.Ien 0.00584f
C6810 XThR.Tn[11] XA.XIR[12].XIC[10].icell.SM 0.00121f
C6811 XA.XIR[2].XIC_15.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Ien 0.00214f
C6812 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C6813 XA.XIR[7].XIC[1].icell.PUM VPWR 0.00937f
C6814 XA.XIR[0].XIC[6].icell.PDM VPWR 0.0078f
C6815 XA.XIR[13].XIC[0].icell.Ien XA.XIR[13].XIC[1].icell.Ien 0.00214f
C6816 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C6817 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.PDM 0.0059f
C6818 XThC.Tn[10] XThR.Tn[3] 0.28739f
C6819 XA.XIR[4].XIC_15.icell.PDM Vbias 0.04401f
C6820 XA.XIR[2].XIC[4].icell.PUM Vbias 0.0031f
C6821 XA.XIR[7].XIC[4].icell.Ien Vbias 0.21098f
C6822 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9] 0.00341f
C6823 XA.XIR[9].XIC[2].icell.PDM Iout 0.00117f
C6824 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11154f
C6825 XThC.Tn[0] XA.XIR[6].XIC_dummy_left.icell.Iout 0.00109f
C6826 XThR.Tn[12] XA.XIR[13].XIC[0].icell.SM 0.00127f
C6827 XA.XIR[9].XIC[10].icell.PUM VPWR 0.00937f
C6828 XA.XIR[10].XIC[2].icell.SM VPWR 0.00158f
C6829 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.Ien 0.00584f
C6830 XA.XIR[1].XIC[6].icell.PUM Vbias 0.0031f
C6831 XThC.Tn[7] VPWR 6.29093f
C6832 XA.XIR[14].XIC[8].icell.SM Vbias 0.00701f
C6833 XA.XIR[15].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.SM 0.0039f
C6834 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C6835 XA.XIR[12].XIC[13].icell.Ien Iout 0.06417f
C6836 XA.XIR[0].XIC[3].icell.PUM VPWR 0.00877f
C6837 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.SM 0.00168f
C6838 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04031f
C6839 XA.XIR[8].XIC[14].icell.PUM Vbias 0.0031f
C6840 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.04036f
C6841 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04031f
C6842 XA.XIR[14].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.SM 0.0039f
C6843 XA.XIR[3].XIC[11].icell.SM VPWR 0.00158f
C6844 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10] 0.00341f
C6845 XThC.Tn[13] XThR.Tn[0] 0.28789f
C6846 XA.XIR[3].XIC_15.icell.SM Vbias 0.00701f
C6847 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C6848 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14] 0.00341f
C6849 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C6850 XA.XIR[3].XIC[7].icell.SM Iout 0.00388f
C6851 XA.XIR[1].XIC[7].icell.PDM Iout 0.00117f
C6852 XA.XIR[2].XIC[4].icell.SM VPWR 0.00158f
C6853 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C6854 XA.XIR[6].XIC[12].icell.Ien Iout 0.06417f
C6855 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C6856 XA.XIR[7].XIC[6].icell.PUM VPWR 0.00937f
C6857 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02762f
C6858 XA.XIR[13].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.SM 0.0039f
C6859 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.03425f
C6860 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C6861 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C6862 XA.XIR[4].XIC[7].icell.PDM Iout 0.00117f
C6863 XA.XIR[1].XIC[6].icell.SM VPWR 0.00158f
C6864 a_5949_10571# VPWR 0.00653f
C6865 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.PDM 0.00591f
C6866 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02827f
C6867 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PUM 0.00465f
C6868 XA.XIR[1].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.SM 0.0039f
C6869 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.Ien 0.00584f
C6870 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C6871 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01451f
C6872 XA.XIR[1].XIC[2].icell.SM Iout 0.00388f
C6873 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02762f
C6874 XA.XIR[3].XIC_15.icell.PDM Iout 0.00133f
C6875 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38997f
C6876 XA.XIR[9].XIC_15.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Ien 0.00214f
C6877 XA.XIR[14].XIC[6].icell.Ien Iout 0.06417f
C6878 XA.XIR[0].XIC_dummy_right.icell.PUM Vbias 0.00223f
C6879 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.Ien 0.00584f
C6880 XA.XIR[8].XIC[14].icell.SM VPWR 0.00207f
C6881 XThC.XTB6.A a_7331_10587# 0.00304f
C6882 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C6883 XA.XIR[12].XIC[14].icell.SM Iout 0.00388f
C6884 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.Ien 0.00584f
C6885 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.15202f
C6886 XA.XIR[5].XIC[0].icell.PDM Vbias 0.04207f
C6887 XThR.XTB7.A a_n1319_5317# 0.0017f
C6888 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04031f
C6889 XA.XIR[13].XIC[8].icell.Ien Iout 0.06417f
C6890 XA.XIR[8].XIC[10].icell.SM Iout 0.00388f
C6891 XThR.Tn[8] XA.XIR[9].XIC[10].icell.SM 0.00121f
C6892 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.03425f
C6893 XA.XIR[6].XIC[1].icell.PUM Vbias 0.0031f
C6894 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C6895 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02762f
C6896 XThR.Tn[2] XA.XIR[3].XIC[5].icell.Ien 0.00338f
C6897 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C6898 XA.XIR[5].XIC[0].icell.PUM VPWR 0.00937f
C6899 XA.XIR[11].XIC[1].icell.Ien XA.XIR[11].XIC[2].icell.Ien 0.00214f
C6900 XThR.Tn[4] XA.XIR[4].XIC[0].icell.PDM 0.00346f
C6901 XThR.Tn[4] XA.XIR[5].XIC[12].icell.Ien 0.00338f
C6902 XThR.XTB3.Y a_n997_3979# 0.00604f
C6903 XThR.XTBN.A XThR.Tn[12] 0.22096f
C6904 XA.XIR[14].XIC_dummy_left.icell.SM VPWR 0.00269f
C6905 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PUM 0.00465f
C6906 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C6907 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PUM 0.00465f
C6908 XThR.Tn[5] XA.XIR[6].XIC_15.icell.PDM 0.00172f
C6909 XThR.Tn[3] XA.XIR[3].XIC[1].icell.PDM 0.00341f
C6910 XThR.Tn[3] XA.XIR[4].XIC[12].icell.Ien 0.00338f
C6911 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.03425f
C6912 a_3773_9615# VPWR 0.70508f
C6913 XThR.Tn[11] XA.XIR[12].XIC[14].icell.Ien 0.00338f
C6914 XThR.Tn[1] XA.XIR[2].XIC[3].icell.SM 0.00121f
C6915 XA.XIR[11].XIC[5].icell.PDM Vbias 0.04261f
C6916 XA.XIR[11].XIC[11].icell.SM Vbias 0.00701f
C6917 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C6918 XThC.Tn[12] XThR.Tn[2] 0.28739f
C6919 XThR.XTB2.Y a_n997_3755# 0.06476f
C6920 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04031f
C6921 XA.XIR[3].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.SM 0.0039f
C6922 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PUM 0.00465f
C6923 XA.XIR[15].XIC[11].icell.SM Iout 0.00388f
C6924 XA.XIR[10].XIC[9].icell.PDM Vbias 0.04261f
C6925 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C6926 XA.XIR[0].XIC[12].icell.SM Iout 0.00367f
C6927 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C6928 XA.XIR[5].XIC[4].icell.PDM VPWR 0.00799f
C6929 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C6930 XThR.Tn[2] XA.XIR[2].XIC[13].icell.PDM 0.00341f
C6931 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C6932 XThC.XTB4.Y a_5155_9615# 0.01546f
C6933 XThR.XTBN.Y a_n1049_8581# 0.0607f
C6934 XThR.Tn[13] XA.XIR[14].XIC[7].icell.SM 0.00121f
C6935 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C6936 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11115f
C6937 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Iout 0.00347f
C6938 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04052f
C6939 XA.XIR[6].XIC[6].icell.PUM Vbias 0.0031f
C6940 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Ien 0.00232f
C6941 XThC.XTB5.Y a_8739_9569# 0.00424f
C6942 XA.XIR[12].XIC[3].icell.PDM VPWR 0.00799f
C6943 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C6944 XA.XIR[15].XIC[7].icell.Ien Vbias 0.17899f
C6945 XA.XIR[2].XIC_15.icell.Ien Iout 0.0642f
C6946 XA.XIR[12].XIC[11].icell.Ien Iout 0.06417f
C6947 XThR.Tn[0] XA.XIR[1].XIC[10].icell.SM 0.00121f
C6948 XA.XIR[5].XIC[7].icell.SM Vbias 0.00701f
C6949 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C6950 XA.XIR[11].XIC[9].icell.PDM VPWR 0.00799f
C6951 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02762f
C6952 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.PUM 0.00121f
C6953 XThR.XTB2.Y a_n1049_5611# 0.00844f
C6954 XA.XIR[7].XIC_dummy_left.icell.Ien Vbias 0.00329f
C6955 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C6956 XA.XIR[4].XIC[10].icell.Ien Vbias 0.21098f
C6957 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PUM 0.00465f
C6958 XA.XIR[14].XIC[0].icell.SM Iout 0.00388f
C6959 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.03425f
C6960 XA.XIR[0].XIC[1].icell.Ien Vbias 0.2113f
C6961 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.SM 0.00168f
C6962 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.03425f
C6963 XA.XIR[2].XIC[1].icell.PDM Vbias 0.04261f
C6964 XThC.Tn[8] XThR.Tn[6] 0.28739f
C6965 XA.XIR[4].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.SM 0.0039f
C6966 XA.XIR[11].XIC[14].icell.PUM Vbias 0.0031f
C6967 XA.XIR[8].XIC[4].icell.Ien Vbias 0.21098f
C6968 XThR.Tn[5] XA.XIR[6].XIC[12].icell.SM 0.00121f
C6969 XA.XIR[3].XIC[3].icell.PUM VPWR 0.00937f
C6970 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.SM 0.00168f
C6971 XA.XIR[10].XIC[1].icell.PDM Iout 0.00117f
C6972 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04031f
C6973 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.0355f
C6974 XA.XIR[6].XIC[6].icell.SM VPWR 0.00158f
C6975 XA.XIR[12].XIC[2].icell.SM Vbias 0.00701f
C6976 XThR.XTB3.Y XThR.Tn[7] 0.00819f
C6977 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C6978 XThR.XTB3.Y a_n997_2891# 0.07285f
C6979 XA.XIR[14].XIC[13].icell.SM Vbias 0.00701f
C6980 XThC.Tn[10] XThR.Tn[11] 0.28739f
C6981 XA.XIR[6].XIC[2].icell.SM Iout 0.00388f
C6982 XA.XIR[15].XIC[9].icell.PUM VPWR 0.00937f
C6983 XA.XIR[11].XIC[5].icell.PUM Vbias 0.0031f
C6984 XA.XIR[5].XIC[9].icell.Ien VPWR 0.1903f
C6985 XThC.XTBN.Y a_8739_9569# 0.22804f
C6986 XA.XIR[9].XIC[13].icell.Ien Vbias 0.21098f
C6987 XThC.Tn[0] XThR.Tn[7] 0.2874f
C6988 XA.XIR[8].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.SM 0.0039f
C6989 XA.XIR[10].XIC[7].icell.PUM Vbias 0.0031f
C6990 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.15222f
C6991 XA.XIR[5].XIC[5].icell.Ien Iout 0.06417f
C6992 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.03425f
C6993 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C6994 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C6995 XA.XIR[8].XIC[1].icell.PDM VPWR 0.00799f
C6996 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C6997 XA.XIR[4].XIC[12].icell.PUM VPWR 0.00937f
C6998 a_n1049_5317# XThR.Tn[6] 0.26047f
C6999 XA.XIR[3].XIC[10].icell.Ien XA.XIR[3].XIC[11].icell.Ien 0.00214f
C7000 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.15202f
C7001 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.15235f
C7002 XA.XIR[2].XIC[5].icell.PDM VPWR 0.00799f
C7003 XA.XIR[0].XIC[6].icell.Ien Vbias 0.21134f
C7004 XThR.Tn[1] a_n1049_7493# 0.00444f
C7005 XA.XIR[13].XIC[2].icell.SM VPWR 0.00158f
C7006 XThC.XTB7.B XThC.Tn[7] 0.08407f
C7007 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C7008 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C7009 XA.XIR[8].XIC[6].icell.PUM VPWR 0.00937f
C7010 XThR.Tn[6] XA.XIR[7].XIC[4].icell.Ien 0.00338f
C7011 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.Ien 0.00584f
C7012 XThC.XTB5.Y XThC.Tn[11] 0.02206f
C7013 XA.XIR[3].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7014 XA.XIR[12].XIC[4].icell.Ien VPWR 0.1903f
C7015 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12] 0.00341f
C7016 XThC.Tn[6] Vbias 2.22871f
C7017 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C7018 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.SM 0.00168f
C7019 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.Ien 0.00256f
C7020 XThR.Tn[5] Iout 1.16233f
C7021 a_8739_9569# XThC.Tn[10] 0.19671f
C7022 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C7023 XA.XIR[11].XIC[5].icell.SM VPWR 0.00158f
C7024 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04031f
C7025 XA.XIR[7].XIC[9].icell.Ien Vbias 0.21098f
C7026 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C7027 XThR.Tn[8] data[4] 0.01643f
C7028 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C7029 XA.XIR[2].XIC[3].icell.Ien XA.XIR[2].XIC[4].icell.Ien 0.00214f
C7030 XA.XIR[2].XIC[9].icell.PUM Vbias 0.0031f
C7031 a_n997_3979# VPWR 0.01662f
C7032 XThR.Tn[11] XA.XIR[12].XIC[12].icell.Ien 0.00338f
C7033 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.SM 0.0039f
C7034 XA.XIR[2].XIC[0].icell.SM Iout 0.00388f
C7035 XThR.Tn[4] XA.XIR[5].XIC[2].icell.SM 0.00121f
C7036 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.03425f
C7037 XA.XIR[11].XIC[9].icell.SM Vbias 0.00701f
C7038 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.04617f
C7039 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01577f
C7040 XThC.Tn[13] XThR.Tn[1] 0.2874f
C7041 XA.XIR[11].XIC[1].icell.SM Iout 0.00388f
C7042 XA.XIR[10].XIC[7].icell.SM VPWR 0.00158f
C7043 XA.XIR[15].XIC[9].icell.SM Iout 0.00388f
C7044 XA.XIR[1].XIC[11].icell.PUM Vbias 0.0031f
C7045 XThR.Tn[3] XA.XIR[4].XIC[2].icell.SM 0.00121f
C7046 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.15202f
C7047 XThR.Tn[14] XA.XIR[15].XIC[4].icell.Ien 0.00338f
C7048 XThR.XTBN.A data[7] 0.07741f
C7049 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.03425f
C7050 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7051 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C7052 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C7053 XThC.XTB2.Y a_5155_9615# 0.00847f
C7054 XA.XIR[10].XIC[3].icell.SM Iout 0.00388f
C7055 XA.XIR[0].XIC[8].icell.PUM VPWR 0.00881f
C7056 XThR.Tn[9] XA.XIR[10].XIC[3].icell.SM 0.00121f
C7057 XA.XIR[1].XIC[5].icell.Ien XA.XIR[1].XIC[6].icell.Ien 0.00214f
C7058 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C7059 XThC.Tn[13] XThR.Tn[12] 0.2874f
C7060 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04031f
C7061 XThR.XTB7.B a_n1319_5317# 0.00108f
C7062 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C7063 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04031f
C7064 XThC.XTB7.A data[2] 0.00198f
C7065 XThC.XTB6.A XThC.XTBN.A 0.0513f
C7066 XA.XIR[2].XIC[0].icell.Ien Vbias 0.20951f
C7067 XThC.XTBN.Y XThC.Tn[11] 0.53369f
C7068 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02762f
C7069 XA.XIR[3].XIC[12].icell.SM Iout 0.00388f
C7070 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.03425f
C7071 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8] 0.00341f
C7072 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04031f
C7073 XThC.Tn[8] XThR.Tn[4] 0.28739f
C7074 a_n1049_7787# XThR.Tn[2] 0.00158f
C7075 XA.XIR[2].XIC[9].icell.SM VPWR 0.00158f
C7076 XA.XIR[0].XIC[8].icell.Ien XA.XIR[0].XIC[8].icell.SM 0.0039f
C7077 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38936f
C7078 XA.XIR[7].XIC[11].icell.PUM VPWR 0.00937f
C7079 XA.XIR[11].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.SM 0.0039f
C7080 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02762f
C7081 XA.XIR[8].XIC[13].icell.Ien XA.XIR[8].XIC[14].icell.Ien 0.00214f
C7082 XA.XIR[1].XIC[11].icell.SM VPWR 0.00158f
C7083 XA.XIR[2].XIC[5].icell.SM Iout 0.00388f
C7084 XA.XIR[10].XIC[1].icell.Ien Vbias 0.21098f
C7085 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04031f
C7086 XA.XIR[7].XIC[1].icell.PDM Vbias 0.04261f
C7087 XA.XIR[5].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.SM 0.0039f
C7088 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.SM 0.00168f
C7089 XThR.Tn[12] XA.XIR[13].XIC[1].icell.SM 0.00121f
C7090 XA.XIR[1].XIC_15.icell.SM Vbias 0.00704f
C7091 XA.XIR[11].XIC[12].icell.PUM Vbias 0.0031f
C7092 XA.XIR[1].XIC[7].icell.SM Iout 0.00388f
C7093 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.SM 0.00168f
C7094 XA.XIR[9].XIC_15.icell.SM Iout 0.0047f
C7095 XThC.Tn[2] XThR.Tn[0] 0.28882f
C7096 XThC.Tn[12] XThR.Tn[10] 0.28739f
C7097 XA.XIR[6].XIC[8].icell.PDM Vbias 0.04261f
C7098 XThC.Tn[4] XThR.Tn[5] 0.28739f
C7099 XA.XIR[15].XIC[14].icell.Ien XA.XIR[15].XIC_15.icell.Ien 0.00214f
C7100 XA.XIR[9].XIC[3].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00214f
C7101 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.15202f
C7102 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.SM 0.0039f
C7103 XA.XIR[8].XIC[1].icell.PUM VPWR 0.00937f
C7104 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PUM 0.00465f
C7105 XA.XIR[14].XIC[5].icell.PDM Vbias 0.04261f
C7106 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.15202f
C7107 XA.XIR[5].XIC_15.icell.PDM Vbias 0.04401f
C7108 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C7109 XA.XIR[14].XIC[11].icell.SM Vbias 0.00701f
C7110 XThC.Tn[10] XThC.Tn[11] 0.09949f
C7111 XThR.Tn[11] XA.XIR[12].XIC[4].icell.SM 0.00121f
C7112 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02762f
C7113 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.SM 0.00168f
C7114 XThC.XTB6.Y a_7875_9569# 0.0046f
C7115 XA.XIR[13].XIC[9].icell.PDM Vbias 0.04261f
C7116 XThR.Tn[2] XA.XIR[3].XIC[10].icell.Ien 0.00338f
C7117 XThR.Tn[7] VPWR 6.97893f
C7118 a_n997_2891# VPWR 0.01347f
C7119 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PUM 0.00465f
C7120 XThR.Tn[4] XA.XIR[4].XIC_15.icell.PDM 0.00341f
C7121 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04031f
C7122 XA.XIR[7].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.SM 0.0039f
C7123 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C7124 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C7125 XA.XIR[7].XIC_15.icell.SM VPWR 0.00275f
C7126 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.03425f
C7127 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.03425f
C7128 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PUM 0.00429f
C7129 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10] 0.00341f
C7130 XA.XIR[7].XIC[5].icell.PDM VPWR 0.00799f
C7131 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.15202f
C7132 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C7133 XA.XIR[9].XIC[3].icell.SM Vbias 0.00701f
C7134 XThR.Tn[1] XA.XIR[2].XIC[8].icell.SM 0.00121f
C7135 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Iout 0.00347f
C7136 XA.XIR[15].XIC[3].icell.PDM VPWR 0.0114f
C7137 XThR.XTB6.Y a_n1049_5317# 0.01199f
C7138 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C7139 XA.XIR[6].XIC[12].icell.PDM VPWR 0.00799f
C7140 XA.XIR[4].XIC[2].icell.Ien VPWR 0.1903f
C7141 XA.XIR[11].XIC[13].icell.Ien Vbias 0.21098f
C7142 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PUM 0.00465f
C7143 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.03425f
C7144 XA.XIR[6].XIC[0].icell.PDM Iout 0.00117f
C7145 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C7146 XA.XIR[14].XIC[9].icell.PDM VPWR 0.00799f
C7147 XA.XIR[15].XIC[13].icell.Ien Iout 0.06807f
C7148 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.03425f
C7149 XA.XIR[5].XIC[7].icell.PDM Iout 0.00117f
C7150 XA.XIR[1].XIC[2].icell.PDM Vbias 0.04261f
C7151 XA.XIR[3].XIC[6].icell.Ien Vbias 0.21098f
C7152 XThR.Tn[11] XA.XIR[12].XIC[10].icell.Ien 0.00338f
C7153 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C7154 XA.XIR[6].XIC[11].icell.PUM Vbias 0.0031f
C7155 XA.XIR[14].XIC[14].icell.PUM Vbias 0.0031f
C7156 XA.XIR[9].XIC[1].icell.PDM VPWR 0.00799f
C7157 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Ien 0.00232f
C7158 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02762f
C7159 XA.XIR[13].XIC[1].icell.PDM Iout 0.00117f
C7160 XThC.Tn[1] XThR.Tn[2] 0.28739f
C7161 XA.XIR[5].XIC[12].icell.SM Vbias 0.00701f
C7162 XA.XIR[3].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.SM 0.0039f
C7163 XA.XIR[4].XIC[2].icell.PDM Vbias 0.04261f
C7164 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.SM 0.00168f
C7165 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.SM 0.00168f
C7166 XA.XIR[5].XIC[12].icell.Ien XA.XIR[5].XIC[13].icell.Ien 0.00214f
C7167 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PUM 0.00465f
C7168 XA.XIR[9].XIC[5].icell.Ien VPWR 0.1903f
C7169 XA.XIR[12].XIC[12].icell.SM VPWR 0.00158f
C7170 XA.XIR[12].XIC[6].icell.PDM Iout 0.00117f
C7171 XA.XIR[4].XIC_15.icell.Ien Vbias 0.21234f
C7172 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.Ien 0.00584f
C7173 XThR.XTB5.A data[5] 0.11096f
C7174 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.SM 0.00168f
C7175 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00584f
C7176 XA.XIR[3].XIC[10].icell.PDM Vbias 0.04261f
C7177 XThC.Tn[10] XThR.Tn[14] 0.28739f
C7178 XThC.XTB4.Y a_7875_9569# 0.00497f
C7179 XA.XIR[8].XIC[12].icell.PDM Vbias 0.04261f
C7180 XA.XIR[14].XIC[5].icell.PUM Vbias 0.0031f
C7181 XA.XIR[1].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.SM 0.0039f
C7182 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02762f
C7183 XThR.XTBN.Y a_n1049_7787# 0.08456f
C7184 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C7185 XThC.XTB1.Y a_3299_10575# 0.0097f
C7186 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C7187 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C7188 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.Ien 0.00584f
C7189 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.04036f
C7190 XA.XIR[13].XIC[7].icell.PUM Vbias 0.0031f
C7191 XThR.XTB7.Y a_n997_3755# 0.00476f
C7192 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C7193 XThR.XTB2.Y data[4] 0.00267f
C7194 XA.XIR[8].XIC[9].icell.Ien Vbias 0.21098f
C7195 XA.XIR[6].XIC[0].icell.Ien XA.XIR[6].XIC[1].icell.Ien 0.00214f
C7196 XA.XIR[3].XIC[8].icell.PUM VPWR 0.00937f
C7197 XA.XIR[11].XIC[14].icell.SM Vbias 0.00701f
C7198 XThC.XTB6.A XThC.Tn[2] 0.00108f
C7199 XA.XIR[1].XIC[6].icell.PDM VPWR 0.00799f
C7200 XThR.Tn[14] XA.XIR[15].XIC[12].icell.SM 0.00121f
C7201 XA.XIR[12].XIC[7].icell.SM Vbias 0.00701f
C7202 XA.XIR[6].XIC[11].icell.SM VPWR 0.00158f
C7203 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02762f
C7204 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.SM 0.00168f
C7205 a_n1049_6405# XThR.Tn[4] 0.26564f
C7206 XA.XIR[6].XIC_15.icell.SM Vbias 0.00701f
C7207 XA.XIR[15].XIC[14].icell.SM Iout 0.00388f
C7208 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C7209 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.15202f
C7210 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7211 a_5155_9615# XThC.Tn[4] 0.26653f
C7212 XA.XIR[11].XIC[10].icell.PUM Vbias 0.0031f
C7213 XA.XIR[4].XIC[6].icell.PDM VPWR 0.00799f
C7214 XA.XIR[6].XIC[7].icell.SM Iout 0.00388f
C7215 XA.XIR[5].XIC[14].icell.Ien VPWR 0.19036f
C7216 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7] 0.00341f
C7217 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04031f
C7218 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.0353f
C7219 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.SM 0.00168f
C7220 XA.XIR[3].XIC[14].icell.PDM VPWR 0.00809f
C7221 XA.XIR[5].XIC[10].icell.Ien Iout 0.06417f
C7222 XA.XIR[1].XIC[3].icell.PUM VPWR 0.00937f
C7223 XA.XIR[14].XIC[5].icell.SM VPWR 0.00158f
C7224 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C7225 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13] 0.00341f
C7226 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.SM 0.00168f
C7227 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.SM 0.00168f
C7228 XA.XIR[14].XIC[9].icell.SM Vbias 0.00701f
C7229 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C7230 XA.XIR[8].XIC[4].icell.PDM Iout 0.00117f
C7231 XA.XIR[3].XIC[2].icell.PDM Iout 0.00117f
C7232 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01577f
C7233 XThC.XTBN.A XThC.Tn[8] 0.1369f
C7234 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.SM 0.00168f
C7235 XA.XIR[0].XIC[11].icell.Ien Vbias 0.2113f
C7236 XThC.Tn[6] XThR.Tn[6] 0.28739f
C7237 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04031f
C7238 XA.XIR[14].XIC[1].icell.SM Iout 0.00388f
C7239 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.Ien 0.00584f
C7240 XA.XIR[13].XIC[7].icell.SM VPWR 0.00158f
C7241 a_n1049_5611# XThR.XTB7.Y 0.00153f
C7242 XA.XIR[12].XIC[7].icell.Ien XA.XIR[12].XIC[8].icell.Ien 0.00214f
C7243 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04031f
C7244 XA.XIR[8].XIC[11].icell.PUM VPWR 0.00937f
C7245 XThR.Tn[6] XA.XIR[7].XIC[9].icell.Ien 0.00338f
C7246 XA.XIR[2].XIC[8].icell.PDM Iout 0.00117f
C7247 XA.XIR[13].XIC[3].icell.SM Iout 0.00388f
C7248 XA.XIR[12].XIC[9].icell.Ien VPWR 0.1903f
C7249 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C7250 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.Ien 0.00584f
C7251 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7252 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02762f
C7253 XThR.Tn[0] XA.XIR[0].XIC[5].icell.PDM 0.00341f
C7254 XA.XIR[12].XIC[5].icell.Ien Iout 0.06417f
C7255 XThR.Tn[14] XA.XIR[15].XIC_15.icell.PUM 0.00186f
C7256 XA.XIR[2].XIC[14].icell.PUM Vbias 0.0031f
C7257 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.SM 0.00168f
C7258 XA.XIR[7].XIC[14].icell.Ien Vbias 0.21098f
C7259 XA.XIR[12].XIC_15.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Ien 0.00214f
C7260 XThR.Tn[4] XA.XIR[5].XIC[7].icell.SM 0.00121f
C7261 XThR.Tn[1] XA.XIR[1].XIC[3].icell.PDM 0.00341f
C7262 XA.XIR[9].XIC[0].icell.Ien VPWR 0.1903f
C7263 XA.XIR[11].XIC[6].icell.SM Iout 0.00388f
C7264 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.Ien 0.00584f
C7265 XA.XIR[11].XIC[11].icell.Ien Vbias 0.21098f
C7266 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C7267 XA.XIR[1].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7268 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.SM 0.00168f
C7269 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04031f
C7270 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.15202f
C7271 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02762f
C7272 XThR.Tn[3] XA.XIR[4].XIC[7].icell.SM 0.00121f
C7273 XThR.Tn[14] XA.XIR[15].XIC[9].icell.Ien 0.00338f
C7274 XA.XIR[10].XIC[8].icell.SM Iout 0.00388f
C7275 XA.XIR[4].XIC[0].icell.SM Vbias 0.00675f
C7276 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02762f
C7277 XThR.Tn[9] XA.XIR[10].XIC[8].icell.SM 0.00121f
C7278 XA.XIR[0].XIC[13].icell.PUM VPWR 0.00877f
C7279 XA.XIR[15].XIC[11].icell.Ien Iout 0.06807f
C7280 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PUM 0.00465f
C7281 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5] 0.00341f
C7282 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.15202f
C7283 XA.XIR[10].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.SM 0.0039f
C7284 XThC.XTB6.Y XThC.Tn[4] 0.00264f
C7285 XA.XIR[13].XIC[1].icell.Ien Vbias 0.21098f
C7286 XThC.XTB7.A a_5949_9615# 0.01824f
C7287 XA.XIR[14].XIC[1].icell.Ien XA.XIR[14].XIC[2].icell.Ien 0.00214f
C7288 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PUM 0.00465f
C7289 XA.XIR[14].XIC[12].icell.PUM Vbias 0.0031f
C7290 XA.XIR[8].XIC_15.icell.SM VPWR 0.00275f
C7291 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.03425f
C7292 XThR.Tn[2] XA.XIR[2].XIC[0].icell.PDM 0.00347f
C7293 XThC.Tn[12] XThR.Tn[13] 0.28739f
C7294 XA.XIR[12].XIC_15.icell.SM Iout 0.0047f
C7295 XA.XIR[6].XIC[5].icell.Ien XA.XIR[6].XIC[6].icell.Ien 0.00214f
C7296 XThC.Tn[2] XThR.Tn[1] 0.28742f
C7297 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04031f
C7298 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C7299 XA.XIR[2].XIC[14].icell.SM VPWR 0.00207f
C7300 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02762f
C7301 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.15202f
C7302 XA.XIR[12].XIC[10].icell.SM VPWR 0.00158f
C7303 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7304 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10] 0.00341f
C7305 XThC.XTB2.Y a_7875_9569# 0.06476f
C7306 XA.XIR[5].XIC[1].icell.PUM VPWR 0.00937f
C7307 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6] 0.00341f
C7308 XA.XIR[2].XIC[10].icell.SM Iout 0.00388f
C7309 XA.XIR[15].XIC[2].icell.SM Vbias 0.00701f
C7310 XA.XIR[5].XIC[4].icell.PUM Vbias 0.0031f
C7311 XThC.Tn[2] XThR.Tn[12] 0.28739f
C7312 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.SM 0.00168f
C7313 XThC.Tn[11] XThR.Tn[8] 0.28739f
C7314 a_n997_1579# VPWR 0.02417f
C7315 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C7316 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.SM 0.00168f
C7317 XThC.XTB5.A XThC.XTB7.A 0.07824f
C7318 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.SM 0.00168f
C7319 XThR.Tn[12] XA.XIR[13].XIC[6].icell.SM 0.00121f
C7320 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C7321 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.Ien 0.00584f
C7322 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.03425f
C7323 XA.XIR[1].XIC[12].icell.SM Iout 0.00388f
C7324 XA.XIR[4].XIC[5].icell.SM Vbias 0.00701f
C7325 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.Ien 0.00584f
C7326 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.SM 0.00168f
C7327 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC[0].icell.Ien 0.00214f
C7328 XThR.Tn[11] XA.XIR[12].XIC_15.icell.Ien 0.00117f
C7329 XThR.XTB3.Y a_n1049_6699# 0.0093f
C7330 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C7331 XThR.Tn[14] XA.XIR[15].XIC[10].icell.SM 0.00121f
C7332 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.15202f
C7333 XThC.XTBN.Y XThC.Tn[0] 0.53577f
C7334 XA.XIR[10].XIC[0].icell.PDM VPWR 0.00799f
C7335 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.03023f
C7336 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C7337 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.Ien 0.00584f
C7338 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.15202f
C7339 XThC.Tn[6] XThR.Tn[4] 0.28739f
C7340 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PUM 0.00465f
C7341 XThR.Tn[2] XA.XIR[3].XIC_15.icell.Ien 0.00117f
C7342 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PUM 0.00465f
C7343 XA.XIR[14].XIC[13].icell.Ien Vbias 0.21098f
C7344 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C7345 XA.XIR[6].XIC[3].icell.PUM VPWR 0.00937f
C7346 XA.XIR[9].XIC[12].icell.PDM Vbias 0.04261f
C7347 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.03425f
C7348 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.SM 0.00168f
C7349 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C7350 XA.XIR[15].XIC[4].icell.Ien VPWR 0.32895f
C7351 XThC.XTB4.Y XThC.Tn[4] 0.00758f
C7352 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C7353 XA.XIR[0].XIC[4].icell.PDM Vbias 0.04271f
C7354 XThC.Tn[1] XThR.Tn[10] 0.28739f
C7355 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02762f
C7356 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.03425f
C7357 XA.XIR[5].XIC[4].icell.SM VPWR 0.00158f
C7358 XA.XIR[12].XIC[13].icell.PUM VPWR 0.00937f
C7359 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.15202f
C7360 XThC.XTB3.Y XThC.Tn[8] 0.00178f
C7361 XA.XIR[11].XIC[13].icell.Ien XA.XIR[11].XIC[14].icell.Ien 0.00214f
C7362 XA.XIR[1].XIC[1].icell.Ien Vbias 0.21104f
C7363 XA.XIR[9].XIC[8].icell.SM Vbias 0.00701f
C7364 XThR.Tn[1] XA.XIR[2].XIC[13].icell.SM 0.00121f
C7365 XA.XIR[10].XIC[2].icell.Ien Vbias 0.21098f
C7366 XA.XIR[7].XIC[8].icell.PDM Iout 0.00117f
C7367 XA.XIR[4].XIC[7].icell.Ien VPWR 0.1903f
C7368 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02762f
C7369 XA.XIR[9].XIC[1].icell.Ien Iout 0.06417f
C7370 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.15202f
C7371 XA.XIR[3].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.SM 0.0039f
C7372 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02823f
C7373 XA.XIR[15].XIC[6].icell.PDM Iout 0.00117f
C7374 XA.XIR[6].XIC_15.icell.PDM Iout 0.00133f
C7375 XA.XIR[0].XIC[1].icell.SM Vbias 0.00716f
C7376 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.PDM 0.00591f
C7377 XThR.XTB7.Y a_n997_715# 0.06874f
C7378 XA.XIR[4].XIC[3].icell.Ien Iout 0.06417f
C7379 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.0343f
C7380 XA.XIR[4].XIC[0].icell.Ien XA.XIR[4].XIC[1].icell.Ien 0.00214f
C7381 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02762f
C7382 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02762f
C7383 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.03425f
C7384 XA.XIR[3].XIC[11].icell.Ien Vbias 0.21098f
C7385 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.Ien 0.00584f
C7386 XA.XIR[6].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7387 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C7388 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C7389 XA.XIR[7].XIC[1].icell.Ien VPWR 0.1903f
C7390 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01093f
C7391 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.SM 0.00168f
C7392 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.15202f
C7393 XA.XIR[2].XIC[4].icell.Ien Vbias 0.21098f
C7394 XThC.XTB5.Y VPWR 1.01191f
C7395 XA.XIR[11].XIC[4].icell.Ien XA.XIR[11].XIC[5].icell.Ien 0.00214f
C7396 XA.XIR[14].XIC[14].icell.SM Vbias 0.00701f
C7397 XA.XIR[7].XIC[4].icell.SM Vbias 0.00701f
C7398 XA.XIR[9].XIC[4].icell.PDM Iout 0.00117f
C7399 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9] 0.00341f
C7400 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02762f
C7401 XA.XIR[9].XIC[10].icell.Ien VPWR 0.1903f
C7402 XA.XIR[10].XIC[4].icell.PUM VPWR 0.00937f
C7403 XA.XIR[1].XIC[6].icell.Ien Vbias 0.21104f
C7404 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PUM 0.00465f
C7405 XA.XIR[14].XIC[10].icell.PUM Vbias 0.0031f
C7406 XA.XIR[9].XIC[6].icell.Ien Iout 0.06417f
C7407 XA.XIR[11].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.SM 0.0039f
C7408 XA.XIR[12].XIC[14].icell.Ien VPWR 0.19036f
C7409 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.15202f
C7410 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.0353f
C7411 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04031f
C7412 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C7413 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18966f
C7414 XA.XIR[10].XIC[6].icell.Ien XA.XIR[10].XIC[7].icell.Ien 0.00214f
C7415 XA.XIR[1].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.SM 0.0039f
C7416 XThR.Tn[4] XA.XIR[5].XIC_15.icell.PDM 0.00172f
C7417 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04031f
C7418 XA.XIR[8].XIC[14].icell.Ien Vbias 0.21098f
C7419 XA.XIR[3].XIC[13].icell.PUM VPWR 0.00937f
C7420 XA.XIR[6].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.SM 0.0039f
C7421 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10] 0.00341f
C7422 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PUM 0.00465f
C7423 XA.XIR[11].XIC_dummy_left.icell.Ien Vbias 0.00329f
C7424 XThR.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.00338f
C7425 XA.XIR[1].XIC[9].icell.PDM Iout 0.00117f
C7426 XA.XIR[6].XIC[12].icell.SM Iout 0.00388f
C7427 XA.XIR[2].XIC[6].icell.PUM VPWR 0.00937f
C7428 XA.XIR[7].XIC[6].icell.Ien VPWR 0.1903f
C7429 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.Ien 0.00584f
C7430 XA.XIR[10].XIC[13].icell.SM Iout 0.00388f
C7431 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.Ien 0.00584f
C7432 XThR.Tn[9] XA.XIR[10].XIC[13].icell.SM 0.00121f
C7433 XA.XIR[9].XIC_dummy_left.icell.SM VPWR 0.00269f
C7434 XA.XIR[15].XIC[2].icell.Ien XA.XIR[15].XIC[3].icell.Ien 0.00214f
C7435 XA.XIR[8].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.SM 0.0039f
C7436 XA.XIR[1].XIC[8].icell.PUM VPWR 0.00937f
C7437 XA.XIR[4].XIC[9].icell.PDM Iout 0.00117f
C7438 XA.XIR[7].XIC[2].icell.Ien Iout 0.06417f
C7439 XA.XIR[5].XIC_15.icell.Ien Iout 0.0642f
C7440 XThC.XTBN.Y VPWR 4.08849f
C7441 XThC.XTB6.Y a_6243_9615# 0.01199f
C7442 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.03425f
C7443 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C7444 a_n1049_6699# VPWR 0.72162f
C7445 XThR.XTB7.A XThR.XTBN.A 0.19736f
C7446 XA.XIR[14].XIC[6].icell.SM Iout 0.00388f
C7447 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C7448 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02762f
C7449 XA.XIR[14].XIC[11].icell.Ien Vbias 0.21098f
C7450 XThR.Tn[7] XA.XIR[8].XIC[3].icell.Ien 0.00338f
C7451 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7452 XA.XIR[12].XIC_15.icell.PDM Iout 0.00133f
C7453 XThR.Tn[6] XA.XIR[7].XIC[14].icell.Ien 0.00338f
C7454 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.Ien 0.00584f
C7455 XA.XIR[14].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.SM 0.0039f
C7456 XA.XIR[13].XIC[8].icell.SM Iout 0.00388f
C7457 XA.XIR[5].XIC[2].icell.PDM Vbias 0.04261f
C7458 XA.XIR[4].XIC[5].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00214f
C7459 XThR.XTB7.A XThR.Tn[6] 0.1056f
C7460 XThC.XTB1.Y XThC.Tn[8] 0.29191f
C7461 XA.XIR[12].XIC[11].icell.PUM VPWR 0.00937f
C7462 XA.XIR[11].XIC[12].icell.Ien XA.XIR[11].XIC[13].icell.Ien 0.00214f
C7463 XA.XIR[6].XIC[1].icell.Ien Vbias 0.21098f
C7464 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10] 0.00341f
C7465 XThR.Tn[2] XA.XIR[3].XIC[5].icell.SM 0.00121f
C7466 XA.XIR[2].XIC[8].icell.Ien XA.XIR[2].XIC[9].icell.Ien 0.00214f
C7467 XThR.Tn[4] XA.XIR[5].XIC[12].icell.SM 0.00121f
C7468 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.15202f
C7469 XThR.Tn[4] XA.XIR[4].XIC[2].icell.PDM 0.00341f
C7470 XThC.Tn[10] VPWR 6.83631f
C7471 XA.XIR[12].XIC[1].icell.PDM Vbias 0.04261f
C7472 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.03425f
C7473 XThR.Tn[2] Vbias 3.74868f
C7474 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.SM 0.0039f
C7475 XThR.Tn[10] XA.XIR[11].XIC[4].icell.Ien 0.00338f
C7476 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C7477 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.03425f
C7478 XThR.Tn[3] XA.XIR[4].XIC[12].icell.SM 0.00121f
C7479 XThR.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.00341f
C7480 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.03425f
C7481 XThC.XTBN.A XThC.Tn[6] 0.00131f
C7482 XA.XIR[11].XIC[7].icell.PDM Vbias 0.04261f
C7483 a_4861_9615# VPWR 0.70525f
C7484 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PUM 0.00465f
C7485 XThR.Tn[9] Iout 1.16233f
C7486 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.SM 0.0039f
C7487 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.15202f
C7488 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C7489 XA.XIR[1].XIC[10].icell.Ien XA.XIR[1].XIC[11].icell.Ien 0.00214f
C7490 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.SM 0.00168f
C7491 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.15202f
C7492 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04031f
C7493 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Ien 0.00584f
C7494 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C7495 XA.XIR[15].XIC[12].icell.SM VPWR 0.00158f
C7496 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PUM 0.0044f
C7497 XA.XIR[5].XIC[6].icell.PDM VPWR 0.00799f
C7498 XThR.Tn[2] XA.XIR[2].XIC_15.icell.PDM 0.00341f
C7499 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.03425f
C7500 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13] 0.00341f
C7501 XThC.XTB4.Y a_6243_9615# 0.00463f
C7502 XA.XIR[3].XIC[1].icell.SM Vbias 0.00701f
C7503 XA.XIR[13].XIC[0].icell.PDM VPWR 0.00799f
C7504 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PUM 0.00465f
C7505 XA.XIR[0].XIC[13].icell.Ien XA.XIR[0].XIC[13].icell.SM 0.0039f
C7506 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.Ien 0.00584f
C7507 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.15202f
C7508 XA.XIR[6].XIC[6].icell.Ien Vbias 0.21098f
C7509 XThC.XTB5.Y a_9827_9569# 0.06458f
C7510 XA.XIR[12].XIC[5].icell.PDM VPWR 0.00799f
C7511 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.SM 0.00168f
C7512 XA.XIR[15].XIC[7].icell.SM Vbias 0.00701f
C7513 XA.XIR[12].XIC[12].icell.Ien VPWR 0.1903f
C7514 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C7515 XA.XIR[5].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.SM 0.0039f
C7516 XA.XIR[5].XIC[9].icell.PUM Vbias 0.0031f
C7517 XThC.XTB7.A a_8739_9569# 0.00342f
C7518 XA.XIR[15].XIC[0].icell.Ien Iout 0.06801f
C7519 XA.XIR[5].XIC[0].icell.SM Iout 0.00388f
C7520 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.SM 0.00168f
C7521 XA.XIR[4].XIC[10].icell.SM Vbias 0.00701f
C7522 XThC.Tn[1] XThR.Tn[13] 0.28739f
C7523 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.03425f
C7524 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.SM 0.00168f
C7525 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02762f
C7526 XA.XIR[0].XIC_dummy_left.icell.Iout Vbias 0.00803f
C7527 XA.XIR[9].XIC[8].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00214f
C7528 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C7529 XA.XIR[2].XIC[3].icell.PDM Vbias 0.04261f
C7530 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PUM 0.00465f
C7531 XA.XIR[8].XIC[1].icell.Ien VPWR 0.1903f
C7532 XThR.XTB3.Y XThR.Tn[8] 0.00178f
C7533 XA.XIR[13].XIC[2].icell.Ien Vbias 0.21098f
C7534 XThR.Tn[14] XA.XIR[15].XIC[12].icell.Ien 0.00338f
C7535 XA.XIR[8].XIC[4].icell.SM Vbias 0.00701f
C7536 XA.XIR[10].XIC[3].icell.PDM Iout 0.00117f
C7537 XA.XIR[3].XIC[3].icell.Ien VPWR 0.1903f
C7538 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04031f
C7539 XA.XIR[10].XIC[11].icell.SM Iout 0.00388f
C7540 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.Ien 0.00584f
C7541 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01577f
C7542 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.Ien 0.00584f
C7543 XThR.Tn[9] XA.XIR[10].XIC[11].icell.SM 0.00121f
C7544 XThC.Tn[4] Iout 0.83918f
C7545 XThC.Tn[4] XThR.Tn[9] 0.28739f
C7546 XA.XIR[12].XIC[4].icell.PUM Vbias 0.0031f
C7547 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02762f
C7548 XA.XIR[6].XIC[8].icell.PUM VPWR 0.00937f
C7549 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.03425f
C7550 XThC.Tn[0] XThR.Tn[8] 0.2874f
C7551 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.Ien 0.00584f
C7552 a_5155_10571# VPWR 0.00653f
C7553 XThR.XTB7.Y a_n997_2667# 0.00474f
C7554 XA.XIR[15].XIC[9].icell.Ien VPWR 0.32895f
C7555 XA.XIR[2].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.SM 0.0039f
C7556 XThR.XTB7.A XThR.Tn[4] 0.02736f
C7557 XA.XIR[11].XIC[5].icell.Ien Vbias 0.21098f
C7558 XA.XIR[5].XIC[9].icell.SM VPWR 0.00158f
C7559 XThC.XTBN.Y a_9827_9569# 0.22873f
C7560 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.15202f
C7561 XA.XIR[15].XIC[5].icell.Ien Iout 0.06807f
C7562 XThR.XTB7.A a_n1049_7493# 0.0127f
C7563 XA.XIR[9].XIC[13].icell.SM Vbias 0.00701f
C7564 XA.XIR[5].XIC[5].icell.SM Iout 0.00388f
C7565 XA.XIR[3].XIC[1].icell.PDM VPWR 0.00799f
C7566 XA.XIR[10].XIC[7].icell.Ien Vbias 0.21098f
C7567 XA.XIR[4].XIC[12].icell.Ien VPWR 0.1903f
C7568 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C7569 XA.XIR[8].XIC[3].icell.PDM VPWR 0.00799f
C7570 XA.XIR[4].XIC_dummy_right.icell.Ien Vbias 0.00288f
C7571 data[1] data[2] 0.01393f
C7572 XA.XIR[2].XIC[7].icell.PDM VPWR 0.00799f
C7573 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.15202f
C7574 XA.XIR[4].XIC[8].icell.Ien Iout 0.06417f
C7575 XA.XIR[0].XIC[6].icell.SM Vbias 0.00716f
C7576 XA.XIR[13].XIC[4].icell.PUM VPWR 0.00937f
C7577 XA.XIR[11].XIC[11].icell.Ien XA.XIR[11].XIC[12].icell.Ien 0.00214f
C7578 XA.XIR[12].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.SM 0.0039f
C7579 XA.XIR[8].XIC[6].icell.Ien VPWR 0.1903f
C7580 XA.XIR[4].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.SM 0.0039f
C7581 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C7582 XThR.Tn[6] XA.XIR[7].XIC[4].icell.SM 0.00121f
C7583 XA.XIR[12].XIC[4].icell.SM VPWR 0.00158f
C7584 XThR.XTBN.Y Vbias 0.01055f
C7585 XA.XIR[11].XIC_15.icell.SM Vbias 0.00701f
C7586 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12] 0.00341f
C7587 XA.XIR[8].XIC[2].icell.Ien Iout 0.06417f
C7588 XThR.Tn[8] XA.XIR[9].XIC[2].icell.Ien 0.00338f
C7589 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PUM 0.00465f
C7590 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.SM 0.00168f
C7591 XA.XIR[11].XIC[7].icell.PUM VPWR 0.00937f
C7592 XA.XIR[2].XIC[9].icell.Ien Vbias 0.21098f
C7593 XA.XIR[15].XIC_15.icell.SM Iout 0.0047f
C7594 XThC.XTB3.Y XThC.Tn[6] 0.00301f
C7595 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04031f
C7596 XA.XIR[7].XIC[9].icell.SM Vbias 0.00701f
C7597 XA.XIR[7].XIC[4].icell.Ien XA.XIR[7].XIC[5].icell.Ien 0.00214f
C7598 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C7599 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.Ien 0.00256f
C7600 XA.XIR[9].XIC_15.icell.Ien VPWR 0.25566f
C7601 XA.XIR[10].XIC[9].icell.PUM VPWR 0.00937f
C7602 XA.XIR[1].XIC[11].icell.Ien Vbias 0.21104f
C7603 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.Ien 0.00584f
C7604 XA.XIR[15].XIC[10].icell.SM VPWR 0.00158f
C7605 XThC.Tn[3] XThC.Tn[5] 0.00492f
C7606 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C7607 XThR.Tn[14] XA.XIR[15].XIC[4].icell.SM 0.00121f
C7608 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C7609 XThR.XTB7.B XThR.XTBN.A 0.35142f
C7610 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C7611 XA.XIR[13].XIC[13].icell.SM Iout 0.00388f
C7612 XA.XIR[9].XIC[11].icell.Ien Iout 0.06417f
C7613 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C7614 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.15202f
C7615 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.SM 0.00168f
C7616 XThC.XTB2.Y a_6243_9615# 0.00844f
C7617 XA.XIR[0].XIC[8].icell.Ien VPWR 0.19149f
C7618 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C7619 XA.XIR[9].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.SM 0.0039f
C7620 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.SM 0.00168f
C7621 XA.XIR[12].XIC[14].icell.PDM Iout 0.00117f
C7622 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PUM 0.00465f
C7623 XThR.XTB7.B XThR.Tn[6] 0.04822f
C7624 XA.XIR[0].XIC[4].icell.Ien Iout 0.06389f
C7625 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04031f
C7626 XThR.Tn[10] XA.XIR[11].XIC[12].icell.SM 0.00121f
C7627 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C7628 XA.XIR[6].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.SM 0.0039f
C7629 XA.XIR[12].XIC[10].icell.Ien VPWR 0.1903f
C7630 XThC.XTB3.Y a_4387_10575# 0.00941f
C7631 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PUM 0.00465f
C7632 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10] 0.00341f
C7633 XA.XIR[15].XIC_15.icell.PDM Iout 0.00133f
C7634 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8] 0.00341f
C7635 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04031f
C7636 XA.XIR[2].XIC[11].icell.PUM VPWR 0.00937f
C7637 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PUM 0.00465f
C7638 XA.XIR[7].XIC[11].icell.Ien VPWR 0.1903f
C7639 XA.XIR[11].XIC[1].icell.PUM Vbias 0.0031f
C7640 XA.XIR[13].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.SM 0.0039f
C7641 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.SM 0.00168f
C7642 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C7643 XThC.Tn[12] XThR.Tn[7] 0.28739f
C7644 XA.XIR[1].XIC[13].icell.PUM VPWR 0.00937f
C7645 XA.XIR[7].XIC[7].icell.Ien Iout 0.06417f
C7646 XThR.Tn[0] XA.XIR[1].XIC[2].icell.Ien 0.00338f
C7647 XThR.Tn[10] Vbias 3.7463f
C7648 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04031f
C7649 XA.XIR[7].XIC[3].icell.PDM Vbias 0.04261f
C7650 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02762f
C7651 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C7652 XThC.XTB7.B XThC.Tn[10] 0.14845f
C7653 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.SM 0.00168f
C7654 XThR.Tn[14] XA.XIR[15].XIC[10].icell.Ien 0.00338f
C7655 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C7656 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C7657 XA.XIR[10].XIC[9].icell.SM Iout 0.00388f
C7658 XA.XIR[15].XIC[1].icell.PDM Vbias 0.04261f
C7659 XA.XIR[6].XIC[10].icell.PDM Vbias 0.04261f
C7660 XA.XIR[15].XIC[13].icell.PUM VPWR 0.00937f
C7661 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C7662 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Iout 0.00347f
C7663 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.Ien 0.00584f
C7664 XThR.Tn[9] XA.XIR[10].XIC[9].icell.SM 0.00121f
C7665 XThC.Tn[9] Vbias 2.3038f
C7666 XA.XIR[3].XIC[0].icell.Ien VPWR 0.1903f
C7667 XThR.Tn[7] XA.XIR[8].XIC[8].icell.Ien 0.00338f
C7668 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.15202f
C7669 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C7670 XThC.XTB7.B a_4861_9615# 0.0036f
C7671 XThR.Tn[8] VPWR 7.51456f
C7672 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02762f
C7673 XA.XIR[14].XIC[7].icell.PDM Vbias 0.04261f
C7674 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.03425f
C7675 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13] 0.00341f
C7676 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.SM 0.00168f
C7677 XThR.Tn[5] XA.XIR[6].XIC[4].icell.Ien 0.00338f
C7678 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C7679 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C7680 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C7681 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02762f
C7682 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C7683 XThC.XTB6.Y a_8963_9569# 0.00468f
C7684 XThR.Tn[10] XA.XIR[11].XIC_15.icell.PUM 0.00186f
C7685 XThR.Tn[2] XA.XIR[3].XIC[10].icell.SM 0.00121f
C7686 XA.XIR[11].XIC[1].icell.Ien VPWR 0.1903f
C7687 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.15202f
C7688 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04031f
C7689 XA.XIR[2].XIC_15.icell.SM VPWR 0.00275f
C7690 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.03023f
C7691 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.03529f
C7692 XA.XIR[7].XIC[7].icell.PDM VPWR 0.00799f
C7693 XThR.Tn[10] XA.XIR[11].XIC[9].icell.Ien 0.00338f
C7694 XThC.XTB7.A data[1] 0.06544f
C7695 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.Ien 0.00584f
C7696 XA.XIR[9].XIC[0].icell.SM VPWR 0.00158f
C7697 XThR.XTB3.Y a_n997_3755# 0.0061f
C7698 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C7699 a_3773_9615# XThC.Tn[1] 0.27139f
C7700 XA.XIR[9].XIC[5].icell.PUM Vbias 0.0031f
C7701 XA.XIR[11].XIC[10].icell.Ien XA.XIR[11].XIC[11].icell.Ien 0.00214f
C7702 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC[0].icell.Ien 0.00214f
C7703 XThR.Tn[14] a_n997_715# 0.1927f
C7704 XA.XIR[4].XIC[2].icell.SM VPWR 0.00158f
C7705 XA.XIR[6].XIC[14].icell.PDM VPWR 0.00809f
C7706 XA.XIR[15].XIC[5].icell.PDM VPWR 0.0114f
C7707 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.15202f
C7708 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.Ien 0.00584f
C7709 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.03425f
C7710 XThR.Tn[11] a_n997_2667# 0.19413f
C7711 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.15202f
C7712 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C7713 XA.XIR[6].XIC[2].icell.PDM Iout 0.00117f
C7714 XThC.Tn[11] XThR.Tn[3] 0.28739f
C7715 XA.XIR[10].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.SM 0.0039f
C7716 XA.XIR[15].XIC[14].icell.Ien VPWR 0.329f
C7717 XA.XIR[6].XIC[10].icell.Ien XA.XIR[6].XIC[11].icell.Ien 0.00214f
C7718 XA.XIR[3].XIC[6].icell.SM Vbias 0.00701f
C7719 XA.XIR[14].XIC[13].icell.Ien XA.XIR[14].XIC[14].icell.Ien 0.00214f
C7720 XA.XIR[1].XIC[4].icell.PDM Vbias 0.04261f
C7721 XA.XIR[5].XIC[9].icell.PDM Iout 0.00117f
C7722 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01757f
C7723 XA.XIR[6].XIC[11].icell.Ien Vbias 0.21098f
C7724 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.15202f
C7725 XThR.XTB7.B XThR.Tn[4] 0.00356f
C7726 XA.XIR[0].XIC[1].icell.Ien XA.XIR[0].XIC[2].icell.Ien 0.00214f
C7727 a_7651_9569# VPWR 0.00385f
C7728 XA.XIR[9].XIC[3].icell.PDM VPWR 0.00799f
C7729 XA.XIR[13].XIC[3].icell.PDM Iout 0.00117f
C7730 XA.XIR[13].XIC[11].icell.SM Iout 0.00388f
C7731 XA.XIR[4].XIC[4].icell.PDM Vbias 0.04261f
C7732 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.SM 0.00168f
C7733 XA.XIR[11].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.SM 0.0039f
C7734 XA.XIR[5].XIC[14].icell.PUM Vbias 0.0031f
C7735 XThR.XTB3.Y a_n1049_5611# 0.009f
C7736 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C7737 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C7738 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PUM 0.00465f
C7739 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.SM 0.00168f
C7740 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.03425f
C7741 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PUM 0.00102f
C7742 XA.XIR[12].XIC[8].icell.PDM Iout 0.00117f
C7743 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02787f
C7744 XA.XIR[9].XIC[5].icell.SM VPWR 0.00158f
C7745 XA.XIR[1].XIC[1].icell.SM Vbias 0.00704f
C7746 XA.XIR[3].XIC[12].icell.PDM Vbias 0.04261f
C7747 XThC.Tn[14] XThR.Tn[0] 0.28766f
C7748 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.Ien 0.00584f
C7749 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C7750 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C7751 XA.XIR[14].XIC[5].icell.Ien Vbias 0.21098f
C7752 XA.XIR[8].XIC[14].icell.PDM Vbias 0.04261f
C7753 XThC.XTB4.Y a_8963_9569# 0.07199f
C7754 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C7755 XThR.Tn[10] XA.XIR[11].XIC[10].icell.SM 0.00121f
C7756 XA.XIR[9].XIC[1].icell.SM Iout 0.00388f
C7757 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C7758 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02762f
C7759 XA.XIR[10].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.SM 0.0039f
C7760 XA.XIR[13].XIC[7].icell.Ien Vbias 0.21098f
C7761 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.SM 0.00168f
C7762 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.SM 0.00168f
C7763 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04031f
C7764 XA.XIR[14].XIC[4].icell.Ien XA.XIR[14].XIC[5].icell.Ien 0.00214f
C7765 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C7766 XA.XIR[8].XIC[9].icell.SM Vbias 0.00701f
C7767 XThR.Tn[11] XA.XIR[12].XIC[0].icell.Ien 0.0037f
C7768 XA.XIR[3].XIC[8].icell.Ien VPWR 0.1903f
C7769 XA.XIR[11].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7770 XA.XIR[1].XIC[8].icell.PDM VPWR 0.00799f
C7771 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C7772 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PUM 0.00465f
C7773 XA.XIR[12].XIC[9].icell.PUM Vbias 0.0031f
C7774 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C7775 XA.XIR[6].XIC[13].icell.PUM VPWR 0.00937f
C7776 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.SM 0.00168f
C7777 XA.XIR[10].XIC[13].icell.Ien Iout 0.06417f
C7778 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Iout 0.00347f
C7779 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C7780 XThR.Tn[9] XA.XIR[10].XIC[13].icell.Ien 0.00338f
C7781 XA.XIR[3].XIC[4].icell.Ien Iout 0.06417f
C7782 XA.XIR[14].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.SM 0.0039f
C7783 XA.XIR[4].XIC[8].icell.PDM VPWR 0.00799f
C7784 XA.XIR[5].XIC[14].icell.SM VPWR 0.00207f
C7785 XA.XIR[7].XIC[1].icell.SM VPWR 0.00158f
C7786 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7] 0.00341f
C7787 XA.XIR[13].XIC[6].icell.Ien XA.XIR[13].XIC[7].icell.Ien 0.00214f
C7788 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C7789 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04031f
C7790 XA.XIR[14].XIC_15.icell.SM Vbias 0.00701f
C7791 XA.XIR[15].XIC[11].icell.PUM VPWR 0.00937f
C7792 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C7793 XA.XIR[5].XIC_15.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Ien 0.00214f
C7794 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C7795 XA.XIR[1].XIC[3].icell.Ien VPWR 0.1903f
C7796 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C7797 XA.XIR[5].XIC[10].icell.SM Iout 0.00388f
C7798 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02762f
C7799 XThC.XTB7.Y a_6243_10571# 0.01283f
C7800 XA.XIR[14].XIC[7].icell.PUM VPWR 0.00937f
C7801 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C7802 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13] 0.00341f
C7803 a_n1049_7493# XThR.Tn[2] 0.26564f
C7804 XA.XIR[3].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.SM 0.0039f
C7805 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C7806 XA.XIR[12].XIC[13].icell.PDM Iout 0.00117f
C7807 XThR.XTBN.Y XThR.Tn[6] 0.59882f
C7808 XA.XIR[3].XIC[4].icell.PDM Iout 0.00117f
C7809 XA.XIR[8].XIC[6].icell.PDM Iout 0.00117f
C7810 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C7811 XA.XIR[0].XIC[11].icell.SM Vbias 0.00716f
C7812 XA.XIR[4].XIC[13].icell.Ien Iout 0.06417f
C7813 XA.XIR[12].XIC_15.icell.Ien VPWR 0.25566f
C7814 XA.XIR[13].XIC[9].icell.PUM VPWR 0.00937f
C7815 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04031f
C7816 XA.XIR[8].XIC[11].icell.Ien VPWR 0.1903f
C7817 XA.XIR[2].XIC[10].icell.PDM Iout 0.00117f
C7818 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C7819 XThR.Tn[6] XA.XIR[7].XIC[9].icell.SM 0.00121f
C7820 XA.XIR[4].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.SM 0.0039f
C7821 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.SM 0.00168f
C7822 XA.XIR[8].XIC[7].icell.Ien Iout 0.06417f
C7823 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10] 0.00341f
C7824 XThR.Tn[8] XA.XIR[9].XIC[7].icell.Ien 0.00338f
C7825 XA.XIR[15].XIC[14].icell.PDM Iout 0.00117f
C7826 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C7827 XThC.XTB5.A data[1] 0.11102f
C7828 XA.XIR[12].XIC[5].icell.SM Iout 0.00388f
C7829 XThR.Tn[0] XA.XIR[0].XIC[7].icell.PDM 0.00341f
C7830 XA.XIR[2].XIC[14].icell.Ien Vbias 0.21098f
C7831 XThC.Tn[13] XThR.Tn[2] 0.2874f
C7832 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C7833 XA.XIR[2].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.SM 0.0039f
C7834 XA.XIR[7].XIC[14].icell.SM Vbias 0.00701f
C7835 XThR.Tn[14] XA.XIR[15].XIC_15.icell.Ien 0.00117f
C7836 XThR.Tn[1] XA.XIR[1].XIC[5].icell.PDM 0.00341f
C7837 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Ien 0.00584f
C7838 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Ien 0.00584f
C7839 XA.XIR[10].XIC[14].icell.SM Iout 0.00388f
C7840 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C7841 XThR.Tn[9] XA.XIR[10].XIC[14].icell.SM 0.00121f
C7842 XThR.XTB2.Y VPWR 0.98845f
C7843 a_n997_3755# VPWR 0.0133f
C7844 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04031f
C7845 XA.XIR[14].XIC[0].icell.Ien Vbias 0.20951f
C7846 XA.XIR[9].XIC_dummy_right.icell.SM VPWR 0.00123f
C7847 XThC.Tn[0] XA.XIR[7].XIC_dummy_left.icell.Iout 0.00109f
C7848 XA.XIR[10].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.SM 0.0039f
C7849 XA.XIR[4].XIC[2].icell.PUM Vbias 0.0031f
C7850 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C7851 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02762f
C7852 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.03425f
C7853 XA.XIR[15].XIC[12].icell.Ien VPWR 0.32895f
C7854 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18966f
C7855 XA.XIR[1].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.SM 0.0039f
C7856 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C7857 XA.XIR[3].XIC_dummy_left.icell.SM VPWR 0.00269f
C7858 XThR.XTB4.Y XThR.Tn[6] 0.00605f
C7859 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5] 0.00341f
C7860 XA.XIR[14].XIC[12].icell.Ien XA.XIR[14].XIC[13].icell.Ien 0.00214f
C7861 XThR.Tn[13] Vbias 3.74874f
C7862 VPWR data[2] 0.21031f
C7863 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02762f
C7864 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13] 0.00341f
C7865 XThR.XTBN.A XThR.Tn[10] 0.12147f
C7866 XA.XIR[0].XIC[9].icell.Ien Iout 0.06389f
C7867 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.03425f
C7868 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.15202f
C7869 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.15202f
C7870 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C7871 XThR.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.00341f
C7872 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PUM 0.00465f
C7873 XA.XIR[13].XIC[9].icell.SM Iout 0.00388f
C7874 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02762f
C7875 XThR.Tn[13] XA.XIR[14].XIC[4].icell.Ien 0.00338f
C7876 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04031f
C7877 XThR.Tn[10] XA.XIR[11].XIC[14].icell.Ien 0.00338f
C7878 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02762f
C7879 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.SM 0.00168f
C7880 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C7881 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02762f
C7882 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.Ien 0.00584f
C7883 XA.XIR[6].XIC[1].icell.SM Vbias 0.00701f
C7884 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C7885 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.15202f
C7886 a_n1049_5611# VPWR 0.71817f
C7887 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6] 0.00341f
C7888 XA.XIR[15].XIC[4].icell.PUM Vbias 0.0031f
C7889 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.Ien 0.00584f
C7890 XA.XIR[15].XIC[7].icell.Ien XA.XIR[15].XIC[8].icell.Ien 0.00214f
C7891 XThC.XTB2.Y data[0] 0.00267f
C7892 XA.XIR[7].XIC[12].icell.Ien Iout 0.06417f
C7893 XThR.Tn[0] XA.XIR[1].XIC[7].icell.Ien 0.00338f
C7894 XThC.Tn[9] XThR.Tn[6] 0.28739f
C7895 XA.XIR[5].XIC[4].icell.Ien Vbias 0.21098f
C7896 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C7897 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C7898 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.SM 0.0039f
C7899 XA.XIR[14].XIC[1].icell.Ien VPWR 0.19084f
C7900 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PUM 0.0047f
C7901 XA.XIR[4].XIC[7].icell.PUM Vbias 0.0031f
C7902 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C7903 XThR.Tn[7] XA.XIR[8].XIC[13].icell.Ien 0.00338f
C7904 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PUM 0.00465f
C7905 XA.XIR[9].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.SM 0.0039f
C7906 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.Ien 0.00584f
C7907 XA.XIR[10].XIC[2].icell.PDM VPWR 0.00799f
C7908 XA.XIR[15].XIC_15.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Ien 0.00214f
C7909 XA.XIR[10].XIC[11].icell.Ien Iout 0.06417f
C7910 XThC.Tn[11] XThR.Tn[11] 0.28739f
C7911 XA.XIR[4].XIC[10].icell.Ien XA.XIR[4].XIC[11].icell.Ien 0.00214f
C7912 XThR.Tn[9] XA.XIR[10].XIC[11].icell.Ien 0.00338f
C7913 XThR.Tn[5] XA.XIR[6].XIC[9].icell.Ien 0.00338f
C7914 XA.XIR[3].XIC[1].icell.Ien Iout 0.06417f
C7915 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C7916 XThR.XTBN.Y XThR.Tn[4] 0.60351f
C7917 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.03425f
C7918 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC[0].icell.Ien 0.00214f
C7919 XThC.Tn[1] XThR.Tn[7] 0.28739f
C7920 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C7921 XA.XIR[6].XIC[3].icell.Ien VPWR 0.1903f
C7922 XA.XIR[2].XIC[13].icell.Ien XA.XIR[2].XIC[14].icell.Ien 0.00214f
C7923 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.SM 0.00168f
C7924 XA.XIR[9].XIC[14].icell.PDM Vbias 0.04261f
C7925 XThR.XTBN.Y a_n1049_7493# 0.08456f
C7926 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C7927 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C7928 XA.XIR[15].XIC[4].icell.SM VPWR 0.00158f
C7929 XA.XIR[7].XIC[1].icell.PUM Vbias 0.0031f
C7930 XA.XIR[0].XIC[6].icell.PDM Vbias 0.04282f
C7931 XA.XIR[5].XIC[6].icell.PUM VPWR 0.00937f
C7932 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Ien 0.00618f
C7933 XThC.XTB7.B a_7651_9569# 0.01152f
C7934 XA.XIR[9].XIC[10].icell.PUM Vbias 0.0031f
C7935 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PUM 0.00465f
C7936 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C7937 XA.XIR[10].XIC[2].icell.SM Vbias 0.00701f
C7938 XThC.XTB5.Y XThC.Tn[12] 0.32495f
C7939 XA.XIR[4].XIC[7].icell.SM VPWR 0.00158f
C7940 XThR.Tn[1] XA.XIR[2].XIC_15.icell.PUM 0.00186f
C7941 XA.XIR[8].XIC[4].icell.Ien XA.XIR[8].XIC[5].icell.Ien 0.00214f
C7942 XA.XIR[7].XIC[10].icell.PDM Iout 0.00117f
C7943 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.0353f
C7944 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PUM 0.00465f
C7945 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.Ien 0.00584f
C7946 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.04041f
C7947 XThC.Tn[7] Vbias 2.28836f
C7948 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PUM 0.00465f
C7949 XThC.Tn[2] XA.XIR[0].XIC[4].icell.PDM 0.00353f
C7950 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.15202f
C7951 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C7952 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C7953 XA.XIR[15].XIC[8].icell.PDM Iout 0.00117f
C7954 XA.XIR[0].XIC[3].icell.PUM Vbias 0.0031f
C7955 XA.XIR[4].XIC[3].icell.SM Iout 0.00388f
C7956 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Iout 0.00347f
C7957 XA.XIR[8].XIC[1].icell.SM VPWR 0.00158f
C7958 XA.XIR[3].XIC[11].icell.SM Vbias 0.00701f
C7959 XThC.Tn[14] XThR.Tn[1] 0.28745f
C7960 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C7961 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.03425f
C7962 XThR.XTB4.Y XThR.Tn[4] 0.00757f
C7963 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C7964 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.Ien 0.00584f
C7965 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02762f
C7966 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.Ien 0.00584f
C7967 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.1106f
C7968 XA.XIR[2].XIC[1].icell.Ien VPWR 0.1903f
C7969 XThR.XTBN.Y XA.XIR[10].XIC_dummy_left.icell.Iout 0.00376f
C7970 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C7971 XA.XIR[0].XIC[10].icell.PDM VPWR 0.00774f
C7972 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C7973 XA.XIR[11].XIC[2].icell.Ien VPWR 0.1903f
C7974 XA.XIR[10].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.SM 0.0039f
C7975 XA.XIR[2].XIC[4].icell.SM Vbias 0.00701f
C7976 XA.XIR[14].XIC_dummy_right.icell.PUM Vbias 0.00223f
C7977 XA.XIR[15].XIC[10].icell.Ien VPWR 0.32895f
C7978 XA.XIR[7].XIC[6].icell.PUM Vbias 0.0031f
C7979 XThC.Tn[14] XThR.Tn[12] 0.28745f
C7980 XA.XIR[9].XIC[6].icell.PDM Iout 0.00117f
C7981 XA.XIR[7].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.SM 0.0039f
C7982 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9] 0.00341f
C7983 XA.XIR[13].XIC[13].icell.Ien Iout 0.06417f
C7984 XA.XIR[14].XIC[11].icell.Ien XA.XIR[14].XIC[12].icell.Ien 0.00214f
C7985 XA.XIR[9].XIC[10].icell.SM VPWR 0.00158f
C7986 XThC.XTB7.A VPWR 0.87301f
C7987 XA.XIR[10].XIC[4].icell.Ien VPWR 0.1903f
C7988 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11] 0.00341f
C7989 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PUM 0.00465f
C7990 XA.XIR[1].XIC[6].icell.SM Vbias 0.00704f
C7991 XThC.Tn[0] XThR.Tn[3] 0.28747f
C7992 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.SM 0.00168f
C7993 XA.XIR[12].XIC[12].icell.PDM Iout 0.00117f
C7994 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.03425f
C7995 data[7] VGND 0.49949f
C7996 data[6] VGND 0.47974f
C7997 data[4] VGND 0.59317f
C7998 data[5] VGND 1.17814f
C7999 Iout VGND 0.32054p
C8000 bias[2] VGND 0.8011f
C8001 bias[0] VGND 2.64942f
C8002 Vbias VGND 0.23088p
C8003 bias[1] VGND 0.72457f
C8004 data[3] VGND 0.49912f
C8005 data[2] VGND 0.48064f
C8006 data[0] VGND 0.59421f
C8007 data[1] VGND 1.17844f
C8008 VPWR VGND 0.34092p
C8009 a_n997_715# VGND 0.5638f
C8010 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C8011 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C8012 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64514f
C8013 XA.XIR[15].XIC_15.icell.SM VGND 0.00474f
C8014 XA.XIR[15].XIC_dummy_right.icell.PUM VGND 0.00215f
C8015 XA.XIR[15].XIC_15.icell.Ien VGND 0.44292f
C8016 XA.XIR[15].XIC[14].icell.SM VGND 0.00502f
C8017 XA.XIR[15].XIC_15.icell.PUM VGND 0.00282f
C8018 XA.XIR[15].XIC[14].icell.Ien VGND 0.44322f
C8019 XA.XIR[15].XIC[13].icell.SM VGND 0.00502f
C8020 XA.XIR[15].XIC[14].icell.PUM VGND 0.00293f
C8021 XA.XIR[15].XIC[13].icell.Ien VGND 0.44322f
C8022 XA.XIR[15].XIC[12].icell.SM VGND 0.00502f
C8023 XA.XIR[15].XIC[13].icell.PUM VGND 0.00293f
C8024 XA.XIR[15].XIC[12].icell.Ien VGND 0.44322f
C8025 XA.XIR[15].XIC[11].icell.SM VGND 0.00502f
C8026 XA.XIR[15].XIC[12].icell.PUM VGND 0.00293f
C8027 XA.XIR[15].XIC[11].icell.Ien VGND 0.44322f
C8028 XA.XIR[15].XIC[10].icell.SM VGND 0.00502f
C8029 XA.XIR[15].XIC[11].icell.PUM VGND 0.00293f
C8030 XA.XIR[15].XIC[10].icell.Ien VGND 0.44322f
C8031 XA.XIR[15].XIC[9].icell.SM VGND 0.00502f
C8032 XA.XIR[15].XIC[10].icell.PUM VGND 0.00293f
C8033 XA.XIR[15].XIC[9].icell.Ien VGND 0.44322f
C8034 XA.XIR[15].XIC[8].icell.SM VGND 0.00502f
C8035 XA.XIR[15].XIC[9].icell.PUM VGND 0.00293f
C8036 XA.XIR[15].XIC[8].icell.Ien VGND 0.44322f
C8037 XA.XIR[15].XIC[7].icell.SM VGND 0.00502f
C8038 XA.XIR[15].XIC[8].icell.PUM VGND 0.00293f
C8039 XA.XIR[15].XIC[7].icell.Ien VGND 0.44322f
C8040 XA.XIR[15].XIC[6].icell.SM VGND 0.00502f
C8041 XA.XIR[15].XIC[7].icell.PUM VGND 0.00293f
C8042 XA.XIR[15].XIC[6].icell.Ien VGND 0.44322f
C8043 XA.XIR[15].XIC[5].icell.SM VGND 0.00502f
C8044 XA.XIR[15].XIC[6].icell.PUM VGND 0.00293f
C8045 XA.XIR[15].XIC[5].icell.Ien VGND 0.44322f
C8046 XA.XIR[15].XIC[4].icell.SM VGND 0.00502f
C8047 XA.XIR[15].XIC[5].icell.PUM VGND 0.00293f
C8048 XA.XIR[15].XIC[4].icell.Ien VGND 0.44322f
C8049 XA.XIR[15].XIC[3].icell.SM VGND 0.00502f
C8050 XA.XIR[15].XIC[4].icell.PUM VGND 0.00293f
C8051 XA.XIR[15].XIC[3].icell.Ien VGND 0.44322f
C8052 XA.XIR[15].XIC[2].icell.SM VGND 0.00502f
C8053 XA.XIR[15].XIC[3].icell.PUM VGND 0.00293f
C8054 XA.XIR[15].XIC[2].icell.Ien VGND 0.44322f
C8055 XA.XIR[15].XIC[1].icell.SM VGND 0.00502f
C8056 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70718f
C8057 XA.XIR[15].XIC[2].icell.PUM VGND 0.00293f
C8058 XA.XIR[15].XIC[1].icell.Ien VGND 0.44322f
C8059 XA.XIR[15].XIC[0].icell.SM VGND 0.00502f
C8060 XA.XIR[15].XIC[1].icell.PUM VGND 0.00293f
C8061 XA.XIR[15].XIC[0].icell.Ien VGND 0.44356f
C8062 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01044f
C8063 XA.XIR[15].XIC[0].icell.PUM VGND 0.00516f
C8064 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.61163f
C8065 XA.XIR[15].XIC_dummy_left.icell.PUM VGND 0.00215f
C8066 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C8067 XA.XIR[15].XIC_15.icell.PDM VGND 0.18779f
C8068 XA.XIR[15].XIC[14].icell.PDM VGND 0.18733f
C8069 XA.XIR[15].XIC[13].icell.PDM VGND 0.18733f
C8070 XA.XIR[15].XIC[12].icell.PDM VGND 0.18733f
C8071 XA.XIR[15].XIC[11].icell.PDM VGND 0.18733f
C8072 XA.XIR[15].XIC[10].icell.PDM VGND 0.18733f
C8073 XA.XIR[15].XIC[9].icell.PDM VGND 0.18733f
C8074 XA.XIR[15].XIC[8].icell.PDM VGND 0.18733f
C8075 XA.XIR[15].XIC[7].icell.PDM VGND 0.18733f
C8076 XA.XIR[15].XIC[6].icell.PDM VGND 0.18733f
C8077 XA.XIR[15].XIC[5].icell.PDM VGND 0.18733f
C8078 XA.XIR[15].XIC[4].icell.PDM VGND 0.18733f
C8079 XA.XIR[15].XIC[3].icell.PDM VGND 0.18733f
C8080 XA.XIR[15].XIC[2].icell.PDM VGND 0.18733f
C8081 XA.XIR[15].XIC[1].icell.PDM VGND 0.18733f
C8082 XA.XIR[15].XIC[0].icell.PDM VGND 0.18741f
C8083 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C8084 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C8085 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C8086 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.608f
C8087 XA.XIR[14].XIC_15.icell.SM VGND 0.00474f
C8088 XA.XIR[14].XIC_dummy_right.icell.PUM VGND 0.00215f
C8089 XA.XIR[14].XIC_15.icell.Ien VGND 0.37063f
C8090 XA.XIR[14].XIC[14].icell.SM VGND 0.00502f
C8091 XA.XIR[14].XIC_15.icell.PUM VGND 0.00282f
C8092 XA.XIR[14].XIC[14].icell.Ien VGND 0.37144f
C8093 XA.XIR[14].XIC[13].icell.SM VGND 0.00502f
C8094 XA.XIR[14].XIC[14].icell.PUM VGND 0.00293f
C8095 XA.XIR[14].XIC[13].icell.Ien VGND 0.37144f
C8096 XA.XIR[14].XIC[12].icell.SM VGND 0.00502f
C8097 XA.XIR[14].XIC[13].icell.PUM VGND 0.00293f
C8098 XA.XIR[14].XIC[12].icell.Ien VGND 0.37144f
C8099 XA.XIR[14].XIC[11].icell.SM VGND 0.00502f
C8100 XA.XIR[14].XIC[12].icell.PUM VGND 0.00293f
C8101 XA.XIR[14].XIC[11].icell.Ien VGND 0.37144f
C8102 XA.XIR[14].XIC[10].icell.SM VGND 0.00502f
C8103 XA.XIR[14].XIC[11].icell.PUM VGND 0.00293f
C8104 XA.XIR[14].XIC[10].icell.Ien VGND 0.37144f
C8105 XA.XIR[14].XIC[9].icell.SM VGND 0.00502f
C8106 XA.XIR[14].XIC[10].icell.PUM VGND 0.00293f
C8107 XA.XIR[14].XIC[9].icell.Ien VGND 0.37144f
C8108 XA.XIR[14].XIC[8].icell.SM VGND 0.00502f
C8109 XA.XIR[14].XIC[9].icell.PUM VGND 0.00293f
C8110 XA.XIR[14].XIC[8].icell.Ien VGND 0.37144f
C8111 XA.XIR[14].XIC[7].icell.SM VGND 0.00502f
C8112 XA.XIR[14].XIC[8].icell.PUM VGND 0.00293f
C8113 XA.XIR[14].XIC[7].icell.Ien VGND 0.37144f
C8114 XA.XIR[14].XIC[6].icell.SM VGND 0.00502f
C8115 XA.XIR[14].XIC[7].icell.PUM VGND 0.00293f
C8116 XA.XIR[14].XIC[6].icell.Ien VGND 0.37144f
C8117 XA.XIR[14].XIC[5].icell.SM VGND 0.00502f
C8118 XA.XIR[14].XIC[6].icell.PUM VGND 0.00293f
C8119 XA.XIR[14].XIC[5].icell.Ien VGND 0.37144f
C8120 XA.XIR[14].XIC[4].icell.SM VGND 0.00502f
C8121 XA.XIR[14].XIC[5].icell.PUM VGND 0.00293f
C8122 XA.XIR[14].XIC[4].icell.Ien VGND 0.37144f
C8123 XA.XIR[14].XIC[3].icell.SM VGND 0.00502f
C8124 XA.XIR[14].XIC[4].icell.PUM VGND 0.00293f
C8125 XA.XIR[14].XIC[3].icell.Ien VGND 0.37144f
C8126 XA.XIR[14].XIC[2].icell.SM VGND 0.00502f
C8127 XA.XIR[14].XIC[3].icell.PUM VGND 0.00293f
C8128 XA.XIR[14].XIC[2].icell.Ien VGND 0.37144f
C8129 XA.XIR[14].XIC[1].icell.SM VGND 0.00502f
C8130 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80696f
C8131 XThR.Tn[14] VGND 14.14128f
C8132 XA.XIR[14].XIC[2].icell.PUM VGND 0.00293f
C8133 XA.XIR[14].XIC[1].icell.Ien VGND 0.37144f
C8134 XA.XIR[14].XIC[0].icell.SM VGND 0.00502f
C8135 a_n997_1579# VGND 0.54776f
C8136 XA.XIR[14].XIC[1].icell.PUM VGND 0.00293f
C8137 XA.XIR[14].XIC[0].icell.Ien VGND 0.37178f
C8138 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01044f
C8139 XA.XIR[14].XIC[0].icell.PUM VGND 0.00516f
C8140 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57579f
C8141 XA.XIR[14].XIC_dummy_left.icell.PUM VGND 0.00215f
C8142 a_n997_1803# VGND 0.53619f
C8143 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C8144 XA.XIR[14].XIC_15.icell.PDM VGND 0.18855f
C8145 XA.XIR[14].XIC[14].icell.PDM VGND 0.18809f
C8146 XA.XIR[14].XIC[13].icell.PDM VGND 0.18809f
C8147 XA.XIR[14].XIC[12].icell.PDM VGND 0.18809f
C8148 XA.XIR[14].XIC[11].icell.PDM VGND 0.18809f
C8149 XA.XIR[14].XIC[10].icell.PDM VGND 0.18809f
C8150 XA.XIR[14].XIC[9].icell.PDM VGND 0.18809f
C8151 XA.XIR[14].XIC[8].icell.PDM VGND 0.18809f
C8152 XA.XIR[14].XIC[7].icell.PDM VGND 0.18809f
C8153 XA.XIR[14].XIC[6].icell.PDM VGND 0.18809f
C8154 XA.XIR[14].XIC[5].icell.PDM VGND 0.18809f
C8155 XA.XIR[14].XIC[4].icell.PDM VGND 0.18809f
C8156 XA.XIR[14].XIC[3].icell.PDM VGND 0.18809f
C8157 XA.XIR[14].XIC[2].icell.PDM VGND 0.18809f
C8158 XA.XIR[14].XIC[1].icell.PDM VGND 0.18809f
C8159 XA.XIR[14].XIC[0].icell.PDM VGND 0.18817f
C8160 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C8161 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C8162 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C8163 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.608f
C8164 XA.XIR[13].XIC_15.icell.SM VGND 0.00474f
C8165 XA.XIR[13].XIC_dummy_right.icell.PUM VGND 0.00215f
C8166 XA.XIR[13].XIC_15.icell.Ien VGND 0.37063f
C8167 XA.XIR[13].XIC[14].icell.SM VGND 0.00502f
C8168 XA.XIR[13].XIC_15.icell.PUM VGND 0.00282f
C8169 XA.XIR[13].XIC[14].icell.Ien VGND 0.37144f
C8170 XA.XIR[13].XIC[13].icell.SM VGND 0.00502f
C8171 XA.XIR[13].XIC[14].icell.PUM VGND 0.00293f
C8172 XA.XIR[13].XIC[13].icell.Ien VGND 0.37144f
C8173 XA.XIR[13].XIC[12].icell.SM VGND 0.00502f
C8174 XA.XIR[13].XIC[13].icell.PUM VGND 0.00293f
C8175 XA.XIR[13].XIC[12].icell.Ien VGND 0.37144f
C8176 XA.XIR[13].XIC[11].icell.SM VGND 0.00502f
C8177 XA.XIR[13].XIC[12].icell.PUM VGND 0.00293f
C8178 XA.XIR[13].XIC[11].icell.Ien VGND 0.37144f
C8179 XA.XIR[13].XIC[10].icell.SM VGND 0.00502f
C8180 XA.XIR[13].XIC[11].icell.PUM VGND 0.00293f
C8181 XA.XIR[13].XIC[10].icell.Ien VGND 0.37144f
C8182 XA.XIR[13].XIC[9].icell.SM VGND 0.00502f
C8183 XA.XIR[13].XIC[10].icell.PUM VGND 0.00293f
C8184 XA.XIR[13].XIC[9].icell.Ien VGND 0.37144f
C8185 XA.XIR[13].XIC[8].icell.SM VGND 0.00502f
C8186 XA.XIR[13].XIC[9].icell.PUM VGND 0.00293f
C8187 XA.XIR[13].XIC[8].icell.Ien VGND 0.37144f
C8188 XA.XIR[13].XIC[7].icell.SM VGND 0.00502f
C8189 XA.XIR[13].XIC[8].icell.PUM VGND 0.00293f
C8190 XA.XIR[13].XIC[7].icell.Ien VGND 0.37144f
C8191 XA.XIR[13].XIC[6].icell.SM VGND 0.00502f
C8192 XA.XIR[13].XIC[7].icell.PUM VGND 0.00293f
C8193 XA.XIR[13].XIC[6].icell.Ien VGND 0.37144f
C8194 XA.XIR[13].XIC[5].icell.SM VGND 0.00502f
C8195 XA.XIR[13].XIC[6].icell.PUM VGND 0.00293f
C8196 XA.XIR[13].XIC[5].icell.Ien VGND 0.37144f
C8197 XA.XIR[13].XIC[4].icell.SM VGND 0.00502f
C8198 XA.XIR[13].XIC[5].icell.PUM VGND 0.00293f
C8199 XA.XIR[13].XIC[4].icell.Ien VGND 0.37144f
C8200 XA.XIR[13].XIC[3].icell.SM VGND 0.00502f
C8201 XA.XIR[13].XIC[4].icell.PUM VGND 0.00293f
C8202 XA.XIR[13].XIC[3].icell.Ien VGND 0.37144f
C8203 XA.XIR[13].XIC[2].icell.SM VGND 0.00502f
C8204 XA.XIR[13].XIC[3].icell.PUM VGND 0.00293f
C8205 XA.XIR[13].XIC[2].icell.Ien VGND 0.37144f
C8206 XA.XIR[13].XIC[1].icell.SM VGND 0.00502f
C8207 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.807f
C8208 XThR.Tn[13] VGND 14.01892f
C8209 XA.XIR[13].XIC[2].icell.PUM VGND 0.00293f
C8210 XA.XIR[13].XIC[1].icell.Ien VGND 0.37144f
C8211 XA.XIR[13].XIC[0].icell.SM VGND 0.00502f
C8212 XA.XIR[13].XIC[1].icell.PUM VGND 0.00293f
C8213 XA.XIR[13].XIC[0].icell.Ien VGND 0.37178f
C8214 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01044f
C8215 XA.XIR[13].XIC[0].icell.PUM VGND 0.00516f
C8216 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57425f
C8217 XA.XIR[13].XIC_dummy_left.icell.PUM VGND 0.00215f
C8218 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C8219 XA.XIR[13].XIC_15.icell.PDM VGND 0.18855f
C8220 XA.XIR[13].XIC[14].icell.PDM VGND 0.18809f
C8221 XA.XIR[13].XIC[13].icell.PDM VGND 0.18809f
C8222 XA.XIR[13].XIC[12].icell.PDM VGND 0.18809f
C8223 XA.XIR[13].XIC[11].icell.PDM VGND 0.18809f
C8224 XA.XIR[13].XIC[10].icell.PDM VGND 0.18809f
C8225 XA.XIR[13].XIC[9].icell.PDM VGND 0.18809f
C8226 XA.XIR[13].XIC[8].icell.PDM VGND 0.18809f
C8227 XA.XIR[13].XIC[7].icell.PDM VGND 0.18809f
C8228 XA.XIR[13].XIC[6].icell.PDM VGND 0.18809f
C8229 XA.XIR[13].XIC[5].icell.PDM VGND 0.18809f
C8230 XA.XIR[13].XIC[4].icell.PDM VGND 0.18809f
C8231 XA.XIR[13].XIC[3].icell.PDM VGND 0.18809f
C8232 XA.XIR[13].XIC[2].icell.PDM VGND 0.18809f
C8233 XA.XIR[13].XIC[1].icell.PDM VGND 0.18809f
C8234 XA.XIR[13].XIC[0].icell.PDM VGND 0.18817f
C8235 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C8236 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C8237 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C8238 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.608f
C8239 XA.XIR[12].XIC_15.icell.SM VGND 0.00474f
C8240 XA.XIR[12].XIC_dummy_right.icell.PUM VGND 0.00215f
C8241 XA.XIR[12].XIC_15.icell.Ien VGND 0.37063f
C8242 XA.XIR[12].XIC[14].icell.SM VGND 0.00502f
C8243 XA.XIR[12].XIC_15.icell.PUM VGND 0.00282f
C8244 XA.XIR[12].XIC[14].icell.Ien VGND 0.37144f
C8245 XA.XIR[12].XIC[13].icell.SM VGND 0.00502f
C8246 XA.XIR[12].XIC[14].icell.PUM VGND 0.00293f
C8247 XA.XIR[12].XIC[13].icell.Ien VGND 0.37144f
C8248 XA.XIR[12].XIC[12].icell.SM VGND 0.00502f
C8249 XA.XIR[12].XIC[13].icell.PUM VGND 0.00293f
C8250 XA.XIR[12].XIC[12].icell.Ien VGND 0.37144f
C8251 XA.XIR[12].XIC[11].icell.SM VGND 0.00502f
C8252 XA.XIR[12].XIC[12].icell.PUM VGND 0.00293f
C8253 XA.XIR[12].XIC[11].icell.Ien VGND 0.37144f
C8254 XA.XIR[12].XIC[10].icell.SM VGND 0.00502f
C8255 XA.XIR[12].XIC[11].icell.PUM VGND 0.00293f
C8256 XA.XIR[12].XIC[10].icell.Ien VGND 0.37144f
C8257 XA.XIR[12].XIC[9].icell.SM VGND 0.00502f
C8258 XA.XIR[12].XIC[10].icell.PUM VGND 0.00293f
C8259 XA.XIR[12].XIC[9].icell.Ien VGND 0.37144f
C8260 XA.XIR[12].XIC[8].icell.SM VGND 0.00502f
C8261 XA.XIR[12].XIC[9].icell.PUM VGND 0.00293f
C8262 XA.XIR[12].XIC[8].icell.Ien VGND 0.37144f
C8263 XA.XIR[12].XIC[7].icell.SM VGND 0.00502f
C8264 XA.XIR[12].XIC[8].icell.PUM VGND 0.00293f
C8265 XA.XIR[12].XIC[7].icell.Ien VGND 0.37144f
C8266 XA.XIR[12].XIC[6].icell.SM VGND 0.00502f
C8267 XA.XIR[12].XIC[7].icell.PUM VGND 0.00293f
C8268 XA.XIR[12].XIC[6].icell.Ien VGND 0.37144f
C8269 XA.XIR[12].XIC[5].icell.SM VGND 0.00502f
C8270 XA.XIR[12].XIC[6].icell.PUM VGND 0.00293f
C8271 XA.XIR[12].XIC[5].icell.Ien VGND 0.37144f
C8272 XA.XIR[12].XIC[4].icell.SM VGND 0.00502f
C8273 XA.XIR[12].XIC[5].icell.PUM VGND 0.00293f
C8274 XA.XIR[12].XIC[4].icell.Ien VGND 0.37144f
C8275 XA.XIR[12].XIC[3].icell.SM VGND 0.00502f
C8276 XA.XIR[12].XIC[4].icell.PUM VGND 0.00293f
C8277 XA.XIR[12].XIC[3].icell.Ien VGND 0.37144f
C8278 XA.XIR[12].XIC[2].icell.SM VGND 0.00502f
C8279 XA.XIR[12].XIC[3].icell.PUM VGND 0.00293f
C8280 XA.XIR[12].XIC[2].icell.Ien VGND 0.37144f
C8281 XA.XIR[12].XIC[1].icell.SM VGND 0.00502f
C8282 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80565f
C8283 XThR.Tn[12] VGND 13.90987f
C8284 XA.XIR[12].XIC[2].icell.PUM VGND 0.00293f
C8285 XA.XIR[12].XIC[1].icell.Ien VGND 0.37144f
C8286 XA.XIR[12].XIC[0].icell.SM VGND 0.00502f
C8287 XA.XIR[12].XIC[1].icell.PUM VGND 0.00293f
C8288 XA.XIR[12].XIC[0].icell.Ien VGND 0.37178f
C8289 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01044f
C8290 XA.XIR[12].XIC[0].icell.PUM VGND 0.00516f
C8291 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.57283f
C8292 XA.XIR[12].XIC_dummy_left.icell.PUM VGND 0.00215f
C8293 a_n997_2667# VGND 0.5457f
C8294 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C8295 XA.XIR[12].XIC_15.icell.PDM VGND 0.18855f
C8296 XA.XIR[12].XIC[14].icell.PDM VGND 0.18809f
C8297 XA.XIR[12].XIC[13].icell.PDM VGND 0.18809f
C8298 XA.XIR[12].XIC[12].icell.PDM VGND 0.18809f
C8299 XA.XIR[12].XIC[11].icell.PDM VGND 0.18809f
C8300 XA.XIR[12].XIC[10].icell.PDM VGND 0.18809f
C8301 XA.XIR[12].XIC[9].icell.PDM VGND 0.18809f
C8302 XA.XIR[12].XIC[8].icell.PDM VGND 0.18809f
C8303 XA.XIR[12].XIC[7].icell.PDM VGND 0.18809f
C8304 XA.XIR[12].XIC[6].icell.PDM VGND 0.18809f
C8305 XA.XIR[12].XIC[5].icell.PDM VGND 0.18809f
C8306 XA.XIR[12].XIC[4].icell.PDM VGND 0.18809f
C8307 XA.XIR[12].XIC[3].icell.PDM VGND 0.18809f
C8308 XA.XIR[12].XIC[2].icell.PDM VGND 0.18809f
C8309 XA.XIR[12].XIC[1].icell.PDM VGND 0.18809f
C8310 XA.XIR[12].XIC[0].icell.PDM VGND 0.18817f
C8311 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C8312 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C8313 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C8314 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.608f
C8315 XA.XIR[11].XIC_15.icell.SM VGND 0.00474f
C8316 XA.XIR[11].XIC_dummy_right.icell.PUM VGND 0.00215f
C8317 XA.XIR[11].XIC_15.icell.Ien VGND 0.37063f
C8318 XA.XIR[11].XIC[14].icell.SM VGND 0.00502f
C8319 XA.XIR[11].XIC_15.icell.PUM VGND 0.00282f
C8320 XA.XIR[11].XIC[14].icell.Ien VGND 0.37144f
C8321 XA.XIR[11].XIC[13].icell.SM VGND 0.00502f
C8322 XA.XIR[11].XIC[14].icell.PUM VGND 0.00293f
C8323 XA.XIR[11].XIC[13].icell.Ien VGND 0.37144f
C8324 XA.XIR[11].XIC[12].icell.SM VGND 0.00502f
C8325 XA.XIR[11].XIC[13].icell.PUM VGND 0.00293f
C8326 XA.XIR[11].XIC[12].icell.Ien VGND 0.37144f
C8327 XA.XIR[11].XIC[11].icell.SM VGND 0.00502f
C8328 XA.XIR[11].XIC[12].icell.PUM VGND 0.00293f
C8329 XA.XIR[11].XIC[11].icell.Ien VGND 0.37144f
C8330 XA.XIR[11].XIC[10].icell.SM VGND 0.00502f
C8331 XA.XIR[11].XIC[11].icell.PUM VGND 0.00293f
C8332 XA.XIR[11].XIC[10].icell.Ien VGND 0.37144f
C8333 XA.XIR[11].XIC[9].icell.SM VGND 0.00502f
C8334 XA.XIR[11].XIC[10].icell.PUM VGND 0.00293f
C8335 XA.XIR[11].XIC[9].icell.Ien VGND 0.37144f
C8336 XA.XIR[11].XIC[8].icell.SM VGND 0.00502f
C8337 XA.XIR[11].XIC[9].icell.PUM VGND 0.00293f
C8338 XA.XIR[11].XIC[8].icell.Ien VGND 0.37144f
C8339 XA.XIR[11].XIC[7].icell.SM VGND 0.00502f
C8340 XA.XIR[11].XIC[8].icell.PUM VGND 0.00293f
C8341 XA.XIR[11].XIC[7].icell.Ien VGND 0.37144f
C8342 XA.XIR[11].XIC[6].icell.SM VGND 0.00502f
C8343 XA.XIR[11].XIC[7].icell.PUM VGND 0.00293f
C8344 XA.XIR[11].XIC[6].icell.Ien VGND 0.37144f
C8345 XA.XIR[11].XIC[5].icell.SM VGND 0.00502f
C8346 XA.XIR[11].XIC[6].icell.PUM VGND 0.00293f
C8347 XA.XIR[11].XIC[5].icell.Ien VGND 0.37144f
C8348 XA.XIR[11].XIC[4].icell.SM VGND 0.00502f
C8349 XA.XIR[11].XIC[5].icell.PUM VGND 0.00293f
C8350 XA.XIR[11].XIC[4].icell.Ien VGND 0.37144f
C8351 XA.XIR[11].XIC[3].icell.SM VGND 0.00502f
C8352 XA.XIR[11].XIC[4].icell.PUM VGND 0.00293f
C8353 XA.XIR[11].XIC[3].icell.Ien VGND 0.37144f
C8354 XA.XIR[11].XIC[2].icell.SM VGND 0.00502f
C8355 XA.XIR[11].XIC[3].icell.PUM VGND 0.00293f
C8356 XA.XIR[11].XIC[2].icell.Ien VGND 0.37144f
C8357 XA.XIR[11].XIC[1].icell.SM VGND 0.00502f
C8358 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.808f
C8359 XThR.Tn[11] VGND 13.97038f
C8360 XA.XIR[11].XIC[2].icell.PUM VGND 0.00293f
C8361 XA.XIR[11].XIC[1].icell.Ien VGND 0.37144f
C8362 XA.XIR[11].XIC[0].icell.SM VGND 0.00502f
C8363 a_n997_2891# VGND 0.54795f
C8364 a_n1331_2891# VGND 0.00194f
C8365 XA.XIR[11].XIC[1].icell.PUM VGND 0.00293f
C8366 XA.XIR[11].XIC[0].icell.Ien VGND 0.37178f
C8367 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01044f
C8368 XA.XIR[11].XIC[0].icell.PUM VGND 0.00516f
C8369 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57297f
C8370 XA.XIR[11].XIC_dummy_left.icell.PUM VGND 0.00215f
C8371 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C8372 XA.XIR[11].XIC_15.icell.PDM VGND 0.18855f
C8373 XA.XIR[11].XIC[14].icell.PDM VGND 0.18809f
C8374 XA.XIR[11].XIC[13].icell.PDM VGND 0.18809f
C8375 XA.XIR[11].XIC[12].icell.PDM VGND 0.18809f
C8376 XA.XIR[11].XIC[11].icell.PDM VGND 0.18809f
C8377 XA.XIR[11].XIC[10].icell.PDM VGND 0.18809f
C8378 XA.XIR[11].XIC[9].icell.PDM VGND 0.18809f
C8379 XA.XIR[11].XIC[8].icell.PDM VGND 0.18809f
C8380 XA.XIR[11].XIC[7].icell.PDM VGND 0.18809f
C8381 XA.XIR[11].XIC[6].icell.PDM VGND 0.18809f
C8382 XA.XIR[11].XIC[5].icell.PDM VGND 0.18809f
C8383 XA.XIR[11].XIC[4].icell.PDM VGND 0.18809f
C8384 XA.XIR[11].XIC[3].icell.PDM VGND 0.18809f
C8385 XA.XIR[11].XIC[2].icell.PDM VGND 0.18809f
C8386 XA.XIR[11].XIC[1].icell.PDM VGND 0.18809f
C8387 XA.XIR[11].XIC[0].icell.PDM VGND 0.18817f
C8388 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C8389 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C8390 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C8391 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.608f
C8392 XA.XIR[10].XIC_15.icell.SM VGND 0.00474f
C8393 XA.XIR[10].XIC_dummy_right.icell.PUM VGND 0.00215f
C8394 XA.XIR[10].XIC_15.icell.Ien VGND 0.37063f
C8395 XA.XIR[10].XIC[14].icell.SM VGND 0.00502f
C8396 XA.XIR[10].XIC_15.icell.PUM VGND 0.00282f
C8397 XA.XIR[10].XIC[14].icell.Ien VGND 0.37144f
C8398 XA.XIR[10].XIC[13].icell.SM VGND 0.00502f
C8399 XA.XIR[10].XIC[14].icell.PUM VGND 0.00293f
C8400 XA.XIR[10].XIC[13].icell.Ien VGND 0.37144f
C8401 XA.XIR[10].XIC[12].icell.SM VGND 0.00502f
C8402 XA.XIR[10].XIC[13].icell.PUM VGND 0.00293f
C8403 XA.XIR[10].XIC[12].icell.Ien VGND 0.37144f
C8404 XA.XIR[10].XIC[11].icell.SM VGND 0.00502f
C8405 XA.XIR[10].XIC[12].icell.PUM VGND 0.00293f
C8406 XA.XIR[10].XIC[11].icell.Ien VGND 0.37144f
C8407 XA.XIR[10].XIC[10].icell.SM VGND 0.00502f
C8408 XA.XIR[10].XIC[11].icell.PUM VGND 0.00293f
C8409 XA.XIR[10].XIC[10].icell.Ien VGND 0.37144f
C8410 XA.XIR[10].XIC[9].icell.SM VGND 0.00502f
C8411 XA.XIR[10].XIC[10].icell.PUM VGND 0.00293f
C8412 XA.XIR[10].XIC[9].icell.Ien VGND 0.37144f
C8413 XA.XIR[10].XIC[8].icell.SM VGND 0.00502f
C8414 XA.XIR[10].XIC[9].icell.PUM VGND 0.00293f
C8415 XA.XIR[10].XIC[8].icell.Ien VGND 0.37144f
C8416 XA.XIR[10].XIC[7].icell.SM VGND 0.00502f
C8417 XA.XIR[10].XIC[8].icell.PUM VGND 0.00293f
C8418 XA.XIR[10].XIC[7].icell.Ien VGND 0.37144f
C8419 XA.XIR[10].XIC[6].icell.SM VGND 0.00502f
C8420 XA.XIR[10].XIC[7].icell.PUM VGND 0.00293f
C8421 XA.XIR[10].XIC[6].icell.Ien VGND 0.37144f
C8422 XA.XIR[10].XIC[5].icell.SM VGND 0.00502f
C8423 XA.XIR[10].XIC[6].icell.PUM VGND 0.00293f
C8424 XA.XIR[10].XIC[5].icell.Ien VGND 0.37144f
C8425 XA.XIR[10].XIC[4].icell.SM VGND 0.00502f
C8426 XA.XIR[10].XIC[5].icell.PUM VGND 0.00293f
C8427 XA.XIR[10].XIC[4].icell.Ien VGND 0.37144f
C8428 XA.XIR[10].XIC[3].icell.SM VGND 0.00502f
C8429 XA.XIR[10].XIC[4].icell.PUM VGND 0.00293f
C8430 XA.XIR[10].XIC[3].icell.Ien VGND 0.37144f
C8431 XA.XIR[10].XIC[2].icell.SM VGND 0.00502f
C8432 XA.XIR[10].XIC[3].icell.PUM VGND 0.00293f
C8433 XA.XIR[10].XIC[2].icell.Ien VGND 0.37144f
C8434 XA.XIR[10].XIC[1].icell.SM VGND 0.00502f
C8435 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80684f
C8436 XThR.Tn[10] VGND 13.91105f
C8437 XA.XIR[10].XIC[2].icell.PUM VGND 0.00293f
C8438 XA.XIR[10].XIC[1].icell.Ien VGND 0.37144f
C8439 XA.XIR[10].XIC[0].icell.SM VGND 0.00502f
C8440 XA.XIR[10].XIC[1].icell.PUM VGND 0.00293f
C8441 XA.XIR[10].XIC[0].icell.Ien VGND 0.37178f
C8442 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01044f
C8443 XA.XIR[10].XIC[0].icell.PUM VGND 0.00516f
C8444 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57425f
C8445 XA.XIR[10].XIC_dummy_left.icell.PUM VGND 0.00215f
C8446 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C8447 XA.XIR[10].XIC_15.icell.PDM VGND 0.18855f
C8448 XA.XIR[10].XIC[14].icell.PDM VGND 0.18809f
C8449 XA.XIR[10].XIC[13].icell.PDM VGND 0.18809f
C8450 XA.XIR[10].XIC[12].icell.PDM VGND 0.18809f
C8451 XA.XIR[10].XIC[11].icell.PDM VGND 0.18809f
C8452 XA.XIR[10].XIC[10].icell.PDM VGND 0.18809f
C8453 XA.XIR[10].XIC[9].icell.PDM VGND 0.18809f
C8454 XA.XIR[10].XIC[8].icell.PDM VGND 0.18809f
C8455 XA.XIR[10].XIC[7].icell.PDM VGND 0.18809f
C8456 XA.XIR[10].XIC[6].icell.PDM VGND 0.18809f
C8457 XA.XIR[10].XIC[5].icell.PDM VGND 0.18809f
C8458 XA.XIR[10].XIC[4].icell.PDM VGND 0.18809f
C8459 XA.XIR[10].XIC[3].icell.PDM VGND 0.18809f
C8460 XA.XIR[10].XIC[2].icell.PDM VGND 0.18809f
C8461 XA.XIR[10].XIC[1].icell.PDM VGND 0.18809f
C8462 XA.XIR[10].XIC[0].icell.PDM VGND 0.18817f
C8463 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C8464 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C8465 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C8466 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.608f
C8467 XA.XIR[9].XIC_15.icell.SM VGND 0.00474f
C8468 XA.XIR[9].XIC_dummy_right.icell.PUM VGND 0.00215f
C8469 XA.XIR[9].XIC_15.icell.Ien VGND 0.37063f
C8470 XA.XIR[9].XIC[14].icell.SM VGND 0.00502f
C8471 XA.XIR[9].XIC_15.icell.PUM VGND 0.00282f
C8472 XA.XIR[9].XIC[14].icell.Ien VGND 0.37144f
C8473 XA.XIR[9].XIC[13].icell.SM VGND 0.00502f
C8474 XA.XIR[9].XIC[14].icell.PUM VGND 0.00293f
C8475 XA.XIR[9].XIC[13].icell.Ien VGND 0.37144f
C8476 XA.XIR[9].XIC[12].icell.SM VGND 0.00502f
C8477 XA.XIR[9].XIC[13].icell.PUM VGND 0.00293f
C8478 XA.XIR[9].XIC[12].icell.Ien VGND 0.37144f
C8479 XA.XIR[9].XIC[11].icell.SM VGND 0.00502f
C8480 XA.XIR[9].XIC[12].icell.PUM VGND 0.00293f
C8481 XA.XIR[9].XIC[11].icell.Ien VGND 0.37144f
C8482 XA.XIR[9].XIC[10].icell.SM VGND 0.00502f
C8483 XA.XIR[9].XIC[11].icell.PUM VGND 0.00293f
C8484 XA.XIR[9].XIC[10].icell.Ien VGND 0.37144f
C8485 XA.XIR[9].XIC[9].icell.SM VGND 0.00502f
C8486 XA.XIR[9].XIC[10].icell.PUM VGND 0.00293f
C8487 XA.XIR[9].XIC[9].icell.Ien VGND 0.37144f
C8488 XA.XIR[9].XIC[8].icell.SM VGND 0.00502f
C8489 XA.XIR[9].XIC[9].icell.PUM VGND 0.00293f
C8490 XA.XIR[9].XIC[8].icell.Ien VGND 0.37144f
C8491 XA.XIR[9].XIC[7].icell.SM VGND 0.00502f
C8492 XA.XIR[9].XIC[8].icell.PUM VGND 0.00293f
C8493 XA.XIR[9].XIC[7].icell.Ien VGND 0.37144f
C8494 XA.XIR[9].XIC[6].icell.SM VGND 0.00502f
C8495 XA.XIR[9].XIC[7].icell.PUM VGND 0.00293f
C8496 XA.XIR[9].XIC[6].icell.Ien VGND 0.37144f
C8497 XA.XIR[9].XIC[5].icell.SM VGND 0.00502f
C8498 XA.XIR[9].XIC[6].icell.PUM VGND 0.00293f
C8499 XA.XIR[9].XIC[5].icell.Ien VGND 0.37144f
C8500 XA.XIR[9].XIC[4].icell.SM VGND 0.00502f
C8501 XA.XIR[9].XIC[5].icell.PUM VGND 0.00293f
C8502 XA.XIR[9].XIC[4].icell.Ien VGND 0.37144f
C8503 XA.XIR[9].XIC[3].icell.SM VGND 0.00502f
C8504 XA.XIR[9].XIC[4].icell.PUM VGND 0.00293f
C8505 XA.XIR[9].XIC[3].icell.Ien VGND 0.37144f
C8506 XA.XIR[9].XIC[2].icell.SM VGND 0.00502f
C8507 XA.XIR[9].XIC[3].icell.PUM VGND 0.00293f
C8508 XA.XIR[9].XIC[2].icell.Ien VGND 0.37144f
C8509 XA.XIR[9].XIC[1].icell.SM VGND 0.00502f
C8510 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.8087f
C8511 XA.XIR[9].XIC[2].icell.PUM VGND 0.00293f
C8512 XA.XIR[9].XIC[1].icell.Ien VGND 0.37144f
C8513 XA.XIR[9].XIC[0].icell.SM VGND 0.00502f
C8514 XThR.Tn[9] VGND 13.95272f
C8515 a_n997_3755# VGND 0.54861f
C8516 XA.XIR[9].XIC[1].icell.PUM VGND 0.00293f
C8517 XA.XIR[9].XIC[0].icell.Ien VGND 0.37178f
C8518 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01044f
C8519 XA.XIR[9].XIC[0].icell.PUM VGND 0.00516f
C8520 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.57323f
C8521 a_n997_3979# VGND 0.54721f
C8522 XA.XIR[9].XIC_dummy_left.icell.PUM VGND 0.00215f
C8523 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C8524 XA.XIR[9].XIC_15.icell.PDM VGND 0.18855f
C8525 XA.XIR[9].XIC[14].icell.PDM VGND 0.18809f
C8526 XA.XIR[9].XIC[13].icell.PDM VGND 0.18809f
C8527 XA.XIR[9].XIC[12].icell.PDM VGND 0.18809f
C8528 XA.XIR[9].XIC[11].icell.PDM VGND 0.18809f
C8529 XA.XIR[9].XIC[10].icell.PDM VGND 0.18809f
C8530 XA.XIR[9].XIC[9].icell.PDM VGND 0.18809f
C8531 XA.XIR[9].XIC[8].icell.PDM VGND 0.18809f
C8532 XA.XIR[9].XIC[7].icell.PDM VGND 0.18809f
C8533 XA.XIR[9].XIC[6].icell.PDM VGND 0.18809f
C8534 XA.XIR[9].XIC[5].icell.PDM VGND 0.18809f
C8535 XA.XIR[9].XIC[4].icell.PDM VGND 0.18809f
C8536 XA.XIR[9].XIC[3].icell.PDM VGND 0.18809f
C8537 XA.XIR[9].XIC[2].icell.PDM VGND 0.18809f
C8538 XA.XIR[9].XIC[1].icell.PDM VGND 0.18809f
C8539 XA.XIR[9].XIC[0].icell.PDM VGND 0.18817f
C8540 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C8541 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C8542 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C8543 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.608f
C8544 XA.XIR[8].XIC_15.icell.SM VGND 0.00474f
C8545 XA.XIR[8].XIC_dummy_right.icell.PUM VGND 0.00215f
C8546 XA.XIR[8].XIC_15.icell.Ien VGND 0.37063f
C8547 XA.XIR[8].XIC[14].icell.SM VGND 0.00502f
C8548 XA.XIR[8].XIC_15.icell.PUM VGND 0.00282f
C8549 XA.XIR[8].XIC[14].icell.Ien VGND 0.37144f
C8550 XA.XIR[8].XIC[13].icell.SM VGND 0.00502f
C8551 XA.XIR[8].XIC[14].icell.PUM VGND 0.00293f
C8552 XA.XIR[8].XIC[13].icell.Ien VGND 0.37144f
C8553 XA.XIR[8].XIC[12].icell.SM VGND 0.00502f
C8554 XA.XIR[8].XIC[13].icell.PUM VGND 0.00293f
C8555 XA.XIR[8].XIC[12].icell.Ien VGND 0.37144f
C8556 XA.XIR[8].XIC[11].icell.SM VGND 0.00502f
C8557 XA.XIR[8].XIC[12].icell.PUM VGND 0.00293f
C8558 XA.XIR[8].XIC[11].icell.Ien VGND 0.37144f
C8559 XA.XIR[8].XIC[10].icell.SM VGND 0.00502f
C8560 XA.XIR[8].XIC[11].icell.PUM VGND 0.00293f
C8561 XA.XIR[8].XIC[10].icell.Ien VGND 0.37144f
C8562 XA.XIR[8].XIC[9].icell.SM VGND 0.00502f
C8563 XA.XIR[8].XIC[10].icell.PUM VGND 0.00293f
C8564 XA.XIR[8].XIC[9].icell.Ien VGND 0.37144f
C8565 XA.XIR[8].XIC[8].icell.SM VGND 0.00502f
C8566 XA.XIR[8].XIC[9].icell.PUM VGND 0.00293f
C8567 XA.XIR[8].XIC[8].icell.Ien VGND 0.37144f
C8568 XA.XIR[8].XIC[7].icell.SM VGND 0.00502f
C8569 XA.XIR[8].XIC[8].icell.PUM VGND 0.00293f
C8570 XA.XIR[8].XIC[7].icell.Ien VGND 0.37144f
C8571 XA.XIR[8].XIC[6].icell.SM VGND 0.00502f
C8572 XA.XIR[8].XIC[7].icell.PUM VGND 0.00293f
C8573 XA.XIR[8].XIC[6].icell.Ien VGND 0.37144f
C8574 XA.XIR[8].XIC[5].icell.SM VGND 0.00502f
C8575 XA.XIR[8].XIC[6].icell.PUM VGND 0.00293f
C8576 XA.XIR[8].XIC[5].icell.Ien VGND 0.37144f
C8577 XA.XIR[8].XIC[4].icell.SM VGND 0.00502f
C8578 XA.XIR[8].XIC[5].icell.PUM VGND 0.00293f
C8579 XA.XIR[8].XIC[4].icell.Ien VGND 0.37144f
C8580 XA.XIR[8].XIC[3].icell.SM VGND 0.00502f
C8581 XA.XIR[8].XIC[4].icell.PUM VGND 0.00293f
C8582 XA.XIR[8].XIC[3].icell.Ien VGND 0.37144f
C8583 XA.XIR[8].XIC[2].icell.SM VGND 0.00502f
C8584 XA.XIR[8].XIC[3].icell.PUM VGND 0.00293f
C8585 XA.XIR[8].XIC[2].icell.Ien VGND 0.37144f
C8586 XA.XIR[8].XIC[1].icell.SM VGND 0.00502f
C8587 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80602f
C8588 XA.XIR[8].XIC[2].icell.PUM VGND 0.00293f
C8589 XA.XIR[8].XIC[1].icell.Ien VGND 0.37144f
C8590 XA.XIR[8].XIC[0].icell.SM VGND 0.00502f
C8591 XThR.Tn[8] VGND 13.8971f
C8592 XA.XIR[8].XIC[1].icell.PUM VGND 0.00293f
C8593 XA.XIR[8].XIC[0].icell.Ien VGND 0.37178f
C8594 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01044f
C8595 XA.XIR[8].XIC[0].icell.PUM VGND 0.00516f
C8596 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57311f
C8597 XA.XIR[8].XIC_dummy_left.icell.PUM VGND 0.00215f
C8598 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C8599 XA.XIR[8].XIC_15.icell.PDM VGND 0.18855f
C8600 XA.XIR[8].XIC[14].icell.PDM VGND 0.18809f
C8601 XA.XIR[8].XIC[13].icell.PDM VGND 0.18809f
C8602 XA.XIR[8].XIC[12].icell.PDM VGND 0.18809f
C8603 XA.XIR[8].XIC[11].icell.PDM VGND 0.18809f
C8604 XA.XIR[8].XIC[10].icell.PDM VGND 0.18809f
C8605 XA.XIR[8].XIC[9].icell.PDM VGND 0.18809f
C8606 XA.XIR[8].XIC[8].icell.PDM VGND 0.18809f
C8607 XA.XIR[8].XIC[7].icell.PDM VGND 0.18809f
C8608 XA.XIR[8].XIC[6].icell.PDM VGND 0.18809f
C8609 XA.XIR[8].XIC[5].icell.PDM VGND 0.18809f
C8610 XA.XIR[8].XIC[4].icell.PDM VGND 0.18809f
C8611 XA.XIR[8].XIC[3].icell.PDM VGND 0.18809f
C8612 XA.XIR[8].XIC[2].icell.PDM VGND 0.18809f
C8613 XA.XIR[8].XIC[1].icell.PDM VGND 0.18809f
C8614 XA.XIR[8].XIC[0].icell.PDM VGND 0.18817f
C8615 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C8616 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C8617 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C8618 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.608f
C8619 XA.XIR[7].XIC_15.icell.SM VGND 0.00474f
C8620 XA.XIR[7].XIC_dummy_right.icell.PUM VGND 0.00215f
C8621 XA.XIR[7].XIC_15.icell.Ien VGND 0.37063f
C8622 XA.XIR[7].XIC[14].icell.SM VGND 0.00502f
C8623 XA.XIR[7].XIC_15.icell.PUM VGND 0.00282f
C8624 XA.XIR[7].XIC[14].icell.Ien VGND 0.37144f
C8625 XA.XIR[7].XIC[13].icell.SM VGND 0.00502f
C8626 XA.XIR[7].XIC[14].icell.PUM VGND 0.00293f
C8627 XA.XIR[7].XIC[13].icell.Ien VGND 0.37144f
C8628 XA.XIR[7].XIC[12].icell.SM VGND 0.00502f
C8629 XA.XIR[7].XIC[13].icell.PUM VGND 0.00293f
C8630 XA.XIR[7].XIC[12].icell.Ien VGND 0.37144f
C8631 XA.XIR[7].XIC[11].icell.SM VGND 0.00502f
C8632 XA.XIR[7].XIC[12].icell.PUM VGND 0.00293f
C8633 XA.XIR[7].XIC[11].icell.Ien VGND 0.37144f
C8634 XA.XIR[7].XIC[10].icell.SM VGND 0.00502f
C8635 XA.XIR[7].XIC[11].icell.PUM VGND 0.00293f
C8636 XA.XIR[7].XIC[10].icell.Ien VGND 0.37144f
C8637 XA.XIR[7].XIC[9].icell.SM VGND 0.00502f
C8638 XA.XIR[7].XIC[10].icell.PUM VGND 0.00293f
C8639 XA.XIR[7].XIC[9].icell.Ien VGND 0.37144f
C8640 XA.XIR[7].XIC[8].icell.SM VGND 0.00502f
C8641 XA.XIR[7].XIC[9].icell.PUM VGND 0.00293f
C8642 XA.XIR[7].XIC[8].icell.Ien VGND 0.37144f
C8643 XA.XIR[7].XIC[7].icell.SM VGND 0.00502f
C8644 XA.XIR[7].XIC[8].icell.PUM VGND 0.00293f
C8645 XA.XIR[7].XIC[7].icell.Ien VGND 0.37144f
C8646 XA.XIR[7].XIC[6].icell.SM VGND 0.00502f
C8647 XA.XIR[7].XIC[7].icell.PUM VGND 0.00293f
C8648 XA.XIR[7].XIC[6].icell.Ien VGND 0.37144f
C8649 XA.XIR[7].XIC[5].icell.SM VGND 0.00502f
C8650 XA.XIR[7].XIC[6].icell.PUM VGND 0.00293f
C8651 XA.XIR[7].XIC[5].icell.Ien VGND 0.37144f
C8652 XA.XIR[7].XIC[4].icell.SM VGND 0.00502f
C8653 XA.XIR[7].XIC[5].icell.PUM VGND 0.00293f
C8654 XA.XIR[7].XIC[4].icell.Ien VGND 0.37144f
C8655 XA.XIR[7].XIC[3].icell.SM VGND 0.00502f
C8656 XA.XIR[7].XIC[4].icell.PUM VGND 0.00293f
C8657 XA.XIR[7].XIC[3].icell.Ien VGND 0.37144f
C8658 XA.XIR[7].XIC[2].icell.SM VGND 0.00502f
C8659 XA.XIR[7].XIC[3].icell.PUM VGND 0.00293f
C8660 XA.XIR[7].XIC[2].icell.Ien VGND 0.37144f
C8661 XA.XIR[7].XIC[1].icell.SM VGND 0.00502f
C8662 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80634f
C8663 XA.XIR[7].XIC[2].icell.PUM VGND 0.00293f
C8664 XA.XIR[7].XIC[1].icell.Ien VGND 0.37144f
C8665 XA.XIR[7].XIC[0].icell.SM VGND 0.00502f
C8666 XA.XIR[7].XIC[1].icell.PUM VGND 0.00293f
C8667 XA.XIR[7].XIC[0].icell.Ien VGND 0.37178f
C8668 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01044f
C8669 XThR.Tn[7] VGND 14.38144f
C8670 XThR.XTBN.A VGND 1.22814f
C8671 XA.XIR[7].XIC[0].icell.PUM VGND 0.00516f
C8672 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57579f
C8673 XA.XIR[7].XIC_dummy_left.icell.PUM VGND 0.00222f
C8674 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C8675 XA.XIR[7].XIC_15.icell.PDM VGND 0.18855f
C8676 XA.XIR[7].XIC[14].icell.PDM VGND 0.18809f
C8677 XA.XIR[7].XIC[13].icell.PDM VGND 0.18809f
C8678 XA.XIR[7].XIC[12].icell.PDM VGND 0.18809f
C8679 XA.XIR[7].XIC[11].icell.PDM VGND 0.18809f
C8680 XA.XIR[7].XIC[10].icell.PDM VGND 0.18809f
C8681 XA.XIR[7].XIC[9].icell.PDM VGND 0.18809f
C8682 XA.XIR[7].XIC[8].icell.PDM VGND 0.18809f
C8683 XA.XIR[7].XIC[7].icell.PDM VGND 0.18809f
C8684 XA.XIR[7].XIC[6].icell.PDM VGND 0.18809f
C8685 XA.XIR[7].XIC[5].icell.PDM VGND 0.18809f
C8686 XA.XIR[7].XIC[4].icell.PDM VGND 0.18809f
C8687 XA.XIR[7].XIC[3].icell.PDM VGND 0.18809f
C8688 XA.XIR[7].XIC[2].icell.PDM VGND 0.18809f
C8689 XA.XIR[7].XIC[1].icell.PDM VGND 0.18809f
C8690 XA.XIR[7].XIC[0].icell.PDM VGND 0.18817f
C8691 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C8692 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C8693 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C8694 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.608f
C8695 XA.XIR[6].XIC_15.icell.SM VGND 0.00474f
C8696 XA.XIR[6].XIC_dummy_right.icell.PUM VGND 0.00215f
C8697 XA.XIR[6].XIC_15.icell.Ien VGND 0.37063f
C8698 XA.XIR[6].XIC[14].icell.SM VGND 0.00502f
C8699 XA.XIR[6].XIC_15.icell.PUM VGND 0.00282f
C8700 XA.XIR[6].XIC[14].icell.Ien VGND 0.37144f
C8701 XA.XIR[6].XIC[13].icell.SM VGND 0.00502f
C8702 XA.XIR[6].XIC[14].icell.PUM VGND 0.00293f
C8703 XA.XIR[6].XIC[13].icell.Ien VGND 0.37144f
C8704 XA.XIR[6].XIC[12].icell.SM VGND 0.00502f
C8705 XA.XIR[6].XIC[13].icell.PUM VGND 0.00293f
C8706 XA.XIR[6].XIC[12].icell.Ien VGND 0.37144f
C8707 XA.XIR[6].XIC[11].icell.SM VGND 0.00502f
C8708 XA.XIR[6].XIC[12].icell.PUM VGND 0.00293f
C8709 XA.XIR[6].XIC[11].icell.Ien VGND 0.37144f
C8710 XA.XIR[6].XIC[10].icell.SM VGND 0.00502f
C8711 XA.XIR[6].XIC[11].icell.PUM VGND 0.00293f
C8712 XA.XIR[6].XIC[10].icell.Ien VGND 0.37144f
C8713 XA.XIR[6].XIC[9].icell.SM VGND 0.00502f
C8714 XA.XIR[6].XIC[10].icell.PUM VGND 0.00293f
C8715 XA.XIR[6].XIC[9].icell.Ien VGND 0.37144f
C8716 XA.XIR[6].XIC[8].icell.SM VGND 0.00502f
C8717 XA.XIR[6].XIC[9].icell.PUM VGND 0.00293f
C8718 XA.XIR[6].XIC[8].icell.Ien VGND 0.37144f
C8719 XA.XIR[6].XIC[7].icell.SM VGND 0.00502f
C8720 XA.XIR[6].XIC[8].icell.PUM VGND 0.00293f
C8721 XA.XIR[6].XIC[7].icell.Ien VGND 0.37144f
C8722 XA.XIR[6].XIC[6].icell.SM VGND 0.00502f
C8723 XA.XIR[6].XIC[7].icell.PUM VGND 0.00293f
C8724 XA.XIR[6].XIC[6].icell.Ien VGND 0.37144f
C8725 XA.XIR[6].XIC[5].icell.SM VGND 0.00502f
C8726 XA.XIR[6].XIC[6].icell.PUM VGND 0.00293f
C8727 XA.XIR[6].XIC[5].icell.Ien VGND 0.37144f
C8728 XA.XIR[6].XIC[4].icell.SM VGND 0.00502f
C8729 XA.XIR[6].XIC[5].icell.PUM VGND 0.00293f
C8730 XA.XIR[6].XIC[4].icell.Ien VGND 0.37144f
C8731 XA.XIR[6].XIC[3].icell.SM VGND 0.00502f
C8732 XA.XIR[6].XIC[4].icell.PUM VGND 0.00293f
C8733 XA.XIR[6].XIC[3].icell.Ien VGND 0.37144f
C8734 XA.XIR[6].XIC[2].icell.SM VGND 0.00502f
C8735 XA.XIR[6].XIC[3].icell.PUM VGND 0.00293f
C8736 XA.XIR[6].XIC[2].icell.Ien VGND 0.37144f
C8737 XA.XIR[6].XIC[1].icell.SM VGND 0.00502f
C8738 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80729f
C8739 XA.XIR[6].XIC[2].icell.PUM VGND 0.00293f
C8740 XA.XIR[6].XIC[1].icell.Ien VGND 0.37144f
C8741 XA.XIR[6].XIC[0].icell.SM VGND 0.00502f
C8742 XA.XIR[6].XIC[1].icell.PUM VGND 0.00293f
C8743 XA.XIR[6].XIC[0].icell.Ien VGND 0.37178f
C8744 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01044f
C8745 XA.XIR[6].XIC[0].icell.PUM VGND 0.00516f
C8746 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57425f
C8747 XThR.Tn[6] VGND 13.98754f
C8748 a_n1049_5317# VGND 0.02283f
C8749 XA.XIR[6].XIC_dummy_left.icell.PUM VGND 0.00215f
C8750 XThR.XTB7.Y VGND 1.36132f
C8751 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C8752 XA.XIR[6].XIC_15.icell.PDM VGND 0.18855f
C8753 XA.XIR[6].XIC[14].icell.PDM VGND 0.18809f
C8754 XA.XIR[6].XIC[13].icell.PDM VGND 0.18809f
C8755 XA.XIR[6].XIC[12].icell.PDM VGND 0.18809f
C8756 XA.XIR[6].XIC[11].icell.PDM VGND 0.18809f
C8757 XA.XIR[6].XIC[10].icell.PDM VGND 0.18809f
C8758 XA.XIR[6].XIC[9].icell.PDM VGND 0.18809f
C8759 XA.XIR[6].XIC[8].icell.PDM VGND 0.18809f
C8760 XA.XIR[6].XIC[7].icell.PDM VGND 0.18809f
C8761 XA.XIR[6].XIC[6].icell.PDM VGND 0.18809f
C8762 XA.XIR[6].XIC[5].icell.PDM VGND 0.18809f
C8763 XA.XIR[6].XIC[4].icell.PDM VGND 0.18809f
C8764 XA.XIR[6].XIC[3].icell.PDM VGND 0.18809f
C8765 XA.XIR[6].XIC[2].icell.PDM VGND 0.18809f
C8766 XA.XIR[6].XIC[1].icell.PDM VGND 0.18809f
C8767 XA.XIR[6].XIC[0].icell.PDM VGND 0.18817f
C8768 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C8769 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C8770 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C8771 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.608f
C8772 XA.XIR[5].XIC_15.icell.SM VGND 0.00474f
C8773 XA.XIR[5].XIC_dummy_right.icell.PUM VGND 0.00215f
C8774 XA.XIR[5].XIC_15.icell.Ien VGND 0.37063f
C8775 XA.XIR[5].XIC[14].icell.SM VGND 0.00502f
C8776 XA.XIR[5].XIC_15.icell.PUM VGND 0.00282f
C8777 XA.XIR[5].XIC[14].icell.Ien VGND 0.37144f
C8778 XA.XIR[5].XIC[13].icell.SM VGND 0.00502f
C8779 XA.XIR[5].XIC[14].icell.PUM VGND 0.00293f
C8780 XA.XIR[5].XIC[13].icell.Ien VGND 0.37144f
C8781 XA.XIR[5].XIC[12].icell.SM VGND 0.00502f
C8782 XA.XIR[5].XIC[13].icell.PUM VGND 0.00293f
C8783 XA.XIR[5].XIC[12].icell.Ien VGND 0.37144f
C8784 XA.XIR[5].XIC[11].icell.SM VGND 0.00502f
C8785 XA.XIR[5].XIC[12].icell.PUM VGND 0.00293f
C8786 XA.XIR[5].XIC[11].icell.Ien VGND 0.37144f
C8787 XA.XIR[5].XIC[10].icell.SM VGND 0.00502f
C8788 XA.XIR[5].XIC[11].icell.PUM VGND 0.00293f
C8789 XA.XIR[5].XIC[10].icell.Ien VGND 0.37144f
C8790 XA.XIR[5].XIC[9].icell.SM VGND 0.00502f
C8791 XA.XIR[5].XIC[10].icell.PUM VGND 0.00293f
C8792 XA.XIR[5].XIC[9].icell.Ien VGND 0.37144f
C8793 XA.XIR[5].XIC[8].icell.SM VGND 0.00502f
C8794 XA.XIR[5].XIC[9].icell.PUM VGND 0.00293f
C8795 XA.XIR[5].XIC[8].icell.Ien VGND 0.37144f
C8796 XA.XIR[5].XIC[7].icell.SM VGND 0.00502f
C8797 XA.XIR[5].XIC[8].icell.PUM VGND 0.00293f
C8798 XA.XIR[5].XIC[7].icell.Ien VGND 0.37144f
C8799 XA.XIR[5].XIC[6].icell.SM VGND 0.00502f
C8800 XA.XIR[5].XIC[7].icell.PUM VGND 0.00293f
C8801 XA.XIR[5].XIC[6].icell.Ien VGND 0.37144f
C8802 XA.XIR[5].XIC[5].icell.SM VGND 0.00502f
C8803 XA.XIR[5].XIC[6].icell.PUM VGND 0.00293f
C8804 XA.XIR[5].XIC[5].icell.Ien VGND 0.37144f
C8805 XA.XIR[5].XIC[4].icell.SM VGND 0.00502f
C8806 XA.XIR[5].XIC[5].icell.PUM VGND 0.00293f
C8807 XA.XIR[5].XIC[4].icell.Ien VGND 0.37144f
C8808 XA.XIR[5].XIC[3].icell.SM VGND 0.00502f
C8809 XA.XIR[5].XIC[4].icell.PUM VGND 0.00293f
C8810 XA.XIR[5].XIC[3].icell.Ien VGND 0.37144f
C8811 XA.XIR[5].XIC[2].icell.SM VGND 0.00502f
C8812 XA.XIR[5].XIC[3].icell.PUM VGND 0.00293f
C8813 XA.XIR[5].XIC[2].icell.Ien VGND 0.37144f
C8814 XA.XIR[5].XIC[1].icell.SM VGND 0.00502f
C8815 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80598f
C8816 XA.XIR[5].XIC[2].icell.PUM VGND 0.00293f
C8817 XA.XIR[5].XIC[1].icell.Ien VGND 0.37144f
C8818 XA.XIR[5].XIC[0].icell.SM VGND 0.00502f
C8819 a_n1049_5611# VGND 0.02888f
C8820 XA.XIR[5].XIC[1].icell.PUM VGND 0.00293f
C8821 XA.XIR[5].XIC[0].icell.Ien VGND 0.37178f
C8822 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01044f
C8823 XA.XIR[5].XIC[0].icell.PUM VGND 0.00516f
C8824 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57291f
C8825 XA.XIR[5].XIC_dummy_left.icell.PUM VGND 0.00215f
C8826 XThR.Tn[5] VGND 13.96673f
C8827 XThR.XTB6.Y VGND 1.38212f
C8828 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C8829 XA.XIR[5].XIC_15.icell.PDM VGND 0.18855f
C8830 XA.XIR[5].XIC[14].icell.PDM VGND 0.18809f
C8831 XA.XIR[5].XIC[13].icell.PDM VGND 0.18809f
C8832 XA.XIR[5].XIC[12].icell.PDM VGND 0.18809f
C8833 XA.XIR[5].XIC[11].icell.PDM VGND 0.18809f
C8834 XA.XIR[5].XIC[10].icell.PDM VGND 0.18809f
C8835 XA.XIR[5].XIC[9].icell.PDM VGND 0.18809f
C8836 XA.XIR[5].XIC[8].icell.PDM VGND 0.18809f
C8837 XA.XIR[5].XIC[7].icell.PDM VGND 0.18809f
C8838 XA.XIR[5].XIC[6].icell.PDM VGND 0.18809f
C8839 XA.XIR[5].XIC[5].icell.PDM VGND 0.18809f
C8840 XA.XIR[5].XIC[4].icell.PDM VGND 0.18809f
C8841 XA.XIR[5].XIC[3].icell.PDM VGND 0.18809f
C8842 XA.XIR[5].XIC[2].icell.PDM VGND 0.18809f
C8843 XA.XIR[5].XIC[1].icell.PDM VGND 0.18809f
C8844 XA.XIR[5].XIC[0].icell.PDM VGND 0.18817f
C8845 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C8846 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C8847 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C8848 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.608f
C8849 XA.XIR[4].XIC_15.icell.SM VGND 0.00474f
C8850 XA.XIR[4].XIC_dummy_right.icell.PUM VGND 0.00215f
C8851 XA.XIR[4].XIC_15.icell.Ien VGND 0.37063f
C8852 XA.XIR[4].XIC[14].icell.SM VGND 0.00502f
C8853 XA.XIR[4].XIC_15.icell.PUM VGND 0.00282f
C8854 XA.XIR[4].XIC[14].icell.Ien VGND 0.37144f
C8855 XA.XIR[4].XIC[13].icell.SM VGND 0.00502f
C8856 XA.XIR[4].XIC[14].icell.PUM VGND 0.00293f
C8857 XA.XIR[4].XIC[13].icell.Ien VGND 0.37144f
C8858 XA.XIR[4].XIC[12].icell.SM VGND 0.00502f
C8859 XA.XIR[4].XIC[13].icell.PUM VGND 0.00293f
C8860 XA.XIR[4].XIC[12].icell.Ien VGND 0.37144f
C8861 XA.XIR[4].XIC[11].icell.SM VGND 0.00502f
C8862 XA.XIR[4].XIC[12].icell.PUM VGND 0.00293f
C8863 XA.XIR[4].XIC[11].icell.Ien VGND 0.37144f
C8864 XA.XIR[4].XIC[10].icell.SM VGND 0.00502f
C8865 XA.XIR[4].XIC[11].icell.PUM VGND 0.00293f
C8866 XA.XIR[4].XIC[10].icell.Ien VGND 0.37144f
C8867 XA.XIR[4].XIC[9].icell.SM VGND 0.00502f
C8868 XA.XIR[4].XIC[10].icell.PUM VGND 0.00293f
C8869 XA.XIR[4].XIC[9].icell.Ien VGND 0.37144f
C8870 XA.XIR[4].XIC[8].icell.SM VGND 0.00502f
C8871 XA.XIR[4].XIC[9].icell.PUM VGND 0.00293f
C8872 XA.XIR[4].XIC[8].icell.Ien VGND 0.37144f
C8873 XA.XIR[4].XIC[7].icell.SM VGND 0.00502f
C8874 XA.XIR[4].XIC[8].icell.PUM VGND 0.00293f
C8875 XA.XIR[4].XIC[7].icell.Ien VGND 0.37144f
C8876 XA.XIR[4].XIC[6].icell.SM VGND 0.00502f
C8877 XA.XIR[4].XIC[7].icell.PUM VGND 0.00293f
C8878 XA.XIR[4].XIC[6].icell.Ien VGND 0.37144f
C8879 XA.XIR[4].XIC[5].icell.SM VGND 0.00502f
C8880 XA.XIR[4].XIC[6].icell.PUM VGND 0.00293f
C8881 XA.XIR[4].XIC[5].icell.Ien VGND 0.37144f
C8882 XA.XIR[4].XIC[4].icell.SM VGND 0.00502f
C8883 XA.XIR[4].XIC[5].icell.PUM VGND 0.00293f
C8884 XA.XIR[4].XIC[4].icell.Ien VGND 0.37144f
C8885 XA.XIR[4].XIC[3].icell.SM VGND 0.00502f
C8886 XA.XIR[4].XIC[4].icell.PUM VGND 0.00293f
C8887 XA.XIR[4].XIC[3].icell.Ien VGND 0.37144f
C8888 XA.XIR[4].XIC[2].icell.SM VGND 0.00502f
C8889 XA.XIR[4].XIC[3].icell.PUM VGND 0.00293f
C8890 XA.XIR[4].XIC[2].icell.Ien VGND 0.37144f
C8891 XA.XIR[4].XIC[1].icell.SM VGND 0.00502f
C8892 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.8077f
C8893 XA.XIR[4].XIC[2].icell.PUM VGND 0.00293f
C8894 XA.XIR[4].XIC[1].icell.Ien VGND 0.37144f
C8895 XA.XIR[4].XIC[0].icell.SM VGND 0.00502f
C8896 XA.XIR[4].XIC[1].icell.PUM VGND 0.00293f
C8897 XA.XIR[4].XIC[0].icell.Ien VGND 0.37178f
C8898 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01044f
C8899 XA.XIR[4].XIC[0].icell.PUM VGND 0.00516f
C8900 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57336f
C8901 XA.XIR[4].XIC_dummy_left.icell.PUM VGND 0.00215f
C8902 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C8903 XA.XIR[4].XIC_15.icell.PDM VGND 0.18855f
C8904 XA.XIR[4].XIC[14].icell.PDM VGND 0.18809f
C8905 XA.XIR[4].XIC[13].icell.PDM VGND 0.18809f
C8906 XA.XIR[4].XIC[12].icell.PDM VGND 0.18809f
C8907 XA.XIR[4].XIC[11].icell.PDM VGND 0.18809f
C8908 XA.XIR[4].XIC[10].icell.PDM VGND 0.18809f
C8909 XA.XIR[4].XIC[9].icell.PDM VGND 0.18809f
C8910 XA.XIR[4].XIC[8].icell.PDM VGND 0.18809f
C8911 XA.XIR[4].XIC[7].icell.PDM VGND 0.18809f
C8912 XA.XIR[4].XIC[6].icell.PDM VGND 0.18809f
C8913 XA.XIR[4].XIC[5].icell.PDM VGND 0.18809f
C8914 XA.XIR[4].XIC[4].icell.PDM VGND 0.18809f
C8915 XA.XIR[4].XIC[3].icell.PDM VGND 0.18809f
C8916 XA.XIR[4].XIC[2].icell.PDM VGND 0.18809f
C8917 XA.XIR[4].XIC[1].icell.PDM VGND 0.18809f
C8918 XA.XIR[4].XIC[0].icell.PDM VGND 0.18817f
C8919 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C8920 XThR.Tn[4] VGND 14.03736f
C8921 a_n1049_6405# VGND 0.02935f
C8922 a_n1319_6405# VGND 0.00166f
C8923 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C8924 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C8925 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.608f
C8926 XA.XIR[3].XIC_15.icell.SM VGND 0.00474f
C8927 XA.XIR[3].XIC_dummy_right.icell.PUM VGND 0.00215f
C8928 XA.XIR[3].XIC_15.icell.Ien VGND 0.37063f
C8929 XA.XIR[3].XIC[14].icell.SM VGND 0.00502f
C8930 XA.XIR[3].XIC_15.icell.PUM VGND 0.00282f
C8931 XA.XIR[3].XIC[14].icell.Ien VGND 0.37144f
C8932 XA.XIR[3].XIC[13].icell.SM VGND 0.00502f
C8933 XA.XIR[3].XIC[14].icell.PUM VGND 0.00293f
C8934 XA.XIR[3].XIC[13].icell.Ien VGND 0.37144f
C8935 XA.XIR[3].XIC[12].icell.SM VGND 0.00502f
C8936 XA.XIR[3].XIC[13].icell.PUM VGND 0.00293f
C8937 XA.XIR[3].XIC[12].icell.Ien VGND 0.37144f
C8938 XA.XIR[3].XIC[11].icell.SM VGND 0.00502f
C8939 XA.XIR[3].XIC[12].icell.PUM VGND 0.00293f
C8940 XA.XIR[3].XIC[11].icell.Ien VGND 0.37144f
C8941 XA.XIR[3].XIC[10].icell.SM VGND 0.00502f
C8942 XA.XIR[3].XIC[11].icell.PUM VGND 0.00293f
C8943 XA.XIR[3].XIC[10].icell.Ien VGND 0.37144f
C8944 XA.XIR[3].XIC[9].icell.SM VGND 0.00502f
C8945 XA.XIR[3].XIC[10].icell.PUM VGND 0.00293f
C8946 XA.XIR[3].XIC[9].icell.Ien VGND 0.37144f
C8947 XA.XIR[3].XIC[8].icell.SM VGND 0.00502f
C8948 XA.XIR[3].XIC[9].icell.PUM VGND 0.00293f
C8949 XA.XIR[3].XIC[8].icell.Ien VGND 0.37144f
C8950 XA.XIR[3].XIC[7].icell.SM VGND 0.00502f
C8951 XA.XIR[3].XIC[8].icell.PUM VGND 0.00293f
C8952 XA.XIR[3].XIC[7].icell.Ien VGND 0.37144f
C8953 XA.XIR[3].XIC[6].icell.SM VGND 0.00502f
C8954 XA.XIR[3].XIC[7].icell.PUM VGND 0.00293f
C8955 XA.XIR[3].XIC[6].icell.Ien VGND 0.37144f
C8956 XA.XIR[3].XIC[5].icell.SM VGND 0.00502f
C8957 XA.XIR[3].XIC[6].icell.PUM VGND 0.00293f
C8958 XA.XIR[3].XIC[5].icell.Ien VGND 0.37144f
C8959 XA.XIR[3].XIC[4].icell.SM VGND 0.00502f
C8960 XA.XIR[3].XIC[5].icell.PUM VGND 0.00293f
C8961 XA.XIR[3].XIC[4].icell.Ien VGND 0.37144f
C8962 XA.XIR[3].XIC[3].icell.SM VGND 0.00502f
C8963 XA.XIR[3].XIC[4].icell.PUM VGND 0.00293f
C8964 XA.XIR[3].XIC[3].icell.Ien VGND 0.37144f
C8965 XA.XIR[3].XIC[2].icell.SM VGND 0.00502f
C8966 XA.XIR[3].XIC[3].icell.PUM VGND 0.00293f
C8967 XA.XIR[3].XIC[2].icell.Ien VGND 0.37144f
C8968 XA.XIR[3].XIC[1].icell.SM VGND 0.00502f
C8969 XThR.XTB5.Y VGND 1.32753f
C8970 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80611f
C8971 XA.XIR[3].XIC[2].icell.PUM VGND 0.00293f
C8972 XA.XIR[3].XIC[1].icell.Ien VGND 0.37144f
C8973 XA.XIR[3].XIC[0].icell.SM VGND 0.00502f
C8974 XA.XIR[3].XIC[1].icell.PUM VGND 0.00293f
C8975 XA.XIR[3].XIC[0].icell.Ien VGND 0.37178f
C8976 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01044f
C8977 XA.XIR[3].XIC[0].icell.PUM VGND 0.00516f
C8978 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57425f
C8979 a_n1049_6699# VGND 0.02979f
C8980 XA.XIR[3].XIC_dummy_left.icell.PUM VGND 0.00215f
C8981 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C8982 XA.XIR[3].XIC_15.icell.PDM VGND 0.18855f
C8983 XA.XIR[3].XIC[14].icell.PDM VGND 0.18809f
C8984 XA.XIR[3].XIC[13].icell.PDM VGND 0.18809f
C8985 XA.XIR[3].XIC[12].icell.PDM VGND 0.18809f
C8986 XA.XIR[3].XIC[11].icell.PDM VGND 0.18809f
C8987 XA.XIR[3].XIC[10].icell.PDM VGND 0.18809f
C8988 XA.XIR[3].XIC[9].icell.PDM VGND 0.18809f
C8989 XA.XIR[3].XIC[8].icell.PDM VGND 0.18809f
C8990 XA.XIR[3].XIC[7].icell.PDM VGND 0.18809f
C8991 XA.XIR[3].XIC[6].icell.PDM VGND 0.18809f
C8992 XA.XIR[3].XIC[5].icell.PDM VGND 0.18809f
C8993 XA.XIR[3].XIC[4].icell.PDM VGND 0.18809f
C8994 XA.XIR[3].XIC[3].icell.PDM VGND 0.18809f
C8995 XA.XIR[3].XIC[2].icell.PDM VGND 0.18809f
C8996 XA.XIR[3].XIC[1].icell.PDM VGND 0.18809f
C8997 XA.XIR[3].XIC[0].icell.PDM VGND 0.18817f
C8998 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C8999 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C9000 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C9001 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.608f
C9002 XA.XIR[2].XIC_15.icell.SM VGND 0.00474f
C9003 XA.XIR[2].XIC_dummy_right.icell.PUM VGND 0.00215f
C9004 XA.XIR[2].XIC_15.icell.Ien VGND 0.37063f
C9005 XA.XIR[2].XIC[14].icell.SM VGND 0.00502f
C9006 XA.XIR[2].XIC_15.icell.PUM VGND 0.00282f
C9007 XA.XIR[2].XIC[14].icell.Ien VGND 0.37144f
C9008 XA.XIR[2].XIC[13].icell.SM VGND 0.00502f
C9009 XA.XIR[2].XIC[14].icell.PUM VGND 0.00293f
C9010 XA.XIR[2].XIC[13].icell.Ien VGND 0.37144f
C9011 XA.XIR[2].XIC[12].icell.SM VGND 0.00502f
C9012 XA.XIR[2].XIC[13].icell.PUM VGND 0.00293f
C9013 XA.XIR[2].XIC[12].icell.Ien VGND 0.37144f
C9014 XA.XIR[2].XIC[11].icell.SM VGND 0.00502f
C9015 XA.XIR[2].XIC[12].icell.PUM VGND 0.00293f
C9016 XA.XIR[2].XIC[11].icell.Ien VGND 0.37144f
C9017 XA.XIR[2].XIC[10].icell.SM VGND 0.00502f
C9018 XA.XIR[2].XIC[11].icell.PUM VGND 0.00293f
C9019 XA.XIR[2].XIC[10].icell.Ien VGND 0.37144f
C9020 XA.XIR[2].XIC[9].icell.SM VGND 0.00502f
C9021 XA.XIR[2].XIC[10].icell.PUM VGND 0.00293f
C9022 XA.XIR[2].XIC[9].icell.Ien VGND 0.37144f
C9023 XA.XIR[2].XIC[8].icell.SM VGND 0.00502f
C9024 XA.XIR[2].XIC[9].icell.PUM VGND 0.00293f
C9025 XA.XIR[2].XIC[8].icell.Ien VGND 0.37144f
C9026 XA.XIR[2].XIC[7].icell.SM VGND 0.00502f
C9027 XA.XIR[2].XIC[8].icell.PUM VGND 0.00293f
C9028 XA.XIR[2].XIC[7].icell.Ien VGND 0.37144f
C9029 XA.XIR[2].XIC[6].icell.SM VGND 0.00502f
C9030 XA.XIR[2].XIC[7].icell.PUM VGND 0.00293f
C9031 XA.XIR[2].XIC[6].icell.Ien VGND 0.37144f
C9032 XA.XIR[2].XIC[5].icell.SM VGND 0.00502f
C9033 XA.XIR[2].XIC[6].icell.PUM VGND 0.00293f
C9034 XA.XIR[2].XIC[5].icell.Ien VGND 0.37144f
C9035 XA.XIR[2].XIC[4].icell.SM VGND 0.00502f
C9036 XA.XIR[2].XIC[5].icell.PUM VGND 0.00293f
C9037 XA.XIR[2].XIC[4].icell.Ien VGND 0.37144f
C9038 XA.XIR[2].XIC[3].icell.SM VGND 0.00502f
C9039 XA.XIR[2].XIC[4].icell.PUM VGND 0.00293f
C9040 XA.XIR[2].XIC[3].icell.Ien VGND 0.37144f
C9041 XA.XIR[2].XIC[2].icell.SM VGND 0.00502f
C9042 XA.XIR[2].XIC[3].icell.PUM VGND 0.00293f
C9043 XA.XIR[2].XIC[2].icell.Ien VGND 0.37144f
C9044 XA.XIR[2].XIC[1].icell.SM VGND 0.00502f
C9045 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80825f
C9046 XA.XIR[2].XIC[2].icell.PUM VGND 0.00293f
C9047 XA.XIR[2].XIC[1].icell.Ien VGND 0.37144f
C9048 XA.XIR[2].XIC[0].icell.SM VGND 0.00502f
C9049 XThR.Tn[3] VGND 13.98256f
C9050 XThR.XTB4.Y VGND 1.76953f
C9051 XA.XIR[2].XIC[1].icell.PUM VGND 0.00293f
C9052 XA.XIR[2].XIC[0].icell.Ien VGND 0.37178f
C9053 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01044f
C9054 XA.XIR[2].XIC[0].icell.PUM VGND 0.00516f
C9055 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57559f
C9056 a_n1335_7243# VGND 0.00179f
C9057 XA.XIR[2].XIC_dummy_left.icell.PUM VGND 0.00215f
C9058 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C9059 XA.XIR[2].XIC_15.icell.PDM VGND 0.18855f
C9060 XA.XIR[2].XIC[14].icell.PDM VGND 0.18809f
C9061 XA.XIR[2].XIC[13].icell.PDM VGND 0.18809f
C9062 XA.XIR[2].XIC[12].icell.PDM VGND 0.18809f
C9063 XA.XIR[2].XIC[11].icell.PDM VGND 0.18809f
C9064 XA.XIR[2].XIC[10].icell.PDM VGND 0.18809f
C9065 XA.XIR[2].XIC[9].icell.PDM VGND 0.18809f
C9066 XA.XIR[2].XIC[8].icell.PDM VGND 0.18809f
C9067 XA.XIR[2].XIC[7].icell.PDM VGND 0.18809f
C9068 XA.XIR[2].XIC[6].icell.PDM VGND 0.18809f
C9069 XA.XIR[2].XIC[5].icell.PDM VGND 0.18809f
C9070 XA.XIR[2].XIC[4].icell.PDM VGND 0.18809f
C9071 XA.XIR[2].XIC[3].icell.PDM VGND 0.18809f
C9072 XA.XIR[2].XIC[2].icell.PDM VGND 0.18809f
C9073 XA.XIR[2].XIC[1].icell.PDM VGND 0.18809f
C9074 XA.XIR[2].XIC[0].icell.PDM VGND 0.18817f
C9075 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C9076 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C9077 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C9078 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.608f
C9079 XA.XIR[1].XIC_15.icell.SM VGND 0.00474f
C9080 XA.XIR[1].XIC_dummy_right.icell.PUM VGND 0.00215f
C9081 XA.XIR[1].XIC_15.icell.Ien VGND 0.37063f
C9082 XA.XIR[1].XIC[14].icell.SM VGND 0.00502f
C9083 XA.XIR[1].XIC_15.icell.PUM VGND 0.00282f
C9084 XA.XIR[1].XIC[14].icell.Ien VGND 0.37144f
C9085 XA.XIR[1].XIC[13].icell.SM VGND 0.00502f
C9086 XA.XIR[1].XIC[14].icell.PUM VGND 0.00293f
C9087 XA.XIR[1].XIC[13].icell.Ien VGND 0.37144f
C9088 XA.XIR[1].XIC[12].icell.SM VGND 0.00502f
C9089 XA.XIR[1].XIC[13].icell.PUM VGND 0.00293f
C9090 XA.XIR[1].XIC[12].icell.Ien VGND 0.37144f
C9091 XA.XIR[1].XIC[11].icell.SM VGND 0.00502f
C9092 XA.XIR[1].XIC[12].icell.PUM VGND 0.00293f
C9093 XA.XIR[1].XIC[11].icell.Ien VGND 0.37144f
C9094 XA.XIR[1].XIC[10].icell.SM VGND 0.00502f
C9095 XA.XIR[1].XIC[11].icell.PUM VGND 0.00293f
C9096 XA.XIR[1].XIC[10].icell.Ien VGND 0.37144f
C9097 XA.XIR[1].XIC[9].icell.SM VGND 0.00502f
C9098 XA.XIR[1].XIC[10].icell.PUM VGND 0.00293f
C9099 XA.XIR[1].XIC[9].icell.Ien VGND 0.37144f
C9100 XA.XIR[1].XIC[8].icell.SM VGND 0.00502f
C9101 XA.XIR[1].XIC[9].icell.PUM VGND 0.00293f
C9102 XA.XIR[1].XIC[8].icell.Ien VGND 0.37144f
C9103 XA.XIR[1].XIC[7].icell.SM VGND 0.00502f
C9104 XA.XIR[1].XIC[8].icell.PUM VGND 0.00293f
C9105 XA.XIR[1].XIC[7].icell.Ien VGND 0.37144f
C9106 XA.XIR[1].XIC[6].icell.SM VGND 0.00502f
C9107 XA.XIR[1].XIC[7].icell.PUM VGND 0.00293f
C9108 XA.XIR[1].XIC[6].icell.Ien VGND 0.37144f
C9109 XA.XIR[1].XIC[5].icell.SM VGND 0.00502f
C9110 XA.XIR[1].XIC[6].icell.PUM VGND 0.00293f
C9111 XA.XIR[1].XIC[5].icell.Ien VGND 0.37144f
C9112 XA.XIR[1].XIC[4].icell.SM VGND 0.00502f
C9113 XA.XIR[1].XIC[5].icell.PUM VGND 0.00293f
C9114 XA.XIR[1].XIC[4].icell.Ien VGND 0.37144f
C9115 XA.XIR[1].XIC[3].icell.SM VGND 0.00502f
C9116 XA.XIR[1].XIC[4].icell.PUM VGND 0.00293f
C9117 XA.XIR[1].XIC[3].icell.Ien VGND 0.37144f
C9118 XA.XIR[1].XIC[2].icell.SM VGND 0.00502f
C9119 XA.XIR[1].XIC[3].icell.PUM VGND 0.00293f
C9120 XA.XIR[1].XIC[2].icell.Ien VGND 0.37144f
C9121 XA.XIR[1].XIC[1].icell.SM VGND 0.00502f
C9122 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80611f
C9123 XA.XIR[1].XIC[2].icell.PUM VGND 0.00293f
C9124 XA.XIR[1].XIC[1].icell.Ien VGND 0.37144f
C9125 XA.XIR[1].XIC[0].icell.SM VGND 0.00502f
C9126 XThR.Tn[2] VGND 14.03476f
C9127 a_n1049_7493# VGND 0.02484f
C9128 XThR.XTB3.Y VGND 2.09162f
C9129 XThR.XTB7.A VGND 1.95537f
C9130 XA.XIR[1].XIC[1].icell.PUM VGND 0.00293f
C9131 XA.XIR[1].XIC[0].icell.Ien VGND 0.37178f
C9132 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01044f
C9133 XA.XIR[1].XIC[0].icell.PUM VGND 0.00516f
C9134 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57379f
C9135 XA.XIR[1].XIC_dummy_left.icell.PUM VGND 0.00215f
C9136 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C9137 XA.XIR[1].XIC_15.icell.PDM VGND 0.18855f
C9138 XA.XIR[1].XIC[14].icell.PDM VGND 0.18809f
C9139 XA.XIR[1].XIC[13].icell.PDM VGND 0.18809f
C9140 XA.XIR[1].XIC[12].icell.PDM VGND 0.18809f
C9141 XA.XIR[1].XIC[11].icell.PDM VGND 0.18809f
C9142 XA.XIR[1].XIC[10].icell.PDM VGND 0.18809f
C9143 XA.XIR[1].XIC[9].icell.PDM VGND 0.18809f
C9144 XA.XIR[1].XIC[8].icell.PDM VGND 0.18809f
C9145 XA.XIR[1].XIC[7].icell.PDM VGND 0.18809f
C9146 XA.XIR[1].XIC[6].icell.PDM VGND 0.18809f
C9147 XA.XIR[1].XIC[5].icell.PDM VGND 0.18809f
C9148 XA.XIR[1].XIC[4].icell.PDM VGND 0.18809f
C9149 XA.XIR[1].XIC[3].icell.PDM VGND 0.18809f
C9150 XA.XIR[1].XIC[2].icell.PDM VGND 0.18809f
C9151 XA.XIR[1].XIC[1].icell.PDM VGND 0.18809f
C9152 XA.XIR[1].XIC[0].icell.PDM VGND 0.18817f
C9153 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C9154 a_n1049_7787# VGND 0.03397f
C9155 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87403f
C9156 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C9157 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61779f
C9158 XA.XIR[0].XIC_15.icell.SM VGND 0.00474f
C9159 XA.XIR[0].XIC_dummy_right.icell.PUM VGND 0.00207f
C9160 XA.XIR[0].XIC_15.icell.Ien VGND 0.37673f
C9161 XA.XIR[0].XIC[14].icell.SM VGND 0.00624f
C9162 XA.XIR[0].XIC_15.icell.PUM VGND 0.00468f
C9163 XA.XIR[0].XIC[14].icell.Ien VGND 0.38432f
C9164 XA.XIR[0].XIC[13].icell.SM VGND 0.00624f
C9165 XA.XIR[0].XIC[14].icell.PUM VGND 0.00392f
C9166 XA.XIR[0].XIC[13].icell.Ien VGND 0.38436f
C9167 XA.XIR[0].XIC[12].icell.SM VGND 0.00624f
C9168 XA.XIR[0].XIC[13].icell.PUM VGND 0.00397f
C9169 XA.XIR[0].XIC[12].icell.Ien VGND 0.381f
C9170 XA.XIR[0].XIC[11].icell.SM VGND 0.00624f
C9171 XA.XIR[0].XIC[12].icell.PUM VGND 0.00392f
C9172 XA.XIR[0].XIC[11].icell.Ien VGND 0.38167f
C9173 XA.XIR[0].XIC[10].icell.SM VGND 0.00624f
C9174 XA.XIR[0].XIC[11].icell.PUM VGND 0.00392f
C9175 XA.XIR[0].XIC[10].icell.Ien VGND 0.38301f
C9176 XA.XIR[0].XIC[9].icell.SM VGND 0.00624f
C9177 XA.XIR[0].XIC[10].icell.PUM VGND 0.00392f
C9178 XA.XIR[0].XIC[9].icell.Ien VGND 0.38128f
C9179 XA.XIR[0].XIC[8].icell.SM VGND 0.00624f
C9180 XA.XIR[0].XIC[9].icell.PUM VGND 0.00392f
C9181 XA.XIR[0].XIC[8].icell.Ien VGND 0.38176f
C9182 XA.XIR[0].XIC[7].icell.SM VGND 0.00624f
C9183 XA.XIR[0].XIC[8].icell.PUM VGND 0.00392f
C9184 XA.XIR[0].XIC[7].icell.Ien VGND 0.382f
C9185 XA.XIR[0].XIC[6].icell.SM VGND 0.00624f
C9186 XA.XIR[0].XIC[7].icell.PUM VGND 0.00392f
C9187 XA.XIR[0].XIC[6].icell.Ien VGND 0.38192f
C9188 XA.XIR[0].XIC[5].icell.SM VGND 0.00624f
C9189 XA.XIR[0].XIC[6].icell.PUM VGND 0.00403f
C9190 XA.XIR[0].XIC[5].icell.Ien VGND 0.38091f
C9191 XA.XIR[0].XIC[4].icell.SM VGND 0.00624f
C9192 XA.XIR[0].XIC[5].icell.PUM VGND 0.00392f
C9193 XA.XIR[0].XIC[4].icell.Ien VGND 0.38104f
C9194 XA.XIR[0].XIC[3].icell.SM VGND 0.00624f
C9195 XA.XIR[0].XIC[4].icell.PUM VGND 0.00392f
C9196 XA.XIR[0].XIC[3].icell.Ien VGND 0.38229f
C9197 XA.XIR[0].XIC[2].icell.SM VGND 0.00624f
C9198 XA.XIR[0].XIC[3].icell.PUM VGND 0.00392f
C9199 XA.XIR[0].XIC[2].icell.Ien VGND 0.38432f
C9200 XA.XIR[0].XIC[1].icell.SM VGND 0.00624f
C9201 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83227f
C9202 XA.XIR[0].XIC[2].icell.PUM VGND 0.00392f
C9203 XA.XIR[0].XIC[1].icell.Ien VGND 0.38432f
C9204 XA.XIR[0].XIC[0].icell.SM VGND 0.00624f
C9205 XA.XIR[0].XIC[1].icell.PUM VGND 0.00394f
C9206 XA.XIR[0].XIC[0].icell.Ien VGND 0.38384f
C9207 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01044f
C9208 XThR.Tn[1] VGND 14.06885f
C9209 a_n1335_8107# VGND 0.00163f
C9210 XThR.XTB2.Y VGND 1.47619f
C9211 XThR.XTB6.A VGND 0.95635f
C9212 XA.XIR[0].XIC[0].icell.PUM VGND 0.00623f
C9213 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58434f
C9214 XA.XIR[0].XIC_dummy_left.icell.PUM VGND 0.00355f
C9215 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.251f
C9216 XA.XIR[0].XIC_15.icell.PDM VGND 0.20765f
C9217 XA.XIR[0].XIC[14].icell.PDM VGND 0.24599f
C9218 XA.XIR[0].XIC[13].icell.PDM VGND 0.24583f
C9219 XA.XIR[0].XIC[12].icell.PDM VGND 0.24144f
C9220 XA.XIR[0].XIC[11].icell.PDM VGND 0.24182f
C9221 XA.XIR[0].XIC[10].icell.PDM VGND 0.24172f
C9222 XA.XIR[0].XIC[9].icell.PDM VGND 0.24144f
C9223 XA.XIR[0].XIC[8].icell.PDM VGND 0.24144f
C9224 XA.XIR[0].XIC[7].icell.PDM VGND 0.24388f
C9225 XA.XIR[0].XIC[6].icell.PDM VGND 0.24108f
C9226 XA.XIR[0].XIC[5].icell.PDM VGND 0.24297f
C9227 XA.XIR[0].XIC[4].icell.PDM VGND 0.24156f
C9228 XA.XIR[0].XIC[3].icell.PDM VGND 0.24455f
C9229 XA.XIR[0].XIC[2].icell.PDM VGND 0.24578f
C9230 XA.XIR[0].XIC[1].icell.PDM VGND 0.24578f
C9231 XA.XIR[0].XIC[0].icell.PDM VGND 0.24457f
C9232 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.24577f
C9233 a_n1335_8331# VGND 0.00203f
C9234 XThR.Tn[0] VGND 14.40233f
C9235 a_n1049_8581# VGND 0.04333f
C9236 XThR.XTBN.Y VGND 7.53702f
C9237 XThR.XTB1.Y VGND 1.80911f
C9238 XThR.XTB7.B VGND 2.61063f
C9239 XThR.XTB5.A VGND 1.75777f
C9240 XThC.Tn[14] VGND 9.98563f
C9241 XThC.Tn[13] VGND 9.79145f
C9242 XThC.Tn[12] VGND 9.63534f
C9243 XThC.Tn[11] VGND 9.46598f
C9244 XThC.Tn[10] VGND 9.29745f
C9245 XThC.Tn[9] VGND 9.27278f
C9246 XThC.Tn[8] VGND 9.24802f
C9247 a_10915_9569# VGND 0.55837f
C9248 a_10051_9569# VGND 0.55761f
C9249 a_9827_9569# VGND 0.54461f
C9250 a_8963_9569# VGND 0.55448f
C9251 a_8739_9569# VGND 0.55288f
C9252 a_7875_9569# VGND 0.55432f
C9253 a_7651_9569# VGND 0.55717f
C9254 XThC.Tn[7] VGND 10.56205f
C9255 XThC.Tn[6] VGND 10.35711f
C9256 XThC.Tn[5] VGND 10.62787f
C9257 XThC.Tn[4] VGND 10.6808f
C9258 XThC.Tn[3] VGND 9.9249f
C9259 XThC.Tn[2] VGND 10.45573f
C9260 XThC.Tn[1] VGND 10.32305f
C9261 XThC.Tn[0] VGND 10.84166f
C9262 a_6243_9615# VGND 0.0299f
C9263 a_5949_9615# VGND 0.03432f
C9264 a_5155_9615# VGND 0.03615f
C9265 a_4861_9615# VGND 0.03632f
C9266 a_4067_9615# VGND 0.03071f
C9267 a_3773_9615# VGND 0.03867f
C9268 a_2979_9615# VGND 0.04107f
C9269 a_8739_10571# VGND 0.00194f
C9270 XThC.XTBN.Y VGND 7.90394f
C9271 XThC.XTB7.Y VGND 1.36247f
C9272 XThC.XTB6.Y VGND 1.3829f
C9273 a_5155_10571# VGND 0.00165f
C9274 XThC.XTB7.B VGND 2.73083f
C9275 XThC.XTB5.Y VGND 1.32591f
C9276 XThC.XTBN.A VGND 1.23171f
C9277 a_4387_10575# VGND 0.00179f
C9278 a_3523_10575# VGND 0.00163f
C9279 a_3299_10575# VGND 0.00202f
C9280 XThC.XTB4.Y VGND 1.69875f
C9281 XThC.XTB3.Y VGND 1.96765f
C9282 XThC.XTB7.A VGND 1.96056f
C9283 XThC.XTB6.A VGND 0.95757f
C9284 XThC.XTB2.Y VGND 1.47589f
C9285 XThC.XTB1.Y VGND 1.77676f
C9286 XThC.XTB5.A VGND 1.75974f
C9287 bias[0].t0 VGND 0.94587f
C9288 XThR.XTB3.Y.t1 VGND 0.06176f
C9289 XThR.XTB3.Y.n0 VGND 0.01521f
C9290 XThR.XTB3.Y.t8 VGND 0.04903f
C9291 XThR.XTB3.Y.t15 VGND 0.02889f
C9292 XThR.XTB3.Y.t13 VGND 0.04903f
C9293 XThR.XTB3.Y.t6 VGND 0.02889f
C9294 XThR.XTB3.Y.t9 VGND 0.04903f
C9295 XThR.XTB3.Y.t17 VGND 0.02889f
C9296 XThR.XTB3.Y.n1 VGND 0.08226f
C9297 XThR.XTB3.Y.n2 VGND 0.08688f
C9298 XThR.XTB3.Y.n3 VGND 0.03573f
C9299 XThR.XTB3.Y.n4 VGND 0.0707f
C9300 XThR.XTB3.Y.t12 VGND 0.04903f
C9301 XThR.XTB3.Y.t4 VGND 0.02889f
C9302 XThR.XTB3.Y.n5 VGND 0.06608f
C9303 XThR.XTB3.Y.n6 VGND 0.03236f
C9304 XThR.XTB3.Y.n7 VGND 0.02685f
C9305 XThR.XTB3.Y.t18 VGND 0.04903f
C9306 XThR.XTB3.Y.t5 VGND 0.02889f
C9307 XThR.XTB3.Y.n8 VGND 0.03005f
C9308 XThR.XTB3.Y.t7 VGND 0.04903f
C9309 XThR.XTB3.Y.t10 VGND 0.02889f
C9310 XThR.XTB3.Y.n9 VGND 0.05992f
C9311 XThR.XTB3.Y.t11 VGND 0.04903f
C9312 XThR.XTB3.Y.t16 VGND 0.02889f
C9313 XThR.XTB3.Y.n10 VGND 0.06454f
C9314 XThR.XTB3.Y.n11 VGND 0.03645f
C9315 XThR.XTB3.Y.n12 VGND 0.06034f
C9316 XThR.XTB3.Y.n13 VGND 0.03128f
C9317 XThR.XTB3.Y.n14 VGND 0.02851f
C9318 XThR.XTB3.Y.n15 VGND 0.06454f
C9319 XThR.XTB3.Y.t14 VGND 0.04903f
C9320 XThR.XTB3.Y.t3 VGND 0.02889f
C9321 XThR.XTB3.Y.n16 VGND 0.05838f
C9322 XThR.XTB3.Y.n17 VGND 0.03236f
C9323 XThR.XTB3.Y.n18 VGND 0.04707f
C9324 XThR.XTB3.Y.n19 VGND 1.31347f
C9325 XThR.XTB3.Y.t0 VGND 0.03152f
C9326 XThR.XTB3.Y.t2 VGND 0.03152f
C9327 XThR.XTB3.Y.n20 VGND 0.06766f
C9328 XThR.XTB3.Y.n21 VGND 0.157f
C9329 XThR.XTB3.Y.n22 VGND 0.03296f
C9330 XThR.XTB1.Y.t1 VGND 0.03165f
C9331 XThR.XTB1.Y.n0 VGND 0.0078f
C9332 XThR.XTB1.Y.t8 VGND 0.02512f
C9333 XThR.XTB1.Y.t15 VGND 0.0148f
C9334 XThR.XTB1.Y.t14 VGND 0.02512f
C9335 XThR.XTB1.Y.t7 VGND 0.0148f
C9336 XThR.XTB1.Y.t10 VGND 0.02512f
C9337 XThR.XTB1.Y.t18 VGND 0.0148f
C9338 XThR.XTB1.Y.n1 VGND 0.04215f
C9339 XThR.XTB1.Y.n2 VGND 0.04452f
C9340 XThR.XTB1.Y.n3 VGND 0.01831f
C9341 XThR.XTB1.Y.n4 VGND 0.03623f
C9342 XThR.XTB1.Y.t13 VGND 0.02512f
C9343 XThR.XTB1.Y.t4 VGND 0.0148f
C9344 XThR.XTB1.Y.n5 VGND 0.03386f
C9345 XThR.XTB1.Y.n6 VGND 0.01658f
C9346 XThR.XTB1.Y.n7 VGND 0.01376f
C9347 XThR.XTB1.Y.t6 VGND 0.02512f
C9348 XThR.XTB1.Y.t11 VGND 0.0148f
C9349 XThR.XTB1.Y.n8 VGND 0.0154f
C9350 XThR.XTB1.Y.t12 VGND 0.02512f
C9351 XThR.XTB1.Y.t16 VGND 0.0148f
C9352 XThR.XTB1.Y.n9 VGND 0.0307f
C9353 XThR.XTB1.Y.t17 VGND 0.02512f
C9354 XThR.XTB1.Y.t5 VGND 0.0148f
C9355 XThR.XTB1.Y.n10 VGND 0.03307f
C9356 XThR.XTB1.Y.n11 VGND 0.01868f
C9357 XThR.XTB1.Y.n12 VGND 0.03092f
C9358 XThR.XTB1.Y.n13 VGND 0.01603f
C9359 XThR.XTB1.Y.n14 VGND 0.01461f
C9360 XThR.XTB1.Y.n15 VGND 0.03307f
C9361 XThR.XTB1.Y.t3 VGND 0.02512f
C9362 XThR.XTB1.Y.t9 VGND 0.0148f
C9363 XThR.XTB1.Y.n16 VGND 0.02991f
C9364 XThR.XTB1.Y.n17 VGND 0.01658f
C9365 XThR.XTB1.Y.n18 VGND 0.02412f
C9366 XThR.XTB1.Y.n19 VGND 0.75219f
C9367 XThR.XTB1.Y.t0 VGND 0.01615f
C9368 XThR.XTB1.Y.t2 VGND 0.01615f
C9369 XThR.XTB1.Y.n20 VGND 0.03467f
C9370 XThR.XTB1.Y.n21 VGND 0.08068f
C9371 XThR.XTB1.Y.n22 VGND 0.01689f
C9372 XThR.XTB4.Y.t8 VGND 0.02956f
C9373 XThR.XTB4.Y.t15 VGND 0.05016f
C9374 XThR.XTB4.Y.t16 VGND 0.02956f
C9375 XThR.XTB4.Y.t5 VGND 0.05016f
C9376 XThR.XTB4.Y.t10 VGND 0.02956f
C9377 XThR.XTB4.Y.t17 VGND 0.05016f
C9378 XThR.XTB4.Y.n0 VGND 0.08416f
C9379 XThR.XTB4.Y.n1 VGND 0.08889f
C9380 XThR.XTB4.Y.n2 VGND 0.03656f
C9381 XThR.XTB4.Y.n3 VGND 0.07234f
C9382 XThR.XTB4.Y.t13 VGND 0.02956f
C9383 XThR.XTB4.Y.t4 VGND 0.05016f
C9384 XThR.XTB4.Y.n4 VGND 0.06761f
C9385 XThR.XTB4.Y.n5 VGND 0.0331f
C9386 XThR.XTB4.Y.n6 VGND 0.01685f
C9387 XThR.XTB4.Y.n7 VGND 0.05355f
C9388 XThR.XTB4.Y.n8 VGND 0.64921f
C9389 XThR.XTB4.Y.t14 VGND 0.02956f
C9390 XThR.XTB4.Y.t7 VGND 0.05016f
C9391 XThR.XTB4.Y.n9 VGND 0.03074f
C9392 XThR.XTB4.Y.t3 VGND 0.02956f
C9393 XThR.XTB4.Y.t12 VGND 0.05016f
C9394 XThR.XTB4.Y.n10 VGND 0.0613f
C9395 XThR.XTB4.Y.t9 VGND 0.02956f
C9396 XThR.XTB4.Y.t2 VGND 0.05016f
C9397 XThR.XTB4.Y.n11 VGND 0.06603f
C9398 XThR.XTB4.Y.n12 VGND 0.03729f
C9399 XThR.XTB4.Y.n13 VGND 0.06174f
C9400 XThR.XTB4.Y.n14 VGND 0.03201f
C9401 XThR.XTB4.Y.n15 VGND 0.02916f
C9402 XThR.XTB4.Y.n16 VGND 0.06603f
C9403 XThR.XTB4.Y.t11 VGND 0.02956f
C9404 XThR.XTB4.Y.t6 VGND 0.05016f
C9405 XThR.XTB4.Y.n17 VGND 0.05972f
C9406 XThR.XTB4.Y.n18 VGND 0.0331f
C9407 XThR.XTB4.Y.n19 VGND 0.05647f
C9408 XThR.XTB4.Y.n20 VGND 1.3092f
C9409 XThR.XTB4.Y.t1 VGND 0.06491f
C9410 XThR.XTB4.Y.n21 VGND 0.12281f
C9411 XThR.XTB4.Y.n22 VGND 0.02892f
C9412 XThR.XTB4.Y.t0 VGND 0.11919f
C9413 XThR.Tn[13].t2 VGND 0.02397f
C9414 XThR.Tn[13].t0 VGND 0.02397f
C9415 XThR.Tn[13].n0 VGND 0.05327f
C9416 XThR.Tn[13].t1 VGND 0.02397f
C9417 XThR.Tn[13].t3 VGND 0.02397f
C9418 XThR.Tn[13].n1 VGND 0.07277f
C9419 XThR.Tn[13].n2 VGND 0.24224f
C9420 XThR.Tn[13].t7 VGND 0.01558f
C9421 XThR.Tn[13].t5 VGND 0.01558f
C9422 XThR.Tn[13].n3 VGND 0.03885f
C9423 XThR.Tn[13].t6 VGND 0.01558f
C9424 XThR.Tn[13].t4 VGND 0.01558f
C9425 XThR.Tn[13].n4 VGND 0.03116f
C9426 XThR.Tn[13].n5 VGND 0.07837f
C9427 XThR.Tn[13].t72 VGND 0.01873f
C9428 XThR.Tn[13].t64 VGND 0.02051f
C9429 XThR.Tn[13].n6 VGND 0.05008f
C9430 XThR.Tn[13].n7 VGND 0.09621f
C9431 XThR.Tn[13].t28 VGND 0.01873f
C9432 XThR.Tn[13].t21 VGND 0.02051f
C9433 XThR.Tn[13].n8 VGND 0.05008f
C9434 XThR.Tn[13].t44 VGND 0.01867f
C9435 XThR.Tn[13].t12 VGND 0.02044f
C9436 XThR.Tn[13].n9 VGND 0.05211f
C9437 XThR.Tn[13].n10 VGND 0.03661f
C9438 XThR.Tn[13].n11 VGND 0.00669f
C9439 XThR.Tn[13].n12 VGND 0.11748f
C9440 XThR.Tn[13].t65 VGND 0.01873f
C9441 XThR.Tn[13].t57 VGND 0.02051f
C9442 XThR.Tn[13].n13 VGND 0.05008f
C9443 XThR.Tn[13].t19 VGND 0.01867f
C9444 XThR.Tn[13].t52 VGND 0.02044f
C9445 XThR.Tn[13].n14 VGND 0.05211f
C9446 XThR.Tn[13].n15 VGND 0.03661f
C9447 XThR.Tn[13].n16 VGND 0.00669f
C9448 XThR.Tn[13].n17 VGND 0.11748f
C9449 XThR.Tn[13].t22 VGND 0.01873f
C9450 XThR.Tn[13].t14 VGND 0.02051f
C9451 XThR.Tn[13].n18 VGND 0.05008f
C9452 XThR.Tn[13].t34 VGND 0.01867f
C9453 XThR.Tn[13].t70 VGND 0.02044f
C9454 XThR.Tn[13].n19 VGND 0.05211f
C9455 XThR.Tn[13].n20 VGND 0.03661f
C9456 XThR.Tn[13].n21 VGND 0.00669f
C9457 XThR.Tn[13].n22 VGND 0.11748f
C9458 XThR.Tn[13].t49 VGND 0.01873f
C9459 XThR.Tn[13].t39 VGND 0.02051f
C9460 XThR.Tn[13].n23 VGND 0.05008f
C9461 XThR.Tn[13].t66 VGND 0.01867f
C9462 XThR.Tn[13].t35 VGND 0.02044f
C9463 XThR.Tn[13].n24 VGND 0.05211f
C9464 XThR.Tn[13].n25 VGND 0.03661f
C9465 XThR.Tn[13].n26 VGND 0.00669f
C9466 XThR.Tn[13].n27 VGND 0.11748f
C9467 XThR.Tn[13].t24 VGND 0.01873f
C9468 XThR.Tn[13].t16 VGND 0.02051f
C9469 XThR.Tn[13].n28 VGND 0.05008f
C9470 XThR.Tn[13].t37 VGND 0.01867f
C9471 XThR.Tn[13].t71 VGND 0.02044f
C9472 XThR.Tn[13].n29 VGND 0.05211f
C9473 XThR.Tn[13].n30 VGND 0.03661f
C9474 XThR.Tn[13].n31 VGND 0.00669f
C9475 XThR.Tn[13].n32 VGND 0.11748f
C9476 XThR.Tn[13].t60 VGND 0.01873f
C9477 XThR.Tn[13].t30 VGND 0.02051f
C9478 XThR.Tn[13].n33 VGND 0.05008f
C9479 XThR.Tn[13].t13 VGND 0.01867f
C9480 XThR.Tn[13].t26 VGND 0.02044f
C9481 XThR.Tn[13].n34 VGND 0.05211f
C9482 XThR.Tn[13].n35 VGND 0.03661f
C9483 XThR.Tn[13].n36 VGND 0.00669f
C9484 XThR.Tn[13].n37 VGND 0.11748f
C9485 XThR.Tn[13].t29 VGND 0.01873f
C9486 XThR.Tn[13].t25 VGND 0.02051f
C9487 XThR.Tn[13].n38 VGND 0.05008f
C9488 XThR.Tn[13].t43 VGND 0.01867f
C9489 XThR.Tn[13].t18 VGND 0.02044f
C9490 XThR.Tn[13].n39 VGND 0.05211f
C9491 XThR.Tn[13].n40 VGND 0.03661f
C9492 XThR.Tn[13].n41 VGND 0.00669f
C9493 XThR.Tn[13].n42 VGND 0.11748f
C9494 XThR.Tn[13].t32 VGND 0.01873f
C9495 XThR.Tn[13].t38 VGND 0.02051f
C9496 XThR.Tn[13].n43 VGND 0.05008f
C9497 XThR.Tn[13].t48 VGND 0.01867f
C9498 XThR.Tn[13].t33 VGND 0.02044f
C9499 XThR.Tn[13].n44 VGND 0.05211f
C9500 XThR.Tn[13].n45 VGND 0.03661f
C9501 XThR.Tn[13].n46 VGND 0.00669f
C9502 XThR.Tn[13].n47 VGND 0.11748f
C9503 XThR.Tn[13].t51 VGND 0.01873f
C9504 XThR.Tn[13].t59 VGND 0.02051f
C9505 XThR.Tn[13].n48 VGND 0.05008f
C9506 XThR.Tn[13].t68 VGND 0.01867f
C9507 XThR.Tn[13].t53 VGND 0.02044f
C9508 XThR.Tn[13].n49 VGND 0.05211f
C9509 XThR.Tn[13].n50 VGND 0.03661f
C9510 XThR.Tn[13].n51 VGND 0.00669f
C9511 XThR.Tn[13].n52 VGND 0.11748f
C9512 XThR.Tn[13].t41 VGND 0.01873f
C9513 XThR.Tn[13].t17 VGND 0.02051f
C9514 XThR.Tn[13].n53 VGND 0.05008f
C9515 XThR.Tn[13].t58 VGND 0.01867f
C9516 XThR.Tn[13].t73 VGND 0.02044f
C9517 XThR.Tn[13].n54 VGND 0.05211f
C9518 XThR.Tn[13].n55 VGND 0.03661f
C9519 XThR.Tn[13].n56 VGND 0.00669f
C9520 XThR.Tn[13].n57 VGND 0.11748f
C9521 XThR.Tn[13].t63 VGND 0.01873f
C9522 XThR.Tn[13].t55 VGND 0.02051f
C9523 XThR.Tn[13].n58 VGND 0.05008f
C9524 XThR.Tn[13].t15 VGND 0.01867f
C9525 XThR.Tn[13].t45 VGND 0.02044f
C9526 XThR.Tn[13].n59 VGND 0.05211f
C9527 XThR.Tn[13].n60 VGND 0.03661f
C9528 XThR.Tn[13].n61 VGND 0.00669f
C9529 XThR.Tn[13].n62 VGND 0.11748f
C9530 XThR.Tn[13].t31 VGND 0.01873f
C9531 XThR.Tn[13].t27 VGND 0.02051f
C9532 XThR.Tn[13].n63 VGND 0.05008f
C9533 XThR.Tn[13].t46 VGND 0.01867f
C9534 XThR.Tn[13].t20 VGND 0.02044f
C9535 XThR.Tn[13].n64 VGND 0.05211f
C9536 XThR.Tn[13].n65 VGND 0.03661f
C9537 XThR.Tn[13].n66 VGND 0.00669f
C9538 XThR.Tn[13].n67 VGND 0.11748f
C9539 XThR.Tn[13].t50 VGND 0.01873f
C9540 XThR.Tn[13].t40 VGND 0.02051f
C9541 XThR.Tn[13].n68 VGND 0.05008f
C9542 XThR.Tn[13].t67 VGND 0.01867f
C9543 XThR.Tn[13].t36 VGND 0.02044f
C9544 XThR.Tn[13].n69 VGND 0.05211f
C9545 XThR.Tn[13].n70 VGND 0.03661f
C9546 XThR.Tn[13].n71 VGND 0.00669f
C9547 XThR.Tn[13].n72 VGND 0.11748f
C9548 XThR.Tn[13].t69 VGND 0.01873f
C9549 XThR.Tn[13].t62 VGND 0.02051f
C9550 XThR.Tn[13].n73 VGND 0.05008f
C9551 XThR.Tn[13].t23 VGND 0.01867f
C9552 XThR.Tn[13].t54 VGND 0.02044f
C9553 XThR.Tn[13].n74 VGND 0.05211f
C9554 XThR.Tn[13].n75 VGND 0.03661f
C9555 XThR.Tn[13].n76 VGND 0.00669f
C9556 XThR.Tn[13].n77 VGND 0.11748f
C9557 XThR.Tn[13].t42 VGND 0.01873f
C9558 XThR.Tn[13].t56 VGND 0.02051f
C9559 XThR.Tn[13].n78 VGND 0.05008f
C9560 XThR.Tn[13].t61 VGND 0.01867f
C9561 XThR.Tn[13].t47 VGND 0.02044f
C9562 XThR.Tn[13].n79 VGND 0.05211f
C9563 XThR.Tn[13].n80 VGND 0.03661f
C9564 XThR.Tn[13].n81 VGND 0.00669f
C9565 XThR.Tn[13].n82 VGND 0.11748f
C9566 XThR.Tn[13].n83 VGND 0.10676f
C9567 XThR.Tn[13].n84 VGND 0.41858f
C9568 XThR.Tn[13].t10 VGND 0.02397f
C9569 XThR.Tn[13].t8 VGND 0.02397f
C9570 XThR.Tn[13].n85 VGND 0.05178f
C9571 XThR.Tn[13].t11 VGND 0.02397f
C9572 XThR.Tn[13].t9 VGND 0.02397f
C9573 XThR.Tn[13].n86 VGND 0.07881f
C9574 XThR.Tn[13].n87 VGND 0.21883f
C9575 XThR.Tn[13].n88 VGND 0.0293f
C9576 XThC.XTB3.Y.t1 VGND 0.06296f
C9577 XThC.XTB3.Y.n0 VGND 0.04069f
C9578 XThC.XTB3.Y.n1 VGND 0.05192f
C9579 XThC.XTB3.Y.t2 VGND 0.03159f
C9580 XThC.XTB3.Y.t0 VGND 0.03159f
C9581 XThC.XTB3.Y.n2 VGND 0.06782f
C9582 XThC.XTB3.Y.t10 VGND 0.04914f
C9583 XThC.XTB3.Y.t17 VGND 0.02896f
C9584 XThC.XTB3.Y.n3 VGND 0.05852f
C9585 XThC.XTB3.Y.t14 VGND 0.04914f
C9586 XThC.XTB3.Y.t5 VGND 0.02896f
C9587 XThC.XTB3.Y.n4 VGND 0.03012f
C9588 XThC.XTB3.Y.t15 VGND 0.04914f
C9589 XThC.XTB3.Y.t6 VGND 0.02896f
C9590 XThC.XTB3.Y.n5 VGND 0.06469f
C9591 XThC.XTB3.Y.t3 VGND 0.04914f
C9592 XThC.XTB3.Y.t9 VGND 0.02896f
C9593 XThC.XTB3.Y.n6 VGND 0.06006f
C9594 XThC.XTB3.Y.n7 VGND 0.03654f
C9595 XThC.XTB3.Y.n8 VGND 0.06049f
C9596 XThC.XTB3.Y.n9 VGND 0.0234f
C9597 XThC.XTB3.Y.n10 VGND 0.02857f
C9598 XThC.XTB3.Y.n11 VGND 0.06469f
C9599 XThC.XTB3.Y.n12 VGND 0.03243f
C9600 XThC.XTB3.Y.n13 VGND 0.05514f
C9601 XThC.XTB3.Y.t16 VGND 0.04914f
C9602 XThC.XTB3.Y.t7 VGND 0.02896f
C9603 XThC.XTB3.Y.n14 VGND 0.06624f
C9604 XThC.XTB3.Y.t4 VGND 0.04914f
C9605 XThC.XTB3.Y.t13 VGND 0.02896f
C9606 XThC.XTB3.Y.t12 VGND 0.04914f
C9607 XThC.XTB3.Y.t18 VGND 0.02896f
C9608 XThC.XTB3.Y.t11 VGND 0.04914f
C9609 XThC.XTB3.Y.t8 VGND 0.02896f
C9610 XThC.XTB3.Y.n15 VGND 0.08245f
C9611 XThC.XTB3.Y.n16 VGND 0.08709f
C9612 XThC.XTB3.Y.n17 VGND 0.03356f
C9613 XThC.XTB3.Y.n18 VGND 0.07087f
C9614 XThC.XTB3.Y.n19 VGND 0.03243f
C9615 XThC.XTB3.Y.n20 VGND 0.02691f
C9616 XThC.XTB3.Y.n21 VGND 1.39635f
C9617 XThC.XTB3.Y.n22 VGND 0.14933f
C9618 XThR.Tn[8].t5 VGND 0.02415f
C9619 XThR.Tn[8].t3 VGND 0.02415f
C9620 XThR.Tn[8].n0 VGND 0.07334f
C9621 XThR.Tn[8].t6 VGND 0.02415f
C9622 XThR.Tn[8].t4 VGND 0.02415f
C9623 XThR.Tn[8].n1 VGND 0.05369f
C9624 XThR.Tn[8].n2 VGND 0.24415f
C9625 XThR.Tn[8].t9 VGND 0.02415f
C9626 XThR.Tn[8].t7 VGND 0.02415f
C9627 XThR.Tn[8].n3 VGND 0.05219f
C9628 XThR.Tn[8].t11 VGND 0.02415f
C9629 XThR.Tn[8].t2 VGND 0.02415f
C9630 XThR.Tn[8].n4 VGND 0.07943f
C9631 XThR.Tn[8].n5 VGND 0.22055f
C9632 XThR.Tn[8].n6 VGND 0.01087f
C9633 XThR.Tn[8].t39 VGND 0.01888f
C9634 XThR.Tn[8].t33 VGND 0.02067f
C9635 XThR.Tn[8].n7 VGND 0.05048f
C9636 XThR.Tn[8].n8 VGND 0.09697f
C9637 XThR.Tn[8].t59 VGND 0.01888f
C9638 XThR.Tn[8].t49 VGND 0.02067f
C9639 XThR.Tn[8].n9 VGND 0.05048f
C9640 XThR.Tn[8].t13 VGND 0.01882f
C9641 XThR.Tn[8].t45 VGND 0.02061f
C9642 XThR.Tn[8].n10 VGND 0.05252f
C9643 XThR.Tn[8].n11 VGND 0.0369f
C9644 XThR.Tn[8].n12 VGND 0.00675f
C9645 XThR.Tn[8].n13 VGND 0.11841f
C9646 XThR.Tn[8].t34 VGND 0.01888f
C9647 XThR.Tn[8].t26 VGND 0.02067f
C9648 XThR.Tn[8].n14 VGND 0.05048f
C9649 XThR.Tn[8].t53 VGND 0.01882f
C9650 XThR.Tn[8].t22 VGND 0.02061f
C9651 XThR.Tn[8].n15 VGND 0.05252f
C9652 XThR.Tn[8].n16 VGND 0.0369f
C9653 XThR.Tn[8].n17 VGND 0.00675f
C9654 XThR.Tn[8].n18 VGND 0.11841f
C9655 XThR.Tn[8].t50 VGND 0.01888f
C9656 XThR.Tn[8].t43 VGND 0.02067f
C9657 XThR.Tn[8].n19 VGND 0.05048f
C9658 XThR.Tn[8].t65 VGND 0.01882f
C9659 XThR.Tn[8].t40 VGND 0.02061f
C9660 XThR.Tn[8].n20 VGND 0.05252f
C9661 XThR.Tn[8].n21 VGND 0.0369f
C9662 XThR.Tn[8].n22 VGND 0.00675f
C9663 XThR.Tn[8].n23 VGND 0.11841f
C9664 XThR.Tn[8].t12 VGND 0.01888f
C9665 XThR.Tn[8].t70 VGND 0.02067f
C9666 XThR.Tn[8].n24 VGND 0.05048f
C9667 XThR.Tn[8].t36 VGND 0.01882f
C9668 XThR.Tn[8].t66 VGND 0.02061f
C9669 XThR.Tn[8].n25 VGND 0.05252f
C9670 XThR.Tn[8].n26 VGND 0.0369f
C9671 XThR.Tn[8].n27 VGND 0.00675f
C9672 XThR.Tn[8].n28 VGND 0.11841f
C9673 XThR.Tn[8].t52 VGND 0.01888f
C9674 XThR.Tn[8].t44 VGND 0.02067f
C9675 XThR.Tn[8].n29 VGND 0.05048f
C9676 XThR.Tn[8].t68 VGND 0.01882f
C9677 XThR.Tn[8].t41 VGND 0.02061f
C9678 XThR.Tn[8].n30 VGND 0.05252f
C9679 XThR.Tn[8].n31 VGND 0.0369f
C9680 XThR.Tn[8].n32 VGND 0.00675f
C9681 XThR.Tn[8].n33 VGND 0.11841f
C9682 XThR.Tn[8].t28 VGND 0.01888f
C9683 XThR.Tn[8].t61 VGND 0.02067f
C9684 XThR.Tn[8].n34 VGND 0.05048f
C9685 XThR.Tn[8].t47 VGND 0.01882f
C9686 XThR.Tn[8].t58 VGND 0.02061f
C9687 XThR.Tn[8].n35 VGND 0.05252f
C9688 XThR.Tn[8].n36 VGND 0.0369f
C9689 XThR.Tn[8].n37 VGND 0.00675f
C9690 XThR.Tn[8].n38 VGND 0.11841f
C9691 XThR.Tn[8].t60 VGND 0.01888f
C9692 XThR.Tn[8].t56 VGND 0.02067f
C9693 XThR.Tn[8].n39 VGND 0.05048f
C9694 XThR.Tn[8].t14 VGND 0.01882f
C9695 XThR.Tn[8].t51 VGND 0.02061f
C9696 XThR.Tn[8].n40 VGND 0.05252f
C9697 XThR.Tn[8].n41 VGND 0.0369f
C9698 XThR.Tn[8].n42 VGND 0.00675f
C9699 XThR.Tn[8].n43 VGND 0.11841f
C9700 XThR.Tn[8].t63 VGND 0.01888f
C9701 XThR.Tn[8].t69 VGND 0.02067f
C9702 XThR.Tn[8].n44 VGND 0.05048f
C9703 XThR.Tn[8].t20 VGND 0.01882f
C9704 XThR.Tn[8].t64 VGND 0.02061f
C9705 XThR.Tn[8].n45 VGND 0.05252f
C9706 XThR.Tn[8].n46 VGND 0.0369f
C9707 XThR.Tn[8].n47 VGND 0.00675f
C9708 XThR.Tn[8].n48 VGND 0.11841f
C9709 XThR.Tn[8].t17 VGND 0.01888f
C9710 XThR.Tn[8].t27 VGND 0.02067f
C9711 XThR.Tn[8].n49 VGND 0.05048f
C9712 XThR.Tn[8].t38 VGND 0.01882f
C9713 XThR.Tn[8].t24 VGND 0.02061f
C9714 XThR.Tn[8].n50 VGND 0.05252f
C9715 XThR.Tn[8].n51 VGND 0.0369f
C9716 XThR.Tn[8].n52 VGND 0.00675f
C9717 XThR.Tn[8].n53 VGND 0.11841f
C9718 XThR.Tn[8].t72 VGND 0.01888f
C9719 XThR.Tn[8].t46 VGND 0.02067f
C9720 XThR.Tn[8].n54 VGND 0.05048f
C9721 XThR.Tn[8].t31 VGND 0.01882f
C9722 XThR.Tn[8].t42 VGND 0.02061f
C9723 XThR.Tn[8].n55 VGND 0.05252f
C9724 XThR.Tn[8].n56 VGND 0.0369f
C9725 XThR.Tn[8].n57 VGND 0.00675f
C9726 XThR.Tn[8].n58 VGND 0.11841f
C9727 XThR.Tn[8].t30 VGND 0.01888f
C9728 XThR.Tn[8].t21 VGND 0.02067f
C9729 XThR.Tn[8].n59 VGND 0.05048f
C9730 XThR.Tn[8].t48 VGND 0.01882f
C9731 XThR.Tn[8].t16 VGND 0.02061f
C9732 XThR.Tn[8].n60 VGND 0.05252f
C9733 XThR.Tn[8].n61 VGND 0.0369f
C9734 XThR.Tn[8].n62 VGND 0.00675f
C9735 XThR.Tn[8].n63 VGND 0.11841f
C9736 XThR.Tn[8].t62 VGND 0.01888f
C9737 XThR.Tn[8].t57 VGND 0.02067f
C9738 XThR.Tn[8].n64 VGND 0.05048f
C9739 XThR.Tn[8].t18 VGND 0.01882f
C9740 XThR.Tn[8].t54 VGND 0.02061f
C9741 XThR.Tn[8].n65 VGND 0.05252f
C9742 XThR.Tn[8].n66 VGND 0.0369f
C9743 XThR.Tn[8].n67 VGND 0.00675f
C9744 XThR.Tn[8].n68 VGND 0.11841f
C9745 XThR.Tn[8].t15 VGND 0.01888f
C9746 XThR.Tn[8].t71 VGND 0.02067f
C9747 XThR.Tn[8].n69 VGND 0.05048f
C9748 XThR.Tn[8].t37 VGND 0.01882f
C9749 XThR.Tn[8].t67 VGND 0.02061f
C9750 XThR.Tn[8].n70 VGND 0.05252f
C9751 XThR.Tn[8].n71 VGND 0.0369f
C9752 XThR.Tn[8].n72 VGND 0.00675f
C9753 XThR.Tn[8].n73 VGND 0.11841f
C9754 XThR.Tn[8].t35 VGND 0.01888f
C9755 XThR.Tn[8].t29 VGND 0.02067f
C9756 XThR.Tn[8].n74 VGND 0.05048f
C9757 XThR.Tn[8].t55 VGND 0.01882f
C9758 XThR.Tn[8].t25 VGND 0.02061f
C9759 XThR.Tn[8].n75 VGND 0.05252f
C9760 XThR.Tn[8].n76 VGND 0.0369f
C9761 XThR.Tn[8].n77 VGND 0.00675f
C9762 XThR.Tn[8].n78 VGND 0.11841f
C9763 XThR.Tn[8].t73 VGND 0.01888f
C9764 XThR.Tn[8].t23 VGND 0.02067f
C9765 XThR.Tn[8].n79 VGND 0.05048f
C9766 XThR.Tn[8].t32 VGND 0.01882f
C9767 XThR.Tn[8].t19 VGND 0.02061f
C9768 XThR.Tn[8].n80 VGND 0.05252f
C9769 XThR.Tn[8].n81 VGND 0.0369f
C9770 XThR.Tn[8].n82 VGND 0.00675f
C9771 XThR.Tn[8].n83 VGND 0.11841f
C9772 XThR.Tn[8].n84 VGND 0.10761f
C9773 XThR.Tn[8].n85 VGND 0.32972f
C9774 XThR.Tn[8].t1 VGND 0.0157f
C9775 XThR.Tn[8].t10 VGND 0.0157f
C9776 XThR.Tn[8].n86 VGND 0.0314f
C9777 XThR.Tn[8].t0 VGND 0.0157f
C9778 XThR.Tn[8].t8 VGND 0.0157f
C9779 XThR.Tn[8].n87 VGND 0.03916f
C9780 XThR.Tn[8].n88 VGND 0.07241f
C9781 XThR.Tn[0].t4 VGND 0.02293f
C9782 XThR.Tn[0].t5 VGND 0.02293f
C9783 XThR.Tn[0].n0 VGND 0.04628f
C9784 XThR.Tn[0].t3 VGND 0.02293f
C9785 XThR.Tn[0].t2 VGND 0.02293f
C9786 XThR.Tn[0].n1 VGND 0.05416f
C9787 XThR.Tn[0].n2 VGND 0.16245f
C9788 XThR.Tn[0].t7 VGND 0.0149f
C9789 XThR.Tn[0].t8 VGND 0.0149f
C9790 XThR.Tn[0].n3 VGND 0.03394f
C9791 XThR.Tn[0].t6 VGND 0.0149f
C9792 XThR.Tn[0].t9 VGND 0.0149f
C9793 XThR.Tn[0].n4 VGND 0.03394f
C9794 XThR.Tn[0].t11 VGND 0.0149f
C9795 XThR.Tn[0].t10 VGND 0.0149f
C9796 XThR.Tn[0].n5 VGND 0.05655f
C9797 XThR.Tn[0].t0 VGND 0.0149f
C9798 XThR.Tn[0].t1 VGND 0.0149f
C9799 XThR.Tn[0].n6 VGND 0.03394f
C9800 XThR.Tn[0].n7 VGND 0.16164f
C9801 XThR.Tn[0].n8 VGND 0.09992f
C9802 XThR.Tn[0].n9 VGND 0.11277f
C9803 XThR.Tn[0].t48 VGND 0.01792f
C9804 XThR.Tn[0].t40 VGND 0.01962f
C9805 XThR.Tn[0].n10 VGND 0.04792f
C9806 XThR.Tn[0].n11 VGND 0.09205f
C9807 XThR.Tn[0].t67 VGND 0.01792f
C9808 XThR.Tn[0].t58 VGND 0.01962f
C9809 XThR.Tn[0].n12 VGND 0.04792f
C9810 XThR.Tn[0].t24 VGND 0.01786f
C9811 XThR.Tn[0].t50 VGND 0.01956f
C9812 XThR.Tn[0].n13 VGND 0.04986f
C9813 XThR.Tn[0].n14 VGND 0.03503f
C9814 XThR.Tn[0].n15 VGND 0.0064f
C9815 XThR.Tn[0].n16 VGND 0.11241f
C9816 XThR.Tn[0].t41 VGND 0.01792f
C9817 XThR.Tn[0].t33 VGND 0.01962f
C9818 XThR.Tn[0].n17 VGND 0.04792f
C9819 XThR.Tn[0].t61 VGND 0.01786f
C9820 XThR.Tn[0].t26 VGND 0.01956f
C9821 XThR.Tn[0].n18 VGND 0.04986f
C9822 XThR.Tn[0].n19 VGND 0.03503f
C9823 XThR.Tn[0].n20 VGND 0.0064f
C9824 XThR.Tn[0].n21 VGND 0.11241f
C9825 XThR.Tn[0].t59 VGND 0.01792f
C9826 XThR.Tn[0].t51 VGND 0.01962f
C9827 XThR.Tn[0].n22 VGND 0.04792f
C9828 XThR.Tn[0].t12 VGND 0.01786f
C9829 XThR.Tn[0].t44 VGND 0.01956f
C9830 XThR.Tn[0].n23 VGND 0.04986f
C9831 XThR.Tn[0].n24 VGND 0.03503f
C9832 XThR.Tn[0].n25 VGND 0.0064f
C9833 XThR.Tn[0].n26 VGND 0.11241f
C9834 XThR.Tn[0].t21 VGND 0.01792f
C9835 XThR.Tn[0].t15 VGND 0.01962f
C9836 XThR.Tn[0].n27 VGND 0.04792f
C9837 XThR.Tn[0].t43 VGND 0.01786f
C9838 XThR.Tn[0].t72 VGND 0.01956f
C9839 XThR.Tn[0].n28 VGND 0.04986f
C9840 XThR.Tn[0].n29 VGND 0.03503f
C9841 XThR.Tn[0].n30 VGND 0.0064f
C9842 XThR.Tn[0].n31 VGND 0.11241f
C9843 XThR.Tn[0].t60 VGND 0.01792f
C9844 XThR.Tn[0].t52 VGND 0.01962f
C9845 XThR.Tn[0].n32 VGND 0.04792f
C9846 XThR.Tn[0].t13 VGND 0.01786f
C9847 XThR.Tn[0].t46 VGND 0.01956f
C9848 XThR.Tn[0].n33 VGND 0.04986f
C9849 XThR.Tn[0].n34 VGND 0.03503f
C9850 XThR.Tn[0].n35 VGND 0.0064f
C9851 XThR.Tn[0].n36 VGND 0.11241f
C9852 XThR.Tn[0].t35 VGND 0.01792f
C9853 XThR.Tn[0].t68 VGND 0.01962f
C9854 XThR.Tn[0].n37 VGND 0.04792f
C9855 XThR.Tn[0].t54 VGND 0.01786f
C9856 XThR.Tn[0].t64 VGND 0.01956f
C9857 XThR.Tn[0].n38 VGND 0.04986f
C9858 XThR.Tn[0].n39 VGND 0.03503f
C9859 XThR.Tn[0].n40 VGND 0.0064f
C9860 XThR.Tn[0].n41 VGND 0.11241f
C9861 XThR.Tn[0].t66 VGND 0.01792f
C9862 XThR.Tn[0].t63 VGND 0.01962f
C9863 XThR.Tn[0].n42 VGND 0.04792f
C9864 XThR.Tn[0].t23 VGND 0.01786f
C9865 XThR.Tn[0].t55 VGND 0.01956f
C9866 XThR.Tn[0].n43 VGND 0.04986f
C9867 XThR.Tn[0].n44 VGND 0.03503f
C9868 XThR.Tn[0].n45 VGND 0.0064f
C9869 XThR.Tn[0].n46 VGND 0.11241f
C9870 XThR.Tn[0].t70 VGND 0.01792f
C9871 XThR.Tn[0].t14 VGND 0.01962f
C9872 XThR.Tn[0].n47 VGND 0.04792f
C9873 XThR.Tn[0].t28 VGND 0.01786f
C9874 XThR.Tn[0].t71 VGND 0.01956f
C9875 XThR.Tn[0].n48 VGND 0.04986f
C9876 XThR.Tn[0].n49 VGND 0.03503f
C9877 XThR.Tn[0].n50 VGND 0.0064f
C9878 XThR.Tn[0].n51 VGND 0.11241f
C9879 XThR.Tn[0].t25 VGND 0.01792f
C9880 XThR.Tn[0].t34 VGND 0.01962f
C9881 XThR.Tn[0].n52 VGND 0.04792f
C9882 XThR.Tn[0].t47 VGND 0.01786f
C9883 XThR.Tn[0].t29 VGND 0.01956f
C9884 XThR.Tn[0].n53 VGND 0.04986f
C9885 XThR.Tn[0].n54 VGND 0.03503f
C9886 XThR.Tn[0].n55 VGND 0.0064f
C9887 XThR.Tn[0].n56 VGND 0.11241f
C9888 XThR.Tn[0].t17 VGND 0.01792f
C9889 XThR.Tn[0].t53 VGND 0.01962f
C9890 XThR.Tn[0].n57 VGND 0.04792f
C9891 XThR.Tn[0].t38 VGND 0.01786f
C9892 XThR.Tn[0].t49 VGND 0.01956f
C9893 XThR.Tn[0].n58 VGND 0.04986f
C9894 XThR.Tn[0].n59 VGND 0.03503f
C9895 XThR.Tn[0].n60 VGND 0.0064f
C9896 XThR.Tn[0].n61 VGND 0.11241f
C9897 XThR.Tn[0].t37 VGND 0.01792f
C9898 XThR.Tn[0].t31 VGND 0.01962f
C9899 XThR.Tn[0].n62 VGND 0.04792f
C9900 XThR.Tn[0].t56 VGND 0.01786f
C9901 XThR.Tn[0].t19 VGND 0.01956f
C9902 XThR.Tn[0].n63 VGND 0.04986f
C9903 XThR.Tn[0].n64 VGND 0.03503f
C9904 XThR.Tn[0].n65 VGND 0.0064f
C9905 XThR.Tn[0].n66 VGND 0.11241f
C9906 XThR.Tn[0].t69 VGND 0.01792f
C9907 XThR.Tn[0].t65 VGND 0.01962f
C9908 XThR.Tn[0].n67 VGND 0.04792f
C9909 XThR.Tn[0].t27 VGND 0.01786f
C9910 XThR.Tn[0].t57 VGND 0.01956f
C9911 XThR.Tn[0].n68 VGND 0.04986f
C9912 XThR.Tn[0].n69 VGND 0.03503f
C9913 XThR.Tn[0].n70 VGND 0.0064f
C9914 XThR.Tn[0].n71 VGND 0.11241f
C9915 XThR.Tn[0].t22 VGND 0.01792f
C9916 XThR.Tn[0].t16 VGND 0.01962f
C9917 XThR.Tn[0].n72 VGND 0.04792f
C9918 XThR.Tn[0].t45 VGND 0.01786f
C9919 XThR.Tn[0].t73 VGND 0.01956f
C9920 XThR.Tn[0].n73 VGND 0.04986f
C9921 XThR.Tn[0].n74 VGND 0.03503f
C9922 XThR.Tn[0].n75 VGND 0.0064f
C9923 XThR.Tn[0].n76 VGND 0.11241f
C9924 XThR.Tn[0].t42 VGND 0.01792f
C9925 XThR.Tn[0].t36 VGND 0.01962f
C9926 XThR.Tn[0].n77 VGND 0.04792f
C9927 XThR.Tn[0].t62 VGND 0.01786f
C9928 XThR.Tn[0].t30 VGND 0.01956f
C9929 XThR.Tn[0].n78 VGND 0.04986f
C9930 XThR.Tn[0].n79 VGND 0.03503f
C9931 XThR.Tn[0].n80 VGND 0.0064f
C9932 XThR.Tn[0].n81 VGND 0.11241f
C9933 XThR.Tn[0].t18 VGND 0.01792f
C9934 XThR.Tn[0].t32 VGND 0.01962f
C9935 XThR.Tn[0].n82 VGND 0.04792f
C9936 XThR.Tn[0].t39 VGND 0.01786f
C9937 XThR.Tn[0].t20 VGND 0.01956f
C9938 XThR.Tn[0].n83 VGND 0.04986f
C9939 XThR.Tn[0].n84 VGND 0.03503f
C9940 XThR.Tn[0].n85 VGND 0.0064f
C9941 XThR.Tn[0].n86 VGND 0.11241f
C9942 XThR.Tn[0].n87 VGND 0.10215f
C9943 XThR.Tn[0].n88 VGND 0.29249f
C9944 XThR.Tn[7].t7 VGND 0.01503f
C9945 XThR.Tn[7].t4 VGND 0.01503f
C9946 XThR.Tn[7].n0 VGND 0.04638f
C9947 XThR.Tn[7].t6 VGND 0.01503f
C9948 XThR.Tn[7].t5 VGND 0.01503f
C9949 XThR.Tn[7].n1 VGND 0.03319f
C9950 XThR.Tn[7].n2 VGND 0.17022f
C9951 XThR.Tn[7].t2 VGND 0.02312f
C9952 XThR.Tn[7].t3 VGND 0.02312f
C9953 XThR.Tn[7].n3 VGND 0.0704f
C9954 XThR.Tn[7].t1 VGND 0.02312f
C9955 XThR.Tn[7].t0 VGND 0.02312f
C9956 XThR.Tn[7].n4 VGND 0.05122f
C9957 XThR.Tn[7].n5 VGND 0.22538f
C9958 XThR.Tn[7].n6 VGND 0.02809f
C9959 XThR.Tn[7].t53 VGND 0.01807f
C9960 XThR.Tn[7].t45 VGND 0.01979f
C9961 XThR.Tn[7].n7 VGND 0.04832f
C9962 XThR.Tn[7].n8 VGND 0.09282f
C9963 XThR.Tn[7].t8 VGND 0.01807f
C9964 XThR.Tn[7].t60 VGND 0.01979f
C9965 XThR.Tn[7].n9 VGND 0.04832f
C9966 XThR.Tn[7].t26 VGND 0.01801f
C9967 XThR.Tn[7].t38 VGND 0.01972f
C9968 XThR.Tn[7].n10 VGND 0.05027f
C9969 XThR.Tn[7].n11 VGND 0.03532f
C9970 XThR.Tn[7].n12 VGND 0.00646f
C9971 XThR.Tn[7].n13 VGND 0.11334f
C9972 XThR.Tn[7].t47 VGND 0.01807f
C9973 XThR.Tn[7].t37 VGND 0.01979f
C9974 XThR.Tn[7].n14 VGND 0.04832f
C9975 XThR.Tn[7].t66 VGND 0.01801f
C9976 XThR.Tn[7].t15 VGND 0.01972f
C9977 XThR.Tn[7].n15 VGND 0.05027f
C9978 XThR.Tn[7].n16 VGND 0.03532f
C9979 XThR.Tn[7].n17 VGND 0.00646f
C9980 XThR.Tn[7].n18 VGND 0.11334f
C9981 XThR.Tn[7].t62 VGND 0.01807f
C9982 XThR.Tn[7].t55 VGND 0.01979f
C9983 XThR.Tn[7].n19 VGND 0.04832f
C9984 XThR.Tn[7].t18 VGND 0.01801f
C9985 XThR.Tn[7].t32 VGND 0.01972f
C9986 XThR.Tn[7].n20 VGND 0.05027f
C9987 XThR.Tn[7].n21 VGND 0.03532f
C9988 XThR.Tn[7].n22 VGND 0.00646f
C9989 XThR.Tn[7].n23 VGND 0.11334f
C9990 XThR.Tn[7].t25 VGND 0.01807f
C9991 XThR.Tn[7].t21 VGND 0.01979f
C9992 XThR.Tn[7].n24 VGND 0.04832f
C9993 XThR.Tn[7].t50 VGND 0.01801f
C9994 XThR.Tn[7].t63 VGND 0.01972f
C9995 XThR.Tn[7].n25 VGND 0.05027f
C9996 XThR.Tn[7].n26 VGND 0.03532f
C9997 XThR.Tn[7].n27 VGND 0.00646f
C9998 XThR.Tn[7].n28 VGND 0.11334f
C9999 XThR.Tn[7].t65 VGND 0.01807f
C10000 XThR.Tn[7].t56 VGND 0.01979f
C10001 XThR.Tn[7].n29 VGND 0.04832f
C10002 XThR.Tn[7].t19 VGND 0.01801f
C10003 XThR.Tn[7].t34 VGND 0.01972f
C10004 XThR.Tn[7].n30 VGND 0.05027f
C10005 XThR.Tn[7].n31 VGND 0.03532f
C10006 XThR.Tn[7].n32 VGND 0.00646f
C10007 XThR.Tn[7].n33 VGND 0.11334f
C10008 XThR.Tn[7].t40 VGND 0.01807f
C10009 XThR.Tn[7].t11 VGND 0.01979f
C10010 XThR.Tn[7].n34 VGND 0.04832f
C10011 XThR.Tn[7].t58 VGND 0.01801f
C10012 XThR.Tn[7].t54 VGND 0.01972f
C10013 XThR.Tn[7].n35 VGND 0.05027f
C10014 XThR.Tn[7].n36 VGND 0.03532f
C10015 XThR.Tn[7].n37 VGND 0.00646f
C10016 XThR.Tn[7].n38 VGND 0.11334f
C10017 XThR.Tn[7].t9 VGND 0.01807f
C10018 XThR.Tn[7].t68 VGND 0.01979f
C10019 XThR.Tn[7].n39 VGND 0.04832f
C10020 XThR.Tn[7].t27 VGND 0.01801f
C10021 XThR.Tn[7].t46 VGND 0.01972f
C10022 XThR.Tn[7].n40 VGND 0.05027f
C10023 XThR.Tn[7].n41 VGND 0.03532f
C10024 XThR.Tn[7].n42 VGND 0.00646f
C10025 XThR.Tn[7].n43 VGND 0.11334f
C10026 XThR.Tn[7].t14 VGND 0.01807f
C10027 XThR.Tn[7].t20 VGND 0.01979f
C10028 XThR.Tn[7].n44 VGND 0.04832f
C10029 XThR.Tn[7].t31 VGND 0.01801f
C10030 XThR.Tn[7].t61 VGND 0.01972f
C10031 XThR.Tn[7].n45 VGND 0.05027f
C10032 XThR.Tn[7].n46 VGND 0.03532f
C10033 XThR.Tn[7].n47 VGND 0.00646f
C10034 XThR.Tn[7].n48 VGND 0.11334f
C10035 XThR.Tn[7].t29 VGND 0.01807f
C10036 XThR.Tn[7].t39 VGND 0.01979f
C10037 XThR.Tn[7].n49 VGND 0.04832f
C10038 XThR.Tn[7].t52 VGND 0.01801f
C10039 XThR.Tn[7].t16 VGND 0.01972f
C10040 XThR.Tn[7].n50 VGND 0.05027f
C10041 XThR.Tn[7].n51 VGND 0.03532f
C10042 XThR.Tn[7].n52 VGND 0.00646f
C10043 XThR.Tn[7].n53 VGND 0.11334f
C10044 XThR.Tn[7].t23 VGND 0.01807f
C10045 XThR.Tn[7].t57 VGND 0.01979f
C10046 XThR.Tn[7].n54 VGND 0.04832f
C10047 XThR.Tn[7].t43 VGND 0.01801f
C10048 XThR.Tn[7].t36 VGND 0.01972f
C10049 XThR.Tn[7].n55 VGND 0.05027f
C10050 XThR.Tn[7].n56 VGND 0.03532f
C10051 XThR.Tn[7].n57 VGND 0.00646f
C10052 XThR.Tn[7].n58 VGND 0.11334f
C10053 XThR.Tn[7].t42 VGND 0.01807f
C10054 XThR.Tn[7].t33 VGND 0.01979f
C10055 XThR.Tn[7].n59 VGND 0.04832f
C10056 XThR.Tn[7].t59 VGND 0.01801f
C10057 XThR.Tn[7].t10 VGND 0.01972f
C10058 XThR.Tn[7].n60 VGND 0.05027f
C10059 XThR.Tn[7].n61 VGND 0.03532f
C10060 XThR.Tn[7].n62 VGND 0.00646f
C10061 XThR.Tn[7].n63 VGND 0.11334f
C10062 XThR.Tn[7].t12 VGND 0.01807f
C10063 XThR.Tn[7].t69 VGND 0.01979f
C10064 XThR.Tn[7].n64 VGND 0.04832f
C10065 XThR.Tn[7].t30 VGND 0.01801f
C10066 XThR.Tn[7].t48 VGND 0.01972f
C10067 XThR.Tn[7].n65 VGND 0.05027f
C10068 XThR.Tn[7].n66 VGND 0.03532f
C10069 XThR.Tn[7].n67 VGND 0.00646f
C10070 XThR.Tn[7].n68 VGND 0.11334f
C10071 XThR.Tn[7].t28 VGND 0.01807f
C10072 XThR.Tn[7].t22 VGND 0.01979f
C10073 XThR.Tn[7].n69 VGND 0.04832f
C10074 XThR.Tn[7].t51 VGND 0.01801f
C10075 XThR.Tn[7].t64 VGND 0.01972f
C10076 XThR.Tn[7].n70 VGND 0.05027f
C10077 XThR.Tn[7].n71 VGND 0.03532f
C10078 XThR.Tn[7].n72 VGND 0.00646f
C10079 XThR.Tn[7].n73 VGND 0.11334f
C10080 XThR.Tn[7].t49 VGND 0.01807f
C10081 XThR.Tn[7].t41 VGND 0.01979f
C10082 XThR.Tn[7].n74 VGND 0.04832f
C10083 XThR.Tn[7].t67 VGND 0.01801f
C10084 XThR.Tn[7].t17 VGND 0.01972f
C10085 XThR.Tn[7].n75 VGND 0.05027f
C10086 XThR.Tn[7].n76 VGND 0.03532f
C10087 XThR.Tn[7].n77 VGND 0.00646f
C10088 XThR.Tn[7].n78 VGND 0.11334f
C10089 XThR.Tn[7].t24 VGND 0.01807f
C10090 XThR.Tn[7].t35 VGND 0.01979f
C10091 XThR.Tn[7].n79 VGND 0.04832f
C10092 XThR.Tn[7].t44 VGND 0.01801f
C10093 XThR.Tn[7].t13 VGND 0.01972f
C10094 XThR.Tn[7].n80 VGND 0.05027f
C10095 XThR.Tn[7].n81 VGND 0.03532f
C10096 XThR.Tn[7].n82 VGND 0.00646f
C10097 XThR.Tn[7].n83 VGND 0.11334f
C10098 XThR.Tn[7].n84 VGND 0.103f
C10099 XThR.Tn[7].n85 VGND 0.41812f
C10100 XThR.Tn[11].t1 VGND 0.01567f
C10101 XThR.Tn[11].t10 VGND 0.01567f
C10102 XThR.Tn[11].n0 VGND 0.03134f
C10103 XThR.Tn[11].t0 VGND 0.01567f
C10104 XThR.Tn[11].t8 VGND 0.01567f
C10105 XThR.Tn[11].n1 VGND 0.03908f
C10106 XThR.Tn[11].n2 VGND 0.07883f
C10107 XThR.Tn[11].t4 VGND 0.0241f
C10108 XThR.Tn[11].t6 VGND 0.0241f
C10109 XThR.Tn[11].n3 VGND 0.07319f
C10110 XThR.Tn[11].t5 VGND 0.0241f
C10111 XThR.Tn[11].t7 VGND 0.0241f
C10112 XThR.Tn[11].n4 VGND 0.05358f
C10113 XThR.Tn[11].n5 VGND 0.24365f
C10114 XThR.Tn[11].t11 VGND 0.0241f
C10115 XThR.Tn[11].t3 VGND 0.0241f
C10116 XThR.Tn[11].n6 VGND 0.05208f
C10117 XThR.Tn[11].t9 VGND 0.0241f
C10118 XThR.Tn[11].t2 VGND 0.0241f
C10119 XThR.Tn[11].n7 VGND 0.07927f
C10120 XThR.Tn[11].n8 VGND 0.2201f
C10121 XThR.Tn[11].n9 VGND 0.02947f
C10122 XThR.Tn[11].t56 VGND 0.01884f
C10123 XThR.Tn[11].t48 VGND 0.02063f
C10124 XThR.Tn[11].n10 VGND 0.05037f
C10125 XThR.Tn[11].n11 VGND 0.09677f
C10126 XThR.Tn[11].t12 VGND 0.01884f
C10127 XThR.Tn[11].t67 VGND 0.02063f
C10128 XThR.Tn[11].n12 VGND 0.05037f
C10129 XThR.Tn[11].t27 VGND 0.01878f
C10130 XThR.Tn[11].t58 VGND 0.02056f
C10131 XThR.Tn[11].n13 VGND 0.05241f
C10132 XThR.Tn[11].n14 VGND 0.03682f
C10133 XThR.Tn[11].n15 VGND 0.00673f
C10134 XThR.Tn[11].n16 VGND 0.11816f
C10135 XThR.Tn[11].t49 VGND 0.01884f
C10136 XThR.Tn[11].t41 VGND 0.02063f
C10137 XThR.Tn[11].n17 VGND 0.05037f
C10138 XThR.Tn[11].t65 VGND 0.01878f
C10139 XThR.Tn[11].t36 VGND 0.02056f
C10140 XThR.Tn[11].n18 VGND 0.05241f
C10141 XThR.Tn[11].n19 VGND 0.03682f
C10142 XThR.Tn[11].n20 VGND 0.00673f
C10143 XThR.Tn[11].n21 VGND 0.11816f
C10144 XThR.Tn[11].t68 VGND 0.01884f
C10145 XThR.Tn[11].t60 VGND 0.02063f
C10146 XThR.Tn[11].n22 VGND 0.05037f
C10147 XThR.Tn[11].t18 VGND 0.01878f
C10148 XThR.Tn[11].t54 VGND 0.02056f
C10149 XThR.Tn[11].n23 VGND 0.05241f
C10150 XThR.Tn[11].n24 VGND 0.03682f
C10151 XThR.Tn[11].n25 VGND 0.00673f
C10152 XThR.Tn[11].n26 VGND 0.11816f
C10153 XThR.Tn[11].t33 VGND 0.01884f
C10154 XThR.Tn[11].t23 VGND 0.02063f
C10155 XThR.Tn[11].n27 VGND 0.05037f
C10156 XThR.Tn[11].t50 VGND 0.01878f
C10157 XThR.Tn[11].t19 VGND 0.02056f
C10158 XThR.Tn[11].n28 VGND 0.05241f
C10159 XThR.Tn[11].n29 VGND 0.03682f
C10160 XThR.Tn[11].n30 VGND 0.00673f
C10161 XThR.Tn[11].n31 VGND 0.11816f
C10162 XThR.Tn[11].t70 VGND 0.01884f
C10163 XThR.Tn[11].t62 VGND 0.02063f
C10164 XThR.Tn[11].n32 VGND 0.05037f
C10165 XThR.Tn[11].t21 VGND 0.01878f
C10166 XThR.Tn[11].t55 VGND 0.02056f
C10167 XThR.Tn[11].n33 VGND 0.05241f
C10168 XThR.Tn[11].n34 VGND 0.03682f
C10169 XThR.Tn[11].n35 VGND 0.00673f
C10170 XThR.Tn[11].n36 VGND 0.11816f
C10171 XThR.Tn[11].t44 VGND 0.01884f
C10172 XThR.Tn[11].t14 VGND 0.02063f
C10173 XThR.Tn[11].n37 VGND 0.05037f
C10174 XThR.Tn[11].t59 VGND 0.01878f
C10175 XThR.Tn[11].t72 VGND 0.02056f
C10176 XThR.Tn[11].n38 VGND 0.05241f
C10177 XThR.Tn[11].n39 VGND 0.03682f
C10178 XThR.Tn[11].n40 VGND 0.00673f
C10179 XThR.Tn[11].n41 VGND 0.11816f
C10180 XThR.Tn[11].t13 VGND 0.01884f
C10181 XThR.Tn[11].t71 VGND 0.02063f
C10182 XThR.Tn[11].n42 VGND 0.05037f
C10183 XThR.Tn[11].t28 VGND 0.01878f
C10184 XThR.Tn[11].t64 VGND 0.02056f
C10185 XThR.Tn[11].n43 VGND 0.05241f
C10186 XThR.Tn[11].n44 VGND 0.03682f
C10187 XThR.Tn[11].n45 VGND 0.00673f
C10188 XThR.Tn[11].n46 VGND 0.11816f
C10189 XThR.Tn[11].t16 VGND 0.01884f
C10190 XThR.Tn[11].t22 VGND 0.02063f
C10191 XThR.Tn[11].n47 VGND 0.05037f
C10192 XThR.Tn[11].t32 VGND 0.01878f
C10193 XThR.Tn[11].t17 VGND 0.02056f
C10194 XThR.Tn[11].n48 VGND 0.05241f
C10195 XThR.Tn[11].n49 VGND 0.03682f
C10196 XThR.Tn[11].n50 VGND 0.00673f
C10197 XThR.Tn[11].n51 VGND 0.11816f
C10198 XThR.Tn[11].t35 VGND 0.01884f
C10199 XThR.Tn[11].t43 VGND 0.02063f
C10200 XThR.Tn[11].n52 VGND 0.05037f
C10201 XThR.Tn[11].t52 VGND 0.01878f
C10202 XThR.Tn[11].t37 VGND 0.02056f
C10203 XThR.Tn[11].n53 VGND 0.05241f
C10204 XThR.Tn[11].n54 VGND 0.03682f
C10205 XThR.Tn[11].n55 VGND 0.00673f
C10206 XThR.Tn[11].n56 VGND 0.11816f
C10207 XThR.Tn[11].t25 VGND 0.01884f
C10208 XThR.Tn[11].t63 VGND 0.02063f
C10209 XThR.Tn[11].n57 VGND 0.05037f
C10210 XThR.Tn[11].t42 VGND 0.01878f
C10211 XThR.Tn[11].t57 VGND 0.02056f
C10212 XThR.Tn[11].n58 VGND 0.05241f
C10213 XThR.Tn[11].n59 VGND 0.03682f
C10214 XThR.Tn[11].n60 VGND 0.00673f
C10215 XThR.Tn[11].n61 VGND 0.11816f
C10216 XThR.Tn[11].t47 VGND 0.01884f
C10217 XThR.Tn[11].t39 VGND 0.02063f
C10218 XThR.Tn[11].n62 VGND 0.05037f
C10219 XThR.Tn[11].t61 VGND 0.01878f
C10220 XThR.Tn[11].t29 VGND 0.02056f
C10221 XThR.Tn[11].n63 VGND 0.05241f
C10222 XThR.Tn[11].n64 VGND 0.03682f
C10223 XThR.Tn[11].n65 VGND 0.00673f
C10224 XThR.Tn[11].n66 VGND 0.11816f
C10225 XThR.Tn[11].t15 VGND 0.01884f
C10226 XThR.Tn[11].t73 VGND 0.02063f
C10227 XThR.Tn[11].n67 VGND 0.05037f
C10228 XThR.Tn[11].t30 VGND 0.01878f
C10229 XThR.Tn[11].t66 VGND 0.02056f
C10230 XThR.Tn[11].n68 VGND 0.05241f
C10231 XThR.Tn[11].n69 VGND 0.03682f
C10232 XThR.Tn[11].n70 VGND 0.00673f
C10233 XThR.Tn[11].n71 VGND 0.11816f
C10234 XThR.Tn[11].t34 VGND 0.01884f
C10235 XThR.Tn[11].t24 VGND 0.02063f
C10236 XThR.Tn[11].n72 VGND 0.05037f
C10237 XThR.Tn[11].t51 VGND 0.01878f
C10238 XThR.Tn[11].t20 VGND 0.02056f
C10239 XThR.Tn[11].n73 VGND 0.05241f
C10240 XThR.Tn[11].n74 VGND 0.03682f
C10241 XThR.Tn[11].n75 VGND 0.00673f
C10242 XThR.Tn[11].n76 VGND 0.11816f
C10243 XThR.Tn[11].t53 VGND 0.01884f
C10244 XThR.Tn[11].t46 VGND 0.02063f
C10245 XThR.Tn[11].n77 VGND 0.05037f
C10246 XThR.Tn[11].t69 VGND 0.01878f
C10247 XThR.Tn[11].t38 VGND 0.02056f
C10248 XThR.Tn[11].n78 VGND 0.05241f
C10249 XThR.Tn[11].n79 VGND 0.03682f
C10250 XThR.Tn[11].n80 VGND 0.00673f
C10251 XThR.Tn[11].n81 VGND 0.11816f
C10252 XThR.Tn[11].t26 VGND 0.01884f
C10253 XThR.Tn[11].t40 VGND 0.02063f
C10254 XThR.Tn[11].n82 VGND 0.05037f
C10255 XThR.Tn[11].t45 VGND 0.01878f
C10256 XThR.Tn[11].t31 VGND 0.02056f
C10257 XThR.Tn[11].n83 VGND 0.05241f
C10258 XThR.Tn[11].n84 VGND 0.03682f
C10259 XThR.Tn[11].n85 VGND 0.00673f
C10260 XThR.Tn[11].n86 VGND 0.11816f
C10261 XThR.Tn[11].n87 VGND 0.10738f
C10262 XThR.Tn[11].n88 VGND 0.38486f
C10263 XThR.Tn[4].t5 VGND 0.02325f
C10264 XThR.Tn[4].t6 VGND 0.02325f
C10265 XThR.Tn[4].n0 VGND 0.04693f
C10266 XThR.Tn[4].t4 VGND 0.02325f
C10267 XThR.Tn[4].t7 VGND 0.02325f
C10268 XThR.Tn[4].n1 VGND 0.05491f
C10269 XThR.Tn[4].n2 VGND 0.16472f
C10270 XThR.Tn[4].t8 VGND 0.01511f
C10271 XThR.Tn[4].t9 VGND 0.01511f
C10272 XThR.Tn[4].n3 VGND 0.05735f
C10273 XThR.Tn[4].t11 VGND 0.01511f
C10274 XThR.Tn[4].t10 VGND 0.01511f
C10275 XThR.Tn[4].n4 VGND 0.03442f
C10276 XThR.Tn[4].n5 VGND 0.1639f
C10277 XThR.Tn[4].t2 VGND 0.01511f
C10278 XThR.Tn[4].t1 VGND 0.01511f
C10279 XThR.Tn[4].n6 VGND 0.03442f
C10280 XThR.Tn[4].n7 VGND 0.10132f
C10281 XThR.Tn[4].t3 VGND 0.01511f
C10282 XThR.Tn[4].t0 VGND 0.01511f
C10283 XThR.Tn[4].n8 VGND 0.03442f
C10284 XThR.Tn[4].n9 VGND 0.11435f
C10285 XThR.Tn[4].t44 VGND 0.01817f
C10286 XThR.Tn[4].t38 VGND 0.0199f
C10287 XThR.Tn[4].n10 VGND 0.04859f
C10288 XThR.Tn[4].n11 VGND 0.09334f
C10289 XThR.Tn[4].t65 VGND 0.01817f
C10290 XThR.Tn[4].t54 VGND 0.0199f
C10291 XThR.Tn[4].n12 VGND 0.04859f
C10292 XThR.Tn[4].t19 VGND 0.01811f
C10293 XThR.Tn[4].t50 VGND 0.01983f
C10294 XThR.Tn[4].n13 VGND 0.05056f
C10295 XThR.Tn[4].n14 VGND 0.03552f
C10296 XThR.Tn[4].n15 VGND 0.00649f
C10297 XThR.Tn[4].n16 VGND 0.11398f
C10298 XThR.Tn[4].t39 VGND 0.01817f
C10299 XThR.Tn[4].t31 VGND 0.0199f
C10300 XThR.Tn[4].n17 VGND 0.04859f
C10301 XThR.Tn[4].t58 VGND 0.01811f
C10302 XThR.Tn[4].t27 VGND 0.01983f
C10303 XThR.Tn[4].n18 VGND 0.05056f
C10304 XThR.Tn[4].n19 VGND 0.03552f
C10305 XThR.Tn[4].n20 VGND 0.00649f
C10306 XThR.Tn[4].n21 VGND 0.11398f
C10307 XThR.Tn[4].t55 VGND 0.01817f
C10308 XThR.Tn[4].t48 VGND 0.0199f
C10309 XThR.Tn[4].n22 VGND 0.04859f
C10310 XThR.Tn[4].t70 VGND 0.01811f
C10311 XThR.Tn[4].t45 VGND 0.01983f
C10312 XThR.Tn[4].n23 VGND 0.05056f
C10313 XThR.Tn[4].n24 VGND 0.03552f
C10314 XThR.Tn[4].n25 VGND 0.00649f
C10315 XThR.Tn[4].n26 VGND 0.11398f
C10316 XThR.Tn[4].t17 VGND 0.01817f
C10317 XThR.Tn[4].t13 VGND 0.0199f
C10318 XThR.Tn[4].n27 VGND 0.04859f
C10319 XThR.Tn[4].t41 VGND 0.01811f
C10320 XThR.Tn[4].t71 VGND 0.01983f
C10321 XThR.Tn[4].n28 VGND 0.05056f
C10322 XThR.Tn[4].n29 VGND 0.03552f
C10323 XThR.Tn[4].n30 VGND 0.00649f
C10324 XThR.Tn[4].n31 VGND 0.11398f
C10325 XThR.Tn[4].t57 VGND 0.01817f
C10326 XThR.Tn[4].t49 VGND 0.0199f
C10327 XThR.Tn[4].n32 VGND 0.04859f
C10328 XThR.Tn[4].t73 VGND 0.01811f
C10329 XThR.Tn[4].t46 VGND 0.01983f
C10330 XThR.Tn[4].n33 VGND 0.05056f
C10331 XThR.Tn[4].n34 VGND 0.03552f
C10332 XThR.Tn[4].n35 VGND 0.00649f
C10333 XThR.Tn[4].n36 VGND 0.11398f
C10334 XThR.Tn[4].t33 VGND 0.01817f
C10335 XThR.Tn[4].t66 VGND 0.0199f
C10336 XThR.Tn[4].n37 VGND 0.04859f
C10337 XThR.Tn[4].t52 VGND 0.01811f
C10338 XThR.Tn[4].t63 VGND 0.01983f
C10339 XThR.Tn[4].n38 VGND 0.05056f
C10340 XThR.Tn[4].n39 VGND 0.03552f
C10341 XThR.Tn[4].n40 VGND 0.00649f
C10342 XThR.Tn[4].n41 VGND 0.11398f
C10343 XThR.Tn[4].t64 VGND 0.01817f
C10344 XThR.Tn[4].t61 VGND 0.0199f
C10345 XThR.Tn[4].n42 VGND 0.04859f
C10346 XThR.Tn[4].t18 VGND 0.01811f
C10347 XThR.Tn[4].t56 VGND 0.01983f
C10348 XThR.Tn[4].n43 VGND 0.05056f
C10349 XThR.Tn[4].n44 VGND 0.03552f
C10350 XThR.Tn[4].n45 VGND 0.00649f
C10351 XThR.Tn[4].n46 VGND 0.11398f
C10352 XThR.Tn[4].t68 VGND 0.01817f
C10353 XThR.Tn[4].t12 VGND 0.0199f
C10354 XThR.Tn[4].n47 VGND 0.04859f
C10355 XThR.Tn[4].t25 VGND 0.01811f
C10356 XThR.Tn[4].t69 VGND 0.01983f
C10357 XThR.Tn[4].n48 VGND 0.05056f
C10358 XThR.Tn[4].n49 VGND 0.03552f
C10359 XThR.Tn[4].n50 VGND 0.00649f
C10360 XThR.Tn[4].n51 VGND 0.11398f
C10361 XThR.Tn[4].t22 VGND 0.01817f
C10362 XThR.Tn[4].t32 VGND 0.0199f
C10363 XThR.Tn[4].n52 VGND 0.04859f
C10364 XThR.Tn[4].t43 VGND 0.01811f
C10365 XThR.Tn[4].t29 VGND 0.01983f
C10366 XThR.Tn[4].n53 VGND 0.05056f
C10367 XThR.Tn[4].n54 VGND 0.03552f
C10368 XThR.Tn[4].n55 VGND 0.00649f
C10369 XThR.Tn[4].n56 VGND 0.11398f
C10370 XThR.Tn[4].t15 VGND 0.01817f
C10371 XThR.Tn[4].t51 VGND 0.0199f
C10372 XThR.Tn[4].n57 VGND 0.04859f
C10373 XThR.Tn[4].t36 VGND 0.01811f
C10374 XThR.Tn[4].t47 VGND 0.01983f
C10375 XThR.Tn[4].n58 VGND 0.05056f
C10376 XThR.Tn[4].n59 VGND 0.03552f
C10377 XThR.Tn[4].n60 VGND 0.00649f
C10378 XThR.Tn[4].n61 VGND 0.11398f
C10379 XThR.Tn[4].t35 VGND 0.01817f
C10380 XThR.Tn[4].t26 VGND 0.0199f
C10381 XThR.Tn[4].n62 VGND 0.04859f
C10382 XThR.Tn[4].t53 VGND 0.01811f
C10383 XThR.Tn[4].t21 VGND 0.01983f
C10384 XThR.Tn[4].n63 VGND 0.05056f
C10385 XThR.Tn[4].n64 VGND 0.03552f
C10386 XThR.Tn[4].n65 VGND 0.00649f
C10387 XThR.Tn[4].n66 VGND 0.11398f
C10388 XThR.Tn[4].t67 VGND 0.01817f
C10389 XThR.Tn[4].t62 VGND 0.0199f
C10390 XThR.Tn[4].n67 VGND 0.04859f
C10391 XThR.Tn[4].t23 VGND 0.01811f
C10392 XThR.Tn[4].t59 VGND 0.01983f
C10393 XThR.Tn[4].n68 VGND 0.05056f
C10394 XThR.Tn[4].n69 VGND 0.03552f
C10395 XThR.Tn[4].n70 VGND 0.00649f
C10396 XThR.Tn[4].n71 VGND 0.11398f
C10397 XThR.Tn[4].t20 VGND 0.01817f
C10398 XThR.Tn[4].t14 VGND 0.0199f
C10399 XThR.Tn[4].n72 VGND 0.04859f
C10400 XThR.Tn[4].t42 VGND 0.01811f
C10401 XThR.Tn[4].t72 VGND 0.01983f
C10402 XThR.Tn[4].n73 VGND 0.05056f
C10403 XThR.Tn[4].n74 VGND 0.03552f
C10404 XThR.Tn[4].n75 VGND 0.00649f
C10405 XThR.Tn[4].n76 VGND 0.11398f
C10406 XThR.Tn[4].t40 VGND 0.01817f
C10407 XThR.Tn[4].t34 VGND 0.0199f
C10408 XThR.Tn[4].n77 VGND 0.04859f
C10409 XThR.Tn[4].t60 VGND 0.01811f
C10410 XThR.Tn[4].t30 VGND 0.01983f
C10411 XThR.Tn[4].n78 VGND 0.05056f
C10412 XThR.Tn[4].n79 VGND 0.03552f
C10413 XThR.Tn[4].n80 VGND 0.00649f
C10414 XThR.Tn[4].n81 VGND 0.11398f
C10415 XThR.Tn[4].t16 VGND 0.01817f
C10416 XThR.Tn[4].t28 VGND 0.0199f
C10417 XThR.Tn[4].n82 VGND 0.04859f
C10418 XThR.Tn[4].t37 VGND 0.01811f
C10419 XThR.Tn[4].t24 VGND 0.01983f
C10420 XThR.Tn[4].n83 VGND 0.05056f
C10421 XThR.Tn[4].n84 VGND 0.03552f
C10422 XThR.Tn[4].n85 VGND 0.00649f
C10423 XThR.Tn[4].n86 VGND 0.11398f
C10424 XThR.Tn[4].n87 VGND 0.10358f
C10425 XThR.Tn[4].n88 VGND 0.19569f
C10426 XThC.Tn[7].t6 VGND 0.01228f
C10427 XThC.Tn[7].t5 VGND 0.01228f
C10428 XThC.Tn[7].n0 VGND 0.03791f
C10429 XThC.Tn[7].t4 VGND 0.01228f
C10430 XThC.Tn[7].t7 VGND 0.01228f
C10431 XThC.Tn[7].n1 VGND 0.02713f
C10432 XThC.Tn[7].n2 VGND 0.13418f
C10433 XThC.Tn[7].t0 VGND 0.0189f
C10434 XThC.Tn[7].t3 VGND 0.0189f
C10435 XThC.Tn[7].n3 VGND 0.0407f
C10436 XThC.Tn[7].t2 VGND 0.0189f
C10437 XThC.Tn[7].t1 VGND 0.0189f
C10438 XThC.Tn[7].n4 VGND 0.06179f
C10439 XThC.Tn[7].n5 VGND 0.18167f
C10440 XThC.Tn[7].t8 VGND 0.01498f
C10441 XThC.Tn[7].t11 VGND 0.01636f
C10442 XThC.Tn[7].n6 VGND 0.03652f
C10443 XThC.Tn[7].n7 VGND 0.02502f
C10444 XThC.Tn[7].n8 VGND 0.08213f
C10445 XThC.Tn[7].t25 VGND 0.01498f
C10446 XThC.Tn[7].t30 VGND 0.01636f
C10447 XThC.Tn[7].n9 VGND 0.03652f
C10448 XThC.Tn[7].n10 VGND 0.02502f
C10449 XThC.Tn[7].n11 VGND 0.08235f
C10450 XThC.Tn[7].n12 VGND 0.13573f
C10451 XThC.Tn[7].t27 VGND 0.01498f
C10452 XThC.Tn[7].t34 VGND 0.01636f
C10453 XThC.Tn[7].n13 VGND 0.03652f
C10454 XThC.Tn[7].n14 VGND 0.02502f
C10455 XThC.Tn[7].n15 VGND 0.08235f
C10456 XThC.Tn[7].n16 VGND 0.13573f
C10457 XThC.Tn[7].t29 VGND 0.01498f
C10458 XThC.Tn[7].t35 VGND 0.01636f
C10459 XThC.Tn[7].n17 VGND 0.03652f
C10460 XThC.Tn[7].n18 VGND 0.02502f
C10461 XThC.Tn[7].n19 VGND 0.08235f
C10462 XThC.Tn[7].n20 VGND 0.13573f
C10463 XThC.Tn[7].t18 VGND 0.01498f
C10464 XThC.Tn[7].t22 VGND 0.01636f
C10465 XThC.Tn[7].n21 VGND 0.03652f
C10466 XThC.Tn[7].n22 VGND 0.02502f
C10467 XThC.Tn[7].n23 VGND 0.08235f
C10468 XThC.Tn[7].n24 VGND 0.13573f
C10469 XThC.Tn[7].t20 VGND 0.01498f
C10470 XThC.Tn[7].t23 VGND 0.01636f
C10471 XThC.Tn[7].n25 VGND 0.03652f
C10472 XThC.Tn[7].n26 VGND 0.02502f
C10473 XThC.Tn[7].n27 VGND 0.08235f
C10474 XThC.Tn[7].n28 VGND 0.13573f
C10475 XThC.Tn[7].t33 VGND 0.01498f
C10476 XThC.Tn[7].t39 VGND 0.01636f
C10477 XThC.Tn[7].n29 VGND 0.03652f
C10478 XThC.Tn[7].n30 VGND 0.02502f
C10479 XThC.Tn[7].n31 VGND 0.08235f
C10480 XThC.Tn[7].n32 VGND 0.13573f
C10481 XThC.Tn[7].t10 VGND 0.01498f
C10482 XThC.Tn[7].t14 VGND 0.01636f
C10483 XThC.Tn[7].n33 VGND 0.03652f
C10484 XThC.Tn[7].n34 VGND 0.02502f
C10485 XThC.Tn[7].n35 VGND 0.08235f
C10486 XThC.Tn[7].n36 VGND 0.13573f
C10487 XThC.Tn[7].t12 VGND 0.01498f
C10488 XThC.Tn[7].t16 VGND 0.01636f
C10489 XThC.Tn[7].n37 VGND 0.03652f
C10490 XThC.Tn[7].n38 VGND 0.02502f
C10491 XThC.Tn[7].n39 VGND 0.08235f
C10492 XThC.Tn[7].n40 VGND 0.13573f
C10493 XThC.Tn[7].t31 VGND 0.01498f
C10494 XThC.Tn[7].t36 VGND 0.01636f
C10495 XThC.Tn[7].n41 VGND 0.03652f
C10496 XThC.Tn[7].n42 VGND 0.02502f
C10497 XThC.Tn[7].n43 VGND 0.08235f
C10498 XThC.Tn[7].n44 VGND 0.13573f
C10499 XThC.Tn[7].t32 VGND 0.01498f
C10500 XThC.Tn[7].t38 VGND 0.01636f
C10501 XThC.Tn[7].n45 VGND 0.03652f
C10502 XThC.Tn[7].n46 VGND 0.02502f
C10503 XThC.Tn[7].n47 VGND 0.08235f
C10504 XThC.Tn[7].n48 VGND 0.13573f
C10505 XThC.Tn[7].t13 VGND 0.01498f
C10506 XThC.Tn[7].t17 VGND 0.01636f
C10507 XThC.Tn[7].n49 VGND 0.03652f
C10508 XThC.Tn[7].n50 VGND 0.02502f
C10509 XThC.Tn[7].n51 VGND 0.08235f
C10510 XThC.Tn[7].n52 VGND 0.13573f
C10511 XThC.Tn[7].t21 VGND 0.01498f
C10512 XThC.Tn[7].t26 VGND 0.01636f
C10513 XThC.Tn[7].n53 VGND 0.03652f
C10514 XThC.Tn[7].n54 VGND 0.02502f
C10515 XThC.Tn[7].n55 VGND 0.08235f
C10516 XThC.Tn[7].n56 VGND 0.13573f
C10517 XThC.Tn[7].t24 VGND 0.01498f
C10518 XThC.Tn[7].t28 VGND 0.01636f
C10519 XThC.Tn[7].n57 VGND 0.03652f
C10520 XThC.Tn[7].n58 VGND 0.02502f
C10521 XThC.Tn[7].n59 VGND 0.08235f
C10522 XThC.Tn[7].n60 VGND 0.13573f
C10523 XThC.Tn[7].t37 VGND 0.01498f
C10524 XThC.Tn[7].t9 VGND 0.01636f
C10525 XThC.Tn[7].n61 VGND 0.03652f
C10526 XThC.Tn[7].n62 VGND 0.02502f
C10527 XThC.Tn[7].n63 VGND 0.08235f
C10528 XThC.Tn[7].n64 VGND 0.13573f
C10529 XThC.Tn[7].t15 VGND 0.01498f
C10530 XThC.Tn[7].t19 VGND 0.01636f
C10531 XThC.Tn[7].n65 VGND 0.03652f
C10532 XThC.Tn[7].n66 VGND 0.02502f
C10533 XThC.Tn[7].n67 VGND 0.08235f
C10534 XThC.Tn[7].n68 VGND 0.13573f
C10535 XThC.Tn[7].n69 VGND 0.34086f
C10536 XThC.Tn[7].n70 VGND 0.02261f
C10537 XThR.Tn[1].t4 VGND 0.02304f
C10538 XThR.Tn[1].t5 VGND 0.02304f
C10539 XThR.Tn[1].n0 VGND 0.0465f
C10540 XThR.Tn[1].t7 VGND 0.02304f
C10541 XThR.Tn[1].t6 VGND 0.02304f
C10542 XThR.Tn[1].n1 VGND 0.05441f
C10543 XThR.Tn[1].n2 VGND 0.15232f
C10544 XThR.Tn[1].t11 VGND 0.01497f
C10545 XThR.Tn[1].t8 VGND 0.01497f
C10546 XThR.Tn[1].n3 VGND 0.05682f
C10547 XThR.Tn[1].t10 VGND 0.01497f
C10548 XThR.Tn[1].t9 VGND 0.01497f
C10549 XThR.Tn[1].n4 VGND 0.0341f
C10550 XThR.Tn[1].n5 VGND 0.16239f
C10551 XThR.Tn[1].t2 VGND 0.01497f
C10552 XThR.Tn[1].t1 VGND 0.01497f
C10553 XThR.Tn[1].n6 VGND 0.0341f
C10554 XThR.Tn[1].n7 VGND 0.10039f
C10555 XThR.Tn[1].t3 VGND 0.01497f
C10556 XThR.Tn[1].t0 VGND 0.01497f
C10557 XThR.Tn[1].n8 VGND 0.0341f
C10558 XThR.Tn[1].n9 VGND 0.11329f
C10559 XThR.Tn[1].t24 VGND 0.01801f
C10560 XThR.Tn[1].t18 VGND 0.01972f
C10561 XThR.Tn[1].n10 VGND 0.04814f
C10562 XThR.Tn[1].n11 VGND 0.09248f
C10563 XThR.Tn[1].t44 VGND 0.01801f
C10564 XThR.Tn[1].t34 VGND 0.01972f
C10565 XThR.Tn[1].n12 VGND 0.04814f
C10566 XThR.Tn[1].t61 VGND 0.01795f
C10567 XThR.Tn[1].t30 VGND 0.01965f
C10568 XThR.Tn[1].n13 VGND 0.05009f
C10569 XThR.Tn[1].n14 VGND 0.03519f
C10570 XThR.Tn[1].n15 VGND 0.00643f
C10571 XThR.Tn[1].n16 VGND 0.11293f
C10572 XThR.Tn[1].t19 VGND 0.01801f
C10573 XThR.Tn[1].t73 VGND 0.01972f
C10574 XThR.Tn[1].n17 VGND 0.04814f
C10575 XThR.Tn[1].t38 VGND 0.01795f
C10576 XThR.Tn[1].t69 VGND 0.01965f
C10577 XThR.Tn[1].n18 VGND 0.05009f
C10578 XThR.Tn[1].n19 VGND 0.03519f
C10579 XThR.Tn[1].n20 VGND 0.00643f
C10580 XThR.Tn[1].n21 VGND 0.11293f
C10581 XThR.Tn[1].t35 VGND 0.01801f
C10582 XThR.Tn[1].t28 VGND 0.01972f
C10583 XThR.Tn[1].n22 VGND 0.04814f
C10584 XThR.Tn[1].t50 VGND 0.01795f
C10585 XThR.Tn[1].t25 VGND 0.01965f
C10586 XThR.Tn[1].n23 VGND 0.05009f
C10587 XThR.Tn[1].n24 VGND 0.03519f
C10588 XThR.Tn[1].n25 VGND 0.00643f
C10589 XThR.Tn[1].n26 VGND 0.11293f
C10590 XThR.Tn[1].t59 VGND 0.01801f
C10591 XThR.Tn[1].t55 VGND 0.01972f
C10592 XThR.Tn[1].n27 VGND 0.04814f
C10593 XThR.Tn[1].t21 VGND 0.01795f
C10594 XThR.Tn[1].t51 VGND 0.01965f
C10595 XThR.Tn[1].n28 VGND 0.05009f
C10596 XThR.Tn[1].n29 VGND 0.03519f
C10597 XThR.Tn[1].n30 VGND 0.00643f
C10598 XThR.Tn[1].n31 VGND 0.11293f
C10599 XThR.Tn[1].t37 VGND 0.01801f
C10600 XThR.Tn[1].t29 VGND 0.01972f
C10601 XThR.Tn[1].n32 VGND 0.04814f
C10602 XThR.Tn[1].t53 VGND 0.01795f
C10603 XThR.Tn[1].t26 VGND 0.01965f
C10604 XThR.Tn[1].n33 VGND 0.05009f
C10605 XThR.Tn[1].n34 VGND 0.03519f
C10606 XThR.Tn[1].n35 VGND 0.00643f
C10607 XThR.Tn[1].n36 VGND 0.11293f
C10608 XThR.Tn[1].t13 VGND 0.01801f
C10609 XThR.Tn[1].t46 VGND 0.01972f
C10610 XThR.Tn[1].n37 VGND 0.04814f
C10611 XThR.Tn[1].t32 VGND 0.01795f
C10612 XThR.Tn[1].t43 VGND 0.01965f
C10613 XThR.Tn[1].n38 VGND 0.05009f
C10614 XThR.Tn[1].n39 VGND 0.03519f
C10615 XThR.Tn[1].n40 VGND 0.00643f
C10616 XThR.Tn[1].n41 VGND 0.11293f
C10617 XThR.Tn[1].t45 VGND 0.01801f
C10618 XThR.Tn[1].t41 VGND 0.01972f
C10619 XThR.Tn[1].n42 VGND 0.04814f
C10620 XThR.Tn[1].t60 VGND 0.01795f
C10621 XThR.Tn[1].t36 VGND 0.01965f
C10622 XThR.Tn[1].n43 VGND 0.05009f
C10623 XThR.Tn[1].n44 VGND 0.03519f
C10624 XThR.Tn[1].n45 VGND 0.00643f
C10625 XThR.Tn[1].n46 VGND 0.11293f
C10626 XThR.Tn[1].t48 VGND 0.01801f
C10627 XThR.Tn[1].t54 VGND 0.01972f
C10628 XThR.Tn[1].n47 VGND 0.04814f
C10629 XThR.Tn[1].t67 VGND 0.01795f
C10630 XThR.Tn[1].t49 VGND 0.01965f
C10631 XThR.Tn[1].n48 VGND 0.05009f
C10632 XThR.Tn[1].n49 VGND 0.03519f
C10633 XThR.Tn[1].n50 VGND 0.00643f
C10634 XThR.Tn[1].n51 VGND 0.11293f
C10635 XThR.Tn[1].t64 VGND 0.01801f
C10636 XThR.Tn[1].t12 VGND 0.01972f
C10637 XThR.Tn[1].n52 VGND 0.04814f
C10638 XThR.Tn[1].t23 VGND 0.01795f
C10639 XThR.Tn[1].t71 VGND 0.01965f
C10640 XThR.Tn[1].n53 VGND 0.05009f
C10641 XThR.Tn[1].n54 VGND 0.03519f
C10642 XThR.Tn[1].n55 VGND 0.00643f
C10643 XThR.Tn[1].n56 VGND 0.11293f
C10644 XThR.Tn[1].t57 VGND 0.01801f
C10645 XThR.Tn[1].t31 VGND 0.01972f
C10646 XThR.Tn[1].n57 VGND 0.04814f
C10647 XThR.Tn[1].t16 VGND 0.01795f
C10648 XThR.Tn[1].t27 VGND 0.01965f
C10649 XThR.Tn[1].n58 VGND 0.05009f
C10650 XThR.Tn[1].n59 VGND 0.03519f
C10651 XThR.Tn[1].n60 VGND 0.00643f
C10652 XThR.Tn[1].n61 VGND 0.11293f
C10653 XThR.Tn[1].t15 VGND 0.01801f
C10654 XThR.Tn[1].t68 VGND 0.01972f
C10655 XThR.Tn[1].n62 VGND 0.04814f
C10656 XThR.Tn[1].t33 VGND 0.01795f
C10657 XThR.Tn[1].t63 VGND 0.01965f
C10658 XThR.Tn[1].n63 VGND 0.05009f
C10659 XThR.Tn[1].n64 VGND 0.03519f
C10660 XThR.Tn[1].n65 VGND 0.00643f
C10661 XThR.Tn[1].n66 VGND 0.11293f
C10662 XThR.Tn[1].t47 VGND 0.01801f
C10663 XThR.Tn[1].t42 VGND 0.01972f
C10664 XThR.Tn[1].n67 VGND 0.04814f
C10665 XThR.Tn[1].t65 VGND 0.01795f
C10666 XThR.Tn[1].t39 VGND 0.01965f
C10667 XThR.Tn[1].n68 VGND 0.05009f
C10668 XThR.Tn[1].n69 VGND 0.03519f
C10669 XThR.Tn[1].n70 VGND 0.00643f
C10670 XThR.Tn[1].n71 VGND 0.11293f
C10671 XThR.Tn[1].t62 VGND 0.01801f
C10672 XThR.Tn[1].t56 VGND 0.01972f
C10673 XThR.Tn[1].n72 VGND 0.04814f
C10674 XThR.Tn[1].t22 VGND 0.01795f
C10675 XThR.Tn[1].t52 VGND 0.01965f
C10676 XThR.Tn[1].n73 VGND 0.05009f
C10677 XThR.Tn[1].n74 VGND 0.03519f
C10678 XThR.Tn[1].n75 VGND 0.00643f
C10679 XThR.Tn[1].n76 VGND 0.11293f
C10680 XThR.Tn[1].t20 VGND 0.01801f
C10681 XThR.Tn[1].t14 VGND 0.01972f
C10682 XThR.Tn[1].n77 VGND 0.04814f
C10683 XThR.Tn[1].t40 VGND 0.01795f
C10684 XThR.Tn[1].t72 VGND 0.01965f
C10685 XThR.Tn[1].n78 VGND 0.05009f
C10686 XThR.Tn[1].n79 VGND 0.03519f
C10687 XThR.Tn[1].n80 VGND 0.00643f
C10688 XThR.Tn[1].n81 VGND 0.11293f
C10689 XThR.Tn[1].t58 VGND 0.01801f
C10690 XThR.Tn[1].t70 VGND 0.01972f
C10691 XThR.Tn[1].n82 VGND 0.04814f
C10692 XThR.Tn[1].t17 VGND 0.01795f
C10693 XThR.Tn[1].t66 VGND 0.01965f
C10694 XThR.Tn[1].n83 VGND 0.05009f
C10695 XThR.Tn[1].n84 VGND 0.03519f
C10696 XThR.Tn[1].n85 VGND 0.00643f
C10697 XThR.Tn[1].n86 VGND 0.11293f
C10698 XThR.Tn[1].n87 VGND 0.10263f
C10699 XThR.Tn[1].n88 VGND 0.29541f
C10700 XThR.Tn[1].n89 VGND 0.04821f
C10701 XThC.Tn[8].t5 VGND 0.01304f
C10702 XThC.Tn[8].t4 VGND 0.01304f
C10703 XThC.Tn[8].n0 VGND 0.03253f
C10704 XThC.Tn[8].t7 VGND 0.01304f
C10705 XThC.Tn[8].t6 VGND 0.01304f
C10706 XThC.Tn[8].n1 VGND 0.02608f
C10707 XThC.Tn[8].n2 VGND 0.06561f
C10708 XThC.Tn[8].n3 VGND 0.02453f
C10709 XThC.Tn[8].t43 VGND 0.0159f
C10710 XThC.Tn[8].t41 VGND 0.01737f
C10711 XThC.Tn[8].n4 VGND 0.03878f
C10712 XThC.Tn[8].n5 VGND 0.02657f
C10713 XThC.Tn[8].n6 VGND 0.0872f
C10714 XThC.Tn[8].t29 VGND 0.0159f
C10715 XThC.Tn[8].t26 VGND 0.01737f
C10716 XThC.Tn[8].n7 VGND 0.03878f
C10717 XThC.Tn[8].n8 VGND 0.02657f
C10718 XThC.Tn[8].n9 VGND 0.08744f
C10719 XThC.Tn[8].n10 VGND 0.1441f
C10720 XThC.Tn[8].t34 VGND 0.0159f
C10721 XThC.Tn[8].t28 VGND 0.01737f
C10722 XThC.Tn[8].n11 VGND 0.03878f
C10723 XThC.Tn[8].n12 VGND 0.02657f
C10724 XThC.Tn[8].n13 VGND 0.08744f
C10725 XThC.Tn[8].n14 VGND 0.1441f
C10726 XThC.Tn[8].t35 VGND 0.0159f
C10727 XThC.Tn[8].t30 VGND 0.01737f
C10728 XThC.Tn[8].n15 VGND 0.03878f
C10729 XThC.Tn[8].n16 VGND 0.02657f
C10730 XThC.Tn[8].n17 VGND 0.08744f
C10731 XThC.Tn[8].n18 VGND 0.1441f
C10732 XThC.Tn[8].t22 VGND 0.0159f
C10733 XThC.Tn[8].t19 VGND 0.01737f
C10734 XThC.Tn[8].n19 VGND 0.03878f
C10735 XThC.Tn[8].n20 VGND 0.02657f
C10736 XThC.Tn[8].n21 VGND 0.08744f
C10737 XThC.Tn[8].n22 VGND 0.1441f
C10738 XThC.Tn[8].t23 VGND 0.0159f
C10739 XThC.Tn[8].t20 VGND 0.01737f
C10740 XThC.Tn[8].n23 VGND 0.03878f
C10741 XThC.Tn[8].n24 VGND 0.02657f
C10742 XThC.Tn[8].n25 VGND 0.08744f
C10743 XThC.Tn[8].n26 VGND 0.1441f
C10744 XThC.Tn[8].t39 VGND 0.0159f
C10745 XThC.Tn[8].t33 VGND 0.01737f
C10746 XThC.Tn[8].n27 VGND 0.03878f
C10747 XThC.Tn[8].n28 VGND 0.02657f
C10748 XThC.Tn[8].n29 VGND 0.08744f
C10749 XThC.Tn[8].n30 VGND 0.1441f
C10750 XThC.Tn[8].t14 VGND 0.0159f
C10751 XThC.Tn[8].t42 VGND 0.01737f
C10752 XThC.Tn[8].n31 VGND 0.03878f
C10753 XThC.Tn[8].n32 VGND 0.02657f
C10754 XThC.Tn[8].n33 VGND 0.08744f
C10755 XThC.Tn[8].n34 VGND 0.1441f
C10756 XThC.Tn[8].t16 VGND 0.0159f
C10757 XThC.Tn[8].t12 VGND 0.01737f
C10758 XThC.Tn[8].n35 VGND 0.03878f
C10759 XThC.Tn[8].n36 VGND 0.02657f
C10760 XThC.Tn[8].n37 VGND 0.08744f
C10761 XThC.Tn[8].n38 VGND 0.1441f
C10762 XThC.Tn[8].t36 VGND 0.0159f
C10763 XThC.Tn[8].t31 VGND 0.01737f
C10764 XThC.Tn[8].n39 VGND 0.03878f
C10765 XThC.Tn[8].n40 VGND 0.02657f
C10766 XThC.Tn[8].n41 VGND 0.08744f
C10767 XThC.Tn[8].n42 VGND 0.1441f
C10768 XThC.Tn[8].t38 VGND 0.0159f
C10769 XThC.Tn[8].t32 VGND 0.01737f
C10770 XThC.Tn[8].n43 VGND 0.03878f
C10771 XThC.Tn[8].n44 VGND 0.02657f
C10772 XThC.Tn[8].n45 VGND 0.08744f
C10773 XThC.Tn[8].n46 VGND 0.1441f
C10774 XThC.Tn[8].t17 VGND 0.0159f
C10775 XThC.Tn[8].t13 VGND 0.01737f
C10776 XThC.Tn[8].n47 VGND 0.03878f
C10777 XThC.Tn[8].n48 VGND 0.02657f
C10778 XThC.Tn[8].n49 VGND 0.08744f
C10779 XThC.Tn[8].n50 VGND 0.1441f
C10780 XThC.Tn[8].t25 VGND 0.0159f
C10781 XThC.Tn[8].t21 VGND 0.01737f
C10782 XThC.Tn[8].n51 VGND 0.03878f
C10783 XThC.Tn[8].n52 VGND 0.02657f
C10784 XThC.Tn[8].n53 VGND 0.08744f
C10785 XThC.Tn[8].n54 VGND 0.1441f
C10786 XThC.Tn[8].t27 VGND 0.0159f
C10787 XThC.Tn[8].t24 VGND 0.01737f
C10788 XThC.Tn[8].n55 VGND 0.03878f
C10789 XThC.Tn[8].n56 VGND 0.02657f
C10790 XThC.Tn[8].n57 VGND 0.08744f
C10791 XThC.Tn[8].n58 VGND 0.1441f
C10792 XThC.Tn[8].t40 VGND 0.0159f
C10793 XThC.Tn[8].t37 VGND 0.01737f
C10794 XThC.Tn[8].n59 VGND 0.03878f
C10795 XThC.Tn[8].n60 VGND 0.02657f
C10796 XThC.Tn[8].n61 VGND 0.08744f
C10797 XThC.Tn[8].n62 VGND 0.1441f
C10798 XThC.Tn[8].t18 VGND 0.0159f
C10799 XThC.Tn[8].t15 VGND 0.01737f
C10800 XThC.Tn[8].n63 VGND 0.03878f
C10801 XThC.Tn[8].n64 VGND 0.02657f
C10802 XThC.Tn[8].n65 VGND 0.08744f
C10803 XThC.Tn[8].n66 VGND 0.1441f
C10804 XThC.Tn[8].n67 VGND 0.60346f
C10805 XThC.Tn[8].n68 VGND 0.23618f
C10806 XThC.Tn[8].t9 VGND 0.02006f
C10807 XThC.Tn[8].t10 VGND 0.02006f
C10808 XThC.Tn[8].n69 VGND 0.04335f
C10809 XThC.Tn[8].t8 VGND 0.02006f
C10810 XThC.Tn[8].t11 VGND 0.02006f
C10811 XThC.Tn[8].n70 VGND 0.06598f
C10812 XThC.Tn[8].n71 VGND 0.18333f
C10813 XThC.Tn[8].n72 VGND 0.02883f
C10814 XThC.Tn[8].t2 VGND 0.02006f
C10815 XThC.Tn[8].t1 VGND 0.02006f
C10816 XThC.Tn[8].n73 VGND 0.0446f
C10817 XThC.Tn[8].t0 VGND 0.02006f
C10818 XThC.Tn[8].t3 VGND 0.02006f
C10819 XThC.Tn[8].n74 VGND 0.06092f
C10820 XThC.Tn[8].n75 VGND 0.1985f
C10821 XThC.XTB1.Y.t2 VGND 0.03224f
C10822 XThC.XTB1.Y.n0 VGND 0.02084f
C10823 XThC.XTB1.Y.n1 VGND 0.02659f
C10824 XThC.XTB1.Y.t1 VGND 0.01618f
C10825 XThC.XTB1.Y.t0 VGND 0.01618f
C10826 XThC.XTB1.Y.n2 VGND 0.03473f
C10827 XThC.XTB1.Y.t17 VGND 0.02517f
C10828 XThC.XTB1.Y.t5 VGND 0.01483f
C10829 XThC.XTB1.Y.n3 VGND 0.02997f
C10830 XThC.XTB1.Y.t6 VGND 0.02517f
C10831 XThC.XTB1.Y.t12 VGND 0.01483f
C10832 XThC.XTB1.Y.n4 VGND 0.01542f
C10833 XThC.XTB1.Y.t8 VGND 0.02517f
C10834 XThC.XTB1.Y.t13 VGND 0.01483f
C10835 XThC.XTB1.Y.n5 VGND 0.03313f
C10836 XThC.XTB1.Y.t11 VGND 0.02517f
C10837 XThC.XTB1.Y.t16 VGND 0.01483f
C10838 XThC.XTB1.Y.n6 VGND 0.03076f
C10839 XThC.XTB1.Y.n7 VGND 0.01871f
C10840 XThC.XTB1.Y.n8 VGND 0.03098f
C10841 XThC.XTB1.Y.n9 VGND 0.01198f
C10842 XThC.XTB1.Y.n10 VGND 0.01463f
C10843 XThC.XTB1.Y.n11 VGND 0.03313f
C10844 XThC.XTB1.Y.n12 VGND 0.01661f
C10845 XThC.XTB1.Y.n13 VGND 0.02824f
C10846 XThC.XTB1.Y.t18 VGND 0.02517f
C10847 XThC.XTB1.Y.t9 VGND 0.01483f
C10848 XThC.XTB1.Y.n14 VGND 0.03392f
C10849 XThC.XTB1.Y.t7 VGND 0.02517f
C10850 XThC.XTB1.Y.t15 VGND 0.01483f
C10851 XThC.XTB1.Y.t14 VGND 0.02517f
C10852 XThC.XTB1.Y.t3 VGND 0.01483f
C10853 XThC.XTB1.Y.t10 VGND 0.02517f
C10854 XThC.XTB1.Y.t4 VGND 0.01483f
C10855 XThC.XTB1.Y.n15 VGND 0.04223f
C10856 XThC.XTB1.Y.n16 VGND 0.0446f
C10857 XThC.XTB1.Y.n17 VGND 0.01719f
C10858 XThC.XTB1.Y.n18 VGND 0.0363f
C10859 XThC.XTB1.Y.n19 VGND 0.01661f
C10860 XThC.XTB1.Y.n20 VGND 0.01378f
C10861 XThC.XTB1.Y.n21 VGND 0.77148f
C10862 XThC.XTB1.Y.n22 VGND 0.07634f
C10863 XThC.Tn[14].t4 VGND 0.01262f
C10864 XThC.Tn[14].t6 VGND 0.01262f
C10865 XThC.Tn[14].n0 VGND 0.03148f
C10866 XThC.Tn[14].t5 VGND 0.01262f
C10867 XThC.Tn[14].t7 VGND 0.01262f
C10868 XThC.Tn[14].n1 VGND 0.02524f
C10869 XThC.Tn[14].n2 VGND 0.06349f
C10870 XThC.Tn[14].t43 VGND 0.01539f
C10871 XThC.Tn[14].t38 VGND 0.01681f
C10872 XThC.Tn[14].n3 VGND 0.03752f
C10873 XThC.Tn[14].n4 VGND 0.02571f
C10874 XThC.Tn[14].n5 VGND 0.08438f
C10875 XThC.Tn[14].t29 VGND 0.01539f
C10876 XThC.Tn[14].t22 VGND 0.01681f
C10877 XThC.Tn[14].n6 VGND 0.03752f
C10878 XThC.Tn[14].n7 VGND 0.02571f
C10879 XThC.Tn[14].n8 VGND 0.08461f
C10880 XThC.Tn[14].n9 VGND 0.13945f
C10881 XThC.Tn[14].t32 VGND 0.01539f
C10882 XThC.Tn[14].t25 VGND 0.01681f
C10883 XThC.Tn[14].n10 VGND 0.03752f
C10884 XThC.Tn[14].n11 VGND 0.02571f
C10885 XThC.Tn[14].n12 VGND 0.08461f
C10886 XThC.Tn[14].n13 VGND 0.13945f
C10887 XThC.Tn[14].t34 VGND 0.01539f
C10888 XThC.Tn[14].t26 VGND 0.01681f
C10889 XThC.Tn[14].n14 VGND 0.03752f
C10890 XThC.Tn[14].n15 VGND 0.02571f
C10891 XThC.Tn[14].n16 VGND 0.08461f
C10892 XThC.Tn[14].n17 VGND 0.13945f
C10893 XThC.Tn[14].t20 VGND 0.01539f
C10894 XThC.Tn[14].t14 VGND 0.01681f
C10895 XThC.Tn[14].n18 VGND 0.03752f
C10896 XThC.Tn[14].n19 VGND 0.02571f
C10897 XThC.Tn[14].n20 VGND 0.08461f
C10898 XThC.Tn[14].n21 VGND 0.13945f
C10899 XThC.Tn[14].t23 VGND 0.01539f
C10900 XThC.Tn[14].t17 VGND 0.01681f
C10901 XThC.Tn[14].n22 VGND 0.03752f
C10902 XThC.Tn[14].n23 VGND 0.02571f
C10903 XThC.Tn[14].n24 VGND 0.08461f
C10904 XThC.Tn[14].n25 VGND 0.13945f
C10905 XThC.Tn[14].t37 VGND 0.01539f
C10906 XThC.Tn[14].t31 VGND 0.01681f
C10907 XThC.Tn[14].n26 VGND 0.03752f
C10908 XThC.Tn[14].n27 VGND 0.02571f
C10909 XThC.Tn[14].n28 VGND 0.08461f
C10910 XThC.Tn[14].n29 VGND 0.13945f
C10911 XThC.Tn[14].t13 VGND 0.01539f
C10912 XThC.Tn[14].t39 VGND 0.01681f
C10913 XThC.Tn[14].n30 VGND 0.03752f
C10914 XThC.Tn[14].n31 VGND 0.02571f
C10915 XThC.Tn[14].n32 VGND 0.08461f
C10916 XThC.Tn[14].n33 VGND 0.13945f
C10917 XThC.Tn[14].t15 VGND 0.01539f
C10918 XThC.Tn[14].t41 VGND 0.01681f
C10919 XThC.Tn[14].n34 VGND 0.03752f
C10920 XThC.Tn[14].n35 VGND 0.02571f
C10921 XThC.Tn[14].n36 VGND 0.08461f
C10922 XThC.Tn[14].n37 VGND 0.13945f
C10923 XThC.Tn[14].t35 VGND 0.01539f
C10924 XThC.Tn[14].t27 VGND 0.01681f
C10925 XThC.Tn[14].n38 VGND 0.03752f
C10926 XThC.Tn[14].n39 VGND 0.02571f
C10927 XThC.Tn[14].n40 VGND 0.08461f
C10928 XThC.Tn[14].n41 VGND 0.13945f
C10929 XThC.Tn[14].t36 VGND 0.01539f
C10930 XThC.Tn[14].t30 VGND 0.01681f
C10931 XThC.Tn[14].n42 VGND 0.03752f
C10932 XThC.Tn[14].n43 VGND 0.02571f
C10933 XThC.Tn[14].n44 VGND 0.08461f
C10934 XThC.Tn[14].n45 VGND 0.13945f
C10935 XThC.Tn[14].t16 VGND 0.01539f
C10936 XThC.Tn[14].t42 VGND 0.01681f
C10937 XThC.Tn[14].n46 VGND 0.03752f
C10938 XThC.Tn[14].n47 VGND 0.02571f
C10939 XThC.Tn[14].n48 VGND 0.08461f
C10940 XThC.Tn[14].n49 VGND 0.13945f
C10941 XThC.Tn[14].t24 VGND 0.01539f
C10942 XThC.Tn[14].t19 VGND 0.01681f
C10943 XThC.Tn[14].n50 VGND 0.03752f
C10944 XThC.Tn[14].n51 VGND 0.02571f
C10945 XThC.Tn[14].n52 VGND 0.08461f
C10946 XThC.Tn[14].n53 VGND 0.13945f
C10947 XThC.Tn[14].t28 VGND 0.01539f
C10948 XThC.Tn[14].t21 VGND 0.01681f
C10949 XThC.Tn[14].n54 VGND 0.03752f
C10950 XThC.Tn[14].n55 VGND 0.02571f
C10951 XThC.Tn[14].n56 VGND 0.08461f
C10952 XThC.Tn[14].n57 VGND 0.13945f
C10953 XThC.Tn[14].t40 VGND 0.01539f
C10954 XThC.Tn[14].t33 VGND 0.01681f
C10955 XThC.Tn[14].n58 VGND 0.03752f
C10956 XThC.Tn[14].n59 VGND 0.02571f
C10957 XThC.Tn[14].n60 VGND 0.08461f
C10958 XThC.Tn[14].n61 VGND 0.13945f
C10959 XThC.Tn[14].t18 VGND 0.01539f
C10960 XThC.Tn[14].t12 VGND 0.01681f
C10961 XThC.Tn[14].n62 VGND 0.03752f
C10962 XThC.Tn[14].n63 VGND 0.02571f
C10963 XThC.Tn[14].n64 VGND 0.08461f
C10964 XThC.Tn[14].n65 VGND 0.13945f
C10965 XThC.Tn[14].n66 VGND 0.91462f
C10966 XThC.Tn[14].n67 VGND 0.26906f
C10967 XThC.Tn[14].t8 VGND 0.01942f
C10968 XThC.Tn[14].t9 VGND 0.01942f
C10969 XThC.Tn[14].n68 VGND 0.04195f
C10970 XThC.Tn[14].t11 VGND 0.01942f
C10971 XThC.Tn[14].t10 VGND 0.01942f
C10972 XThC.Tn[14].n69 VGND 0.06385f
C10973 XThC.Tn[14].n70 VGND 0.1774f
C10974 XThC.Tn[14].n71 VGND 0.02789f
C10975 XThC.Tn[14].t1 VGND 0.01942f
C10976 XThC.Tn[14].t0 VGND 0.01942f
C10977 XThC.Tn[14].n72 VGND 0.04316f
C10978 XThC.Tn[14].t3 VGND 0.01942f
C10979 XThC.Tn[14].t2 VGND 0.01942f
C10980 XThC.Tn[14].n73 VGND 0.05895f
C10981 XThC.Tn[14].n74 VGND 0.19209f
C10982 XThR.Tn[10].t6 VGND 0.02415f
C10983 XThR.Tn[10].t4 VGND 0.02415f
C10984 XThR.Tn[10].n0 VGND 0.07333f
C10985 XThR.Tn[10].t7 VGND 0.02415f
C10986 XThR.Tn[10].t5 VGND 0.02415f
C10987 XThR.Tn[10].n1 VGND 0.05368f
C10988 XThR.Tn[10].n2 VGND 0.2441f
C10989 XThR.Tn[10].t3 VGND 0.02415f
C10990 XThR.Tn[10].t8 VGND 0.02415f
C10991 XThR.Tn[10].n3 VGND 0.05218f
C10992 XThR.Tn[10].t10 VGND 0.02415f
C10993 XThR.Tn[10].t1 VGND 0.02415f
C10994 XThR.Tn[10].n4 VGND 0.07942f
C10995 XThR.Tn[10].n5 VGND 0.22051f
C10996 XThR.Tn[10].n6 VGND 0.01087f
C10997 XThR.Tn[10].t54 VGND 0.01887f
C10998 XThR.Tn[10].t47 VGND 0.02067f
C10999 XThR.Tn[10].n7 VGND 0.05047f
C11000 XThR.Tn[10].n8 VGND 0.09695f
C11001 XThR.Tn[10].t13 VGND 0.01887f
C11002 XThR.Tn[10].t63 VGND 0.02067f
C11003 XThR.Tn[10].n9 VGND 0.05047f
C11004 XThR.Tn[10].t50 VGND 0.01881f
C11005 XThR.Tn[10].t60 VGND 0.0206f
C11006 XThR.Tn[10].n10 VGND 0.05251f
C11007 XThR.Tn[10].n11 VGND 0.03689f
C11008 XThR.Tn[10].n12 VGND 0.00674f
C11009 XThR.Tn[10].n13 VGND 0.11838f
C11010 XThR.Tn[10].t48 VGND 0.01887f
C11011 XThR.Tn[10].t41 VGND 0.02067f
C11012 XThR.Tn[10].n14 VGND 0.05047f
C11013 XThR.Tn[10].t23 VGND 0.01881f
C11014 XThR.Tn[10].t36 VGND 0.0206f
C11015 XThR.Tn[10].n15 VGND 0.05251f
C11016 XThR.Tn[10].n16 VGND 0.03689f
C11017 XThR.Tn[10].n17 VGND 0.00674f
C11018 XThR.Tn[10].n18 VGND 0.11838f
C11019 XThR.Tn[10].t65 VGND 0.01887f
C11020 XThR.Tn[10].t58 VGND 0.02067f
C11021 XThR.Tn[10].n19 VGND 0.05047f
C11022 XThR.Tn[10].t40 VGND 0.01881f
C11023 XThR.Tn[10].t55 VGND 0.0206f
C11024 XThR.Tn[10].n20 VGND 0.05251f
C11025 XThR.Tn[10].n21 VGND 0.03689f
C11026 XThR.Tn[10].n22 VGND 0.00674f
C11027 XThR.Tn[10].n23 VGND 0.11838f
C11028 XThR.Tn[10].t30 VGND 0.01887f
C11029 XThR.Tn[10].t26 VGND 0.02067f
C11030 XThR.Tn[10].n24 VGND 0.05047f
C11031 XThR.Tn[10].t70 VGND 0.01881f
C11032 XThR.Tn[10].t21 VGND 0.0206f
C11033 XThR.Tn[10].n25 VGND 0.05251f
C11034 XThR.Tn[10].n26 VGND 0.03689f
C11035 XThR.Tn[10].n27 VGND 0.00674f
C11036 XThR.Tn[10].n28 VGND 0.11838f
C11037 XThR.Tn[10].t67 VGND 0.01887f
C11038 XThR.Tn[10].t59 VGND 0.02067f
C11039 XThR.Tn[10].n29 VGND 0.05047f
C11040 XThR.Tn[10].t42 VGND 0.01881f
C11041 XThR.Tn[10].t56 VGND 0.0206f
C11042 XThR.Tn[10].n30 VGND 0.05251f
C11043 XThR.Tn[10].n31 VGND 0.03689f
C11044 XThR.Tn[10].n32 VGND 0.00674f
C11045 XThR.Tn[10].n33 VGND 0.11838f
C11046 XThR.Tn[10].t44 VGND 0.01887f
C11047 XThR.Tn[10].t15 VGND 0.02067f
C11048 XThR.Tn[10].n34 VGND 0.05047f
C11049 XThR.Tn[10].t18 VGND 0.01881f
C11050 XThR.Tn[10].t12 VGND 0.0206f
C11051 XThR.Tn[10].n35 VGND 0.05251f
C11052 XThR.Tn[10].n36 VGND 0.03689f
C11053 XThR.Tn[10].n37 VGND 0.00674f
C11054 XThR.Tn[10].n38 VGND 0.11838f
C11055 XThR.Tn[10].t14 VGND 0.01887f
C11056 XThR.Tn[10].t69 VGND 0.02067f
C11057 XThR.Tn[10].n39 VGND 0.05047f
C11058 XThR.Tn[10].t51 VGND 0.01881f
C11059 XThR.Tn[10].t66 VGND 0.0206f
C11060 XThR.Tn[10].n40 VGND 0.05251f
C11061 XThR.Tn[10].n41 VGND 0.03689f
C11062 XThR.Tn[10].n42 VGND 0.00674f
C11063 XThR.Tn[10].n43 VGND 0.11838f
C11064 XThR.Tn[10].t17 VGND 0.01887f
C11065 XThR.Tn[10].t24 VGND 0.02067f
C11066 XThR.Tn[10].n44 VGND 0.05047f
C11067 XThR.Tn[10].t53 VGND 0.01881f
C11068 XThR.Tn[10].t20 VGND 0.0206f
C11069 XThR.Tn[10].n45 VGND 0.05251f
C11070 XThR.Tn[10].n46 VGND 0.03689f
C11071 XThR.Tn[10].n47 VGND 0.00674f
C11072 XThR.Tn[10].n48 VGND 0.11838f
C11073 XThR.Tn[10].t33 VGND 0.01887f
C11074 XThR.Tn[10].t43 VGND 0.02067f
C11075 XThR.Tn[10].n49 VGND 0.05047f
C11076 XThR.Tn[10].t73 VGND 0.01881f
C11077 XThR.Tn[10].t38 VGND 0.0206f
C11078 XThR.Tn[10].n50 VGND 0.05251f
C11079 XThR.Tn[10].n51 VGND 0.03689f
C11080 XThR.Tn[10].n52 VGND 0.00674f
C11081 XThR.Tn[10].n53 VGND 0.11838f
C11082 XThR.Tn[10].t28 VGND 0.01887f
C11083 XThR.Tn[10].t61 VGND 0.02067f
C11084 XThR.Tn[10].n54 VGND 0.05047f
C11085 XThR.Tn[10].t62 VGND 0.01881f
C11086 XThR.Tn[10].t57 VGND 0.0206f
C11087 XThR.Tn[10].n55 VGND 0.05251f
C11088 XThR.Tn[10].n56 VGND 0.03689f
C11089 XThR.Tn[10].n57 VGND 0.00674f
C11090 XThR.Tn[10].n58 VGND 0.11838f
C11091 XThR.Tn[10].t46 VGND 0.01887f
C11092 XThR.Tn[10].t35 VGND 0.02067f
C11093 XThR.Tn[10].n59 VGND 0.05047f
C11094 XThR.Tn[10].t19 VGND 0.01881f
C11095 XThR.Tn[10].t32 VGND 0.0206f
C11096 XThR.Tn[10].n60 VGND 0.05251f
C11097 XThR.Tn[10].n61 VGND 0.03689f
C11098 XThR.Tn[10].n62 VGND 0.00674f
C11099 XThR.Tn[10].n63 VGND 0.11838f
C11100 XThR.Tn[10].t16 VGND 0.01887f
C11101 XThR.Tn[10].t72 VGND 0.02067f
C11102 XThR.Tn[10].n64 VGND 0.05047f
C11103 XThR.Tn[10].t52 VGND 0.01881f
C11104 XThR.Tn[10].t68 VGND 0.0206f
C11105 XThR.Tn[10].n65 VGND 0.05251f
C11106 XThR.Tn[10].n66 VGND 0.03689f
C11107 XThR.Tn[10].n67 VGND 0.00674f
C11108 XThR.Tn[10].n68 VGND 0.11838f
C11109 XThR.Tn[10].t31 VGND 0.01887f
C11110 XThR.Tn[10].t27 VGND 0.02067f
C11111 XThR.Tn[10].n69 VGND 0.05047f
C11112 XThR.Tn[10].t71 VGND 0.01881f
C11113 XThR.Tn[10].t22 VGND 0.0206f
C11114 XThR.Tn[10].n70 VGND 0.05251f
C11115 XThR.Tn[10].n71 VGND 0.03689f
C11116 XThR.Tn[10].n72 VGND 0.00674f
C11117 XThR.Tn[10].n73 VGND 0.11838f
C11118 XThR.Tn[10].t49 VGND 0.01887f
C11119 XThR.Tn[10].t45 VGND 0.02067f
C11120 XThR.Tn[10].n74 VGND 0.05047f
C11121 XThR.Tn[10].t25 VGND 0.01881f
C11122 XThR.Tn[10].t39 VGND 0.0206f
C11123 XThR.Tn[10].n75 VGND 0.05251f
C11124 XThR.Tn[10].n76 VGND 0.03689f
C11125 XThR.Tn[10].n77 VGND 0.00674f
C11126 XThR.Tn[10].n78 VGND 0.11838f
C11127 XThR.Tn[10].t29 VGND 0.01887f
C11128 XThR.Tn[10].t37 VGND 0.02067f
C11129 XThR.Tn[10].n79 VGND 0.05047f
C11130 XThR.Tn[10].t64 VGND 0.01881f
C11131 XThR.Tn[10].t34 VGND 0.0206f
C11132 XThR.Tn[10].n80 VGND 0.05251f
C11133 XThR.Tn[10].n81 VGND 0.03689f
C11134 XThR.Tn[10].n82 VGND 0.00674f
C11135 XThR.Tn[10].n83 VGND 0.11838f
C11136 XThR.Tn[10].n84 VGND 0.10758f
C11137 XThR.Tn[10].n85 VGND 0.3312f
C11138 XThR.Tn[10].t2 VGND 0.0157f
C11139 XThR.Tn[10].t11 VGND 0.0157f
C11140 XThR.Tn[10].n86 VGND 0.03915f
C11141 XThR.Tn[10].t9 VGND 0.0157f
C11142 XThR.Tn[10].t0 VGND 0.0157f
C11143 XThR.Tn[10].n87 VGND 0.0314f
C11144 XThR.Tn[10].n88 VGND 0.07239f
C11145 XThC.Tn[3].t5 VGND 0.01826f
C11146 XThC.Tn[3].t4 VGND 0.01826f
C11147 XThC.Tn[3].n0 VGND 0.03685f
C11148 XThC.Tn[3].t7 VGND 0.01826f
C11149 XThC.Tn[3].t6 VGND 0.01826f
C11150 XThC.Tn[3].n1 VGND 0.04312f
C11151 XThC.Tn[3].n2 VGND 0.12934f
C11152 XThC.Tn[3].t1 VGND 0.01187f
C11153 XThC.Tn[3].t0 VGND 0.01187f
C11154 XThC.Tn[3].n3 VGND 0.02703f
C11155 XThC.Tn[3].t11 VGND 0.01187f
C11156 XThC.Tn[3].t10 VGND 0.01187f
C11157 XThC.Tn[3].n4 VGND 0.04503f
C11158 XThC.Tn[3].t9 VGND 0.01187f
C11159 XThC.Tn[3].t8 VGND 0.01187f
C11160 XThC.Tn[3].n5 VGND 0.02703f
C11161 XThC.Tn[3].n6 VGND 0.1287f
C11162 XThC.Tn[3].t3 VGND 0.01187f
C11163 XThC.Tn[3].t2 VGND 0.01187f
C11164 XThC.Tn[3].n7 VGND 0.02703f
C11165 XThC.Tn[3].n8 VGND 0.07956f
C11166 XThC.Tn[3].n9 VGND 0.08979f
C11167 XThC.Tn[3].t12 VGND 0.01447f
C11168 XThC.Tn[3].t42 VGND 0.01581f
C11169 XThC.Tn[3].n10 VGND 0.03529f
C11170 XThC.Tn[3].n11 VGND 0.02417f
C11171 XThC.Tn[3].n12 VGND 0.07935f
C11172 XThC.Tn[3].t30 VGND 0.01447f
C11173 XThC.Tn[3].t27 VGND 0.01581f
C11174 XThC.Tn[3].n13 VGND 0.03529f
C11175 XThC.Tn[3].n14 VGND 0.02417f
C11176 XThC.Tn[3].n15 VGND 0.07957f
C11177 XThC.Tn[3].n16 VGND 0.13113f
C11178 XThC.Tn[3].t35 VGND 0.01447f
C11179 XThC.Tn[3].t29 VGND 0.01581f
C11180 XThC.Tn[3].n17 VGND 0.03529f
C11181 XThC.Tn[3].n18 VGND 0.02417f
C11182 XThC.Tn[3].n19 VGND 0.07957f
C11183 XThC.Tn[3].n20 VGND 0.13113f
C11184 XThC.Tn[3].t36 VGND 0.01447f
C11185 XThC.Tn[3].t31 VGND 0.01581f
C11186 XThC.Tn[3].n21 VGND 0.03529f
C11187 XThC.Tn[3].n22 VGND 0.02417f
C11188 XThC.Tn[3].n23 VGND 0.07957f
C11189 XThC.Tn[3].n24 VGND 0.13113f
C11190 XThC.Tn[3].t23 VGND 0.01447f
C11191 XThC.Tn[3].t20 VGND 0.01581f
C11192 XThC.Tn[3].n25 VGND 0.03529f
C11193 XThC.Tn[3].n26 VGND 0.02417f
C11194 XThC.Tn[3].n27 VGND 0.07957f
C11195 XThC.Tn[3].n28 VGND 0.13113f
C11196 XThC.Tn[3].t24 VGND 0.01447f
C11197 XThC.Tn[3].t21 VGND 0.01581f
C11198 XThC.Tn[3].n29 VGND 0.03529f
C11199 XThC.Tn[3].n30 VGND 0.02417f
C11200 XThC.Tn[3].n31 VGND 0.07957f
C11201 XThC.Tn[3].n32 VGND 0.13113f
C11202 XThC.Tn[3].t40 VGND 0.01447f
C11203 XThC.Tn[3].t34 VGND 0.01581f
C11204 XThC.Tn[3].n33 VGND 0.03529f
C11205 XThC.Tn[3].n34 VGND 0.02417f
C11206 XThC.Tn[3].n35 VGND 0.07957f
C11207 XThC.Tn[3].n36 VGND 0.13113f
C11208 XThC.Tn[3].t15 VGND 0.01447f
C11209 XThC.Tn[3].t43 VGND 0.01581f
C11210 XThC.Tn[3].n37 VGND 0.03529f
C11211 XThC.Tn[3].n38 VGND 0.02417f
C11212 XThC.Tn[3].n39 VGND 0.07957f
C11213 XThC.Tn[3].n40 VGND 0.13113f
C11214 XThC.Tn[3].t17 VGND 0.01447f
C11215 XThC.Tn[3].t13 VGND 0.01581f
C11216 XThC.Tn[3].n41 VGND 0.03529f
C11217 XThC.Tn[3].n42 VGND 0.02417f
C11218 XThC.Tn[3].n43 VGND 0.07957f
C11219 XThC.Tn[3].n44 VGND 0.13113f
C11220 XThC.Tn[3].t37 VGND 0.01447f
C11221 XThC.Tn[3].t32 VGND 0.01581f
C11222 XThC.Tn[3].n45 VGND 0.03529f
C11223 XThC.Tn[3].n46 VGND 0.02417f
C11224 XThC.Tn[3].n47 VGND 0.07957f
C11225 XThC.Tn[3].n48 VGND 0.13113f
C11226 XThC.Tn[3].t39 VGND 0.01447f
C11227 XThC.Tn[3].t33 VGND 0.01581f
C11228 XThC.Tn[3].n49 VGND 0.03529f
C11229 XThC.Tn[3].n50 VGND 0.02417f
C11230 XThC.Tn[3].n51 VGND 0.07957f
C11231 XThC.Tn[3].n52 VGND 0.13113f
C11232 XThC.Tn[3].t18 VGND 0.01447f
C11233 XThC.Tn[3].t14 VGND 0.01581f
C11234 XThC.Tn[3].n53 VGND 0.03529f
C11235 XThC.Tn[3].n54 VGND 0.02417f
C11236 XThC.Tn[3].n55 VGND 0.07957f
C11237 XThC.Tn[3].n56 VGND 0.13113f
C11238 XThC.Tn[3].t26 VGND 0.01447f
C11239 XThC.Tn[3].t22 VGND 0.01581f
C11240 XThC.Tn[3].n57 VGND 0.03529f
C11241 XThC.Tn[3].n58 VGND 0.02417f
C11242 XThC.Tn[3].n59 VGND 0.07957f
C11243 XThC.Tn[3].n60 VGND 0.13113f
C11244 XThC.Tn[3].t28 VGND 0.01447f
C11245 XThC.Tn[3].t25 VGND 0.01581f
C11246 XThC.Tn[3].n61 VGND 0.03529f
C11247 XThC.Tn[3].n62 VGND 0.02417f
C11248 XThC.Tn[3].n63 VGND 0.07957f
C11249 XThC.Tn[3].n64 VGND 0.13113f
C11250 XThC.Tn[3].t41 VGND 0.01447f
C11251 XThC.Tn[3].t38 VGND 0.01581f
C11252 XThC.Tn[3].n65 VGND 0.03529f
C11253 XThC.Tn[3].n66 VGND 0.02417f
C11254 XThC.Tn[3].n67 VGND 0.07957f
C11255 XThC.Tn[3].n68 VGND 0.13113f
C11256 XThC.Tn[3].t19 VGND 0.01447f
C11257 XThC.Tn[3].t16 VGND 0.01581f
C11258 XThC.Tn[3].n69 VGND 0.03529f
C11259 XThC.Tn[3].n70 VGND 0.02417f
C11260 XThC.Tn[3].n71 VGND 0.07957f
C11261 XThC.Tn[3].n72 VGND 0.13113f
C11262 XThC.Tn[3].n73 VGND 0.77119f
C11263 XThC.Tn[3].n74 VGND 0.1112f
C11264 XThC.Tn[1].t3 VGND 0.01715f
C11265 XThC.Tn[1].t2 VGND 0.01715f
C11266 XThC.Tn[1].n0 VGND 0.03462f
C11267 XThC.Tn[1].t1 VGND 0.01715f
C11268 XThC.Tn[1].t0 VGND 0.01715f
C11269 XThC.Tn[1].n1 VGND 0.04051f
C11270 XThC.Tn[1].n2 VGND 0.12152f
C11271 XThC.Tn[1].t11 VGND 0.01115f
C11272 XThC.Tn[1].t10 VGND 0.01115f
C11273 XThC.Tn[1].n3 VGND 0.04231f
C11274 XThC.Tn[1].t9 VGND 0.01115f
C11275 XThC.Tn[1].t8 VGND 0.01115f
C11276 XThC.Tn[1].n4 VGND 0.02539f
C11277 XThC.Tn[1].n5 VGND 0.12091f
C11278 XThC.Tn[1].t7 VGND 0.01115f
C11279 XThC.Tn[1].t6 VGND 0.01115f
C11280 XThC.Tn[1].n6 VGND 0.02539f
C11281 XThC.Tn[1].n7 VGND 0.07475f
C11282 XThC.Tn[1].t5 VGND 0.01115f
C11283 XThC.Tn[1].t4 VGND 0.01115f
C11284 XThC.Tn[1].n8 VGND 0.02539f
C11285 XThC.Tn[1].n9 VGND 0.08436f
C11286 XThC.Tn[1].t31 VGND 0.0136f
C11287 XThC.Tn[1].t29 VGND 0.01485f
C11288 XThC.Tn[1].n10 VGND 0.03315f
C11289 XThC.Tn[1].n11 VGND 0.02271f
C11290 XThC.Tn[1].n12 VGND 0.07455f
C11291 XThC.Tn[1].t17 VGND 0.0136f
C11292 XThC.Tn[1].t14 VGND 0.01485f
C11293 XThC.Tn[1].n13 VGND 0.03315f
C11294 XThC.Tn[1].n14 VGND 0.02271f
C11295 XThC.Tn[1].n15 VGND 0.07475f
C11296 XThC.Tn[1].n16 VGND 0.1232f
C11297 XThC.Tn[1].t22 VGND 0.0136f
C11298 XThC.Tn[1].t16 VGND 0.01485f
C11299 XThC.Tn[1].n17 VGND 0.03315f
C11300 XThC.Tn[1].n18 VGND 0.02271f
C11301 XThC.Tn[1].n19 VGND 0.07475f
C11302 XThC.Tn[1].n20 VGND 0.1232f
C11303 XThC.Tn[1].t23 VGND 0.0136f
C11304 XThC.Tn[1].t18 VGND 0.01485f
C11305 XThC.Tn[1].n21 VGND 0.03315f
C11306 XThC.Tn[1].n22 VGND 0.02271f
C11307 XThC.Tn[1].n23 VGND 0.07475f
C11308 XThC.Tn[1].n24 VGND 0.1232f
C11309 XThC.Tn[1].t42 VGND 0.0136f
C11310 XThC.Tn[1].t39 VGND 0.01485f
C11311 XThC.Tn[1].n25 VGND 0.03315f
C11312 XThC.Tn[1].n26 VGND 0.02271f
C11313 XThC.Tn[1].n27 VGND 0.07475f
C11314 XThC.Tn[1].n28 VGND 0.1232f
C11315 XThC.Tn[1].t43 VGND 0.0136f
C11316 XThC.Tn[1].t40 VGND 0.01485f
C11317 XThC.Tn[1].n29 VGND 0.03315f
C11318 XThC.Tn[1].n30 VGND 0.02271f
C11319 XThC.Tn[1].n31 VGND 0.07475f
C11320 XThC.Tn[1].n32 VGND 0.1232f
C11321 XThC.Tn[1].t27 VGND 0.0136f
C11322 XThC.Tn[1].t21 VGND 0.01485f
C11323 XThC.Tn[1].n33 VGND 0.03315f
C11324 XThC.Tn[1].n34 VGND 0.02271f
C11325 XThC.Tn[1].n35 VGND 0.07475f
C11326 XThC.Tn[1].n36 VGND 0.1232f
C11327 XThC.Tn[1].t34 VGND 0.0136f
C11328 XThC.Tn[1].t30 VGND 0.01485f
C11329 XThC.Tn[1].n37 VGND 0.03315f
C11330 XThC.Tn[1].n38 VGND 0.02271f
C11331 XThC.Tn[1].n39 VGND 0.07475f
C11332 XThC.Tn[1].n40 VGND 0.1232f
C11333 XThC.Tn[1].t36 VGND 0.0136f
C11334 XThC.Tn[1].t32 VGND 0.01485f
C11335 XThC.Tn[1].n41 VGND 0.03315f
C11336 XThC.Tn[1].n42 VGND 0.02271f
C11337 XThC.Tn[1].n43 VGND 0.07475f
C11338 XThC.Tn[1].n44 VGND 0.1232f
C11339 XThC.Tn[1].t24 VGND 0.0136f
C11340 XThC.Tn[1].t19 VGND 0.01485f
C11341 XThC.Tn[1].n45 VGND 0.03315f
C11342 XThC.Tn[1].n46 VGND 0.02271f
C11343 XThC.Tn[1].n47 VGND 0.07475f
C11344 XThC.Tn[1].n48 VGND 0.1232f
C11345 XThC.Tn[1].t26 VGND 0.0136f
C11346 XThC.Tn[1].t20 VGND 0.01485f
C11347 XThC.Tn[1].n49 VGND 0.03315f
C11348 XThC.Tn[1].n50 VGND 0.02271f
C11349 XThC.Tn[1].n51 VGND 0.07475f
C11350 XThC.Tn[1].n52 VGND 0.1232f
C11351 XThC.Tn[1].t37 VGND 0.0136f
C11352 XThC.Tn[1].t33 VGND 0.01485f
C11353 XThC.Tn[1].n53 VGND 0.03315f
C11354 XThC.Tn[1].n54 VGND 0.02271f
C11355 XThC.Tn[1].n55 VGND 0.07475f
C11356 XThC.Tn[1].n56 VGND 0.1232f
C11357 XThC.Tn[1].t13 VGND 0.0136f
C11358 XThC.Tn[1].t41 VGND 0.01485f
C11359 XThC.Tn[1].n57 VGND 0.03315f
C11360 XThC.Tn[1].n58 VGND 0.02271f
C11361 XThC.Tn[1].n59 VGND 0.07475f
C11362 XThC.Tn[1].n60 VGND 0.1232f
C11363 XThC.Tn[1].t15 VGND 0.0136f
C11364 XThC.Tn[1].t12 VGND 0.01485f
C11365 XThC.Tn[1].n61 VGND 0.03315f
C11366 XThC.Tn[1].n62 VGND 0.02271f
C11367 XThC.Tn[1].n63 VGND 0.07475f
C11368 XThC.Tn[1].n64 VGND 0.1232f
C11369 XThC.Tn[1].t28 VGND 0.0136f
C11370 XThC.Tn[1].t25 VGND 0.01485f
C11371 XThC.Tn[1].n65 VGND 0.03315f
C11372 XThC.Tn[1].n66 VGND 0.02271f
C11373 XThC.Tn[1].n67 VGND 0.07475f
C11374 XThC.Tn[1].n68 VGND 0.1232f
C11375 XThC.Tn[1].t38 VGND 0.0136f
C11376 XThC.Tn[1].t35 VGND 0.01485f
C11377 XThC.Tn[1].n69 VGND 0.03315f
C11378 XThC.Tn[1].n70 VGND 0.02271f
C11379 XThC.Tn[1].n71 VGND 0.07475f
C11380 XThC.Tn[1].n72 VGND 0.1232f
C11381 XThC.Tn[1].n73 VGND 0.62603f
C11382 XThC.Tn[1].n74 VGND 0.11896f
C11383 XThC.Tn[2].t11 VGND 0.0117f
C11384 XThC.Tn[2].t8 VGND 0.0117f
C11385 XThC.Tn[2].n0 VGND 0.04439f
C11386 XThC.Tn[2].t9 VGND 0.0117f
C11387 XThC.Tn[2].t10 VGND 0.0117f
C11388 XThC.Tn[2].n1 VGND 0.02664f
C11389 XThC.Tn[2].n2 VGND 0.12687f
C11390 XThC.Tn[2].t5 VGND 0.0117f
C11391 XThC.Tn[2].t4 VGND 0.0117f
C11392 XThC.Tn[2].n3 VGND 0.02664f
C11393 XThC.Tn[2].n4 VGND 0.07843f
C11394 XThC.Tn[2].t7 VGND 0.0117f
C11395 XThC.Tn[2].t6 VGND 0.0117f
C11396 XThC.Tn[2].n5 VGND 0.02664f
C11397 XThC.Tn[2].n6 VGND 0.08852f
C11398 XThC.Tn[2].t20 VGND 0.01427f
C11399 XThC.Tn[2].t18 VGND 0.01558f
C11400 XThC.Tn[2].n7 VGND 0.03478f
C11401 XThC.Tn[2].n8 VGND 0.02383f
C11402 XThC.Tn[2].n9 VGND 0.07822f
C11403 XThC.Tn[2].t38 VGND 0.01427f
C11404 XThC.Tn[2].t35 VGND 0.01558f
C11405 XThC.Tn[2].n10 VGND 0.03478f
C11406 XThC.Tn[2].n11 VGND 0.02383f
C11407 XThC.Tn[2].n12 VGND 0.07844f
C11408 XThC.Tn[2].n13 VGND 0.12927f
C11409 XThC.Tn[2].t43 VGND 0.01427f
C11410 XThC.Tn[2].t37 VGND 0.01558f
C11411 XThC.Tn[2].n14 VGND 0.03478f
C11412 XThC.Tn[2].n15 VGND 0.02383f
C11413 XThC.Tn[2].n16 VGND 0.07844f
C11414 XThC.Tn[2].n17 VGND 0.12927f
C11415 XThC.Tn[2].t12 VGND 0.01427f
C11416 XThC.Tn[2].t39 VGND 0.01558f
C11417 XThC.Tn[2].n18 VGND 0.03478f
C11418 XThC.Tn[2].n19 VGND 0.02383f
C11419 XThC.Tn[2].n20 VGND 0.07844f
C11420 XThC.Tn[2].n21 VGND 0.12927f
C11421 XThC.Tn[2].t31 VGND 0.01427f
C11422 XThC.Tn[2].t28 VGND 0.01558f
C11423 XThC.Tn[2].n22 VGND 0.03478f
C11424 XThC.Tn[2].n23 VGND 0.02383f
C11425 XThC.Tn[2].n24 VGND 0.07844f
C11426 XThC.Tn[2].n25 VGND 0.12927f
C11427 XThC.Tn[2].t32 VGND 0.01427f
C11428 XThC.Tn[2].t29 VGND 0.01558f
C11429 XThC.Tn[2].n26 VGND 0.03478f
C11430 XThC.Tn[2].n27 VGND 0.02383f
C11431 XThC.Tn[2].n28 VGND 0.07844f
C11432 XThC.Tn[2].n29 VGND 0.12927f
C11433 XThC.Tn[2].t16 VGND 0.01427f
C11434 XThC.Tn[2].t42 VGND 0.01558f
C11435 XThC.Tn[2].n30 VGND 0.03478f
C11436 XThC.Tn[2].n31 VGND 0.02383f
C11437 XThC.Tn[2].n32 VGND 0.07844f
C11438 XThC.Tn[2].n33 VGND 0.12927f
C11439 XThC.Tn[2].t23 VGND 0.01427f
C11440 XThC.Tn[2].t19 VGND 0.01558f
C11441 XThC.Tn[2].n34 VGND 0.03478f
C11442 XThC.Tn[2].n35 VGND 0.02383f
C11443 XThC.Tn[2].n36 VGND 0.07844f
C11444 XThC.Tn[2].n37 VGND 0.12927f
C11445 XThC.Tn[2].t25 VGND 0.01427f
C11446 XThC.Tn[2].t21 VGND 0.01558f
C11447 XThC.Tn[2].n38 VGND 0.03478f
C11448 XThC.Tn[2].n39 VGND 0.02383f
C11449 XThC.Tn[2].n40 VGND 0.07844f
C11450 XThC.Tn[2].n41 VGND 0.12927f
C11451 XThC.Tn[2].t13 VGND 0.01427f
C11452 XThC.Tn[2].t40 VGND 0.01558f
C11453 XThC.Tn[2].n42 VGND 0.03478f
C11454 XThC.Tn[2].n43 VGND 0.02383f
C11455 XThC.Tn[2].n44 VGND 0.07844f
C11456 XThC.Tn[2].n45 VGND 0.12927f
C11457 XThC.Tn[2].t15 VGND 0.01427f
C11458 XThC.Tn[2].t41 VGND 0.01558f
C11459 XThC.Tn[2].n46 VGND 0.03478f
C11460 XThC.Tn[2].n47 VGND 0.02383f
C11461 XThC.Tn[2].n48 VGND 0.07844f
C11462 XThC.Tn[2].n49 VGND 0.12927f
C11463 XThC.Tn[2].t26 VGND 0.01427f
C11464 XThC.Tn[2].t22 VGND 0.01558f
C11465 XThC.Tn[2].n50 VGND 0.03478f
C11466 XThC.Tn[2].n51 VGND 0.02383f
C11467 XThC.Tn[2].n52 VGND 0.07844f
C11468 XThC.Tn[2].n53 VGND 0.12927f
C11469 XThC.Tn[2].t34 VGND 0.01427f
C11470 XThC.Tn[2].t30 VGND 0.01558f
C11471 XThC.Tn[2].n54 VGND 0.03478f
C11472 XThC.Tn[2].n55 VGND 0.02383f
C11473 XThC.Tn[2].n56 VGND 0.07844f
C11474 XThC.Tn[2].n57 VGND 0.12927f
C11475 XThC.Tn[2].t36 VGND 0.01427f
C11476 XThC.Tn[2].t33 VGND 0.01558f
C11477 XThC.Tn[2].n58 VGND 0.03478f
C11478 XThC.Tn[2].n59 VGND 0.02383f
C11479 XThC.Tn[2].n60 VGND 0.07844f
C11480 XThC.Tn[2].n61 VGND 0.12927f
C11481 XThC.Tn[2].t17 VGND 0.01427f
C11482 XThC.Tn[2].t14 VGND 0.01558f
C11483 XThC.Tn[2].n62 VGND 0.03478f
C11484 XThC.Tn[2].n63 VGND 0.02383f
C11485 XThC.Tn[2].n64 VGND 0.07844f
C11486 XThC.Tn[2].n65 VGND 0.12927f
C11487 XThC.Tn[2].t27 VGND 0.01427f
C11488 XThC.Tn[2].t24 VGND 0.01558f
C11489 XThC.Tn[2].n66 VGND 0.03478f
C11490 XThC.Tn[2].n67 VGND 0.02383f
C11491 XThC.Tn[2].n68 VGND 0.07844f
C11492 XThC.Tn[2].n69 VGND 0.12927f
C11493 XThC.Tn[2].n70 VGND 0.50031f
C11494 XThC.Tn[2].n71 VGND 0.1061f
C11495 XThC.Tn[2].t1 VGND 0.018f
C11496 XThC.Tn[2].t0 VGND 0.018f
C11497 XThC.Tn[2].n72 VGND 0.04251f
C11498 XThC.Tn[2].t3 VGND 0.018f
C11499 XThC.Tn[2].t2 VGND 0.018f
C11500 XThC.Tn[2].n73 VGND 0.03633f
C11501 XThC.Tn[2].n74 VGND 0.119f
C11502 XThC.Tn[2].n75 VGND 0.03766f
C11503 Iout.n0 VGND 0.23929f
C11504 Iout.n1 VGND 1.25122f
C11505 Iout.n2 VGND 0.23929f
C11506 Iout.n3 VGND 0.23929f
C11507 Iout.t218 VGND 0.02304f
C11508 Iout.n4 VGND 0.05124f
C11509 Iout.n5 VGND 0.20242f
C11510 Iout.n6 VGND 0.23929f
C11511 Iout.n7 VGND 1.25122f
C11512 Iout.n8 VGND 0.23929f
C11513 Iout.t0 VGND 0.02304f
C11514 Iout.n9 VGND 0.05124f
C11515 Iout.n10 VGND 0.20242f
C11516 Iout.n11 VGND 0.23929f
C11517 Iout.n12 VGND 1.25122f
C11518 Iout.n13 VGND 0.23929f
C11519 Iout.t142 VGND 0.02304f
C11520 Iout.n14 VGND 0.05124f
C11521 Iout.n15 VGND 0.20242f
C11522 Iout.n16 VGND 0.23929f
C11523 Iout.n17 VGND 1.25122f
C11524 Iout.n18 VGND 0.23929f
C11525 Iout.t85 VGND 0.02304f
C11526 Iout.n19 VGND 0.05124f
C11527 Iout.n20 VGND 0.20242f
C11528 Iout.n21 VGND 0.49611f
C11529 Iout.t224 VGND 0.02304f
C11530 Iout.n22 VGND 0.05124f
C11531 Iout.n23 VGND 0.29851f
C11532 Iout.n24 VGND 0.23929f
C11533 Iout.n25 VGND 0.23929f
C11534 Iout.n26 VGND 0.23929f
C11535 Iout.n27 VGND 0.23929f
C11536 Iout.n28 VGND 0.23929f
C11537 Iout.n29 VGND 0.23929f
C11538 Iout.n30 VGND 0.23929f
C11539 Iout.n31 VGND 0.23929f
C11540 Iout.n32 VGND 0.23929f
C11541 Iout.n33 VGND 0.23929f
C11542 Iout.n34 VGND 0.23929f
C11543 Iout.n35 VGND 0.23929f
C11544 Iout.n36 VGND 0.23929f
C11545 Iout.n37 VGND 0.23929f
C11546 Iout.t92 VGND 0.02304f
C11547 Iout.n38 VGND 0.05124f
C11548 Iout.n39 VGND 0.02606f
C11549 Iout.n40 VGND 0.23929f
C11550 Iout.n41 VGND 0.04775f
C11551 Iout.t30 VGND 0.02304f
C11552 Iout.n42 VGND 0.05124f
C11553 Iout.n43 VGND 0.02606f
C11554 Iout.t100 VGND 0.02304f
C11555 Iout.n44 VGND 0.05124f
C11556 Iout.n45 VGND 0.02606f
C11557 Iout.n46 VGND 0.23929f
C11558 Iout.t168 VGND 0.02304f
C11559 Iout.n47 VGND 0.05124f
C11560 Iout.n48 VGND 0.02606f
C11561 Iout.n49 VGND 0.23929f
C11562 Iout.t56 VGND 0.02304f
C11563 Iout.n50 VGND 0.05124f
C11564 Iout.n51 VGND 0.02606f
C11565 Iout.n52 VGND 0.23929f
C11566 Iout.t145 VGND 0.02304f
C11567 Iout.n53 VGND 0.05124f
C11568 Iout.n54 VGND 0.02606f
C11569 Iout.n55 VGND 0.23929f
C11570 Iout.t32 VGND 0.02304f
C11571 Iout.n56 VGND 0.05124f
C11572 Iout.n57 VGND 0.02606f
C11573 Iout.n58 VGND 0.23929f
C11574 Iout.t5 VGND 0.02304f
C11575 Iout.n59 VGND 0.05124f
C11576 Iout.n60 VGND 0.02606f
C11577 Iout.n61 VGND 0.23929f
C11578 Iout.t68 VGND 0.02304f
C11579 Iout.n62 VGND 0.05124f
C11580 Iout.n63 VGND 0.02606f
C11581 Iout.n64 VGND 0.23929f
C11582 Iout.t82 VGND 0.02304f
C11583 Iout.n65 VGND 0.05124f
C11584 Iout.n66 VGND 0.02606f
C11585 Iout.n67 VGND 0.23929f
C11586 Iout.t242 VGND 0.02304f
C11587 Iout.n68 VGND 0.05124f
C11588 Iout.n69 VGND 0.02606f
C11589 Iout.n70 VGND 0.23929f
C11590 Iout.t136 VGND 0.02304f
C11591 Iout.n71 VGND 0.05124f
C11592 Iout.n72 VGND 0.02606f
C11593 Iout.n73 VGND 0.23929f
C11594 Iout.t223 VGND 0.02304f
C11595 Iout.n74 VGND 0.05124f
C11596 Iout.n75 VGND 0.02606f
C11597 Iout.n76 VGND 0.23929f
C11598 Iout.t128 VGND 0.02304f
C11599 Iout.n77 VGND 0.05124f
C11600 Iout.n78 VGND 0.02606f
C11601 Iout.n79 VGND 0.23929f
C11602 Iout.n80 VGND 0.23929f
C11603 Iout.t110 VGND 0.02304f
C11604 Iout.n81 VGND 0.05124f
C11605 Iout.n82 VGND 0.02606f
C11606 Iout.n83 VGND 0.23929f
C11607 Iout.n84 VGND 0.04775f
C11608 Iout.t60 VGND 0.02304f
C11609 Iout.n85 VGND 0.05124f
C11610 Iout.n86 VGND 0.02606f
C11611 Iout.t138 VGND 0.02304f
C11612 Iout.n87 VGND 0.05124f
C11613 Iout.n88 VGND 0.02606f
C11614 Iout.n89 VGND 0.23929f
C11615 Iout.t254 VGND 0.02304f
C11616 Iout.n90 VGND 0.05124f
C11617 Iout.n91 VGND 0.02606f
C11618 Iout.n92 VGND 0.23929f
C11619 Iout.t42 VGND 0.02304f
C11620 Iout.n93 VGND 0.05124f
C11621 Iout.n94 VGND 0.02606f
C11622 Iout.n95 VGND 0.23929f
C11623 Iout.t1 VGND 0.02304f
C11624 Iout.n96 VGND 0.05124f
C11625 Iout.n97 VGND 0.02606f
C11626 Iout.n98 VGND 0.23929f
C11627 Iout.t246 VGND 0.02304f
C11628 Iout.n99 VGND 0.05124f
C11629 Iout.n100 VGND 0.02606f
C11630 Iout.n101 VGND 0.23929f
C11631 Iout.t240 VGND 0.02304f
C11632 Iout.n102 VGND 0.05124f
C11633 Iout.n103 VGND 0.02606f
C11634 Iout.n104 VGND 0.23929f
C11635 Iout.t251 VGND 0.02304f
C11636 Iout.n105 VGND 0.05124f
C11637 Iout.n106 VGND 0.02606f
C11638 Iout.n107 VGND 0.23929f
C11639 Iout.t9 VGND 0.02304f
C11640 Iout.n108 VGND 0.05124f
C11641 Iout.n109 VGND 0.02606f
C11642 Iout.n110 VGND 0.23929f
C11643 Iout.t105 VGND 0.02304f
C11644 Iout.n111 VGND 0.05124f
C11645 Iout.n112 VGND 0.02606f
C11646 Iout.n113 VGND 0.23929f
C11647 Iout.t133 VGND 0.02304f
C11648 Iout.n114 VGND 0.05124f
C11649 Iout.n115 VGND 0.02606f
C11650 Iout.n116 VGND 0.23929f
C11651 Iout.t124 VGND 0.02304f
C11652 Iout.n117 VGND 0.05124f
C11653 Iout.n118 VGND 0.02606f
C11654 Iout.n119 VGND 0.23929f
C11655 Iout.t21 VGND 0.02304f
C11656 Iout.n120 VGND 0.05124f
C11657 Iout.n121 VGND 0.02606f
C11658 Iout.n122 VGND 0.04775f
C11659 Iout.t96 VGND 0.02304f
C11660 Iout.n123 VGND 0.05124f
C11661 Iout.n124 VGND 0.02606f
C11662 Iout.n125 VGND 0.23929f
C11663 Iout.n126 VGND 0.23929f
C11664 Iout.t160 VGND 0.02304f
C11665 Iout.n127 VGND 0.05124f
C11666 Iout.n128 VGND 0.02606f
C11667 Iout.n129 VGND 0.04775f
C11668 Iout.t87 VGND 0.02304f
C11669 Iout.n130 VGND 0.05124f
C11670 Iout.n131 VGND 0.02606f
C11671 Iout.n132 VGND 0.23929f
C11672 Iout.t113 VGND 0.02304f
C11673 Iout.n133 VGND 0.05124f
C11674 Iout.n134 VGND 0.02606f
C11675 Iout.n135 VGND 0.04775f
C11676 Iout.t91 VGND 0.02304f
C11677 Iout.n136 VGND 0.05124f
C11678 Iout.n137 VGND 0.02606f
C11679 Iout.n138 VGND 0.23929f
C11680 Iout.n139 VGND 0.23929f
C11681 Iout.t86 VGND 0.02304f
C11682 Iout.n140 VGND 0.05124f
C11683 Iout.n141 VGND 0.02606f
C11684 Iout.n142 VGND 0.04775f
C11685 Iout.t239 VGND 0.02304f
C11686 Iout.n143 VGND 0.05124f
C11687 Iout.n144 VGND 0.02606f
C11688 Iout.n145 VGND 0.14126f
C11689 Iout.t227 VGND 0.02304f
C11690 Iout.n146 VGND 0.05124f
C11691 Iout.n147 VGND 0.02606f
C11692 Iout.n148 VGND 0.04775f
C11693 Iout.t228 VGND 0.02304f
C11694 Iout.n149 VGND 0.05124f
C11695 Iout.n150 VGND 0.02606f
C11696 Iout.n151 VGND 0.23929f
C11697 Iout.n152 VGND 0.14126f
C11698 Iout.n153 VGND 0.23929f
C11699 Iout.n154 VGND 0.23929f
C11700 Iout.n155 VGND 0.23929f
C11701 Iout.t220 VGND 0.02304f
C11702 Iout.n156 VGND 0.05124f
C11703 Iout.n157 VGND 0.02606f
C11704 Iout.n158 VGND 0.23929f
C11705 Iout.n159 VGND 0.23929f
C11706 Iout.n160 VGND 0.23929f
C11707 Iout.n161 VGND 0.23929f
C11708 Iout.n162 VGND 0.23929f
C11709 Iout.n163 VGND 0.23929f
C11710 Iout.n164 VGND 0.23929f
C11711 Iout.n165 VGND 0.23929f
C11712 Iout.n166 VGND 0.23929f
C11713 Iout.n167 VGND 0.23929f
C11714 Iout.t203 VGND 0.02304f
C11715 Iout.n168 VGND 0.05124f
C11716 Iout.n169 VGND 0.02606f
C11717 Iout.n170 VGND 0.23929f
C11718 Iout.n171 VGND 0.04775f
C11719 Iout.t183 VGND 0.02304f
C11720 Iout.n172 VGND 0.05124f
C11721 Iout.n173 VGND 0.02606f
C11722 Iout.t4 VGND 0.02304f
C11723 Iout.n174 VGND 0.05124f
C11724 Iout.n175 VGND 0.02606f
C11725 Iout.n176 VGND 0.23929f
C11726 Iout.t78 VGND 0.02304f
C11727 Iout.n177 VGND 0.05124f
C11728 Iout.n178 VGND 0.02606f
C11729 Iout.n179 VGND 0.23929f
C11730 Iout.t43 VGND 0.02304f
C11731 Iout.n180 VGND 0.05124f
C11732 Iout.n181 VGND 0.02606f
C11733 Iout.n182 VGND 0.23929f
C11734 Iout.t174 VGND 0.02304f
C11735 Iout.n183 VGND 0.05124f
C11736 Iout.n184 VGND 0.02606f
C11737 Iout.n185 VGND 0.23929f
C11738 Iout.t19 VGND 0.02304f
C11739 Iout.n186 VGND 0.05124f
C11740 Iout.n187 VGND 0.02606f
C11741 Iout.n188 VGND 0.23929f
C11742 Iout.t255 VGND 0.02304f
C11743 Iout.n189 VGND 0.05124f
C11744 Iout.n190 VGND 0.02606f
C11745 Iout.n191 VGND 0.14126f
C11746 Iout.t157 VGND 0.02304f
C11747 Iout.n192 VGND 0.05124f
C11748 Iout.n193 VGND 0.02606f
C11749 Iout.n194 VGND 0.04775f
C11750 Iout.t253 VGND 0.02304f
C11751 Iout.n195 VGND 0.05124f
C11752 Iout.n196 VGND 0.02606f
C11753 Iout.n197 VGND 0.14126f
C11754 Iout.n198 VGND 0.04775f
C11755 Iout.t140 VGND 0.02304f
C11756 Iout.n199 VGND 0.05124f
C11757 Iout.n200 VGND 0.02606f
C11758 Iout.n201 VGND 0.04775f
C11759 Iout.t231 VGND 0.02304f
C11760 Iout.n202 VGND 0.05124f
C11761 Iout.n203 VGND 0.02606f
C11762 Iout.n204 VGND 0.14126f
C11763 Iout.n205 VGND 0.04775f
C11764 Iout.t194 VGND 0.02304f
C11765 Iout.n206 VGND 0.05124f
C11766 Iout.n207 VGND 0.02606f
C11767 Iout.n208 VGND 0.14126f
C11768 Iout.n209 VGND 0.04775f
C11769 Iout.t83 VGND 0.02304f
C11770 Iout.n210 VGND 0.05124f
C11771 Iout.n211 VGND 0.02606f
C11772 Iout.n212 VGND 0.14126f
C11773 Iout.n213 VGND 0.04775f
C11774 Iout.t90 VGND 0.02304f
C11775 Iout.n214 VGND 0.05124f
C11776 Iout.n215 VGND 0.02606f
C11777 Iout.n216 VGND 0.14126f
C11778 Iout.n217 VGND 0.04775f
C11779 Iout.t33 VGND 0.02304f
C11780 Iout.n218 VGND 0.05124f
C11781 Iout.n219 VGND 0.02606f
C11782 Iout.n220 VGND 0.14126f
C11783 Iout.n221 VGND 0.04775f
C11784 Iout.t206 VGND 0.02304f
C11785 Iout.n222 VGND 0.05124f
C11786 Iout.n223 VGND 0.02606f
C11787 Iout.n224 VGND 0.14126f
C11788 Iout.n225 VGND 0.04775f
C11789 Iout.t208 VGND 0.02304f
C11790 Iout.n226 VGND 0.05124f
C11791 Iout.n227 VGND 0.02606f
C11792 Iout.n228 VGND 0.04775f
C11793 Iout.n229 VGND 0.14126f
C11794 Iout.n230 VGND 0.23929f
C11795 Iout.n231 VGND 0.04775f
C11796 Iout.t159 VGND 0.02304f
C11797 Iout.n232 VGND 0.05124f
C11798 Iout.n233 VGND 0.02606f
C11799 Iout.n234 VGND 0.04775f
C11800 Iout.t114 VGND 0.02304f
C11801 Iout.n235 VGND 0.05124f
C11802 Iout.n236 VGND 0.02606f
C11803 Iout.n237 VGND 0.04775f
C11804 Iout.t143 VGND 0.02304f
C11805 Iout.n238 VGND 0.05124f
C11806 Iout.n239 VGND 0.02606f
C11807 Iout.n240 VGND 0.04775f
C11808 Iout.t18 VGND 0.02304f
C11809 Iout.n241 VGND 0.05124f
C11810 Iout.n242 VGND 0.02606f
C11811 Iout.n243 VGND 0.04775f
C11812 Iout.t131 VGND 0.02304f
C11813 Iout.n244 VGND 0.05124f
C11814 Iout.n245 VGND 0.02606f
C11815 Iout.n246 VGND 0.04775f
C11816 Iout.t215 VGND 0.02304f
C11817 Iout.n247 VGND 0.05124f
C11818 Iout.n248 VGND 0.02606f
C11819 Iout.n249 VGND 0.04775f
C11820 Iout.t173 VGND 0.02304f
C11821 Iout.n250 VGND 0.05124f
C11822 Iout.n251 VGND 0.02606f
C11823 Iout.t29 VGND 0.02304f
C11824 Iout.n252 VGND 0.05124f
C11825 Iout.n253 VGND 0.02606f
C11826 Iout.n254 VGND 0.04775f
C11827 Iout.t47 VGND 0.02304f
C11828 Iout.n255 VGND 0.05124f
C11829 Iout.n256 VGND 0.02606f
C11830 Iout.n257 VGND 0.04775f
C11831 Iout.n258 VGND 0.23929f
C11832 Iout.t134 VGND 0.02304f
C11833 Iout.n259 VGND 0.05124f
C11834 Iout.n260 VGND 0.02606f
C11835 Iout.n261 VGND 0.04775f
C11836 Iout.n262 VGND 0.23929f
C11837 Iout.n263 VGND 0.23929f
C11838 Iout.n264 VGND 0.04775f
C11839 Iout.t117 VGND 0.02304f
C11840 Iout.n265 VGND 0.05124f
C11841 Iout.n266 VGND 0.02606f
C11842 Iout.n267 VGND 0.04775f
C11843 Iout.n268 VGND 0.23929f
C11844 Iout.n269 VGND 0.23929f
C11845 Iout.n270 VGND 0.04775f
C11846 Iout.t45 VGND 0.02304f
C11847 Iout.n271 VGND 0.05124f
C11848 Iout.n272 VGND 0.02606f
C11849 Iout.n273 VGND 0.04775f
C11850 Iout.n274 VGND 0.23929f
C11851 Iout.n275 VGND 0.23929f
C11852 Iout.n276 VGND 0.04775f
C11853 Iout.t195 VGND 0.02304f
C11854 Iout.n277 VGND 0.05124f
C11855 Iout.n278 VGND 0.02606f
C11856 Iout.n279 VGND 0.04775f
C11857 Iout.n280 VGND 0.23929f
C11858 Iout.n281 VGND 0.23929f
C11859 Iout.n282 VGND 0.04775f
C11860 Iout.t101 VGND 0.02304f
C11861 Iout.n283 VGND 0.05124f
C11862 Iout.n284 VGND 0.02606f
C11863 Iout.n285 VGND 0.04775f
C11864 Iout.n286 VGND 0.23929f
C11865 Iout.n287 VGND 0.23929f
C11866 Iout.n288 VGND 0.04775f
C11867 Iout.t74 VGND 0.02304f
C11868 Iout.n289 VGND 0.05124f
C11869 Iout.n290 VGND 0.02606f
C11870 Iout.n291 VGND 0.04775f
C11871 Iout.n292 VGND 0.23929f
C11872 Iout.n293 VGND 0.23929f
C11873 Iout.n294 VGND 0.04775f
C11874 Iout.t66 VGND 0.02304f
C11875 Iout.n295 VGND 0.05124f
C11876 Iout.n296 VGND 0.02606f
C11877 Iout.n297 VGND 0.04775f
C11878 Iout.n298 VGND 0.23929f
C11879 Iout.n299 VGND 0.23929f
C11880 Iout.n300 VGND 0.04775f
C11881 Iout.t153 VGND 0.02304f
C11882 Iout.n301 VGND 0.05124f
C11883 Iout.n302 VGND 0.02606f
C11884 Iout.n303 VGND 0.04775f
C11885 Iout.n304 VGND 0.23929f
C11886 Iout.t181 VGND 0.02304f
C11887 Iout.n305 VGND 0.05124f
C11888 Iout.n306 VGND 0.02606f
C11889 Iout.n307 VGND 0.04775f
C11890 Iout.t237 VGND 0.02304f
C11891 Iout.n308 VGND 0.05124f
C11892 Iout.n309 VGND 0.02606f
C11893 Iout.n310 VGND 0.04775f
C11894 Iout.t154 VGND 0.02304f
C11895 Iout.n311 VGND 0.05124f
C11896 Iout.n312 VGND 0.02606f
C11897 Iout.n313 VGND 0.04775f
C11898 Iout.t10 VGND 0.02304f
C11899 Iout.n314 VGND 0.05124f
C11900 Iout.n315 VGND 0.02606f
C11901 Iout.n316 VGND 0.04775f
C11902 Iout.t250 VGND 0.02304f
C11903 Iout.n317 VGND 0.05124f
C11904 Iout.n318 VGND 0.02606f
C11905 Iout.n319 VGND 0.04775f
C11906 Iout.t7 VGND 0.02304f
C11907 Iout.n320 VGND 0.05124f
C11908 Iout.n321 VGND 0.02606f
C11909 Iout.n322 VGND 0.04775f
C11910 Iout.t212 VGND 0.02304f
C11911 Iout.n323 VGND 0.05124f
C11912 Iout.n324 VGND 0.02606f
C11913 Iout.n325 VGND 0.04775f
C11914 Iout.t229 VGND 0.02304f
C11915 Iout.n326 VGND 0.05124f
C11916 Iout.n327 VGND 0.02606f
C11917 Iout.n328 VGND 0.04775f
C11918 Iout.t193 VGND 0.02304f
C11919 Iout.n329 VGND 0.05124f
C11920 Iout.n330 VGND 0.02606f
C11921 Iout.n331 VGND 0.04775f
C11922 Iout.n332 VGND 0.23929f
C11923 Iout.t234 VGND 0.02304f
C11924 Iout.n333 VGND 0.05124f
C11925 Iout.n334 VGND 0.02606f
C11926 Iout.n335 VGND 0.04775f
C11927 Iout.t17 VGND 0.02304f
C11928 Iout.n336 VGND 0.05124f
C11929 Iout.n337 VGND 0.02606f
C11930 Iout.n338 VGND 0.04775f
C11931 Iout.t230 VGND 0.02304f
C11932 Iout.n339 VGND 0.05124f
C11933 Iout.n340 VGND 0.02606f
C11934 Iout.n341 VGND 0.04775f
C11935 Iout.t205 VGND 0.02304f
C11936 Iout.n342 VGND 0.05124f
C11937 Iout.n343 VGND 0.02606f
C11938 Iout.n344 VGND 0.04775f
C11939 Iout.t210 VGND 0.02304f
C11940 Iout.n345 VGND 0.05124f
C11941 Iout.n346 VGND 0.02606f
C11942 Iout.n347 VGND 0.04775f
C11943 Iout.t213 VGND 0.02304f
C11944 Iout.n348 VGND 0.05124f
C11945 Iout.n349 VGND 0.02606f
C11946 Iout.n350 VGND 0.04775f
C11947 Iout.t13 VGND 0.02304f
C11948 Iout.n351 VGND 0.05124f
C11949 Iout.n352 VGND 0.02606f
C11950 Iout.n353 VGND 0.04775f
C11951 Iout.t209 VGND 0.02304f
C11952 Iout.n354 VGND 0.05124f
C11953 Iout.n355 VGND 0.02606f
C11954 Iout.n356 VGND 0.04775f
C11955 Iout.t107 VGND 0.02304f
C11956 Iout.n357 VGND 0.05124f
C11957 Iout.n358 VGND 0.02606f
C11958 Iout.n359 VGND 0.04775f
C11959 Iout.t147 VGND 0.02304f
C11960 Iout.n360 VGND 0.05124f
C11961 Iout.n361 VGND 0.02606f
C11962 Iout.n362 VGND 0.04775f
C11963 Iout.t31 VGND 0.02304f
C11964 Iout.n363 VGND 0.05124f
C11965 Iout.n364 VGND 0.02606f
C11966 Iout.n365 VGND 0.04775f
C11967 Iout.t226 VGND 0.02304f
C11968 Iout.n366 VGND 0.05124f
C11969 Iout.n367 VGND 0.02606f
C11970 Iout.n368 VGND 0.04775f
C11971 Iout.n369 VGND 0.23929f
C11972 Iout.t139 VGND 0.02304f
C11973 Iout.n370 VGND 0.05124f
C11974 Iout.n371 VGND 0.02606f
C11975 Iout.n372 VGND 0.04775f
C11976 Iout.n373 VGND 0.23929f
C11977 Iout.n374 VGND 0.23929f
C11978 Iout.n375 VGND 0.04775f
C11979 Iout.t121 VGND 0.02304f
C11980 Iout.n376 VGND 0.05124f
C11981 Iout.n377 VGND 0.02606f
C11982 Iout.t12 VGND 0.02304f
C11983 Iout.n378 VGND 0.05124f
C11984 Iout.n379 VGND 0.02606f
C11985 Iout.n380 VGND 0.04775f
C11986 Iout.n381 VGND 0.23929f
C11987 Iout.n382 VGND 0.23929f
C11988 Iout.n383 VGND 0.04775f
C11989 Iout.t24 VGND 0.02304f
C11990 Iout.n384 VGND 0.05124f
C11991 Iout.n385 VGND 0.02606f
C11992 Iout.t99 VGND 0.02304f
C11993 Iout.n386 VGND 0.05124f
C11994 Iout.n387 VGND 0.02606f
C11995 Iout.n388 VGND 0.04775f
C11996 Iout.n389 VGND 0.23929f
C11997 Iout.n390 VGND 0.23929f
C11998 Iout.n391 VGND 0.04775f
C11999 Iout.t152 VGND 0.02304f
C12000 Iout.n392 VGND 0.05124f
C12001 Iout.n393 VGND 0.02606f
C12002 Iout.t165 VGND 0.02304f
C12003 Iout.n394 VGND 0.05124f
C12004 Iout.n395 VGND 0.02606f
C12005 Iout.n396 VGND 0.04775f
C12006 Iout.n397 VGND 0.23929f
C12007 Iout.n398 VGND 0.23929f
C12008 Iout.n399 VGND 0.04775f
C12009 Iout.t50 VGND 0.02304f
C12010 Iout.n400 VGND 0.05124f
C12011 Iout.n401 VGND 0.02606f
C12012 Iout.t172 VGND 0.02304f
C12013 Iout.n402 VGND 0.05124f
C12014 Iout.n403 VGND 0.02606f
C12015 Iout.n404 VGND 0.04775f
C12016 Iout.n405 VGND 0.23929f
C12017 Iout.n406 VGND 0.23929f
C12018 Iout.n407 VGND 0.04775f
C12019 Iout.t61 VGND 0.02304f
C12020 Iout.n408 VGND 0.05124f
C12021 Iout.n409 VGND 0.02606f
C12022 Iout.t199 VGND 0.02304f
C12023 Iout.n410 VGND 0.05124f
C12024 Iout.n411 VGND 0.02606f
C12025 Iout.n412 VGND 0.04775f
C12026 Iout.n413 VGND 0.23929f
C12027 Iout.n414 VGND 0.23929f
C12028 Iout.n415 VGND 0.04775f
C12029 Iout.t51 VGND 0.02304f
C12030 Iout.n416 VGND 0.05124f
C12031 Iout.n417 VGND 0.02606f
C12032 Iout.t198 VGND 0.02304f
C12033 Iout.n418 VGND 0.05124f
C12034 Iout.n419 VGND 0.02606f
C12035 Iout.n420 VGND 0.04775f
C12036 Iout.n421 VGND 0.23929f
C12037 Iout.n422 VGND 0.23929f
C12038 Iout.n423 VGND 0.04775f
C12039 Iout.t190 VGND 0.02304f
C12040 Iout.n424 VGND 0.05124f
C12041 Iout.n425 VGND 0.02606f
C12042 Iout.t88 VGND 0.02304f
C12043 Iout.n426 VGND 0.05124f
C12044 Iout.n427 VGND 0.02606f
C12045 Iout.n428 VGND 0.04775f
C12046 Iout.n429 VGND 0.23929f
C12047 Iout.n430 VGND 0.23929f
C12048 Iout.n431 VGND 0.04775f
C12049 Iout.t106 VGND 0.02304f
C12050 Iout.n432 VGND 0.05124f
C12051 Iout.n433 VGND 0.02606f
C12052 Iout.t155 VGND 0.02304f
C12053 Iout.n434 VGND 0.05124f
C12054 Iout.n435 VGND 0.02606f
C12055 Iout.n436 VGND 0.23929f
C12056 Iout.n437 VGND 0.04775f
C12057 Iout.t6 VGND 0.02304f
C12058 Iout.n438 VGND 0.05124f
C12059 Iout.n439 VGND 0.02606f
C12060 Iout.n440 VGND 0.04775f
C12061 Iout.t214 VGND 0.02304f
C12062 Iout.n441 VGND 0.05124f
C12063 Iout.n442 VGND 0.02606f
C12064 Iout.n443 VGND 0.04775f
C12065 Iout.n444 VGND 0.23929f
C12066 Iout.n445 VGND 0.23929f
C12067 Iout.n446 VGND 0.04775f
C12068 Iout.t232 VGND 0.02304f
C12069 Iout.n447 VGND 0.05124f
C12070 Iout.n448 VGND 0.02606f
C12071 Iout.t252 VGND 0.02304f
C12072 Iout.n449 VGND 0.05124f
C12073 Iout.n450 VGND 0.02606f
C12074 Iout.n451 VGND 0.04775f
C12075 Iout.t129 VGND 0.02304f
C12076 Iout.n452 VGND 0.05124f
C12077 Iout.n453 VGND 0.02606f
C12078 Iout.n454 VGND 0.04775f
C12079 Iout.n455 VGND 0.23929f
C12080 Iout.n456 VGND 0.23929f
C12081 Iout.n457 VGND 0.04775f
C12082 Iout.t27 VGND 0.02304f
C12083 Iout.n458 VGND 0.05124f
C12084 Iout.n459 VGND 0.02606f
C12085 Iout.t186 VGND 0.02304f
C12086 Iout.n460 VGND 0.05124f
C12087 Iout.n461 VGND 0.02606f
C12088 Iout.n462 VGND 0.04775f
C12089 Iout.t158 VGND 0.02304f
C12090 Iout.n463 VGND 0.05124f
C12091 Iout.n464 VGND 0.02606f
C12092 Iout.n465 VGND 0.04775f
C12093 Iout.n466 VGND 0.23929f
C12094 Iout.n467 VGND 0.23929f
C12095 Iout.n468 VGND 0.04775f
C12096 Iout.t166 VGND 0.02304f
C12097 Iout.n469 VGND 0.05124f
C12098 Iout.n470 VGND 0.02606f
C12099 Iout.n471 VGND 0.04775f
C12100 Iout.t201 VGND 0.02304f
C12101 Iout.n472 VGND 0.05124f
C12102 Iout.n473 VGND 0.02606f
C12103 Iout.n474 VGND 0.04775f
C12104 Iout.n475 VGND 0.23929f
C12105 Iout.n476 VGND 0.23929f
C12106 Iout.n477 VGND 0.04775f
C12107 Iout.t167 VGND 0.02304f
C12108 Iout.n478 VGND 0.05124f
C12109 Iout.n479 VGND 0.02606f
C12110 Iout.t58 VGND 0.02304f
C12111 Iout.n480 VGND 0.05124f
C12112 Iout.n481 VGND 0.02606f
C12113 Iout.n482 VGND 0.04775f
C12114 Iout.t243 VGND 0.02304f
C12115 Iout.n483 VGND 0.05124f
C12116 Iout.n484 VGND 0.02606f
C12117 Iout.n485 VGND 0.04775f
C12118 Iout.n486 VGND 0.23929f
C12119 Iout.n487 VGND 0.23929f
C12120 Iout.n488 VGND 0.04775f
C12121 Iout.t38 VGND 0.02304f
C12122 Iout.n489 VGND 0.05124f
C12123 Iout.n490 VGND 0.02606f
C12124 Iout.t55 VGND 0.02304f
C12125 Iout.n491 VGND 0.05124f
C12126 Iout.n492 VGND 0.02606f
C12127 Iout.n493 VGND 0.04775f
C12128 Iout.t34 VGND 0.02304f
C12129 Iout.n494 VGND 0.05124f
C12130 Iout.n495 VGND 0.02606f
C12131 Iout.n496 VGND 0.04775f
C12132 Iout.n497 VGND 0.23929f
C12133 Iout.n498 VGND 0.14126f
C12134 Iout.n499 VGND 0.04775f
C12135 Iout.t197 VGND 0.02304f
C12136 Iout.n500 VGND 0.05124f
C12137 Iout.n501 VGND 0.02606f
C12138 Iout.n502 VGND 0.14126f
C12139 Iout.n503 VGND 0.04775f
C12140 Iout.t241 VGND 0.02304f
C12141 Iout.n504 VGND 0.05124f
C12142 Iout.n505 VGND 0.02606f
C12143 Iout.n506 VGND 0.04775f
C12144 Iout.t112 VGND 0.02304f
C12145 Iout.n507 VGND 0.05124f
C12146 Iout.n508 VGND 0.02606f
C12147 Iout.t20 VGND 0.02304f
C12148 Iout.n509 VGND 0.05124f
C12149 Iout.n510 VGND 0.02606f
C12150 Iout.n511 VGND 0.14126f
C12151 Iout.n512 VGND 0.04775f
C12152 Iout.t65 VGND 0.02304f
C12153 Iout.n513 VGND 0.05124f
C12154 Iout.n514 VGND 0.02606f
C12155 Iout.n515 VGND 0.04775f
C12156 Iout.n516 VGND 0.14126f
C12157 Iout.n517 VGND 0.23929f
C12158 Iout.n518 VGND 0.04775f
C12159 Iout.t2 VGND 0.02304f
C12160 Iout.n519 VGND 0.05124f
C12161 Iout.n520 VGND 0.02606f
C12162 Iout.n521 VGND 0.04775f
C12163 Iout.n522 VGND 0.23929f
C12164 Iout.n523 VGND 0.23929f
C12165 Iout.n524 VGND 0.04775f
C12166 Iout.t130 VGND 0.02304f
C12167 Iout.n525 VGND 0.05124f
C12168 Iout.n526 VGND 0.02606f
C12169 Iout.n527 VGND 0.04775f
C12170 Iout.n528 VGND 0.23929f
C12171 Iout.n529 VGND 0.23929f
C12172 Iout.n530 VGND 0.04775f
C12173 Iout.t59 VGND 0.02304f
C12174 Iout.n531 VGND 0.05124f
C12175 Iout.n532 VGND 0.02606f
C12176 Iout.n533 VGND 0.04775f
C12177 Iout.t146 VGND 0.02304f
C12178 Iout.n534 VGND 0.05124f
C12179 Iout.n535 VGND 0.02606f
C12180 Iout.t75 VGND 0.02304f
C12181 Iout.n536 VGND 0.05124f
C12182 Iout.n537 VGND 0.02606f
C12183 Iout.n538 VGND 0.04775f
C12184 Iout.n539 VGND 0.23929f
C12185 Iout.n540 VGND 0.23929f
C12186 Iout.n541 VGND 0.04775f
C12187 Iout.t119 VGND 0.02304f
C12188 Iout.n542 VGND 0.05124f
C12189 Iout.n543 VGND 0.02606f
C12190 Iout.n544 VGND 0.04775f
C12191 Iout.n545 VGND 0.23929f
C12192 Iout.n546 VGND 0.23929f
C12193 Iout.n547 VGND 0.04775f
C12194 Iout.t122 VGND 0.02304f
C12195 Iout.n548 VGND 0.05124f
C12196 Iout.n549 VGND 0.02606f
C12197 Iout.n550 VGND 0.04775f
C12198 Iout.n551 VGND 0.23929f
C12199 Iout.n552 VGND 0.23929f
C12200 Iout.n553 VGND 0.04775f
C12201 Iout.t171 VGND 0.02304f
C12202 Iout.n554 VGND 0.05124f
C12203 Iout.n555 VGND 0.02606f
C12204 Iout.n556 VGND 0.04775f
C12205 Iout.t178 VGND 0.02304f
C12206 Iout.n557 VGND 0.05124f
C12207 Iout.n558 VGND 0.02606f
C12208 Iout.t14 VGND 0.02304f
C12209 Iout.n559 VGND 0.05124f
C12210 Iout.n560 VGND 0.02606f
C12211 Iout.n561 VGND 0.04775f
C12212 Iout.n562 VGND 0.23929f
C12213 Iout.t15 VGND 0.02304f
C12214 Iout.n563 VGND 0.05124f
C12215 Iout.n564 VGND 0.02606f
C12216 Iout.n565 VGND 0.04775f
C12217 Iout.n566 VGND 0.23929f
C12218 Iout.n567 VGND 0.23929f
C12219 Iout.n568 VGND 0.04775f
C12220 Iout.t79 VGND 0.02304f
C12221 Iout.n569 VGND 0.05124f
C12222 Iout.n570 VGND 0.02606f
C12223 Iout.n571 VGND 0.04775f
C12224 Iout.n572 VGND 0.23929f
C12225 Iout.t161 VGND 0.02304f
C12226 Iout.n573 VGND 0.05124f
C12227 Iout.n574 VGND 0.02606f
C12228 Iout.n575 VGND 0.04775f
C12229 Iout.t177 VGND 0.02304f
C12230 Iout.n576 VGND 0.05124f
C12231 Iout.n577 VGND 0.02606f
C12232 Iout.n578 VGND 0.04775f
C12233 Iout.n579 VGND 0.23929f
C12234 Iout.n580 VGND 0.23929f
C12235 Iout.n581 VGND 0.04775f
C12236 Iout.t222 VGND 0.02304f
C12237 Iout.n582 VGND 0.05124f
C12238 Iout.n583 VGND 0.02606f
C12239 Iout.n584 VGND 0.04775f
C12240 Iout.n585 VGND 0.23929f
C12241 Iout.n586 VGND 0.23929f
C12242 Iout.n587 VGND 0.04775f
C12243 Iout.t179 VGND 0.02304f
C12244 Iout.n588 VGND 0.05124f
C12245 Iout.n589 VGND 0.02606f
C12246 Iout.n590 VGND 0.04775f
C12247 Iout.n591 VGND 0.23929f
C12248 Iout.n592 VGND 0.23929f
C12249 Iout.n593 VGND 0.04775f
C12250 Iout.t175 VGND 0.02304f
C12251 Iout.n594 VGND 0.05124f
C12252 Iout.n595 VGND 0.02606f
C12253 Iout.n596 VGND 0.04775f
C12254 Iout.n597 VGND 0.23929f
C12255 Iout.n598 VGND 0.23929f
C12256 Iout.n599 VGND 0.04775f
C12257 Iout.t22 VGND 0.02304f
C12258 Iout.n600 VGND 0.05124f
C12259 Iout.n601 VGND 0.02606f
C12260 Iout.n602 VGND 0.04775f
C12261 Iout.n603 VGND 0.23929f
C12262 Iout.n604 VGND 0.23929f
C12263 Iout.n605 VGND 0.04775f
C12264 Iout.t39 VGND 0.02304f
C12265 Iout.n606 VGND 0.05124f
C12266 Iout.n607 VGND 0.02606f
C12267 Iout.n608 VGND 0.04775f
C12268 Iout.n609 VGND 0.23929f
C12269 Iout.n610 VGND 0.23929f
C12270 Iout.n611 VGND 0.04775f
C12271 Iout.t62 VGND 0.02304f
C12272 Iout.n612 VGND 0.05124f
C12273 Iout.n613 VGND 0.02606f
C12274 Iout.n614 VGND 0.04775f
C12275 Iout.n615 VGND 0.23929f
C12276 Iout.n616 VGND 0.23929f
C12277 Iout.n617 VGND 0.04775f
C12278 Iout.t132 VGND 0.02304f
C12279 Iout.n618 VGND 0.05124f
C12280 Iout.n619 VGND 0.02606f
C12281 Iout.n620 VGND 0.04775f
C12282 Iout.n621 VGND 0.23929f
C12283 Iout.n622 VGND 0.23929f
C12284 Iout.n623 VGND 0.04775f
C12285 Iout.t202 VGND 0.02304f
C12286 Iout.n624 VGND 0.05124f
C12287 Iout.n625 VGND 0.02606f
C12288 Iout.n626 VGND 0.04775f
C12289 Iout.n627 VGND 0.23929f
C12290 Iout.n628 VGND 0.23929f
C12291 Iout.n629 VGND 0.04775f
C12292 Iout.t84 VGND 0.02304f
C12293 Iout.n630 VGND 0.05124f
C12294 Iout.n631 VGND 0.02606f
C12295 Iout.n632 VGND 0.04775f
C12296 Iout.n633 VGND 0.23929f
C12297 Iout.n634 VGND 0.23929f
C12298 Iout.n635 VGND 0.04775f
C12299 Iout.t64 VGND 0.02304f
C12300 Iout.n636 VGND 0.05124f
C12301 Iout.n637 VGND 0.02606f
C12302 Iout.n638 VGND 0.04775f
C12303 Iout.n639 VGND 0.23929f
C12304 Iout.n640 VGND 0.23929f
C12305 Iout.n641 VGND 0.04775f
C12306 Iout.t120 VGND 0.02304f
C12307 Iout.n642 VGND 0.05124f
C12308 Iout.n643 VGND 0.02606f
C12309 Iout.n644 VGND 0.04775f
C12310 Iout.n645 VGND 0.23929f
C12311 Iout.n646 VGND 0.23929f
C12312 Iout.n647 VGND 0.04775f
C12313 Iout.t71 VGND 0.02304f
C12314 Iout.n648 VGND 0.05124f
C12315 Iout.n649 VGND 0.02606f
C12316 Iout.n650 VGND 0.04775f
C12317 Iout.n651 VGND 0.23929f
C12318 Iout.n652 VGND 0.23929f
C12319 Iout.n653 VGND 0.04775f
C12320 Iout.t180 VGND 0.02304f
C12321 Iout.n654 VGND 0.05124f
C12322 Iout.n655 VGND 0.02606f
C12323 Iout.n656 VGND 0.04775f
C12324 Iout.t245 VGND 0.02304f
C12325 Iout.n657 VGND 0.05124f
C12326 Iout.n658 VGND 0.02606f
C12327 Iout.n659 VGND 0.04775f
C12328 Iout.t35 VGND 0.02304f
C12329 Iout.n660 VGND 0.05124f
C12330 Iout.n661 VGND 0.02606f
C12331 Iout.n662 VGND 0.04775f
C12332 Iout.t3 VGND 0.02304f
C12333 Iout.n663 VGND 0.05124f
C12334 Iout.n664 VGND 0.02606f
C12335 Iout.n665 VGND 0.04775f
C12336 Iout.t163 VGND 0.02304f
C12337 Iout.n666 VGND 0.05124f
C12338 Iout.n667 VGND 0.02606f
C12339 Iout.n668 VGND 0.04775f
C12340 Iout.t141 VGND 0.02304f
C12341 Iout.n669 VGND 0.05124f
C12342 Iout.n670 VGND 0.02606f
C12343 Iout.n671 VGND 0.04775f
C12344 Iout.t185 VGND 0.02304f
C12345 Iout.n672 VGND 0.05124f
C12346 Iout.n673 VGND 0.02606f
C12347 Iout.n674 VGND 0.04775f
C12348 Iout.t94 VGND 0.02304f
C12349 Iout.n675 VGND 0.05124f
C12350 Iout.n676 VGND 0.02606f
C12351 Iout.n677 VGND 0.04775f
C12352 Iout.t40 VGND 0.02304f
C12353 Iout.n678 VGND 0.05124f
C12354 Iout.n679 VGND 0.02606f
C12355 Iout.n680 VGND 0.04775f
C12356 Iout.t247 VGND 0.02304f
C12357 Iout.n681 VGND 0.05124f
C12358 Iout.n682 VGND 0.02606f
C12359 Iout.n683 VGND 0.04775f
C12360 Iout.t116 VGND 0.02304f
C12361 Iout.n684 VGND 0.05124f
C12362 Iout.n685 VGND 0.02606f
C12363 Iout.n686 VGND 0.04775f
C12364 Iout.t170 VGND 0.02304f
C12365 Iout.n687 VGND 0.05124f
C12366 Iout.n688 VGND 0.02606f
C12367 Iout.n689 VGND 0.04775f
C12368 Iout.t97 VGND 0.02304f
C12369 Iout.n690 VGND 0.05124f
C12370 Iout.n691 VGND 0.02606f
C12371 Iout.t225 VGND 0.02304f
C12372 Iout.n692 VGND 0.05124f
C12373 Iout.n693 VGND 0.02606f
C12374 Iout.n694 VGND 0.04775f
C12375 Iout.t54 VGND 0.02304f
C12376 Iout.n695 VGND 0.05124f
C12377 Iout.n696 VGND 0.02606f
C12378 Iout.n697 VGND 0.04775f
C12379 Iout.n698 VGND 0.23929f
C12380 Iout.t26 VGND 0.02304f
C12381 Iout.n699 VGND 0.05124f
C12382 Iout.n700 VGND 0.02606f
C12383 Iout.n701 VGND 0.04775f
C12384 Iout.n702 VGND 0.23929f
C12385 Iout.n703 VGND 0.23929f
C12386 Iout.n704 VGND 0.04775f
C12387 Iout.t11 VGND 0.02304f
C12388 Iout.n705 VGND 0.05124f
C12389 Iout.n706 VGND 0.02606f
C12390 Iout.n707 VGND 0.04775f
C12391 Iout.n708 VGND 0.23929f
C12392 Iout.n709 VGND 0.23929f
C12393 Iout.n710 VGND 0.04775f
C12394 Iout.t233 VGND 0.02304f
C12395 Iout.n711 VGND 0.05124f
C12396 Iout.n712 VGND 0.02606f
C12397 Iout.n713 VGND 0.04775f
C12398 Iout.n714 VGND 0.23929f
C12399 Iout.n715 VGND 0.23929f
C12400 Iout.n716 VGND 0.04775f
C12401 Iout.t125 VGND 0.02304f
C12402 Iout.n717 VGND 0.05124f
C12403 Iout.n718 VGND 0.02606f
C12404 Iout.n719 VGND 0.04775f
C12405 Iout.n720 VGND 0.23929f
C12406 Iout.n721 VGND 0.23929f
C12407 Iout.n722 VGND 0.04775f
C12408 Iout.t109 VGND 0.02304f
C12409 Iout.n723 VGND 0.05124f
C12410 Iout.n724 VGND 0.02606f
C12411 Iout.n725 VGND 0.04775f
C12412 Iout.n726 VGND 0.23929f
C12413 Iout.n727 VGND 0.23929f
C12414 Iout.n728 VGND 0.04775f
C12415 Iout.t169 VGND 0.02304f
C12416 Iout.n729 VGND 0.05124f
C12417 Iout.n730 VGND 0.02606f
C12418 Iout.n731 VGND 0.04775f
C12419 Iout.n732 VGND 0.23929f
C12420 Iout.n733 VGND 0.23929f
C12421 Iout.n734 VGND 0.04775f
C12422 Iout.t200 VGND 0.02304f
C12423 Iout.n735 VGND 0.05124f
C12424 Iout.n736 VGND 0.02606f
C12425 Iout.n737 VGND 0.04775f
C12426 Iout.n738 VGND 0.23929f
C12427 Iout.n739 VGND 0.23929f
C12428 Iout.n740 VGND 0.04775f
C12429 Iout.t63 VGND 0.02304f
C12430 Iout.n741 VGND 0.05124f
C12431 Iout.n742 VGND 0.02606f
C12432 Iout.n743 VGND 0.04775f
C12433 Iout.n744 VGND 0.23929f
C12434 Iout.n745 VGND 0.23929f
C12435 Iout.n746 VGND 0.04775f
C12436 Iout.t53 VGND 0.02304f
C12437 Iout.n747 VGND 0.05124f
C12438 Iout.n748 VGND 0.02606f
C12439 Iout.n749 VGND 0.04775f
C12440 Iout.n750 VGND 0.23929f
C12441 Iout.n751 VGND 0.23929f
C12442 Iout.n752 VGND 0.04775f
C12443 Iout.t98 VGND 0.02304f
C12444 Iout.n753 VGND 0.05124f
C12445 Iout.n754 VGND 0.02606f
C12446 Iout.n755 VGND 0.04775f
C12447 Iout.n756 VGND 0.23929f
C12448 Iout.n757 VGND 0.23929f
C12449 Iout.n758 VGND 0.04775f
C12450 Iout.t126 VGND 0.02304f
C12451 Iout.n759 VGND 0.05124f
C12452 Iout.n760 VGND 0.02606f
C12453 Iout.n761 VGND 0.04775f
C12454 Iout.n762 VGND 0.23929f
C12455 Iout.n763 VGND 0.23929f
C12456 Iout.n764 VGND 0.04775f
C12457 Iout.t127 VGND 0.02304f
C12458 Iout.n765 VGND 0.05124f
C12459 Iout.n766 VGND 0.02606f
C12460 Iout.n767 VGND 0.04775f
C12461 Iout.n768 VGND 0.23929f
C12462 Iout.n769 VGND 0.23929f
C12463 Iout.n770 VGND 0.04775f
C12464 Iout.t69 VGND 0.02304f
C12465 Iout.n771 VGND 0.05124f
C12466 Iout.n772 VGND 0.02606f
C12467 Iout.n773 VGND 0.04775f
C12468 Iout.n774 VGND 0.23929f
C12469 Iout.n775 VGND 0.23929f
C12470 Iout.n776 VGND 0.04775f
C12471 Iout.t81 VGND 0.02304f
C12472 Iout.n777 VGND 0.05124f
C12473 Iout.n778 VGND 0.02606f
C12474 Iout.n779 VGND 0.04775f
C12475 Iout.n780 VGND 0.23929f
C12476 Iout.t235 VGND 0.02304f
C12477 Iout.n781 VGND 0.05124f
C12478 Iout.n782 VGND 0.02606f
C12479 Iout.n783 VGND 0.04775f
C12480 Iout.t221 VGND 0.02304f
C12481 Iout.n784 VGND 0.05124f
C12482 Iout.n785 VGND 0.02606f
C12483 Iout.n786 VGND 0.04775f
C12484 Iout.t28 VGND 0.02304f
C12485 Iout.n787 VGND 0.05124f
C12486 Iout.n788 VGND 0.02606f
C12487 Iout.n789 VGND 0.04775f
C12488 Iout.t144 VGND 0.02304f
C12489 Iout.n790 VGND 0.05124f
C12490 Iout.n791 VGND 0.02606f
C12491 Iout.n792 VGND 0.04775f
C12492 Iout.t111 VGND 0.02304f
C12493 Iout.n793 VGND 0.05124f
C12494 Iout.n794 VGND 0.02606f
C12495 Iout.n795 VGND 0.04775f
C12496 Iout.t77 VGND 0.02304f
C12497 Iout.n796 VGND 0.05124f
C12498 Iout.n797 VGND 0.02606f
C12499 Iout.n798 VGND 0.04775f
C12500 Iout.t23 VGND 0.02304f
C12501 Iout.n799 VGND 0.05124f
C12502 Iout.n800 VGND 0.02606f
C12503 Iout.n801 VGND 0.04775f
C12504 Iout.t238 VGND 0.02304f
C12505 Iout.n802 VGND 0.05124f
C12506 Iout.n803 VGND 0.02606f
C12507 Iout.n804 VGND 0.04775f
C12508 Iout.t123 VGND 0.02304f
C12509 Iout.n805 VGND 0.05124f
C12510 Iout.n806 VGND 0.02606f
C12511 Iout.n807 VGND 0.04775f
C12512 Iout.t80 VGND 0.02304f
C12513 Iout.n808 VGND 0.05124f
C12514 Iout.n809 VGND 0.02606f
C12515 Iout.n810 VGND 0.04775f
C12516 Iout.t70 VGND 0.02304f
C12517 Iout.n811 VGND 0.05124f
C12518 Iout.n812 VGND 0.02606f
C12519 Iout.n813 VGND 0.04775f
C12520 Iout.t8 VGND 0.02304f
C12521 Iout.n814 VGND 0.05124f
C12522 Iout.n815 VGND 0.02606f
C12523 Iout.n816 VGND 0.04775f
C12524 Iout.t211 VGND 0.02304f
C12525 Iout.n817 VGND 0.05124f
C12526 Iout.n818 VGND 0.02606f
C12527 Iout.n819 VGND 0.04775f
C12528 Iout.t36 VGND 0.02304f
C12529 Iout.n820 VGND 0.05124f
C12530 Iout.n821 VGND 0.02606f
C12531 Iout.n822 VGND 0.04775f
C12532 Iout.t156 VGND 0.02304f
C12533 Iout.n823 VGND 0.05124f
C12534 Iout.n824 VGND 0.02606f
C12535 Iout.n825 VGND 0.04775f
C12536 Iout.n826 VGND 0.23929f
C12537 Iout.t176 VGND 0.02304f
C12538 Iout.n827 VGND 0.05124f
C12539 Iout.n828 VGND 0.02606f
C12540 Iout.n829 VGND 0.08168f
C12541 Iout.n830 VGND 0.49611f
C12542 Iout.n831 VGND 0.04775f
C12543 Iout.t52 VGND 0.02304f
C12544 Iout.n832 VGND 0.05124f
C12545 Iout.n833 VGND 0.02606f
C12546 Iout.t25 VGND 0.02304f
C12547 Iout.n834 VGND 0.05124f
C12548 Iout.n835 VGND 0.02606f
C12549 Iout.n836 VGND 0.04775f
C12550 Iout.n837 VGND 0.49611f
C12551 Iout.n838 VGND 0.08168f
C12552 Iout.t46 VGND 0.02304f
C12553 Iout.n839 VGND 0.05124f
C12554 Iout.n840 VGND 0.02606f
C12555 Iout.t41 VGND 0.02304f
C12556 Iout.n841 VGND 0.05124f
C12557 Iout.n842 VGND 0.02606f
C12558 Iout.n843 VGND 0.08168f
C12559 Iout.n844 VGND 0.49611f
C12560 Iout.n845 VGND 0.04775f
C12561 Iout.t151 VGND 0.02304f
C12562 Iout.n846 VGND 0.05124f
C12563 Iout.n847 VGND 0.02606f
C12564 Iout.t236 VGND 0.02304f
C12565 Iout.n848 VGND 0.05124f
C12566 Iout.n849 VGND 0.02606f
C12567 Iout.n850 VGND 0.04775f
C12568 Iout.n851 VGND 0.49611f
C12569 Iout.n852 VGND 0.08168f
C12570 Iout.t150 VGND 0.02304f
C12571 Iout.n853 VGND 0.05124f
C12572 Iout.n854 VGND 0.02606f
C12573 Iout.t72 VGND 0.02304f
C12574 Iout.n855 VGND 0.05124f
C12575 Iout.n856 VGND 0.02606f
C12576 Iout.n857 VGND 0.08168f
C12577 Iout.n858 VGND 0.49611f
C12578 Iout.n859 VGND 0.04775f
C12579 Iout.t164 VGND 0.02304f
C12580 Iout.n860 VGND 0.05124f
C12581 Iout.n861 VGND 0.02606f
C12582 Iout.t188 VGND 0.02304f
C12583 Iout.n862 VGND 0.05124f
C12584 Iout.n863 VGND 0.02606f
C12585 Iout.n864 VGND 0.04775f
C12586 Iout.n865 VGND 0.49611f
C12587 Iout.n866 VGND 0.08168f
C12588 Iout.t37 VGND 0.02304f
C12589 Iout.n867 VGND 0.05124f
C12590 Iout.n868 VGND 0.02606f
C12591 Iout.t49 VGND 0.02304f
C12592 Iout.n869 VGND 0.05124f
C12593 Iout.n870 VGND 0.02606f
C12594 Iout.n871 VGND 0.08168f
C12595 Iout.n872 VGND 0.49611f
C12596 Iout.n873 VGND 0.04775f
C12597 Iout.t182 VGND 0.02304f
C12598 Iout.n874 VGND 0.05124f
C12599 Iout.n875 VGND 0.02606f
C12600 Iout.t104 VGND 0.02304f
C12601 Iout.n876 VGND 0.05124f
C12602 Iout.n877 VGND 0.02606f
C12603 Iout.n878 VGND 0.04775f
C12604 Iout.n879 VGND 0.49611f
C12605 Iout.n880 VGND 0.08168f
C12606 Iout.t103 VGND 0.02304f
C12607 Iout.n881 VGND 0.05124f
C12608 Iout.n882 VGND 0.02606f
C12609 Iout.t162 VGND 0.02304f
C12610 Iout.n883 VGND 0.05124f
C12611 Iout.n884 VGND 0.02606f
C12612 Iout.n885 VGND 0.08168f
C12613 Iout.n886 VGND 0.49611f
C12614 Iout.n887 VGND 0.04775f
C12615 Iout.t192 VGND 0.02304f
C12616 Iout.n888 VGND 0.05124f
C12617 Iout.n889 VGND 0.02606f
C12618 Iout.t76 VGND 0.02304f
C12619 Iout.n890 VGND 0.05124f
C12620 Iout.n891 VGND 0.02606f
C12621 Iout.n892 VGND 0.04775f
C12622 Iout.n893 VGND 0.49611f
C12623 Iout.n894 VGND 0.08168f
C12624 Iout.t219 VGND 0.02304f
C12625 Iout.n895 VGND 0.05124f
C12626 Iout.n896 VGND 0.02606f
C12627 Iout.t44 VGND 0.02304f
C12628 Iout.n897 VGND 0.05124f
C12629 Iout.n898 VGND 0.02606f
C12630 Iout.n899 VGND 0.08168f
C12631 Iout.n900 VGND 0.49611f
C12632 Iout.n901 VGND 0.04775f
C12633 Iout.t137 VGND 0.02304f
C12634 Iout.n902 VGND 0.05124f
C12635 Iout.n903 VGND 0.02606f
C12636 Iout.t248 VGND 0.02304f
C12637 Iout.n904 VGND 0.05124f
C12638 Iout.n905 VGND 0.02606f
C12639 Iout.n906 VGND 0.04775f
C12640 Iout.n907 VGND 0.49611f
C12641 Iout.n908 VGND 0.08168f
C12642 Iout.t16 VGND 0.02304f
C12643 Iout.n909 VGND 0.05124f
C12644 Iout.n910 VGND 0.02606f
C12645 Iout.t95 VGND 0.02304f
C12646 Iout.n911 VGND 0.05124f
C12647 Iout.n912 VGND 0.02606f
C12648 Iout.n913 VGND 0.08168f
C12649 Iout.n914 VGND 0.49611f
C12650 Iout.n915 VGND 0.04775f
C12651 Iout.t249 VGND 0.02304f
C12652 Iout.n916 VGND 0.05124f
C12653 Iout.n917 VGND 0.02606f
C12654 Iout.t184 VGND 0.02304f
C12655 Iout.n918 VGND 0.05124f
C12656 Iout.n919 VGND 0.02606f
C12657 Iout.n920 VGND 0.04775f
C12658 Iout.n921 VGND 0.49611f
C12659 Iout.n922 VGND 0.08168f
C12660 Iout.t135 VGND 0.02304f
C12661 Iout.n923 VGND 0.05124f
C12662 Iout.n924 VGND 0.02606f
C12663 Iout.n925 VGND 0.08168f
C12664 Iout.t108 VGND 0.02304f
C12665 Iout.n926 VGND 0.05124f
C12666 Iout.n927 VGND 0.02606f
C12667 Iout.n928 VGND 0.08168f
C12668 Iout.n929 VGND 0.49611f
C12669 Iout.n930 VGND 0.04775f
C12670 Iout.t67 VGND 0.02304f
C12671 Iout.n931 VGND 0.05124f
C12672 Iout.n932 VGND 0.02606f
C12673 Iout.n933 VGND 0.04775f
C12674 Iout.t73 VGND 0.02304f
C12675 Iout.n934 VGND 0.05124f
C12676 Iout.n935 VGND 0.20242f
C12677 Iout.n936 VGND 2.65139f
C12678 Iout.n937 VGND 1.25122f
C12679 Iout.t244 VGND 0.02304f
C12680 Iout.n938 VGND 0.05124f
C12681 Iout.n939 VGND 0.20242f
C12682 Iout.n940 VGND 0.04775f
C12683 Iout.n941 VGND 0.23929f
C12684 Iout.n942 VGND 0.23929f
C12685 Iout.n943 VGND 0.04775f
C12686 Iout.t216 VGND 0.02304f
C12687 Iout.n944 VGND 0.05124f
C12688 Iout.n945 VGND 0.02606f
C12689 Iout.n946 VGND 0.04775f
C12690 Iout.n947 VGND 0.23929f
C12691 Iout.n948 VGND 0.23929f
C12692 Iout.n949 VGND 0.04775f
C12693 Iout.t187 VGND 0.02304f
C12694 Iout.n950 VGND 0.05124f
C12695 Iout.n951 VGND 0.02606f
C12696 Iout.n952 VGND 0.04775f
C12697 Iout.t204 VGND 0.02304f
C12698 Iout.n953 VGND 0.05124f
C12699 Iout.n954 VGND 0.20242f
C12700 Iout.n955 VGND 1.25122f
C12701 Iout.n956 VGND 1.25122f
C12702 Iout.t89 VGND 0.02304f
C12703 Iout.n957 VGND 0.05124f
C12704 Iout.n958 VGND 0.20242f
C12705 Iout.n959 VGND 0.04775f
C12706 Iout.n960 VGND 0.23929f
C12707 Iout.n961 VGND 0.23929f
C12708 Iout.n962 VGND 0.04775f
C12709 Iout.t48 VGND 0.02304f
C12710 Iout.n963 VGND 0.05124f
C12711 Iout.n964 VGND 0.02606f
C12712 Iout.n965 VGND 0.04775f
C12713 Iout.n966 VGND 0.23929f
C12714 Iout.n967 VGND 0.23929f
C12715 Iout.n968 VGND 0.04775f
C12716 Iout.t189 VGND 0.02304f
C12717 Iout.n969 VGND 0.05124f
C12718 Iout.n970 VGND 0.02606f
C12719 Iout.n971 VGND 0.04775f
C12720 Iout.t118 VGND 0.02304f
C12721 Iout.n972 VGND 0.05124f
C12722 Iout.n973 VGND 0.20242f
C12723 Iout.n974 VGND 1.25122f
C12724 Iout.n975 VGND 1.25122f
C12725 Iout.t207 VGND 0.02304f
C12726 Iout.n976 VGND 0.05124f
C12727 Iout.n977 VGND 0.20242f
C12728 Iout.n978 VGND 0.04775f
C12729 Iout.n979 VGND 0.23929f
C12730 Iout.n980 VGND 0.23929f
C12731 Iout.n981 VGND 0.04775f
C12732 Iout.t115 VGND 0.02304f
C12733 Iout.n982 VGND 0.05124f
C12734 Iout.n983 VGND 0.02606f
C12735 Iout.n984 VGND 0.04775f
C12736 Iout.n985 VGND 0.23929f
C12737 Iout.n986 VGND 0.23929f
C12738 Iout.n987 VGND 0.04775f
C12739 Iout.t102 VGND 0.02304f
C12740 Iout.n988 VGND 0.05124f
C12741 Iout.n989 VGND 0.02606f
C12742 Iout.n990 VGND 0.04775f
C12743 Iout.t196 VGND 0.02304f
C12744 Iout.n991 VGND 0.05124f
C12745 Iout.n992 VGND 0.20242f
C12746 Iout.n993 VGND 1.25122f
C12747 Iout.n994 VGND 1.25122f
C12748 Iout.t57 VGND 0.02304f
C12749 Iout.n995 VGND 0.05124f
C12750 Iout.n996 VGND 0.20242f
C12751 Iout.n997 VGND 0.04775f
C12752 Iout.n998 VGND 0.23929f
C12753 Iout.n999 VGND 0.23929f
C12754 Iout.n1000 VGND 0.04775f
C12755 Iout.t217 VGND 0.02304f
C12756 Iout.n1001 VGND 0.05124f
C12757 Iout.n1002 VGND 0.02606f
C12758 Iout.n1003 VGND 0.04775f
C12759 Iout.n1004 VGND 0.23929f
C12760 Iout.n1005 VGND 0.23929f
C12761 Iout.n1006 VGND 0.04775f
C12762 Iout.t191 VGND 0.02304f
C12763 Iout.n1007 VGND 0.05124f
C12764 Iout.n1008 VGND 0.02606f
C12765 Iout.n1009 VGND 0.04775f
C12766 Iout.t149 VGND 0.02304f
C12767 Iout.n1010 VGND 0.05124f
C12768 Iout.n1011 VGND 0.20242f
C12769 Iout.n1012 VGND 1.25122f
C12770 Iout.n1013 VGND 1.1235f
C12771 Iout.t93 VGND 0.02304f
C12772 Iout.n1014 VGND 0.05124f
C12773 Iout.n1015 VGND 0.20242f
C12774 Iout.n1016 VGND 0.04775f
C12775 Iout.n1017 VGND 0.23929f
C12776 Iout.n1018 VGND 0.14126f
C12777 Iout.n1019 VGND 0.04775f
C12778 Iout.t148 VGND 0.02304f
C12779 Iout.n1020 VGND 0.05124f
C12780 Iout.n1021 VGND 0.20242f
C12781 Iout.n1022 VGND 0.23244f
C12782 XThC.Tn[4].t5 VGND 0.01821f
C12783 XThC.Tn[4].t4 VGND 0.01821f
C12784 XThC.Tn[4].n0 VGND 0.03675f
C12785 XThC.Tn[4].t7 VGND 0.01821f
C12786 XThC.Tn[4].t6 VGND 0.01821f
C12787 XThC.Tn[4].n1 VGND 0.043f
C12788 XThC.Tn[4].n2 VGND 0.12038f
C12789 XThC.Tn[4].t1 VGND 0.01183f
C12790 XThC.Tn[4].t0 VGND 0.01183f
C12791 XThC.Tn[4].n3 VGND 0.02695f
C12792 XThC.Tn[4].t8 VGND 0.01183f
C12793 XThC.Tn[4].t11 VGND 0.01183f
C12794 XThC.Tn[4].n4 VGND 0.0449f
C12795 XThC.Tn[4].t10 VGND 0.01183f
C12796 XThC.Tn[4].t9 VGND 0.01183f
C12797 XThC.Tn[4].n5 VGND 0.02695f
C12798 XThC.Tn[4].n6 VGND 0.12834f
C12799 XThC.Tn[4].t3 VGND 0.01183f
C12800 XThC.Tn[4].t2 VGND 0.01183f
C12801 XThC.Tn[4].n7 VGND 0.02695f
C12802 XThC.Tn[4].n8 VGND 0.07934f
C12803 XThC.Tn[4].n9 VGND 0.08954f
C12804 XThC.Tn[4].t28 VGND 0.01443f
C12805 XThC.Tn[4].t26 VGND 0.01576f
C12806 XThC.Tn[4].n10 VGND 0.03519f
C12807 XThC.Tn[4].n11 VGND 0.02411f
C12808 XThC.Tn[4].n12 VGND 0.07913f
C12809 XThC.Tn[4].t14 VGND 0.01443f
C12810 XThC.Tn[4].t43 VGND 0.01576f
C12811 XThC.Tn[4].n13 VGND 0.03519f
C12812 XThC.Tn[4].n14 VGND 0.02411f
C12813 XThC.Tn[4].n15 VGND 0.07935f
C12814 XThC.Tn[4].n16 VGND 0.13077f
C12815 XThC.Tn[4].t19 VGND 0.01443f
C12816 XThC.Tn[4].t13 VGND 0.01576f
C12817 XThC.Tn[4].n17 VGND 0.03519f
C12818 XThC.Tn[4].n18 VGND 0.02411f
C12819 XThC.Tn[4].n19 VGND 0.07935f
C12820 XThC.Tn[4].n20 VGND 0.13077f
C12821 XThC.Tn[4].t20 VGND 0.01443f
C12822 XThC.Tn[4].t15 VGND 0.01576f
C12823 XThC.Tn[4].n21 VGND 0.03519f
C12824 XThC.Tn[4].n22 VGND 0.02411f
C12825 XThC.Tn[4].n23 VGND 0.07935f
C12826 XThC.Tn[4].n24 VGND 0.13077f
C12827 XThC.Tn[4].t39 VGND 0.01443f
C12828 XThC.Tn[4].t36 VGND 0.01576f
C12829 XThC.Tn[4].n25 VGND 0.03519f
C12830 XThC.Tn[4].n26 VGND 0.02411f
C12831 XThC.Tn[4].n27 VGND 0.07935f
C12832 XThC.Tn[4].n28 VGND 0.13077f
C12833 XThC.Tn[4].t40 VGND 0.01443f
C12834 XThC.Tn[4].t37 VGND 0.01576f
C12835 XThC.Tn[4].n29 VGND 0.03519f
C12836 XThC.Tn[4].n30 VGND 0.02411f
C12837 XThC.Tn[4].n31 VGND 0.07935f
C12838 XThC.Tn[4].n32 VGND 0.13077f
C12839 XThC.Tn[4].t24 VGND 0.01443f
C12840 XThC.Tn[4].t18 VGND 0.01576f
C12841 XThC.Tn[4].n33 VGND 0.03519f
C12842 XThC.Tn[4].n34 VGND 0.02411f
C12843 XThC.Tn[4].n35 VGND 0.07935f
C12844 XThC.Tn[4].n36 VGND 0.13077f
C12845 XThC.Tn[4].t31 VGND 0.01443f
C12846 XThC.Tn[4].t27 VGND 0.01576f
C12847 XThC.Tn[4].n37 VGND 0.03519f
C12848 XThC.Tn[4].n38 VGND 0.02411f
C12849 XThC.Tn[4].n39 VGND 0.07935f
C12850 XThC.Tn[4].n40 VGND 0.13077f
C12851 XThC.Tn[4].t33 VGND 0.01443f
C12852 XThC.Tn[4].t29 VGND 0.01576f
C12853 XThC.Tn[4].n41 VGND 0.03519f
C12854 XThC.Tn[4].n42 VGND 0.02411f
C12855 XThC.Tn[4].n43 VGND 0.07935f
C12856 XThC.Tn[4].n44 VGND 0.13077f
C12857 XThC.Tn[4].t21 VGND 0.01443f
C12858 XThC.Tn[4].t16 VGND 0.01576f
C12859 XThC.Tn[4].n45 VGND 0.03519f
C12860 XThC.Tn[4].n46 VGND 0.02411f
C12861 XThC.Tn[4].n47 VGND 0.07935f
C12862 XThC.Tn[4].n48 VGND 0.13077f
C12863 XThC.Tn[4].t23 VGND 0.01443f
C12864 XThC.Tn[4].t17 VGND 0.01576f
C12865 XThC.Tn[4].n49 VGND 0.03519f
C12866 XThC.Tn[4].n50 VGND 0.02411f
C12867 XThC.Tn[4].n51 VGND 0.07935f
C12868 XThC.Tn[4].n52 VGND 0.13077f
C12869 XThC.Tn[4].t34 VGND 0.01443f
C12870 XThC.Tn[4].t30 VGND 0.01576f
C12871 XThC.Tn[4].n53 VGND 0.03519f
C12872 XThC.Tn[4].n54 VGND 0.02411f
C12873 XThC.Tn[4].n55 VGND 0.07935f
C12874 XThC.Tn[4].n56 VGND 0.13077f
C12875 XThC.Tn[4].t42 VGND 0.01443f
C12876 XThC.Tn[4].t38 VGND 0.01576f
C12877 XThC.Tn[4].n57 VGND 0.03519f
C12878 XThC.Tn[4].n58 VGND 0.02411f
C12879 XThC.Tn[4].n59 VGND 0.07935f
C12880 XThC.Tn[4].n60 VGND 0.13077f
C12881 XThC.Tn[4].t12 VGND 0.01443f
C12882 XThC.Tn[4].t41 VGND 0.01576f
C12883 XThC.Tn[4].n61 VGND 0.03519f
C12884 XThC.Tn[4].n62 VGND 0.02411f
C12885 XThC.Tn[4].n63 VGND 0.07935f
C12886 XThC.Tn[4].n64 VGND 0.13077f
C12887 XThC.Tn[4].t25 VGND 0.01443f
C12888 XThC.Tn[4].t22 VGND 0.01576f
C12889 XThC.Tn[4].n65 VGND 0.03519f
C12890 XThC.Tn[4].n66 VGND 0.02411f
C12891 XThC.Tn[4].n67 VGND 0.07935f
C12892 XThC.Tn[4].n68 VGND 0.13077f
C12893 XThC.Tn[4].t35 VGND 0.01443f
C12894 XThC.Tn[4].t32 VGND 0.01576f
C12895 XThC.Tn[4].n69 VGND 0.03519f
C12896 XThC.Tn[4].n70 VGND 0.02411f
C12897 XThC.Tn[4].n71 VGND 0.07935f
C12898 XThC.Tn[4].n72 VGND 0.13077f
C12899 XThC.Tn[4].n73 VGND 0.16028f
C12900 XThC.Tn[4].n74 VGND 0.0381f
C12901 XThR.Tn[5].t8 VGND 0.01513f
C12902 XThR.Tn[5].t9 VGND 0.01513f
C12903 XThR.Tn[5].n0 VGND 0.0574f
C12904 XThR.Tn[5].t11 VGND 0.01513f
C12905 XThR.Tn[5].t10 VGND 0.01513f
C12906 XThR.Tn[5].n1 VGND 0.03445f
C12907 XThR.Tn[5].n2 VGND 0.16407f
C12908 XThR.Tn[5].t6 VGND 0.01513f
C12909 XThR.Tn[5].t5 VGND 0.01513f
C12910 XThR.Tn[5].n3 VGND 0.03445f
C12911 XThR.Tn[5].n4 VGND 0.10142f
C12912 XThR.Tn[5].t7 VGND 0.01513f
C12913 XThR.Tn[5].t4 VGND 0.01513f
C12914 XThR.Tn[5].n5 VGND 0.03445f
C12915 XThR.Tn[5].n6 VGND 0.11446f
C12916 XThR.Tn[5].t17 VGND 0.01819f
C12917 XThR.Tn[5].t72 VGND 0.01992f
C12918 XThR.Tn[5].n7 VGND 0.04864f
C12919 XThR.Tn[5].n8 VGND 0.09344f
C12920 XThR.Tn[5].t39 VGND 0.01819f
C12921 XThR.Tn[5].t26 VGND 0.01992f
C12922 XThR.Tn[5].n9 VGND 0.04864f
C12923 XThR.Tn[5].t13 VGND 0.01813f
C12924 XThR.Tn[5].t23 VGND 0.01985f
C12925 XThR.Tn[5].n10 VGND 0.05061f
C12926 XThR.Tn[5].n11 VGND 0.03555f
C12927 XThR.Tn[5].n12 VGND 0.0065f
C12928 XThR.Tn[5].n13 VGND 0.11409f
C12929 XThR.Tn[5].t73 VGND 0.01819f
C12930 XThR.Tn[5].t66 VGND 0.01992f
C12931 XThR.Tn[5].n14 VGND 0.04864f
C12932 XThR.Tn[5].t48 VGND 0.01813f
C12933 XThR.Tn[5].t61 VGND 0.01985f
C12934 XThR.Tn[5].n15 VGND 0.05061f
C12935 XThR.Tn[5].n16 VGND 0.03555f
C12936 XThR.Tn[5].n17 VGND 0.0065f
C12937 XThR.Tn[5].n18 VGND 0.11409f
C12938 XThR.Tn[5].t28 VGND 0.01819f
C12939 XThR.Tn[5].t21 VGND 0.01992f
C12940 XThR.Tn[5].n19 VGND 0.04864f
C12941 XThR.Tn[5].t65 VGND 0.01813f
C12942 XThR.Tn[5].t18 VGND 0.01985f
C12943 XThR.Tn[5].n20 VGND 0.05061f
C12944 XThR.Tn[5].n21 VGND 0.03555f
C12945 XThR.Tn[5].n22 VGND 0.0065f
C12946 XThR.Tn[5].n23 VGND 0.11409f
C12947 XThR.Tn[5].t55 VGND 0.01819f
C12948 XThR.Tn[5].t51 VGND 0.01992f
C12949 XThR.Tn[5].n24 VGND 0.04864f
C12950 XThR.Tn[5].t33 VGND 0.01813f
C12951 XThR.Tn[5].t46 VGND 0.01985f
C12952 XThR.Tn[5].n25 VGND 0.05061f
C12953 XThR.Tn[5].n26 VGND 0.03555f
C12954 XThR.Tn[5].n27 VGND 0.0065f
C12955 XThR.Tn[5].n28 VGND 0.11409f
C12956 XThR.Tn[5].t30 VGND 0.01819f
C12957 XThR.Tn[5].t22 VGND 0.01992f
C12958 XThR.Tn[5].n29 VGND 0.04864f
C12959 XThR.Tn[5].t67 VGND 0.01813f
C12960 XThR.Tn[5].t19 VGND 0.01985f
C12961 XThR.Tn[5].n30 VGND 0.05061f
C12962 XThR.Tn[5].n31 VGND 0.03555f
C12963 XThR.Tn[5].n32 VGND 0.0065f
C12964 XThR.Tn[5].n33 VGND 0.11409f
C12965 XThR.Tn[5].t69 VGND 0.01819f
C12966 XThR.Tn[5].t40 VGND 0.01992f
C12967 XThR.Tn[5].n34 VGND 0.04864f
C12968 XThR.Tn[5].t43 VGND 0.01813f
C12969 XThR.Tn[5].t37 VGND 0.01985f
C12970 XThR.Tn[5].n35 VGND 0.05061f
C12971 XThR.Tn[5].n36 VGND 0.03555f
C12972 XThR.Tn[5].n37 VGND 0.0065f
C12973 XThR.Tn[5].n38 VGND 0.11409f
C12974 XThR.Tn[5].t38 VGND 0.01819f
C12975 XThR.Tn[5].t32 VGND 0.01992f
C12976 XThR.Tn[5].n39 VGND 0.04864f
C12977 XThR.Tn[5].t14 VGND 0.01813f
C12978 XThR.Tn[5].t29 VGND 0.01985f
C12979 XThR.Tn[5].n40 VGND 0.05061f
C12980 XThR.Tn[5].n41 VGND 0.03555f
C12981 XThR.Tn[5].n42 VGND 0.0065f
C12982 XThR.Tn[5].n43 VGND 0.11409f
C12983 XThR.Tn[5].t42 VGND 0.01819f
C12984 XThR.Tn[5].t49 VGND 0.01992f
C12985 XThR.Tn[5].n44 VGND 0.04864f
C12986 XThR.Tn[5].t16 VGND 0.01813f
C12987 XThR.Tn[5].t45 VGND 0.01985f
C12988 XThR.Tn[5].n45 VGND 0.05061f
C12989 XThR.Tn[5].n46 VGND 0.03555f
C12990 XThR.Tn[5].n47 VGND 0.0065f
C12991 XThR.Tn[5].n48 VGND 0.11409f
C12992 XThR.Tn[5].t58 VGND 0.01819f
C12993 XThR.Tn[5].t68 VGND 0.01992f
C12994 XThR.Tn[5].n49 VGND 0.04864f
C12995 XThR.Tn[5].t36 VGND 0.01813f
C12996 XThR.Tn[5].t63 VGND 0.01985f
C12997 XThR.Tn[5].n50 VGND 0.05061f
C12998 XThR.Tn[5].n51 VGND 0.03555f
C12999 XThR.Tn[5].n52 VGND 0.0065f
C13000 XThR.Tn[5].n53 VGND 0.11409f
C13001 XThR.Tn[5].t53 VGND 0.01819f
C13002 XThR.Tn[5].t24 VGND 0.01992f
C13003 XThR.Tn[5].n54 VGND 0.04864f
C13004 XThR.Tn[5].t25 VGND 0.01813f
C13005 XThR.Tn[5].t20 VGND 0.01985f
C13006 XThR.Tn[5].n55 VGND 0.05061f
C13007 XThR.Tn[5].n56 VGND 0.03555f
C13008 XThR.Tn[5].n57 VGND 0.0065f
C13009 XThR.Tn[5].n58 VGND 0.11409f
C13010 XThR.Tn[5].t71 VGND 0.01819f
C13011 XThR.Tn[5].t60 VGND 0.01992f
C13012 XThR.Tn[5].n59 VGND 0.04864f
C13013 XThR.Tn[5].t44 VGND 0.01813f
C13014 XThR.Tn[5].t57 VGND 0.01985f
C13015 XThR.Tn[5].n60 VGND 0.05061f
C13016 XThR.Tn[5].n61 VGND 0.03555f
C13017 XThR.Tn[5].n62 VGND 0.0065f
C13018 XThR.Tn[5].n63 VGND 0.11409f
C13019 XThR.Tn[5].t41 VGND 0.01819f
C13020 XThR.Tn[5].t35 VGND 0.01992f
C13021 XThR.Tn[5].n64 VGND 0.04864f
C13022 XThR.Tn[5].t15 VGND 0.01813f
C13023 XThR.Tn[5].t31 VGND 0.01985f
C13024 XThR.Tn[5].n65 VGND 0.05061f
C13025 XThR.Tn[5].n66 VGND 0.03555f
C13026 XThR.Tn[5].n67 VGND 0.0065f
C13027 XThR.Tn[5].n68 VGND 0.11409f
C13028 XThR.Tn[5].t56 VGND 0.01819f
C13029 XThR.Tn[5].t52 VGND 0.01992f
C13030 XThR.Tn[5].n69 VGND 0.04864f
C13031 XThR.Tn[5].t34 VGND 0.01813f
C13032 XThR.Tn[5].t47 VGND 0.01985f
C13033 XThR.Tn[5].n70 VGND 0.05061f
C13034 XThR.Tn[5].n71 VGND 0.03555f
C13035 XThR.Tn[5].n72 VGND 0.0065f
C13036 XThR.Tn[5].n73 VGND 0.11409f
C13037 XThR.Tn[5].t12 VGND 0.01819f
C13038 XThR.Tn[5].t70 VGND 0.01992f
C13039 XThR.Tn[5].n74 VGND 0.04864f
C13040 XThR.Tn[5].t50 VGND 0.01813f
C13041 XThR.Tn[5].t64 VGND 0.01985f
C13042 XThR.Tn[5].n75 VGND 0.05061f
C13043 XThR.Tn[5].n76 VGND 0.03555f
C13044 XThR.Tn[5].n77 VGND 0.0065f
C13045 XThR.Tn[5].n78 VGND 0.11409f
C13046 XThR.Tn[5].t54 VGND 0.01819f
C13047 XThR.Tn[5].t62 VGND 0.01992f
C13048 XThR.Tn[5].n79 VGND 0.04864f
C13049 XThR.Tn[5].t27 VGND 0.01813f
C13050 XThR.Tn[5].t59 VGND 0.01985f
C13051 XThR.Tn[5].n80 VGND 0.05061f
C13052 XThR.Tn[5].n81 VGND 0.03555f
C13053 XThR.Tn[5].n82 VGND 0.0065f
C13054 XThR.Tn[5].n83 VGND 0.11409f
C13055 XThR.Tn[5].n84 VGND 0.10368f
C13056 XThR.Tn[5].n85 VGND 0.20081f
C13057 XThR.Tn[5].t2 VGND 0.02327f
C13058 XThR.Tn[5].t3 VGND 0.02327f
C13059 XThR.Tn[5].n86 VGND 0.04698f
C13060 XThR.Tn[5].t1 VGND 0.02327f
C13061 XThR.Tn[5].t0 VGND 0.02327f
C13062 XThR.Tn[5].n87 VGND 0.05497f
C13063 XThR.Tn[5].n88 VGND 0.15388f
C13064 XThR.Tn[5].n89 VGND 0.0487f
C13065 XThR.Tn[3].t4 VGND 0.02315f
C13066 XThR.Tn[3].t5 VGND 0.02315f
C13067 XThR.Tn[3].n0 VGND 0.04673f
C13068 XThR.Tn[3].t3 VGND 0.02315f
C13069 XThR.Tn[3].t6 VGND 0.02315f
C13070 XThR.Tn[3].n1 VGND 0.05468f
C13071 XThR.Tn[3].n2 VGND 0.15307f
C13072 XThR.Tn[3].t10 VGND 0.01505f
C13073 XThR.Tn[3].t7 VGND 0.01505f
C13074 XThR.Tn[3].n3 VGND 0.03427f
C13075 XThR.Tn[3].t9 VGND 0.01505f
C13076 XThR.Tn[3].t8 VGND 0.01505f
C13077 XThR.Tn[3].n4 VGND 0.03427f
C13078 XThR.Tn[3].t11 VGND 0.01505f
C13079 XThR.Tn[3].t1 VGND 0.01505f
C13080 XThR.Tn[3].n5 VGND 0.0571f
C13081 XThR.Tn[3].t2 VGND 0.01505f
C13082 XThR.Tn[3].t0 VGND 0.01505f
C13083 XThR.Tn[3].n6 VGND 0.03427f
C13084 XThR.Tn[3].n7 VGND 0.16319f
C13085 XThR.Tn[3].n8 VGND 0.10088f
C13086 XThR.Tn[3].n9 VGND 0.11385f
C13087 XThR.Tn[3].t64 VGND 0.01809f
C13088 XThR.Tn[3].t57 VGND 0.01981f
C13089 XThR.Tn[3].n10 VGND 0.04838f
C13090 XThR.Tn[3].n11 VGND 0.09294f
C13091 XThR.Tn[3].t18 VGND 0.01809f
C13092 XThR.Tn[3].t70 VGND 0.01981f
C13093 XThR.Tn[3].n12 VGND 0.04838f
C13094 XThR.Tn[3].t24 VGND 0.01803f
C13095 XThR.Tn[3].t55 VGND 0.01975f
C13096 XThR.Tn[3].n13 VGND 0.05034f
C13097 XThR.Tn[3].n14 VGND 0.03536f
C13098 XThR.Tn[3].n15 VGND 0.00647f
C13099 XThR.Tn[3].n16 VGND 0.11349f
C13100 XThR.Tn[3].t59 VGND 0.01809f
C13101 XThR.Tn[3].t49 VGND 0.01981f
C13102 XThR.Tn[3].n17 VGND 0.04838f
C13103 XThR.Tn[3].t62 VGND 0.01803f
C13104 XThR.Tn[3].t29 VGND 0.01975f
C13105 XThR.Tn[3].n18 VGND 0.05034f
C13106 XThR.Tn[3].n19 VGND 0.03536f
C13107 XThR.Tn[3].n20 VGND 0.00647f
C13108 XThR.Tn[3].n21 VGND 0.11349f
C13109 XThR.Tn[3].t71 VGND 0.01809f
C13110 XThR.Tn[3].t67 VGND 0.01981f
C13111 XThR.Tn[3].n22 VGND 0.04838f
C13112 XThR.Tn[3].t12 VGND 0.01803f
C13113 XThR.Tn[3].t47 VGND 0.01975f
C13114 XThR.Tn[3].n23 VGND 0.05034f
C13115 XThR.Tn[3].n24 VGND 0.03536f
C13116 XThR.Tn[3].n25 VGND 0.00647f
C13117 XThR.Tn[3].n26 VGND 0.11349f
C13118 XThR.Tn[3].t39 VGND 0.01809f
C13119 XThR.Tn[3].t33 VGND 0.01981f
C13120 XThR.Tn[3].n27 VGND 0.04838f
C13121 XThR.Tn[3].t42 VGND 0.01803f
C13122 XThR.Tn[3].t13 VGND 0.01975f
C13123 XThR.Tn[3].n28 VGND 0.05034f
C13124 XThR.Tn[3].n29 VGND 0.03536f
C13125 XThR.Tn[3].n30 VGND 0.00647f
C13126 XThR.Tn[3].n31 VGND 0.11349f
C13127 XThR.Tn[3].t72 VGND 0.01809f
C13128 XThR.Tn[3].t68 VGND 0.01981f
C13129 XThR.Tn[3].n32 VGND 0.04838f
C13130 XThR.Tn[3].t16 VGND 0.01803f
C13131 XThR.Tn[3].t48 VGND 0.01975f
C13132 XThR.Tn[3].n33 VGND 0.05034f
C13133 XThR.Tn[3].n34 VGND 0.03536f
C13134 XThR.Tn[3].n35 VGND 0.00647f
C13135 XThR.Tn[3].n36 VGND 0.11349f
C13136 XThR.Tn[3].t52 VGND 0.01809f
C13137 XThR.Tn[3].t20 VGND 0.01981f
C13138 XThR.Tn[3].n37 VGND 0.04838f
C13139 XThR.Tn[3].t56 VGND 0.01803f
C13140 XThR.Tn[3].t66 VGND 0.01975f
C13141 XThR.Tn[3].n38 VGND 0.05034f
C13142 XThR.Tn[3].n39 VGND 0.03536f
C13143 XThR.Tn[3].n40 VGND 0.00647f
C13144 XThR.Tn[3].n41 VGND 0.11349f
C13145 XThR.Tn[3].t19 VGND 0.01809f
C13146 XThR.Tn[3].t14 VGND 0.01981f
C13147 XThR.Tn[3].n42 VGND 0.04838f
C13148 XThR.Tn[3].t23 VGND 0.01803f
C13149 XThR.Tn[3].t61 VGND 0.01975f
C13150 XThR.Tn[3].n43 VGND 0.05034f
C13151 XThR.Tn[3].n44 VGND 0.03536f
C13152 XThR.Tn[3].n45 VGND 0.00647f
C13153 XThR.Tn[3].n46 VGND 0.11349f
C13154 XThR.Tn[3].t22 VGND 0.01809f
C13155 XThR.Tn[3].t31 VGND 0.01981f
C13156 XThR.Tn[3].n47 VGND 0.04838f
C13157 XThR.Tn[3].t28 VGND 0.01803f
C13158 XThR.Tn[3].t73 VGND 0.01975f
C13159 XThR.Tn[3].n48 VGND 0.05034f
C13160 XThR.Tn[3].n49 VGND 0.03536f
C13161 XThR.Tn[3].n50 VGND 0.00647f
C13162 XThR.Tn[3].n51 VGND 0.11349f
C13163 XThR.Tn[3].t41 VGND 0.01809f
C13164 XThR.Tn[3].t51 VGND 0.01981f
C13165 XThR.Tn[3].n52 VGND 0.04838f
C13166 XThR.Tn[3].t45 VGND 0.01803f
C13167 XThR.Tn[3].t30 VGND 0.01975f
C13168 XThR.Tn[3].n53 VGND 0.05034f
C13169 XThR.Tn[3].n54 VGND 0.03536f
C13170 XThR.Tn[3].n55 VGND 0.00647f
C13171 XThR.Tn[3].n56 VGND 0.11349f
C13172 XThR.Tn[3].t35 VGND 0.01809f
C13173 XThR.Tn[3].t69 VGND 0.01981f
C13174 XThR.Tn[3].n57 VGND 0.04838f
C13175 XThR.Tn[3].t37 VGND 0.01803f
C13176 XThR.Tn[3].t50 VGND 0.01975f
C13177 XThR.Tn[3].n58 VGND 0.05034f
C13178 XThR.Tn[3].n59 VGND 0.03536f
C13179 XThR.Tn[3].n60 VGND 0.00647f
C13180 XThR.Tn[3].n61 VGND 0.11349f
C13181 XThR.Tn[3].t54 VGND 0.01809f
C13182 XThR.Tn[3].t44 VGND 0.01981f
C13183 XThR.Tn[3].n62 VGND 0.04838f
C13184 XThR.Tn[3].t58 VGND 0.01803f
C13185 XThR.Tn[3].t25 VGND 0.01975f
C13186 XThR.Tn[3].n63 VGND 0.05034f
C13187 XThR.Tn[3].n64 VGND 0.03536f
C13188 XThR.Tn[3].n65 VGND 0.00647f
C13189 XThR.Tn[3].n66 VGND 0.11349f
C13190 XThR.Tn[3].t21 VGND 0.01809f
C13191 XThR.Tn[3].t17 VGND 0.01981f
C13192 XThR.Tn[3].n67 VGND 0.04838f
C13193 XThR.Tn[3].t26 VGND 0.01803f
C13194 XThR.Tn[3].t63 VGND 0.01975f
C13195 XThR.Tn[3].n68 VGND 0.05034f
C13196 XThR.Tn[3].n69 VGND 0.03536f
C13197 XThR.Tn[3].n70 VGND 0.00647f
C13198 XThR.Tn[3].n71 VGND 0.11349f
C13199 XThR.Tn[3].t40 VGND 0.01809f
C13200 XThR.Tn[3].t34 VGND 0.01981f
C13201 XThR.Tn[3].n72 VGND 0.04838f
C13202 XThR.Tn[3].t43 VGND 0.01803f
C13203 XThR.Tn[3].t15 VGND 0.01975f
C13204 XThR.Tn[3].n73 VGND 0.05034f
C13205 XThR.Tn[3].n74 VGND 0.03536f
C13206 XThR.Tn[3].n75 VGND 0.00647f
C13207 XThR.Tn[3].n76 VGND 0.11349f
C13208 XThR.Tn[3].t60 VGND 0.01809f
C13209 XThR.Tn[3].t53 VGND 0.01981f
C13210 XThR.Tn[3].n77 VGND 0.04838f
C13211 XThR.Tn[3].t65 VGND 0.01803f
C13212 XThR.Tn[3].t32 VGND 0.01975f
C13213 XThR.Tn[3].n78 VGND 0.05034f
C13214 XThR.Tn[3].n79 VGND 0.03536f
C13215 XThR.Tn[3].n80 VGND 0.00647f
C13216 XThR.Tn[3].n81 VGND 0.11349f
C13217 XThR.Tn[3].t36 VGND 0.01809f
C13218 XThR.Tn[3].t46 VGND 0.01981f
C13219 XThR.Tn[3].n82 VGND 0.04838f
C13220 XThR.Tn[3].t38 VGND 0.01803f
C13221 XThR.Tn[3].t27 VGND 0.01975f
C13222 XThR.Tn[3].n83 VGND 0.05034f
C13223 XThR.Tn[3].n84 VGND 0.03536f
C13224 XThR.Tn[3].n85 VGND 0.00647f
C13225 XThR.Tn[3].n86 VGND 0.11349f
C13226 XThR.Tn[3].n87 VGND 0.10313f
C13227 XThR.Tn[3].n88 VGND 0.22842f
C13228 XThR.Tn[3].n89 VGND 0.04845f
C13229 XThC.XTB4.Y.t4 VGND 0.02956f
C13230 XThC.XTB4.Y.t13 VGND 0.05016f
C13231 XThC.XTB4.Y.n0 VGND 0.05972f
C13232 XThC.XTB4.Y.t7 VGND 0.02956f
C13233 XThC.XTB4.Y.t17 VGND 0.05016f
C13234 XThC.XTB4.Y.n1 VGND 0.03074f
C13235 XThC.XTB4.Y.t10 VGND 0.02956f
C13236 XThC.XTB4.Y.t2 VGND 0.05016f
C13237 XThC.XTB4.Y.n2 VGND 0.06603f
C13238 XThC.XTB4.Y.t14 VGND 0.02956f
C13239 XThC.XTB4.Y.t3 VGND 0.05016f
C13240 XThC.XTB4.Y.n3 VGND 0.0613f
C13241 XThC.XTB4.Y.n4 VGND 0.03729f
C13242 XThC.XTB4.Y.n5 VGND 0.06174f
C13243 XThC.XTB4.Y.n6 VGND 0.02389f
C13244 XThC.XTB4.Y.n7 VGND 0.02916f
C13245 XThC.XTB4.Y.n8 VGND 0.06603f
C13246 XThC.XTB4.Y.n9 VGND 0.0331f
C13247 XThC.XTB4.Y.n10 VGND 0.06459f
C13248 XThC.XTB4.Y.t5 VGND 0.02956f
C13249 XThC.XTB4.Y.t16 VGND 0.05016f
C13250 XThC.XTB4.Y.n11 VGND 0.06761f
C13251 XThC.XTB4.Y.t9 VGND 0.02956f
C13252 XThC.XTB4.Y.t6 VGND 0.05016f
C13253 XThC.XTB4.Y.t15 VGND 0.02956f
C13254 XThC.XTB4.Y.t12 VGND 0.05016f
C13255 XThC.XTB4.Y.t11 VGND 0.02956f
C13256 XThC.XTB4.Y.t8 VGND 0.05016f
C13257 XThC.XTB4.Y.n12 VGND 0.08416f
C13258 XThC.XTB4.Y.n13 VGND 0.08889f
C13259 XThC.XTB4.Y.n14 VGND 0.03426f
C13260 XThC.XTB4.Y.n15 VGND 0.07234f
C13261 XThC.XTB4.Y.n16 VGND 0.0331f
C13262 XThC.XTB4.Y.n17 VGND 0.02701f
C13263 XThC.XTB4.Y.n18 VGND 0.63971f
C13264 XThC.XTB4.Y.n19 VGND 1.30917f
C13265 XThC.XTB4.Y.t1 VGND 0.06491f
C13266 XThC.XTB4.Y.n20 VGND 0.11223f
C13267 XThC.XTB4.Y.t0 VGND 0.12238f
C13268 XThC.XTB4.Y.n21 VGND 0.16166f
C13269 XThC.Tn[0].t11 VGND 0.00786f
C13270 XThC.Tn[0].t10 VGND 0.00786f
C13271 XThC.Tn[0].n0 VGND 0.02982f
C13272 XThC.Tn[0].t8 VGND 0.00786f
C13273 XThC.Tn[0].t9 VGND 0.00786f
C13274 XThC.Tn[0].n1 VGND 0.01789f
C13275 XThC.Tn[0].n2 VGND 0.08522f
C13276 XThC.Tn[0].t7 VGND 0.00786f
C13277 XThC.Tn[0].t6 VGND 0.00786f
C13278 XThC.Tn[0].n3 VGND 0.01789f
C13279 XThC.Tn[0].n4 VGND 0.05268f
C13280 XThC.Tn[0].t5 VGND 0.00786f
C13281 XThC.Tn[0].t4 VGND 0.00786f
C13282 XThC.Tn[0].n5 VGND 0.01789f
C13283 XThC.Tn[0].n6 VGND 0.05945f
C13284 XThC.Tn[0].t18 VGND 0.00958f
C13285 XThC.Tn[0].t22 VGND 0.01047f
C13286 XThC.Tn[0].n7 VGND 0.02336f
C13287 XThC.Tn[0].n8 VGND 0.01601f
C13288 XThC.Tn[0].n9 VGND 0.05254f
C13289 XThC.Tn[0].t35 VGND 0.00958f
C13290 XThC.Tn[0].t41 VGND 0.01047f
C13291 XThC.Tn[0].n10 VGND 0.02336f
C13292 XThC.Tn[0].n11 VGND 0.01601f
C13293 XThC.Tn[0].n12 VGND 0.05268f
C13294 XThC.Tn[0].n13 VGND 0.08683f
C13295 XThC.Tn[0].t37 VGND 0.00958f
C13296 XThC.Tn[0].t12 VGND 0.01047f
C13297 XThC.Tn[0].n14 VGND 0.02336f
C13298 XThC.Tn[0].n15 VGND 0.01601f
C13299 XThC.Tn[0].n16 VGND 0.05268f
C13300 XThC.Tn[0].n17 VGND 0.08683f
C13301 XThC.Tn[0].t39 VGND 0.00958f
C13302 XThC.Tn[0].t13 VGND 0.01047f
C13303 XThC.Tn[0].n18 VGND 0.02336f
C13304 XThC.Tn[0].n19 VGND 0.01601f
C13305 XThC.Tn[0].n20 VGND 0.05268f
C13306 XThC.Tn[0].n21 VGND 0.08683f
C13307 XThC.Tn[0].t28 VGND 0.00958f
C13308 XThC.Tn[0].t32 VGND 0.01047f
C13309 XThC.Tn[0].n22 VGND 0.02336f
C13310 XThC.Tn[0].n23 VGND 0.01601f
C13311 XThC.Tn[0].n24 VGND 0.05268f
C13312 XThC.Tn[0].n25 VGND 0.08683f
C13313 XThC.Tn[0].t30 VGND 0.00958f
C13314 XThC.Tn[0].t34 VGND 0.01047f
C13315 XThC.Tn[0].n26 VGND 0.02336f
C13316 XThC.Tn[0].n27 VGND 0.01601f
C13317 XThC.Tn[0].n28 VGND 0.05268f
C13318 XThC.Tn[0].n29 VGND 0.08683f
C13319 XThC.Tn[0].t43 VGND 0.00958f
C13320 XThC.Tn[0].t17 VGND 0.01047f
C13321 XThC.Tn[0].n30 VGND 0.02336f
C13322 XThC.Tn[0].n31 VGND 0.01601f
C13323 XThC.Tn[0].n32 VGND 0.05268f
C13324 XThC.Tn[0].n33 VGND 0.08683f
C13325 XThC.Tn[0].t20 VGND 0.00958f
C13326 XThC.Tn[0].t25 VGND 0.01047f
C13327 XThC.Tn[0].n34 VGND 0.02336f
C13328 XThC.Tn[0].n35 VGND 0.01601f
C13329 XThC.Tn[0].n36 VGND 0.05268f
C13330 XThC.Tn[0].n37 VGND 0.08683f
C13331 XThC.Tn[0].t21 VGND 0.00958f
C13332 XThC.Tn[0].t26 VGND 0.01047f
C13333 XThC.Tn[0].n38 VGND 0.02336f
C13334 XThC.Tn[0].n39 VGND 0.01601f
C13335 XThC.Tn[0].n40 VGND 0.05268f
C13336 XThC.Tn[0].n41 VGND 0.08683f
C13337 XThC.Tn[0].t40 VGND 0.00958f
C13338 XThC.Tn[0].t15 VGND 0.01047f
C13339 XThC.Tn[0].n42 VGND 0.02336f
C13340 XThC.Tn[0].n43 VGND 0.01601f
C13341 XThC.Tn[0].n44 VGND 0.05268f
C13342 XThC.Tn[0].n45 VGND 0.08683f
C13343 XThC.Tn[0].t42 VGND 0.00958f
C13344 XThC.Tn[0].t16 VGND 0.01047f
C13345 XThC.Tn[0].n46 VGND 0.02336f
C13346 XThC.Tn[0].n47 VGND 0.01601f
C13347 XThC.Tn[0].n48 VGND 0.05268f
C13348 XThC.Tn[0].n49 VGND 0.08683f
C13349 XThC.Tn[0].t23 VGND 0.00958f
C13350 XThC.Tn[0].t27 VGND 0.01047f
C13351 XThC.Tn[0].n50 VGND 0.02336f
C13352 XThC.Tn[0].n51 VGND 0.01601f
C13353 XThC.Tn[0].n52 VGND 0.05268f
C13354 XThC.Tn[0].n53 VGND 0.08683f
C13355 XThC.Tn[0].t31 VGND 0.00958f
C13356 XThC.Tn[0].t36 VGND 0.01047f
C13357 XThC.Tn[0].n54 VGND 0.02336f
C13358 XThC.Tn[0].n55 VGND 0.01601f
C13359 XThC.Tn[0].n56 VGND 0.05268f
C13360 XThC.Tn[0].n57 VGND 0.08683f
C13361 XThC.Tn[0].t33 VGND 0.00958f
C13362 XThC.Tn[0].t38 VGND 0.01047f
C13363 XThC.Tn[0].n58 VGND 0.02336f
C13364 XThC.Tn[0].n59 VGND 0.01601f
C13365 XThC.Tn[0].n60 VGND 0.05268f
C13366 XThC.Tn[0].n61 VGND 0.08683f
C13367 XThC.Tn[0].t14 VGND 0.00958f
C13368 XThC.Tn[0].t19 VGND 0.01047f
C13369 XThC.Tn[0].n62 VGND 0.02336f
C13370 XThC.Tn[0].n63 VGND 0.01601f
C13371 XThC.Tn[0].n64 VGND 0.05268f
C13372 XThC.Tn[0].n65 VGND 0.08683f
C13373 XThC.Tn[0].t24 VGND 0.00958f
C13374 XThC.Tn[0].t29 VGND 0.01047f
C13375 XThC.Tn[0].n66 VGND 0.02336f
C13376 XThC.Tn[0].n67 VGND 0.01601f
C13377 XThC.Tn[0].n68 VGND 0.05268f
C13378 XThC.Tn[0].n69 VGND 0.08683f
C13379 XThC.Tn[0].n70 VGND 0.53339f
C13380 XThC.Tn[0].n71 VGND 0.06506f
C13381 XThC.Tn[0].t1 VGND 0.01209f
C13382 XThC.Tn[0].t0 VGND 0.01209f
C13383 XThC.Tn[0].n72 VGND 0.0244f
C13384 XThC.Tn[0].t3 VGND 0.01209f
C13385 XThC.Tn[0].t2 VGND 0.01209f
C13386 XThC.Tn[0].n73 VGND 0.02855f
C13387 XThC.Tn[0].n74 VGND 0.07993f
C13388 XThC.Tn[0].n75 VGND 0.0253f
C13389 XThC.Tn[13].t11 VGND 0.01267f
C13390 XThC.Tn[13].t9 VGND 0.01267f
C13391 XThC.Tn[13].n0 VGND 0.03161f
C13392 XThC.Tn[13].t8 VGND 0.01267f
C13393 XThC.Tn[13].t10 VGND 0.01267f
C13394 XThC.Tn[13].n1 VGND 0.02535f
C13395 XThC.Tn[13].n2 VGND 0.05845f
C13396 XThC.Tn[13].t29 VGND 0.01546f
C13397 XThC.Tn[13].t27 VGND 0.01688f
C13398 XThC.Tn[13].n3 VGND 0.03768f
C13399 XThC.Tn[13].n4 VGND 0.02582f
C13400 XThC.Tn[13].n5 VGND 0.08475f
C13401 XThC.Tn[13].t15 VGND 0.01546f
C13402 XThC.Tn[13].t12 VGND 0.01688f
C13403 XThC.Tn[13].n6 VGND 0.03768f
C13404 XThC.Tn[13].n7 VGND 0.02582f
C13405 XThC.Tn[13].n8 VGND 0.08498f
C13406 XThC.Tn[13].n9 VGND 0.14005f
C13407 XThC.Tn[13].t20 VGND 0.01546f
C13408 XThC.Tn[13].t14 VGND 0.01688f
C13409 XThC.Tn[13].n10 VGND 0.03768f
C13410 XThC.Tn[13].n11 VGND 0.02582f
C13411 XThC.Tn[13].n12 VGND 0.08498f
C13412 XThC.Tn[13].n13 VGND 0.14005f
C13413 XThC.Tn[13].t21 VGND 0.01546f
C13414 XThC.Tn[13].t16 VGND 0.01688f
C13415 XThC.Tn[13].n14 VGND 0.03768f
C13416 XThC.Tn[13].n15 VGND 0.02582f
C13417 XThC.Tn[13].n16 VGND 0.08498f
C13418 XThC.Tn[13].n17 VGND 0.14005f
C13419 XThC.Tn[13].t40 VGND 0.01546f
C13420 XThC.Tn[13].t37 VGND 0.01688f
C13421 XThC.Tn[13].n18 VGND 0.03768f
C13422 XThC.Tn[13].n19 VGND 0.02582f
C13423 XThC.Tn[13].n20 VGND 0.08498f
C13424 XThC.Tn[13].n21 VGND 0.14005f
C13425 XThC.Tn[13].t41 VGND 0.01546f
C13426 XThC.Tn[13].t38 VGND 0.01688f
C13427 XThC.Tn[13].n22 VGND 0.03768f
C13428 XThC.Tn[13].n23 VGND 0.02582f
C13429 XThC.Tn[13].n24 VGND 0.08498f
C13430 XThC.Tn[13].n25 VGND 0.14005f
C13431 XThC.Tn[13].t25 VGND 0.01546f
C13432 XThC.Tn[13].t19 VGND 0.01688f
C13433 XThC.Tn[13].n26 VGND 0.03768f
C13434 XThC.Tn[13].n27 VGND 0.02582f
C13435 XThC.Tn[13].n28 VGND 0.08498f
C13436 XThC.Tn[13].n29 VGND 0.14005f
C13437 XThC.Tn[13].t32 VGND 0.01546f
C13438 XThC.Tn[13].t28 VGND 0.01688f
C13439 XThC.Tn[13].n30 VGND 0.03768f
C13440 XThC.Tn[13].n31 VGND 0.02582f
C13441 XThC.Tn[13].n32 VGND 0.08498f
C13442 XThC.Tn[13].n33 VGND 0.14005f
C13443 XThC.Tn[13].t34 VGND 0.01546f
C13444 XThC.Tn[13].t30 VGND 0.01688f
C13445 XThC.Tn[13].n34 VGND 0.03768f
C13446 XThC.Tn[13].n35 VGND 0.02582f
C13447 XThC.Tn[13].n36 VGND 0.08498f
C13448 XThC.Tn[13].n37 VGND 0.14005f
C13449 XThC.Tn[13].t22 VGND 0.01546f
C13450 XThC.Tn[13].t17 VGND 0.01688f
C13451 XThC.Tn[13].n38 VGND 0.03768f
C13452 XThC.Tn[13].n39 VGND 0.02582f
C13453 XThC.Tn[13].n40 VGND 0.08498f
C13454 XThC.Tn[13].n41 VGND 0.14005f
C13455 XThC.Tn[13].t24 VGND 0.01546f
C13456 XThC.Tn[13].t18 VGND 0.01688f
C13457 XThC.Tn[13].n42 VGND 0.03768f
C13458 XThC.Tn[13].n43 VGND 0.02582f
C13459 XThC.Tn[13].n44 VGND 0.08498f
C13460 XThC.Tn[13].n45 VGND 0.14005f
C13461 XThC.Tn[13].t35 VGND 0.01546f
C13462 XThC.Tn[13].t31 VGND 0.01688f
C13463 XThC.Tn[13].n46 VGND 0.03768f
C13464 XThC.Tn[13].n47 VGND 0.02582f
C13465 XThC.Tn[13].n48 VGND 0.08498f
C13466 XThC.Tn[13].n49 VGND 0.14005f
C13467 XThC.Tn[13].t43 VGND 0.01546f
C13468 XThC.Tn[13].t39 VGND 0.01688f
C13469 XThC.Tn[13].n50 VGND 0.03768f
C13470 XThC.Tn[13].n51 VGND 0.02582f
C13471 XThC.Tn[13].n52 VGND 0.08498f
C13472 XThC.Tn[13].n53 VGND 0.14005f
C13473 XThC.Tn[13].t13 VGND 0.01546f
C13474 XThC.Tn[13].t42 VGND 0.01688f
C13475 XThC.Tn[13].n54 VGND 0.03768f
C13476 XThC.Tn[13].n55 VGND 0.02582f
C13477 XThC.Tn[13].n56 VGND 0.08498f
C13478 XThC.Tn[13].n57 VGND 0.14005f
C13479 XThC.Tn[13].t26 VGND 0.01546f
C13480 XThC.Tn[13].t23 VGND 0.01688f
C13481 XThC.Tn[13].n58 VGND 0.03768f
C13482 XThC.Tn[13].n59 VGND 0.02582f
C13483 XThC.Tn[13].n60 VGND 0.08498f
C13484 XThC.Tn[13].n61 VGND 0.14005f
C13485 XThC.Tn[13].t36 VGND 0.01546f
C13486 XThC.Tn[13].t33 VGND 0.01688f
C13487 XThC.Tn[13].n62 VGND 0.03768f
C13488 XThC.Tn[13].n63 VGND 0.02582f
C13489 XThC.Tn[13].n64 VGND 0.08498f
C13490 XThC.Tn[13].n65 VGND 0.14005f
C13491 XThC.Tn[13].n66 VGND 0.72631f
C13492 XThC.Tn[13].n67 VGND 0.25541f
C13493 XThC.Tn[13].t6 VGND 0.0195f
C13494 XThC.Tn[13].t5 VGND 0.0195f
C13495 XThC.Tn[13].n68 VGND 0.04213f
C13496 XThC.Tn[13].t4 VGND 0.0195f
C13497 XThC.Tn[13].t7 VGND 0.0195f
C13498 XThC.Tn[13].n69 VGND 0.06641f
C13499 XThC.Tn[13].n70 VGND 0.17588f
C13500 XThC.Tn[13].n71 VGND 0.01295f
C13501 XThC.Tn[13].t1 VGND 0.0195f
C13502 XThC.Tn[13].t0 VGND 0.0195f
C13503 XThC.Tn[13].n72 VGND 0.05921f
C13504 XThC.Tn[13].t3 VGND 0.0195f
C13505 XThC.Tn[13].t2 VGND 0.0195f
C13506 XThC.Tn[13].n73 VGND 0.04335f
C13507 XThC.Tn[13].n74 VGND 0.19292f
C13508 XThC.Tn[12].t11 VGND 0.01298f
C13509 XThC.Tn[12].t10 VGND 0.01298f
C13510 XThC.Tn[12].n0 VGND 0.03236f
C13511 XThC.Tn[12].t9 VGND 0.01298f
C13512 XThC.Tn[12].t8 VGND 0.01298f
C13513 XThC.Tn[12].n1 VGND 0.02595f
C13514 XThC.Tn[12].n2 VGND 0.06529f
C13515 XThC.Tn[12].t37 VGND 0.01582f
C13516 XThC.Tn[12].t35 VGND 0.01728f
C13517 XThC.Tn[12].n3 VGND 0.03858f
C13518 XThC.Tn[12].n4 VGND 0.02643f
C13519 XThC.Tn[12].n5 VGND 0.08676f
C13520 XThC.Tn[12].t23 VGND 0.01582f
C13521 XThC.Tn[12].t20 VGND 0.01728f
C13522 XThC.Tn[12].n6 VGND 0.03858f
C13523 XThC.Tn[12].n7 VGND 0.02643f
C13524 XThC.Tn[12].n8 VGND 0.087f
C13525 XThC.Tn[12].n9 VGND 0.14339f
C13526 XThC.Tn[12].t28 VGND 0.01582f
C13527 XThC.Tn[12].t22 VGND 0.01728f
C13528 XThC.Tn[12].n10 VGND 0.03858f
C13529 XThC.Tn[12].n11 VGND 0.02643f
C13530 XThC.Tn[12].n12 VGND 0.087f
C13531 XThC.Tn[12].n13 VGND 0.14339f
C13532 XThC.Tn[12].t29 VGND 0.01582f
C13533 XThC.Tn[12].t24 VGND 0.01728f
C13534 XThC.Tn[12].n14 VGND 0.03858f
C13535 XThC.Tn[12].n15 VGND 0.02643f
C13536 XThC.Tn[12].n16 VGND 0.087f
C13537 XThC.Tn[12].n17 VGND 0.14339f
C13538 XThC.Tn[12].t16 VGND 0.01582f
C13539 XThC.Tn[12].t13 VGND 0.01728f
C13540 XThC.Tn[12].n18 VGND 0.03858f
C13541 XThC.Tn[12].n19 VGND 0.02643f
C13542 XThC.Tn[12].n20 VGND 0.087f
C13543 XThC.Tn[12].n21 VGND 0.14339f
C13544 XThC.Tn[12].t17 VGND 0.01582f
C13545 XThC.Tn[12].t14 VGND 0.01728f
C13546 XThC.Tn[12].n22 VGND 0.03858f
C13547 XThC.Tn[12].n23 VGND 0.02643f
C13548 XThC.Tn[12].n24 VGND 0.087f
C13549 XThC.Tn[12].n25 VGND 0.14339f
C13550 XThC.Tn[12].t33 VGND 0.01582f
C13551 XThC.Tn[12].t27 VGND 0.01728f
C13552 XThC.Tn[12].n26 VGND 0.03858f
C13553 XThC.Tn[12].n27 VGND 0.02643f
C13554 XThC.Tn[12].n28 VGND 0.087f
C13555 XThC.Tn[12].n29 VGND 0.14339f
C13556 XThC.Tn[12].t40 VGND 0.01582f
C13557 XThC.Tn[12].t36 VGND 0.01728f
C13558 XThC.Tn[12].n30 VGND 0.03858f
C13559 XThC.Tn[12].n31 VGND 0.02643f
C13560 XThC.Tn[12].n32 VGND 0.087f
C13561 XThC.Tn[12].n33 VGND 0.14339f
C13562 XThC.Tn[12].t42 VGND 0.01582f
C13563 XThC.Tn[12].t38 VGND 0.01728f
C13564 XThC.Tn[12].n34 VGND 0.03858f
C13565 XThC.Tn[12].n35 VGND 0.02643f
C13566 XThC.Tn[12].n36 VGND 0.087f
C13567 XThC.Tn[12].n37 VGND 0.14339f
C13568 XThC.Tn[12].t30 VGND 0.01582f
C13569 XThC.Tn[12].t25 VGND 0.01728f
C13570 XThC.Tn[12].n38 VGND 0.03858f
C13571 XThC.Tn[12].n39 VGND 0.02643f
C13572 XThC.Tn[12].n40 VGND 0.087f
C13573 XThC.Tn[12].n41 VGND 0.14339f
C13574 XThC.Tn[12].t32 VGND 0.01582f
C13575 XThC.Tn[12].t26 VGND 0.01728f
C13576 XThC.Tn[12].n42 VGND 0.03858f
C13577 XThC.Tn[12].n43 VGND 0.02643f
C13578 XThC.Tn[12].n44 VGND 0.087f
C13579 XThC.Tn[12].n45 VGND 0.14339f
C13580 XThC.Tn[12].t43 VGND 0.01582f
C13581 XThC.Tn[12].t39 VGND 0.01728f
C13582 XThC.Tn[12].n46 VGND 0.03858f
C13583 XThC.Tn[12].n47 VGND 0.02643f
C13584 XThC.Tn[12].n48 VGND 0.087f
C13585 XThC.Tn[12].n49 VGND 0.14339f
C13586 XThC.Tn[12].t19 VGND 0.01582f
C13587 XThC.Tn[12].t15 VGND 0.01728f
C13588 XThC.Tn[12].n50 VGND 0.03858f
C13589 XThC.Tn[12].n51 VGND 0.02643f
C13590 XThC.Tn[12].n52 VGND 0.087f
C13591 XThC.Tn[12].n53 VGND 0.14339f
C13592 XThC.Tn[12].t21 VGND 0.01582f
C13593 XThC.Tn[12].t18 VGND 0.01728f
C13594 XThC.Tn[12].n54 VGND 0.03858f
C13595 XThC.Tn[12].n55 VGND 0.02643f
C13596 XThC.Tn[12].n56 VGND 0.087f
C13597 XThC.Tn[12].n57 VGND 0.14339f
C13598 XThC.Tn[12].t34 VGND 0.01582f
C13599 XThC.Tn[12].t31 VGND 0.01728f
C13600 XThC.Tn[12].n58 VGND 0.03858f
C13601 XThC.Tn[12].n59 VGND 0.02643f
C13602 XThC.Tn[12].n60 VGND 0.087f
C13603 XThC.Tn[12].n61 VGND 0.14339f
C13604 XThC.Tn[12].t12 VGND 0.01582f
C13605 XThC.Tn[12].t41 VGND 0.01728f
C13606 XThC.Tn[12].n62 VGND 0.03858f
C13607 XThC.Tn[12].n63 VGND 0.02643f
C13608 XThC.Tn[12].n64 VGND 0.087f
C13609 XThC.Tn[12].n65 VGND 0.14339f
C13610 XThC.Tn[12].n66 VGND 0.68185f
C13611 XThC.Tn[12].n67 VGND 0.24221f
C13612 XThC.Tn[12].t5 VGND 0.01996f
C13613 XThC.Tn[12].t6 VGND 0.01996f
C13614 XThC.Tn[12].n68 VGND 0.04313f
C13615 XThC.Tn[12].t4 VGND 0.01996f
C13616 XThC.Tn[12].t7 VGND 0.01996f
C13617 XThC.Tn[12].n69 VGND 0.06565f
C13618 XThC.Tn[12].n70 VGND 0.18241f
C13619 XThC.Tn[12].n71 VGND 0.02868f
C13620 XThC.Tn[12].t1 VGND 0.01996f
C13621 XThC.Tn[12].t0 VGND 0.01996f
C13622 XThC.Tn[12].n72 VGND 0.06062f
C13623 XThC.Tn[12].t3 VGND 0.01996f
C13624 XThC.Tn[12].t2 VGND 0.01996f
C13625 XThC.Tn[12].n73 VGND 0.04438f
C13626 XThC.Tn[12].n74 VGND 0.19752f
C13627 XThC.Tn[11].t8 VGND 0.01319f
C13628 XThC.Tn[11].t1 VGND 0.01319f
C13629 XThC.Tn[11].n0 VGND 0.0329f
C13630 XThC.Tn[11].t6 VGND 0.01319f
C13631 XThC.Tn[11].t10 VGND 0.01319f
C13632 XThC.Tn[11].n1 VGND 0.02638f
C13633 XThC.Tn[11].n2 VGND 0.06083f
C13634 XThC.Tn[11].t20 VGND 0.01608f
C13635 XThC.Tn[11].t18 VGND 0.01757f
C13636 XThC.Tn[11].n3 VGND 0.03922f
C13637 XThC.Tn[11].n4 VGND 0.02687f
C13638 XThC.Tn[11].n5 VGND 0.08819f
C13639 XThC.Tn[11].t38 VGND 0.01608f
C13640 XThC.Tn[11].t35 VGND 0.01757f
C13641 XThC.Tn[11].n6 VGND 0.03922f
C13642 XThC.Tn[11].n7 VGND 0.02687f
C13643 XThC.Tn[11].n8 VGND 0.08843f
C13644 XThC.Tn[11].n9 VGND 0.14574f
C13645 XThC.Tn[11].t43 VGND 0.01608f
C13646 XThC.Tn[11].t37 VGND 0.01757f
C13647 XThC.Tn[11].n10 VGND 0.03922f
C13648 XThC.Tn[11].n11 VGND 0.02687f
C13649 XThC.Tn[11].n12 VGND 0.08843f
C13650 XThC.Tn[11].n13 VGND 0.14574f
C13651 XThC.Tn[11].t12 VGND 0.01608f
C13652 XThC.Tn[11].t39 VGND 0.01757f
C13653 XThC.Tn[11].n14 VGND 0.03922f
C13654 XThC.Tn[11].n15 VGND 0.02687f
C13655 XThC.Tn[11].n16 VGND 0.08843f
C13656 XThC.Tn[11].n17 VGND 0.14574f
C13657 XThC.Tn[11].t31 VGND 0.01608f
C13658 XThC.Tn[11].t28 VGND 0.01757f
C13659 XThC.Tn[11].n18 VGND 0.03922f
C13660 XThC.Tn[11].n19 VGND 0.02687f
C13661 XThC.Tn[11].n20 VGND 0.08843f
C13662 XThC.Tn[11].n21 VGND 0.14574f
C13663 XThC.Tn[11].t32 VGND 0.01608f
C13664 XThC.Tn[11].t29 VGND 0.01757f
C13665 XThC.Tn[11].n22 VGND 0.03922f
C13666 XThC.Tn[11].n23 VGND 0.02687f
C13667 XThC.Tn[11].n24 VGND 0.08843f
C13668 XThC.Tn[11].n25 VGND 0.14574f
C13669 XThC.Tn[11].t16 VGND 0.01608f
C13670 XThC.Tn[11].t42 VGND 0.01757f
C13671 XThC.Tn[11].n26 VGND 0.03922f
C13672 XThC.Tn[11].n27 VGND 0.02687f
C13673 XThC.Tn[11].n28 VGND 0.08843f
C13674 XThC.Tn[11].n29 VGND 0.14574f
C13675 XThC.Tn[11].t23 VGND 0.01608f
C13676 XThC.Tn[11].t19 VGND 0.01757f
C13677 XThC.Tn[11].n30 VGND 0.03922f
C13678 XThC.Tn[11].n31 VGND 0.02687f
C13679 XThC.Tn[11].n32 VGND 0.08843f
C13680 XThC.Tn[11].n33 VGND 0.14574f
C13681 XThC.Tn[11].t25 VGND 0.01608f
C13682 XThC.Tn[11].t21 VGND 0.01757f
C13683 XThC.Tn[11].n34 VGND 0.03922f
C13684 XThC.Tn[11].n35 VGND 0.02687f
C13685 XThC.Tn[11].n36 VGND 0.08843f
C13686 XThC.Tn[11].n37 VGND 0.14574f
C13687 XThC.Tn[11].t13 VGND 0.01608f
C13688 XThC.Tn[11].t40 VGND 0.01757f
C13689 XThC.Tn[11].n38 VGND 0.03922f
C13690 XThC.Tn[11].n39 VGND 0.02687f
C13691 XThC.Tn[11].n40 VGND 0.08843f
C13692 XThC.Tn[11].n41 VGND 0.14574f
C13693 XThC.Tn[11].t15 VGND 0.01608f
C13694 XThC.Tn[11].t41 VGND 0.01757f
C13695 XThC.Tn[11].n42 VGND 0.03922f
C13696 XThC.Tn[11].n43 VGND 0.02687f
C13697 XThC.Tn[11].n44 VGND 0.08843f
C13698 XThC.Tn[11].n45 VGND 0.14574f
C13699 XThC.Tn[11].t26 VGND 0.01608f
C13700 XThC.Tn[11].t22 VGND 0.01757f
C13701 XThC.Tn[11].n46 VGND 0.03922f
C13702 XThC.Tn[11].n47 VGND 0.02687f
C13703 XThC.Tn[11].n48 VGND 0.08843f
C13704 XThC.Tn[11].n49 VGND 0.14574f
C13705 XThC.Tn[11].t34 VGND 0.01608f
C13706 XThC.Tn[11].t30 VGND 0.01757f
C13707 XThC.Tn[11].n50 VGND 0.03922f
C13708 XThC.Tn[11].n51 VGND 0.02687f
C13709 XThC.Tn[11].n52 VGND 0.08843f
C13710 XThC.Tn[11].n53 VGND 0.14574f
C13711 XThC.Tn[11].t36 VGND 0.01608f
C13712 XThC.Tn[11].t33 VGND 0.01757f
C13713 XThC.Tn[11].n54 VGND 0.03922f
C13714 XThC.Tn[11].n55 VGND 0.02687f
C13715 XThC.Tn[11].n56 VGND 0.08843f
C13716 XThC.Tn[11].n57 VGND 0.14574f
C13717 XThC.Tn[11].t17 VGND 0.01608f
C13718 XThC.Tn[11].t14 VGND 0.01757f
C13719 XThC.Tn[11].n58 VGND 0.03922f
C13720 XThC.Tn[11].n59 VGND 0.02687f
C13721 XThC.Tn[11].n60 VGND 0.08843f
C13722 XThC.Tn[11].n61 VGND 0.14574f
C13723 XThC.Tn[11].t27 VGND 0.01608f
C13724 XThC.Tn[11].t24 VGND 0.01757f
C13725 XThC.Tn[11].n62 VGND 0.03922f
C13726 XThC.Tn[11].n63 VGND 0.02687f
C13727 XThC.Tn[11].n64 VGND 0.08843f
C13728 XThC.Tn[11].n65 VGND 0.14574f
C13729 XThC.Tn[11].n66 VGND 0.6764f
C13730 XThC.Tn[11].n67 VGND 0.26496f
C13731 XThC.Tn[11].t11 VGND 0.02029f
C13732 XThC.Tn[11].t0 VGND 0.02029f
C13733 XThC.Tn[11].n68 VGND 0.04384f
C13734 XThC.Tn[11].t7 VGND 0.02029f
C13735 XThC.Tn[11].t9 VGND 0.02029f
C13736 XThC.Tn[11].n69 VGND 0.06911f
C13737 XThC.Tn[11].n70 VGND 0.18303f
C13738 XThC.Tn[11].n71 VGND 0.01348f
C13739 XThC.Tn[11].t2 VGND 0.02029f
C13740 XThC.Tn[11].t5 VGND 0.02029f
C13741 XThC.Tn[11].n72 VGND 0.06161f
C13742 XThC.Tn[11].t4 VGND 0.02029f
C13743 XThC.Tn[11].t3 VGND 0.02029f
C13744 XThC.Tn[11].n73 VGND 0.04511f
C13745 XThC.Tn[11].n74 VGND 0.20076f
C13746 XThC.Tn[9].t5 VGND 0.013f
C13747 XThC.Tn[9].t4 VGND 0.013f
C13748 XThC.Tn[9].n0 VGND 0.03242f
C13749 XThC.Tn[9].t6 VGND 0.013f
C13750 XThC.Tn[9].t7 VGND 0.013f
C13751 XThC.Tn[9].n1 VGND 0.026f
C13752 XThC.Tn[9].n2 VGND 0.05995f
C13753 XThC.Tn[9].t26 VGND 0.01585f
C13754 XThC.Tn[9].t12 VGND 0.01732f
C13755 XThC.Tn[9].n3 VGND 0.03865f
C13756 XThC.Tn[9].n4 VGND 0.02648f
C13757 XThC.Tn[9].n5 VGND 0.08692f
C13758 XThC.Tn[9].t13 VGND 0.01585f
C13759 XThC.Tn[9].t30 VGND 0.01732f
C13760 XThC.Tn[9].n6 VGND 0.03865f
C13761 XThC.Tn[9].n7 VGND 0.02648f
C13762 XThC.Tn[9].n8 VGND 0.08716f
C13763 XThC.Tn[9].n9 VGND 0.14365f
C13764 XThC.Tn[9].t15 VGND 0.01585f
C13765 XThC.Tn[9].t34 VGND 0.01732f
C13766 XThC.Tn[9].n10 VGND 0.03865f
C13767 XThC.Tn[9].n11 VGND 0.02648f
C13768 XThC.Tn[9].n12 VGND 0.08716f
C13769 XThC.Tn[9].n13 VGND 0.14365f
C13770 XThC.Tn[9].t17 VGND 0.01585f
C13771 XThC.Tn[9].t35 VGND 0.01732f
C13772 XThC.Tn[9].n14 VGND 0.03865f
C13773 XThC.Tn[9].n15 VGND 0.02648f
C13774 XThC.Tn[9].n16 VGND 0.08716f
C13775 XThC.Tn[9].n17 VGND 0.14365f
C13776 XThC.Tn[9].t39 VGND 0.01585f
C13777 XThC.Tn[9].t24 VGND 0.01732f
C13778 XThC.Tn[9].n18 VGND 0.03865f
C13779 XThC.Tn[9].n19 VGND 0.02648f
C13780 XThC.Tn[9].n20 VGND 0.08716f
C13781 XThC.Tn[9].n21 VGND 0.14365f
C13782 XThC.Tn[9].t40 VGND 0.01585f
C13783 XThC.Tn[9].t25 VGND 0.01732f
C13784 XThC.Tn[9].n22 VGND 0.03865f
C13785 XThC.Tn[9].n23 VGND 0.02648f
C13786 XThC.Tn[9].n24 VGND 0.08716f
C13787 XThC.Tn[9].n25 VGND 0.14365f
C13788 XThC.Tn[9].t22 VGND 0.01585f
C13789 XThC.Tn[9].t38 VGND 0.01732f
C13790 XThC.Tn[9].n26 VGND 0.03865f
C13791 XThC.Tn[9].n27 VGND 0.02648f
C13792 XThC.Tn[9].n28 VGND 0.08716f
C13793 XThC.Tn[9].n29 VGND 0.14365f
C13794 XThC.Tn[9].t28 VGND 0.01585f
C13795 XThC.Tn[9].t14 VGND 0.01732f
C13796 XThC.Tn[9].n30 VGND 0.03865f
C13797 XThC.Tn[9].n31 VGND 0.02648f
C13798 XThC.Tn[9].n32 VGND 0.08716f
C13799 XThC.Tn[9].n33 VGND 0.14365f
C13800 XThC.Tn[9].t31 VGND 0.01585f
C13801 XThC.Tn[9].t16 VGND 0.01732f
C13802 XThC.Tn[9].n34 VGND 0.03865f
C13803 XThC.Tn[9].n35 VGND 0.02648f
C13804 XThC.Tn[9].n36 VGND 0.08716f
C13805 XThC.Tn[9].n37 VGND 0.14365f
C13806 XThC.Tn[9].t19 VGND 0.01585f
C13807 XThC.Tn[9].t36 VGND 0.01732f
C13808 XThC.Tn[9].n38 VGND 0.03865f
C13809 XThC.Tn[9].n39 VGND 0.02648f
C13810 XThC.Tn[9].n40 VGND 0.08716f
C13811 XThC.Tn[9].n41 VGND 0.14365f
C13812 XThC.Tn[9].t21 VGND 0.01585f
C13813 XThC.Tn[9].t37 VGND 0.01732f
C13814 XThC.Tn[9].n42 VGND 0.03865f
C13815 XThC.Tn[9].n43 VGND 0.02648f
C13816 XThC.Tn[9].n44 VGND 0.08716f
C13817 XThC.Tn[9].n45 VGND 0.14365f
C13818 XThC.Tn[9].t32 VGND 0.01585f
C13819 XThC.Tn[9].t18 VGND 0.01732f
C13820 XThC.Tn[9].n46 VGND 0.03865f
C13821 XThC.Tn[9].n47 VGND 0.02648f
C13822 XThC.Tn[9].n48 VGND 0.08716f
C13823 XThC.Tn[9].n49 VGND 0.14365f
C13824 XThC.Tn[9].t42 VGND 0.01585f
C13825 XThC.Tn[9].t27 VGND 0.01732f
C13826 XThC.Tn[9].n50 VGND 0.03865f
C13827 XThC.Tn[9].n51 VGND 0.02648f
C13828 XThC.Tn[9].n52 VGND 0.08716f
C13829 XThC.Tn[9].n53 VGND 0.14365f
C13830 XThC.Tn[9].t43 VGND 0.01585f
C13831 XThC.Tn[9].t29 VGND 0.01732f
C13832 XThC.Tn[9].n54 VGND 0.03865f
C13833 XThC.Tn[9].n55 VGND 0.02648f
C13834 XThC.Tn[9].n56 VGND 0.08716f
C13835 XThC.Tn[9].n57 VGND 0.14365f
C13836 XThC.Tn[9].t23 VGND 0.01585f
C13837 XThC.Tn[9].t41 VGND 0.01732f
C13838 XThC.Tn[9].n58 VGND 0.03865f
C13839 XThC.Tn[9].n59 VGND 0.02648f
C13840 XThC.Tn[9].n60 VGND 0.08716f
C13841 XThC.Tn[9].n61 VGND 0.14365f
C13842 XThC.Tn[9].t33 VGND 0.01585f
C13843 XThC.Tn[9].t20 VGND 0.01732f
C13844 XThC.Tn[9].n62 VGND 0.03865f
C13845 XThC.Tn[9].n63 VGND 0.02648f
C13846 XThC.Tn[9].n64 VGND 0.08716f
C13847 XThC.Tn[9].n65 VGND 0.14365f
C13848 XThC.Tn[9].n66 VGND 0.61747f
C13849 XThC.Tn[9].n67 VGND 0.26115f
C13850 XThC.Tn[9].t8 VGND 0.02f
C13851 XThC.Tn[9].t11 VGND 0.02f
C13852 XThC.Tn[9].n68 VGND 0.04321f
C13853 XThC.Tn[9].t10 VGND 0.02f
C13854 XThC.Tn[9].t9 VGND 0.02f
C13855 XThC.Tn[9].n69 VGND 0.06812f
C13856 XThC.Tn[9].n70 VGND 0.1804f
C13857 XThC.Tn[9].n71 VGND 0.01328f
C13858 XThC.Tn[9].t1 VGND 0.02f
C13859 XThC.Tn[9].t0 VGND 0.02f
C13860 XThC.Tn[9].n72 VGND 0.06073f
C13861 XThC.Tn[9].t3 VGND 0.02f
C13862 XThC.Tn[9].t2 VGND 0.02f
C13863 XThC.Tn[9].n73 VGND 0.04446f
C13864 XThC.Tn[9].n74 VGND 0.19787f
C13865 XThC.Tn[5].t7 VGND 0.01807f
C13866 XThC.Tn[5].t6 VGND 0.01807f
C13867 XThC.Tn[5].n0 VGND 0.03647f
C13868 XThC.Tn[5].t5 VGND 0.01807f
C13869 XThC.Tn[5].t4 VGND 0.01807f
C13870 XThC.Tn[5].n1 VGND 0.04267f
C13871 XThC.Tn[5].n2 VGND 0.12799f
C13872 XThC.Tn[5].t1 VGND 0.01174f
C13873 XThC.Tn[5].t0 VGND 0.01174f
C13874 XThC.Tn[5].n3 VGND 0.02674f
C13875 XThC.Tn[5].t8 VGND 0.01174f
C13876 XThC.Tn[5].t11 VGND 0.01174f
C13877 XThC.Tn[5].n4 VGND 0.04456f
C13878 XThC.Tn[5].t10 VGND 0.01174f
C13879 XThC.Tn[5].t9 VGND 0.01174f
C13880 XThC.Tn[5].n5 VGND 0.02674f
C13881 XThC.Tn[5].n6 VGND 0.12735f
C13882 XThC.Tn[5].t3 VGND 0.01174f
C13883 XThC.Tn[5].t2 VGND 0.01174f
C13884 XThC.Tn[5].n7 VGND 0.02674f
C13885 XThC.Tn[5].n8 VGND 0.07873f
C13886 XThC.Tn[5].n9 VGND 0.08885f
C13887 XThC.Tn[5].t15 VGND 0.01432f
C13888 XThC.Tn[5].t33 VGND 0.01564f
C13889 XThC.Tn[5].n10 VGND 0.03492f
C13890 XThC.Tn[5].n11 VGND 0.02392f
C13891 XThC.Tn[5].n12 VGND 0.07852f
C13892 XThC.Tn[5].t34 VGND 0.01432f
C13893 XThC.Tn[5].t19 VGND 0.01564f
C13894 XThC.Tn[5].n13 VGND 0.03492f
C13895 XThC.Tn[5].n14 VGND 0.02392f
C13896 XThC.Tn[5].n15 VGND 0.07873f
C13897 XThC.Tn[5].n16 VGND 0.12976f
C13898 XThC.Tn[5].t36 VGND 0.01432f
C13899 XThC.Tn[5].t23 VGND 0.01564f
C13900 XThC.Tn[5].n17 VGND 0.03492f
C13901 XThC.Tn[5].n18 VGND 0.02392f
C13902 XThC.Tn[5].n19 VGND 0.07873f
C13903 XThC.Tn[5].n20 VGND 0.12976f
C13904 XThC.Tn[5].t38 VGND 0.01432f
C13905 XThC.Tn[5].t24 VGND 0.01564f
C13906 XThC.Tn[5].n21 VGND 0.03492f
C13907 XThC.Tn[5].n22 VGND 0.02392f
C13908 XThC.Tn[5].n23 VGND 0.07873f
C13909 XThC.Tn[5].n24 VGND 0.12976f
C13910 XThC.Tn[5].t28 VGND 0.01432f
C13911 XThC.Tn[5].t13 VGND 0.01564f
C13912 XThC.Tn[5].n25 VGND 0.03492f
C13913 XThC.Tn[5].n26 VGND 0.02392f
C13914 XThC.Tn[5].n27 VGND 0.07873f
C13915 XThC.Tn[5].n28 VGND 0.12976f
C13916 XThC.Tn[5].t29 VGND 0.01432f
C13917 XThC.Tn[5].t14 VGND 0.01564f
C13918 XThC.Tn[5].n29 VGND 0.03492f
C13919 XThC.Tn[5].n30 VGND 0.02392f
C13920 XThC.Tn[5].n31 VGND 0.07873f
C13921 XThC.Tn[5].n32 VGND 0.12976f
C13922 XThC.Tn[5].t43 VGND 0.01432f
C13923 XThC.Tn[5].t27 VGND 0.01564f
C13924 XThC.Tn[5].n33 VGND 0.03492f
C13925 XThC.Tn[5].n34 VGND 0.02392f
C13926 XThC.Tn[5].n35 VGND 0.07873f
C13927 XThC.Tn[5].n36 VGND 0.12976f
C13928 XThC.Tn[5].t17 VGND 0.01432f
C13929 XThC.Tn[5].t35 VGND 0.01564f
C13930 XThC.Tn[5].n37 VGND 0.03492f
C13931 XThC.Tn[5].n38 VGND 0.02392f
C13932 XThC.Tn[5].n39 VGND 0.07873f
C13933 XThC.Tn[5].n40 VGND 0.12976f
C13934 XThC.Tn[5].t20 VGND 0.01432f
C13935 XThC.Tn[5].t37 VGND 0.01564f
C13936 XThC.Tn[5].n41 VGND 0.03492f
C13937 XThC.Tn[5].n42 VGND 0.02392f
C13938 XThC.Tn[5].n43 VGND 0.07873f
C13939 XThC.Tn[5].n44 VGND 0.12976f
C13940 XThC.Tn[5].t40 VGND 0.01432f
C13941 XThC.Tn[5].t25 VGND 0.01564f
C13942 XThC.Tn[5].n45 VGND 0.03492f
C13943 XThC.Tn[5].n46 VGND 0.02392f
C13944 XThC.Tn[5].n47 VGND 0.07873f
C13945 XThC.Tn[5].n48 VGND 0.12976f
C13946 XThC.Tn[5].t42 VGND 0.01432f
C13947 XThC.Tn[5].t26 VGND 0.01564f
C13948 XThC.Tn[5].n49 VGND 0.03492f
C13949 XThC.Tn[5].n50 VGND 0.02392f
C13950 XThC.Tn[5].n51 VGND 0.07873f
C13951 XThC.Tn[5].n52 VGND 0.12976f
C13952 XThC.Tn[5].t21 VGND 0.01432f
C13953 XThC.Tn[5].t39 VGND 0.01564f
C13954 XThC.Tn[5].n53 VGND 0.03492f
C13955 XThC.Tn[5].n54 VGND 0.02392f
C13956 XThC.Tn[5].n55 VGND 0.07873f
C13957 XThC.Tn[5].n56 VGND 0.12976f
C13958 XThC.Tn[5].t31 VGND 0.01432f
C13959 XThC.Tn[5].t16 VGND 0.01564f
C13960 XThC.Tn[5].n57 VGND 0.03492f
C13961 XThC.Tn[5].n58 VGND 0.02392f
C13962 XThC.Tn[5].n59 VGND 0.07873f
C13963 XThC.Tn[5].n60 VGND 0.12976f
C13964 XThC.Tn[5].t32 VGND 0.01432f
C13965 XThC.Tn[5].t18 VGND 0.01564f
C13966 XThC.Tn[5].n61 VGND 0.03492f
C13967 XThC.Tn[5].n62 VGND 0.02392f
C13968 XThC.Tn[5].n63 VGND 0.07873f
C13969 XThC.Tn[5].n64 VGND 0.12976f
C13970 XThC.Tn[5].t12 VGND 0.01432f
C13971 XThC.Tn[5].t30 VGND 0.01564f
C13972 XThC.Tn[5].n65 VGND 0.03492f
C13973 XThC.Tn[5].n66 VGND 0.02392f
C13974 XThC.Tn[5].n67 VGND 0.07873f
C13975 XThC.Tn[5].n68 VGND 0.12976f
C13976 XThC.Tn[5].t22 VGND 0.01432f
C13977 XThC.Tn[5].t41 VGND 0.01564f
C13978 XThC.Tn[5].n69 VGND 0.03492f
C13979 XThC.Tn[5].n70 VGND 0.02392f
C13980 XThC.Tn[5].n71 VGND 0.07873f
C13981 XThC.Tn[5].n72 VGND 0.12976f
C13982 XThC.Tn[5].n73 VGND 0.14766f
C13983 XThR.Tn[9].t2 VGND 0.02425f
C13984 XThR.Tn[9].t0 VGND 0.02425f
C13985 XThR.Tn[9].n0 VGND 0.07362f
C13986 XThR.Tn[9].t3 VGND 0.02425f
C13987 XThR.Tn[9].t1 VGND 0.02425f
C13988 XThR.Tn[9].n1 VGND 0.0539f
C13989 XThR.Tn[9].n2 VGND 0.24507f
C13990 XThR.Tn[9].t5 VGND 0.01576f
C13991 XThR.Tn[9].t7 VGND 0.01576f
C13992 XThR.Tn[9].n3 VGND 0.03931f
C13993 XThR.Tn[9].t4 VGND 0.01576f
C13994 XThR.Tn[9].t6 VGND 0.01576f
C13995 XThR.Tn[9].n4 VGND 0.03152f
C13996 XThR.Tn[9].n5 VGND 0.07929f
C13997 XThR.Tn[9].t17 VGND 0.01895f
C13998 XThR.Tn[9].t71 VGND 0.02075f
C13999 XThR.Tn[9].n6 VGND 0.05067f
C14000 XThR.Tn[9].n7 VGND 0.09733f
C14001 XThR.Tn[9].t35 VGND 0.01895f
C14002 XThR.Tn[9].t28 VGND 0.02075f
C14003 XThR.Tn[9].n8 VGND 0.05067f
C14004 XThR.Tn[9].t50 VGND 0.01889f
C14005 XThR.Tn[9].t19 VGND 0.02068f
C14006 XThR.Tn[9].n9 VGND 0.05272f
C14007 XThR.Tn[9].n10 VGND 0.03704f
C14008 XThR.Tn[9].n11 VGND 0.00677f
C14009 XThR.Tn[9].n12 VGND 0.11885f
C14010 XThR.Tn[9].t72 VGND 0.01895f
C14011 XThR.Tn[9].t64 VGND 0.02075f
C14012 XThR.Tn[9].n13 VGND 0.05067f
C14013 XThR.Tn[9].t26 VGND 0.01889f
C14014 XThR.Tn[9].t59 VGND 0.02068f
C14015 XThR.Tn[9].n14 VGND 0.05272f
C14016 XThR.Tn[9].n15 VGND 0.03704f
C14017 XThR.Tn[9].n16 VGND 0.00677f
C14018 XThR.Tn[9].n17 VGND 0.11885f
C14019 XThR.Tn[9].t29 VGND 0.01895f
C14020 XThR.Tn[9].t21 VGND 0.02075f
C14021 XThR.Tn[9].n18 VGND 0.05067f
C14022 XThR.Tn[9].t41 VGND 0.01889f
C14023 XThR.Tn[9].t15 VGND 0.02068f
C14024 XThR.Tn[9].n19 VGND 0.05272f
C14025 XThR.Tn[9].n20 VGND 0.03704f
C14026 XThR.Tn[9].n21 VGND 0.00677f
C14027 XThR.Tn[9].n22 VGND 0.11885f
C14028 XThR.Tn[9].t56 VGND 0.01895f
C14029 XThR.Tn[9].t46 VGND 0.02075f
C14030 XThR.Tn[9].n23 VGND 0.05067f
C14031 XThR.Tn[9].t73 VGND 0.01889f
C14032 XThR.Tn[9].t42 VGND 0.02068f
C14033 XThR.Tn[9].n24 VGND 0.05272f
C14034 XThR.Tn[9].n25 VGND 0.03704f
C14035 XThR.Tn[9].n26 VGND 0.00677f
C14036 XThR.Tn[9].n27 VGND 0.11885f
C14037 XThR.Tn[9].t31 VGND 0.01895f
C14038 XThR.Tn[9].t23 VGND 0.02075f
C14039 XThR.Tn[9].n28 VGND 0.05067f
C14040 XThR.Tn[9].t44 VGND 0.01889f
C14041 XThR.Tn[9].t16 VGND 0.02068f
C14042 XThR.Tn[9].n29 VGND 0.05272f
C14043 XThR.Tn[9].n30 VGND 0.03704f
C14044 XThR.Tn[9].n31 VGND 0.00677f
C14045 XThR.Tn[9].n32 VGND 0.11885f
C14046 XThR.Tn[9].t67 VGND 0.01895f
C14047 XThR.Tn[9].t37 VGND 0.02075f
C14048 XThR.Tn[9].n33 VGND 0.05067f
C14049 XThR.Tn[9].t20 VGND 0.01889f
C14050 XThR.Tn[9].t33 VGND 0.02068f
C14051 XThR.Tn[9].n34 VGND 0.05272f
C14052 XThR.Tn[9].n35 VGND 0.03704f
C14053 XThR.Tn[9].n36 VGND 0.00677f
C14054 XThR.Tn[9].n37 VGND 0.11885f
C14055 XThR.Tn[9].t36 VGND 0.01895f
C14056 XThR.Tn[9].t32 VGND 0.02075f
C14057 XThR.Tn[9].n38 VGND 0.05067f
C14058 XThR.Tn[9].t51 VGND 0.01889f
C14059 XThR.Tn[9].t25 VGND 0.02068f
C14060 XThR.Tn[9].n39 VGND 0.05272f
C14061 XThR.Tn[9].n40 VGND 0.03704f
C14062 XThR.Tn[9].n41 VGND 0.00677f
C14063 XThR.Tn[9].n42 VGND 0.11885f
C14064 XThR.Tn[9].t39 VGND 0.01895f
C14065 XThR.Tn[9].t45 VGND 0.02075f
C14066 XThR.Tn[9].n43 VGND 0.05067f
C14067 XThR.Tn[9].t55 VGND 0.01889f
C14068 XThR.Tn[9].t40 VGND 0.02068f
C14069 XThR.Tn[9].n44 VGND 0.05272f
C14070 XThR.Tn[9].n45 VGND 0.03704f
C14071 XThR.Tn[9].n46 VGND 0.00677f
C14072 XThR.Tn[9].n47 VGND 0.11885f
C14073 XThR.Tn[9].t58 VGND 0.01895f
C14074 XThR.Tn[9].t66 VGND 0.02075f
C14075 XThR.Tn[9].n48 VGND 0.05067f
C14076 XThR.Tn[9].t13 VGND 0.01889f
C14077 XThR.Tn[9].t60 VGND 0.02068f
C14078 XThR.Tn[9].n49 VGND 0.05272f
C14079 XThR.Tn[9].n50 VGND 0.03704f
C14080 XThR.Tn[9].n51 VGND 0.00677f
C14081 XThR.Tn[9].n52 VGND 0.11885f
C14082 XThR.Tn[9].t48 VGND 0.01895f
C14083 XThR.Tn[9].t24 VGND 0.02075f
C14084 XThR.Tn[9].n53 VGND 0.05067f
C14085 XThR.Tn[9].t65 VGND 0.01889f
C14086 XThR.Tn[9].t18 VGND 0.02068f
C14087 XThR.Tn[9].n54 VGND 0.05272f
C14088 XThR.Tn[9].n55 VGND 0.03704f
C14089 XThR.Tn[9].n56 VGND 0.00677f
C14090 XThR.Tn[9].n57 VGND 0.11885f
C14091 XThR.Tn[9].t70 VGND 0.01895f
C14092 XThR.Tn[9].t62 VGND 0.02075f
C14093 XThR.Tn[9].n58 VGND 0.05067f
C14094 XThR.Tn[9].t22 VGND 0.01889f
C14095 XThR.Tn[9].t52 VGND 0.02068f
C14096 XThR.Tn[9].n59 VGND 0.05272f
C14097 XThR.Tn[9].n60 VGND 0.03704f
C14098 XThR.Tn[9].n61 VGND 0.00677f
C14099 XThR.Tn[9].n62 VGND 0.11885f
C14100 XThR.Tn[9].t38 VGND 0.01895f
C14101 XThR.Tn[9].t34 VGND 0.02075f
C14102 XThR.Tn[9].n63 VGND 0.05067f
C14103 XThR.Tn[9].t53 VGND 0.01889f
C14104 XThR.Tn[9].t27 VGND 0.02068f
C14105 XThR.Tn[9].n64 VGND 0.05272f
C14106 XThR.Tn[9].n65 VGND 0.03704f
C14107 XThR.Tn[9].n66 VGND 0.00677f
C14108 XThR.Tn[9].n67 VGND 0.11885f
C14109 XThR.Tn[9].t57 VGND 0.01895f
C14110 XThR.Tn[9].t47 VGND 0.02075f
C14111 XThR.Tn[9].n68 VGND 0.05067f
C14112 XThR.Tn[9].t12 VGND 0.01889f
C14113 XThR.Tn[9].t43 VGND 0.02068f
C14114 XThR.Tn[9].n69 VGND 0.05272f
C14115 XThR.Tn[9].n70 VGND 0.03704f
C14116 XThR.Tn[9].n71 VGND 0.00677f
C14117 XThR.Tn[9].n72 VGND 0.11885f
C14118 XThR.Tn[9].t14 VGND 0.01895f
C14119 XThR.Tn[9].t69 VGND 0.02075f
C14120 XThR.Tn[9].n73 VGND 0.05067f
C14121 XThR.Tn[9].t30 VGND 0.01889f
C14122 XThR.Tn[9].t61 VGND 0.02068f
C14123 XThR.Tn[9].n74 VGND 0.05272f
C14124 XThR.Tn[9].n75 VGND 0.03704f
C14125 XThR.Tn[9].n76 VGND 0.00677f
C14126 XThR.Tn[9].n77 VGND 0.11885f
C14127 XThR.Tn[9].t49 VGND 0.01895f
C14128 XThR.Tn[9].t63 VGND 0.02075f
C14129 XThR.Tn[9].n78 VGND 0.05067f
C14130 XThR.Tn[9].t68 VGND 0.01889f
C14131 XThR.Tn[9].t54 VGND 0.02068f
C14132 XThR.Tn[9].n79 VGND 0.05272f
C14133 XThR.Tn[9].n80 VGND 0.03704f
C14134 XThR.Tn[9].n81 VGND 0.00677f
C14135 XThR.Tn[9].n82 VGND 0.11885f
C14136 XThR.Tn[9].n83 VGND 0.10801f
C14137 XThR.Tn[9].n84 VGND 0.35039f
C14138 XThR.Tn[9].t10 VGND 0.02425f
C14139 XThR.Tn[9].t8 VGND 0.02425f
C14140 XThR.Tn[9].n85 VGND 0.05239f
C14141 XThR.Tn[9].t11 VGND 0.02425f
C14142 XThR.Tn[9].t9 VGND 0.02425f
C14143 XThR.Tn[9].n86 VGND 0.07973f
C14144 XThR.Tn[9].n87 VGND 0.22139f
C14145 XThR.Tn[9].n88 VGND 0.02964f
C14146 XThC.Tn[6].t11 VGND 0.01183f
C14147 XThC.Tn[6].t10 VGND 0.01183f
C14148 XThC.Tn[6].n0 VGND 0.04489f
C14149 XThC.Tn[6].t9 VGND 0.01183f
C14150 XThC.Tn[6].t8 VGND 0.01183f
C14151 XThC.Tn[6].n1 VGND 0.02694f
C14152 XThC.Tn[6].n2 VGND 0.12829f
C14153 XThC.Tn[6].t6 VGND 0.01183f
C14154 XThC.Tn[6].t5 VGND 0.01183f
C14155 XThC.Tn[6].n3 VGND 0.02694f
C14156 XThC.Tn[6].n4 VGND 0.07931f
C14157 XThC.Tn[6].t4 VGND 0.01183f
C14158 XThC.Tn[6].t7 VGND 0.01183f
C14159 XThC.Tn[6].n5 VGND 0.02694f
C14160 XThC.Tn[6].n6 VGND 0.0895f
C14161 XThC.Tn[6].t23 VGND 0.01443f
C14162 XThC.Tn[6].t26 VGND 0.01576f
C14163 XThC.Tn[6].n7 VGND 0.03517f
C14164 XThC.Tn[6].n8 VGND 0.0241f
C14165 XThC.Tn[6].n9 VGND 0.0791f
C14166 XThC.Tn[6].t40 VGND 0.01443f
C14167 XThC.Tn[6].t13 VGND 0.01576f
C14168 XThC.Tn[6].n10 VGND 0.03517f
C14169 XThC.Tn[6].n11 VGND 0.0241f
C14170 XThC.Tn[6].n12 VGND 0.07932f
C14171 XThC.Tn[6].n13 VGND 0.13072f
C14172 XThC.Tn[6].t42 VGND 0.01443f
C14173 XThC.Tn[6].t17 VGND 0.01576f
C14174 XThC.Tn[6].n14 VGND 0.03517f
C14175 XThC.Tn[6].n15 VGND 0.0241f
C14176 XThC.Tn[6].n16 VGND 0.07932f
C14177 XThC.Tn[6].n17 VGND 0.13072f
C14178 XThC.Tn[6].t12 VGND 0.01443f
C14179 XThC.Tn[6].t18 VGND 0.01576f
C14180 XThC.Tn[6].n18 VGND 0.03517f
C14181 XThC.Tn[6].n19 VGND 0.0241f
C14182 XThC.Tn[6].n20 VGND 0.07932f
C14183 XThC.Tn[6].n21 VGND 0.13072f
C14184 XThC.Tn[6].t33 VGND 0.01443f
C14185 XThC.Tn[6].t37 VGND 0.01576f
C14186 XThC.Tn[6].n22 VGND 0.03517f
C14187 XThC.Tn[6].n23 VGND 0.0241f
C14188 XThC.Tn[6].n24 VGND 0.07932f
C14189 XThC.Tn[6].n25 VGND 0.13072f
C14190 XThC.Tn[6].t35 VGND 0.01443f
C14191 XThC.Tn[6].t38 VGND 0.01576f
C14192 XThC.Tn[6].n26 VGND 0.03517f
C14193 XThC.Tn[6].n27 VGND 0.0241f
C14194 XThC.Tn[6].n28 VGND 0.07932f
C14195 XThC.Tn[6].n29 VGND 0.13072f
C14196 XThC.Tn[6].t16 VGND 0.01443f
C14197 XThC.Tn[6].t22 VGND 0.01576f
C14198 XThC.Tn[6].n30 VGND 0.03517f
C14199 XThC.Tn[6].n31 VGND 0.0241f
C14200 XThC.Tn[6].n32 VGND 0.07932f
C14201 XThC.Tn[6].n33 VGND 0.13072f
C14202 XThC.Tn[6].t25 VGND 0.01443f
C14203 XThC.Tn[6].t29 VGND 0.01576f
C14204 XThC.Tn[6].n34 VGND 0.03517f
C14205 XThC.Tn[6].n35 VGND 0.0241f
C14206 XThC.Tn[6].n36 VGND 0.07932f
C14207 XThC.Tn[6].n37 VGND 0.13072f
C14208 XThC.Tn[6].t27 VGND 0.01443f
C14209 XThC.Tn[6].t31 VGND 0.01576f
C14210 XThC.Tn[6].n38 VGND 0.03517f
C14211 XThC.Tn[6].n39 VGND 0.0241f
C14212 XThC.Tn[6].n40 VGND 0.07932f
C14213 XThC.Tn[6].n41 VGND 0.13072f
C14214 XThC.Tn[6].t14 VGND 0.01443f
C14215 XThC.Tn[6].t19 VGND 0.01576f
C14216 XThC.Tn[6].n42 VGND 0.03517f
C14217 XThC.Tn[6].n43 VGND 0.0241f
C14218 XThC.Tn[6].n44 VGND 0.07932f
C14219 XThC.Tn[6].n45 VGND 0.13072f
C14220 XThC.Tn[6].t15 VGND 0.01443f
C14221 XThC.Tn[6].t21 VGND 0.01576f
C14222 XThC.Tn[6].n46 VGND 0.03517f
C14223 XThC.Tn[6].n47 VGND 0.0241f
C14224 XThC.Tn[6].n48 VGND 0.07932f
C14225 XThC.Tn[6].n49 VGND 0.13072f
C14226 XThC.Tn[6].t28 VGND 0.01443f
C14227 XThC.Tn[6].t32 VGND 0.01576f
C14228 XThC.Tn[6].n50 VGND 0.03517f
C14229 XThC.Tn[6].n51 VGND 0.0241f
C14230 XThC.Tn[6].n52 VGND 0.07932f
C14231 XThC.Tn[6].n53 VGND 0.13072f
C14232 XThC.Tn[6].t36 VGND 0.01443f
C14233 XThC.Tn[6].t41 VGND 0.01576f
C14234 XThC.Tn[6].n54 VGND 0.03517f
C14235 XThC.Tn[6].n55 VGND 0.0241f
C14236 XThC.Tn[6].n56 VGND 0.07932f
C14237 XThC.Tn[6].n57 VGND 0.13072f
C14238 XThC.Tn[6].t39 VGND 0.01443f
C14239 XThC.Tn[6].t43 VGND 0.01576f
C14240 XThC.Tn[6].n58 VGND 0.03517f
C14241 XThC.Tn[6].n59 VGND 0.0241f
C14242 XThC.Tn[6].n60 VGND 0.07932f
C14243 XThC.Tn[6].n61 VGND 0.13072f
C14244 XThC.Tn[6].t20 VGND 0.01443f
C14245 XThC.Tn[6].t24 VGND 0.01576f
C14246 XThC.Tn[6].n62 VGND 0.03517f
C14247 XThC.Tn[6].n63 VGND 0.0241f
C14248 XThC.Tn[6].n64 VGND 0.07932f
C14249 XThC.Tn[6].n65 VGND 0.13072f
C14250 XThC.Tn[6].t30 VGND 0.01443f
C14251 XThC.Tn[6].t34 VGND 0.01576f
C14252 XThC.Tn[6].n66 VGND 0.03517f
C14253 XThC.Tn[6].n67 VGND 0.0241f
C14254 XThC.Tn[6].n68 VGND 0.07932f
C14255 XThC.Tn[6].n69 VGND 0.13072f
C14256 XThC.Tn[6].n70 VGND 0.14537f
C14257 XThC.Tn[6].t1 VGND 0.0182f
C14258 XThC.Tn[6].t0 VGND 0.0182f
C14259 XThC.Tn[6].n71 VGND 0.04298f
C14260 XThC.Tn[6].t3 VGND 0.0182f
C14261 XThC.Tn[6].t2 VGND 0.0182f
C14262 XThC.Tn[6].n72 VGND 0.03674f
C14263 XThC.Tn[6].n73 VGND 0.12033f
C14264 XThC.Tn[6].n74 VGND 0.03808f
C14265 XThC.XTBN.Y.n0 VGND 0.01531f
C14266 XThC.XTBN.Y.t50 VGND 0.01024f
C14267 XThC.XTBN.Y.t118 VGND 0.00603f
C14268 XThC.XTBN.Y.t18 VGND 0.01024f
C14269 XThC.XTBN.Y.t83 VGND 0.00603f
C14270 XThC.XTBN.Y.n1 VGND 0.01477f
C14271 XThC.XTBN.Y.n2 VGND 0.00524f
C14272 XThC.XTBN.Y.t120 VGND 0.01024f
C14273 XThC.XTBN.Y.t71 VGND 0.00603f
C14274 XThC.XTBN.Y.t114 VGND 0.01024f
C14275 XThC.XTBN.Y.t62 VGND 0.00603f
C14276 XThC.XTBN.Y.n3 VGND 0.0138f
C14277 XThC.XTBN.Y.n4 VGND 0.00676f
C14278 XThC.XTBN.Y.n5 VGND 0.01477f
C14279 XThC.XTBN.Y.n6 VGND 0.00676f
C14280 XThC.XTBN.Y.n7 VGND 0.00548f
C14281 XThC.XTBN.Y.n8 VGND 0.00561f
C14282 XThC.XTBN.Y.n9 VGND 0.00676f
C14283 XThC.XTBN.Y.n10 VGND 0.02164f
C14284 XThC.XTBN.Y.n11 VGND 0.00584f
C14285 XThC.XTBN.Y.n12 VGND 0.00877f
C14286 XThC.XTBN.Y.t121 VGND 0.00603f
C14287 XThC.XTBN.Y.t79 VGND 0.01024f
C14288 XThC.XTBN.Y.t84 VGND 0.00603f
C14289 XThC.XTBN.Y.t36 VGND 0.01024f
C14290 XThC.XTBN.Y.n13 VGND 0.01477f
C14291 XThC.XTBN.Y.n14 VGND 0.00524f
C14292 XThC.XTBN.Y.t73 VGND 0.00603f
C14293 XThC.XTBN.Y.t26 VGND 0.01024f
C14294 XThC.XTBN.Y.t64 VGND 0.00603f
C14295 XThC.XTBN.Y.t21 VGND 0.01024f
C14296 XThC.XTBN.Y.n15 VGND 0.0138f
C14297 XThC.XTBN.Y.n16 VGND 0.00676f
C14298 XThC.XTBN.Y.n17 VGND 0.01477f
C14299 XThC.XTBN.Y.n18 VGND 0.00676f
C14300 XThC.XTBN.Y.n19 VGND 0.00548f
C14301 XThC.XTBN.Y.n20 VGND 0.00561f
C14302 XThC.XTBN.Y.n21 VGND 0.00676f
C14303 XThC.XTBN.Y.n22 VGND 0.02164f
C14304 XThC.XTBN.Y.n23 VGND 0.00584f
C14305 XThC.XTBN.Y.n24 VGND 0.00417f
C14306 XThC.XTBN.Y.n25 VGND 0.11789f
C14307 XThC.XTBN.Y.t106 VGND 0.01024f
C14308 XThC.XTBN.Y.t89 VGND 0.00603f
C14309 XThC.XTBN.Y.t70 VGND 0.01024f
C14310 XThC.XTBN.Y.t41 VGND 0.00603f
C14311 XThC.XTBN.Y.n26 VGND 0.01477f
C14312 XThC.XTBN.Y.n27 VGND 0.00524f
C14313 XThC.XTBN.Y.t56 VGND 0.01024f
C14314 XThC.XTBN.Y.t35 VGND 0.00603f
C14315 XThC.XTBN.Y.t48 VGND 0.01024f
C14316 XThC.XTBN.Y.t32 VGND 0.00603f
C14317 XThC.XTBN.Y.n28 VGND 0.0138f
C14318 XThC.XTBN.Y.n29 VGND 0.00676f
C14319 XThC.XTBN.Y.n30 VGND 0.01477f
C14320 XThC.XTBN.Y.n31 VGND 0.00676f
C14321 XThC.XTBN.Y.n32 VGND 0.00548f
C14322 XThC.XTBN.Y.n33 VGND 0.00561f
C14323 XThC.XTBN.Y.n34 VGND 0.00676f
C14324 XThC.XTBN.Y.n35 VGND 0.02164f
C14325 XThC.XTBN.Y.n36 VGND 0.00584f
C14326 XThC.XTBN.Y.n37 VGND 0.00417f
C14327 XThC.XTBN.Y.n38 VGND 0.07443f
C14328 XThC.XTBN.Y.t43 VGND 0.00603f
C14329 XThC.XTBN.Y.t39 VGND 0.01024f
C14330 XThC.XTBN.Y.t10 VGND 0.00603f
C14331 XThC.XTBN.Y.t122 VGND 0.01024f
C14332 XThC.XTBN.Y.n39 VGND 0.01477f
C14333 XThC.XTBN.Y.n40 VGND 0.00524f
C14334 XThC.XTBN.Y.t112 VGND 0.00603f
C14335 XThC.XTBN.Y.t109 VGND 0.01024f
C14336 XThC.XTBN.Y.t108 VGND 0.00603f
C14337 XThC.XTBN.Y.t102 VGND 0.01024f
C14338 XThC.XTBN.Y.n41 VGND 0.0138f
C14339 XThC.XTBN.Y.n42 VGND 0.00676f
C14340 XThC.XTBN.Y.n43 VGND 0.01477f
C14341 XThC.XTBN.Y.n44 VGND 0.00676f
C14342 XThC.XTBN.Y.n45 VGND 0.00548f
C14343 XThC.XTBN.Y.n46 VGND 0.00561f
C14344 XThC.XTBN.Y.n47 VGND 0.00676f
C14345 XThC.XTBN.Y.n48 VGND 0.02164f
C14346 XThC.XTBN.Y.n49 VGND 0.00584f
C14347 XThC.XTBN.Y.n50 VGND 0.00417f
C14348 XThC.XTBN.Y.n51 VGND 0.07443f
C14349 XThC.XTBN.Y.t47 VGND 0.01024f
C14350 XThC.XTBN.Y.t31 VGND 0.00603f
C14351 XThC.XTBN.Y.t17 VGND 0.01024f
C14352 XThC.XTBN.Y.t104 VGND 0.00603f
C14353 XThC.XTBN.Y.n52 VGND 0.01477f
C14354 XThC.XTBN.Y.n53 VGND 0.00524f
C14355 XThC.XTBN.Y.t116 VGND 0.01024f
C14356 XThC.XTBN.Y.t94 VGND 0.00603f
C14357 XThC.XTBN.Y.t111 VGND 0.01024f
C14358 XThC.XTBN.Y.t92 VGND 0.00603f
C14359 XThC.XTBN.Y.n54 VGND 0.0138f
C14360 XThC.XTBN.Y.n55 VGND 0.00676f
C14361 XThC.XTBN.Y.n56 VGND 0.01477f
C14362 XThC.XTBN.Y.n57 VGND 0.00676f
C14363 XThC.XTBN.Y.n58 VGND 0.00548f
C14364 XThC.XTBN.Y.n59 VGND 0.00561f
C14365 XThC.XTBN.Y.n60 VGND 0.00676f
C14366 XThC.XTBN.Y.n61 VGND 0.02164f
C14367 XThC.XTBN.Y.n62 VGND 0.00584f
C14368 XThC.XTBN.Y.n63 VGND 0.00417f
C14369 XThC.XTBN.Y.n64 VGND 0.07443f
C14370 XThC.XTBN.Y.t107 VGND 0.00603f
C14371 XThC.XTBN.Y.t101 VGND 0.01024f
C14372 XThC.XTBN.Y.t72 VGND 0.00603f
C14373 XThC.XTBN.Y.t63 VGND 0.01024f
C14374 XThC.XTBN.Y.n65 VGND 0.01477f
C14375 XThC.XTBN.Y.n66 VGND 0.00524f
C14376 XThC.XTBN.Y.t57 VGND 0.00603f
C14377 XThC.XTBN.Y.t52 VGND 0.01024f
C14378 XThC.XTBN.Y.t49 VGND 0.00603f
C14379 XThC.XTBN.Y.t44 VGND 0.01024f
C14380 XThC.XTBN.Y.n67 VGND 0.0138f
C14381 XThC.XTBN.Y.n68 VGND 0.00676f
C14382 XThC.XTBN.Y.n69 VGND 0.01477f
C14383 XThC.XTBN.Y.n70 VGND 0.00676f
C14384 XThC.XTBN.Y.n71 VGND 0.00548f
C14385 XThC.XTBN.Y.n72 VGND 0.00561f
C14386 XThC.XTBN.Y.n73 VGND 0.00676f
C14387 XThC.XTBN.Y.n74 VGND 0.02164f
C14388 XThC.XTBN.Y.n75 VGND 0.00584f
C14389 XThC.XTBN.Y.n76 VGND 0.00417f
C14390 XThC.XTBN.Y.n77 VGND 0.07443f
C14391 XThC.XTBN.Y.t25 VGND 0.01024f
C14392 XThC.XTBN.Y.t123 VGND 0.00603f
C14393 XThC.XTBN.Y.t100 VGND 0.01024f
C14394 XThC.XTBN.Y.t85 VGND 0.00603f
C14395 XThC.XTBN.Y.n78 VGND 0.01477f
C14396 XThC.XTBN.Y.n79 VGND 0.00524f
C14397 XThC.XTBN.Y.t93 VGND 0.01024f
C14398 XThC.XTBN.Y.t74 VGND 0.00603f
C14399 XThC.XTBN.Y.t90 VGND 0.01024f
C14400 XThC.XTBN.Y.t65 VGND 0.00603f
C14401 XThC.XTBN.Y.n80 VGND 0.0138f
C14402 XThC.XTBN.Y.n81 VGND 0.00676f
C14403 XThC.XTBN.Y.n82 VGND 0.01477f
C14404 XThC.XTBN.Y.n83 VGND 0.00676f
C14405 XThC.XTBN.Y.n84 VGND 0.00548f
C14406 XThC.XTBN.Y.n85 VGND 0.00561f
C14407 XThC.XTBN.Y.n86 VGND 0.00676f
C14408 XThC.XTBN.Y.n87 VGND 0.02164f
C14409 XThC.XTBN.Y.n88 VGND 0.00584f
C14410 XThC.XTBN.Y.n89 VGND 0.00417f
C14411 XThC.XTBN.Y.n90 VGND 0.06646f
C14412 XThC.XTBN.Y.t46 VGND 0.01024f
C14413 XThC.XTBN.Y.t67 VGND 0.00603f
C14414 XThC.XTBN.Y.n91 VGND 0.00619f
C14415 XThC.XTBN.Y.t6 VGND 0.01024f
C14416 XThC.XTBN.Y.t24 VGND 0.00603f
C14417 XThC.XTBN.Y.n92 VGND 0.01243f
C14418 XThC.XTBN.Y.t12 VGND 0.01024f
C14419 XThC.XTBN.Y.t29 VGND 0.00603f
C14420 XThC.XTBN.Y.n93 VGND 0.01348f
C14421 XThC.XTBN.Y.n94 VGND 0.0076f
C14422 XThC.XTBN.Y.n95 VGND 0.01252f
C14423 XThC.XTBN.Y.n96 VGND 0.00434f
C14424 XThC.XTBN.Y.n97 VGND 0.00603f
C14425 XThC.XTBN.Y.n98 VGND 0.01348f
C14426 XThC.XTBN.Y.t54 VGND 0.01024f
C14427 XThC.XTBN.Y.t76 VGND 0.00603f
C14428 XThC.XTBN.Y.n99 VGND 0.01227f
C14429 XThC.XTBN.Y.n100 VGND 0.00676f
C14430 XThC.XTBN.Y.n101 VGND 0.01009f
C14431 XThC.XTBN.Y.t55 VGND 0.00603f
C14432 XThC.XTBN.Y.t38 VGND 0.01024f
C14433 XThC.XTBN.Y.n102 VGND 0.00619f
C14434 XThC.XTBN.Y.t16 VGND 0.00603f
C14435 XThC.XTBN.Y.t113 VGND 0.01024f
C14436 XThC.XTBN.Y.n103 VGND 0.01243f
C14437 XThC.XTBN.Y.t19 VGND 0.00603f
C14438 XThC.XTBN.Y.t119 VGND 0.01024f
C14439 XThC.XTBN.Y.n104 VGND 0.01348f
C14440 XThC.XTBN.Y.n105 VGND 0.0076f
C14441 XThC.XTBN.Y.n106 VGND 0.01252f
C14442 XThC.XTBN.Y.n107 VGND 0.00434f
C14443 XThC.XTBN.Y.n108 VGND 0.00603f
C14444 XThC.XTBN.Y.n109 VGND 0.01348f
C14445 XThC.XTBN.Y.t59 VGND 0.00603f
C14446 XThC.XTBN.Y.t42 VGND 0.01024f
C14447 XThC.XTBN.Y.n110 VGND 0.01227f
C14448 XThC.XTBN.Y.n111 VGND 0.00676f
C14449 XThC.XTBN.Y.n112 VGND 0.00747f
C14450 XThC.XTBN.Y.n113 VGND 0.11256f
C14451 XThC.XTBN.Y.t30 VGND 0.01024f
C14452 XThC.XTBN.Y.t8 VGND 0.00603f
C14453 XThC.XTBN.Y.n114 VGND 0.00619f
C14454 XThC.XTBN.Y.t98 VGND 0.01024f
C14455 XThC.XTBN.Y.t82 VGND 0.00603f
C14456 XThC.XTBN.Y.n115 VGND 0.01243f
C14457 XThC.XTBN.Y.t103 VGND 0.01024f
C14458 XThC.XTBN.Y.t87 VGND 0.00603f
C14459 XThC.XTBN.Y.n116 VGND 0.01348f
C14460 XThC.XTBN.Y.n117 VGND 0.0076f
C14461 XThC.XTBN.Y.n118 VGND 0.01252f
C14462 XThC.XTBN.Y.n119 VGND 0.00434f
C14463 XThC.XTBN.Y.n120 VGND 0.00603f
C14464 XThC.XTBN.Y.n121 VGND 0.01348f
C14465 XThC.XTBN.Y.t34 VGND 0.01024f
C14466 XThC.XTBN.Y.t15 VGND 0.00603f
C14467 XThC.XTBN.Y.n122 VGND 0.01227f
C14468 XThC.XTBN.Y.n123 VGND 0.00676f
C14469 XThC.XTBN.Y.n124 VGND 0.00747f
C14470 XThC.XTBN.Y.n125 VGND 0.07521f
C14471 XThC.XTBN.Y.t110 VGND 0.00603f
C14472 XThC.XTBN.Y.t96 VGND 0.01024f
C14473 XThC.XTBN.Y.n126 VGND 0.00619f
C14474 XThC.XTBN.Y.t68 VGND 0.00603f
C14475 XThC.XTBN.Y.t51 VGND 0.01024f
C14476 XThC.XTBN.Y.n127 VGND 0.01243f
C14477 XThC.XTBN.Y.t77 VGND 0.00603f
C14478 XThC.XTBN.Y.t58 VGND 0.01024f
C14479 XThC.XTBN.Y.n128 VGND 0.01348f
C14480 XThC.XTBN.Y.n129 VGND 0.0076f
C14481 XThC.XTBN.Y.n130 VGND 0.01252f
C14482 XThC.XTBN.Y.n131 VGND 0.00434f
C14483 XThC.XTBN.Y.n132 VGND 0.00603f
C14484 XThC.XTBN.Y.n133 VGND 0.01348f
C14485 XThC.XTBN.Y.t115 VGND 0.00603f
C14486 XThC.XTBN.Y.t99 VGND 0.01024f
C14487 XThC.XTBN.Y.n134 VGND 0.01227f
C14488 XThC.XTBN.Y.n135 VGND 0.00676f
C14489 XThC.XTBN.Y.n136 VGND 0.00747f
C14490 XThC.XTBN.Y.n137 VGND 0.07521f
C14491 XThC.XTBN.Y.t88 VGND 0.01024f
C14492 XThC.XTBN.Y.t60 VGND 0.00603f
C14493 XThC.XTBN.Y.n138 VGND 0.00619f
C14494 XThC.XTBN.Y.t37 VGND 0.01024f
C14495 XThC.XTBN.Y.t20 VGND 0.00603f
C14496 XThC.XTBN.Y.n139 VGND 0.01243f
C14497 XThC.XTBN.Y.t40 VGND 0.01024f
C14498 XThC.XTBN.Y.t22 VGND 0.00603f
C14499 XThC.XTBN.Y.n140 VGND 0.01348f
C14500 XThC.XTBN.Y.n141 VGND 0.0076f
C14501 XThC.XTBN.Y.n142 VGND 0.01252f
C14502 XThC.XTBN.Y.n143 VGND 0.00434f
C14503 XThC.XTBN.Y.n144 VGND 0.00603f
C14504 XThC.XTBN.Y.n145 VGND 0.01348f
C14505 XThC.XTBN.Y.t91 VGND 0.01024f
C14506 XThC.XTBN.Y.t66 VGND 0.00603f
C14507 XThC.XTBN.Y.n146 VGND 0.01227f
C14508 XThC.XTBN.Y.n147 VGND 0.00676f
C14509 XThC.XTBN.Y.n148 VGND 0.00747f
C14510 XThC.XTBN.Y.n149 VGND 0.07534f
C14511 XThC.XTBN.Y.t45 VGND 0.00603f
C14512 XThC.XTBN.Y.t7 VGND 0.01024f
C14513 XThC.XTBN.Y.n150 VGND 0.00619f
C14514 XThC.XTBN.Y.t5 VGND 0.00603f
C14515 XThC.XTBN.Y.t81 VGND 0.01024f
C14516 XThC.XTBN.Y.n151 VGND 0.01243f
C14517 XThC.XTBN.Y.t11 VGND 0.00603f
C14518 XThC.XTBN.Y.t86 VGND 0.01024f
C14519 XThC.XTBN.Y.n152 VGND 0.01348f
C14520 XThC.XTBN.Y.n153 VGND 0.0076f
C14521 XThC.XTBN.Y.n154 VGND 0.01252f
C14522 XThC.XTBN.Y.n155 VGND 0.00434f
C14523 XThC.XTBN.Y.n156 VGND 0.00603f
C14524 XThC.XTBN.Y.n157 VGND 0.01348f
C14525 XThC.XTBN.Y.t53 VGND 0.00603f
C14526 XThC.XTBN.Y.t13 VGND 0.01024f
C14527 XThC.XTBN.Y.n158 VGND 0.01227f
C14528 XThC.XTBN.Y.n159 VGND 0.00676f
C14529 XThC.XTBN.Y.n160 VGND 0.00747f
C14530 XThC.XTBN.Y.n161 VGND 0.07521f
C14531 XThC.XTBN.Y.t23 VGND 0.01024f
C14532 XThC.XTBN.Y.t117 VGND 0.00603f
C14533 XThC.XTBN.Y.n162 VGND 0.00619f
C14534 XThC.XTBN.Y.t95 VGND 0.01024f
C14535 XThC.XTBN.Y.t78 VGND 0.00603f
C14536 XThC.XTBN.Y.n163 VGND 0.01243f
C14537 XThC.XTBN.Y.t97 VGND 0.01024f
C14538 XThC.XTBN.Y.t80 VGND 0.00603f
C14539 XThC.XTBN.Y.n164 VGND 0.01348f
C14540 XThC.XTBN.Y.n165 VGND 0.0076f
C14541 XThC.XTBN.Y.n166 VGND 0.01252f
C14542 XThC.XTBN.Y.n167 VGND 0.00434f
C14543 XThC.XTBN.Y.n168 VGND 0.00603f
C14544 XThC.XTBN.Y.n169 VGND 0.01348f
C14545 XThC.XTBN.Y.t28 VGND 0.01024f
C14546 XThC.XTBN.Y.t4 VGND 0.00603f
C14547 XThC.XTBN.Y.n170 VGND 0.01227f
C14548 XThC.XTBN.Y.n171 VGND 0.00676f
C14549 XThC.XTBN.Y.n172 VGND 0.00747f
C14550 XThC.XTBN.Y.n173 VGND 0.08751f
C14551 XThC.XTBN.Y.n174 VGND 0.11019f
C14552 XThC.XTBN.Y.t105 VGND 0.00603f
C14553 XThC.XTBN.Y.t75 VGND 0.01024f
C14554 XThC.XTBN.Y.t69 VGND 0.00603f
C14555 XThC.XTBN.Y.t33 VGND 0.01024f
C14556 XThC.XTBN.Y.n175 VGND 0.01477f
C14557 XThC.XTBN.Y.t61 VGND 0.00603f
C14558 XThC.XTBN.Y.t27 VGND 0.01024f
C14559 XThC.XTBN.Y.n176 VGND 0.02293f
C14560 XThC.XTBN.Y.n177 VGND 0.00676f
C14561 XThC.XTBN.Y.n178 VGND 0.00561f
C14562 XThC.XTBN.Y.n179 VGND 0.00561f
C14563 XThC.XTBN.Y.n180 VGND 0.00676f
C14564 XThC.XTBN.Y.n181 VGND 0.01477f
C14565 XThC.XTBN.Y.t14 VGND 0.00603f
C14566 XThC.XTBN.Y.t9 VGND 0.01024f
C14567 XThC.XTBN.Y.n182 VGND 0.0138f
C14568 XThC.XTBN.Y.n183 VGND 0.00676f
C14569 XThC.XTBN.Y.n184 VGND 0.00372f
C14570 XThC.XTBN.Y.n185 VGND 0.00408f
C14571 XThC.XTBN.Y.n186 VGND 0.11129f
C14572 XThC.XTBN.Y.n187 VGND 0.02169f
C14573 XThC.XTBN.Y.t3 VGND 0.00428f
C14574 XThC.XTBN.Y.t2 VGND 0.00428f
C14575 XThC.XTBN.Y.n188 VGND 0.0094f
C14576 XThC.XTBN.Y.n189 VGND 0.00607f
C14577 XThC.XTBN.Y.n190 VGND 0.00526f
C14578 XThC.XTBN.Y.t0 VGND 0.00658f
C14579 XThC.XTBN.Y.t1 VGND 0.00658f
C14580 XThC.XTBN.Y.n191 VGND 0.01513f
C14581 XThC.XTBN.Y.n192 VGND 0.0307f
C14582 XThR.Tn[12].t0 VGND 0.02425f
C14583 XThR.Tn[12].t2 VGND 0.02425f
C14584 XThR.Tn[12].n0 VGND 0.0539f
C14585 XThR.Tn[12].t3 VGND 0.02425f
C14586 XThR.Tn[12].t1 VGND 0.02425f
C14587 XThR.Tn[12].n1 VGND 0.07362f
C14588 XThR.Tn[12].n2 VGND 0.24508f
C14589 XThR.Tn[12].t11 VGND 0.01576f
C14590 XThR.Tn[12].t9 VGND 0.01576f
C14591 XThR.Tn[12].n3 VGND 0.03931f
C14592 XThR.Tn[12].t10 VGND 0.01576f
C14593 XThR.Tn[12].t8 VGND 0.01576f
C14594 XThR.Tn[12].n4 VGND 0.03152f
C14595 XThR.Tn[12].n5 VGND 0.07268f
C14596 XThR.Tn[12].t36 VGND 0.01895f
C14597 XThR.Tn[12].t28 VGND 0.02075f
C14598 XThR.Tn[12].n6 VGND 0.05067f
C14599 XThR.Tn[12].n7 VGND 0.09734f
C14600 XThR.Tn[12].t53 VGND 0.01895f
C14601 XThR.Tn[12].t43 VGND 0.02075f
C14602 XThR.Tn[12].n8 VGND 0.05067f
C14603 XThR.Tn[12].t71 VGND 0.01889f
C14604 XThR.Tn[12].t21 VGND 0.02068f
C14605 XThR.Tn[12].n9 VGND 0.05272f
C14606 XThR.Tn[12].n10 VGND 0.03704f
C14607 XThR.Tn[12].n11 VGND 0.00677f
C14608 XThR.Tn[12].n12 VGND 0.11886f
C14609 XThR.Tn[12].t30 VGND 0.01895f
C14610 XThR.Tn[12].t20 VGND 0.02075f
C14611 XThR.Tn[12].n13 VGND 0.05067f
C14612 XThR.Tn[12].t49 VGND 0.01889f
C14613 XThR.Tn[12].t60 VGND 0.02068f
C14614 XThR.Tn[12].n14 VGND 0.05272f
C14615 XThR.Tn[12].n15 VGND 0.03704f
C14616 XThR.Tn[12].n16 VGND 0.00677f
C14617 XThR.Tn[12].n17 VGND 0.11886f
C14618 XThR.Tn[12].t45 VGND 0.01895f
C14619 XThR.Tn[12].t38 VGND 0.02075f
C14620 XThR.Tn[12].n18 VGND 0.05067f
C14621 XThR.Tn[12].t63 VGND 0.01889f
C14622 XThR.Tn[12].t15 VGND 0.02068f
C14623 XThR.Tn[12].n19 VGND 0.05272f
C14624 XThR.Tn[12].n20 VGND 0.03704f
C14625 XThR.Tn[12].n21 VGND 0.00677f
C14626 XThR.Tn[12].n22 VGND 0.11886f
C14627 XThR.Tn[12].t70 VGND 0.01895f
C14628 XThR.Tn[12].t66 VGND 0.02075f
C14629 XThR.Tn[12].n23 VGND 0.05067f
C14630 XThR.Tn[12].t33 VGND 0.01889f
C14631 XThR.Tn[12].t46 VGND 0.02068f
C14632 XThR.Tn[12].n24 VGND 0.05272f
C14633 XThR.Tn[12].n25 VGND 0.03704f
C14634 XThR.Tn[12].n26 VGND 0.00677f
C14635 XThR.Tn[12].n27 VGND 0.11886f
C14636 XThR.Tn[12].t48 VGND 0.01895f
C14637 XThR.Tn[12].t39 VGND 0.02075f
C14638 XThR.Tn[12].n28 VGND 0.05067f
C14639 XThR.Tn[12].t64 VGND 0.01889f
C14640 XThR.Tn[12].t17 VGND 0.02068f
C14641 XThR.Tn[12].n29 VGND 0.05272f
C14642 XThR.Tn[12].n30 VGND 0.03704f
C14643 XThR.Tn[12].n31 VGND 0.00677f
C14644 XThR.Tn[12].n32 VGND 0.11886f
C14645 XThR.Tn[12].t23 VGND 0.01895f
C14646 XThR.Tn[12].t56 VGND 0.02075f
C14647 XThR.Tn[12].n33 VGND 0.05067f
C14648 XThR.Tn[12].t41 VGND 0.01889f
C14649 XThR.Tn[12].t37 VGND 0.02068f
C14650 XThR.Tn[12].n34 VGND 0.05272f
C14651 XThR.Tn[12].n35 VGND 0.03704f
C14652 XThR.Tn[12].n36 VGND 0.00677f
C14653 XThR.Tn[12].n37 VGND 0.11886f
C14654 XThR.Tn[12].t54 VGND 0.01895f
C14655 XThR.Tn[12].t51 VGND 0.02075f
C14656 XThR.Tn[12].n38 VGND 0.05067f
C14657 XThR.Tn[12].t72 VGND 0.01889f
C14658 XThR.Tn[12].t29 VGND 0.02068f
C14659 XThR.Tn[12].n39 VGND 0.05272f
C14660 XThR.Tn[12].n40 VGND 0.03704f
C14661 XThR.Tn[12].n41 VGND 0.00677f
C14662 XThR.Tn[12].n42 VGND 0.11886f
C14663 XThR.Tn[12].t59 VGND 0.01895f
C14664 XThR.Tn[12].t65 VGND 0.02075f
C14665 XThR.Tn[12].n43 VGND 0.05067f
C14666 XThR.Tn[12].t14 VGND 0.01889f
C14667 XThR.Tn[12].t44 VGND 0.02068f
C14668 XThR.Tn[12].n44 VGND 0.05272f
C14669 XThR.Tn[12].n45 VGND 0.03704f
C14670 XThR.Tn[12].n46 VGND 0.00677f
C14671 XThR.Tn[12].n47 VGND 0.11886f
C14672 XThR.Tn[12].t12 VGND 0.01895f
C14673 XThR.Tn[12].t22 VGND 0.02075f
C14674 XThR.Tn[12].n48 VGND 0.05067f
C14675 XThR.Tn[12].t35 VGND 0.01889f
C14676 XThR.Tn[12].t61 VGND 0.02068f
C14677 XThR.Tn[12].n49 VGND 0.05272f
C14678 XThR.Tn[12].n50 VGND 0.03704f
C14679 XThR.Tn[12].n51 VGND 0.00677f
C14680 XThR.Tn[12].n52 VGND 0.11886f
C14681 XThR.Tn[12].t68 VGND 0.01895f
C14682 XThR.Tn[12].t40 VGND 0.02075f
C14683 XThR.Tn[12].n53 VGND 0.05067f
C14684 XThR.Tn[12].t26 VGND 0.01889f
C14685 XThR.Tn[12].t19 VGND 0.02068f
C14686 XThR.Tn[12].n54 VGND 0.05272f
C14687 XThR.Tn[12].n55 VGND 0.03704f
C14688 XThR.Tn[12].n56 VGND 0.00677f
C14689 XThR.Tn[12].n57 VGND 0.11886f
C14690 XThR.Tn[12].t25 VGND 0.01895f
C14691 XThR.Tn[12].t16 VGND 0.02075f
C14692 XThR.Tn[12].n58 VGND 0.05067f
C14693 XThR.Tn[12].t42 VGND 0.01889f
C14694 XThR.Tn[12].t55 VGND 0.02068f
C14695 XThR.Tn[12].n59 VGND 0.05272f
C14696 XThR.Tn[12].n60 VGND 0.03704f
C14697 XThR.Tn[12].n61 VGND 0.00677f
C14698 XThR.Tn[12].n62 VGND 0.11886f
C14699 XThR.Tn[12].t57 VGND 0.01895f
C14700 XThR.Tn[12].t52 VGND 0.02075f
C14701 XThR.Tn[12].n63 VGND 0.05067f
C14702 XThR.Tn[12].t13 VGND 0.01889f
C14703 XThR.Tn[12].t31 VGND 0.02068f
C14704 XThR.Tn[12].n64 VGND 0.05272f
C14705 XThR.Tn[12].n65 VGND 0.03704f
C14706 XThR.Tn[12].n66 VGND 0.00677f
C14707 XThR.Tn[12].n67 VGND 0.11886f
C14708 XThR.Tn[12].t73 VGND 0.01895f
C14709 XThR.Tn[12].t67 VGND 0.02075f
C14710 XThR.Tn[12].n68 VGND 0.05067f
C14711 XThR.Tn[12].t34 VGND 0.01889f
C14712 XThR.Tn[12].t47 VGND 0.02068f
C14713 XThR.Tn[12].n69 VGND 0.05272f
C14714 XThR.Tn[12].n70 VGND 0.03704f
C14715 XThR.Tn[12].n71 VGND 0.00677f
C14716 XThR.Tn[12].n72 VGND 0.11886f
C14717 XThR.Tn[12].t32 VGND 0.01895f
C14718 XThR.Tn[12].t24 VGND 0.02075f
C14719 XThR.Tn[12].n73 VGND 0.05067f
C14720 XThR.Tn[12].t50 VGND 0.01889f
C14721 XThR.Tn[12].t62 VGND 0.02068f
C14722 XThR.Tn[12].n74 VGND 0.05272f
C14723 XThR.Tn[12].n75 VGND 0.03704f
C14724 XThR.Tn[12].n76 VGND 0.00677f
C14725 XThR.Tn[12].n77 VGND 0.11886f
C14726 XThR.Tn[12].t69 VGND 0.01895f
C14727 XThR.Tn[12].t18 VGND 0.02075f
C14728 XThR.Tn[12].n78 VGND 0.05067f
C14729 XThR.Tn[12].t27 VGND 0.01889f
C14730 XThR.Tn[12].t58 VGND 0.02068f
C14731 XThR.Tn[12].n79 VGND 0.05272f
C14732 XThR.Tn[12].n80 VGND 0.03704f
C14733 XThR.Tn[12].n81 VGND 0.00677f
C14734 XThR.Tn[12].n82 VGND 0.11886f
C14735 XThR.Tn[12].n83 VGND 0.10802f
C14736 XThR.Tn[12].n84 VGND 0.36839f
C14737 XThR.Tn[12].t6 VGND 0.02425f
C14738 XThR.Tn[12].t4 VGND 0.02425f
C14739 XThR.Tn[12].n85 VGND 0.05239f
C14740 XThR.Tn[12].t7 VGND 0.02425f
C14741 XThR.Tn[12].t5 VGND 0.02425f
C14742 XThR.Tn[12].n86 VGND 0.07973f
C14743 XThR.Tn[12].n87 VGND 0.2214f
C14744 XThR.Tn[12].n88 VGND 0.01091f
C14745 Vbias.n0 VGND 0.99957f
C14746 Vbias.t176 VGND 0.32014f
C14747 Vbias.n1 VGND 0.31618f
C14748 Vbias.t105 VGND 0.32014f
C14749 Vbias.n2 VGND 0.31618f
C14750 Vbias.n3 VGND 0.08903f
C14751 Vbias.n4 VGND 0.33651f
C14752 Vbias.t141 VGND 0.32014f
C14753 Vbias.n5 VGND 0.31618f
C14754 Vbias.t233 VGND 0.32014f
C14755 Vbias.n6 VGND 0.31618f
C14756 Vbias.n7 VGND 0.33651f
C14757 Vbias.t205 VGND 0.32014f
C14758 Vbias.n8 VGND 0.31618f
C14759 Vbias.n9 VGND 0.08903f
C14760 Vbias.t19 VGND 0.32014f
C14761 Vbias.n10 VGND 0.31618f
C14762 Vbias.t7 VGND 0.32014f
C14763 Vbias.n11 VGND 0.31618f
C14764 Vbias.n12 VGND 0.33651f
C14765 Vbias.t188 VGND 0.32014f
C14766 Vbias.n13 VGND 0.31618f
C14767 Vbias.n14 VGND 0.18804f
C14768 Vbias.n15 VGND 0.18804f
C14769 Vbias.t168 VGND 0.32014f
C14770 Vbias.n16 VGND 0.31618f
C14771 Vbias.n17 VGND 0.33651f
C14772 Vbias.t243 VGND 0.32014f
C14773 Vbias.n18 VGND 0.31618f
C14774 Vbias.t90 VGND 0.32014f
C14775 Vbias.n19 VGND 0.31618f
C14776 Vbias.n20 VGND 0.33651f
C14777 Vbias.t20 VGND 0.32014f
C14778 Vbias.n21 VGND 0.31618f
C14779 Vbias.t253 VGND 0.32014f
C14780 Vbias.n22 VGND 0.31618f
C14781 Vbias.n23 VGND 0.33651f
C14782 Vbias.t70 VGND 0.32014f
C14783 Vbias.n24 VGND 0.31618f
C14784 Vbias.t241 VGND 0.32014f
C14785 Vbias.n25 VGND 0.31618f
C14786 Vbias.n26 VGND 0.33651f
C14787 Vbias.t166 VGND 0.32014f
C14788 Vbias.n27 VGND 0.31618f
C14789 Vbias.t91 VGND 0.32014f
C14790 Vbias.n28 VGND 0.31618f
C14791 Vbias.n29 VGND 0.33651f
C14792 Vbias.t164 VGND 0.32014f
C14793 Vbias.n30 VGND 0.31618f
C14794 Vbias.t142 VGND 0.32014f
C14795 Vbias.n31 VGND 0.31618f
C14796 Vbias.n32 VGND 0.33651f
C14797 Vbias.t71 VGND 0.32014f
C14798 Vbias.n33 VGND 0.31618f
C14799 Vbias.t242 VGND 0.32014f
C14800 Vbias.n34 VGND 0.31618f
C14801 Vbias.n35 VGND 0.33651f
C14802 Vbias.t55 VGND 0.32014f
C14803 Vbias.n36 VGND 0.31618f
C14804 Vbias.t222 VGND 0.32014f
C14805 Vbias.n37 VGND 0.31618f
C14806 Vbias.n38 VGND 0.33651f
C14807 Vbias.t151 VGND 0.32014f
C14808 Vbias.n39 VGND 0.31618f
C14809 Vbias.t64 VGND 0.32014f
C14810 Vbias.n40 VGND 0.31618f
C14811 Vbias.n41 VGND 0.33651f
C14812 Vbias.t136 VGND 0.32014f
C14813 Vbias.n42 VGND 0.31618f
C14814 Vbias.t51 VGND 0.32014f
C14815 Vbias.n43 VGND 0.31618f
C14816 Vbias.n44 VGND 0.33651f
C14817 Vbias.t238 VGND 0.32014f
C14818 Vbias.n45 VGND 0.31618f
C14819 Vbias.t224 VGND 0.32014f
C14820 Vbias.n46 VGND 0.31618f
C14821 Vbias.n47 VGND 0.33651f
C14822 Vbias.t36 VGND 0.32014f
C14823 Vbias.n48 VGND 0.31618f
C14824 Vbias.t196 VGND 0.32014f
C14825 Vbias.n49 VGND 0.31618f
C14826 Vbias.n50 VGND 0.33651f
C14827 Vbias.t125 VGND 0.32014f
C14828 Vbias.n51 VGND 0.31618f
C14829 Vbias.t52 VGND 0.32014f
C14830 Vbias.n52 VGND 0.31618f
C14831 Vbias.t124 VGND 0.32014f
C14832 Vbias.n53 VGND 0.31618f
C14833 Vbias.n54 VGND 0.04247f
C14834 Vbias.t82 VGND 0.32014f
C14835 Vbias.n55 VGND 0.31618f
C14836 Vbias.t220 VGND 0.32014f
C14837 Vbias.n56 VGND 0.31618f
C14838 Vbias.n57 VGND 0.08903f
C14839 Vbias.n58 VGND 0.18804f
C14840 Vbias.t200 VGND 0.32014f
C14841 Vbias.n59 VGND 0.31618f
C14842 Vbias.n60 VGND 0.08903f
C14843 Vbias.n61 VGND 0.18804f
C14844 Vbias.t47 VGND 0.32014f
C14845 Vbias.n62 VGND 0.31618f
C14846 Vbias.n63 VGND 0.08903f
C14847 Vbias.n64 VGND 0.18804f
C14848 Vbias.t27 VGND 0.32014f
C14849 Vbias.n65 VGND 0.31618f
C14850 Vbias.n66 VGND 0.08903f
C14851 Vbias.n67 VGND 0.18804f
C14852 Vbias.t194 VGND 0.32014f
C14853 Vbias.n68 VGND 0.31618f
C14854 Vbias.n69 VGND 0.08903f
C14855 Vbias.n70 VGND 0.18804f
C14856 Vbias.t120 VGND 0.32014f
C14857 Vbias.n71 VGND 0.31618f
C14858 Vbias.n72 VGND 0.08903f
C14859 Vbias.n73 VGND 0.18804f
C14860 Vbias.t97 VGND 0.32014f
C14861 Vbias.n74 VGND 0.31618f
C14862 Vbias.n75 VGND 0.08903f
C14863 Vbias.n76 VGND 0.18804f
C14864 Vbias.t13 VGND 0.32014f
C14865 Vbias.n77 VGND 0.31618f
C14866 Vbias.n78 VGND 0.08903f
C14867 Vbias.n79 VGND 0.18804f
C14868 Vbias.t178 VGND 0.32014f
C14869 Vbias.n80 VGND 0.31618f
C14870 Vbias.n81 VGND 0.08903f
C14871 Vbias.n82 VGND 0.18804f
C14872 Vbias.t94 VGND 0.32014f
C14873 Vbias.n83 VGND 0.31618f
C14874 Vbias.n84 VGND 0.08903f
C14875 Vbias.n85 VGND 0.18804f
C14876 Vbias.t9 VGND 0.32014f
C14877 Vbias.n86 VGND 0.31618f
C14878 Vbias.n87 VGND 0.08903f
C14879 Vbias.n88 VGND 0.18804f
C14880 Vbias.t256 VGND 0.32014f
C14881 Vbias.n89 VGND 0.31618f
C14882 Vbias.n90 VGND 0.08903f
C14883 Vbias.n91 VGND 0.18804f
C14884 Vbias.t155 VGND 0.32014f
C14885 Vbias.n92 VGND 0.31618f
C14886 Vbias.n93 VGND 0.08903f
C14887 Vbias.n94 VGND 0.18804f
C14888 Vbias.n95 VGND 0.08642f
C14889 Vbias.n96 VGND 0.33651f
C14890 Vbias.t11 VGND 0.32014f
C14891 Vbias.n97 VGND 0.31618f
C14892 Vbias.t83 VGND 0.32014f
C14893 Vbias.n98 VGND 0.31618f
C14894 Vbias.n99 VGND 0.33651f
C14895 Vbias.t12 VGND 0.32014f
C14896 Vbias.n100 VGND 0.31618f
C14897 Vbias.t108 VGND 0.32014f
C14898 Vbias.n101 VGND 0.31618f
C14899 Vbias.n102 VGND 0.33651f
C14900 Vbias.t180 VGND 0.32014f
C14901 Vbias.n103 VGND 0.31618f
C14902 Vbias.t192 VGND 0.32014f
C14903 Vbias.n104 VGND 0.31618f
C14904 Vbias.n105 VGND 0.33651f
C14905 Vbias.t118 VGND 0.32014f
C14906 Vbias.n106 VGND 0.31618f
C14907 Vbias.t208 VGND 0.32014f
C14908 Vbias.n107 VGND 0.31618f
C14909 Vbias.n108 VGND 0.33651f
C14910 Vbias.t24 VGND 0.32014f
C14911 Vbias.n109 VGND 0.31618f
C14912 Vbias.t107 VGND 0.32014f
C14913 Vbias.n110 VGND 0.31618f
C14914 Vbias.n111 VGND 0.33651f
C14915 Vbias.t35 VGND 0.32014f
C14916 Vbias.n112 VGND 0.31618f
C14917 Vbias.t122 VGND 0.32014f
C14918 Vbias.n113 VGND 0.31618f
C14919 Vbias.n114 VGND 0.33651f
C14920 Vbias.t195 VGND 0.32014f
C14921 Vbias.n115 VGND 0.31618f
C14922 Vbias.t28 VGND 0.32014f
C14923 Vbias.n116 VGND 0.31618f
C14924 Vbias.n117 VGND 0.33651f
C14925 Vbias.t214 VGND 0.32014f
C14926 Vbias.n118 VGND 0.31618f
C14927 Vbias.t235 VGND 0.32014f
C14928 Vbias.n119 VGND 0.31618f
C14929 Vbias.n120 VGND 0.33651f
C14930 Vbias.t48 VGND 0.32014f
C14931 Vbias.n121 VGND 0.31618f
C14932 Vbias.t121 VGND 0.32014f
C14933 Vbias.n122 VGND 0.31618f
C14934 Vbias.n123 VGND 0.33651f
C14935 Vbias.t49 VGND 0.32014f
C14936 Vbias.n124 VGND 0.31618f
C14937 Vbias.t139 VGND 0.32014f
C14938 Vbias.n125 VGND 0.31618f
C14939 Vbias.n126 VGND 0.33651f
C14940 Vbias.t212 VGND 0.32014f
C14941 Vbias.n127 VGND 0.31618f
C14942 Vbias.t234 VGND 0.32014f
C14943 Vbias.n128 VGND 0.31618f
C14944 Vbias.n129 VGND 0.33651f
C14945 Vbias.t161 VGND 0.32014f
C14946 Vbias.n130 VGND 0.31618f
C14947 Vbias.t57 VGND 0.32014f
C14948 Vbias.n131 VGND 0.31618f
C14949 Vbias.n132 VGND 0.33651f
C14950 Vbias.t128 VGND 0.32014f
C14951 Vbias.n133 VGND 0.31618f
C14952 Vbias.t148 VGND 0.32014f
C14953 Vbias.n134 VGND 0.31618f
C14954 Vbias.n135 VGND 0.33651f
C14955 Vbias.t76 VGND 0.32014f
C14956 Vbias.n136 VGND 0.31618f
C14957 Vbias.t87 VGND 0.32014f
C14958 Vbias.n137 VGND 0.31618f
C14959 Vbias.n138 VGND 0.33651f
C14960 Vbias.t15 VGND 0.32014f
C14961 Vbias.n139 VGND 0.31618f
C14962 Vbias.t116 VGND 0.32014f
C14963 Vbias.n140 VGND 0.31618f
C14964 Vbias.t44 VGND 0.32014f
C14965 Vbias.n141 VGND 0.31618f
C14966 Vbias.n142 VGND 0.08642f
C14967 Vbias.n143 VGND 0.33651f
C14968 Vbias.t77 VGND 0.32014f
C14969 Vbias.n144 VGND 0.31618f
C14970 Vbias.t149 VGND 0.32014f
C14971 Vbias.n145 VGND 0.31618f
C14972 Vbias.n146 VGND 0.33651f
C14973 Vbias.t117 VGND 0.32014f
C14974 Vbias.n147 VGND 0.31618f
C14975 Vbias.t217 VGND 0.32014f
C14976 Vbias.n148 VGND 0.31618f
C14977 Vbias.n149 VGND 0.33651f
C14978 Vbias.t252 VGND 0.32014f
C14979 Vbias.n150 VGND 0.31618f
C14980 Vbias.t259 VGND 0.32014f
C14981 Vbias.n151 VGND 0.31618f
C14982 Vbias.n152 VGND 0.33651f
C14983 Vbias.t230 VGND 0.32014f
C14984 Vbias.n153 VGND 0.31618f
C14985 Vbias.t58 VGND 0.32014f
C14986 Vbias.n154 VGND 0.31618f
C14987 Vbias.n155 VGND 0.33651f
C14988 Vbias.t88 VGND 0.32014f
C14989 Vbias.n156 VGND 0.31618f
C14990 Vbias.t174 VGND 0.32014f
C14991 Vbias.n157 VGND 0.31618f
C14992 Vbias.n158 VGND 0.33651f
C14993 Vbias.t145 VGND 0.32014f
C14994 Vbias.n159 VGND 0.31618f
C14995 Vbias.t232 VGND 0.32014f
C14996 Vbias.n160 VGND 0.31618f
C14997 Vbias.n161 VGND 0.33651f
C14998 Vbias.t6 VGND 0.32014f
C14999 Vbias.n162 VGND 0.31618f
C15000 Vbias.t93 VGND 0.32014f
C15001 Vbias.n163 VGND 0.31618f
C15002 Vbias.n164 VGND 0.33651f
C15003 Vbias.t62 VGND 0.32014f
C15004 Vbias.n165 VGND 0.31618f
C15005 Vbias.t86 VGND 0.32014f
C15006 Vbias.n166 VGND 0.31618f
C15007 Vbias.n167 VGND 0.33651f
C15008 Vbias.t113 VGND 0.32014f
C15009 Vbias.n168 VGND 0.31618f
C15010 Vbias.t186 VGND 0.32014f
C15011 Vbias.n169 VGND 0.31618f
C15012 Vbias.n170 VGND 0.33651f
C15013 Vbias.t159 VGND 0.32014f
C15014 Vbias.n171 VGND 0.31618f
C15015 Vbias.t246 VGND 0.32014f
C15016 Vbias.n172 VGND 0.31618f
C15017 Vbias.n173 VGND 0.33651f
C15018 Vbias.t22 VGND 0.32014f
C15019 Vbias.n174 VGND 0.31618f
C15020 Vbias.t39 VGND 0.32014f
C15021 Vbias.n175 VGND 0.31618f
C15022 Vbias.n176 VGND 0.33651f
C15023 Vbias.t16 VGND 0.32014f
C15024 Vbias.n177 VGND 0.31618f
C15025 Vbias.t163 VGND 0.32014f
C15026 Vbias.n178 VGND 0.31618f
C15027 Vbias.n179 VGND 0.33651f
C15028 Vbias.t191 VGND 0.32014f
C15029 Vbias.n180 VGND 0.31618f
C15030 Vbias.t215 VGND 0.32014f
C15031 Vbias.n181 VGND 0.31618f
C15032 Vbias.n182 VGND 0.33651f
C15033 Vbias.t182 VGND 0.32014f
C15034 Vbias.n183 VGND 0.31618f
C15035 Vbias.t100 VGND 0.32014f
C15036 Vbias.n184 VGND 0.31618f
C15037 Vbias.n185 VGND 0.33651f
C15038 Vbias.t132 VGND 0.32014f
C15039 Vbias.n186 VGND 0.31618f
C15040 Vbias.n187 VGND 0.08903f
C15041 Vbias.n188 VGND 0.33651f
C15042 Vbias.t59 VGND 0.32014f
C15043 Vbias.n189 VGND 0.31618f
C15044 Vbias.t260 VGND 0.32014f
C15045 Vbias.n190 VGND 0.31618f
C15046 Vbias.n191 VGND 0.08642f
C15047 Vbias.t78 VGND 0.32014f
C15048 Vbias.n192 VGND 0.31618f
C15049 Vbias.n193 VGND 0.08903f
C15050 Vbias.n194 VGND 0.18804f
C15051 Vbias.t175 VGND 0.32014f
C15052 Vbias.n195 VGND 0.31618f
C15053 Vbias.n196 VGND 0.08903f
C15054 Vbias.n197 VGND 0.18804f
C15055 Vbias.t183 VGND 0.32014f
C15056 Vbias.n198 VGND 0.31618f
C15057 Vbias.n199 VGND 0.08903f
C15058 Vbias.n200 VGND 0.18804f
C15059 Vbias.t18 VGND 0.32014f
C15060 Vbias.n201 VGND 0.31618f
C15061 Vbias.n202 VGND 0.08903f
C15062 Vbias.n203 VGND 0.18804f
C15063 Vbias.t102 VGND 0.32014f
C15064 Vbias.n204 VGND 0.31618f
C15065 Vbias.n205 VGND 0.08903f
C15066 Vbias.n206 VGND 0.18804f
C15067 Vbias.t187 VGND 0.32014f
C15068 Vbias.n207 VGND 0.31618f
C15069 Vbias.n208 VGND 0.08903f
C15070 Vbias.n209 VGND 0.18804f
C15071 Vbias.t23 VGND 0.32014f
C15072 Vbias.n210 VGND 0.31618f
C15073 Vbias.n211 VGND 0.08903f
C15074 Vbias.n212 VGND 0.18804f
C15075 Vbias.t40 VGND 0.32014f
C15076 Vbias.n213 VGND 0.31618f
C15077 Vbias.n214 VGND 0.08903f
C15078 Vbias.n215 VGND 0.18804f
C15079 Vbias.t114 VGND 0.32014f
C15080 Vbias.n216 VGND 0.31618f
C15081 Vbias.n217 VGND 0.08903f
C15082 Vbias.n218 VGND 0.18804f
C15083 Vbias.t206 VGND 0.32014f
C15084 Vbias.n219 VGND 0.31618f
C15085 Vbias.n220 VGND 0.08903f
C15086 Vbias.n221 VGND 0.18804f
C15087 Vbias.t228 VGND 0.32014f
C15088 Vbias.n222 VGND 0.31618f
C15089 Vbias.n223 VGND 0.08903f
C15090 Vbias.n224 VGND 0.18804f
C15091 Vbias.t119 VGND 0.32014f
C15092 Vbias.n225 VGND 0.31618f
C15093 Vbias.n226 VGND 0.08903f
C15094 Vbias.n227 VGND 0.18804f
C15095 Vbias.t144 VGND 0.32014f
C15096 Vbias.n228 VGND 0.31618f
C15097 Vbias.n229 VGND 0.08903f
C15098 Vbias.n230 VGND 0.18804f
C15099 Vbias.t156 VGND 0.32014f
C15100 Vbias.n231 VGND 0.31618f
C15101 Vbias.n232 VGND 0.33651f
C15102 Vbias.t227 VGND 0.32014f
C15103 Vbias.n233 VGND 0.31618f
C15104 Vbias.n234 VGND 0.99957f
C15105 Vbias.t75 VGND 0.32014f
C15106 Vbias.n235 VGND 0.31618f
C15107 Vbias.n236 VGND 0.33651f
C15108 Vbias.t185 VGND 0.32014f
C15109 Vbias.n237 VGND 0.31618f
C15110 Vbias.t167 VGND 0.32014f
C15111 Vbias.n238 VGND 0.31618f
C15112 Vbias.n239 VGND 0.33651f
C15113 Vbias.t46 VGND 0.32014f
C15114 Vbias.n240 VGND 0.31618f
C15115 Vbias.t157 VGND 0.32014f
C15116 Vbias.n241 VGND 0.31618f
C15117 Vbias.n242 VGND 0.33651f
C15118 Vbias.t17 VGND 0.32014f
C15119 Vbias.n243 VGND 0.31618f
C15120 Vbias.t251 VGND 0.32014f
C15121 Vbias.n244 VGND 0.31618f
C15122 Vbias.n245 VGND 0.33651f
C15123 Vbias.t131 VGND 0.32014f
C15124 Vbias.n246 VGND 0.31618f
C15125 Vbias.t41 VGND 0.32014f
C15126 Vbias.n247 VGND 0.31618f
C15127 Vbias.n248 VGND 0.33651f
C15128 Vbias.t162 VGND 0.32014f
C15129 Vbias.n249 VGND 0.31618f
C15130 Vbias.t89 VGND 0.32014f
C15131 Vbias.n250 VGND 0.31618f
C15132 Vbias.n251 VGND 0.33651f
C15133 Vbias.t229 VGND 0.32014f
C15134 Vbias.n252 VGND 0.31618f
C15135 Vbias.t207 VGND 0.32014f
C15136 Vbias.n253 VGND 0.31618f
C15137 Vbias.n254 VGND 0.33651f
C15138 Vbias.t69 VGND 0.32014f
C15139 Vbias.n255 VGND 0.31618f
C15140 Vbias.t239 VGND 0.32014f
C15141 Vbias.n256 VGND 0.31618f
C15142 Vbias.n257 VGND 0.33651f
C15143 Vbias.t115 VGND 0.32014f
C15144 Vbias.n258 VGND 0.31618f
C15145 Vbias.t31 VGND 0.32014f
C15146 Vbias.n259 VGND 0.31618f
C15147 Vbias.n260 VGND 0.33651f
C15148 Vbias.t150 VGND 0.32014f
C15149 Vbias.n261 VGND 0.31618f
C15150 Vbias.t61 VGND 0.32014f
C15151 Vbias.n262 VGND 0.31618f
C15152 Vbias.n263 VGND 0.33651f
C15153 Vbias.t203 VGND 0.32014f
C15154 Vbias.n264 VGND 0.31618f
C15155 Vbias.t112 VGND 0.32014f
C15156 Vbias.n265 VGND 0.31618f
C15157 Vbias.n266 VGND 0.33651f
C15158 Vbias.t236 VGND 0.32014f
C15159 Vbias.n267 VGND 0.31618f
C15160 Vbias.t221 VGND 0.32014f
C15161 Vbias.n268 VGND 0.31618f
C15162 Vbias.n269 VGND 0.33651f
C15163 Vbias.t103 VGND 0.32014f
C15164 Vbias.n270 VGND 0.31618f
C15165 Vbias.t261 VGND 0.32014f
C15166 Vbias.n271 VGND 0.31618f
C15167 Vbias.n272 VGND 0.33651f
C15168 Vbias.t123 VGND 0.32014f
C15169 Vbias.n273 VGND 0.31618f
C15170 Vbias.t50 VGND 0.32014f
C15171 Vbias.n274 VGND 0.31618f
C15172 Vbias.t184 VGND 0.32014f
C15173 Vbias.n275 VGND 0.31618f
C15174 Vbias.n276 VGND 0.08642f
C15175 Vbias.n277 VGND 0.33651f
C15176 Vbias.n278 VGND 0.33651f
C15177 Vbias.t181 VGND 0.32014f
C15178 Vbias.n279 VGND 0.31618f
C15179 Vbias.t80 VGND 0.32014f
C15180 Vbias.n280 VGND 0.31618f
C15181 Vbias.n281 VGND 0.33651f
C15182 Vbias.t202 VGND 0.32014f
C15183 Vbias.n282 VGND 0.31618f
C15184 Vbias.t104 VGND 0.32014f
C15185 Vbias.n283 VGND 0.31618f
C15186 Vbias.t244 VGND 0.32014f
C15187 Vbias.n284 VGND 0.31618f
C15188 Vbias.n285 VGND 0.08903f
C15189 Vbias.n286 VGND 0.33651f
C15190 Vbias.t81 VGND 0.32014f
C15191 Vbias.n287 VGND 0.31618f
C15192 Vbias.t165 VGND 0.32014f
C15193 Vbias.n288 VGND 0.31618f
C15194 Vbias.n289 VGND 0.34709f
C15195 Vbias.t92 VGND 0.32014f
C15196 Vbias.n290 VGND 0.31618f
C15197 Vbias.t72 VGND 0.32014f
C15198 Vbias.n291 VGND 0.31618f
C15199 Vbias.n292 VGND 0.34709f
C15200 Vbias.t143 VGND 0.32014f
C15201 Vbias.n293 VGND 0.31618f
C15202 Vbias.t247 VGND 0.32014f
C15203 Vbias.n294 VGND 0.31618f
C15204 Vbias.n295 VGND 0.34709f
C15205 Vbias.t172 VGND 0.32014f
C15206 Vbias.n296 VGND 0.31618f
C15207 Vbias.t152 VGND 0.32014f
C15208 Vbias.n297 VGND 0.31618f
C15209 Vbias.n298 VGND 0.34709f
C15210 Vbias.t223 VGND 0.32014f
C15211 Vbias.n299 VGND 0.31618f
C15212 Vbias.t138 VGND 0.32014f
C15213 Vbias.n300 VGND 0.31618f
C15214 Vbias.n301 VGND 0.34709f
C15215 Vbias.t66 VGND 0.32014f
C15216 Vbias.n302 VGND 0.31618f
C15217 Vbias.t248 VGND 0.32014f
C15218 Vbias.n303 VGND 0.31618f
C15219 Vbias.n304 VGND 0.34709f
C15220 Vbias.t65 VGND 0.32014f
C15221 Vbias.n305 VGND 0.31618f
C15222 Vbias.t37 VGND 0.32014f
C15223 Vbias.n306 VGND 0.31618f
C15224 Vbias.n307 VGND 0.34709f
C15225 Vbias.t225 VGND 0.32014f
C15226 Vbias.n308 VGND 0.31618f
C15227 Vbias.t140 VGND 0.32014f
C15228 Vbias.n309 VGND 0.31618f
C15229 Vbias.n310 VGND 0.34709f
C15230 Vbias.t213 VGND 0.32014f
C15231 Vbias.n311 VGND 0.31618f
C15232 Vbias.t126 VGND 0.32014f
C15233 Vbias.n312 VGND 0.31618f
C15234 Vbias.n313 VGND 0.34709f
C15235 Vbias.t53 VGND 0.32014f
C15236 Vbias.n314 VGND 0.31618f
C15237 Vbias.t219 VGND 0.32014f
C15238 Vbias.n315 VGND 0.31618f
C15239 Vbias.n316 VGND 0.34709f
C15240 Vbias.t33 VGND 0.32014f
C15241 Vbias.n317 VGND 0.31618f
C15242 Vbias.t209 VGND 0.32014f
C15243 Vbias.n318 VGND 0.31618f
C15244 Vbias.n319 VGND 0.34709f
C15245 Vbias.t134 VGND 0.32014f
C15246 Vbias.n320 VGND 0.31618f
C15247 Vbias.t127 VGND 0.32014f
C15248 Vbias.n321 VGND 0.31618f
C15249 Vbias.n322 VGND 0.34709f
C15250 Vbias.t198 VGND 0.32014f
C15251 Vbias.n323 VGND 0.31618f
C15252 Vbias.t25 VGND 0.32014f
C15253 Vbias.n324 VGND 0.31618f
C15254 Vbias.n325 VGND 0.08642f
C15255 Vbias.t95 VGND 0.32014f
C15256 Vbias.n326 VGND 0.31618f
C15257 Vbias.n327 VGND 0.34709f
C15258 Vbias.t26 VGND 0.32014f
C15259 Vbias.n328 VGND 0.31618f
C15260 Vbias.t210 VGND 0.32014f
C15261 Vbias.n329 VGND 0.31618f
C15262 Vbias.t135 VGND 0.32014f
C15263 Vbias.n330 VGND 0.31618f
C15264 Vbias.n331 VGND 0.08642f
C15265 Vbias.t255 VGND 0.32014f
C15266 Vbias.n332 VGND 0.31618f
C15267 Vbias.t146 VGND 0.32014f
C15268 Vbias.n333 VGND 0.31618f
C15269 Vbias.t30 VGND 0.32014f
C15270 Vbias.n334 VGND 0.31618f
C15271 Vbias.n335 VGND 0.08903f
C15272 Vbias.t99 VGND 0.32014f
C15273 Vbias.n336 VGND 0.31618f
C15274 Vbias.n337 VGND 0.9716f
C15275 Vbias.t211 VGND 0.32014f
C15276 Vbias.n338 VGND 0.31618f
C15277 Vbias.n339 VGND 0.08903f
C15278 Vbias.n340 VGND 0.18804f
C15279 Vbias.t54 VGND 0.32014f
C15280 Vbias.n341 VGND 0.31618f
C15281 Vbias.n342 VGND 0.08903f
C15282 Vbias.n343 VGND 0.18804f
C15283 Vbias.t63 VGND 0.32014f
C15284 Vbias.n344 VGND 0.31618f
C15285 Vbias.n345 VGND 0.08903f
C15286 Vbias.n346 VGND 0.18804f
C15287 Vbias.t147 VGND 0.32014f
C15288 Vbias.n347 VGND 0.31618f
C15289 Vbias.n348 VGND 0.08903f
C15290 Vbias.n349 VGND 0.18804f
C15291 Vbias.t240 VGND 0.32014f
C15292 Vbias.n350 VGND 0.31618f
C15293 Vbias.n351 VGND 0.08903f
C15294 Vbias.n352 VGND 0.18804f
C15295 Vbias.t67 VGND 0.32014f
C15296 Vbias.n353 VGND 0.31618f
C15297 Vbias.n354 VGND 0.08903f
C15298 Vbias.n355 VGND 0.18804f
C15299 Vbias.t153 VGND 0.32014f
C15300 Vbias.n356 VGND 0.31618f
C15301 Vbias.n357 VGND 0.08903f
C15302 Vbias.n358 VGND 0.18804f
C15303 Vbias.t173 VGND 0.32014f
C15304 Vbias.n359 VGND 0.31618f
C15305 Vbias.n360 VGND 0.08903f
C15306 Vbias.n361 VGND 0.18804f
C15307 Vbias.t249 VGND 0.32014f
C15308 Vbias.n362 VGND 0.31618f
C15309 Vbias.n363 VGND 0.08903f
C15310 Vbias.n364 VGND 0.18804f
C15311 Vbias.t79 VGND 0.32014f
C15312 Vbias.n365 VGND 0.31618f
C15313 Vbias.n366 VGND 0.08903f
C15314 Vbias.n367 VGND 0.18804f
C15315 Vbias.t101 VGND 0.32014f
C15316 Vbias.n368 VGND 0.31618f
C15317 Vbias.n369 VGND 0.08903f
C15318 Vbias.n370 VGND 0.18804f
C15319 Vbias.t254 VGND 0.32014f
C15320 Vbias.n371 VGND 0.31618f
C15321 Vbias.n372 VGND 0.08903f
C15322 Vbias.n373 VGND 0.18804f
C15323 Vbias.t21 VGND 0.32014f
C15324 Vbias.n374 VGND 0.31618f
C15325 Vbias.n375 VGND 0.08903f
C15326 Vbias.n376 VGND 0.18804f
C15327 Vbias.n377 VGND 0.18804f
C15328 Vbias.t189 VGND 0.32014f
C15329 Vbias.n378 VGND 0.31618f
C15330 Vbias.t56 VGND 0.32014f
C15331 Vbias.n379 VGND 0.31618f
C15332 Vbias.n380 VGND 0.18804f
C15333 Vbias.n381 VGND 0.25661f
C15334 Vbias.n382 VGND 0.34709f
C15335 Vbias.n383 VGND 0.08903f
C15336 Vbias.n384 VGND 0.18804f
C15337 Vbias.n385 VGND 0.99957f
C15338 Vbias.n386 VGND 0.18804f
C15339 Vbias.n387 VGND 0.99957f
C15340 Vbias.n388 VGND 0.99957f
C15341 Vbias.n389 VGND 0.99957f
C15342 Vbias.t8 VGND 0.32014f
C15343 Vbias.n390 VGND 0.31618f
C15344 Vbias.n391 VGND 0.08903f
C15345 Vbias.n392 VGND 0.18804f
C15346 Vbias.n393 VGND 0.18804f
C15347 Vbias.n394 VGND 0.08903f
C15348 Vbias.n395 VGND 0.33651f
C15349 Vbias.n396 VGND 0.34709f
C15350 Vbias.n397 VGND 0.25661f
C15351 Vbias.n398 VGND 0.18804f
C15352 Vbias.t137 VGND 0.32014f
C15353 Vbias.n399 VGND 0.31618f
C15354 Vbias.n400 VGND 0.25661f
C15355 Vbias.n401 VGND 0.18804f
C15356 Vbias.t109 VGND 0.32014f
C15357 Vbias.n402 VGND 0.31618f
C15358 Vbias.n403 VGND 0.25661f
C15359 Vbias.n404 VGND 0.18804f
C15360 Vbias.t218 VGND 0.32014f
C15361 Vbias.n405 VGND 0.31618f
C15362 Vbias.n406 VGND 0.25661f
C15363 Vbias.n407 VGND 0.18804f
C15364 Vbias.t197 VGND 0.32014f
C15365 Vbias.n408 VGND 0.31618f
C15366 Vbias.n409 VGND 0.25661f
C15367 Vbias.n410 VGND 0.18804f
C15368 Vbias.t106 VGND 0.32014f
C15369 Vbias.n411 VGND 0.31618f
C15370 Vbias.n412 VGND 0.25661f
C15371 Vbias.n413 VGND 0.18804f
C15372 Vbias.t34 VGND 0.32014f
C15373 Vbias.n414 VGND 0.31618f
C15374 Vbias.n415 VGND 0.25661f
C15375 Vbias.n416 VGND 0.18804f
C15376 Vbias.t14 VGND 0.32014f
C15377 Vbias.n417 VGND 0.31618f
C15378 Vbias.n418 VGND 0.25661f
C15379 Vbias.n419 VGND 0.18804f
C15380 Vbias.t179 VGND 0.32014f
C15381 Vbias.n420 VGND 0.31618f
C15382 Vbias.n421 VGND 0.25661f
C15383 Vbias.n422 VGND 0.18804f
C15384 Vbias.t96 VGND 0.32014f
C15385 Vbias.n423 VGND 0.31618f
C15386 Vbias.n424 VGND 0.25661f
C15387 Vbias.n425 VGND 0.18804f
C15388 Vbias.t10 VGND 0.32014f
C15389 Vbias.n426 VGND 0.31618f
C15390 Vbias.n427 VGND 0.25661f
C15391 Vbias.n428 VGND 0.18804f
C15392 Vbias.t177 VGND 0.32014f
C15393 Vbias.n429 VGND 0.31618f
C15394 Vbias.n430 VGND 0.25661f
C15395 Vbias.n431 VGND 0.18804f
C15396 Vbias.t169 VGND 0.32014f
C15397 Vbias.n432 VGND 0.31618f
C15398 Vbias.n433 VGND 0.25661f
C15399 Vbias.n434 VGND 0.18804f
C15400 Vbias.t74 VGND 0.32014f
C15401 Vbias.n435 VGND 0.31618f
C15402 Vbias.n436 VGND 0.25661f
C15403 Vbias.n437 VGND 0.18804f
C15404 Vbias.n438 VGND 0.254f
C15405 Vbias.n439 VGND 0.34709f
C15406 Vbias.n440 VGND 0.33651f
C15407 Vbias.n441 VGND 0.08642f
C15408 Vbias.n442 VGND 0.18804f
C15409 Vbias.n443 VGND 0.08903f
C15410 Vbias.n444 VGND 0.33651f
C15411 Vbias.n445 VGND 0.33651f
C15412 Vbias.n446 VGND 0.08903f
C15413 Vbias.n447 VGND 0.18804f
C15414 Vbias.n448 VGND 0.18804f
C15415 Vbias.n449 VGND 0.08903f
C15416 Vbias.n450 VGND 0.33651f
C15417 Vbias.n451 VGND 0.33651f
C15418 Vbias.n452 VGND 0.08903f
C15419 Vbias.n453 VGND 0.18804f
C15420 Vbias.n454 VGND 0.18804f
C15421 Vbias.n455 VGND 0.08903f
C15422 Vbias.n456 VGND 0.33651f
C15423 Vbias.n457 VGND 0.33651f
C15424 Vbias.n458 VGND 0.08903f
C15425 Vbias.n459 VGND 0.18804f
C15426 Vbias.n460 VGND 0.18804f
C15427 Vbias.n461 VGND 0.08903f
C15428 Vbias.n462 VGND 0.33651f
C15429 Vbias.n463 VGND 0.33651f
C15430 Vbias.n464 VGND 0.08903f
C15431 Vbias.n465 VGND 0.18804f
C15432 Vbias.n466 VGND 0.18804f
C15433 Vbias.n467 VGND 0.08903f
C15434 Vbias.n468 VGND 0.33651f
C15435 Vbias.n469 VGND 0.33651f
C15436 Vbias.n470 VGND 0.08903f
C15437 Vbias.n471 VGND 0.18804f
C15438 Vbias.n472 VGND 0.18804f
C15439 Vbias.n473 VGND 0.08903f
C15440 Vbias.n474 VGND 0.33651f
C15441 Vbias.n475 VGND 0.33651f
C15442 Vbias.n476 VGND 0.08903f
C15443 Vbias.n477 VGND 0.18804f
C15444 Vbias.n478 VGND 0.18804f
C15445 Vbias.n479 VGND 0.08903f
C15446 Vbias.n480 VGND 0.33651f
C15447 Vbias.n481 VGND 0.33651f
C15448 Vbias.n482 VGND 0.08903f
C15449 Vbias.n483 VGND 0.18804f
C15450 Vbias.n484 VGND 0.18804f
C15451 Vbias.n485 VGND 0.08903f
C15452 Vbias.n486 VGND 0.33651f
C15453 Vbias.n487 VGND 0.33651f
C15454 Vbias.n488 VGND 0.08903f
C15455 Vbias.n489 VGND 0.18804f
C15456 Vbias.n490 VGND 0.18804f
C15457 Vbias.n491 VGND 0.08903f
C15458 Vbias.n492 VGND 0.33651f
C15459 Vbias.n493 VGND 0.33651f
C15460 Vbias.n494 VGND 0.08903f
C15461 Vbias.n495 VGND 0.18804f
C15462 Vbias.n496 VGND 0.18804f
C15463 Vbias.n497 VGND 0.08903f
C15464 Vbias.n498 VGND 0.33651f
C15465 Vbias.n499 VGND 0.33651f
C15466 Vbias.n500 VGND 0.08903f
C15467 Vbias.n501 VGND 0.18804f
C15468 Vbias.n502 VGND 0.18804f
C15469 Vbias.n503 VGND 0.08903f
C15470 Vbias.n504 VGND 0.33651f
C15471 Vbias.n505 VGND 0.33651f
C15472 Vbias.n506 VGND 0.08903f
C15473 Vbias.n507 VGND 0.18804f
C15474 Vbias.n508 VGND 0.18804f
C15475 Vbias.n509 VGND 0.08903f
C15476 Vbias.n510 VGND 0.33651f
C15477 Vbias.n511 VGND 0.33651f
C15478 Vbias.n512 VGND 0.08903f
C15479 Vbias.n513 VGND 0.18804f
C15480 Vbias.n514 VGND 0.18804f
C15481 Vbias.n515 VGND 0.08903f
C15482 Vbias.n516 VGND 0.33651f
C15483 Vbias.n517 VGND 0.33651f
C15484 Vbias.n518 VGND 0.08903f
C15485 Vbias.n519 VGND 0.18804f
C15486 Vbias.t170 VGND 0.32014f
C15487 Vbias.n520 VGND 0.31618f
C15488 Vbias.n521 VGND 0.08903f
C15489 Vbias.n522 VGND 0.18804f
C15490 Vbias.n523 VGND 0.18804f
C15491 Vbias.n524 VGND 0.08903f
C15492 Vbias.n525 VGND 0.33651f
C15493 Vbias.n526 VGND 0.33651f
C15494 Vbias.n527 VGND 0.33651f
C15495 Vbias.n528 VGND 0.08903f
C15496 Vbias.n529 VGND 0.18804f
C15497 Vbias.n530 VGND 0.18804f
C15498 Vbias.n531 VGND 0.08903f
C15499 Vbias.n532 VGND 0.33651f
C15500 Vbias.n533 VGND 0.33651f
C15501 Vbias.n534 VGND 0.08903f
C15502 Vbias.n535 VGND 0.18804f
C15503 Vbias.t73 VGND 0.32014f
C15504 Vbias.n536 VGND 0.31618f
C15505 Vbias.n537 VGND 0.08903f
C15506 Vbias.n538 VGND 0.18804f
C15507 Vbias.t42 VGND 0.32014f
C15508 Vbias.n539 VGND 0.31618f
C15509 Vbias.n540 VGND 0.08903f
C15510 Vbias.n541 VGND 0.18804f
C15511 Vbias.t154 VGND 0.32014f
C15512 Vbias.n542 VGND 0.31618f
C15513 Vbias.n543 VGND 0.08903f
C15514 Vbias.n544 VGND 0.18804f
C15515 Vbias.t129 VGND 0.32014f
C15516 Vbias.n545 VGND 0.31618f
C15517 Vbias.n546 VGND 0.08903f
C15518 Vbias.n547 VGND 0.18804f
C15519 Vbias.t38 VGND 0.32014f
C15520 Vbias.n548 VGND 0.31618f
C15521 Vbias.n549 VGND 0.08903f
C15522 Vbias.n550 VGND 0.18804f
C15523 Vbias.t226 VGND 0.32014f
C15524 Vbias.n551 VGND 0.31618f
C15525 Vbias.n552 VGND 0.08903f
C15526 Vbias.n553 VGND 0.18804f
C15527 Vbias.t204 VGND 0.32014f
C15528 Vbias.n554 VGND 0.31618f
C15529 Vbias.n555 VGND 0.08903f
C15530 Vbias.n556 VGND 0.18804f
C15531 Vbias.t111 VGND 0.32014f
C15532 Vbias.n557 VGND 0.31618f
C15533 Vbias.n558 VGND 0.08903f
C15534 Vbias.n559 VGND 0.18804f
C15535 Vbias.t29 VGND 0.32014f
C15536 Vbias.n560 VGND 0.31618f
C15537 Vbias.n561 VGND 0.08903f
C15538 Vbias.n562 VGND 0.18804f
C15539 Vbias.t201 VGND 0.32014f
C15540 Vbias.n563 VGND 0.31618f
C15541 Vbias.n564 VGND 0.08903f
C15542 Vbias.n565 VGND 0.18804f
C15543 Vbias.t110 VGND 0.32014f
C15544 Vbias.n566 VGND 0.31618f
C15545 Vbias.n567 VGND 0.08903f
C15546 Vbias.n568 VGND 0.18804f
C15547 Vbias.t98 VGND 0.32014f
C15548 Vbias.n569 VGND 0.31618f
C15549 Vbias.n570 VGND 0.08903f
C15550 Vbias.n571 VGND 0.18804f
C15551 Vbias.t257 VGND 0.32014f
C15552 Vbias.n572 VGND 0.31618f
C15553 Vbias.n573 VGND 0.08903f
C15554 Vbias.n574 VGND 0.18804f
C15555 Vbias.n575 VGND 0.08642f
C15556 Vbias.n576 VGND 0.33651f
C15557 Vbias.n577 VGND 0.33651f
C15558 Vbias.n578 VGND 0.08642f
C15559 Vbias.n579 VGND 0.18804f
C15560 Vbias.n580 VGND 0.08903f
C15561 Vbias.n581 VGND 0.33651f
C15562 Vbias.n582 VGND 0.33651f
C15563 Vbias.n583 VGND 0.08903f
C15564 Vbias.n584 VGND 0.18804f
C15565 Vbias.n585 VGND 0.18804f
C15566 Vbias.n586 VGND 0.08903f
C15567 Vbias.n587 VGND 0.33651f
C15568 Vbias.n588 VGND 0.33651f
C15569 Vbias.n589 VGND 0.08903f
C15570 Vbias.n590 VGND 0.18804f
C15571 Vbias.n591 VGND 0.18804f
C15572 Vbias.n592 VGND 0.08903f
C15573 Vbias.n593 VGND 0.33651f
C15574 Vbias.n594 VGND 0.33651f
C15575 Vbias.n595 VGND 0.08903f
C15576 Vbias.n596 VGND 0.18804f
C15577 Vbias.n597 VGND 0.18804f
C15578 Vbias.n598 VGND 0.08903f
C15579 Vbias.n599 VGND 0.33651f
C15580 Vbias.n600 VGND 0.33651f
C15581 Vbias.n601 VGND 0.08903f
C15582 Vbias.n602 VGND 0.18804f
C15583 Vbias.n603 VGND 0.18804f
C15584 Vbias.n604 VGND 0.08903f
C15585 Vbias.n605 VGND 0.33651f
C15586 Vbias.n606 VGND 0.33651f
C15587 Vbias.n607 VGND 0.08903f
C15588 Vbias.n608 VGND 0.18804f
C15589 Vbias.n609 VGND 0.18804f
C15590 Vbias.n610 VGND 0.08903f
C15591 Vbias.n611 VGND 0.33651f
C15592 Vbias.n612 VGND 0.33651f
C15593 Vbias.n613 VGND 0.08903f
C15594 Vbias.n614 VGND 0.18804f
C15595 Vbias.n615 VGND 0.18804f
C15596 Vbias.n616 VGND 0.08903f
C15597 Vbias.n617 VGND 0.33651f
C15598 Vbias.n618 VGND 0.33651f
C15599 Vbias.n619 VGND 0.08903f
C15600 Vbias.n620 VGND 0.18804f
C15601 Vbias.n621 VGND 0.18804f
C15602 Vbias.n622 VGND 0.08903f
C15603 Vbias.n623 VGND 0.33651f
C15604 Vbias.n624 VGND 0.33651f
C15605 Vbias.n625 VGND 0.08903f
C15606 Vbias.n626 VGND 0.18804f
C15607 Vbias.n627 VGND 0.18804f
C15608 Vbias.n628 VGND 0.08903f
C15609 Vbias.n629 VGND 0.33651f
C15610 Vbias.n630 VGND 0.33651f
C15611 Vbias.n631 VGND 0.08903f
C15612 Vbias.n632 VGND 0.18804f
C15613 Vbias.n633 VGND 0.18804f
C15614 Vbias.n634 VGND 0.08903f
C15615 Vbias.n635 VGND 0.33651f
C15616 Vbias.n636 VGND 0.33651f
C15617 Vbias.n637 VGND 0.08903f
C15618 Vbias.n638 VGND 0.18804f
C15619 Vbias.n639 VGND 0.18804f
C15620 Vbias.n640 VGND 0.08903f
C15621 Vbias.n641 VGND 0.33651f
C15622 Vbias.n642 VGND 0.33651f
C15623 Vbias.n643 VGND 0.08903f
C15624 Vbias.n644 VGND 0.18804f
C15625 Vbias.n645 VGND 0.18804f
C15626 Vbias.n646 VGND 0.08903f
C15627 Vbias.n647 VGND 0.33651f
C15628 Vbias.n648 VGND 0.33651f
C15629 Vbias.n649 VGND 0.08903f
C15630 Vbias.n650 VGND 0.18804f
C15631 Vbias.n651 VGND 0.18804f
C15632 Vbias.n652 VGND 0.08903f
C15633 Vbias.n653 VGND 0.33651f
C15634 Vbias.n654 VGND 0.33651f
C15635 Vbias.n655 VGND 0.08903f
C15636 Vbias.n656 VGND 0.18804f
C15637 Vbias.t84 VGND 0.32014f
C15638 Vbias.n657 VGND 0.31618f
C15639 Vbias.n658 VGND 0.08903f
C15640 Vbias.n659 VGND 0.18804f
C15641 Vbias.t245 VGND 0.32014f
C15642 Vbias.n660 VGND 0.31618f
C15643 Vbias.n661 VGND 0.08903f
C15644 Vbias.n662 VGND 0.18804f
C15645 Vbias.n663 VGND 0.99957f
C15646 Vbias.n664 VGND 0.99957f
C15647 Vbias.n665 VGND 0.99957f
C15648 Vbias.t160 VGND 0.32014f
C15649 Vbias.n666 VGND 0.31618f
C15650 Vbias.n667 VGND 0.08903f
C15651 Vbias.n668 VGND 0.18804f
C15652 Vbias.t68 VGND 0.32014f
C15653 Vbias.n669 VGND 0.31618f
C15654 Vbias.n670 VGND 0.08903f
C15655 Vbias.n671 VGND 0.18804f
C15656 Vbias.n672 VGND 0.99957f
C15657 Vbias.t250 VGND 0.32014f
C15658 Vbias.n673 VGND 0.31618f
C15659 Vbias.n674 VGND 0.33651f
C15660 Vbias.n675 VGND 0.08903f
C15661 Vbias.n676 VGND 0.18804f
C15662 Vbias.n677 VGND 0.99957f
C15663 Vbias.t171 VGND 0.32014f
C15664 Vbias.n678 VGND 0.31618f
C15665 Vbias.n679 VGND 0.08903f
C15666 Vbias.n680 VGND 0.18804f
C15667 Vbias.n681 VGND 0.99957f
C15668 Vbias.n682 VGND 0.99957f
C15669 Vbias.n683 VGND 0.99957f
C15670 Vbias.n684 VGND 0.18804f
C15671 Vbias.n685 VGND 0.18804f
C15672 Vbias.n686 VGND 0.08903f
C15673 Vbias.n687 VGND 0.33651f
C15674 Vbias.n688 VGND 0.33651f
C15675 Vbias.n689 VGND 0.08903f
C15676 Vbias.n690 VGND 0.18804f
C15677 Vbias.n691 VGND 0.18804f
C15678 Vbias.n692 VGND 0.08903f
C15679 Vbias.n693 VGND 0.33651f
C15680 Vbias.n694 VGND 0.33651f
C15681 Vbias.n695 VGND 0.33651f
C15682 Vbias.n696 VGND 0.08903f
C15683 Vbias.n697 VGND 0.18804f
C15684 Vbias.t199 VGND 0.32014f
C15685 Vbias.n698 VGND 0.31618f
C15686 Vbias.n699 VGND 0.08903f
C15687 Vbias.n700 VGND 0.18804f
C15688 Vbias.n701 VGND 0.18804f
C15689 Vbias.n702 VGND 0.08903f
C15690 Vbias.n703 VGND 0.33651f
C15691 Vbias.n704 VGND 0.33651f
C15692 Vbias.n705 VGND 0.08903f
C15693 Vbias.n706 VGND 0.18804f
C15694 Vbias.n707 VGND 0.18804f
C15695 Vbias.n708 VGND 0.08903f
C15696 Vbias.n709 VGND 0.33651f
C15697 Vbias.n710 VGND 0.33651f
C15698 Vbias.n711 VGND 0.08903f
C15699 Vbias.n712 VGND 0.18804f
C15700 Vbias.n713 VGND 0.18804f
C15701 Vbias.n714 VGND 0.08903f
C15702 Vbias.n715 VGND 0.33651f
C15703 Vbias.n716 VGND 0.33651f
C15704 Vbias.n717 VGND 0.08903f
C15705 Vbias.n718 VGND 0.18804f
C15706 Vbias.n719 VGND 0.18804f
C15707 Vbias.n720 VGND 0.08903f
C15708 Vbias.n721 VGND 0.33651f
C15709 Vbias.n722 VGND 0.33651f
C15710 Vbias.n723 VGND 0.08903f
C15711 Vbias.n724 VGND 0.18804f
C15712 Vbias.n725 VGND 0.18804f
C15713 Vbias.n726 VGND 0.08903f
C15714 Vbias.n727 VGND 0.33651f
C15715 Vbias.n728 VGND 0.33651f
C15716 Vbias.n729 VGND 0.08903f
C15717 Vbias.n730 VGND 0.18804f
C15718 Vbias.n731 VGND 0.18804f
C15719 Vbias.n732 VGND 0.08903f
C15720 Vbias.n733 VGND 0.33651f
C15721 Vbias.n734 VGND 0.33651f
C15722 Vbias.n735 VGND 0.08903f
C15723 Vbias.n736 VGND 0.18804f
C15724 Vbias.n737 VGND 0.18804f
C15725 Vbias.n738 VGND 0.08903f
C15726 Vbias.n739 VGND 0.33651f
C15727 Vbias.n740 VGND 0.33651f
C15728 Vbias.n741 VGND 0.08903f
C15729 Vbias.n742 VGND 0.18804f
C15730 Vbias.n743 VGND 0.18804f
C15731 Vbias.n744 VGND 0.08903f
C15732 Vbias.n745 VGND 0.33651f
C15733 Vbias.n746 VGND 0.33651f
C15734 Vbias.n747 VGND 0.08903f
C15735 Vbias.n748 VGND 0.18804f
C15736 Vbias.n749 VGND 0.18804f
C15737 Vbias.n750 VGND 0.08903f
C15738 Vbias.n751 VGND 0.33651f
C15739 Vbias.n752 VGND 0.33651f
C15740 Vbias.n753 VGND 0.08903f
C15741 Vbias.n754 VGND 0.18804f
C15742 Vbias.n755 VGND 0.18804f
C15743 Vbias.n756 VGND 0.08903f
C15744 Vbias.n757 VGND 0.33651f
C15745 Vbias.n758 VGND 0.33651f
C15746 Vbias.n759 VGND 0.08903f
C15747 Vbias.n760 VGND 0.18804f
C15748 Vbias.n761 VGND 0.18804f
C15749 Vbias.n762 VGND 0.08903f
C15750 Vbias.n763 VGND 0.33651f
C15751 Vbias.n764 VGND 0.33651f
C15752 Vbias.n765 VGND 0.08903f
C15753 Vbias.n766 VGND 0.18804f
C15754 Vbias.n767 VGND 0.18804f
C15755 Vbias.n768 VGND 0.08903f
C15756 Vbias.n769 VGND 0.33651f
C15757 Vbias.n770 VGND 0.33651f
C15758 Vbias.n771 VGND 0.08903f
C15759 Vbias.n772 VGND 0.18804f
C15760 Vbias.n773 VGND 0.18804f
C15761 Vbias.n774 VGND 0.08903f
C15762 Vbias.n775 VGND 0.33651f
C15763 Vbias.n776 VGND 0.33651f
C15764 Vbias.n777 VGND 0.08903f
C15765 Vbias.n778 VGND 0.18804f
C15766 Vbias.n779 VGND 0.08642f
C15767 Vbias.n780 VGND 0.33651f
C15768 Vbias.n781 VGND 0.33651f
C15769 Vbias.n782 VGND 0.33651f
C15770 Vbias.n783 VGND 0.08642f
C15771 Vbias.t190 VGND 0.32014f
C15772 Vbias.n784 VGND 0.31618f
C15773 Vbias.n785 VGND 0.08903f
C15774 Vbias.n786 VGND 0.18804f
C15775 Vbias.t32 VGND 0.32014f
C15776 Vbias.n787 VGND 0.31618f
C15777 Vbias.n788 VGND 0.08903f
C15778 Vbias.n789 VGND 0.18804f
C15779 Vbias.t43 VGND 0.32014f
C15780 Vbias.n790 VGND 0.31618f
C15781 Vbias.n791 VGND 0.08903f
C15782 Vbias.n792 VGND 0.18804f
C15783 Vbias.t130 VGND 0.32014f
C15784 Vbias.n793 VGND 0.31618f
C15785 Vbias.n794 VGND 0.08903f
C15786 Vbias.n795 VGND 0.18804f
C15787 Vbias.t216 VGND 0.32014f
C15788 Vbias.n796 VGND 0.31618f
C15789 Vbias.n797 VGND 0.08903f
C15790 Vbias.n798 VGND 0.18804f
C15791 Vbias.t45 VGND 0.32014f
C15792 Vbias.n799 VGND 0.31618f
C15793 Vbias.n800 VGND 0.08903f
C15794 Vbias.n801 VGND 0.18804f
C15795 Vbias.t133 VGND 0.32014f
C15796 Vbias.n802 VGND 0.31618f
C15797 Vbias.n803 VGND 0.08903f
C15798 Vbias.n804 VGND 0.18804f
C15799 Vbias.t158 VGND 0.32014f
C15800 Vbias.n805 VGND 0.31618f
C15801 Vbias.n806 VGND 0.08903f
C15802 Vbias.n807 VGND 0.18804f
C15803 Vbias.t231 VGND 0.32014f
C15804 Vbias.n808 VGND 0.31618f
C15805 Vbias.n809 VGND 0.08903f
C15806 Vbias.n810 VGND 0.18804f
C15807 Vbias.t60 VGND 0.32014f
C15808 Vbias.n811 VGND 0.31618f
C15809 Vbias.n812 VGND 0.08903f
C15810 Vbias.n813 VGND 0.18804f
C15811 Vbias.t85 VGND 0.32014f
C15812 Vbias.n814 VGND 0.31618f
C15813 Vbias.n815 VGND 0.08903f
C15814 Vbias.n816 VGND 0.18804f
C15815 Vbias.t237 VGND 0.32014f
C15816 Vbias.n817 VGND 0.31618f
C15817 Vbias.n818 VGND 0.08903f
C15818 Vbias.n819 VGND 0.18804f
C15819 Vbias.t258 VGND 0.32014f
C15820 Vbias.n820 VGND 0.31618f
C15821 Vbias.n821 VGND 0.08903f
C15822 Vbias.n822 VGND 0.18804f
C15823 Vbias.n823 VGND 0.18804f
C15824 Vbias.n824 VGND 0.08903f
C15825 Vbias.n825 VGND 0.33651f
C15826 Vbias.n826 VGND 0.33651f
C15827 Vbias.n827 VGND 0.08903f
C15828 Vbias.n828 VGND 0.18804f
C15829 Vbias.n829 VGND 0.18804f
C15830 Vbias.n830 VGND 0.08903f
C15831 Vbias.n831 VGND 0.33651f
C15832 Vbias.n832 VGND 0.33651f
C15833 Vbias.n833 VGND 0.08903f
C15834 Vbias.n834 VGND 0.18804f
C15835 Vbias.n835 VGND 0.18804f
C15836 Vbias.n836 VGND 0.08903f
C15837 Vbias.n837 VGND 0.33651f
C15838 Vbias.n838 VGND 0.33651f
C15839 Vbias.n839 VGND 0.08903f
C15840 Vbias.n840 VGND 0.18804f
C15841 Vbias.n841 VGND 0.18804f
C15842 Vbias.n842 VGND 0.08903f
C15843 Vbias.n843 VGND 0.33651f
C15844 Vbias.n844 VGND 0.33651f
C15845 Vbias.n845 VGND 0.08903f
C15846 Vbias.n846 VGND 0.18804f
C15847 Vbias.n847 VGND 0.18804f
C15848 Vbias.n848 VGND 0.08903f
C15849 Vbias.n849 VGND 0.33651f
C15850 Vbias.n850 VGND 0.33651f
C15851 Vbias.n851 VGND 0.08903f
C15852 Vbias.n852 VGND 0.18804f
C15853 Vbias.n853 VGND 0.18804f
C15854 Vbias.n854 VGND 0.08903f
C15855 Vbias.n855 VGND 0.33651f
C15856 Vbias.n856 VGND 0.33651f
C15857 Vbias.n857 VGND 0.08903f
C15858 Vbias.n858 VGND 0.18804f
C15859 Vbias.n859 VGND 0.18804f
C15860 Vbias.n860 VGND 0.08903f
C15861 Vbias.n861 VGND 0.33651f
C15862 Vbias.n862 VGND 0.33651f
C15863 Vbias.n863 VGND 0.08903f
C15864 Vbias.n864 VGND 0.18804f
C15865 Vbias.n865 VGND 0.18804f
C15866 Vbias.n866 VGND 0.08903f
C15867 Vbias.n867 VGND 0.33651f
C15868 Vbias.n868 VGND 0.33651f
C15869 Vbias.n869 VGND 0.08903f
C15870 Vbias.n870 VGND 0.18804f
C15871 Vbias.n871 VGND 0.18804f
C15872 Vbias.n872 VGND 0.08903f
C15873 Vbias.n873 VGND 0.33651f
C15874 Vbias.n874 VGND 0.33651f
C15875 Vbias.n875 VGND 0.08903f
C15876 Vbias.n876 VGND 0.18804f
C15877 Vbias.n877 VGND 0.18804f
C15878 Vbias.n878 VGND 0.08903f
C15879 Vbias.n879 VGND 0.33651f
C15880 Vbias.n880 VGND 0.33651f
C15881 Vbias.n881 VGND 0.08903f
C15882 Vbias.n882 VGND 0.18804f
C15883 Vbias.n883 VGND 0.18804f
C15884 Vbias.n884 VGND 0.08903f
C15885 Vbias.n885 VGND 0.33651f
C15886 Vbias.n886 VGND 0.33651f
C15887 Vbias.n887 VGND 0.08903f
C15888 Vbias.n888 VGND 0.18804f
C15889 Vbias.n889 VGND 0.18804f
C15890 Vbias.n890 VGND 0.08903f
C15891 Vbias.n891 VGND 0.33651f
C15892 Vbias.n892 VGND 0.33651f
C15893 Vbias.n893 VGND 0.08903f
C15894 Vbias.n894 VGND 0.18804f
C15895 Vbias.n895 VGND 0.18804f
C15896 Vbias.n896 VGND 0.08903f
C15897 Vbias.n897 VGND 0.33651f
C15898 Vbias.n898 VGND 0.33651f
C15899 Vbias.n899 VGND 0.08903f
C15900 Vbias.n900 VGND 0.18804f
C15901 Vbias.t193 VGND 0.32014f
C15902 Vbias.n901 VGND 0.31618f
C15903 Vbias.n902 VGND 0.08642f
C15904 Vbias.n903 VGND 0.18804f
C15905 Vbias.n904 VGND 0.08903f
C15906 Vbias.n905 VGND 0.33651f
C15907 Vbias.n906 VGND 0.33651f
C15908 Vbias.n907 VGND 0.08903f
C15909 Vbias.n908 VGND 0.18804f
C15910 Vbias.n909 VGND 0.08642f
C15911 Vbias.n910 VGND 0.33651f
C15912 Vbias.n911 VGND 0.33651f
C15913 Vbias.n912 VGND 0.33373f
C15914 Vbias.n913 VGND 0.08642f
C15915 Vbias.n914 VGND 0.18804f
C15916 Vbias.n915 VGND 0.08903f
C15917 Vbias.n916 VGND 0.33373f
C15918 Vbias.n917 VGND 0.04509f
C15919 Vbias.n918 VGND 0.18804f
C15920 Vbias.n919 VGND 0.18804f
C15921 Vbias.n920 VGND 0.04509f
C15922 Vbias.n921 VGND 0.33373f
C15923 Vbias.n922 VGND 0.08903f
C15924 Vbias.n923 VGND 0.18804f
C15925 Vbias.n924 VGND 0.18804f
C15926 Vbias.n925 VGND 0.08903f
C15927 Vbias.n926 VGND 0.33373f
C15928 Vbias.n927 VGND 0.04509f
C15929 Vbias.n928 VGND 0.18804f
C15930 Vbias.n929 VGND 0.18804f
C15931 Vbias.n930 VGND 0.04509f
C15932 Vbias.n931 VGND 0.33373f
C15933 Vbias.n932 VGND 0.08903f
C15934 Vbias.n933 VGND 0.18804f
C15935 Vbias.n934 VGND 0.18804f
C15936 Vbias.n935 VGND 0.08903f
C15937 Vbias.n936 VGND 0.33373f
C15938 Vbias.n937 VGND 0.04509f
C15939 Vbias.n938 VGND 0.18804f
C15940 Vbias.n939 VGND 0.18804f
C15941 Vbias.n940 VGND 0.04509f
C15942 Vbias.n941 VGND 0.33373f
C15943 Vbias.n942 VGND 0.08903f
C15944 Vbias.n943 VGND 0.18804f
C15945 Vbias.n944 VGND 0.18804f
C15946 Vbias.n945 VGND 0.08903f
C15947 Vbias.n946 VGND 0.33373f
C15948 Vbias.n947 VGND 0.04509f
C15949 Vbias.n948 VGND 0.18804f
C15950 Vbias.n949 VGND 0.18804f
C15951 Vbias.n950 VGND 0.04509f
C15952 Vbias.n951 VGND 0.33373f
C15953 Vbias.n952 VGND 0.08903f
C15954 Vbias.n953 VGND 0.18804f
C15955 Vbias.n954 VGND 0.18804f
C15956 Vbias.n955 VGND 0.08903f
C15957 Vbias.n956 VGND 0.33373f
C15958 Vbias.n957 VGND 0.04509f
C15959 Vbias.n958 VGND 0.18804f
C15960 Vbias.n959 VGND 0.18804f
C15961 Vbias.n960 VGND 0.04509f
C15962 Vbias.n961 VGND 0.33373f
C15963 Vbias.n962 VGND 0.08903f
C15964 Vbias.n963 VGND 0.18804f
C15965 Vbias.n964 VGND 0.18804f
C15966 Vbias.n965 VGND 0.08903f
C15967 Vbias.n966 VGND 0.33373f
C15968 Vbias.n967 VGND 0.04509f
C15969 Vbias.n968 VGND 0.18804f
C15970 Vbias.n969 VGND 0.18804f
C15971 Vbias.n970 VGND 0.04509f
C15972 Vbias.n971 VGND 0.33373f
C15973 Vbias.n972 VGND 0.08903f
C15974 Vbias.n973 VGND 0.18804f
C15975 Vbias.n974 VGND 0.18804f
C15976 Vbias.n975 VGND 0.08903f
C15977 Vbias.n976 VGND 0.33373f
C15978 Vbias.n977 VGND 0.04509f
C15979 Vbias.n978 VGND 0.18804f
C15980 Vbias.n979 VGND 0.18804f
C15981 Vbias.n980 VGND 0.04509f
C15982 Vbias.n981 VGND 0.33373f
C15983 Vbias.n982 VGND 0.33651f
C15984 Vbias.n983 VGND 0.08903f
C15985 Vbias.n984 VGND 0.18804f
C15986 Vbias.n985 VGND 0.18804f
C15987 Vbias.n986 VGND 0.08903f
C15988 Vbias.n987 VGND 0.33651f
C15989 Vbias.n988 VGND 0.33373f
C15990 Vbias.n989 VGND 0.04509f
C15991 Vbias.n990 VGND 0.18804f
C15992 Vbias.n991 VGND 1.16253f
C15993 Vbias.t1 VGND 0.06542f
C15994 Vbias.t0 VGND 0.06542f
C15995 Vbias.n992 VGND 0.44073f
C15996 Vbias.t4 VGND 0.06542f
C15997 Vbias.t5 VGND 0.06542f
C15998 Vbias.n993 VGND 0.44073f
C15999 Vbias.n994 VGND 1.3303f
C16000 Vbias.t3 VGND 0.30514f
C16001 Vbias.t2 VGND 1.1998f
C16002 Vbias.n995 VGND 2.22128f
C16003 Vbias.n996 VGND 0.85437f
C16004 Vbias.n997 VGND 2.00052f
C16005 XThR.Tn[14].t0 VGND 0.02436f
C16006 XThR.Tn[14].t1 VGND 0.02436f
C16007 XThR.Tn[14].n0 VGND 0.07395f
C16008 XThR.Tn[14].t2 VGND 0.02436f
C16009 XThR.Tn[14].t3 VGND 0.02436f
C16010 XThR.Tn[14].n1 VGND 0.05414f
C16011 XThR.Tn[14].n2 VGND 0.24618f
C16012 XThR.Tn[14].t6 VGND 0.01583f
C16013 XThR.Tn[14].t7 VGND 0.01583f
C16014 XThR.Tn[14].n3 VGND 0.03948f
C16015 XThR.Tn[14].t4 VGND 0.01583f
C16016 XThR.Tn[14].t5 VGND 0.01583f
C16017 XThR.Tn[14].n4 VGND 0.03166f
C16018 XThR.Tn[14].n5 VGND 0.07301f
C16019 XThR.Tn[14].t69 VGND 0.01904f
C16020 XThR.Tn[14].t62 VGND 0.02084f
C16021 XThR.Tn[14].n6 VGND 0.0509f
C16022 XThR.Tn[14].n7 VGND 0.09778f
C16023 XThR.Tn[14].t24 VGND 0.01904f
C16024 XThR.Tn[14].t13 VGND 0.02084f
C16025 XThR.Tn[14].n8 VGND 0.0509f
C16026 XThR.Tn[14].t28 VGND 0.01897f
C16027 XThR.Tn[14].t60 VGND 0.02078f
C16028 XThR.Tn[14].n9 VGND 0.05296f
C16029 XThR.Tn[14].n10 VGND 0.03721f
C16030 XThR.Tn[14].n11 VGND 0.0068f
C16031 XThR.Tn[14].n12 VGND 0.11939f
C16032 XThR.Tn[14].t64 VGND 0.01904f
C16033 XThR.Tn[14].t54 VGND 0.02084f
C16034 XThR.Tn[14].n13 VGND 0.0509f
C16035 XThR.Tn[14].t67 VGND 0.01897f
C16036 XThR.Tn[14].t34 VGND 0.02078f
C16037 XThR.Tn[14].n14 VGND 0.05296f
C16038 XThR.Tn[14].n15 VGND 0.03721f
C16039 XThR.Tn[14].n16 VGND 0.0068f
C16040 XThR.Tn[14].n17 VGND 0.11939f
C16041 XThR.Tn[14].t14 VGND 0.01904f
C16042 XThR.Tn[14].t72 VGND 0.02084f
C16043 XThR.Tn[14].n18 VGND 0.0509f
C16044 XThR.Tn[14].t17 VGND 0.01897f
C16045 XThR.Tn[14].t52 VGND 0.02078f
C16046 XThR.Tn[14].n19 VGND 0.05296f
C16047 XThR.Tn[14].n20 VGND 0.03721f
C16048 XThR.Tn[14].n21 VGND 0.0068f
C16049 XThR.Tn[14].n22 VGND 0.11939f
C16050 XThR.Tn[14].t44 VGND 0.01904f
C16051 XThR.Tn[14].t38 VGND 0.02084f
C16052 XThR.Tn[14].n23 VGND 0.0509f
C16053 XThR.Tn[14].t47 VGND 0.01897f
C16054 XThR.Tn[14].t18 VGND 0.02078f
C16055 XThR.Tn[14].n24 VGND 0.05296f
C16056 XThR.Tn[14].n25 VGND 0.03721f
C16057 XThR.Tn[14].n26 VGND 0.0068f
C16058 XThR.Tn[14].n27 VGND 0.11939f
C16059 XThR.Tn[14].t15 VGND 0.01904f
C16060 XThR.Tn[14].t73 VGND 0.02084f
C16061 XThR.Tn[14].n28 VGND 0.0509f
C16062 XThR.Tn[14].t21 VGND 0.01897f
C16063 XThR.Tn[14].t53 VGND 0.02078f
C16064 XThR.Tn[14].n29 VGND 0.05296f
C16065 XThR.Tn[14].n30 VGND 0.03721f
C16066 XThR.Tn[14].n31 VGND 0.0068f
C16067 XThR.Tn[14].n32 VGND 0.11939f
C16068 XThR.Tn[14].t57 VGND 0.01904f
C16069 XThR.Tn[14].t25 VGND 0.02084f
C16070 XThR.Tn[14].n33 VGND 0.0509f
C16071 XThR.Tn[14].t61 VGND 0.01897f
C16072 XThR.Tn[14].t71 VGND 0.02078f
C16073 XThR.Tn[14].n34 VGND 0.05296f
C16074 XThR.Tn[14].n35 VGND 0.03721f
C16075 XThR.Tn[14].n36 VGND 0.0068f
C16076 XThR.Tn[14].n37 VGND 0.11939f
C16077 XThR.Tn[14].t23 VGND 0.01904f
C16078 XThR.Tn[14].t19 VGND 0.02084f
C16079 XThR.Tn[14].n38 VGND 0.0509f
C16080 XThR.Tn[14].t29 VGND 0.01897f
C16081 XThR.Tn[14].t66 VGND 0.02078f
C16082 XThR.Tn[14].n39 VGND 0.05296f
C16083 XThR.Tn[14].n40 VGND 0.03721f
C16084 XThR.Tn[14].n41 VGND 0.0068f
C16085 XThR.Tn[14].n42 VGND 0.11939f
C16086 XThR.Tn[14].t27 VGND 0.01904f
C16087 XThR.Tn[14].t36 VGND 0.02084f
C16088 XThR.Tn[14].n43 VGND 0.0509f
C16089 XThR.Tn[14].t33 VGND 0.01897f
C16090 XThR.Tn[14].t16 VGND 0.02078f
C16091 XThR.Tn[14].n44 VGND 0.05296f
C16092 XThR.Tn[14].n45 VGND 0.03721f
C16093 XThR.Tn[14].n46 VGND 0.0068f
C16094 XThR.Tn[14].n47 VGND 0.11939f
C16095 XThR.Tn[14].t46 VGND 0.01904f
C16096 XThR.Tn[14].t56 VGND 0.02084f
C16097 XThR.Tn[14].n48 VGND 0.0509f
C16098 XThR.Tn[14].t50 VGND 0.01897f
C16099 XThR.Tn[14].t35 VGND 0.02078f
C16100 XThR.Tn[14].n49 VGND 0.05296f
C16101 XThR.Tn[14].n50 VGND 0.03721f
C16102 XThR.Tn[14].n51 VGND 0.0068f
C16103 XThR.Tn[14].n52 VGND 0.11939f
C16104 XThR.Tn[14].t40 VGND 0.01904f
C16105 XThR.Tn[14].t12 VGND 0.02084f
C16106 XThR.Tn[14].n53 VGND 0.0509f
C16107 XThR.Tn[14].t42 VGND 0.01897f
C16108 XThR.Tn[14].t55 VGND 0.02078f
C16109 XThR.Tn[14].n54 VGND 0.05296f
C16110 XThR.Tn[14].n55 VGND 0.03721f
C16111 XThR.Tn[14].n56 VGND 0.0068f
C16112 XThR.Tn[14].n57 VGND 0.11939f
C16113 XThR.Tn[14].t59 VGND 0.01904f
C16114 XThR.Tn[14].t49 VGND 0.02084f
C16115 XThR.Tn[14].n58 VGND 0.0509f
C16116 XThR.Tn[14].t63 VGND 0.01897f
C16117 XThR.Tn[14].t30 VGND 0.02078f
C16118 XThR.Tn[14].n59 VGND 0.05296f
C16119 XThR.Tn[14].n60 VGND 0.03721f
C16120 XThR.Tn[14].n61 VGND 0.0068f
C16121 XThR.Tn[14].n62 VGND 0.11939f
C16122 XThR.Tn[14].t26 VGND 0.01904f
C16123 XThR.Tn[14].t22 VGND 0.02084f
C16124 XThR.Tn[14].n63 VGND 0.0509f
C16125 XThR.Tn[14].t31 VGND 0.01897f
C16126 XThR.Tn[14].t68 VGND 0.02078f
C16127 XThR.Tn[14].n64 VGND 0.05296f
C16128 XThR.Tn[14].n65 VGND 0.03721f
C16129 XThR.Tn[14].n66 VGND 0.0068f
C16130 XThR.Tn[14].n67 VGND 0.11939f
C16131 XThR.Tn[14].t45 VGND 0.01904f
C16132 XThR.Tn[14].t39 VGND 0.02084f
C16133 XThR.Tn[14].n68 VGND 0.0509f
C16134 XThR.Tn[14].t48 VGND 0.01897f
C16135 XThR.Tn[14].t20 VGND 0.02078f
C16136 XThR.Tn[14].n69 VGND 0.05296f
C16137 XThR.Tn[14].n70 VGND 0.03721f
C16138 XThR.Tn[14].n71 VGND 0.0068f
C16139 XThR.Tn[14].n72 VGND 0.11939f
C16140 XThR.Tn[14].t65 VGND 0.01904f
C16141 XThR.Tn[14].t58 VGND 0.02084f
C16142 XThR.Tn[14].n73 VGND 0.0509f
C16143 XThR.Tn[14].t70 VGND 0.01897f
C16144 XThR.Tn[14].t37 VGND 0.02078f
C16145 XThR.Tn[14].n74 VGND 0.05296f
C16146 XThR.Tn[14].n75 VGND 0.03721f
C16147 XThR.Tn[14].n76 VGND 0.0068f
C16148 XThR.Tn[14].n77 VGND 0.11939f
C16149 XThR.Tn[14].t41 VGND 0.01904f
C16150 XThR.Tn[14].t51 VGND 0.02084f
C16151 XThR.Tn[14].n78 VGND 0.0509f
C16152 XThR.Tn[14].t43 VGND 0.01897f
C16153 XThR.Tn[14].t32 VGND 0.02078f
C16154 XThR.Tn[14].n79 VGND 0.05296f
C16155 XThR.Tn[14].n80 VGND 0.03721f
C16156 XThR.Tn[14].n81 VGND 0.0068f
C16157 XThR.Tn[14].n82 VGND 0.11939f
C16158 XThR.Tn[14].n83 VGND 0.1085f
C16159 XThR.Tn[14].n84 VGND 0.43586f
C16160 XThR.Tn[14].t10 VGND 0.02436f
C16161 XThR.Tn[14].t11 VGND 0.02436f
C16162 XThR.Tn[14].n85 VGND 0.05262f
C16163 XThR.Tn[14].t8 VGND 0.02436f
C16164 XThR.Tn[14].t9 VGND 0.02436f
C16165 XThR.Tn[14].n86 VGND 0.08009f
C16166 XThR.Tn[14].n87 VGND 0.22239f
C16167 XThR.Tn[14].n88 VGND 0.01096f
C16168 XThR.Tn[6].t2 VGND 0.02335f
C16169 XThR.Tn[6].t1 VGND 0.02335f
C16170 XThR.Tn[6].n0 VGND 0.05514f
C16171 XThR.Tn[6].t3 VGND 0.02335f
C16172 XThR.Tn[6].t0 VGND 0.02335f
C16173 XThR.Tn[6].n1 VGND 0.04712f
C16174 XThR.Tn[6].n2 VGND 0.16538f
C16175 XThR.Tn[6].t8 VGND 0.01517f
C16176 XThR.Tn[6].t9 VGND 0.01517f
C16177 XThR.Tn[6].n3 VGND 0.05758f
C16178 XThR.Tn[6].t11 VGND 0.01517f
C16179 XThR.Tn[6].t10 VGND 0.01517f
C16180 XThR.Tn[6].n4 VGND 0.03456f
C16181 XThR.Tn[6].n5 VGND 0.16456f
C16182 XThR.Tn[6].t7 VGND 0.01517f
C16183 XThR.Tn[6].t6 VGND 0.01517f
C16184 XThR.Tn[6].n6 VGND 0.03456f
C16185 XThR.Tn[6].n7 VGND 0.10173f
C16186 XThR.Tn[6].t4 VGND 0.01517f
C16187 XThR.Tn[6].t5 VGND 0.01517f
C16188 XThR.Tn[6].n8 VGND 0.03456f
C16189 XThR.Tn[6].n9 VGND 0.11481f
C16190 XThR.Tn[6].t62 VGND 0.01825f
C16191 XThR.Tn[6].t56 VGND 0.01998f
C16192 XThR.Tn[6].n10 VGND 0.04879f
C16193 XThR.Tn[6].n11 VGND 0.09372f
C16194 XThR.Tn[6].t20 VGND 0.01825f
C16195 XThR.Tn[6].t72 VGND 0.01998f
C16196 XThR.Tn[6].n12 VGND 0.04879f
C16197 XThR.Tn[6].t36 VGND 0.01819f
C16198 XThR.Tn[6].t68 VGND 0.01991f
C16199 XThR.Tn[6].n13 VGND 0.05076f
C16200 XThR.Tn[6].n14 VGND 0.03566f
C16201 XThR.Tn[6].n15 VGND 0.00652f
C16202 XThR.Tn[6].n16 VGND 0.11444f
C16203 XThR.Tn[6].t57 VGND 0.01825f
C16204 XThR.Tn[6].t49 VGND 0.01998f
C16205 XThR.Tn[6].n17 VGND 0.04879f
C16206 XThR.Tn[6].t14 VGND 0.01819f
C16207 XThR.Tn[6].t45 VGND 0.01991f
C16208 XThR.Tn[6].n18 VGND 0.05076f
C16209 XThR.Tn[6].n19 VGND 0.03566f
C16210 XThR.Tn[6].n20 VGND 0.00652f
C16211 XThR.Tn[6].n21 VGND 0.11444f
C16212 XThR.Tn[6].t73 VGND 0.01825f
C16213 XThR.Tn[6].t66 VGND 0.01998f
C16214 XThR.Tn[6].n22 VGND 0.04879f
C16215 XThR.Tn[6].t26 VGND 0.01819f
C16216 XThR.Tn[6].t63 VGND 0.01991f
C16217 XThR.Tn[6].n23 VGND 0.05076f
C16218 XThR.Tn[6].n24 VGND 0.03566f
C16219 XThR.Tn[6].n25 VGND 0.00652f
C16220 XThR.Tn[6].n26 VGND 0.11444f
C16221 XThR.Tn[6].t35 VGND 0.01825f
C16222 XThR.Tn[6].t31 VGND 0.01998f
C16223 XThR.Tn[6].n27 VGND 0.04879f
C16224 XThR.Tn[6].t59 VGND 0.01819f
C16225 XThR.Tn[6].t27 VGND 0.01991f
C16226 XThR.Tn[6].n28 VGND 0.05076f
C16227 XThR.Tn[6].n29 VGND 0.03566f
C16228 XThR.Tn[6].n30 VGND 0.00652f
C16229 XThR.Tn[6].n31 VGND 0.11444f
C16230 XThR.Tn[6].t13 VGND 0.01825f
C16231 XThR.Tn[6].t67 VGND 0.01998f
C16232 XThR.Tn[6].n32 VGND 0.04879f
C16233 XThR.Tn[6].t29 VGND 0.01819f
C16234 XThR.Tn[6].t64 VGND 0.01991f
C16235 XThR.Tn[6].n33 VGND 0.05076f
C16236 XThR.Tn[6].n34 VGND 0.03566f
C16237 XThR.Tn[6].n35 VGND 0.00652f
C16238 XThR.Tn[6].n36 VGND 0.11444f
C16239 XThR.Tn[6].t51 VGND 0.01825f
C16240 XThR.Tn[6].t22 VGND 0.01998f
C16241 XThR.Tn[6].n37 VGND 0.04879f
C16242 XThR.Tn[6].t70 VGND 0.01819f
C16243 XThR.Tn[6].t19 VGND 0.01991f
C16244 XThR.Tn[6].n38 VGND 0.05076f
C16245 XThR.Tn[6].n39 VGND 0.03566f
C16246 XThR.Tn[6].n40 VGND 0.00652f
C16247 XThR.Tn[6].n41 VGND 0.11444f
C16248 XThR.Tn[6].t21 VGND 0.01825f
C16249 XThR.Tn[6].t17 VGND 0.01998f
C16250 XThR.Tn[6].n42 VGND 0.04879f
C16251 XThR.Tn[6].t37 VGND 0.01819f
C16252 XThR.Tn[6].t12 VGND 0.01991f
C16253 XThR.Tn[6].n43 VGND 0.05076f
C16254 XThR.Tn[6].n44 VGND 0.03566f
C16255 XThR.Tn[6].n45 VGND 0.00652f
C16256 XThR.Tn[6].n46 VGND 0.11444f
C16257 XThR.Tn[6].t24 VGND 0.01825f
C16258 XThR.Tn[6].t30 VGND 0.01998f
C16259 XThR.Tn[6].n47 VGND 0.04879f
C16260 XThR.Tn[6].t43 VGND 0.01819f
C16261 XThR.Tn[6].t25 VGND 0.01991f
C16262 XThR.Tn[6].n48 VGND 0.05076f
C16263 XThR.Tn[6].n49 VGND 0.03566f
C16264 XThR.Tn[6].n50 VGND 0.00652f
C16265 XThR.Tn[6].n51 VGND 0.11444f
C16266 XThR.Tn[6].t40 VGND 0.01825f
C16267 XThR.Tn[6].t50 VGND 0.01998f
C16268 XThR.Tn[6].n52 VGND 0.04879f
C16269 XThR.Tn[6].t61 VGND 0.01819f
C16270 XThR.Tn[6].t47 VGND 0.01991f
C16271 XThR.Tn[6].n53 VGND 0.05076f
C16272 XThR.Tn[6].n54 VGND 0.03566f
C16273 XThR.Tn[6].n55 VGND 0.00652f
C16274 XThR.Tn[6].n56 VGND 0.11444f
C16275 XThR.Tn[6].t33 VGND 0.01825f
C16276 XThR.Tn[6].t69 VGND 0.01998f
C16277 XThR.Tn[6].n57 VGND 0.04879f
C16278 XThR.Tn[6].t54 VGND 0.01819f
C16279 XThR.Tn[6].t65 VGND 0.01991f
C16280 XThR.Tn[6].n58 VGND 0.05076f
C16281 XThR.Tn[6].n59 VGND 0.03566f
C16282 XThR.Tn[6].n60 VGND 0.00652f
C16283 XThR.Tn[6].n61 VGND 0.11444f
C16284 XThR.Tn[6].t53 VGND 0.01825f
C16285 XThR.Tn[6].t44 VGND 0.01998f
C16286 XThR.Tn[6].n62 VGND 0.04879f
C16287 XThR.Tn[6].t71 VGND 0.01819f
C16288 XThR.Tn[6].t39 VGND 0.01991f
C16289 XThR.Tn[6].n63 VGND 0.05076f
C16290 XThR.Tn[6].n64 VGND 0.03566f
C16291 XThR.Tn[6].n65 VGND 0.00652f
C16292 XThR.Tn[6].n66 VGND 0.11444f
C16293 XThR.Tn[6].t23 VGND 0.01825f
C16294 XThR.Tn[6].t18 VGND 0.01998f
C16295 XThR.Tn[6].n67 VGND 0.04879f
C16296 XThR.Tn[6].t41 VGND 0.01819f
C16297 XThR.Tn[6].t15 VGND 0.01991f
C16298 XThR.Tn[6].n68 VGND 0.05076f
C16299 XThR.Tn[6].n69 VGND 0.03566f
C16300 XThR.Tn[6].n70 VGND 0.00652f
C16301 XThR.Tn[6].n71 VGND 0.11444f
C16302 XThR.Tn[6].t38 VGND 0.01825f
C16303 XThR.Tn[6].t32 VGND 0.01998f
C16304 XThR.Tn[6].n72 VGND 0.04879f
C16305 XThR.Tn[6].t60 VGND 0.01819f
C16306 XThR.Tn[6].t28 VGND 0.01991f
C16307 XThR.Tn[6].n73 VGND 0.05076f
C16308 XThR.Tn[6].n74 VGND 0.03566f
C16309 XThR.Tn[6].n75 VGND 0.00652f
C16310 XThR.Tn[6].n76 VGND 0.11444f
C16311 XThR.Tn[6].t58 VGND 0.01825f
C16312 XThR.Tn[6].t52 VGND 0.01998f
C16313 XThR.Tn[6].n77 VGND 0.04879f
C16314 XThR.Tn[6].t16 VGND 0.01819f
C16315 XThR.Tn[6].t48 VGND 0.01991f
C16316 XThR.Tn[6].n78 VGND 0.05076f
C16317 XThR.Tn[6].n79 VGND 0.03566f
C16318 XThR.Tn[6].n80 VGND 0.00652f
C16319 XThR.Tn[6].n81 VGND 0.11444f
C16320 XThR.Tn[6].t34 VGND 0.01825f
C16321 XThR.Tn[6].t46 VGND 0.01998f
C16322 XThR.Tn[6].n82 VGND 0.04879f
C16323 XThR.Tn[6].t55 VGND 0.01819f
C16324 XThR.Tn[6].t42 VGND 0.01991f
C16325 XThR.Tn[6].n83 VGND 0.05076f
C16326 XThR.Tn[6].n84 VGND 0.03566f
C16327 XThR.Tn[6].n85 VGND 0.00652f
C16328 XThR.Tn[6].n86 VGND 0.11444f
C16329 XThR.Tn[6].n87 VGND 0.104f
C16330 XThR.Tn[6].n88 VGND 0.17311f
C16331 XThC.Tn[10].t2 VGND 0.01306f
C16332 XThC.Tn[10].t8 VGND 0.01306f
C16333 XThC.Tn[10].n0 VGND 0.03258f
C16334 XThC.Tn[10].t10 VGND 0.01306f
C16335 XThC.Tn[10].t3 VGND 0.01306f
C16336 XThC.Tn[10].n1 VGND 0.02613f
C16337 XThC.Tn[10].n2 VGND 0.06572f
C16338 XThC.Tn[10].n3 VGND 0.02851f
C16339 XThC.Tn[10].t38 VGND 0.01593f
C16340 XThC.Tn[10].t36 VGND 0.0174f
C16341 XThC.Tn[10].n4 VGND 0.03884f
C16342 XThC.Tn[10].n5 VGND 0.02661f
C16343 XThC.Tn[10].n6 VGND 0.08734f
C16344 XThC.Tn[10].t24 VGND 0.01593f
C16345 XThC.Tn[10].t21 VGND 0.0174f
C16346 XThC.Tn[10].n7 VGND 0.03884f
C16347 XThC.Tn[10].n8 VGND 0.02661f
C16348 XThC.Tn[10].n9 VGND 0.08758f
C16349 XThC.Tn[10].n10 VGND 0.14434f
C16350 XThC.Tn[10].t29 VGND 0.01593f
C16351 XThC.Tn[10].t23 VGND 0.0174f
C16352 XThC.Tn[10].n11 VGND 0.03884f
C16353 XThC.Tn[10].n12 VGND 0.02661f
C16354 XThC.Tn[10].n13 VGND 0.08758f
C16355 XThC.Tn[10].n14 VGND 0.14434f
C16356 XThC.Tn[10].t30 VGND 0.01593f
C16357 XThC.Tn[10].t25 VGND 0.0174f
C16358 XThC.Tn[10].n15 VGND 0.03884f
C16359 XThC.Tn[10].n16 VGND 0.02661f
C16360 XThC.Tn[10].n17 VGND 0.08758f
C16361 XThC.Tn[10].n18 VGND 0.14434f
C16362 XThC.Tn[10].t17 VGND 0.01593f
C16363 XThC.Tn[10].t14 VGND 0.0174f
C16364 XThC.Tn[10].n19 VGND 0.03884f
C16365 XThC.Tn[10].n20 VGND 0.02661f
C16366 XThC.Tn[10].n21 VGND 0.08758f
C16367 XThC.Tn[10].n22 VGND 0.14434f
C16368 XThC.Tn[10].t18 VGND 0.01593f
C16369 XThC.Tn[10].t15 VGND 0.0174f
C16370 XThC.Tn[10].n23 VGND 0.03884f
C16371 XThC.Tn[10].n24 VGND 0.02661f
C16372 XThC.Tn[10].n25 VGND 0.08758f
C16373 XThC.Tn[10].n26 VGND 0.14434f
C16374 XThC.Tn[10].t34 VGND 0.01593f
C16375 XThC.Tn[10].t28 VGND 0.0174f
C16376 XThC.Tn[10].n27 VGND 0.03884f
C16377 XThC.Tn[10].n28 VGND 0.02661f
C16378 XThC.Tn[10].n29 VGND 0.08758f
C16379 XThC.Tn[10].n30 VGND 0.14434f
C16380 XThC.Tn[10].t41 VGND 0.01593f
C16381 XThC.Tn[10].t37 VGND 0.0174f
C16382 XThC.Tn[10].n31 VGND 0.03884f
C16383 XThC.Tn[10].n32 VGND 0.02661f
C16384 XThC.Tn[10].n33 VGND 0.08758f
C16385 XThC.Tn[10].n34 VGND 0.14434f
C16386 XThC.Tn[10].t43 VGND 0.01593f
C16387 XThC.Tn[10].t39 VGND 0.0174f
C16388 XThC.Tn[10].n35 VGND 0.03884f
C16389 XThC.Tn[10].n36 VGND 0.02661f
C16390 XThC.Tn[10].n37 VGND 0.08758f
C16391 XThC.Tn[10].n38 VGND 0.14434f
C16392 XThC.Tn[10].t31 VGND 0.01593f
C16393 XThC.Tn[10].t26 VGND 0.0174f
C16394 XThC.Tn[10].n39 VGND 0.03884f
C16395 XThC.Tn[10].n40 VGND 0.02661f
C16396 XThC.Tn[10].n41 VGND 0.08758f
C16397 XThC.Tn[10].n42 VGND 0.14434f
C16398 XThC.Tn[10].t33 VGND 0.01593f
C16399 XThC.Tn[10].t27 VGND 0.0174f
C16400 XThC.Tn[10].n43 VGND 0.03884f
C16401 XThC.Tn[10].n44 VGND 0.02661f
C16402 XThC.Tn[10].n45 VGND 0.08758f
C16403 XThC.Tn[10].n46 VGND 0.14434f
C16404 XThC.Tn[10].t12 VGND 0.01593f
C16405 XThC.Tn[10].t40 VGND 0.0174f
C16406 XThC.Tn[10].n47 VGND 0.03884f
C16407 XThC.Tn[10].n48 VGND 0.02661f
C16408 XThC.Tn[10].n49 VGND 0.08758f
C16409 XThC.Tn[10].n50 VGND 0.14434f
C16410 XThC.Tn[10].t20 VGND 0.01593f
C16411 XThC.Tn[10].t16 VGND 0.0174f
C16412 XThC.Tn[10].n51 VGND 0.03884f
C16413 XThC.Tn[10].n52 VGND 0.02661f
C16414 XThC.Tn[10].n53 VGND 0.08758f
C16415 XThC.Tn[10].n54 VGND 0.14434f
C16416 XThC.Tn[10].t22 VGND 0.01593f
C16417 XThC.Tn[10].t19 VGND 0.0174f
C16418 XThC.Tn[10].n55 VGND 0.03884f
C16419 XThC.Tn[10].n56 VGND 0.02661f
C16420 XThC.Tn[10].n57 VGND 0.08758f
C16421 XThC.Tn[10].n58 VGND 0.14434f
C16422 XThC.Tn[10].t35 VGND 0.01593f
C16423 XThC.Tn[10].t32 VGND 0.0174f
C16424 XThC.Tn[10].n59 VGND 0.03884f
C16425 XThC.Tn[10].n60 VGND 0.02661f
C16426 XThC.Tn[10].n61 VGND 0.08758f
C16427 XThC.Tn[10].n62 VGND 0.14434f
C16428 XThC.Tn[10].t13 VGND 0.01593f
C16429 XThC.Tn[10].t42 VGND 0.0174f
C16430 XThC.Tn[10].n63 VGND 0.03884f
C16431 XThC.Tn[10].n64 VGND 0.02661f
C16432 XThC.Tn[10].n65 VGND 0.08758f
C16433 XThC.Tn[10].n66 VGND 0.14434f
C16434 XThC.Tn[10].n67 VGND 0.61921f
C16435 XThC.Tn[10].n68 VGND 0.2357f
C16436 XThC.Tn[10].t5 VGND 0.0201f
C16437 XThC.Tn[10].t4 VGND 0.0201f
C16438 XThC.Tn[10].n69 VGND 0.04342f
C16439 XThC.Tn[10].t9 VGND 0.0201f
C16440 XThC.Tn[10].t1 VGND 0.0201f
C16441 XThC.Tn[10].n70 VGND 0.06609f
C16442 XThC.Tn[10].n71 VGND 0.18363f
C16443 XThC.Tn[10].n72 VGND 0.02887f
C16444 XThC.Tn[10].t7 VGND 0.0201f
C16445 XThC.Tn[10].t6 VGND 0.0201f
C16446 XThC.Tn[10].n73 VGND 0.04468f
C16447 XThC.Tn[10].t11 VGND 0.0201f
C16448 XThC.Tn[10].t0 VGND 0.0201f
C16449 XThC.Tn[10].n74 VGND 0.06102f
C16450 XThC.Tn[10].n75 VGND 0.19884f
C16451 VPWR.n0 VGND 0.0471f
C16452 VPWR.t989 VGND 0.29789f
C16453 VPWR.t105 VGND 0.13182f
C16454 VPWR.t1694 VGND 0.38006f
C16455 VPWR.t37 VGND 0.14381f
C16456 VPWR.t1890 VGND 0.14381f
C16457 VPWR.t368 VGND 0.14381f
C16458 VPWR.t720 VGND 0.14381f
C16459 VPWR.t716 VGND 0.14381f
C16460 VPWR.t712 VGND 0.14381f
C16461 VPWR.t439 VGND 0.10101f
C16462 VPWR.n1 VGND 0.18352f
C16463 VPWR.n2 VGND 0.0971f
C16464 VPWR.t106 VGND 0.05745f
C16465 VPWR.n3 VGND 0.00925f
C16466 VPWR.t440 VGND 0.0144f
C16467 VPWR.t713 VGND 0.0144f
C16468 VPWR.n4 VGND 0.03162f
C16469 VPWR.t717 VGND 0.0144f
C16470 VPWR.t721 VGND 0.0144f
C16471 VPWR.n5 VGND 0.03156f
C16472 VPWR.n6 VGND 0.06483f
C16473 VPWR.n7 VGND 0.18274f
C16474 VPWR.n8 VGND 0.05786f
C16475 VPWR.n9 VGND 0.0425f
C16476 VPWR.n10 VGND 0.07617f
C16477 VPWR.n11 VGND 0.01124f
C16478 VPWR.n12 VGND 0.01638f
C16479 VPWR.n13 VGND 0.0192f
C16480 VPWR.n14 VGND 0.02816f
C16481 VPWR.n15 VGND 0.08524f
C16482 VPWR.n16 VGND 0.01215f
C16483 VPWR.t990 VGND 0.05743f
C16484 VPWR.n17 VGND 0.07387f
C16485 VPWR.n18 VGND 0.33732f
C16486 VPWR.n19 VGND 0.98363f
C16487 VPWR.n20 VGND 0.32018f
C16488 VPWR.n21 VGND 1.02091f
C16489 VPWR.n22 VGND 0.13957f
C16490 VPWR.t1970 VGND 0.01125f
C16491 VPWR.t1375 VGND 0.01232f
C16492 VPWR.n23 VGND 0.03009f
C16493 VPWR.n24 VGND 0.07993f
C16494 VPWR.t2021 VGND 0.01125f
C16495 VPWR.t1264 VGND 0.01232f
C16496 VPWR.n25 VGND 0.03009f
C16497 VPWR.n26 VGND 0.16087f
C16498 VPWR.t1956 VGND 0.01125f
C16499 VPWR.t1412 VGND 0.01232f
C16500 VPWR.n27 VGND 0.03009f
C16501 VPWR.n28 VGND 0.12818f
C16502 VPWR.t1995 VGND 0.01125f
C16503 VPWR.t1304 VGND 0.01232f
C16504 VPWR.n29 VGND 0.03009f
C16505 VPWR.n30 VGND 0.12818f
C16506 VPWR.t2064 VGND 0.01125f
C16507 VPWR.t1120 VGND 0.01232f
C16508 VPWR.n31 VGND 0.03009f
C16509 VPWR.n32 VGND 0.12818f
C16510 VPWR.t1997 VGND 0.01125f
C16511 VPWR.t1297 VGND 0.01232f
C16512 VPWR.n33 VGND 0.03009f
C16513 VPWR.n34 VGND 0.12818f
C16514 VPWR.t1943 VGND 0.01125f
C16515 VPWR.t1192 VGND 0.01232f
C16516 VPWR.n35 VGND 0.03009f
C16517 VPWR.n36 VGND 0.12818f
C16518 VPWR.t2022 VGND 0.01125f
C16519 VPWR.t1232 VGND 0.01232f
C16520 VPWR.n37 VGND 0.03009f
C16521 VPWR.n38 VGND 0.12818f
C16522 VPWR.t2028 VGND 0.01125f
C16523 VPWR.t1125 VGND 0.01232f
C16524 VPWR.n39 VGND 0.03009f
C16525 VPWR.n40 VGND 0.12818f
C16526 VPWR.t2069 VGND 0.01125f
C16527 VPWR.t1399 VGND 0.01232f
C16528 VPWR.n41 VGND 0.03009f
C16529 VPWR.n42 VGND 0.12818f
C16530 VPWR.t2051 VGND 0.01125f
C16531 VPWR.t1291 VGND 0.01232f
C16532 VPWR.n43 VGND 0.03009f
C16533 VPWR.n44 VGND 0.12818f
C16534 VPWR.t1946 VGND 0.01125f
C16535 VPWR.t1442 VGND 0.01232f
C16536 VPWR.n45 VGND 0.03009f
C16537 VPWR.n46 VGND 0.12818f
C16538 VPWR.t2026 VGND 0.01125f
C16539 VPWR.t1224 VGND 0.01232f
C16540 VPWR.n47 VGND 0.03009f
C16541 VPWR.n48 VGND 0.12818f
C16542 VPWR.t2066 VGND 0.01125f
C16543 VPWR.t1112 VGND 0.01232f
C16544 VPWR.n49 VGND 0.03009f
C16545 VPWR.n50 VGND 0.12818f
C16546 VPWR.t1963 VGND 0.01125f
C16547 VPWR.t1394 VGND 0.01232f
C16548 VPWR.n51 VGND 0.03009f
C16549 VPWR.n52 VGND 0.12818f
C16550 VPWR.t2053 VGND 0.01125f
C16551 VPWR.t1434 VGND 0.01232f
C16552 VPWR.n53 VGND 0.03009f
C16553 VPWR.n54 VGND 0.13878f
C16554 VPWR.n55 VGND 0.11587f
C16555 VPWR.t1223 VGND 0.03348f
C16556 VPWR.t1328 VGND 0.02976f
C16557 VPWR.n56 VGND 0.09198f
C16558 VPWR.t1091 VGND 0.09265f
C16559 VPWR.t1098 VGND 0.03348f
C16560 VPWR.t1092 VGND 0.02976f
C16561 VPWR.n57 VGND 0.09198f
C16562 VPWR.n58 VGND 0.03454f
C16563 VPWR.n59 VGND 0.13984f
C16564 VPWR.n60 VGND 0.13984f
C16565 VPWR.n61 VGND 0.03454f
C16566 VPWR.t1079 VGND 0.03348f
C16567 VPWR.t1452 VGND 0.02976f
C16568 VPWR.n62 VGND 0.09198f
C16569 VPWR.t1318 VGND 0.09265f
C16570 VPWR.t1229 VGND 0.03348f
C16571 VPWR.t1319 VGND 0.02976f
C16572 VPWR.n63 VGND 0.09198f
C16573 VPWR.n64 VGND 0.03454f
C16574 VPWR.n65 VGND 0.13984f
C16575 VPWR.n66 VGND 0.13984f
C16576 VPWR.n67 VGND 0.03454f
C16577 VPWR.t1199 VGND 0.03348f
C16578 VPWR.t1191 VGND 0.02976f
C16579 VPWR.n68 VGND 0.09198f
C16580 VPWR.t1172 VGND 0.09265f
C16581 VPWR.t1455 VGND 0.03348f
C16582 VPWR.t1173 VGND 0.02976f
C16583 VPWR.n69 VGND 0.09198f
C16584 VPWR.n70 VGND 0.03454f
C16585 VPWR.n71 VGND 0.13984f
C16586 VPWR.n72 VGND 0.13984f
C16587 VPWR.n73 VGND 0.03454f
C16588 VPWR.t1325 VGND 0.03348f
C16589 VPWR.t1406 VGND 0.02976f
C16590 VPWR.n74 VGND 0.09198f
C16591 VPWR.t1295 VGND 0.09265f
C16592 VPWR.t1309 VGND 0.03348f
C16593 VPWR.t1296 VGND 0.02976f
C16594 VPWR.n75 VGND 0.09198f
C16595 VPWR.n76 VGND 0.03454f
C16596 VPWR.n77 VGND 0.13984f
C16597 VPWR.n78 VGND 0.13984f
C16598 VPWR.n79 VGND 0.03454f
C16599 VPWR.t1149 VGND 0.03348f
C16600 VPWR.t1168 VGND 0.02976f
C16601 VPWR.n80 VGND 0.09198f
C16602 VPWR.t1132 VGND 0.09265f
C16603 VPWR.t1428 VGND 0.03348f
C16604 VPWR.t1133 VGND 0.02976f
C16605 VPWR.n81 VGND 0.09198f
C16606 VPWR.n82 VGND 0.03454f
C16607 VPWR.n83 VGND 0.13984f
C16608 VPWR.n84 VGND 0.13984f
C16609 VPWR.n85 VGND 0.03454f
C16610 VPWR.t1272 VGND 0.03348f
C16611 VPWR.t1409 VGND 0.02976f
C16612 VPWR.n86 VGND 0.09198f
C16613 VPWR.t1253 VGND 0.09265f
C16614 VPWR.t1260 VGND 0.03348f
C16615 VPWR.t1254 VGND 0.02976f
C16616 VPWR.n87 VGND 0.09198f
C16617 VPWR.n88 VGND 0.03454f
C16618 VPWR.n89 VGND 0.13984f
C16619 VPWR.n90 VGND 0.13984f
C16620 VPWR.n91 VGND 0.03454f
C16621 VPWR.t1152 VGND 0.03348f
C16622 VPWR.t1146 VGND 0.02976f
C16623 VPWR.n92 VGND 0.09198f
C16624 VPWR.t1383 VGND 0.09265f
C16625 VPWR.t1387 VGND 0.03348f
C16626 VPWR.t1384 VGND 0.02976f
C16627 VPWR.n93 VGND 0.09198f
C16628 VPWR.n94 VGND 0.03454f
C16629 VPWR.n95 VGND 0.13984f
C16630 VPWR.n96 VGND 0.13984f
C16631 VPWR.n97 VGND 0.03454f
C16632 VPWR.t1275 VGND 0.03348f
C16633 VPWR.t1366 VGND 0.02976f
C16634 VPWR.n98 VGND 0.09198f
C16635 VPWR.t1129 VGND 0.14585f
C16636 VPWR.t1105 VGND 0.07889f
C16637 VPWR.t1236 VGND 0.09265f
C16638 VPWR.t1130 VGND 0.03348f
C16639 VPWR.t1237 VGND 0.02976f
C16640 VPWR.n99 VGND 0.09198f
C16641 VPWR.t1987 VGND 0.01125f
C16642 VPWR.t1364 VGND 0.01232f
C16643 VPWR.n100 VGND 0.03008f
C16644 VPWR.n101 VGND 0.03301f
C16645 VPWR.n102 VGND 0.00701f
C16646 VPWR.n103 VGND 0.01831f
C16647 VPWR.t2032 VGND 0.01125f
C16648 VPWR.t1235 VGND 0.01232f
C16649 VPWR.n104 VGND 0.03008f
C16650 VPWR.n105 VGND 0.03301f
C16651 VPWR.t1981 VGND 0.01122f
C16652 VPWR.t1128 VGND 0.01228f
C16653 VPWR.n106 VGND 0.03131f
C16654 VPWR.n107 VGND 0.01979f
C16655 VPWR.t1934 VGND 0.01141f
C16656 VPWR.t1104 VGND 0.01247f
C16657 VPWR.n108 VGND 0.02782f
C16658 VPWR.n109 VGND 0.02832f
C16659 VPWR.n110 VGND 0.01785f
C16660 VPWR.n111 VGND 0.00701f
C16661 VPWR.n112 VGND 0.01831f
C16662 VPWR.n113 VGND 0.02668f
C16663 VPWR.t2001 VGND 0.01125f
C16664 VPWR.t1326 VGND 0.01232f
C16665 VPWR.n114 VGND 0.03008f
C16666 VPWR.n115 VGND 0.03301f
C16667 VPWR.t1951 VGND 0.01122f
C16668 VPWR.t1221 VGND 0.01228f
C16669 VPWR.n116 VGND 0.03131f
C16670 VPWR.n117 VGND 0.03712f
C16671 VPWR.n118 VGND 0.00837f
C16672 VPWR.t2048 VGND 0.01141f
C16673 VPWR.t1205 VGND 0.01247f
C16674 VPWR.n119 VGND 0.02782f
C16675 VPWR.n120 VGND 0.02832f
C16676 VPWR.n121 VGND 0.01785f
C16677 VPWR.n122 VGND 0.00701f
C16678 VPWR.n123 VGND 0.01831f
C16679 VPWR.n124 VGND 0.02554f
C16680 VPWR.t1940 VGND 0.01125f
C16681 VPWR.t1090 VGND 0.01232f
C16682 VPWR.n125 VGND 0.03008f
C16683 VPWR.n126 VGND 0.03301f
C16684 VPWR.t1991 VGND 0.01122f
C16685 VPWR.t1096 VGND 0.01228f
C16686 VPWR.n127 VGND 0.03131f
C16687 VPWR.n128 VGND 0.03712f
C16688 VPWR.n129 VGND 0.00837f
C16689 VPWR.t1990 VGND 0.01141f
C16690 VPWR.t1354 VGND 0.01247f
C16691 VPWR.n130 VGND 0.02782f
C16692 VPWR.n131 VGND 0.02832f
C16693 VPWR.n132 VGND 0.01785f
C16694 VPWR.n133 VGND 0.00701f
C16695 VPWR.n134 VGND 0.01831f
C16696 VPWR.n135 VGND 0.02396f
C16697 VPWR.n136 VGND 0.2127f
C16698 VPWR.t1954 VGND 0.01125f
C16699 VPWR.t1450 VGND 0.01232f
C16700 VPWR.n137 VGND 0.03008f
C16701 VPWR.n138 VGND 0.03301f
C16702 VPWR.t2046 VGND 0.01122f
C16703 VPWR.t1077 VGND 0.01228f
C16704 VPWR.n139 VGND 0.03131f
C16705 VPWR.n140 VGND 0.03712f
C16706 VPWR.n141 VGND 0.00837f
C16707 VPWR.t1999 VGND 0.01141f
C16708 VPWR.t1329 VGND 0.01247f
C16709 VPWR.n142 VGND 0.02782f
C16710 VPWR.n143 VGND 0.02832f
C16711 VPWR.n144 VGND 0.01785f
C16712 VPWR.n145 VGND 0.00701f
C16713 VPWR.n146 VGND 0.01831f
C16714 VPWR.n147 VGND 0.02396f
C16715 VPWR.n148 VGND 0.17674f
C16716 VPWR.t2004 VGND 0.01125f
C16717 VPWR.t1317 VGND 0.01232f
C16718 VPWR.n149 VGND 0.03008f
C16719 VPWR.n150 VGND 0.03301f
C16720 VPWR.t1942 VGND 0.01122f
C16721 VPWR.t1227 VGND 0.01228f
C16722 VPWR.n151 VGND 0.03131f
C16723 VPWR.n152 VGND 0.03712f
C16724 VPWR.n153 VGND 0.00837f
C16725 VPWR.t2007 VGND 0.01141f
C16726 VPWR.t1310 VGND 0.01247f
C16727 VPWR.n154 VGND 0.02782f
C16728 VPWR.n155 VGND 0.02832f
C16729 VPWR.n156 VGND 0.01785f
C16730 VPWR.n157 VGND 0.00701f
C16731 VPWR.n158 VGND 0.01831f
C16732 VPWR.n159 VGND 0.02396f
C16733 VPWR.n160 VGND 0.17674f
C16734 VPWR.t2052 VGND 0.01125f
C16735 VPWR.t1189 VGND 0.01232f
C16736 VPWR.n161 VGND 0.03008f
C16737 VPWR.n162 VGND 0.03301f
C16738 VPWR.t1998 VGND 0.01122f
C16739 VPWR.t1197 VGND 0.01228f
C16740 VPWR.n163 VGND 0.03131f
C16741 VPWR.n164 VGND 0.03712f
C16742 VPWR.n165 VGND 0.00837f
C16743 VPWR.t1952 VGND 0.01141f
C16744 VPWR.t1456 VGND 0.01247f
C16745 VPWR.n166 VGND 0.02782f
C16746 VPWR.n167 VGND 0.02832f
C16747 VPWR.n168 VGND 0.01785f
C16748 VPWR.n169 VGND 0.00701f
C16749 VPWR.n170 VGND 0.01831f
C16750 VPWR.n171 VGND 0.02396f
C16751 VPWR.n172 VGND 0.17674f
C16752 VPWR.t2058 VGND 0.01125f
C16753 VPWR.t1171 VGND 0.01232f
C16754 VPWR.n173 VGND 0.03008f
C16755 VPWR.n174 VGND 0.03301f
C16756 VPWR.t2006 VGND 0.01122f
C16757 VPWR.t1453 VGND 0.01228f
C16758 VPWR.n175 VGND 0.03131f
C16759 VPWR.n176 VGND 0.03712f
C16760 VPWR.n177 VGND 0.00837f
C16761 VPWR.t1961 VGND 0.01141f
C16762 VPWR.t1437 VGND 0.01247f
C16763 VPWR.n178 VGND 0.02782f
C16764 VPWR.n179 VGND 0.02832f
C16765 VPWR.n180 VGND 0.01785f
C16766 VPWR.n181 VGND 0.00701f
C16767 VPWR.n182 VGND 0.01831f
C16768 VPWR.n183 VGND 0.02396f
C16769 VPWR.n184 VGND 0.17674f
C16770 VPWR.t1973 VGND 0.01125f
C16771 VPWR.t1404 VGND 0.01232f
C16772 VPWR.n185 VGND 0.03008f
C16773 VPWR.n186 VGND 0.03301f
C16774 VPWR.t2054 VGND 0.01122f
C16775 VPWR.t1323 VGND 0.01228f
C16776 VPWR.n187 VGND 0.03131f
C16777 VPWR.n188 VGND 0.03712f
C16778 VPWR.n189 VGND 0.00837f
C16779 VPWR.t2017 VGND 0.01141f
C16780 VPWR.t1276 VGND 0.01247f
C16781 VPWR.n190 VGND 0.02782f
C16782 VPWR.n191 VGND 0.02832f
C16783 VPWR.n192 VGND 0.01785f
C16784 VPWR.n193 VGND 0.00701f
C16785 VPWR.n194 VGND 0.01831f
C16786 VPWR.n195 VGND 0.02396f
C16787 VPWR.n196 VGND 0.17674f
C16788 VPWR.t2009 VGND 0.01125f
C16789 VPWR.t1294 VGND 0.01232f
C16790 VPWR.n197 VGND 0.03008f
C16791 VPWR.n198 VGND 0.03301f
C16792 VPWR.t1960 VGND 0.01122f
C16793 VPWR.t1307 VGND 0.01228f
C16794 VPWR.n199 VGND 0.03131f
C16795 VPWR.n200 VGND 0.03712f
C16796 VPWR.n201 VGND 0.00837f
C16797 VPWR.t2057 VGND 0.01141f
C16798 VPWR.t1174 VGND 0.01247f
C16799 VPWR.n202 VGND 0.02782f
C16800 VPWR.n203 VGND 0.02832f
C16801 VPWR.n204 VGND 0.01785f
C16802 VPWR.n205 VGND 0.00701f
C16803 VPWR.n206 VGND 0.01831f
C16804 VPWR.n207 VGND 0.02396f
C16805 VPWR.n208 VGND 0.17674f
C16806 VPWR.t2060 VGND 0.01125f
C16807 VPWR.t1166 VGND 0.01232f
C16808 VPWR.n209 VGND 0.03008f
C16809 VPWR.n210 VGND 0.03301f
C16810 VPWR.t1974 VGND 0.01122f
C16811 VPWR.t1147 VGND 0.01228f
C16812 VPWR.n211 VGND 0.03131f
C16813 VPWR.n212 VGND 0.03712f
C16814 VPWR.n213 VGND 0.00837f
C16815 VPWR.t1928 VGND 0.01141f
C16816 VPWR.t1139 VGND 0.01247f
C16817 VPWR.n214 VGND 0.02782f
C16818 VPWR.n215 VGND 0.02832f
C16819 VPWR.n216 VGND 0.01785f
C16820 VPWR.n217 VGND 0.00701f
C16821 VPWR.n218 VGND 0.01831f
C16822 VPWR.n219 VGND 0.02396f
C16823 VPWR.n220 VGND 0.17674f
C16824 VPWR.t1931 VGND 0.01125f
C16825 VPWR.t1131 VGND 0.01232f
C16826 VPWR.n221 VGND 0.03008f
C16827 VPWR.n222 VGND 0.03301f
C16828 VPWR.t2056 VGND 0.01122f
C16829 VPWR.t1426 VGND 0.01228f
C16830 VPWR.n223 VGND 0.03131f
C16831 VPWR.n224 VGND 0.03712f
C16832 VPWR.n225 VGND 0.00837f
C16833 VPWR.t2008 VGND 0.01141f
C16834 VPWR.t1302 VGND 0.01247f
C16835 VPWR.n226 VGND 0.02782f
C16836 VPWR.n227 VGND 0.02832f
C16837 VPWR.n228 VGND 0.01785f
C16838 VPWR.n229 VGND 0.00701f
C16839 VPWR.n230 VGND 0.01831f
C16840 VPWR.n231 VGND 0.02396f
C16841 VPWR.n232 VGND 0.17674f
C16842 VPWR.t1972 VGND 0.01125f
C16843 VPWR.t1407 VGND 0.01232f
C16844 VPWR.n233 VGND 0.03008f
C16845 VPWR.n234 VGND 0.03301f
C16846 VPWR.t1926 VGND 0.01122f
C16847 VPWR.t1270 VGND 0.01228f
C16848 VPWR.n235 VGND 0.03131f
C16849 VPWR.n236 VGND 0.03712f
C16850 VPWR.n237 VGND 0.00837f
C16851 VPWR.t2016 VGND 0.01141f
C16852 VPWR.t1278 VGND 0.01247f
C16853 VPWR.n238 VGND 0.02782f
C16854 VPWR.n239 VGND 0.02832f
C16855 VPWR.n240 VGND 0.01785f
C16856 VPWR.n241 VGND 0.00701f
C16857 VPWR.n242 VGND 0.01831f
C16858 VPWR.n243 VGND 0.02396f
C16859 VPWR.n244 VGND 0.17674f
C16860 VPWR.t2027 VGND 0.01125f
C16861 VPWR.t1252 VGND 0.01232f
C16862 VPWR.n245 VGND 0.03008f
C16863 VPWR.n246 VGND 0.03301f
C16864 VPWR.t1932 VGND 0.01122f
C16865 VPWR.t1258 VGND 0.01228f
C16866 VPWR.n247 VGND 0.03131f
C16867 VPWR.n248 VGND 0.03712f
C16868 VPWR.n249 VGND 0.00837f
C16869 VPWR.t1930 VGND 0.01141f
C16870 VPWR.t1134 VGND 0.01247f
C16871 VPWR.n250 VGND 0.02782f
C16872 VPWR.n251 VGND 0.02832f
C16873 VPWR.n252 VGND 0.01785f
C16874 VPWR.n253 VGND 0.00701f
C16875 VPWR.n254 VGND 0.01831f
C16876 VPWR.n255 VGND 0.02396f
C16877 VPWR.n256 VGND 0.17674f
C16878 VPWR.t2068 VGND 0.01125f
C16879 VPWR.t1144 VGND 0.01232f
C16880 VPWR.n257 VGND 0.03008f
C16881 VPWR.n258 VGND 0.03301f
C16882 VPWR.t2015 VGND 0.01122f
C16883 VPWR.t1150 VGND 0.01228f
C16884 VPWR.n259 VGND 0.03131f
C16885 VPWR.n260 VGND 0.03712f
C16886 VPWR.n261 VGND 0.00837f
C16887 VPWR.t1971 VGND 0.01141f
C16888 VPWR.t1410 VGND 0.01247f
C16889 VPWR.n262 VGND 0.02782f
C16890 VPWR.n263 VGND 0.02832f
C16891 VPWR.n264 VGND 0.01785f
C16892 VPWR.n265 VGND 0.00701f
C16893 VPWR.n266 VGND 0.01831f
C16894 VPWR.n267 VGND 0.02396f
C16895 VPWR.n268 VGND 0.17674f
C16896 VPWR.t1980 VGND 0.01125f
C16897 VPWR.t1382 VGND 0.01232f
C16898 VPWR.n269 VGND 0.03008f
C16899 VPWR.n270 VGND 0.03301f
C16900 VPWR.t2029 VGND 0.01122f
C16901 VPWR.t1385 VGND 0.01228f
C16902 VPWR.n271 VGND 0.03131f
C16903 VPWR.n272 VGND 0.03712f
C16904 VPWR.n273 VGND 0.00837f
C16905 VPWR.t1983 VGND 0.01141f
C16906 VPWR.t1370 VGND 0.01247f
C16907 VPWR.n274 VGND 0.02782f
C16908 VPWR.n275 VGND 0.02832f
C16909 VPWR.n276 VGND 0.01785f
C16910 VPWR.n277 VGND 0.00701f
C16911 VPWR.n278 VGND 0.01831f
C16912 VPWR.n279 VGND 0.02396f
C16913 VPWR.n280 VGND 0.17674f
C16914 VPWR.n281 VGND 0.23844f
C16915 VPWR.n282 VGND 0.02396f
C16916 VPWR.n283 VGND 0.01785f
C16917 VPWR.t2030 VGND 0.01141f
C16918 VPWR.t1240 VGND 0.01247f
C16919 VPWR.n284 VGND 0.02782f
C16920 VPWR.n285 VGND 0.02832f
C16921 VPWR.n286 VGND 0.00837f
C16922 VPWR.t1933 VGND 0.01122f
C16923 VPWR.t1273 VGND 0.01228f
C16924 VPWR.n287 VGND 0.03131f
C16925 VPWR.n288 VGND 0.03712f
C16926 VPWR.n289 VGND 0.03454f
C16927 VPWR.t567 VGND 0.03348f
C16928 VPWR.t1748 VGND 0.02976f
C16929 VPWR.n290 VGND 0.09198f
C16930 VPWR.t566 VGND 0.14585f
C16931 VPWR.t1774 VGND 0.07889f
C16932 VPWR.t1747 VGND 0.09265f
C16933 VPWR.t27 VGND 0.03348f
C16934 VPWR.t1436 VGND 0.02976f
C16935 VPWR.n291 VGND 0.09198f
C16936 VPWR.n292 VGND 0.01806f
C16937 VPWR.n293 VGND 0.07657f
C16938 VPWR.t1435 VGND 0.13401f
C16939 VPWR.t242 VGND 0.07889f
C16940 VPWR.t26 VGND 0.12017f
C16941 VPWR.t355 VGND 0.03348f
C16942 VPWR.t176 VGND 0.02976f
C16943 VPWR.n294 VGND 0.09198f
C16944 VPWR.n295 VGND 0.01806f
C16945 VPWR.n296 VGND 0.00732f
C16946 VPWR.n297 VGND 0.10877f
C16947 VPWR.t175 VGND 0.09265f
C16948 VPWR.t1605 VGND 0.07889f
C16949 VPWR.t354 VGND 0.12017f
C16950 VPWR.t1792 VGND 0.03348f
C16951 VPWR.t1045 VGND 0.02976f
C16952 VPWR.n298 VGND 0.09198f
C16953 VPWR.n299 VGND 0.01806f
C16954 VPWR.n300 VGND 0.00732f
C16955 VPWR.n301 VGND 0.10877f
C16956 VPWR.t1044 VGND 0.09265f
C16957 VPWR.t881 VGND 0.07889f
C16958 VPWR.t1791 VGND 0.12017f
C16959 VPWR.t218 VGND 0.03348f
C16960 VPWR.t876 VGND 0.02976f
C16961 VPWR.n302 VGND 0.09198f
C16962 VPWR.n303 VGND 0.01806f
C16963 VPWR.n304 VGND 0.00732f
C16964 VPWR.n305 VGND 0.10877f
C16965 VPWR.t875 VGND 0.09265f
C16966 VPWR.t882 VGND 0.07889f
C16967 VPWR.t217 VGND 0.12017f
C16968 VPWR.t1000 VGND 0.03348f
C16969 VPWR.t896 VGND 0.02976f
C16970 VPWR.n306 VGND 0.09198f
C16971 VPWR.n307 VGND 0.01806f
C16972 VPWR.n308 VGND 0.00732f
C16973 VPWR.n309 VGND 0.10877f
C16974 VPWR.t895 VGND 0.09265f
C16975 VPWR.t1775 VGND 0.07889f
C16976 VPWR.t999 VGND 0.12017f
C16977 VPWR.t331 VGND 0.03348f
C16978 VPWR.t1625 VGND 0.02976f
C16979 VPWR.n310 VGND 0.09198f
C16980 VPWR.n311 VGND 0.01806f
C16981 VPWR.n312 VGND 0.00732f
C16982 VPWR.n313 VGND 0.10877f
C16983 VPWR.t1624 VGND 0.09265f
C16984 VPWR.t1776 VGND 0.07889f
C16985 VPWR.t330 VGND 0.12017f
C16986 VPWR.t452 VGND 0.03348f
C16987 VPWR.t341 VGND 0.02976f
C16988 VPWR.n314 VGND 0.09198f
C16989 VPWR.n315 VGND 0.01806f
C16990 VPWR.n316 VGND 0.00732f
C16991 VPWR.n317 VGND 0.10877f
C16992 VPWR.t340 VGND 0.09265f
C16993 VPWR.t240 VGND 0.07889f
C16994 VPWR.t451 VGND 0.12017f
C16995 VPWR.t1851 VGND 0.03348f
C16996 VPWR.t658 VGND 0.02976f
C16997 VPWR.n318 VGND 0.09198f
C16998 VPWR.n319 VGND 0.01806f
C16999 VPWR.n320 VGND 0.00732f
C17000 VPWR.n321 VGND 0.10877f
C17001 VPWR.t657 VGND 0.09265f
C17002 VPWR.t243 VGND 0.07889f
C17003 VPWR.t1850 VGND 0.12017f
C17004 VPWR.t198 VGND 0.03348f
C17005 VPWR.t1702 VGND 0.02976f
C17006 VPWR.n322 VGND 0.09198f
C17007 VPWR.n323 VGND 0.01806f
C17008 VPWR.n324 VGND 0.00732f
C17009 VPWR.n325 VGND 0.10877f
C17010 VPWR.t1701 VGND 0.09265f
C17011 VPWR.t244 VGND 0.07889f
C17012 VPWR.t197 VGND 0.12017f
C17013 VPWR.t786 VGND 0.03348f
C17014 VPWR.t270 VGND 0.02976f
C17015 VPWR.n326 VGND 0.09198f
C17016 VPWR.n327 VGND 0.01806f
C17017 VPWR.n328 VGND 0.00732f
C17018 VPWR.n329 VGND 0.10877f
C17019 VPWR.t269 VGND 0.09265f
C17020 VPWR.t883 VGND 0.07889f
C17021 VPWR.t785 VGND 0.12017f
C17022 VPWR.t975 VGND 0.03348f
C17023 VPWR.t792 VGND 0.02976f
C17024 VPWR.n330 VGND 0.09198f
C17025 VPWR.n331 VGND 0.01806f
C17026 VPWR.n332 VGND 0.00732f
C17027 VPWR.n333 VGND 0.10877f
C17028 VPWR.t791 VGND 0.09265f
C17029 VPWR.t239 VGND 0.07889f
C17030 VPWR.t974 VGND 0.12017f
C17031 VPWR.t1722 VGND 0.03348f
C17032 VPWR.t981 VGND 0.02976f
C17033 VPWR.n334 VGND 0.09198f
C17034 VPWR.n335 VGND 0.01806f
C17035 VPWR.n336 VGND 0.00732f
C17036 VPWR.n337 VGND 0.10877f
C17037 VPWR.t980 VGND 0.09265f
C17038 VPWR.t1773 VGND 0.07889f
C17039 VPWR.t1721 VGND 0.12017f
C17040 VPWR.t1494 VGND 0.03348f
C17041 VPWR.t313 VGND 0.02976f
C17042 VPWR.n338 VGND 0.09198f
C17043 VPWR.n339 VGND 0.01806f
C17044 VPWR.n340 VGND 0.00732f
C17045 VPWR.n341 VGND 0.10877f
C17046 VPWR.t312 VGND 0.09265f
C17047 VPWR.t1777 VGND 0.07889f
C17048 VPWR.t1493 VGND 0.12017f
C17049 VPWR.t1670 VGND 0.03348f
C17050 VPWR.t1470 VGND 0.02976f
C17051 VPWR.n342 VGND 0.09198f
C17052 VPWR.n343 VGND 0.01806f
C17053 VPWR.n344 VGND 0.00732f
C17054 VPWR.n345 VGND 0.10877f
C17055 VPWR.t1469 VGND 0.09265f
C17056 VPWR.t1604 VGND 0.07889f
C17057 VPWR.t1669 VGND 0.12017f
C17058 VPWR.t924 VGND 0.03348f
C17059 VPWR.t700 VGND 0.02976f
C17060 VPWR.n346 VGND 0.09198f
C17061 VPWR.n347 VGND 0.01806f
C17062 VPWR.n348 VGND 0.00732f
C17063 VPWR.n349 VGND 0.10877f
C17064 VPWR.t699 VGND 0.09265f
C17065 VPWR.t241 VGND 0.07889f
C17066 VPWR.t923 VGND 0.12017f
C17067 VPWR.n350 VGND 0.10877f
C17068 VPWR.n351 VGND 0.00732f
C17069 VPWR.n352 VGND 0.01806f
C17070 VPWR.n353 VGND 0.13984f
C17071 VPWR.n354 VGND 1.01451f
C17072 VPWR.n355 VGND 0.13984f
C17073 VPWR.t573 VGND 0.03348f
C17074 VPWR.t1563 VGND 0.02976f
C17075 VPWR.n356 VGND 0.09198f
C17076 VPWR.t572 VGND 0.14585f
C17077 VPWR.t931 VGND 0.07889f
C17078 VPWR.t1562 VGND 0.09265f
C17079 VPWR.t703 VGND 0.12017f
C17080 VPWR.t1744 VGND 0.03348f
C17081 VPWR.t708 VGND 0.02976f
C17082 VPWR.n357 VGND 0.09198f
C17083 VPWR.n358 VGND 0.13984f
C17084 VPWR.n359 VGND 0.13984f
C17085 VPWR.t704 VGND 0.03348f
C17086 VPWR.t1462 VGND 0.02976f
C17087 VPWR.n360 VGND 0.09198f
C17088 VPWR.t1673 VGND 0.07889f
C17089 VPWR.t1461 VGND 0.09265f
C17090 VPWR.t1729 VGND 0.12017f
C17091 VPWR.t1486 VGND 0.03348f
C17092 VPWR.t325 VGND 0.02976f
C17093 VPWR.n361 VGND 0.09198f
C17094 VPWR.n362 VGND 0.13984f
C17095 VPWR.n363 VGND 0.13984f
C17096 VPWR.t1730 VGND 0.03348f
C17097 VPWR.t757 VGND 0.02976f
C17098 VPWR.n364 VGND 0.09198f
C17099 VPWR.t930 VGND 0.07889f
C17100 VPWR.t756 VGND 0.09265f
C17101 VPWR.t795 VGND 0.12017f
C17102 VPWR.t751 VGND 0.03348f
C17103 VPWR.t810 VGND 0.02976f
C17104 VPWR.n365 VGND 0.09198f
C17105 VPWR.n366 VGND 0.13984f
C17106 VPWR.n367 VGND 0.13984f
C17107 VPWR.t796 VGND 0.03348f
C17108 VPWR.t280 VGND 0.02976f
C17109 VPWR.n368 VGND 0.09198f
C17110 VPWR.t816 VGND 0.07889f
C17111 VPWR.t279 VGND 0.09265f
C17112 VPWR.t1856 VGND 0.12017f
C17113 VPWR.t274 VGND 0.03348f
C17114 VPWR.t200 VGND 0.02976f
C17115 VPWR.n369 VGND 0.09198f
C17116 VPWR.n370 VGND 0.13984f
C17117 VPWR.n371 VGND 0.13984f
C17118 VPWR.t1857 VGND 0.03348f
C17119 VPWR.t668 VGND 0.02976f
C17120 VPWR.n372 VGND 0.09198f
C17121 VPWR.t346 VGND 0.07889f
C17122 VPWR.t667 VGND 0.09265f
C17123 VPWR.t336 VGND 0.12017f
C17124 VPWR.t662 VGND 0.03348f
C17125 VPWR.t538 VGND 0.02976f
C17126 VPWR.n373 VGND 0.09198f
C17127 VPWR.n374 VGND 0.13984f
C17128 VPWR.n375 VGND 0.13984f
C17129 VPWR.t337 VGND 0.03348f
C17130 VPWR.t769 VGND 0.02976f
C17131 VPWR.n376 VGND 0.09198f
C17132 VPWR.t933 VGND 0.07889f
C17133 VPWR.t768 VGND 0.09265f
C17134 VPWR.t891 VGND 0.12017f
C17135 VPWR.t1629 VGND 0.03348f
C17136 VPWR.t994 VGND 0.02976f
C17137 VPWR.n377 VGND 0.09198f
C17138 VPWR.n378 VGND 0.13984f
C17139 VPWR.n379 VGND 0.13984f
C17140 VPWR.t892 VGND 0.03348f
C17141 VPWR.t93 VGND 0.02976f
C17142 VPWR.n380 VGND 0.09198f
C17143 VPWR.t815 VGND 0.07889f
C17144 VPWR.t92 VGND 0.09265f
C17145 VPWR.t639 VGND 0.12017f
C17146 VPWR.t1798 VGND 0.03348f
C17147 VPWR.t1022 VGND 0.02976f
C17148 VPWR.n381 VGND 0.09198f
C17149 VPWR.n382 VGND 0.13984f
C17150 VPWR.n383 VGND 0.13984f
C17151 VPWR.t640 VGND 0.03348f
C17152 VPWR.t230 VGND 0.02976f
C17153 VPWR.n384 VGND 0.09198f
C17154 VPWR.t1674 VGND 0.07889f
C17155 VPWR.t229 VGND 0.09265f
C17156 VPWR.t168 VGND 0.03348f
C17157 VPWR.t1396 VGND 0.02976f
C17158 VPWR.n385 VGND 0.09198f
C17159 VPWR.t19 VGND 0.03348f
C17160 VPWR.t1114 VGND 0.02976f
C17161 VPWR.n386 VGND 0.09198f
C17162 VPWR.t562 VGND 0.14585f
C17163 VPWR.t606 VGND 0.07889f
C17164 VPWR.t919 VGND 0.09265f
C17165 VPWR.t563 VGND 0.03348f
C17166 VPWR.t920 VGND 0.02976f
C17167 VPWR.n387 VGND 0.09198f
C17168 VPWR.n388 VGND 0.01806f
C17169 VPWR.n389 VGND 0.00732f
C17170 VPWR.n390 VGND 0.10877f
C17171 VPWR.t288 VGND 0.12017f
C17172 VPWR.t941 VGND 0.07889f
C17173 VPWR.t781 VGND 0.09265f
C17174 VPWR.t289 VGND 0.03348f
C17175 VPWR.t782 VGND 0.02976f
C17176 VPWR.n391 VGND 0.09198f
C17177 VPWR.n392 VGND 0.01806f
C17178 VPWR.n393 VGND 0.00732f
C17179 VPWR.n394 VGND 0.10877f
C17180 VPWR.t726 VGND 0.12017f
C17181 VPWR.t686 VGND 0.07889f
C17182 VPWR.t1479 VGND 0.09265f
C17183 VPWR.t727 VGND 0.03348f
C17184 VPWR.t1480 VGND 0.02976f
C17185 VPWR.n395 VGND 0.09198f
C17186 VPWR.n396 VGND 0.01806f
C17187 VPWR.n397 VGND 0.00732f
C17188 VPWR.n398 VGND 0.10877f
C17189 VPWR.t1505 VGND 0.12017f
C17190 VPWR.t685 VGND 0.07889f
C17191 VPWR.t1733 VGND 0.09265f
C17192 VPWR.t1506 VGND 0.03348f
C17193 VPWR.t1734 VGND 0.02976f
C17194 VPWR.n399 VGND 0.09198f
C17195 VPWR.n400 VGND 0.01806f
C17196 VPWR.n401 VGND 0.00732f
C17197 VPWR.n402 VGND 0.10877f
C17198 VPWR.t1576 VGND 0.12017f
C17199 VPWR.t605 VGND 0.07889f
C17200 VPWR.t81 VGND 0.09265f
C17201 VPWR.t1577 VGND 0.03348f
C17202 VPWR.t82 VGND 0.02976f
C17203 VPWR.n403 VGND 0.09198f
C17204 VPWR.n404 VGND 0.01806f
C17205 VPWR.n405 VGND 0.00732f
C17206 VPWR.n406 VGND 0.10877f
C17207 VPWR.t296 VGND 0.12017f
C17208 VPWR.t972 VGND 0.07889f
C17209 VPWR.t803 VGND 0.09265f
C17210 VPWR.t297 VGND 0.03348f
C17211 VPWR.t804 VGND 0.02976f
C17212 VPWR.n407 VGND 0.09198f
C17213 VPWR.n408 VGND 0.01806f
C17214 VPWR.n409 VGND 0.00732f
C17215 VPWR.n410 VGND 0.10877f
C17216 VPWR.t797 VGND 0.12017f
C17217 VPWR.t971 VGND 0.07889f
C17218 VPWR.t193 VGND 0.09265f
C17219 VPWR.t798 VGND 0.03348f
C17220 VPWR.t194 VGND 0.02976f
C17221 VPWR.n411 VGND 0.09198f
C17222 VPWR.n412 VGND 0.01806f
C17223 VPWR.n413 VGND 0.00732f
C17224 VPWR.n414 VGND 0.10877f
C17225 VPWR.t187 VGND 0.12017f
C17226 VPWR.t604 VGND 0.07889f
C17227 VPWR.t463 VGND 0.09265f
C17228 VPWR.t188 VGND 0.03348f
C17229 VPWR.t464 VGND 0.02976f
C17230 VPWR.n415 VGND 0.09198f
C17231 VPWR.n416 VGND 0.01806f
C17232 VPWR.n417 VGND 0.00732f
C17233 VPWR.n418 VGND 0.10877f
C17234 VPWR.t420 VGND 0.12017f
C17235 VPWR.t603 VGND 0.07889f
C17236 VPWR.t1825 VGND 0.09265f
C17237 VPWR.t421 VGND 0.03348f
C17238 VPWR.t1826 VGND 0.02976f
C17239 VPWR.n419 VGND 0.09198f
C17240 VPWR.n420 VGND 0.01806f
C17241 VPWR.n421 VGND 0.00732f
C17242 VPWR.n422 VGND 0.10877f
C17243 VPWR.t1819 VGND 0.12017f
C17244 VPWR.t973 VGND 0.07889f
C17245 VPWR.t1541 VGND 0.09265f
C17246 VPWR.t1820 VGND 0.03348f
C17247 VPWR.t1542 VGND 0.02976f
C17248 VPWR.n423 VGND 0.09198f
C17249 VPWR.n424 VGND 0.01806f
C17250 VPWR.n425 VGND 0.00732f
C17251 VPWR.n426 VGND 0.10877f
C17252 VPWR.t1535 VGND 0.12017f
C17253 VPWR.t684 VGND 0.07889f
C17254 VPWR.t835 VGND 0.09265f
C17255 VPWR.t1536 VGND 0.03348f
C17256 VPWR.t836 VGND 0.02976f
C17257 VPWR.n427 VGND 0.09198f
C17258 VPWR.n428 VGND 0.01806f
C17259 VPWR.n429 VGND 0.00732f
C17260 VPWR.n430 VGND 0.10877f
C17261 VPWR.t829 VGND 0.12017f
C17262 VPWR.t683 VGND 0.07889f
C17263 VPWR.t1739 VGND 0.09265f
C17264 VPWR.t830 VGND 0.03348f
C17265 VPWR.t1740 VGND 0.02976f
C17266 VPWR.n431 VGND 0.09198f
C17267 VPWR.n432 VGND 0.01806f
C17268 VPWR.n433 VGND 0.00732f
C17269 VPWR.n434 VGND 0.10877f
C17270 VPWR.t1600 VGND 0.12017f
C17271 VPWR.t970 VGND 0.07889f
C17272 VPWR.t1803 VGND 0.09265f
C17273 VPWR.t1601 VGND 0.03348f
C17274 VPWR.t1804 VGND 0.02976f
C17275 VPWR.n435 VGND 0.09198f
C17276 VPWR.n436 VGND 0.01806f
C17277 VPWR.n437 VGND 0.00732f
C17278 VPWR.n438 VGND 0.10877f
C17279 VPWR.t259 VGND 0.12017f
C17280 VPWR.t969 VGND 0.07889f
C17281 VPWR.t1547 VGND 0.09265f
C17282 VPWR.t260 VGND 0.03348f
C17283 VPWR.t1548 VGND 0.02976f
C17284 VPWR.n439 VGND 0.09198f
C17285 VPWR.n440 VGND 0.01806f
C17286 VPWR.n441 VGND 0.00732f
C17287 VPWR.n442 VGND 0.10877f
C17288 VPWR.t360 VGND 0.12017f
C17289 VPWR.t687 VGND 0.07889f
C17290 VPWR.t171 VGND 0.09265f
C17291 VPWR.t361 VGND 0.03348f
C17292 VPWR.t172 VGND 0.02976f
C17293 VPWR.n443 VGND 0.09198f
C17294 VPWR.n444 VGND 0.01806f
C17295 VPWR.n445 VGND 0.00732f
C17296 VPWR.n446 VGND 0.10877f
C17297 VPWR.t18 VGND 0.12017f
C17298 VPWR.t602 VGND 0.07889f
C17299 VPWR.t1113 VGND 0.13401f
C17300 VPWR.n447 VGND 0.07657f
C17301 VPWR.n448 VGND 0.01806f
C17302 VPWR.n449 VGND 0.13984f
C17303 VPWR.n450 VGND 1.02091f
C17304 VPWR.n451 VGND 0.13984f
C17305 VPWR.t1059 VGND 0.03348f
C17306 VPWR.t1226 VGND 0.02976f
C17307 VPWR.n452 VGND 0.09198f
C17308 VPWR.t20 VGND 0.09265f
C17309 VPWR.t1550 VGND 0.03348f
C17310 VPWR.t21 VGND 0.02976f
C17311 VPWR.n453 VGND 0.09198f
C17312 VPWR.n454 VGND 0.13984f
C17313 VPWR.n455 VGND 0.13984f
C17314 VPWR.t99 VGND 0.03348f
C17315 VPWR.t587 VGND 0.02976f
C17316 VPWR.n456 VGND 0.09198f
C17317 VPWR.t263 VGND 0.09265f
C17318 VPWR.t1008 VGND 0.03348f
C17319 VPWR.t264 VGND 0.02976f
C17320 VPWR.n457 VGND 0.09198f
C17321 VPWR.n458 VGND 0.13984f
C17322 VPWR.n459 VGND 0.13984f
C17323 VPWR.t644 VGND 0.03348f
C17324 VPWR.t210 VGND 0.02976f
C17325 VPWR.n460 VGND 0.09198f
C17326 VPWR.t647 VGND 0.09265f
C17327 VPWR.t65 VGND 0.03348f
C17328 VPWR.t648 VGND 0.02976f
C17329 VPWR.n461 VGND 0.09198f
C17330 VPWR.n462 VGND 0.13984f
C17331 VPWR.n463 VGND 0.13984f
C17332 VPWR.t408 VGND 0.03348f
C17333 VPWR.t73 VGND 0.02976f
C17334 VPWR.n464 VGND 0.09198f
C17335 VPWR.t411 VGND 0.09265f
C17336 VPWR.t458 VGND 0.03348f
C17337 VPWR.t412 VGND 0.02976f
C17338 VPWR.n465 VGND 0.09198f
C17339 VPWR.n466 VGND 0.13984f
C17340 VPWR.n467 VGND 0.13984f
C17341 VPWR.t301 VGND 0.03348f
C17342 VPWR.t214 VGND 0.02976f
C17343 VPWR.n468 VGND 0.09198f
C17344 VPWR.t304 VGND 0.09265f
C17345 VPWR.t945 VGND 0.03348f
C17346 VPWR.t305 VGND 0.02976f
C17347 VPWR.n469 VGND 0.09198f
C17348 VPWR.n470 VGND 0.13984f
C17349 VPWR.n471 VGND 0.13984f
C17350 VPWR.t850 VGND 0.03348f
C17351 VPWR.t949 VGND 0.02976f
C17352 VPWR.n472 VGND 0.09198f
C17353 VPWR.t853 VGND 0.09265f
C17354 VPWR.t154 VGND 0.03348f
C17355 VPWR.t854 VGND 0.02976f
C17356 VPWR.n473 VGND 0.09198f
C17357 VPWR.n474 VGND 0.13984f
C17358 VPWR.n475 VGND 0.13984f
C17359 VPWR.t1520 VGND 0.03348f
C17360 VPWR.t128 VGND 0.02976f
C17361 VPWR.n476 VGND 0.09198f
C17362 VPWR.t1499 VGND 0.09265f
C17363 VPWR.t914 VGND 0.03348f
C17364 VPWR.t1500 VGND 0.02976f
C17365 VPWR.n477 VGND 0.09198f
C17366 VPWR.n478 VGND 0.13984f
C17367 VPWR.n479 VGND 0.13984f
C17368 VPWR.t1843 VGND 0.03348f
C17369 VPWR.t1837 VGND 0.02976f
C17370 VPWR.n480 VGND 0.09198f
C17371 VPWR.t552 VGND 0.14585f
C17372 VPWR.t402 VGND 0.07889f
C17373 VPWR.t821 VGND 0.09265f
C17374 VPWR.t553 VGND 0.03348f
C17375 VPWR.t822 VGND 0.02976f
C17376 VPWR.n481 VGND 0.09198f
C17377 VPWR.t565 VGND 0.03348f
C17378 VPWR.t1746 VGND 0.02976f
C17379 VPWR.n482 VGND 0.09198f
C17380 VPWR.t564 VGND 0.14585f
C17381 VPWR.t1643 VGND 0.07889f
C17382 VPWR.t1745 VGND 0.09265f
C17383 VPWR.t25 VGND 0.03348f
C17384 VPWR.t1444 VGND 0.02976f
C17385 VPWR.n483 VGND 0.09198f
C17386 VPWR.n484 VGND 0.01806f
C17387 VPWR.n485 VGND 0.07657f
C17388 VPWR.t1443 VGND 0.13401f
C17389 VPWR.t76 VGND 0.07889f
C17390 VPWR.t24 VGND 0.12017f
C17391 VPWR.t353 VGND 0.03348f
C17392 VPWR.t174 VGND 0.02976f
C17393 VPWR.n486 VGND 0.09198f
C17394 VPWR.n487 VGND 0.01806f
C17395 VPWR.n488 VGND 0.00732f
C17396 VPWR.n489 VGND 0.10877f
C17397 VPWR.t173 VGND 0.09265f
C17398 VPWR.t739 VGND 0.07889f
C17399 VPWR.t352 VGND 0.12017f
C17400 VPWR.t1788 VGND 0.03348f
C17401 VPWR.t1043 VGND 0.02976f
C17402 VPWR.n490 VGND 0.09198f
C17403 VPWR.n491 VGND 0.01806f
C17404 VPWR.n492 VGND 0.00732f
C17405 VPWR.n493 VGND 0.10877f
C17406 VPWR.t1042 VGND 0.09265f
C17407 VPWR.t935 VGND 0.07889f
C17408 VPWR.t1787 VGND 0.12017f
C17409 VPWR.t216 VGND 0.03348f
C17410 VPWR.t872 VGND 0.02976f
C17411 VPWR.n494 VGND 0.09198f
C17412 VPWR.n495 VGND 0.01806f
C17413 VPWR.n496 VGND 0.00732f
C17414 VPWR.n497 VGND 0.10877f
C17415 VPWR.t871 VGND 0.09265f
C17416 VPWR.t936 VGND 0.07889f
C17417 VPWR.t215 VGND 0.12017f
C17418 VPWR.t998 VGND 0.03348f
C17419 VPWR.t894 VGND 0.02976f
C17420 VPWR.n498 VGND 0.09198f
C17421 VPWR.n499 VGND 0.01806f
C17422 VPWR.n500 VGND 0.00732f
C17423 VPWR.n501 VGND 0.10877f
C17424 VPWR.t893 VGND 0.09265f
C17425 VPWR.t735 VGND 0.07889f
C17426 VPWR.t997 VGND 0.12017f
C17427 VPWR.t329 VGND 0.03348f
C17428 VPWR.t1002 VGND 0.02976f
C17429 VPWR.n502 VGND 0.09198f
C17430 VPWR.n503 VGND 0.01806f
C17431 VPWR.n504 VGND 0.00732f
C17432 VPWR.n505 VGND 0.10877f
C17433 VPWR.t1001 VGND 0.09265f
C17434 VPWR.t736 VGND 0.07889f
C17435 VPWR.t328 VGND 0.12017f
C17436 VPWR.t450 VGND 0.03348f
C17437 VPWR.t339 VGND 0.02976f
C17438 VPWR.n506 VGND 0.09198f
C17439 VPWR.n507 VGND 0.01806f
C17440 VPWR.n508 VGND 0.00732f
C17441 VPWR.n509 VGND 0.10877f
C17442 VPWR.t338 VGND 0.09265f
C17443 VPWR.t74 VGND 0.07889f
C17444 VPWR.t449 VGND 0.12017f
C17445 VPWR.t146 VGND 0.03348f
C17446 VPWR.t454 VGND 0.02976f
C17447 VPWR.n510 VGND 0.09198f
C17448 VPWR.n511 VGND 0.01806f
C17449 VPWR.n512 VGND 0.00732f
C17450 VPWR.n513 VGND 0.10877f
C17451 VPWR.t453 VGND 0.09265f
C17452 VPWR.t1640 VGND 0.07889f
C17453 VPWR.t145 VGND 0.12017f
C17454 VPWR.t196 VGND 0.03348f
C17455 VPWR.t1698 VGND 0.02976f
C17456 VPWR.n514 VGND 0.09198f
C17457 VPWR.n515 VGND 0.01806f
C17458 VPWR.n516 VGND 0.00732f
C17459 VPWR.n517 VGND 0.10877f
C17460 VPWR.t1697 VGND 0.09265f
C17461 VPWR.t1641 VGND 0.07889f
C17462 VPWR.t195 VGND 0.12017f
C17463 VPWR.t784 VGND 0.03348f
C17464 VPWR.t266 VGND 0.02976f
C17465 VPWR.n518 VGND 0.09198f
C17466 VPWR.n519 VGND 0.01806f
C17467 VPWR.n520 VGND 0.00732f
C17468 VPWR.n521 VGND 0.10877f
C17469 VPWR.t265 VGND 0.09265f
C17470 VPWR.t937 VGND 0.07889f
C17471 VPWR.t783 VGND 0.12017f
C17472 VPWR.t404 VGND 0.03348f
C17473 VPWR.t788 VGND 0.02976f
C17474 VPWR.n522 VGND 0.09198f
C17475 VPWR.n523 VGND 0.01806f
C17476 VPWR.n524 VGND 0.00732f
C17477 VPWR.n525 VGND 0.10877f
C17478 VPWR.t787 VGND 0.09265f
C17479 VPWR.t938 VGND 0.07889f
C17480 VPWR.t403 VGND 0.12017f
C17481 VPWR.t132 VGND 0.03348f
C17482 VPWR.t977 VGND 0.02976f
C17483 VPWR.n526 VGND 0.09198f
C17484 VPWR.n527 VGND 0.01806f
C17485 VPWR.n528 VGND 0.00732f
C17486 VPWR.n529 VGND 0.10877f
C17487 VPWR.t976 VGND 0.09265f
C17488 VPWR.t1642 VGND 0.07889f
C17489 VPWR.t131 VGND 0.12017f
C17490 VPWR.t1498 VGND 0.03348f
C17491 VPWR.t1831 VGND 0.02976f
C17492 VPWR.n530 VGND 0.09198f
C17493 VPWR.n531 VGND 0.01806f
C17494 VPWR.n532 VGND 0.00732f
C17495 VPWR.n533 VGND 0.10877f
C17496 VPWR.t1830 VGND 0.09265f
C17497 VPWR.t737 VGND 0.07889f
C17498 VPWR.t1497 VGND 0.12017f
C17499 VPWR.t1668 VGND 0.03348f
C17500 VPWR.t1472 VGND 0.02976f
C17501 VPWR.n534 VGND 0.09198f
C17502 VPWR.n535 VGND 0.01806f
C17503 VPWR.n536 VGND 0.00732f
C17504 VPWR.n537 VGND 0.10877f
C17505 VPWR.t1471 VGND 0.09265f
C17506 VPWR.t738 VGND 0.07889f
C17507 VPWR.t1667 VGND 0.12017f
C17508 VPWR.t922 VGND 0.03348f
C17509 VPWR.t1672 VGND 0.02976f
C17510 VPWR.n538 VGND 0.09198f
C17511 VPWR.n539 VGND 0.01806f
C17512 VPWR.n540 VGND 0.00732f
C17513 VPWR.n541 VGND 0.10877f
C17514 VPWR.t1671 VGND 0.09265f
C17515 VPWR.t75 VGND 0.07889f
C17516 VPWR.t921 VGND 0.12017f
C17517 VPWR.n542 VGND 0.10877f
C17518 VPWR.n543 VGND 0.00732f
C17519 VPWR.n544 VGND 0.01806f
C17520 VPWR.n545 VGND 0.13984f
C17521 VPWR.n546 VGND 1.01451f
C17522 VPWR.n547 VGND 0.13984f
C17523 VPWR.t579 VGND 0.03348f
C17524 VPWR.t632 VGND 0.02976f
C17525 VPWR.n548 VGND 0.09198f
C17526 VPWR.t578 VGND 0.14585f
C17527 VPWR.t1887 VGND 0.07889f
C17528 VPWR.t631 VGND 0.09265f
C17529 VPWR.t1578 VGND 0.12017f
C17530 VPWR.t1558 VGND 0.03348f
C17531 VPWR.t1587 VGND 0.02976f
C17532 VPWR.n549 VGND 0.09198f
C17533 VPWR.n550 VGND 0.13984f
C17534 VPWR.n551 VGND 0.13984f
C17535 VPWR.t1579 VGND 0.03348f
C17536 VPWR.t1512 VGND 0.02976f
C17537 VPWR.n552 VGND 0.09198f
C17538 VPWR.t1655 VGND 0.07889f
C17539 VPWR.t1511 VGND 0.09265f
C17540 VPWR.t320 VGND 0.12017f
C17541 VPWR.t1474 VGND 0.03348f
C17542 VPWR.t1812 VGND 0.02976f
C17543 VPWR.n553 VGND 0.09198f
C17544 VPWR.n554 VGND 0.13984f
C17545 VPWR.n555 VGND 0.13984f
C17546 VPWR.t321 VGND 0.03348f
C17547 VPWR.t743 VGND 0.02976f
C17548 VPWR.n556 VGND 0.09198f
C17549 VPWR.t1886 VGND 0.07889f
C17550 VPWR.t742 VGND 0.09265f
C17551 VPWR.t1753 VGND 0.12017f
C17552 VPWR.t1875 VGND 0.03348f
C17553 VPWR.t1762 VGND 0.02976f
C17554 VPWR.n557 VGND 0.09198f
C17555 VPWR.n558 VGND 0.13984f
C17556 VPWR.n559 VGND 0.13984f
C17557 VPWR.t1754 VGND 0.03348f
C17558 VPWR.t13 VGND 0.02976f
C17559 VPWR.n560 VGND 0.09198f
C17560 VPWR.t1659 VGND 0.07889f
C17561 VPWR.t12 VGND 0.09265f
C17562 VPWR.t1703 VGND 0.12017f
C17563 VPWR.t5 VGND 0.03348f
C17564 VPWR.t162 VGND 0.02976f
C17565 VPWR.n561 VGND 0.09198f
C17566 VPWR.n562 VGND 0.13984f
C17567 VPWR.n563 VGND 0.13984f
C17568 VPWR.t1704 VGND 0.03348f
C17569 VPWR.t182 VGND 0.02976f
C17570 VPWR.n564 VGND 0.09198f
C17571 VPWR.t1884 VGND 0.07889f
C17572 VPWR.t181 VGND 0.09265f
C17573 VPWR.t762 VGND 0.12017f
C17574 VPWR.t140 VGND 0.03348f
C17575 VPWR.t61 VGND 0.02976f
C17576 VPWR.n565 VGND 0.09198f
C17577 VPWR.n566 VGND 0.13984f
C17578 VPWR.n567 VGND 0.13984f
C17579 VPWR.t763 VGND 0.03348f
C17580 VPWR.t593 VGND 0.02976f
C17581 VPWR.n568 VGND 0.09198f
C17582 VPWR.t1923 VGND 0.07889f
C17583 VPWR.t592 VGND 0.09265f
C17584 VPWR.t669 VGND 0.12017f
C17585 VPWR.t393 VGND 0.03348f
C17586 VPWR.t1004 VGND 0.02976f
C17587 VPWR.n569 VGND 0.09198f
C17588 VPWR.n570 VGND 0.13984f
C17589 VPWR.n571 VGND 0.13984f
C17590 VPWR.t670 VGND 0.03348f
C17591 VPWR.t252 VGND 0.02976f
C17592 VPWR.n572 VGND 0.09198f
C17593 VPWR.t1658 VGND 0.07889f
C17594 VPWR.t251 VGND 0.09265f
C17595 VPWR.t598 VGND 0.12017f
C17596 VPWR.t878 VGND 0.03348f
C17597 VPWR.t1055 VGND 0.02976f
C17598 VPWR.n573 VGND 0.09198f
C17599 VPWR.n574 VGND 0.13984f
C17600 VPWR.n575 VGND 0.13984f
C17601 VPWR.t599 VGND 0.03348f
C17602 VPWR.t1712 VGND 0.02976f
C17603 VPWR.n576 VGND 0.09198f
C17604 VPWR.t1656 VGND 0.07889f
C17605 VPWR.t1711 VGND 0.09265f
C17606 VPWR.t226 VGND 0.03348f
C17607 VPWR.t1293 VGND 0.02976f
C17608 VPWR.n577 VGND 0.09198f
C17609 VPWR.t31 VGND 0.03348f
C17610 VPWR.t1401 VGND 0.02976f
C17611 VPWR.n578 VGND 0.09198f
C17612 VPWR.t570 VGND 0.14585f
C17613 VPWR.t367 VGND 0.07889f
C17614 VPWR.t1751 VGND 0.09265f
C17615 VPWR.t571 VGND 0.03348f
C17616 VPWR.t1752 VGND 0.02976f
C17617 VPWR.n579 VGND 0.09198f
C17618 VPWR.n580 VGND 0.01806f
C17619 VPWR.n581 VGND 0.00732f
C17620 VPWR.n582 VGND 0.10877f
C17621 VPWR.t1741 VGND 0.12017f
C17622 VPWR.t362 VGND 0.07889f
C17623 VPWR.t681 VGND 0.09265f
C17624 VPWR.t1742 VGND 0.03348f
C17625 VPWR.t682 VGND 0.02976f
C17626 VPWR.n583 VGND 0.09198f
C17627 VPWR.n584 VGND 0.01806f
C17628 VPWR.n585 VGND 0.00732f
C17629 VPWR.n586 VGND 0.10877f
C17630 VPWR.t701 VGND 0.12017f
C17631 VPWR.t351 VGND 0.07889f
C17632 VPWR.t1463 VGND 0.09265f
C17633 VPWR.t702 VGND 0.03348f
C17634 VPWR.t1464 VGND 0.02976f
C17635 VPWR.n587 VGND 0.09198f
C17636 VPWR.n588 VGND 0.01806f
C17637 VPWR.n589 VGND 0.00732f
C17638 VPWR.n590 VGND 0.10877f
C17639 VPWR.t1487 VGND 0.12017f
C17640 VPWR.t350 VGND 0.07889f
C17641 VPWR.t322 VGND 0.09265f
C17642 VPWR.t1488 VGND 0.03348f
C17643 VPWR.t323 VGND 0.02976f
C17644 VPWR.n591 VGND 0.09198f
C17645 VPWR.n592 VGND 0.01806f
C17646 VPWR.n593 VGND 0.00732f
C17647 VPWR.n594 VGND 0.10877f
C17648 VPWR.t1725 VGND 0.12017f
C17649 VPWR.t366 VGND 0.07889f
C17650 VPWR.t754 VGND 0.09265f
C17651 VPWR.t1726 VGND 0.03348f
C17652 VPWR.t755 VGND 0.02976f
C17653 VPWR.n595 VGND 0.09198f
C17654 VPWR.n596 VGND 0.01806f
C17655 VPWR.n597 VGND 0.00732f
C17656 VPWR.n598 VGND 0.10877f
C17657 VPWR.t748 VGND 0.12017f
C17658 VPWR.t847 VGND 0.07889f
C17659 VPWR.t807 VGND 0.09265f
C17660 VPWR.t749 VGND 0.03348f
C17661 VPWR.t808 VGND 0.02976f
C17662 VPWR.n599 VGND 0.09198f
C17663 VPWR.n600 VGND 0.01806f
C17664 VPWR.n601 VGND 0.00732f
C17665 VPWR.n602 VGND 0.10877f
C17666 VPWR.t793 VGND 0.12017f
C17667 VPWR.t846 VGND 0.07889f
C17668 VPWR.t277 VGND 0.09265f
C17669 VPWR.t794 VGND 0.03348f
C17670 VPWR.t278 VGND 0.02976f
C17671 VPWR.n603 VGND 0.09198f
C17672 VPWR.n604 VGND 0.01806f
C17673 VPWR.n605 VGND 0.00732f
C17674 VPWR.n606 VGND 0.10877f
C17675 VPWR.t271 VGND 0.12017f
C17676 VPWR.t365 VGND 0.07889f
C17677 VPWR.t1709 VGND 0.09265f
C17678 VPWR.t272 VGND 0.03348f
C17679 VPWR.t1710 VGND 0.02976f
C17680 VPWR.n607 VGND 0.09198f
C17681 VPWR.n608 VGND 0.01806f
C17682 VPWR.n609 VGND 0.00732f
C17683 VPWR.n610 VGND 0.10877f
C17684 VPWR.t1854 VGND 0.12017f
C17685 VPWR.t364 VGND 0.07889f
C17686 VPWR.t665 VGND 0.09265f
C17687 VPWR.t1855 VGND 0.03348f
C17688 VPWR.t666 VGND 0.02976f
C17689 VPWR.n611 VGND 0.09198f
C17690 VPWR.n612 VGND 0.01806f
C17691 VPWR.n613 VGND 0.00732f
C17692 VPWR.n614 VGND 0.10877f
C17693 VPWR.t659 VGND 0.12017f
C17694 VPWR.t848 VGND 0.07889f
C17695 VPWR.t535 VGND 0.09265f
C17696 VPWR.t660 VGND 0.03348f
C17697 VPWR.t536 VGND 0.02976f
C17698 VPWR.n615 VGND 0.09198f
C17699 VPWR.n616 VGND 0.01806f
C17700 VPWR.n617 VGND 0.00732f
C17701 VPWR.n618 VGND 0.10877f
C17702 VPWR.t334 VGND 0.12017f
C17703 VPWR.t349 VGND 0.07889f
C17704 VPWR.t1632 VGND 0.09265f
C17705 VPWR.t335 VGND 0.03348f
C17706 VPWR.t1633 VGND 0.02976f
C17707 VPWR.n619 VGND 0.09198f
C17708 VPWR.n620 VGND 0.01806f
C17709 VPWR.n621 VGND 0.00732f
C17710 VPWR.n622 VGND 0.10877f
C17711 VPWR.t1626 VGND 0.12017f
C17712 VPWR.t348 VGND 0.07889f
C17713 VPWR.t991 VGND 0.09265f
C17714 VPWR.t1627 VGND 0.03348f
C17715 VPWR.t992 VGND 0.02976f
C17716 VPWR.n623 VGND 0.09198f
C17717 VPWR.n624 VGND 0.01806f
C17718 VPWR.n625 VGND 0.00732f
C17719 VPWR.n626 VGND 0.10877f
C17720 VPWR.t889 VGND 0.12017f
C17721 VPWR.t845 VGND 0.07889f
C17722 VPWR.t90 VGND 0.09265f
C17723 VPWR.t890 VGND 0.03348f
C17724 VPWR.t91 VGND 0.02976f
C17725 VPWR.n627 VGND 0.09198f
C17726 VPWR.n628 VGND 0.01806f
C17727 VPWR.n629 VGND 0.00732f
C17728 VPWR.n630 VGND 0.10877f
C17729 VPWR.t1795 VGND 0.12017f
C17730 VPWR.t844 VGND 0.07889f
C17731 VPWR.t1048 VGND 0.09265f
C17732 VPWR.t1796 VGND 0.03348f
C17733 VPWR.t1049 VGND 0.02976f
C17734 VPWR.n631 VGND 0.09198f
C17735 VPWR.n632 VGND 0.01806f
C17736 VPWR.n633 VGND 0.00732f
C17737 VPWR.n634 VGND 0.10877f
C17738 VPWR.t637 VGND 0.12017f
C17739 VPWR.t843 VGND 0.07889f
C17740 VPWR.t227 VGND 0.09265f
C17741 VPWR.t638 VGND 0.03348f
C17742 VPWR.t228 VGND 0.02976f
C17743 VPWR.n635 VGND 0.09198f
C17744 VPWR.n636 VGND 0.01806f
C17745 VPWR.n637 VGND 0.00732f
C17746 VPWR.n638 VGND 0.10877f
C17747 VPWR.t30 VGND 0.12017f
C17748 VPWR.t363 VGND 0.07889f
C17749 VPWR.t1400 VGND 0.13401f
C17750 VPWR.n639 VGND 0.07657f
C17751 VPWR.n640 VGND 0.01806f
C17752 VPWR.n641 VGND 0.13984f
C17753 VPWR.n642 VGND 1.02091f
C17754 VPWR.n643 VGND 0.13984f
C17755 VPWR.t1716 VGND 0.03348f
C17756 VPWR.t1127 VGND 0.02976f
C17757 VPWR.n644 VGND 0.09198f
C17758 VPWR.t165 VGND 0.09265f
C17759 VPWR.t357 VGND 0.03348f
C17760 VPWR.t166 VGND 0.02976f
C17761 VPWR.n645 VGND 0.09198f
C17762 VPWR.n646 VGND 0.13984f
C17763 VPWR.n647 VGND 0.13984f
C17764 VPWR.t256 VGND 0.03348f
C17765 VPWR.t1544 VGND 0.02976f
C17766 VPWR.n648 VGND 0.09198f
C17767 VPWR.t1799 VGND 0.09265f
C17768 VPWR.t1597 VGND 0.03348f
C17769 VPWR.t1800 VGND 0.02976f
C17770 VPWR.n649 VGND 0.09198f
C17771 VPWR.n650 VGND 0.13984f
C17772 VPWR.n651 VGND 0.13984f
C17773 VPWR.t826 VGND 0.03348f
C17774 VPWR.t1736 VGND 0.02976f
C17775 VPWR.n652 VGND 0.09198f
C17776 VPWR.t831 VGND 0.09265f
C17777 VPWR.t1532 VGND 0.03348f
C17778 VPWR.t832 VGND 0.02976f
C17779 VPWR.n653 VGND 0.09198f
C17780 VPWR.n654 VGND 0.13984f
C17781 VPWR.n655 VGND 0.13984f
C17782 VPWR.t868 VGND 0.03348f
C17783 VPWR.t1538 VGND 0.02976f
C17784 VPWR.n656 VGND 0.09198f
C17785 VPWR.t1821 VGND 0.09265f
C17786 VPWR.t417 VGND 0.03348f
C17787 VPWR.t1822 VGND 0.02976f
C17788 VPWR.n657 VGND 0.09198f
C17789 VPWR.n658 VGND 0.13984f
C17790 VPWR.n659 VGND 0.13984f
C17791 VPWR.t311 VGND 0.03348f
C17792 VPWR.t460 VGND 0.02976f
C17793 VPWR.n660 VGND 0.09198f
C17794 VPWR.t189 VGND 0.09265f
C17795 VPWR.t1678 VGND 0.03348f
C17796 VPWR.t190 VGND 0.02976f
C17797 VPWR.n661 VGND 0.09198f
C17798 VPWR.n662 VGND 0.13984f
C17799 VPWR.n663 VGND 0.13984f
C17800 VPWR.t1076 VGND 0.03348f
C17801 VPWR.t800 VGND 0.02976f
C17802 VPWR.n664 VGND 0.09198f
C17803 VPWR.t77 VGND 0.09265f
C17804 VPWR.t1816 VGND 0.03348f
C17805 VPWR.t78 VGND 0.02976f
C17806 VPWR.n665 VGND 0.09198f
C17807 VPWR.n666 VGND 0.13984f
C17808 VPWR.n667 VGND 0.13984f
C17809 VPWR.t1510 VGND 0.03348f
C17810 VPWR.t1728 VGND 0.02976f
C17811 VPWR.n668 VGND 0.09198f
C17812 VPWR.t1483 VGND 0.09265f
C17813 VPWR.t723 VGND 0.03348f
C17814 VPWR.t1484 VGND 0.02976f
C17815 VPWR.n669 VGND 0.09198f
C17816 VPWR.n670 VGND 0.13984f
C17817 VPWR.n671 VGND 0.13984f
C17818 VPWR.t285 VGND 0.03348f
C17819 VPWR.t729 VGND 0.02976f
C17820 VPWR.n672 VGND 0.09198f
C17821 VPWR.t558 VGND 0.14585f
C17822 VPWR.t446 VGND 0.07889f
C17823 VPWR.t692 VGND 0.09265f
C17824 VPWR.t559 VGND 0.03348f
C17825 VPWR.t693 VGND 0.02976f
C17826 VPWR.n673 VGND 0.09198f
C17827 VPWR.t551 VGND 0.03348f
C17828 VPWR.t1847 VGND 0.02976f
C17829 VPWR.n674 VGND 0.09198f
C17830 VPWR.t550 VGND 0.14585f
C17831 VPWR.t774 VGND 0.07889f
C17832 VPWR.t1846 VGND 0.09265f
C17833 VPWR.t236 VGND 0.03348f
C17834 VPWR.t1234 VGND 0.02976f
C17835 VPWR.n675 VGND 0.09198f
C17836 VPWR.n676 VGND 0.01806f
C17837 VPWR.n677 VGND 0.07657f
C17838 VPWR.t1233 VGND 0.13401f
C17839 VPWR.t1602 VGND 0.07889f
C17840 VPWR.t235 VGND 0.12017f
C17841 VPWR.t1057 VGND 0.03348f
C17842 VPWR.t1720 VGND 0.02976f
C17843 VPWR.n678 VGND 0.09198f
C17844 VPWR.n679 VGND 0.01806f
C17845 VPWR.n680 VGND 0.00732f
C17846 VPWR.n681 VGND 0.10877f
C17847 VPWR.t1719 VGND 0.09265f
C17848 VPWR.t83 VGND 0.07889f
C17849 VPWR.t1056 VGND 0.12017f
C17850 VPWR.t97 VGND 0.03348f
C17851 VPWR.t583 VGND 0.02976f
C17852 VPWR.n682 VGND 0.09198f
C17853 VPWR.n683 VGND 0.01806f
C17854 VPWR.n684 VGND 0.00732f
C17855 VPWR.n685 VGND 0.10877f
C17856 VPWR.t582 VGND 0.09265f
C17857 VPWR.t84 VGND 0.07889f
C17858 VPWR.t96 VGND 0.12017f
C17859 VPWR.t1006 VGND 0.03348f
C17860 VPWR.t262 VGND 0.02976f
C17861 VPWR.n686 VGND 0.09198f
C17862 VPWR.n687 VGND 0.01806f
C17863 VPWR.n688 VGND 0.00732f
C17864 VPWR.n689 VGND 0.10877f
C17865 VPWR.t261 VGND 0.09265f
C17866 VPWR.t85 VGND 0.07889f
C17867 VPWR.t1005 VGND 0.12017f
C17868 VPWR.t597 VGND 0.03348f
C17869 VPWR.t206 VGND 0.02976f
C17870 VPWR.n690 VGND 0.09198f
C17871 VPWR.n691 VGND 0.01806f
C17872 VPWR.n692 VGND 0.00732f
C17873 VPWR.n693 VGND 0.10877f
C17874 VPWR.t205 VGND 0.09265f
C17875 VPWR.t653 VGND 0.07889f
C17876 VPWR.t596 VGND 0.12017f
C17877 VPWR.t63 VGND 0.03348f
C17878 VPWR.t646 VGND 0.02976f
C17879 VPWR.n694 VGND 0.09198f
C17880 VPWR.n695 VGND 0.01806f
C17881 VPWR.n696 VGND 0.00732f
C17882 VPWR.n697 VGND 0.10877f
C17883 VPWR.t645 VGND 0.09265f
C17884 VPWR.t654 VGND 0.07889f
C17885 VPWR.t62 VGND 0.12017f
C17886 VPWR.t406 VGND 0.03348f
C17887 VPWR.t69 VGND 0.02976f
C17888 VPWR.n698 VGND 0.09198f
C17889 VPWR.n699 VGND 0.01806f
C17890 VPWR.n700 VGND 0.00732f
C17891 VPWR.n701 VGND 0.10877f
C17892 VPWR.t68 VGND 0.09265f
C17893 VPWR.t939 VGND 0.07889f
C17894 VPWR.t405 VGND 0.12017f
C17895 VPWR.t204 VGND 0.03348f
C17896 VPWR.t410 VGND 0.02976f
C17897 VPWR.n702 VGND 0.09198f
C17898 VPWR.n703 VGND 0.01806f
C17899 VPWR.n704 VGND 0.00732f
C17900 VPWR.n705 VGND 0.10877f
C17901 VPWR.t409 VGND 0.09265f
C17902 VPWR.t1603 VGND 0.07889f
C17903 VPWR.t203 VGND 0.12017f
C17904 VPWR.t299 VGND 0.03348f
C17905 VPWR.t212 VGND 0.02976f
C17906 VPWR.n706 VGND 0.09198f
C17907 VPWR.n707 VGND 0.01806f
C17908 VPWR.n708 VGND 0.00732f
C17909 VPWR.n709 VGND 0.10877f
C17910 VPWR.t211 VGND 0.09265f
C17911 VPWR.t772 VGND 0.07889f
C17912 VPWR.t298 VGND 0.12017f
C17913 VPWR.t943 VGND 0.03348f
C17914 VPWR.t303 VGND 0.02976f
C17915 VPWR.n710 VGND 0.09198f
C17916 VPWR.n711 VGND 0.01806f
C17917 VPWR.n712 VGND 0.00732f
C17918 VPWR.n713 VGND 0.10877f
C17919 VPWR.t302 VGND 0.09265f
C17920 VPWR.t86 VGND 0.07889f
C17921 VPWR.t942 VGND 0.12017f
C17922 VPWR.t747 VGND 0.03348f
C17923 VPWR.t947 VGND 0.02976f
C17924 VPWR.n714 VGND 0.09198f
C17925 VPWR.n715 VGND 0.01806f
C17926 VPWR.n716 VGND 0.00732f
C17927 VPWR.n717 VGND 0.10877f
C17928 VPWR.t946 VGND 0.09265f
C17929 VPWR.t87 VGND 0.07889f
C17930 VPWR.t746 VGND 0.12017f
C17931 VPWR.t152 VGND 0.03348f
C17932 VPWR.t852 VGND 0.02976f
C17933 VPWR.n718 VGND 0.09198f
C17934 VPWR.n719 VGND 0.01806f
C17935 VPWR.n720 VGND 0.00732f
C17936 VPWR.n721 VGND 0.10877f
C17937 VPWR.t851 VGND 0.09265f
C17938 VPWR.t773 VGND 0.07889f
C17939 VPWR.t151 VGND 0.12017f
C17940 VPWR.t1522 VGND 0.03348f
C17941 VPWR.t1575 VGND 0.02976f
C17942 VPWR.n722 VGND 0.09198f
C17943 VPWR.n723 VGND 0.01806f
C17944 VPWR.n724 VGND 0.00732f
C17945 VPWR.n725 VGND 0.10877f
C17946 VPWR.t1574 VGND 0.09265f
C17947 VPWR.t655 VGND 0.07889f
C17948 VPWR.t1521 VGND 0.12017f
C17949 VPWR.t912 VGND 0.03348f
C17950 VPWR.t1502 VGND 0.02976f
C17951 VPWR.n726 VGND 0.09198f
C17952 VPWR.n727 VGND 0.01806f
C17953 VPWR.n728 VGND 0.00732f
C17954 VPWR.n729 VGND 0.10877f
C17955 VPWR.t1501 VGND 0.09265f
C17956 VPWR.t656 VGND 0.07889f
C17957 VPWR.t911 VGND 0.12017f
C17958 VPWR.t634 VGND 0.03348f
C17959 VPWR.t1835 VGND 0.02976f
C17960 VPWR.n730 VGND 0.09198f
C17961 VPWR.n731 VGND 0.01806f
C17962 VPWR.n732 VGND 0.00732f
C17963 VPWR.n733 VGND 0.10877f
C17964 VPWR.t1834 VGND 0.09265f
C17965 VPWR.t940 VGND 0.07889f
C17966 VPWR.t633 VGND 0.12017f
C17967 VPWR.n734 VGND 0.10877f
C17968 VPWR.n735 VGND 0.00732f
C17969 VPWR.n736 VGND 0.01806f
C17970 VPWR.n737 VGND 0.13984f
C17971 VPWR.n738 VGND 1.01451f
C17972 VPWR.n739 VGND 0.13984f
C17973 VPWR.t555 VGND 0.03348f
C17974 VPWR.t824 VGND 0.02976f
C17975 VPWR.n740 VGND 0.09198f
C17976 VPWR.t554 VGND 0.14585f
C17977 VPWR.t1036 VGND 0.07889f
C17978 VPWR.t823 VGND 0.09265f
C17979 VPWR.t1838 VGND 0.12017f
C17980 VPWR.t820 VGND 0.03348f
C17981 VPWR.t1841 VGND 0.02976f
C17982 VPWR.n741 VGND 0.09198f
C17983 VPWR.n742 VGND 0.13984f
C17984 VPWR.n743 VGND 0.13984f
C17985 VPWR.t1839 VGND 0.03348f
C17986 VPWR.t1492 VGND 0.02976f
C17987 VPWR.n744 VGND 0.09198f
C17988 VPWR.t985 VGND 0.07889f
C17989 VPWR.t1491 VGND 0.09265f
C17990 VPWR.t1805 VGND 0.12017f
C17991 VPWR.t1516 VGND 0.03348f
C17992 VPWR.t130 VGND 0.02976f
C17993 VPWR.n745 VGND 0.09198f
C17994 VPWR.n746 VGND 0.13984f
C17995 VPWR.n747 VGND 0.13984f
C17996 VPWR.t1806 VGND 0.03348f
C17997 VPWR.t1074 VGND 0.02976f
C17998 VPWR.n748 VGND 0.09198f
C17999 VPWR.t1035 VGND 0.07889f
C18000 VPWR.t1073 VGND 0.09265f
C18001 VPWR.t950 VGND 0.12017f
C18002 VPWR.t856 VGND 0.03348f
C18003 VPWR.t1676 VGND 0.02976f
C18004 VPWR.n749 VGND 0.09198f
C18005 VPWR.n750 VGND 0.13984f
C18006 VPWR.n751 VGND 0.13984f
C18007 VPWR.t951 VGND 0.03348f
C18008 VPWR.t309 VGND 0.02976f
C18009 VPWR.n752 VGND 0.09198f
C18010 VPWR.t1038 VGND 0.07889f
C18011 VPWR.t308 VGND 0.09265f
C18012 VPWR.t155 VGND 0.12017f
C18013 VPWR.t307 VGND 0.03348f
C18014 VPWR.t148 VGND 0.02976f
C18015 VPWR.n753 VGND 0.09198f
C18016 VPWR.n754 VGND 0.13984f
C18017 VPWR.n755 VGND 0.13984f
C18018 VPWR.t156 VGND 0.03348f
C18019 VPWR.t866 VGND 0.02976f
C18020 VPWR.n756 VGND 0.09198f
C18021 VPWR.t1033 VGND 0.07889f
C18022 VPWR.t865 VGND 0.09265f
C18023 VPWR.t70 VGND 0.12017f
C18024 VPWR.t864 VGND 0.03348f
C18025 VPWR.t1530 VGND 0.02976f
C18026 VPWR.n757 VGND 0.09198f
C18027 VPWR.n758 VGND 0.13984f
C18028 VPWR.n759 VGND 0.13984f
C18029 VPWR.t71 VGND 0.03348f
C18030 VPWR.t1917 VGND 0.02976f
C18031 VPWR.n760 VGND 0.09198f
C18032 VPWR.t983 VGND 0.07889f
C18033 VPWR.t1916 VGND 0.09265f
C18034 VPWR.t207 VGND 0.12017f
C18035 VPWR.t1915 VGND 0.03348f
C18036 VPWR.t1595 VGND 0.02976f
C18037 VPWR.n761 VGND 0.09198f
C18038 VPWR.n762 VGND 0.13984f
C18039 VPWR.n763 VGND 0.13984f
C18040 VPWR.t208 VGND 0.03348f
C18041 VPWR.t1790 VGND 0.02976f
C18042 VPWR.n764 VGND 0.09198f
C18043 VPWR.t1037 VGND 0.07889f
C18044 VPWR.t1789 VGND 0.09265f
C18045 VPWR.t584 VGND 0.12017f
C18046 VPWR.t246 VGND 0.03348f
C18047 VPWR.t589 VGND 0.02976f
C18048 VPWR.n765 VGND 0.09198f
C18049 VPWR.n766 VGND 0.13984f
C18050 VPWR.n767 VGND 0.13984f
C18051 VPWR.t585 VGND 0.03348f
C18052 VPWR.t23 VGND 0.02976f
C18053 VPWR.n768 VGND 0.09198f
C18054 VPWR.t986 VGND 0.07889f
C18055 VPWR.t22 VGND 0.09265f
C18056 VPWR.t1061 VGND 0.03348f
C18057 VPWR.t1194 VGND 0.02976f
C18058 VPWR.n769 VGND 0.09198f
C18059 VPWR.t222 VGND 0.03348f
C18060 VPWR.t1299 VGND 0.02976f
C18061 VPWR.n770 VGND 0.09198f
C18062 VPWR.t576 VGND 0.14585f
C18063 VPWR.t1897 VGND 0.07889f
C18064 VPWR.t629 VGND 0.09265f
C18065 VPWR.t577 VGND 0.03348f
C18066 VPWR.t630 VGND 0.02976f
C18067 VPWR.n771 VGND 0.09198f
C18068 VPWR.n772 VGND 0.01806f
C18069 VPWR.n773 VGND 0.00732f
C18070 VPWR.n774 VGND 0.10877f
C18071 VPWR.t1555 VGND 0.12017f
C18072 VPWR.t1895 VGND 0.07889f
C18073 VPWR.t1582 VGND 0.09265f
C18074 VPWR.t1556 VGND 0.03348f
C18075 VPWR.t1583 VGND 0.02976f
C18076 VPWR.n775 VGND 0.09198f
C18077 VPWR.n776 VGND 0.01806f
C18078 VPWR.n777 VGND 0.00732f
C18079 VPWR.n778 VGND 0.10877f
C18080 VPWR.t679 VGND 0.12017f
C18081 VPWR.t119 VGND 0.07889f
C18082 VPWR.t1495 VGND 0.09265f
C18083 VPWR.t680 VGND 0.03348f
C18084 VPWR.t1496 VGND 0.02976f
C18085 VPWR.n779 VGND 0.09198f
C18086 VPWR.n780 VGND 0.01806f
C18087 VPWR.n781 VGND 0.00732f
C18088 VPWR.n782 VGND 0.10877f
C18089 VPWR.t1475 VGND 0.12017f
C18090 VPWR.t120 VGND 0.07889f
C18091 VPWR.t1809 VGND 0.09265f
C18092 VPWR.t1476 VGND 0.03348f
C18093 VPWR.t1810 VGND 0.02976f
C18094 VPWR.n783 VGND 0.09198f
C18095 VPWR.n784 VGND 0.01806f
C18096 VPWR.n785 VGND 0.00732f
C18097 VPWR.n786 VGND 0.10877f
C18098 VPWR.t316 VGND 0.12017f
C18099 VPWR.t610 VGND 0.07889f
C18100 VPWR.t1878 VGND 0.09265f
C18101 VPWR.t317 VGND 0.03348f
C18102 VPWR.t1879 VGND 0.02976f
C18103 VPWR.n787 VGND 0.09198f
C18104 VPWR.n788 VGND 0.01806f
C18105 VPWR.n789 VGND 0.00732f
C18106 VPWR.n790 VGND 0.10877f
C18107 VPWR.t1872 VGND 0.12017f
C18108 VPWR.t123 VGND 0.07889f
C18109 VPWR.t1757 VGND 0.09265f
C18110 VPWR.t1873 VGND 0.03348f
C18111 VPWR.t1758 VGND 0.02976f
C18112 VPWR.n791 VGND 0.09198f
C18113 VPWR.n792 VGND 0.01806f
C18114 VPWR.n793 VGND 0.00732f
C18115 VPWR.n794 VGND 0.10877f
C18116 VPWR.t959 VGND 0.12017f
C18117 VPWR.t124 VGND 0.07889f
C18118 VPWR.t8 VGND 0.09265f
C18119 VPWR.t960 VGND 0.03348f
C18120 VPWR.t9 VGND 0.02976f
C18121 VPWR.n795 VGND 0.09198f
C18122 VPWR.n796 VGND 0.01806f
C18123 VPWR.n797 VGND 0.00732f
C18124 VPWR.n798 VGND 0.10877f
C18125 VPWR.t2 VGND 0.12017f
C18126 VPWR.t1896 VGND 0.07889f
C18127 VPWR.t159 VGND 0.09265f
C18128 VPWR.t3 VGND 0.03348f
C18129 VPWR.t160 VGND 0.02976f
C18130 VPWR.n799 VGND 0.09198f
C18131 VPWR.n800 VGND 0.01806f
C18132 VPWR.n801 VGND 0.00732f
C18133 VPWR.n802 VGND 0.10877f
C18134 VPWR.t1699 VGND 0.12017f
C18135 VPWR.t126 VGND 0.07889f
C18136 VPWR.t177 VGND 0.09265f
C18137 VPWR.t1700 VGND 0.03348f
C18138 VPWR.t178 VGND 0.02976f
C18139 VPWR.n803 VGND 0.09198f
C18140 VPWR.n804 VGND 0.01806f
C18141 VPWR.n805 VGND 0.00732f
C18142 VPWR.n806 VGND 0.10877f
C18143 VPWR.t137 VGND 0.12017f
C18144 VPWR.t122 VGND 0.07889f
C18145 VPWR.t58 VGND 0.09265f
C18146 VPWR.t138 VGND 0.03348f
C18147 VPWR.t59 VGND 0.02976f
C18148 VPWR.n807 VGND 0.09198f
C18149 VPWR.n808 VGND 0.01806f
C18150 VPWR.n809 VGND 0.00732f
C18151 VPWR.n810 VGND 0.10877f
C18152 VPWR.t760 VGND 0.12017f
C18153 VPWR.t113 VGND 0.07889f
C18154 VPWR.t396 VGND 0.09265f
C18155 VPWR.t761 VGND 0.03348f
C18156 VPWR.t397 VGND 0.02976f
C18157 VPWR.n811 VGND 0.09198f
C18158 VPWR.n812 VGND 0.01806f
C18159 VPWR.n813 VGND 0.00732f
C18160 VPWR.n814 VGND 0.10877f
C18161 VPWR.t390 VGND 0.12017f
C18162 VPWR.t112 VGND 0.07889f
C18163 VPWR.t675 VGND 0.09265f
C18164 VPWR.t391 VGND 0.03348f
C18165 VPWR.t676 VGND 0.02976f
C18166 VPWR.n815 VGND 0.09198f
C18167 VPWR.n816 VGND 0.01806f
C18168 VPWR.n817 VGND 0.00732f
C18169 VPWR.n818 VGND 0.10877f
C18170 VPWR.t777 VGND 0.12017f
C18171 VPWR.t125 VGND 0.07889f
C18172 VPWR.t249 VGND 0.09265f
C18173 VPWR.t778 VGND 0.03348f
C18174 VPWR.t250 VGND 0.02976f
C18175 VPWR.n819 VGND 0.09198f
C18176 VPWR.n820 VGND 0.01806f
C18177 VPWR.n821 VGND 0.00732f
C18178 VPWR.n822 VGND 0.10877f
C18179 VPWR.t873 VGND 0.12017f
C18180 VPWR.t121 VGND 0.07889f
C18181 VPWR.t1052 VGND 0.09265f
C18182 VPWR.t874 VGND 0.03348f
C18183 VPWR.t1053 VGND 0.02976f
C18184 VPWR.n823 VGND 0.09198f
C18185 VPWR.n824 VGND 0.01806f
C18186 VPWR.n825 VGND 0.00732f
C18187 VPWR.n826 VGND 0.10877f
C18188 VPWR.t386 VGND 0.12017f
C18189 VPWR.t118 VGND 0.07889f
C18190 VPWR.t1064 VGND 0.09265f
C18191 VPWR.t387 VGND 0.03348f
C18192 VPWR.t1065 VGND 0.02976f
C18193 VPWR.n827 VGND 0.09198f
C18194 VPWR.n828 VGND 0.01806f
C18195 VPWR.n829 VGND 0.00732f
C18196 VPWR.n830 VGND 0.10877f
C18197 VPWR.t221 VGND 0.12017f
C18198 VPWR.t1894 VGND 0.07889f
C18199 VPWR.t1298 VGND 0.13401f
C18200 VPWR.n831 VGND 0.07657f
C18201 VPWR.n832 VGND 0.01806f
C18202 VPWR.n833 VGND 0.13984f
C18203 VPWR.n834 VGND 1.02091f
C18204 VPWR.n835 VGND 0.13984f
C18205 VPWR.t1718 VGND 0.03348f
C18206 VPWR.t1122 VGND 0.02976f
C18207 VPWR.n836 VGND 0.09198f
C18208 VPWR.t169 VGND 0.09265f
C18209 VPWR.t359 VGND 0.03348f
C18210 VPWR.t170 VGND 0.02976f
C18211 VPWR.n837 VGND 0.09198f
C18212 VPWR.n838 VGND 0.13984f
C18213 VPWR.n839 VGND 0.13984f
C18214 VPWR.t258 VGND 0.03348f
C18215 VPWR.t1546 VGND 0.02976f
C18216 VPWR.n840 VGND 0.09198f
C18217 VPWR.t1801 VGND 0.09265f
C18218 VPWR.t1599 VGND 0.03348f
C18219 VPWR.t1802 VGND 0.02976f
C18220 VPWR.n841 VGND 0.09198f
C18221 VPWR.n842 VGND 0.13984f
C18222 VPWR.n843 VGND 0.13984f
C18223 VPWR.t828 VGND 0.03348f
C18224 VPWR.t1738 VGND 0.02976f
C18225 VPWR.n844 VGND 0.09198f
C18226 VPWR.t833 VGND 0.09265f
C18227 VPWR.t1534 VGND 0.03348f
C18228 VPWR.t834 VGND 0.02976f
C18229 VPWR.n845 VGND 0.09198f
C18230 VPWR.n846 VGND 0.13984f
C18231 VPWR.n847 VGND 0.13984f
C18232 VPWR.t1818 VGND 0.03348f
C18233 VPWR.t1540 VGND 0.02976f
C18234 VPWR.n848 VGND 0.09198f
C18235 VPWR.t1823 VGND 0.09265f
C18236 VPWR.t419 VGND 0.03348f
C18237 VPWR.t1824 VGND 0.02976f
C18238 VPWR.n849 VGND 0.09198f
C18239 VPWR.n850 VGND 0.13984f
C18240 VPWR.n851 VGND 0.13984f
C18241 VPWR.t186 VGND 0.03348f
C18242 VPWR.t462 VGND 0.02976f
C18243 VPWR.n852 VGND 0.09198f
C18244 VPWR.t191 VGND 0.09265f
C18245 VPWR.t1680 VGND 0.03348f
C18246 VPWR.t192 VGND 0.02976f
C18247 VPWR.n853 VGND 0.09198f
C18248 VPWR.n854 VGND 0.13984f
C18249 VPWR.n855 VGND 0.13984f
C18250 VPWR.t295 VGND 0.03348f
C18251 VPWR.t802 VGND 0.02976f
C18252 VPWR.n856 VGND 0.09198f
C18253 VPWR.t79 VGND 0.09265f
C18254 VPWR.t1573 VGND 0.03348f
C18255 VPWR.t80 VGND 0.02976f
C18256 VPWR.n857 VGND 0.09198f
C18257 VPWR.n858 VGND 0.13984f
C18258 VPWR.n859 VGND 0.13984f
C18259 VPWR.t1508 VGND 0.03348f
C18260 VPWR.t1732 VGND 0.02976f
C18261 VPWR.n860 VGND 0.09198f
C18262 VPWR.t1481 VGND 0.09265f
C18263 VPWR.t725 VGND 0.03348f
C18264 VPWR.t1482 VGND 0.02976f
C18265 VPWR.n861 VGND 0.09198f
C18266 VPWR.n862 VGND 0.13984f
C18267 VPWR.n863 VGND 0.13984f
C18268 VPWR.t287 VGND 0.03348f
C18269 VPWR.t780 VGND 0.02976f
C18270 VPWR.n864 VGND 0.09198f
C18271 VPWR.t560 VGND 0.14585f
C18272 VPWR.t1907 VGND 0.07889f
C18273 VPWR.t917 VGND 0.09265f
C18274 VPWR.t561 VGND 0.03348f
C18275 VPWR.t918 VGND 0.02976f
C18276 VPWR.n865 VGND 0.09198f
C18277 VPWR.t575 VGND 0.03348f
C18278 VPWR.t628 VGND 0.02976f
C18279 VPWR.n866 VGND 0.09198f
C18280 VPWR.t574 VGND 0.14585f
C18281 VPWR.t956 VGND 0.07889f
C18282 VPWR.t627 VGND 0.09265f
C18283 VPWR.t220 VGND 0.03348f
C18284 VPWR.t1306 VGND 0.02976f
C18285 VPWR.n867 VGND 0.09198f
C18286 VPWR.n868 VGND 0.01806f
C18287 VPWR.n869 VGND 0.07657f
C18288 VPWR.t1305 VGND 0.13401f
C18289 VPWR.t952 VGND 0.07889f
C18290 VPWR.t219 VGND 0.12017f
C18291 VPWR.t385 VGND 0.03348f
C18292 VPWR.t1063 VGND 0.02976f
C18293 VPWR.n870 VGND 0.09198f
C18294 VPWR.n871 VGND 0.01806f
C18295 VPWR.n872 VGND 0.00732f
C18296 VPWR.n873 VGND 0.10877f
C18297 VPWR.t1062 VGND 0.09265f
C18298 VPWR.t929 VGND 0.07889f
C18299 VPWR.t384 VGND 0.12017f
C18300 VPWR.t870 VGND 0.03348f
C18301 VPWR.t1051 VGND 0.02976f
C18302 VPWR.n874 VGND 0.09198f
C18303 VPWR.n875 VGND 0.01806f
C18304 VPWR.n876 VGND 0.00732f
C18305 VPWR.n877 VGND 0.10877f
C18306 VPWR.t1050 VGND 0.09265f
C18307 VPWR.t1634 VGND 0.07889f
C18308 VPWR.t869 VGND 0.12017f
C18309 VPWR.t776 VGND 0.03348f
C18310 VPWR.t248 VGND 0.02976f
C18311 VPWR.n878 VGND 0.09198f
C18312 VPWR.n879 VGND 0.01806f
C18313 VPWR.n880 VGND 0.00732f
C18314 VPWR.n881 VGND 0.10877f
C18315 VPWR.t247 VGND 0.09265f
C18316 VPWR.t1635 VGND 0.07889f
C18317 VPWR.t775 VGND 0.12017f
C18318 VPWR.t389 VGND 0.03348f
C18319 VPWR.t674 VGND 0.02976f
C18320 VPWR.n882 VGND 0.09198f
C18321 VPWR.n883 VGND 0.01806f
C18322 VPWR.n884 VGND 0.00732f
C18323 VPWR.n885 VGND 0.10877f
C18324 VPWR.t673 VGND 0.09265f
C18325 VPWR.t925 VGND 0.07889f
C18326 VPWR.t388 VGND 0.12017f
C18327 VPWR.t759 VGND 0.03348f
C18328 VPWR.t395 VGND 0.02976f
C18329 VPWR.n886 VGND 0.09198f
C18330 VPWR.n887 VGND 0.01806f
C18331 VPWR.n888 VGND 0.00732f
C18332 VPWR.n889 VGND 0.10877f
C18333 VPWR.t394 VGND 0.09265f
C18334 VPWR.t926 VGND 0.07889f
C18335 VPWR.t758 VGND 0.12017f
C18336 VPWR.t136 VGND 0.03348f
C18337 VPWR.t767 VGND 0.02976f
C18338 VPWR.n890 VGND 0.09198f
C18339 VPWR.n891 VGND 0.01806f
C18340 VPWR.n892 VGND 0.00732f
C18341 VPWR.n893 VGND 0.10877f
C18342 VPWR.t766 VGND 0.09265f
C18343 VPWR.t1638 VGND 0.07889f
C18344 VPWR.t135 VGND 0.12017f
C18345 VPWR.t1859 VGND 0.03348f
C18346 VPWR.t142 VGND 0.02976f
C18347 VPWR.n894 VGND 0.09198f
C18348 VPWR.n895 VGND 0.01806f
C18349 VPWR.n896 VGND 0.00732f
C18350 VPWR.n897 VGND 0.10877f
C18351 VPWR.t141 VGND 0.09265f
C18352 VPWR.t953 VGND 0.07889f
C18353 VPWR.t1858 VGND 0.12017f
C18354 VPWR.t1 VGND 0.03348f
C18355 VPWR.t158 VGND 0.02976f
C18356 VPWR.n898 VGND 0.09198f
C18357 VPWR.n899 VGND 0.01806f
C18358 VPWR.n900 VGND 0.00732f
C18359 VPWR.n901 VGND 0.10877f
C18360 VPWR.t157 VGND 0.09265f
C18361 VPWR.t954 VGND 0.07889f
C18362 VPWR.t0 VGND 0.12017f
C18363 VPWR.t958 VGND 0.03348f
C18364 VPWR.t7 VGND 0.02976f
C18365 VPWR.n902 VGND 0.09198f
C18366 VPWR.n903 VGND 0.01806f
C18367 VPWR.n904 VGND 0.00732f
C18368 VPWR.n905 VGND 0.10877f
C18369 VPWR.t6 VGND 0.09265f
C18370 VPWR.t1636 VGND 0.07889f
C18371 VPWR.t957 VGND 0.12017f
C18372 VPWR.t1871 VGND 0.03348f
C18373 VPWR.t1756 VGND 0.02976f
C18374 VPWR.n906 VGND 0.09198f
C18375 VPWR.n907 VGND 0.01806f
C18376 VPWR.n908 VGND 0.00732f
C18377 VPWR.n909 VGND 0.10877f
C18378 VPWR.t1755 VGND 0.09265f
C18379 VPWR.t1637 VGND 0.07889f
C18380 VPWR.t1870 VGND 0.12017f
C18381 VPWR.t315 VGND 0.03348f
C18382 VPWR.t1877 VGND 0.02976f
C18383 VPWR.n910 VGND 0.09198f
C18384 VPWR.n911 VGND 0.01806f
C18385 VPWR.n912 VGND 0.00732f
C18386 VPWR.n913 VGND 0.10877f
C18387 VPWR.t1876 VGND 0.09265f
C18388 VPWR.t955 VGND 0.07889f
C18389 VPWR.t314 VGND 0.12017f
C18390 VPWR.t1478 VGND 0.03348f
C18391 VPWR.t1808 VGND 0.02976f
C18392 VPWR.n914 VGND 0.09198f
C18393 VPWR.n915 VGND 0.01806f
C18394 VPWR.n916 VGND 0.00732f
C18395 VPWR.n917 VGND 0.10877f
C18396 VPWR.t1807 VGND 0.09265f
C18397 VPWR.t927 VGND 0.07889f
C18398 VPWR.t1477 VGND 0.12017f
C18399 VPWR.t678 VGND 0.03348f
C18400 VPWR.t1514 VGND 0.02976f
C18401 VPWR.n918 VGND 0.09198f
C18402 VPWR.n919 VGND 0.01806f
C18403 VPWR.n920 VGND 0.00732f
C18404 VPWR.n921 VGND 0.10877f
C18405 VPWR.t1513 VGND 0.09265f
C18406 VPWR.t928 VGND 0.07889f
C18407 VPWR.t677 VGND 0.12017f
C18408 VPWR.t1554 VGND 0.03348f
C18409 VPWR.t1581 VGND 0.02976f
C18410 VPWR.n922 VGND 0.09198f
C18411 VPWR.n923 VGND 0.01806f
C18412 VPWR.n924 VGND 0.00732f
C18413 VPWR.n925 VGND 0.10877f
C18414 VPWR.t1580 VGND 0.09265f
C18415 VPWR.t1639 VGND 0.07889f
C18416 VPWR.t1553 VGND 0.12017f
C18417 VPWR.n926 VGND 0.10877f
C18418 VPWR.n927 VGND 0.00732f
C18419 VPWR.n928 VGND 0.01806f
C18420 VPWR.n929 VGND 0.13984f
C18421 VPWR.n930 VGND 1.01451f
C18422 VPWR.n931 VGND 0.13984f
C18423 VPWR.t569 VGND 0.03348f
C18424 VPWR.t1750 VGND 0.02976f
C18425 VPWR.n932 VGND 0.09198f
C18426 VPWR.t568 VGND 0.14585f
C18427 VPWR.t908 VGND 0.07889f
C18428 VPWR.t1749 VGND 0.09265f
C18429 VPWR.t697 VGND 0.12017f
C18430 VPWR.t436 VGND 0.03348f
C18431 VPWR.t706 VGND 0.02976f
C18432 VPWR.n933 VGND 0.09198f
C18433 VPWR.n934 VGND 0.13984f
C18434 VPWR.n935 VGND 0.13984f
C18435 VPWR.t698 VGND 0.03348f
C18436 VPWR.t1466 VGND 0.02976f
C18437 VPWR.n936 VGND 0.09198f
C18438 VPWR.t1031 VGND 0.07889f
C18439 VPWR.t1465 VGND 0.09265f
C18440 VPWR.t1723 VGND 0.12017f
C18441 VPWR.t1490 VGND 0.03348f
C18442 VPWR.t319 VGND 0.02976f
C18443 VPWR.n937 VGND 0.09198f
C18444 VPWR.n938 VGND 0.13984f
C18445 VPWR.n939 VGND 0.13984f
C18446 VPWR.t1724 VGND 0.03348f
C18447 VPWR.t753 VGND 0.02976f
C18448 VPWR.n940 VGND 0.09198f
C18449 VPWR.t907 VGND 0.07889f
C18450 VPWR.t752 VGND 0.09265f
C18451 VPWR.t789 VGND 0.12017f
C18452 VPWR.t979 VGND 0.03348f
C18453 VPWR.t806 VGND 0.02976f
C18454 VPWR.n941 VGND 0.09198f
C18455 VPWR.n942 VGND 0.13984f
C18456 VPWR.n943 VGND 0.13984f
C18457 VPWR.t790 VGND 0.03348f
C18458 VPWR.t276 VGND 0.02976f
C18459 VPWR.n944 VGND 0.09198f
C18460 VPWR.t860 VGND 0.07889f
C18461 VPWR.t275 VGND 0.09265f
C18462 VPWR.t1852 VGND 0.12017f
C18463 VPWR.t268 VGND 0.03348f
C18464 VPWR.t1706 VGND 0.02976f
C18465 VPWR.n945 VGND 0.09198f
C18466 VPWR.n946 VGND 0.13984f
C18467 VPWR.n947 VGND 0.13984f
C18468 VPWR.t1853 VGND 0.03348f
C18469 VPWR.t664 VGND 0.02976f
C18470 VPWR.n948 VGND 0.09198f
C18471 VPWR.t905 VGND 0.07889f
C18472 VPWR.t663 VGND 0.09265f
C18473 VPWR.t332 VGND 0.12017f
C18474 VPWR.t456 VGND 0.03348f
C18475 VPWR.t534 VGND 0.02976f
C18476 VPWR.n949 VGND 0.09198f
C18477 VPWR.n950 VGND 0.13984f
C18478 VPWR.n951 VGND 0.13984f
C18479 VPWR.t333 VGND 0.03348f
C18480 VPWR.t1631 VGND 0.02976f
C18481 VPWR.n952 VGND 0.09198f
C18482 VPWR.t1029 VGND 0.07889f
C18483 VPWR.t1630 VGND 0.09265f
C18484 VPWR.t887 VGND 0.12017f
C18485 VPWR.t1623 VGND 0.03348f
C18486 VPWR.t898 VGND 0.02976f
C18487 VPWR.n953 VGND 0.09198f
C18488 VPWR.n954 VGND 0.13984f
C18489 VPWR.n955 VGND 0.13984f
C18490 VPWR.t888 VGND 0.03348f
C18491 VPWR.t880 VGND 0.02976f
C18492 VPWR.n956 VGND 0.09198f
C18493 VPWR.t859 VGND 0.07889f
C18494 VPWR.t879 VGND 0.09265f
C18495 VPWR.t635 VGND 0.12017f
C18496 VPWR.t1794 VGND 0.03348f
C18497 VPWR.t1047 VGND 0.02976f
C18498 VPWR.n957 VGND 0.09198f
C18499 VPWR.n958 VGND 0.13984f
C18500 VPWR.n959 VGND 0.13984f
C18501 VPWR.t636 VGND 0.03348f
C18502 VPWR.t224 VGND 0.02976f
C18503 VPWR.n960 VGND 0.09198f
C18504 VPWR.t857 VGND 0.07889f
C18505 VPWR.t223 VGND 0.09265f
C18506 VPWR.t29 VGND 0.03348f
C18507 VPWR.t1414 VGND 0.02976f
C18508 VPWR.n961 VGND 0.09198f
C18509 VPWR.t232 VGND 0.03348f
C18510 VPWR.t1266 VGND 0.02976f
C18511 VPWR.n962 VGND 0.09198f
C18512 VPWR.t580 VGND 0.14585f
C18513 VPWR.t1025 VGND 0.07889f
C18514 VPWR.t1844 VGND 0.09265f
C18515 VPWR.t581 VGND 0.03348f
C18516 VPWR.t1845 VGND 0.02976f
C18517 VPWR.n963 VGND 0.09198f
C18518 VPWR.n964 VGND 0.01806f
C18519 VPWR.n965 VGND 0.00732f
C18520 VPWR.n966 VGND 0.10877f
C18521 VPWR.t625 VGND 0.12017f
C18522 VPWR.t1588 VGND 0.07889f
C18523 VPWR.t909 VGND 0.09265f
C18524 VPWR.t626 VGND 0.03348f
C18525 VPWR.t910 VGND 0.02976f
C18526 VPWR.n967 VGND 0.09198f
C18527 VPWR.n968 VGND 0.01806f
C18528 VPWR.n969 VGND 0.00732f
C18529 VPWR.n970 VGND 0.10877f
C18530 VPWR.t1584 VGND 0.12017f
C18531 VPWR.t1664 VGND 0.07889f
C18532 VPWR.t1503 VGND 0.09265f
C18533 VPWR.t1585 VGND 0.03348f
C18534 VPWR.t1504 VGND 0.02976f
C18535 VPWR.n971 VGND 0.09198f
C18536 VPWR.n972 VGND 0.01806f
C18537 VPWR.n973 VGND 0.00732f
C18538 VPWR.n974 VGND 0.10877f
C18539 VPWR.t1467 VGND 0.12017f
C18540 VPWR.t1663 VGND 0.07889f
C18541 VPWR.t1813 VGND 0.09265f
C18542 VPWR.t1468 VGND 0.03348f
C18543 VPWR.t1814 VGND 0.02976f
C18544 VPWR.n975 VGND 0.09198f
C18545 VPWR.n976 VGND 0.01806f
C18546 VPWR.n977 VGND 0.00732f
C18547 VPWR.n978 VGND 0.10877f
C18548 VPWR.t326 VGND 0.12017f
C18549 VPWR.t601 VGND 0.07889f
C18550 VPWR.t744 VGND 0.09265f
C18551 VPWR.t327 VGND 0.03348f
C18552 VPWR.t745 VGND 0.02976f
C18553 VPWR.n979 VGND 0.09198f
C18554 VPWR.n980 VGND 0.01806f
C18555 VPWR.n981 VGND 0.00732f
C18556 VPWR.n982 VGND 0.10877f
C18557 VPWR.t740 VGND 0.12017f
C18558 VPWR.t424 VGND 0.07889f
C18559 VPWR.t1763 VGND 0.09265f
C18560 VPWR.t741 VGND 0.03348f
C18561 VPWR.t1764 VGND 0.02976f
C18562 VPWR.n983 VGND 0.09198f
C18563 VPWR.n984 VGND 0.01806f
C18564 VPWR.n985 VGND 0.00732f
C18565 VPWR.n986 VGND 0.10877f
C18566 VPWR.t1759 VGND 0.12017f
C18567 VPWR.t423 VGND 0.07889f
C18568 VPWR.t14 VGND 0.09265f
C18569 VPWR.t1760 VGND 0.03348f
C18570 VPWR.t15 VGND 0.02976f
C18571 VPWR.n987 VGND 0.09198f
C18572 VPWR.n988 VGND 0.01806f
C18573 VPWR.n989 VGND 0.00732f
C18574 VPWR.n990 VGND 0.10877f
C18575 VPWR.t10 VGND 0.12017f
C18576 VPWR.t600 VGND 0.07889f
C18577 VPWR.t163 VGND 0.09265f
C18578 VPWR.t11 VGND 0.03348f
C18579 VPWR.t164 VGND 0.02976f
C18580 VPWR.n991 VGND 0.09198f
C18581 VPWR.n992 VGND 0.01806f
C18582 VPWR.n993 VGND 0.00732f
C18583 VPWR.n994 VGND 0.10877f
C18584 VPWR.t1707 VGND 0.12017f
C18585 VPWR.t1590 VGND 0.07889f
C18586 VPWR.t183 VGND 0.09265f
C18587 VPWR.t1708 VGND 0.03348f
C18588 VPWR.t184 VGND 0.02976f
C18589 VPWR.n995 VGND 0.09198f
C18590 VPWR.n996 VGND 0.01806f
C18591 VPWR.n997 VGND 0.00732f
C18592 VPWR.n998 VGND 0.10877f
C18593 VPWR.t179 VGND 0.12017f
C18594 VPWR.t425 VGND 0.07889f
C18595 VPWR.t66 VGND 0.09265f
C18596 VPWR.t180 VGND 0.03348f
C18597 VPWR.t67 VGND 0.02976f
C18598 VPWR.n999 VGND 0.09198f
C18599 VPWR.n1000 VGND 0.01806f
C18600 VPWR.n1001 VGND 0.00732f
C18601 VPWR.n1002 VGND 0.10877f
C18602 VPWR.t764 VGND 0.12017f
C18603 VPWR.t1027 VGND 0.07889f
C18604 VPWR.t594 VGND 0.09265f
C18605 VPWR.t765 VGND 0.03348f
C18606 VPWR.t595 VGND 0.02976f
C18607 VPWR.n1003 VGND 0.09198f
C18608 VPWR.n1004 VGND 0.01806f
C18609 VPWR.n1005 VGND 0.00732f
C18610 VPWR.n1006 VGND 0.10877f
C18611 VPWR.t590 VGND 0.12017f
C18612 VPWR.t1026 VGND 0.07889f
C18613 VPWR.t1009 VGND 0.09265f
C18614 VPWR.t591 VGND 0.03348f
C18615 VPWR.t1010 VGND 0.02976f
C18616 VPWR.n1007 VGND 0.09198f
C18617 VPWR.n1008 VGND 0.01806f
C18618 VPWR.n1009 VGND 0.00732f
C18619 VPWR.n1010 VGND 0.10877f
C18620 VPWR.t671 VGND 0.12017f
C18621 VPWR.t422 VGND 0.07889f
C18622 VPWR.t253 VGND 0.09265f
C18623 VPWR.t672 VGND 0.03348f
C18624 VPWR.t254 VGND 0.02976f
C18625 VPWR.n1011 VGND 0.09198f
C18626 VPWR.n1012 VGND 0.01806f
C18627 VPWR.n1013 VGND 0.00732f
C18628 VPWR.n1014 VGND 0.10877f
C18629 VPWR.t88 VGND 0.12017f
C18630 VPWR.t1666 VGND 0.07889f
C18631 VPWR.t1551 VGND 0.09265f
C18632 VPWR.t89 VGND 0.03348f
C18633 VPWR.t1552 VGND 0.02976f
C18634 VPWR.n1015 VGND 0.09198f
C18635 VPWR.n1016 VGND 0.01806f
C18636 VPWR.n1017 VGND 0.00732f
C18637 VPWR.n1018 VGND 0.10877f
C18638 VPWR.t641 VGND 0.12017f
C18639 VPWR.t1665 VGND 0.07889f
C18640 VPWR.t1713 VGND 0.09265f
C18641 VPWR.t642 VGND 0.03348f
C18642 VPWR.t1714 VGND 0.02976f
C18643 VPWR.n1019 VGND 0.09198f
C18644 VPWR.n1020 VGND 0.01806f
C18645 VPWR.n1021 VGND 0.00732f
C18646 VPWR.n1022 VGND 0.10877f
C18647 VPWR.t231 VGND 0.12017f
C18648 VPWR.t1589 VGND 0.07889f
C18649 VPWR.t1265 VGND 0.13401f
C18650 VPWR.n1023 VGND 0.07657f
C18651 VPWR.n1024 VGND 0.01806f
C18652 VPWR.n1025 VGND 0.13984f
C18653 VPWR.n1026 VGND 5.87665f
C18654 VPWR.n1027 VGND 0.066f
C18655 VPWR.n1028 VGND -0.01875f
C18656 VPWR.t2061 VGND 0.01122f
C18657 VPWR.t1267 VGND 0.01228f
C18658 VPWR.n1029 VGND 0.03058f
C18659 VPWR.n1030 VGND 0.00584f
C18660 VPWR.t1269 VGND 0.02693f
C18661 VPWR.n1031 VGND 0.05753f
C18662 VPWR.t1377 VGND 0.02976f
C18663 VPWR.n1032 VGND 0.04716f
C18664 VPWR.t233 VGND 0.09265f
C18665 VPWR.t1957 VGND 0.01122f
C18666 VPWR.t1159 VGND 0.01228f
C18667 VPWR.n1033 VGND 0.03058f
C18668 VPWR.n1034 VGND 0.00584f
C18669 VPWR.t1161 VGND 0.02693f
C18670 VPWR.n1035 VGND 0.05753f
C18671 VPWR.t234 VGND 0.02976f
C18672 VPWR.n1036 VGND 0.04716f
C18673 VPWR.n1037 VGND -0.01875f
C18674 VPWR.n1038 VGND 0.066f
C18675 VPWR.t2065 VGND 0.01141f
C18676 VPWR.t1118 VGND 0.01247f
C18677 VPWR.n1039 VGND 0.02783f
C18678 VPWR.n1040 VGND 0.01907f
C18679 VPWR.n1041 VGND 0.06276f
C18680 VPWR.n1042 VGND 0.09795f
C18681 VPWR.n1043 VGND 0.05468f
C18682 VPWR.n1044 VGND 0.066f
C18683 VPWR.n1045 VGND -0.01875f
C18684 VPWR.t1967 VGND 0.01122f
C18685 VPWR.t1245 VGND 0.01228f
C18686 VPWR.n1046 VGND 0.03058f
C18687 VPWR.n1047 VGND 0.00584f
C18688 VPWR.t1247 VGND 0.02693f
C18689 VPWR.n1048 VGND 0.05753f
C18690 VPWR.t996 VGND 0.02976f
C18691 VPWR.n1049 VGND 0.04716f
C18692 VPWR.t995 VGND 0.09265f
C18693 VPWR.t1110 VGND 0.12017f
C18694 VPWR.t2055 VGND 0.01122f
C18695 VPWR.t1286 VGND 0.01228f
C18696 VPWR.n1050 VGND 0.03058f
C18697 VPWR.n1051 VGND 0.00584f
C18698 VPWR.t1288 VGND 0.02693f
C18699 VPWR.n1052 VGND 0.05753f
C18700 VPWR.t95 VGND 0.02976f
C18701 VPWR.n1053 VGND 0.04716f
C18702 VPWR.n1054 VGND 0.00809f
C18703 VPWR.n1055 VGND 0.19469f
C18704 VPWR.n1056 VGND 0.08393f
C18705 VPWR.n1057 VGND 0.03454f
C18706 VPWR.t1341 VGND 0.03348f
C18707 VPWR.t1333 VGND 0.02976f
C18708 VPWR.n1058 VGND 0.09198f
C18709 VPWR.t1332 VGND 0.09265f
C18710 VPWR.t1084 VGND 0.12017f
C18711 VPWR.t1369 VGND 0.03348f
C18712 VPWR.t1361 VGND 0.02976f
C18713 VPWR.n1059 VGND 0.09198f
C18714 VPWR.n1060 VGND 0.00809f
C18715 VPWR.t1085 VGND 0.03348f
C18716 VPWR.t1212 VGND 0.02976f
C18717 VPWR.n1061 VGND 0.09198f
C18718 VPWR.t1087 VGND 0.07889f
C18719 VPWR.t1211 VGND 0.13401f
C18720 VPWR.n1062 VGND 0.07653f
C18721 VPWR.n1063 VGND 0.01707f
C18722 VPWR.t2034 VGND 0.01125f
C18723 VPWR.t1210 VGND 0.01232f
C18724 VPWR.n1064 VGND 0.03008f
C18725 VPWR.n1065 VGND 0.03301f
C18726 VPWR.n1066 VGND 0.00701f
C18727 VPWR.n1067 VGND 0.01831f
C18728 VPWR.n1068 VGND 0.17674f
C18729 VPWR.t1989 VGND 0.01125f
C18730 VPWR.t1331 VGND 0.01232f
C18731 VPWR.n1069 VGND 0.03008f
C18732 VPWR.n1070 VGND 0.03301f
C18733 VPWR.n1071 VGND 0.01723f
C18734 VPWR.n1072 VGND 0.00701f
C18735 VPWR.n1073 VGND 0.00809f
C18736 VPWR.n1074 VGND 0.01723f
C18737 VPWR.n1075 VGND 0.00701f
C18738 VPWR.t1988 VGND 0.01141f
C18739 VPWR.t1337 VGND 0.01247f
C18740 VPWR.n1076 VGND 0.02782f
C18741 VPWR.n1077 VGND 0.02832f
C18742 VPWR.n1078 VGND 0.01831f
C18743 VPWR.n1079 VGND 0.17674f
C18744 VPWR.t1947 VGND 0.01125f
C18745 VPWR.t1439 VGND 0.01232f
C18746 VPWR.n1080 VGND 0.03008f
C18747 VPWR.n1081 VGND 0.03301f
C18748 VPWR.n1082 VGND 0.01723f
C18749 VPWR.n1083 VGND 0.00701f
C18750 VPWR.n1084 VGND 0.01723f
C18751 VPWR.n1085 VGND 0.00701f
C18752 VPWR.t1945 VGND 0.01141f
C18753 VPWR.t1445 VGND 0.01247f
C18754 VPWR.n1086 VGND 0.02782f
C18755 VPWR.n1087 VGND 0.02832f
C18756 VPWR.n1088 VGND 0.01831f
C18757 VPWR.n1089 VGND 0.17674f
C18758 VPWR.t1949 VGND 0.01125f
C18759 VPWR.t1431 VGND 0.01232f
C18760 VPWR.n1090 VGND 0.03008f
C18761 VPWR.n1091 VGND 0.03301f
C18762 VPWR.n1092 VGND 0.01723f
C18763 VPWR.n1093 VGND 0.00701f
C18764 VPWR.n1094 VGND 0.01723f
C18765 VPWR.n1095 VGND 0.00701f
C18766 VPWR.t2049 VGND 0.01141f
C18767 VPWR.t1164 VGND 0.01247f
C18768 VPWR.n1096 VGND 0.02782f
C18769 VPWR.n1097 VGND 0.02832f
C18770 VPWR.n1098 VGND 0.01831f
C18771 VPWR.n1099 VGND 0.17674f
C18772 VPWR.t2059 VGND 0.01125f
C18773 VPWR.t1136 VGND 0.01232f
C18774 VPWR.n1100 VGND 0.03008f
C18775 VPWR.n1101 VGND 0.03301f
C18776 VPWR.n1102 VGND 0.01723f
C18777 VPWR.n1103 VGND 0.00701f
C18778 VPWR.n1104 VGND 0.01723f
C18779 VPWR.n1105 VGND 0.00701f
C18780 VPWR.t2014 VGND 0.01141f
C18781 VPWR.t1248 VGND 0.01247f
C18782 VPWR.n1106 VGND 0.02782f
C18783 VPWR.n1107 VGND 0.02832f
C18784 VPWR.n1108 VGND 0.01831f
C18785 VPWR.n1109 VGND 0.02668f
C18786 VPWR.t2018 VGND 0.01125f
C18787 VPWR.t1242 VGND 0.01232f
C18788 VPWR.n1110 VGND 0.03008f
C18789 VPWR.n1111 VGND 0.03301f
C18790 VPWR.n1112 VGND 0.01831f
C18791 VPWR.n1113 VGND 0.00701f
C18792 VPWR.t2012 VGND 0.01122f
C18793 VPWR.t1388 VGND 0.01228f
C18794 VPWR.n1114 VGND 0.03131f
C18795 VPWR.n1115 VGND 0.01979f
C18796 VPWR.t1969 VGND 0.01141f
C18797 VPWR.t1378 VGND 0.01247f
C18798 VPWR.n1116 VGND 0.02782f
C18799 VPWR.n1117 VGND 0.02832f
C18800 VPWR.n1118 VGND 0.01785f
C18801 VPWR.t2067 VGND 0.01125f
C18802 VPWR.t1106 VGND 0.01232f
C18803 VPWR.n1119 VGND 0.03008f
C18804 VPWR.n1120 VGND 0.03301f
C18805 VPWR.n1121 VGND 0.00809f
C18806 VPWR.t1390 VGND 0.03348f
C18807 VPWR.t1108 VGND 0.02976f
C18808 VPWR.n1122 VGND 0.09198f
C18809 VPWR.t1389 VGND 0.14585f
C18810 VPWR.t1379 VGND 0.07889f
C18811 VPWR.t1107 VGND 0.09265f
C18812 VPWR.t1262 VGND 0.12017f
C18813 VPWR.t1158 VGND 0.03348f
C18814 VPWR.t1244 VGND 0.02976f
C18815 VPWR.n1123 VGND 0.09198f
C18816 VPWR.n1124 VGND 0.00837f
C18817 VPWR.t2062 VGND 0.01122f
C18818 VPWR.t1261 VGND 0.01228f
C18819 VPWR.n1125 VGND 0.03131f
C18820 VPWR.n1126 VGND 0.03712f
C18821 VPWR.n1127 VGND 0.03454f
C18822 VPWR.n1128 VGND 0.13984f
C18823 VPWR.n1129 VGND 0.00809f
C18824 VPWR.n1130 VGND 0.01806f
C18825 VPWR.n1131 VGND 0.066f
C18826 VPWR.n1132 VGND 0.05468f
C18827 VPWR.t1950 VGND 0.01141f
C18828 VPWR.t1429 VGND 0.01247f
C18829 VPWR.n1133 VGND 0.02783f
C18830 VPWR.n1134 VGND 0.01907f
C18831 VPWR.n1135 VGND 0.06276f
C18832 VPWR.n1136 VGND 0.09795f
C18833 VPWR.n1137 VGND 0.066f
C18834 VPWR.n1138 VGND 0.066f
C18835 VPWR.n1139 VGND 0.066f
C18836 VPWR.n1140 VGND 0.066f
C18837 VPWR.n1141 VGND 0.066f
C18838 VPWR.n1142 VGND 0.066f
C18839 VPWR.n1143 VGND 0.05468f
C18840 VPWR.n1144 VGND 0.00809f
C18841 VPWR.n1145 VGND -0.01875f
C18842 VPWR.t2020 VGND 0.01122f
C18843 VPWR.t1372 VGND 0.01228f
C18844 VPWR.n1146 VGND 0.03058f
C18845 VPWR.n1147 VGND 0.00584f
C18846 VPWR.t1374 VGND 0.02693f
C18847 VPWR.n1148 VGND 0.05753f
C18848 VPWR.t540 VGND 0.02976f
C18849 VPWR.n1149 VGND 0.04716f
C18850 VPWR.t539 VGND 0.09265f
C18851 VPWR.t1119 VGND 0.07889f
C18852 VPWR.t1246 VGND 0.12017f
C18853 VPWR.t1975 VGND 0.01122f
C18854 VPWR.t1115 VGND 0.01228f
C18855 VPWR.n1150 VGND 0.03058f
C18856 VPWR.n1151 VGND 0.00584f
C18857 VPWR.t1117 VGND 0.02693f
C18858 VPWR.n1152 VGND 0.05753f
C18859 VPWR.t771 VGND 0.02976f
C18860 VPWR.n1153 VGND 0.04716f
C18861 VPWR.n1154 VGND 0.00809f
C18862 VPWR.n1155 VGND 0.00809f
C18863 VPWR.t1927 VGND 0.01122f
C18864 VPWR.t1356 VGND 0.01228f
C18865 VPWR.n1156 VGND 0.03058f
C18866 VPWR.n1157 VGND 0.00584f
C18867 VPWR.t1358 VGND 0.02693f
C18868 VPWR.n1158 VGND 0.05753f
C18869 VPWR.t1069 VGND 0.02976f
C18870 VPWR.n1159 VGND 0.04716f
C18871 VPWR.t201 VGND 0.09265f
C18872 VPWR.t1938 VGND 0.01122f
C18873 VPWR.t1215 VGND 0.01228f
C18874 VPWR.n1160 VGND 0.03058f
C18875 VPWR.n1161 VGND 0.00584f
C18876 VPWR.t1217 VGND 0.02693f
C18877 VPWR.n1162 VGND 0.05753f
C18878 VPWR.t202 VGND 0.02976f
C18879 VPWR.n1163 VGND 0.04716f
C18880 VPWR.n1164 VGND 0.00809f
C18881 VPWR.n1165 VGND 0.00809f
C18882 VPWR.t2023 VGND 0.01122f
C18883 VPWR.t1093 VGND 0.01228f
C18884 VPWR.n1166 VGND 0.03058f
C18885 VPWR.n1167 VGND 0.00584f
C18886 VPWR.t1095 VGND 0.02693f
C18887 VPWR.n1168 VGND 0.05753f
C18888 VPWR.t282 VGND 0.02976f
C18889 VPWR.n1169 VGND 0.04716f
C18890 VPWR.t811 VGND 0.09265f
C18891 VPWR.t2035 VGND 0.01122f
C18892 VPWR.t1342 VGND 0.01228f
C18893 VPWR.n1170 VGND 0.03058f
C18894 VPWR.n1171 VGND 0.00584f
C18895 VPWR.t1344 VGND 0.02693f
C18896 VPWR.n1172 VGND 0.05753f
C18897 VPWR.t812 VGND 0.02976f
C18898 VPWR.n1173 VGND 0.04716f
C18899 VPWR.n1174 VGND 0.00809f
C18900 VPWR.n1175 VGND 0.00837f
C18901 VPWR.t1958 VGND 0.01122f
C18902 VPWR.t1153 VGND 0.01228f
C18903 VPWR.n1176 VGND 0.03131f
C18904 VPWR.n1177 VGND 0.03712f
C18905 VPWR.n1178 VGND 0.03454f
C18906 VPWR.t1143 VGND 0.03348f
C18907 VPWR.t1138 VGND 0.02976f
C18908 VPWR.n1179 VGND 0.09198f
C18909 VPWR.t1249 VGND 0.07889f
C18910 VPWR.t1256 VGND 0.09265f
C18911 VPWR.t1263 VGND 0.03348f
C18912 VPWR.t1257 VGND 0.02976f
C18913 VPWR.n1180 VGND 0.09198f
C18914 VPWR.n1181 VGND 0.00728f
C18915 VPWR.n1182 VGND 0.10877f
C18916 VPWR.t1424 VGND 0.12017f
C18917 VPWR.t1290 VGND 0.07889f
C18918 VPWR.t1416 VGND 0.09265f
C18919 VPWR.t1425 VGND 0.03348f
C18920 VPWR.t1417 VGND 0.02976f
C18921 VPWR.n1183 VGND 0.09198f
C18922 VPWR.n1184 VGND 0.00728f
C18923 VPWR.n1185 VGND 0.10877f
C18924 VPWR.t1142 VGND 0.12017f
C18925 VPWR.t1398 VGND 0.07889f
C18926 VPWR.t1137 VGND 0.09265f
C18927 VPWR.t1214 VGND 0.07889f
C18928 VPWR.t1340 VGND 0.12017f
C18929 VPWR.t1103 VGND 0.03348f
C18930 VPWR.t1204 VGND 0.02976f
C18931 VPWR.n1186 VGND 0.09198f
C18932 VPWR.n1187 VGND 0.00728f
C18933 VPWR.n1188 VGND 0.10877f
C18934 VPWR.t1203 VGND 0.09265f
C18935 VPWR.t1188 VGND 0.07889f
C18936 VPWR.t1102 VGND 0.12017f
C18937 VPWR.t1082 VGND 0.03348f
C18938 VPWR.t1460 VGND 0.02976f
C18939 VPWR.n1189 VGND 0.09198f
C18940 VPWR.n1190 VGND 0.00728f
C18941 VPWR.n1191 VGND 0.10877f
C18942 VPWR.t1459 VGND 0.09265f
C18943 VPWR.t1338 VGND 0.07889f
C18944 VPWR.t1081 VGND 0.12017f
C18945 VPWR.t1336 VGND 0.03348f
C18946 VPWR.t1441 VGND 0.02976f
C18947 VPWR.n1192 VGND 0.09198f
C18948 VPWR.n1193 VGND 0.00837f
C18949 VPWR.t2031 VGND 0.01122f
C18950 VPWR.t1080 VGND 0.01228f
C18951 VPWR.n1194 VGND 0.03131f
C18952 VPWR.n1195 VGND 0.03712f
C18953 VPWR.n1196 VGND 0.03454f
C18954 VPWR.n1197 VGND 0.01723f
C18955 VPWR.n1198 VGND 0.00728f
C18956 VPWR.n1199 VGND 0.10877f
C18957 VPWR.t1440 VGND 0.09265f
C18958 VPWR.t1316 VGND 0.07889f
C18959 VPWR.t1335 VGND 0.12017f
C18960 VPWR.t1209 VGND 0.03348f
C18961 VPWR.t1282 VGND 0.02976f
C18962 VPWR.n1200 VGND 0.09198f
C18963 VPWR.n1201 VGND 0.00728f
C18964 VPWR.n1202 VGND 0.10877f
C18965 VPWR.t1281 VGND 0.09265f
C18966 VPWR.t1163 VGND 0.07889f
C18967 VPWR.t1208 VGND 0.12017f
C18968 VPWR.t1183 VGND 0.03348f
C18969 VPWR.t1178 VGND 0.02976f
C18970 VPWR.n1203 VGND 0.09198f
C18971 VPWR.n1204 VGND 0.00728f
C18972 VPWR.n1205 VGND 0.10877f
C18973 VPWR.t1177 VGND 0.09265f
C18974 VPWR.t1446 VGND 0.07889f
C18975 VPWR.t1182 VGND 0.12017f
C18976 VPWR.t1422 VGND 0.03348f
C18977 VPWR.t1433 VGND 0.02976f
C18978 VPWR.n1206 VGND 0.09198f
C18979 VPWR.n1207 VGND 0.00837f
C18980 VPWR.t1992 VGND 0.01122f
C18981 VPWR.t1181 VGND 0.01228f
C18982 VPWR.n1208 VGND 0.03131f
C18983 VPWR.n1209 VGND 0.03712f
C18984 VPWR.n1210 VGND 0.03454f
C18985 VPWR.n1211 VGND 0.01723f
C18986 VPWR.n1212 VGND 0.00728f
C18987 VPWR.n1213 VGND 0.10877f
C18988 VPWR.t1432 VGND 0.09265f
C18989 VPWR.t1403 VGND 0.07889f
C18990 VPWR.t1421 VGND 0.12017f
C18991 VPWR.t1314 VGND 0.03348f
C18992 VPWR.t1393 VGND 0.02976f
C18993 VPWR.n1214 VGND 0.09198f
C18994 VPWR.n1215 VGND 0.00728f
C18995 VPWR.n1216 VGND 0.10877f
C18996 VPWR.t1392 VGND 0.09265f
C18997 VPWR.t1180 VGND 0.07889f
C18998 VPWR.t1313 VGND 0.12017f
C18999 VPWR.t1155 VGND 0.03348f
C19000 VPWR.t1285 VGND 0.02976f
C19001 VPWR.n1217 VGND 0.09198f
C19002 VPWR.n1218 VGND 0.00728f
C19003 VPWR.n1219 VGND 0.10877f
C19004 VPWR.t1284 VGND 0.09265f
C19005 VPWR.t1165 VGND 0.07889f
C19006 VPWR.t1154 VGND 0.12017f
C19007 VPWR.n1220 VGND 0.10877f
C19008 VPWR.n1221 VGND 0.00728f
C19009 VPWR.n1222 VGND 0.01723f
C19010 VPWR.n1223 VGND 0.00809f
C19011 VPWR.t2041 VGND 0.01122f
C19012 VPWR.t1320 VGND 0.01228f
C19013 VPWR.n1224 VGND 0.03058f
C19014 VPWR.n1225 VGND 0.00584f
C19015 VPWR.t1322 VGND 0.02693f
C19016 VPWR.n1226 VGND 0.05753f
C19017 VPWR.t1881 VGND 0.02976f
C19018 VPWR.n1227 VGND 0.04716f
C19019 VPWR.t1185 VGND 0.14585f
C19020 VPWR.t1170 VGND 0.07889f
C19021 VPWR.t1564 VGND 0.09265f
C19022 VPWR.t1948 VGND 0.01122f
C19023 VPWR.t1184 VGND 0.01228f
C19024 VPWR.n1228 VGND 0.03058f
C19025 VPWR.n1229 VGND 0.00584f
C19026 VPWR.t1186 VGND 0.02693f
C19027 VPWR.n1230 VGND 0.05753f
C19028 VPWR.t1565 VGND 0.02976f
C19029 VPWR.n1231 VGND 0.04716f
C19030 VPWR.n1232 VGND -0.01875f
C19031 VPWR.n1233 VGND 0.0471f
C19032 VPWR.t109 VGND 0.98059f
C19033 VPWR.n1234 VGND 0.53482f
C19034 VPWR.t32 VGND 0.98059f
C19035 VPWR.n1235 VGND 0.41593f
C19036 VPWR.n1236 VGND 0.29227f
C19037 VPWR.t110 VGND 0.05745f
C19038 VPWR.n1237 VGND 0.00925f
C19039 VPWR.t694 VGND 0.0144f
C19040 VPWR.t1827 VGND 0.0144f
C19041 VPWR.n1238 VGND 0.03162f
C19042 VPWR.t1828 VGND 0.0144f
C19043 VPWR.t611 VGND 0.0144f
C19044 VPWR.n1239 VGND 0.03156f
C19045 VPWR.t1769 VGND 0.0144f
C19046 VPWR.t1768 VGND 0.0144f
C19047 VPWR.n1240 VGND 0.03156f
C19048 VPWR.n1241 VGND 0.10473f
C19049 VPWR.n1242 VGND 0.18274f
C19050 VPWR.n1243 VGND 0.05786f
C19051 VPWR.n1244 VGND 0.0425f
C19052 VPWR.t1765 VGND 0.0144f
C19053 VPWR.t1770 VGND 0.0144f
C19054 VPWR.n1245 VGND 0.03162f
C19055 VPWR.n1246 VGND 0.12967f
C19056 VPWR.n1247 VGND 0.01124f
C19057 VPWR.n1248 VGND 0.01638f
C19058 VPWR.n1249 VGND 0.0192f
C19059 VPWR.n1250 VGND 0.02816f
C19060 VPWR.t107 VGND 0.05745f
C19061 VPWR.n1251 VGND 0.15135f
C19062 VPWR.n1252 VGND 0.01215f
C19063 VPWR.t1832 VGND 0.05743f
C19064 VPWR.t1848 VGND 0.05743f
C19065 VPWR.n1253 VGND 0.13514f
C19066 VPWR.n1254 VGND 0.33732f
C19067 VPWR.n1255 VGND 1.64922f
C19068 VPWR.n1256 VGND 0.0471f
C19069 VPWR.t34 VGND 0.98059f
C19070 VPWR.n1257 VGND 0.53482f
C19071 VPWR.t44 VGND 0.98059f
C19072 VPWR.n1258 VGND 0.41593f
C19073 VPWR.n1259 VGND 0.2949f
C19074 VPWR.n1260 VGND 0.00925f
C19075 VPWR.t1686 VGND 0.0144f
C19076 VPWR.t1684 VGND 0.0144f
C19077 VPWR.n1261 VGND 0.03162f
C19078 VPWR.t1683 VGND 0.0144f
C19079 VPWR.t1681 VGND 0.0144f
C19080 VPWR.n1262 VGND 0.03156f
C19081 VPWR.t813 VGND 0.0144f
C19082 VPWR.t915 VGND 0.0144f
C19083 VPWR.n1263 VGND 0.03156f
C19084 VPWR.n1264 VGND 0.10473f
C19085 VPWR.n1265 VGND 0.18274f
C19086 VPWR.n1266 VGND 0.05786f
C19087 VPWR.n1267 VGND 0.0425f
C19088 VPWR.t1925 VGND 0.0144f
C19089 VPWR.t102 VGND 0.0144f
C19090 VPWR.n1268 VGND 0.03162f
C19091 VPWR.n1269 VGND 0.12967f
C19092 VPWR.n1270 VGND 0.01124f
C19093 VPWR.n1271 VGND 0.01638f
C19094 VPWR.n1272 VGND 0.0192f
C19095 VPWR.n1273 VGND 0.02765f
C19096 VPWR.n1274 VGND 0.00771f
C19097 VPWR.t111 VGND 0.05737f
C19098 VPWR.n1275 VGND 0.06132f
C19099 VPWR.n1276 VGND 0.00734f
C19100 VPWR.t988 VGND 0.05749f
C19101 VPWR.n1277 VGND 0.09156f
C19102 VPWR.n1278 VGND 0.33732f
C19103 VPWR.n1279 VGND 1.64922f
C19104 VPWR.n1280 VGND 0.0471f
C19105 VPWR.t108 VGND 0.98059f
C19106 VPWR.n1281 VGND 0.53482f
C19107 VPWR.t104 VGND 0.98059f
C19108 VPWR.n1282 VGND 0.41593f
C19109 VPWR.n1283 VGND 0.2949f
C19110 VPWR.n1284 VGND 0.00925f
C19111 VPWR.t968 VGND 0.0144f
C19112 VPWR.t966 VGND 0.0144f
C19113 VPWR.n1285 VGND 0.03162f
C19114 VPWR.t965 VGND 0.0144f
C19115 VPWR.t964 VGND 0.0144f
C19116 VPWR.n1286 VGND 0.03156f
C19117 VPWR.t617 VGND 0.0144f
C19118 VPWR.t624 VGND 0.0144f
C19119 VPWR.n1287 VGND 0.03156f
C19120 VPWR.n1288 VGND 0.10473f
C19121 VPWR.n1289 VGND 0.18274f
C19122 VPWR.n1290 VGND 0.05786f
C19123 VPWR.n1291 VGND 0.0425f
C19124 VPWR.t621 VGND 0.0144f
C19125 VPWR.t618 VGND 0.0144f
C19126 VPWR.n1292 VGND 0.03162f
C19127 VPWR.n1293 VGND 0.12967f
C19128 VPWR.n1294 VGND 0.01124f
C19129 VPWR.n1295 VGND 0.01638f
C19130 VPWR.n1296 VGND 0.0192f
C19131 VPWR.n1297 VGND 0.02765f
C19132 VPWR.n1298 VGND 0.01405f
C19133 VPWR.n1299 VGND 0.01315f
C19134 VPWR.t1833 VGND 0.05749f
C19135 VPWR.t1849 VGND 0.05749f
C19136 VPWR.n1300 VGND 0.16979f
C19137 VPWR.n1301 VGND 0.33732f
C19138 VPWR.n1302 VGND 1.64922f
C19139 VPWR.t838 VGND 0.0574f
C19140 VPWR.t1869 VGND 0.05749f
C19141 VPWR.t840 VGND 0.057f
C19142 VPWR.n1303 VGND 0.1478f
C19143 VPWR.t380 VGND 0.05635f
C19144 VPWR.n1304 VGND 0.0681f
C19145 VPWR.n1305 VGND 0.0471f
C19146 VPWR.t442 VGND 0.05425f
C19147 VPWR.n1306 VGND 0.05159f
C19148 VPWR.t719 VGND 0.0144f
C19149 VPWR.t370 VGND 0.0144f
C19150 VPWR.n1307 VGND 0.03147f
C19151 VPWR.t1889 VGND 0.0504f
C19152 VPWR.n1308 VGND 0.07559f
C19153 VPWR.n1309 VGND 0.0471f
C19154 VPWR.t376 VGND 0.05743f
C19155 VPWR.n1310 VGND 0.0723f
C19156 VPWR.n1311 VGND 0.02765f
C19157 VPWR.n1312 VGND 0.0471f
C19158 VPWR.n1313 VGND 0.01215f
C19159 VPWR.t372 VGND 0.0144f
C19160 VPWR.t374 VGND 0.0144f
C19161 VPWR.n1314 VGND 0.03147f
C19162 VPWR.n1315 VGND 0.04611f
C19163 VPWR.n1316 VGND 0.01215f
C19164 VPWR.n1317 VGND 0.03533f
C19165 VPWR.n1318 VGND 0.03533f
C19166 VPWR.n1319 VGND 0.0471f
C19167 VPWR.n1320 VGND 0.00834f
C19168 VPWR.t715 VGND 0.0144f
C19169 VPWR.t438 VGND 0.0144f
C19170 VPWR.n1321 VGND 0.03147f
C19171 VPWR.n1322 VGND 0.03623f
C19172 VPWR.t382 VGND 0.0144f
C19173 VPWR.t609 VGND 0.0144f
C19174 VPWR.n1323 VGND 0.03147f
C19175 VPWR.n1324 VGND 0.04004f
C19176 VPWR.n1325 VGND 0.01061f
C19177 VPWR.n1326 VGND 0.04275f
C19178 VPWR.n1327 VGND 0.01613f
C19179 VPWR.n1328 VGND 0.00635f
C19180 VPWR.t415 VGND 0.0483f
C19181 VPWR.t837 VGND 0.10867f
C19182 VPWR.t1868 VGND 0.12678f
C19183 VPWR.t839 VGND 0.23545f
C19184 VPWR.t375 VGND 0.12669f
C19185 VPWR.t373 VGND 0.14381f
C19186 VPWR.t371 VGND 0.13981f
C19187 VPWR.t369 VGND 0.22359f
C19188 VPWR.t718 VGND 0.19017f
C19189 VPWR.t1888 VGND 0.12678f
C19190 VPWR.t437 VGND 0.12678f
C19191 VPWR.t608 VGND 0.12678f
C19192 VPWR.t714 VGND 0.12678f
C19193 VPWR.t381 VGND 0.12678f
C19194 VPWR.t441 VGND 0.12678f
C19195 VPWR.t379 VGND 0.12527f
C19196 VPWR.n1329 VGND 0.43087f
C19197 VPWR.n1330 VGND 0.17507f
C19198 VPWR.n1331 VGND 0.0192f
C19199 VPWR.n1332 VGND 0.03533f
C19200 VPWR.n1333 VGND 0.0425f
C19201 VPWR.n1334 VGND 0.01088f
C19202 VPWR.n1335 VGND 0.06389f
C19203 VPWR.n1336 VGND 0.31812f
C19204 VPWR.n1337 VGND 1.64922f
C19205 VPWR.t100 VGND 0.05647f
C19206 VPWR.t711 VGND 0.05631f
C19207 VPWR.t283 VGND 0.05743f
C19208 VPWR.n1338 VGND 0.08004f
C19209 VPWR.t1829 VGND 0.05483f
C19210 VPWR.t1771 VGND 0.05483f
C19211 VPWR.n1339 VGND 0.09948f
C19212 VPWR.n1340 VGND 0.0471f
C19213 VPWR.n1341 VGND 0.00916f
C19214 VPWR.n1342 VGND 0.0471f
C19215 VPWR.t695 VGND 0.0144f
C19216 VPWR.t1693 VGND 0.0144f
C19217 VPWR.n1343 VGND 0.03147f
C19218 VPWR.t1772 VGND 0.0144f
C19219 VPWR.t36 VGND 0.0144f
C19220 VPWR.n1344 VGND 0.03147f
C19221 VPWR.n1345 VGND 0.06411f
C19222 VPWR.t39 VGND 0.05743f
C19223 VPWR.t1689 VGND 0.05743f
C19224 VPWR.n1346 VGND 0.13235f
C19225 VPWR.n1347 VGND 0.02765f
C19226 VPWR.n1348 VGND 0.0471f
C19227 VPWR.n1349 VGND 0.01215f
C19228 VPWR.t731 VGND 0.0144f
C19229 VPWR.t1891 VGND 0.0144f
C19230 VPWR.n1350 VGND 0.03147f
C19231 VPWR.t45 VGND 0.0144f
C19232 VPWR.t1696 VGND 0.0144f
C19233 VPWR.n1351 VGND 0.03147f
C19234 VPWR.n1352 VGND 0.07246f
C19235 VPWR.n1353 VGND 0.01215f
C19236 VPWR.n1354 VGND 0.0471f
C19237 VPWR.n1355 VGND 0.0471f
C19238 VPWR.n1356 VGND 0.0471f
C19239 VPWR.n1357 VGND 0.01133f
C19240 VPWR.t612 VGND 0.0144f
C19241 VPWR.t696 VGND 0.0144f
C19242 VPWR.n1358 VGND 0.03147f
C19243 VPWR.t1767 VGND 0.0144f
C19244 VPWR.t1766 VGND 0.0144f
C19245 VPWR.n1359 VGND 0.03147f
C19246 VPWR.n1360 VGND 0.06411f
C19247 VPWR.n1361 VGND 0.01061f
C19248 VPWR.n1362 VGND 0.00988f
C19249 VPWR.n1363 VGND 0.0471f
C19250 VPWR.n1364 VGND 0.03533f
C19251 VPWR.n1365 VGND 0.00798f
C19252 VPWR.t38 VGND 0.98059f
C19253 VPWR.n1366 VGND 0.53482f
C19254 VPWR.t35 VGND 0.98059f
C19255 VPWR.n1367 VGND 0.41593f
C19256 VPWR.n1368 VGND 0.29227f
C19257 VPWR.n1369 VGND 0.0192f
C19258 VPWR.n1370 VGND 0.03533f
C19259 VPWR.n1371 VGND 0.04275f
C19260 VPWR.n1372 VGND 0.0107f
C19261 VPWR.n1373 VGND 0.05857f
C19262 VPWR.n1374 VGND 0.07933f
C19263 VPWR.n1375 VGND 0.31787f
C19264 VPWR.n1376 VGND 1.64922f
C19265 VPWR.t547 VGND 0.05737f
C19266 VPWR.t1653 VGND 0.05737f
C19267 VPWR.n1377 VGND 0.01405f
C19268 VPWR.t1682 VGND 0.05483f
C19269 VPWR.t101 VGND 0.05483f
C19270 VPWR.n1378 VGND 0.09948f
C19271 VPWR.n1379 VGND 0.0471f
C19272 VPWR.n1380 VGND 0.00916f
C19273 VPWR.n1381 VGND 0.0471f
C19274 VPWR.t1687 VGND 0.0144f
C19275 VPWR.t41 VGND 0.0144f
C19276 VPWR.n1382 VGND 0.03147f
C19277 VPWR.t17 VGND 0.0144f
C19278 VPWR.t1690 VGND 0.0144f
C19279 VPWR.n1383 VGND 0.03147f
C19280 VPWR.n1384 VGND 0.06411f
C19281 VPWR.t1691 VGND 0.05743f
C19282 VPWR.t33 VGND 0.05743f
C19283 VPWR.n1385 VGND 0.13235f
C19284 VPWR.n1386 VGND 0.02765f
C19285 VPWR.n1387 VGND 0.0471f
C19286 VPWR.n1388 VGND 0.01215f
C19287 VPWR.t1695 VGND 0.0144f
C19288 VPWR.t607 VGND 0.0144f
C19289 VPWR.n1389 VGND 0.03147f
C19290 VPWR.t1692 VGND 0.0144f
C19291 VPWR.t733 VGND 0.0144f
C19292 VPWR.n1390 VGND 0.03147f
C19293 VPWR.n1391 VGND 0.07246f
C19294 VPWR.n1392 VGND 0.01215f
C19295 VPWR.n1393 VGND 0.0471f
C19296 VPWR.n1394 VGND 0.0471f
C19297 VPWR.n1395 VGND 0.0471f
C19298 VPWR.n1396 VGND 0.01133f
C19299 VPWR.t1688 VGND 0.0144f
C19300 VPWR.t1685 VGND 0.0144f
C19301 VPWR.n1397 VGND 0.03147f
C19302 VPWR.t916 VGND 0.0144f
C19303 VPWR.t1924 VGND 0.0144f
C19304 VPWR.n1398 VGND 0.03147f
C19305 VPWR.n1399 VGND 0.06411f
C19306 VPWR.n1400 VGND 0.01061f
C19307 VPWR.n1401 VGND 0.00988f
C19308 VPWR.n1402 VGND 0.0471f
C19309 VPWR.n1403 VGND 0.03533f
C19310 VPWR.n1404 VGND 0.00798f
C19311 VPWR.t40 VGND 0.98059f
C19312 VPWR.n1405 VGND 0.53482f
C19313 VPWR.t16 VGND 0.98059f
C19314 VPWR.n1406 VGND 0.41593f
C19315 VPWR.n1407 VGND 0.2949f
C19316 VPWR.n1408 VGND 0.0192f
C19317 VPWR.n1409 VGND 0.03533f
C19318 VPWR.n1410 VGND 0.04275f
C19319 VPWR.n1411 VGND 0.01088f
C19320 VPWR.n1412 VGND 0.11596f
C19321 VPWR.n1413 VGND 0.32299f
C19322 VPWR.n1414 VGND 1.64922f
C19323 VPWR.t967 VGND 0.05483f
C19324 VPWR.t619 VGND 0.05483f
C19325 VPWR.n1415 VGND 0.09948f
C19326 VPWR.n1416 VGND 0.0471f
C19327 VPWR.n1417 VGND 0.00916f
C19328 VPWR.n1418 VGND 0.0471f
C19329 VPWR.t962 VGND 0.0144f
C19330 VPWR.t730 VGND 0.0144f
C19331 VPWR.n1419 VGND 0.03147f
C19332 VPWR.t620 VGND 0.0144f
C19333 VPWR.t1893 VGND 0.0144f
C19334 VPWR.n1420 VGND 0.03147f
C19335 VPWR.n1421 VGND 0.06411f
C19336 VPWR.t43 VGND 0.05743f
C19337 VPWR.t1072 VGND 0.05743f
C19338 VPWR.n1422 VGND 0.13235f
C19339 VPWR.n1423 VGND 0.02765f
C19340 VPWR.n1424 VGND 0.0471f
C19341 VPWR.n1425 VGND 0.01215f
C19342 VPWR.t732 VGND 0.0144f
C19343 VPWR.t1892 VGND 0.0144f
C19344 VPWR.n1426 VGND 0.03147f
C19345 VPWR.t378 VGND 0.0144f
C19346 VPWR.t383 VGND 0.0144f
C19347 VPWR.n1427 VGND 0.03147f
C19348 VPWR.n1428 VGND 0.07246f
C19349 VPWR.n1429 VGND 0.01215f
C19350 VPWR.n1430 VGND 0.0471f
C19351 VPWR.n1431 VGND 0.0471f
C19352 VPWR.n1432 VGND 0.0471f
C19353 VPWR.n1433 VGND 0.01133f
C19354 VPWR.t963 VGND 0.0144f
C19355 VPWR.t961 VGND 0.0144f
C19356 VPWR.n1434 VGND 0.03147f
C19357 VPWR.t623 VGND 0.0144f
C19358 VPWR.t622 VGND 0.0144f
C19359 VPWR.n1435 VGND 0.03147f
C19360 VPWR.n1436 VGND 0.06411f
C19361 VPWR.n1437 VGND 0.01061f
C19362 VPWR.n1438 VGND 0.00988f
C19363 VPWR.n1439 VGND 0.0471f
C19364 VPWR.n1440 VGND 0.03533f
C19365 VPWR.n1441 VGND 0.00798f
C19366 VPWR.t42 VGND 0.75221f
C19367 VPWR.n1442 VGND 0.43036f
C19368 VPWR.t377 VGND 0.75221f
C19369 VPWR.n1443 VGND 0.33723f
C19370 VPWR.n1444 VGND 0.28271f
C19371 VPWR.n1445 VGND 0.4322f
C19372 VPWR.n1446 VGND 6.28433f
C19373 VPWR.n1447 VGND 9.20004f
C19374 VPWR.n1448 VGND 0.08393f
C19375 VPWR.n1449 VGND 1.10545f
C19376 VPWR.n1450 VGND 1.01451f
C19377 VPWR.n1451 VGND 0.06515f
C19378 VPWR.n1452 VGND 0.05468f
C19379 VPWR.t2045 VGND 0.01141f
C19380 VPWR.t1169 VGND 0.01247f
C19381 VPWR.n1453 VGND 0.02783f
C19382 VPWR.n1454 VGND 0.01907f
C19383 VPWR.n1455 VGND 0.06276f
C19384 VPWR.n1456 VGND 0.07802f
C19385 VPWR.n1457 VGND 0.09221f
C19386 VPWR.t1996 VGND 0.01141f
C19387 VPWR.t1300 VGND 0.01247f
C19388 VPWR.n1458 VGND 0.02783f
C19389 VPWR.n1459 VGND 0.01907f
C19390 VPWR.n1460 VGND 0.06276f
C19391 VPWR.n1461 VGND 0.09795f
C19392 VPWR.n1462 VGND 0.09221f
C19393 VPWR.n1463 VGND 0.066f
C19394 VPWR.n1464 VGND 0.05468f
C19395 VPWR.n1465 VGND 0.13984f
C19396 VPWR.n1466 VGND 0.01806f
C19397 VPWR.n1467 VGND 0.00732f
C19398 VPWR.n1468 VGND 0.10877f
C19399 VPWR.t1346 VGND 0.12017f
C19400 VPWR.t1301 VGND 0.07889f
C19401 VPWR.t709 VGND 0.09265f
C19402 VPWR.t2044 VGND 0.01122f
C19403 VPWR.t1345 VGND 0.01228f
C19404 VPWR.n1469 VGND 0.03058f
C19405 VPWR.n1470 VGND 0.00584f
C19406 VPWR.t1347 VGND 0.02693f
C19407 VPWR.n1471 VGND 0.05753f
C19408 VPWR.t710 VGND 0.02976f
C19409 VPWR.n1472 VGND 0.04716f
C19410 VPWR.n1473 VGND 0.01806f
C19411 VPWR.n1474 VGND 0.00732f
C19412 VPWR.n1475 VGND 0.10877f
C19413 VPWR.t1448 VGND 0.12017f
C19414 VPWR.t1430 VGND 0.07889f
C19415 VPWR.t1517 VGND 0.09265f
C19416 VPWR.t1994 VGND 0.01122f
C19417 VPWR.t1447 VGND 0.01228f
C19418 VPWR.n1476 VGND 0.03058f
C19419 VPWR.n1477 VGND 0.00584f
C19420 VPWR.t1449 VGND 0.02693f
C19421 VPWR.n1478 VGND 0.05753f
C19422 VPWR.t1518 VGND 0.02976f
C19423 VPWR.n1479 VGND 0.04716f
C19424 VPWR.n1480 VGND 0.00732f
C19425 VPWR.n1481 VGND 0.10877f
C19426 VPWR.t1219 VGND 0.12017f
C19427 VPWR.t1089 VGND 0.07889f
C19428 VPWR.t149 VGND 0.09265f
C19429 VPWR.t1982 VGND 0.01122f
C19430 VPWR.t1218 VGND 0.01228f
C19431 VPWR.n1482 VGND 0.03058f
C19432 VPWR.n1483 VGND 0.00584f
C19433 VPWR.t1220 VGND 0.02693f
C19434 VPWR.n1484 VGND 0.05753f
C19435 VPWR.t150 VGND 0.02976f
C19436 VPWR.n1485 VGND 0.04716f
C19437 VPWR.n1486 VGND 0.00809f
C19438 VPWR.n1487 VGND 0.08393f
C19439 VPWR.n1488 VGND -0.01875f
C19440 VPWR.n1489 VGND 0.13984f
C19441 VPWR.n1490 VGND 0.01806f
C19442 VPWR.n1491 VGND 0.00732f
C19443 VPWR.n1492 VGND 0.10877f
C19444 VPWR.t1321 VGND 0.12017f
C19445 VPWR.t1196 VGND 0.07889f
C19446 VPWR.t1880 VGND 0.09265f
C19447 VPWR.t1351 VGND 0.07889f
C19448 VPWR.t1343 VGND 0.12017f
C19449 VPWR.n1493 VGND 0.10877f
C19450 VPWR.n1494 VGND 0.00732f
C19451 VPWR.n1495 VGND 0.01806f
C19452 VPWR.n1496 VGND 0.05468f
C19453 VPWR.n1497 VGND 0.13984f
C19454 VPWR.n1498 VGND -0.01875f
C19455 VPWR.n1499 VGND 0.08393f
C19456 VPWR.n1500 VGND 0.08393f
C19457 VPWR.n1501 VGND -0.01875f
C19458 VPWR.n1502 VGND 0.05468f
C19459 VPWR.n1503 VGND 0.13984f
C19460 VPWR.n1504 VGND 0.01806f
C19461 VPWR.n1505 VGND 0.00732f
C19462 VPWR.n1506 VGND 0.10877f
C19463 VPWR.t1094 VGND 0.12017f
C19464 VPWR.t1353 VGND 0.07889f
C19465 VPWR.t281 VGND 0.09265f
C19466 VPWR.t1201 VGND 0.07889f
C19467 VPWR.t1216 VGND 0.12017f
C19468 VPWR.n1507 VGND 0.10877f
C19469 VPWR.n1508 VGND 0.00732f
C19470 VPWR.n1509 VGND 0.01806f
C19471 VPWR.n1510 VGND 0.05468f
C19472 VPWR.n1511 VGND 0.13984f
C19473 VPWR.n1512 VGND -0.01875f
C19474 VPWR.n1513 VGND 0.08393f
C19475 VPWR.n1514 VGND 0.08393f
C19476 VPWR.n1515 VGND -0.01875f
C19477 VPWR.n1516 VGND 0.05468f
C19478 VPWR.n1517 VGND 0.13984f
C19479 VPWR.n1518 VGND 0.01806f
C19480 VPWR.n1519 VGND 0.00732f
C19481 VPWR.n1520 VGND 0.10877f
C19482 VPWR.t1357 VGND 0.12017f
C19483 VPWR.t1231 VGND 0.07889f
C19484 VPWR.t1068 VGND 0.09265f
C19485 VPWR.t1349 VGND 0.07889f
C19486 VPWR.t1373 VGND 0.12017f
C19487 VPWR.n1521 VGND 0.10877f
C19488 VPWR.n1522 VGND 0.00732f
C19489 VPWR.n1523 VGND 0.01806f
C19490 VPWR.n1524 VGND 0.05468f
C19491 VPWR.n1525 VGND 0.13984f
C19492 VPWR.n1526 VGND -0.01875f
C19493 VPWR.n1527 VGND 0.08393f
C19494 VPWR.n1528 VGND 0.08393f
C19495 VPWR.n1529 VGND 0.08393f
C19496 VPWR.n1530 VGND 0.08393f
C19497 VPWR.n1531 VGND -0.01875f
C19498 VPWR.n1532 VGND 0.13984f
C19499 VPWR.n1533 VGND 0.01806f
C19500 VPWR.n1534 VGND 0.00732f
C19501 VPWR.n1535 VGND 0.10877f
C19502 VPWR.t770 VGND 0.09265f
C19503 VPWR.t1100 VGND 0.07889f
C19504 VPWR.t1116 VGND 0.12017f
C19505 VPWR.n1536 VGND 0.10877f
C19506 VPWR.n1537 VGND 0.00732f
C19507 VPWR.n1538 VGND 0.01806f
C19508 VPWR.n1539 VGND 0.13984f
C19509 VPWR.n1540 VGND 0.05468f
C19510 VPWR.n1541 VGND 0.066f
C19511 VPWR.n1542 VGND 0.09221f
C19512 VPWR.t1929 VGND 0.01141f
C19513 VPWR.t1099 VGND 0.01247f
C19514 VPWR.n1543 VGND 0.02783f
C19515 VPWR.n1544 VGND 0.01907f
C19516 VPWR.n1545 VGND 0.06276f
C19517 VPWR.n1546 VGND 0.09795f
C19518 VPWR.n1547 VGND 0.09221f
C19519 VPWR.t1986 VGND 0.01141f
C19520 VPWR.t1348 VGND 0.01247f
C19521 VPWR.n1548 VGND 0.02783f
C19522 VPWR.n1549 VGND 0.01907f
C19523 VPWR.n1550 VGND 0.06276f
C19524 VPWR.n1551 VGND 0.09795f
C19525 VPWR.n1552 VGND 0.09221f
C19526 VPWR.t2025 VGND 0.01141f
C19527 VPWR.t1230 VGND 0.01247f
C19528 VPWR.n1553 VGND 0.02783f
C19529 VPWR.n1554 VGND 0.01907f
C19530 VPWR.n1555 VGND 0.06276f
C19531 VPWR.n1556 VGND 0.09795f
C19532 VPWR.n1557 VGND 0.09221f
C19533 VPWR.t2037 VGND 0.01141f
C19534 VPWR.t1200 VGND 0.01247f
C19535 VPWR.n1558 VGND 0.02783f
C19536 VPWR.n1559 VGND 0.01907f
C19537 VPWR.n1560 VGND 0.06276f
C19538 VPWR.n1561 VGND 0.09795f
C19539 VPWR.n1562 VGND 0.09221f
C19540 VPWR.t1979 VGND 0.01141f
C19541 VPWR.t1352 VGND 0.01247f
C19542 VPWR.n1563 VGND 0.02783f
C19543 VPWR.n1564 VGND 0.01907f
C19544 VPWR.n1565 VGND 0.06276f
C19545 VPWR.n1566 VGND 0.09795f
C19546 VPWR.n1567 VGND 0.09221f
C19547 VPWR.t1985 VGND 0.01141f
C19548 VPWR.t1350 VGND 0.01247f
C19549 VPWR.n1568 VGND 0.02783f
C19550 VPWR.n1569 VGND 0.01907f
C19551 VPWR.n1570 VGND 0.06276f
C19552 VPWR.n1571 VGND 0.09795f
C19553 VPWR.n1572 VGND 0.09221f
C19554 VPWR.t2039 VGND 0.01141f
C19555 VPWR.t1195 VGND 0.01247f
C19556 VPWR.n1573 VGND 0.02783f
C19557 VPWR.n1574 VGND 0.01907f
C19558 VPWR.n1575 VGND 0.06276f
C19559 VPWR.n1576 VGND 0.09795f
C19560 VPWR.n1577 VGND 0.09221f
C19561 VPWR.t1936 VGND 0.01141f
C19562 VPWR.t1088 VGND 0.01247f
C19563 VPWR.n1578 VGND 0.02783f
C19564 VPWR.n1579 VGND 0.01907f
C19565 VPWR.n1580 VGND 0.06276f
C19566 VPWR.n1581 VGND 0.09795f
C19567 VPWR.n1582 VGND 0.09221f
C19568 VPWR.n1583 VGND 0.066f
C19569 VPWR.n1584 VGND 0.05468f
C19570 VPWR.n1585 VGND 0.13984f
C19571 VPWR.n1586 VGND -0.01875f
C19572 VPWR.n1587 VGND 0.08393f
C19573 VPWR.n1588 VGND 0.08393f
C19574 VPWR.n1589 VGND -0.01875f
C19575 VPWR.n1590 VGND 0.00809f
C19576 VPWR.n1591 VGND 0.01723f
C19577 VPWR.n1592 VGND 0.00728f
C19578 VPWR.n1593 VGND 0.10877f
C19579 VPWR.t1243 VGND 0.09265f
C19580 VPWR.t1124 VGND 0.07889f
C19581 VPWR.t1157 VGND 0.12017f
C19582 VPWR.n1594 VGND 0.10877f
C19583 VPWR.n1595 VGND 0.00728f
C19584 VPWR.n1596 VGND 0.01723f
C19585 VPWR.n1597 VGND 0.03454f
C19586 VPWR.t1966 VGND 0.01122f
C19587 VPWR.t1156 VGND 0.01228f
C19588 VPWR.n1598 VGND 0.03131f
C19589 VPWR.n1599 VGND 0.03712f
C19590 VPWR.n1600 VGND 0.00837f
C19591 VPWR.t2063 VGND 0.01141f
C19592 VPWR.t1123 VGND 0.01247f
C19593 VPWR.n1601 VGND 0.02782f
C19594 VPWR.n1602 VGND 0.02832f
C19595 VPWR.n1603 VGND 0.01785f
C19596 VPWR.n1604 VGND 0.00701f
C19597 VPWR.n1605 VGND 0.01831f
C19598 VPWR.n1606 VGND 0.02396f
C19599 VPWR.n1607 VGND 0.23844f
C19600 VPWR.n1608 VGND 0.17674f
C19601 VPWR.n1609 VGND 0.02396f
C19602 VPWR.n1610 VGND 0.01785f
C19603 VPWR.t2010 VGND 0.01125f
C19604 VPWR.t1255 VGND 0.01232f
C19605 VPWR.n1611 VGND 0.03008f
C19606 VPWR.n1612 VGND 0.03301f
C19607 VPWR.n1613 VGND 0.03454f
C19608 VPWR.t2047 VGND 0.01122f
C19609 VPWR.t1423 VGND 0.01228f
C19610 VPWR.n1614 VGND 0.03131f
C19611 VPWR.n1615 VGND 0.03712f
C19612 VPWR.n1616 VGND 0.00837f
C19613 VPWR.t2000 VGND 0.01141f
C19614 VPWR.t1289 VGND 0.01247f
C19615 VPWR.n1617 VGND 0.02782f
C19616 VPWR.n1618 VGND 0.02832f
C19617 VPWR.n1619 VGND 0.01831f
C19618 VPWR.n1620 VGND 0.02396f
C19619 VPWR.n1621 VGND 0.01785f
C19620 VPWR.t1955 VGND 0.01125f
C19621 VPWR.t1415 VGND 0.01232f
C19622 VPWR.n1622 VGND 0.03008f
C19623 VPWR.n1623 VGND 0.03301f
C19624 VPWR.n1624 VGND 0.03454f
C19625 VPWR.t1965 VGND 0.01122f
C19626 VPWR.t1141 VGND 0.01228f
C19627 VPWR.n1625 VGND 0.03131f
C19628 VPWR.n1626 VGND 0.03712f
C19629 VPWR.n1627 VGND 0.00837f
C19630 VPWR.t1962 VGND 0.01141f
C19631 VPWR.t1397 VGND 0.01247f
C19632 VPWR.n1628 VGND 0.02782f
C19633 VPWR.n1629 VGND 0.02832f
C19634 VPWR.n1630 VGND 0.01785f
C19635 VPWR.n1631 VGND 0.00701f
C19636 VPWR.n1632 VGND 0.01831f
C19637 VPWR.n1633 VGND 0.02396f
C19638 VPWR.n1634 VGND 0.17674f
C19639 VPWR.n1635 VGND 0.17674f
C19640 VPWR.n1636 VGND 0.02396f
C19641 VPWR.n1637 VGND 0.01785f
C19642 VPWR.t2002 VGND 0.01125f
C19643 VPWR.t1283 VGND 0.01232f
C19644 VPWR.n1638 VGND 0.03008f
C19645 VPWR.n1639 VGND 0.03301f
C19646 VPWR.n1640 VGND 0.03454f
C19647 VPWR.t1944 VGND 0.01122f
C19648 VPWR.t1312 VGND 0.01228f
C19649 VPWR.n1641 VGND 0.03131f
C19650 VPWR.n1642 VGND 0.03712f
C19651 VPWR.n1643 VGND 0.00837f
C19652 VPWR.t2042 VGND 0.01141f
C19653 VPWR.t1179 VGND 0.01247f
C19654 VPWR.n1644 VGND 0.02782f
C19655 VPWR.n1645 VGND 0.02832f
C19656 VPWR.n1646 VGND 0.01831f
C19657 VPWR.n1647 VGND 0.02396f
C19658 VPWR.n1648 VGND 0.01785f
C19659 VPWR.t1964 VGND 0.01125f
C19660 VPWR.t1391 VGND 0.01232f
C19661 VPWR.n1649 VGND 0.03008f
C19662 VPWR.n1650 VGND 0.03301f
C19663 VPWR.n1651 VGND 0.03454f
C19664 VPWR.t2005 VGND 0.01122f
C19665 VPWR.t1420 VGND 0.01228f
C19666 VPWR.n1652 VGND 0.03131f
C19667 VPWR.n1653 VGND 0.03712f
C19668 VPWR.n1654 VGND 0.00837f
C19669 VPWR.t1959 VGND 0.01141f
C19670 VPWR.t1402 VGND 0.01247f
C19671 VPWR.n1655 VGND 0.02782f
C19672 VPWR.n1656 VGND 0.02832f
C19673 VPWR.n1657 VGND 0.01785f
C19674 VPWR.n1658 VGND 0.00701f
C19675 VPWR.n1659 VGND 0.01831f
C19676 VPWR.n1660 VGND 0.02396f
C19677 VPWR.n1661 VGND 0.17674f
C19678 VPWR.n1662 VGND 0.17674f
C19679 VPWR.n1663 VGND 0.02396f
C19680 VPWR.n1664 VGND 0.01785f
C19681 VPWR.t2043 VGND 0.01125f
C19682 VPWR.t1176 VGND 0.01232f
C19683 VPWR.n1665 VGND 0.03008f
C19684 VPWR.n1666 VGND 0.03301f
C19685 VPWR.n1667 VGND 0.03454f
C19686 VPWR.t1941 VGND 0.01122f
C19687 VPWR.t1207 VGND 0.01228f
C19688 VPWR.n1668 VGND 0.03131f
C19689 VPWR.n1669 VGND 0.03712f
C19690 VPWR.n1670 VGND 0.00837f
C19691 VPWR.t2050 VGND 0.01141f
C19692 VPWR.t1162 VGND 0.01247f
C19693 VPWR.n1671 VGND 0.02782f
C19694 VPWR.n1672 VGND 0.02832f
C19695 VPWR.n1673 VGND 0.01831f
C19696 VPWR.n1674 VGND 0.02396f
C19697 VPWR.n1675 VGND 0.01785f
C19698 VPWR.t2003 VGND 0.01125f
C19699 VPWR.t1280 VGND 0.01232f
C19700 VPWR.n1676 VGND 0.03008f
C19701 VPWR.n1677 VGND 0.03301f
C19702 VPWR.n1678 VGND 0.03454f
C19703 VPWR.t2038 VGND 0.01122f
C19704 VPWR.t1334 VGND 0.01228f
C19705 VPWR.n1679 VGND 0.03131f
C19706 VPWR.n1680 VGND 0.03712f
C19707 VPWR.n1681 VGND 0.00837f
C19708 VPWR.t1993 VGND 0.01141f
C19709 VPWR.t1315 VGND 0.01247f
C19710 VPWR.n1682 VGND 0.02782f
C19711 VPWR.n1683 VGND 0.02832f
C19712 VPWR.n1684 VGND 0.01785f
C19713 VPWR.n1685 VGND 0.00701f
C19714 VPWR.n1686 VGND 0.01831f
C19715 VPWR.n1687 VGND 0.02396f
C19716 VPWR.n1688 VGND 0.17674f
C19717 VPWR.n1689 VGND 0.17674f
C19718 VPWR.n1690 VGND 0.02396f
C19719 VPWR.n1691 VGND 0.01785f
C19720 VPWR.t1939 VGND 0.01125f
C19721 VPWR.t1458 VGND 0.01232f
C19722 VPWR.n1692 VGND 0.03008f
C19723 VPWR.n1693 VGND 0.03301f
C19724 VPWR.n1694 VGND 0.03454f
C19725 VPWR.t1978 VGND 0.01122f
C19726 VPWR.t1101 VGND 0.01228f
C19727 VPWR.n1695 VGND 0.03131f
C19728 VPWR.n1696 VGND 0.03712f
C19729 VPWR.n1697 VGND 0.00837f
C19730 VPWR.t2040 VGND 0.01141f
C19731 VPWR.t1187 VGND 0.01247f
C19732 VPWR.n1698 VGND 0.02782f
C19733 VPWR.n1699 VGND 0.02832f
C19734 VPWR.n1700 VGND 0.01831f
C19735 VPWR.n1701 VGND 0.02396f
C19736 VPWR.n1702 VGND 0.01785f
C19737 VPWR.t2036 VGND 0.01125f
C19738 VPWR.t1202 VGND 0.01232f
C19739 VPWR.n1703 VGND 0.03008f
C19740 VPWR.n1704 VGND 0.03301f
C19741 VPWR.n1705 VGND 0.03454f
C19742 VPWR.t1935 VGND 0.01122f
C19743 VPWR.t1339 VGND 0.01228f
C19744 VPWR.n1706 VGND 0.03131f
C19745 VPWR.n1707 VGND 0.03712f
C19746 VPWR.n1708 VGND 0.00837f
C19747 VPWR.t2033 VGND 0.01141f
C19748 VPWR.t1213 VGND 0.01247f
C19749 VPWR.n1709 VGND 0.02782f
C19750 VPWR.n1710 VGND 0.02832f
C19751 VPWR.n1711 VGND 0.01785f
C19752 VPWR.n1712 VGND 0.00701f
C19753 VPWR.n1713 VGND 0.01831f
C19754 VPWR.n1714 VGND 0.02396f
C19755 VPWR.n1715 VGND 0.17674f
C19756 VPWR.t1977 VGND 0.01125f
C19757 VPWR.t1359 VGND 0.01232f
C19758 VPWR.n1716 VGND 0.03008f
C19759 VPWR.n1717 VGND 0.03301f
C19760 VPWR.t2024 VGND 0.01122f
C19761 VPWR.t1367 VGND 0.01228f
C19762 VPWR.n1718 VGND 0.03131f
C19763 VPWR.n1719 VGND 0.03712f
C19764 VPWR.n1720 VGND 0.00837f
C19765 VPWR.t2019 VGND 0.01141f
C19766 VPWR.t1238 VGND 0.01247f
C19767 VPWR.n1721 VGND 0.02782f
C19768 VPWR.n1722 VGND 0.02832f
C19769 VPWR.n1723 VGND 0.01785f
C19770 VPWR.n1724 VGND 0.00701f
C19771 VPWR.n1725 VGND 0.01831f
C19772 VPWR.n1726 VGND 0.02396f
C19773 VPWR.n1727 VGND 0.2127f
C19774 VPWR.n1728 VGND 0.02554f
C19775 VPWR.n1729 VGND 0.01785f
C19776 VPWR.t1937 VGND 0.01141f
C19777 VPWR.t1086 VGND 0.01247f
C19778 VPWR.n1730 VGND 0.02782f
C19779 VPWR.n1731 VGND 0.02832f
C19780 VPWR.n1732 VGND 0.00837f
C19781 VPWR.t1984 VGND 0.01122f
C19782 VPWR.t1083 VGND 0.01228f
C19783 VPWR.n1733 VGND 0.03131f
C19784 VPWR.n1734 VGND 0.03712f
C19785 VPWR.n1735 VGND 0.03454f
C19786 VPWR.n1736 VGND 0.00809f
C19787 VPWR.n1737 VGND 0.01723f
C19788 VPWR.n1738 VGND 0.00728f
C19789 VPWR.n1739 VGND 0.10877f
C19790 VPWR.t1360 VGND 0.09265f
C19791 VPWR.t1239 VGND 0.07889f
C19792 VPWR.t1368 VGND 0.12017f
C19793 VPWR.n1740 VGND 0.10877f
C19794 VPWR.n1741 VGND 0.00728f
C19795 VPWR.n1742 VGND 0.01723f
C19796 VPWR.n1743 VGND 0.00809f
C19797 VPWR.n1744 VGND 0.05468f
C19798 VPWR.t2011 VGND 0.01122f
C19799 VPWR.t1109 VGND 0.01228f
C19800 VPWR.n1745 VGND 0.03058f
C19801 VPWR.n1746 VGND 0.00584f
C19802 VPWR.t1111 VGND 0.02693f
C19803 VPWR.n1747 VGND 0.05753f
C19804 VPWR.t1024 VGND 0.02976f
C19805 VPWR.n1748 VGND 0.04716f
C19806 VPWR.t1381 VGND 0.07889f
C19807 VPWR.t1023 VGND 0.09265f
C19808 VPWR.t1419 VGND 0.07889f
C19809 VPWR.t1160 VGND 0.12017f
C19810 VPWR.n1749 VGND 0.10877f
C19811 VPWR.n1750 VGND 0.00732f
C19812 VPWR.n1751 VGND 0.01806f
C19813 VPWR.n1752 VGND 0.13984f
C19814 VPWR.n1753 VGND -0.01875f
C19815 VPWR.n1754 VGND 0.08393f
C19816 VPWR.n1755 VGND 0.08393f
C19817 VPWR.n1756 VGND -0.01875f
C19818 VPWR.n1757 VGND 0.13984f
C19819 VPWR.n1758 VGND 0.01806f
C19820 VPWR.n1759 VGND 0.00732f
C19821 VPWR.n1760 VGND 0.10877f
C19822 VPWR.t94 VGND 0.09265f
C19823 VPWR.t1363 VGND 0.07889f
C19824 VPWR.t1287 VGND 0.12017f
C19825 VPWR.n1761 VGND 0.10877f
C19826 VPWR.n1762 VGND 0.00732f
C19827 VPWR.n1763 VGND 0.01806f
C19828 VPWR.n1764 VGND 0.13984f
C19829 VPWR.n1765 VGND 0.05468f
C19830 VPWR.n1766 VGND 0.066f
C19831 VPWR.n1767 VGND 0.09221f
C19832 VPWR.t1976 VGND 0.01141f
C19833 VPWR.t1362 VGND 0.01247f
C19834 VPWR.n1768 VGND 0.02783f
C19835 VPWR.n1769 VGND 0.01907f
C19836 VPWR.n1770 VGND 0.06276f
C19837 VPWR.n1771 VGND 0.09795f
C19838 VPWR.n1772 VGND 0.09221f
C19839 VPWR.t1968 VGND 0.01141f
C19840 VPWR.t1380 VGND 0.01247f
C19841 VPWR.n1773 VGND 0.02783f
C19842 VPWR.n1774 VGND 0.01907f
C19843 VPWR.n1775 VGND 0.06276f
C19844 VPWR.n1776 VGND 0.09795f
C19845 VPWR.t2013 VGND 0.01141f
C19846 VPWR.t1250 VGND 0.01247f
C19847 VPWR.n1777 VGND 0.02783f
C19848 VPWR.n1778 VGND 0.01907f
C19849 VPWR.n1779 VGND 0.06274f
C19850 VPWR.n1780 VGND 0.05165f
C19851 VPWR.t1953 VGND 0.01141f
C19852 VPWR.t1418 VGND 0.01247f
C19853 VPWR.n1781 VGND 0.02783f
C19854 VPWR.n1782 VGND 0.01907f
C19855 VPWR.n1783 VGND 0.06276f
C19856 VPWR.n1784 VGND 0.09795f
C19857 VPWR.n1785 VGND 0.09221f
C19858 VPWR.n1786 VGND 0.066f
C19859 VPWR.n1787 VGND 0.05468f
C19860 VPWR.n1788 VGND 0.13984f
C19861 VPWR.n1789 VGND 0.01806f
C19862 VPWR.n1790 VGND 0.00732f
C19863 VPWR.n1791 VGND 0.10877f
C19864 VPWR.t1268 VGND 0.12017f
C19865 VPWR.t1251 VGND 0.07889f
C19866 VPWR.t1376 VGND 0.13401f
C19867 VPWR.n1792 VGND 0.07657f
C19868 VPWR.n1793 VGND 0.01806f
C19869 VPWR.n1794 VGND 0.13984f
C19870 VPWR.n1795 VGND 0.16543f
C19871 VPWR.n1796 VGND 1.02091f
C19872 VPWR.n1797 VGND 0.08393f
C19873 VPWR.n1798 VGND 0.08393f
C19874 VPWR.n1799 VGND 0.08393f
C19875 VPWR.n1800 VGND 0.08393f
C19876 VPWR.n1801 VGND 0.08393f
C19877 VPWR.n1802 VGND 0.08393f
C19878 VPWR.n1803 VGND 0.08393f
C19879 VPWR.n1804 VGND 0.08393f
C19880 VPWR.n1805 VGND 0.08393f
C19881 VPWR.n1806 VGND 0.08393f
C19882 VPWR.n1807 VGND 0.08393f
C19883 VPWR.n1808 VGND 0.08393f
C19884 VPWR.n1809 VGND 0.08393f
C19885 VPWR.n1810 VGND 0.08393f
C19886 VPWR.n1811 VGND 0.08393f
C19887 VPWR.n1812 VGND 0.19469f
C19888 VPWR.n1813 VGND 1.02091f
C19889 VPWR.n1814 VGND 1.02091f
C19890 VPWR.n1815 VGND 0.19469f
C19891 VPWR.n1816 VGND 0.13984f
C19892 VPWR.n1817 VGND 0.01806f
C19893 VPWR.n1818 VGND 0.07657f
C19894 VPWR.t1413 VGND 0.13401f
C19895 VPWR.t904 VGND 0.07889f
C19896 VPWR.t28 VGND 0.12017f
C19897 VPWR.n1819 VGND 0.10877f
C19898 VPWR.n1820 VGND 0.00732f
C19899 VPWR.n1821 VGND 0.01806f
C19900 VPWR.n1822 VGND 0.13984f
C19901 VPWR.n1823 VGND 0.08393f
C19902 VPWR.n1824 VGND 0.08393f
C19903 VPWR.n1825 VGND 0.13984f
C19904 VPWR.n1826 VGND 0.01806f
C19905 VPWR.n1827 VGND 0.00732f
C19906 VPWR.n1828 VGND 0.10877f
C19907 VPWR.t1046 VGND 0.09265f
C19908 VPWR.t858 VGND 0.07889f
C19909 VPWR.t1793 VGND 0.12017f
C19910 VPWR.n1829 VGND 0.10877f
C19911 VPWR.n1830 VGND 0.00732f
C19912 VPWR.n1831 VGND 0.01806f
C19913 VPWR.n1832 VGND 0.13984f
C19914 VPWR.n1833 VGND 0.08393f
C19915 VPWR.n1834 VGND 0.08393f
C19916 VPWR.n1835 VGND 0.13984f
C19917 VPWR.n1836 VGND 0.01806f
C19918 VPWR.n1837 VGND 0.00732f
C19919 VPWR.n1838 VGND 0.10877f
C19920 VPWR.t897 VGND 0.09265f
C19921 VPWR.t1028 VGND 0.07889f
C19922 VPWR.t1622 VGND 0.12017f
C19923 VPWR.n1839 VGND 0.10877f
C19924 VPWR.n1840 VGND 0.00732f
C19925 VPWR.n1841 VGND 0.01806f
C19926 VPWR.n1842 VGND 0.13984f
C19927 VPWR.n1843 VGND 0.08393f
C19928 VPWR.n1844 VGND 0.08393f
C19929 VPWR.n1845 VGND 0.13984f
C19930 VPWR.n1846 VGND 0.01806f
C19931 VPWR.n1847 VGND 0.00732f
C19932 VPWR.n1848 VGND 0.10877f
C19933 VPWR.t533 VGND 0.09265f
C19934 VPWR.t862 VGND 0.07889f
C19935 VPWR.t455 VGND 0.12017f
C19936 VPWR.n1849 VGND 0.10877f
C19937 VPWR.n1850 VGND 0.00732f
C19938 VPWR.n1851 VGND 0.01806f
C19939 VPWR.n1852 VGND 0.13984f
C19940 VPWR.n1853 VGND 0.08393f
C19941 VPWR.n1854 VGND 0.08393f
C19942 VPWR.n1855 VGND 0.13984f
C19943 VPWR.n1856 VGND 0.01806f
C19944 VPWR.n1857 VGND 0.00732f
C19945 VPWR.n1858 VGND 0.10877f
C19946 VPWR.t1705 VGND 0.09265f
C19947 VPWR.t906 VGND 0.07889f
C19948 VPWR.t267 VGND 0.12017f
C19949 VPWR.n1859 VGND 0.10877f
C19950 VPWR.n1860 VGND 0.00732f
C19951 VPWR.n1861 VGND 0.01806f
C19952 VPWR.n1862 VGND 0.13984f
C19953 VPWR.n1863 VGND 0.08393f
C19954 VPWR.n1864 VGND 0.08393f
C19955 VPWR.n1865 VGND 0.13984f
C19956 VPWR.n1866 VGND 0.01806f
C19957 VPWR.n1867 VGND 0.00732f
C19958 VPWR.n1868 VGND 0.10877f
C19959 VPWR.t805 VGND 0.09265f
C19960 VPWR.t861 VGND 0.07889f
C19961 VPWR.t978 VGND 0.12017f
C19962 VPWR.n1869 VGND 0.10877f
C19963 VPWR.n1870 VGND 0.00732f
C19964 VPWR.n1871 VGND 0.01806f
C19965 VPWR.n1872 VGND 0.13984f
C19966 VPWR.n1873 VGND 0.08393f
C19967 VPWR.n1874 VGND 0.08393f
C19968 VPWR.n1875 VGND 0.13984f
C19969 VPWR.n1876 VGND 0.01806f
C19970 VPWR.n1877 VGND 0.00732f
C19971 VPWR.n1878 VGND 0.10877f
C19972 VPWR.t318 VGND 0.09265f
C19973 VPWR.t1030 VGND 0.07889f
C19974 VPWR.t1489 VGND 0.12017f
C19975 VPWR.n1879 VGND 0.10877f
C19976 VPWR.n1880 VGND 0.00732f
C19977 VPWR.n1881 VGND 0.01806f
C19978 VPWR.n1882 VGND 0.13984f
C19979 VPWR.n1883 VGND 0.08393f
C19980 VPWR.n1884 VGND 0.08393f
C19981 VPWR.n1885 VGND 0.13984f
C19982 VPWR.n1886 VGND 0.01806f
C19983 VPWR.n1887 VGND 0.00732f
C19984 VPWR.n1888 VGND 0.10877f
C19985 VPWR.t705 VGND 0.09265f
C19986 VPWR.t903 VGND 0.07889f
C19987 VPWR.t435 VGND 0.12017f
C19988 VPWR.n1889 VGND 0.10877f
C19989 VPWR.n1890 VGND 0.00732f
C19990 VPWR.n1891 VGND 0.01806f
C19991 VPWR.n1892 VGND 0.13984f
C19992 VPWR.n1893 VGND 0.08393f
C19993 VPWR.n1894 VGND 1.01451f
C19994 VPWR.n1895 VGND 0.19469f
C19995 VPWR.n1896 VGND 0.08393f
C19996 VPWR.n1897 VGND 0.08393f
C19997 VPWR.n1898 VGND 0.08393f
C19998 VPWR.n1899 VGND 0.08393f
C19999 VPWR.n1900 VGND 0.08393f
C20000 VPWR.n1901 VGND 0.08393f
C20001 VPWR.n1902 VGND 0.08393f
C20002 VPWR.n1903 VGND 0.08393f
C20003 VPWR.n1904 VGND 0.08393f
C20004 VPWR.n1905 VGND 0.08393f
C20005 VPWR.n1906 VGND 0.08393f
C20006 VPWR.n1907 VGND 0.08393f
C20007 VPWR.n1908 VGND 0.08393f
C20008 VPWR.n1909 VGND 0.08393f
C20009 VPWR.n1910 VGND 0.08393f
C20010 VPWR.n1911 VGND 1.01451f
C20011 VPWR.n1912 VGND 1.01451f
C20012 VPWR.n1913 VGND 0.08393f
C20013 VPWR.n1914 VGND 0.13984f
C20014 VPWR.n1915 VGND 0.01806f
C20015 VPWR.n1916 VGND 0.00732f
C20016 VPWR.n1917 VGND 0.10877f
C20017 VPWR.t286 VGND 0.12017f
C20018 VPWR.t899 VGND 0.07889f
C20019 VPWR.t779 VGND 0.09265f
C20020 VPWR.t1911 VGND 0.07889f
C20021 VPWR.t724 VGND 0.12017f
C20022 VPWR.n1918 VGND 0.10877f
C20023 VPWR.n1919 VGND 0.00732f
C20024 VPWR.n1920 VGND 0.01806f
C20025 VPWR.n1921 VGND 0.13984f
C20026 VPWR.n1922 VGND 0.08393f
C20027 VPWR.n1923 VGND 0.08393f
C20028 VPWR.n1924 VGND 0.13984f
C20029 VPWR.n1925 VGND 0.01806f
C20030 VPWR.n1926 VGND 0.00732f
C20031 VPWR.n1927 VGND 0.10877f
C20032 VPWR.t1507 VGND 0.12017f
C20033 VPWR.t1910 VGND 0.07889f
C20034 VPWR.t1731 VGND 0.09265f
C20035 VPWR.t1906 VGND 0.07889f
C20036 VPWR.t1572 VGND 0.12017f
C20037 VPWR.n1928 VGND 0.10877f
C20038 VPWR.n1929 VGND 0.00732f
C20039 VPWR.n1930 VGND 0.01806f
C20040 VPWR.n1931 VGND 0.13984f
C20041 VPWR.n1932 VGND 0.08393f
C20042 VPWR.n1933 VGND 0.08393f
C20043 VPWR.n1934 VGND 0.13984f
C20044 VPWR.n1935 VGND 0.01806f
C20045 VPWR.n1936 VGND 0.00732f
C20046 VPWR.n1937 VGND 0.10877f
C20047 VPWR.t294 VGND 0.12017f
C20048 VPWR.t1570 VGND 0.07889f
C20049 VPWR.t801 VGND 0.09265f
C20050 VPWR.t1569 VGND 0.07889f
C20051 VPWR.t1679 VGND 0.12017f
C20052 VPWR.n1938 VGND 0.10877f
C20053 VPWR.n1939 VGND 0.00732f
C20054 VPWR.n1940 VGND 0.01806f
C20055 VPWR.n1941 VGND 0.13984f
C20056 VPWR.n1942 VGND 0.08393f
C20057 VPWR.n1943 VGND 0.08393f
C20058 VPWR.n1944 VGND 0.13984f
C20059 VPWR.n1945 VGND 0.01806f
C20060 VPWR.n1946 VGND 0.00732f
C20061 VPWR.n1947 VGND 0.10877f
C20062 VPWR.t185 VGND 0.12017f
C20063 VPWR.t902 VGND 0.07889f
C20064 VPWR.t461 VGND 0.09265f
C20065 VPWR.t901 VGND 0.07889f
C20066 VPWR.t418 VGND 0.12017f
C20067 VPWR.n1948 VGND 0.10877f
C20068 VPWR.n1949 VGND 0.00732f
C20069 VPWR.n1950 VGND 0.01806f
C20070 VPWR.n1951 VGND 0.13984f
C20071 VPWR.n1952 VGND 0.08393f
C20072 VPWR.n1953 VGND 0.08393f
C20073 VPWR.n1954 VGND 0.13984f
C20074 VPWR.n1955 VGND 0.01806f
C20075 VPWR.n1956 VGND 0.00732f
C20076 VPWR.n1957 VGND 0.10877f
C20077 VPWR.t1817 VGND 0.12017f
C20078 VPWR.t1571 VGND 0.07889f
C20079 VPWR.t1539 VGND 0.09265f
C20080 VPWR.t1909 VGND 0.07889f
C20081 VPWR.t1533 VGND 0.12017f
C20082 VPWR.n1958 VGND 0.10877f
C20083 VPWR.n1959 VGND 0.00732f
C20084 VPWR.n1960 VGND 0.01806f
C20085 VPWR.n1961 VGND 0.13984f
C20086 VPWR.n1962 VGND 0.08393f
C20087 VPWR.n1963 VGND 0.08393f
C20088 VPWR.n1964 VGND 0.13984f
C20089 VPWR.n1965 VGND 0.01806f
C20090 VPWR.n1966 VGND 0.00732f
C20091 VPWR.n1967 VGND 0.10877f
C20092 VPWR.t827 VGND 0.12017f
C20093 VPWR.t1908 VGND 0.07889f
C20094 VPWR.t1737 VGND 0.09265f
C20095 VPWR.t1568 VGND 0.07889f
C20096 VPWR.t1598 VGND 0.12017f
C20097 VPWR.n1968 VGND 0.10877f
C20098 VPWR.n1969 VGND 0.00732f
C20099 VPWR.n1970 VGND 0.01806f
C20100 VPWR.n1971 VGND 0.13984f
C20101 VPWR.n1972 VGND 0.08393f
C20102 VPWR.n1973 VGND 0.08393f
C20103 VPWR.n1974 VGND 0.13984f
C20104 VPWR.n1975 VGND 0.01806f
C20105 VPWR.n1976 VGND 0.00732f
C20106 VPWR.n1977 VGND 0.10877f
C20107 VPWR.t257 VGND 0.12017f
C20108 VPWR.t1567 VGND 0.07889f
C20109 VPWR.t1545 VGND 0.09265f
C20110 VPWR.t1566 VGND 0.07889f
C20111 VPWR.t358 VGND 0.12017f
C20112 VPWR.n1978 VGND 0.10877f
C20113 VPWR.n1979 VGND 0.00732f
C20114 VPWR.n1980 VGND 0.01806f
C20115 VPWR.n1981 VGND 0.13984f
C20116 VPWR.n1982 VGND 0.08393f
C20117 VPWR.n1983 VGND 0.08393f
C20118 VPWR.n1984 VGND 0.13984f
C20119 VPWR.n1985 VGND 0.01806f
C20120 VPWR.n1986 VGND 0.00732f
C20121 VPWR.n1987 VGND 0.10877f
C20122 VPWR.t1717 VGND 0.12017f
C20123 VPWR.t900 VGND 0.07889f
C20124 VPWR.t1121 VGND 0.13401f
C20125 VPWR.n1988 VGND 0.07657f
C20126 VPWR.n1989 VGND 0.01806f
C20127 VPWR.n1990 VGND 0.13984f
C20128 VPWR.n1991 VGND 0.19469f
C20129 VPWR.n1992 VGND 1.02091f
C20130 VPWR.n1993 VGND 0.08393f
C20131 VPWR.n1994 VGND 0.08393f
C20132 VPWR.n1995 VGND 0.08393f
C20133 VPWR.n1996 VGND 0.08393f
C20134 VPWR.n1997 VGND 0.08393f
C20135 VPWR.n1998 VGND 0.08393f
C20136 VPWR.n1999 VGND 0.08393f
C20137 VPWR.n2000 VGND 0.08393f
C20138 VPWR.n2001 VGND 0.08393f
C20139 VPWR.n2002 VGND 0.08393f
C20140 VPWR.n2003 VGND 0.08393f
C20141 VPWR.n2004 VGND 0.08393f
C20142 VPWR.n2005 VGND 0.08393f
C20143 VPWR.n2006 VGND 0.08393f
C20144 VPWR.n2007 VGND 0.08393f
C20145 VPWR.n2008 VGND 0.19469f
C20146 VPWR.n2009 VGND 1.02091f
C20147 VPWR.n2010 VGND 1.02091f
C20148 VPWR.n2011 VGND 0.19469f
C20149 VPWR.n2012 VGND 0.13984f
C20150 VPWR.n2013 VGND 0.01806f
C20151 VPWR.n2014 VGND 0.07657f
C20152 VPWR.t1193 VGND 0.13401f
C20153 VPWR.t1032 VGND 0.07889f
C20154 VPWR.t1060 VGND 0.12017f
C20155 VPWR.n2015 VGND 0.10877f
C20156 VPWR.n2016 VGND 0.00732f
C20157 VPWR.n2017 VGND 0.01806f
C20158 VPWR.n2018 VGND 0.13984f
C20159 VPWR.n2019 VGND 0.08393f
C20160 VPWR.n2020 VGND 0.08393f
C20161 VPWR.n2021 VGND 0.13984f
C20162 VPWR.n2022 VGND 0.01806f
C20163 VPWR.n2023 VGND 0.00732f
C20164 VPWR.n2024 VGND 0.10877f
C20165 VPWR.t588 VGND 0.09265f
C20166 VPWR.t987 VGND 0.07889f
C20167 VPWR.t245 VGND 0.12017f
C20168 VPWR.n2025 VGND 0.10877f
C20169 VPWR.n2026 VGND 0.00732f
C20170 VPWR.n2027 VGND 0.01806f
C20171 VPWR.n2028 VGND 0.13984f
C20172 VPWR.n2029 VGND 0.08393f
C20173 VPWR.n2030 VGND 0.08393f
C20174 VPWR.n2031 VGND 0.13984f
C20175 VPWR.n2032 VGND 0.01806f
C20176 VPWR.n2033 VGND 0.00732f
C20177 VPWR.n2034 VGND 0.10877f
C20178 VPWR.t1594 VGND 0.09265f
C20179 VPWR.t982 VGND 0.07889f
C20180 VPWR.t1914 VGND 0.12017f
C20181 VPWR.n2035 VGND 0.10877f
C20182 VPWR.n2036 VGND 0.00732f
C20183 VPWR.n2037 VGND 0.01806f
C20184 VPWR.n2038 VGND 0.13984f
C20185 VPWR.n2039 VGND 0.08393f
C20186 VPWR.n2040 VGND 0.08393f
C20187 VPWR.n2041 VGND 0.13984f
C20188 VPWR.n2042 VGND 0.01806f
C20189 VPWR.n2043 VGND 0.00732f
C20190 VPWR.n2044 VGND 0.10877f
C20191 VPWR.t1529 VGND 0.09265f
C20192 VPWR.t1040 VGND 0.07889f
C20193 VPWR.t863 VGND 0.12017f
C20194 VPWR.n2045 VGND 0.10877f
C20195 VPWR.n2046 VGND 0.00732f
C20196 VPWR.n2047 VGND 0.01806f
C20197 VPWR.n2048 VGND 0.13984f
C20198 VPWR.n2049 VGND 0.08393f
C20199 VPWR.n2050 VGND 0.08393f
C20200 VPWR.n2051 VGND 0.13984f
C20201 VPWR.n2052 VGND 0.01806f
C20202 VPWR.n2053 VGND 0.00732f
C20203 VPWR.n2054 VGND 0.10877f
C20204 VPWR.t147 VGND 0.09265f
C20205 VPWR.t1034 VGND 0.07889f
C20206 VPWR.t306 VGND 0.12017f
C20207 VPWR.n2055 VGND 0.10877f
C20208 VPWR.n2056 VGND 0.00732f
C20209 VPWR.n2057 VGND 0.01806f
C20210 VPWR.n2058 VGND 0.13984f
C20211 VPWR.n2059 VGND 0.08393f
C20212 VPWR.n2060 VGND 0.08393f
C20213 VPWR.n2061 VGND 0.13984f
C20214 VPWR.n2062 VGND 0.01806f
C20215 VPWR.n2063 VGND 0.00732f
C20216 VPWR.n2064 VGND 0.10877f
C20217 VPWR.t1675 VGND 0.09265f
C20218 VPWR.t1039 VGND 0.07889f
C20219 VPWR.t855 VGND 0.12017f
C20220 VPWR.n2065 VGND 0.10877f
C20221 VPWR.n2066 VGND 0.00732f
C20222 VPWR.n2067 VGND 0.01806f
C20223 VPWR.n2068 VGND 0.13984f
C20224 VPWR.n2069 VGND 0.08393f
C20225 VPWR.n2070 VGND 0.08393f
C20226 VPWR.n2071 VGND 0.13984f
C20227 VPWR.n2072 VGND 0.01806f
C20228 VPWR.n2073 VGND 0.00732f
C20229 VPWR.n2074 VGND 0.10877f
C20230 VPWR.t129 VGND 0.09265f
C20231 VPWR.t984 VGND 0.07889f
C20232 VPWR.t1515 VGND 0.12017f
C20233 VPWR.n2075 VGND 0.10877f
C20234 VPWR.n2076 VGND 0.00732f
C20235 VPWR.n2077 VGND 0.01806f
C20236 VPWR.n2078 VGND 0.13984f
C20237 VPWR.n2079 VGND 0.08393f
C20238 VPWR.n2080 VGND 0.08393f
C20239 VPWR.n2081 VGND 0.13984f
C20240 VPWR.n2082 VGND 0.01806f
C20241 VPWR.n2083 VGND 0.00732f
C20242 VPWR.n2084 VGND 0.10877f
C20243 VPWR.t1840 VGND 0.09265f
C20244 VPWR.t1041 VGND 0.07889f
C20245 VPWR.t819 VGND 0.12017f
C20246 VPWR.n2085 VGND 0.10877f
C20247 VPWR.n2086 VGND 0.00732f
C20248 VPWR.n2087 VGND 0.01806f
C20249 VPWR.n2088 VGND 0.13984f
C20250 VPWR.n2089 VGND 0.08393f
C20251 VPWR.n2090 VGND 1.01451f
C20252 VPWR.n2091 VGND 0.19469f
C20253 VPWR.n2092 VGND 0.08393f
C20254 VPWR.n2093 VGND 0.08393f
C20255 VPWR.n2094 VGND 0.08393f
C20256 VPWR.n2095 VGND 0.08393f
C20257 VPWR.n2096 VGND 0.08393f
C20258 VPWR.n2097 VGND 0.08393f
C20259 VPWR.n2098 VGND 0.08393f
C20260 VPWR.n2099 VGND 0.08393f
C20261 VPWR.n2100 VGND 0.08393f
C20262 VPWR.n2101 VGND 0.08393f
C20263 VPWR.n2102 VGND 0.08393f
C20264 VPWR.n2103 VGND 0.08393f
C20265 VPWR.n2104 VGND 0.08393f
C20266 VPWR.n2105 VGND 0.08393f
C20267 VPWR.n2106 VGND 0.08393f
C20268 VPWR.n2107 VGND 1.01451f
C20269 VPWR.n2108 VGND 1.01451f
C20270 VPWR.n2109 VGND 0.08393f
C20271 VPWR.n2110 VGND 0.13984f
C20272 VPWR.n2111 VGND 0.01806f
C20273 VPWR.n2112 VGND 0.00732f
C20274 VPWR.n2113 VGND 0.10877f
C20275 VPWR.t284 VGND 0.12017f
C20276 VPWR.t841 VGND 0.07889f
C20277 VPWR.t728 VGND 0.09265f
C20278 VPWR.t1648 VGND 0.07889f
C20279 VPWR.t722 VGND 0.12017f
C20280 VPWR.n2114 VGND 0.10877f
C20281 VPWR.n2115 VGND 0.00732f
C20282 VPWR.n2116 VGND 0.01806f
C20283 VPWR.n2117 VGND 0.13984f
C20284 VPWR.n2118 VGND 0.08393f
C20285 VPWR.n2119 VGND 0.08393f
C20286 VPWR.n2120 VGND 0.13984f
C20287 VPWR.n2121 VGND 0.01806f
C20288 VPWR.n2122 VGND 0.00732f
C20289 VPWR.n2123 VGND 0.10877f
C20290 VPWR.t1509 VGND 0.12017f
C20291 VPWR.t1593 VGND 0.07889f
C20292 VPWR.t1727 VGND 0.09265f
C20293 VPWR.t445 VGND 0.07889f
C20294 VPWR.t1815 VGND 0.12017f
C20295 VPWR.n2124 VGND 0.10877f
C20296 VPWR.n2125 VGND 0.00732f
C20297 VPWR.n2126 VGND 0.01806f
C20298 VPWR.n2127 VGND 0.13984f
C20299 VPWR.n2128 VGND 0.08393f
C20300 VPWR.n2129 VGND 0.08393f
C20301 VPWR.n2130 VGND 0.13984f
C20302 VPWR.n2131 VGND 0.01806f
C20303 VPWR.n2132 VGND 0.00732f
C20304 VPWR.n2133 VGND 0.10877f
C20305 VPWR.t1075 VGND 0.12017f
C20306 VPWR.t116 VGND 0.07889f
C20307 VPWR.t799 VGND 0.09265f
C20308 VPWR.t115 VGND 0.07889f
C20309 VPWR.t1677 VGND 0.12017f
C20310 VPWR.n2134 VGND 0.10877f
C20311 VPWR.n2135 VGND 0.00732f
C20312 VPWR.n2136 VGND 0.01806f
C20313 VPWR.n2137 VGND 0.13984f
C20314 VPWR.n2138 VGND 0.08393f
C20315 VPWR.n2139 VGND 0.08393f
C20316 VPWR.n2140 VGND 0.13984f
C20317 VPWR.n2141 VGND 0.01806f
C20318 VPWR.n2142 VGND 0.00732f
C20319 VPWR.n2143 VGND 0.10877f
C20320 VPWR.t310 VGND 0.12017f
C20321 VPWR.t444 VGND 0.07889f
C20322 VPWR.t459 VGND 0.09265f
C20323 VPWR.t443 VGND 0.07889f
C20324 VPWR.t416 VGND 0.12017f
C20325 VPWR.n2144 VGND 0.10877f
C20326 VPWR.n2145 VGND 0.00732f
C20327 VPWR.n2146 VGND 0.01806f
C20328 VPWR.n2147 VGND 0.13984f
C20329 VPWR.n2148 VGND 0.08393f
C20330 VPWR.n2149 VGND 0.08393f
C20331 VPWR.n2150 VGND 0.13984f
C20332 VPWR.n2151 VGND 0.01806f
C20333 VPWR.n2152 VGND 0.00732f
C20334 VPWR.n2153 VGND 0.10877f
C20335 VPWR.t867 VGND 0.12017f
C20336 VPWR.t117 VGND 0.07889f
C20337 VPWR.t1537 VGND 0.09265f
C20338 VPWR.t1592 VGND 0.07889f
C20339 VPWR.t1531 VGND 0.12017f
C20340 VPWR.n2154 VGND 0.10877f
C20341 VPWR.n2155 VGND 0.00732f
C20342 VPWR.n2156 VGND 0.01806f
C20343 VPWR.n2157 VGND 0.13984f
C20344 VPWR.n2158 VGND 0.08393f
C20345 VPWR.n2159 VGND 0.08393f
C20346 VPWR.n2160 VGND 0.13984f
C20347 VPWR.n2161 VGND 0.01806f
C20348 VPWR.n2162 VGND 0.00732f
C20349 VPWR.n2163 VGND 0.10877f
C20350 VPWR.t825 VGND 0.12017f
C20351 VPWR.t1591 VGND 0.07889f
C20352 VPWR.t1735 VGND 0.09265f
C20353 VPWR.t114 VGND 0.07889f
C20354 VPWR.t1596 VGND 0.12017f
C20355 VPWR.n2164 VGND 0.10877f
C20356 VPWR.n2165 VGND 0.00732f
C20357 VPWR.n2166 VGND 0.01806f
C20358 VPWR.n2167 VGND 0.13984f
C20359 VPWR.n2168 VGND 0.08393f
C20360 VPWR.n2169 VGND 0.08393f
C20361 VPWR.n2170 VGND 0.13984f
C20362 VPWR.n2171 VGND 0.01806f
C20363 VPWR.n2172 VGND 0.00732f
C20364 VPWR.n2173 VGND 0.10877f
C20365 VPWR.t255 VGND 0.12017f
C20366 VPWR.t1650 VGND 0.07889f
C20367 VPWR.t1543 VGND 0.09265f
C20368 VPWR.t1649 VGND 0.07889f
C20369 VPWR.t356 VGND 0.12017f
C20370 VPWR.n2174 VGND 0.10877f
C20371 VPWR.n2175 VGND 0.00732f
C20372 VPWR.n2176 VGND 0.01806f
C20373 VPWR.n2177 VGND 0.13984f
C20374 VPWR.n2178 VGND 0.08393f
C20375 VPWR.n2179 VGND 0.08393f
C20376 VPWR.n2180 VGND 0.13984f
C20377 VPWR.n2181 VGND 0.01806f
C20378 VPWR.n2182 VGND 0.00732f
C20379 VPWR.n2183 VGND 0.10877f
C20380 VPWR.t1715 VGND 0.12017f
C20381 VPWR.t842 VGND 0.07889f
C20382 VPWR.t1126 VGND 0.13401f
C20383 VPWR.n2184 VGND 0.07657f
C20384 VPWR.n2185 VGND 0.01806f
C20385 VPWR.n2186 VGND 0.13984f
C20386 VPWR.n2187 VGND 0.19469f
C20387 VPWR.n2188 VGND 1.02091f
C20388 VPWR.n2189 VGND 0.08393f
C20389 VPWR.n2190 VGND 0.08393f
C20390 VPWR.n2191 VGND 0.08393f
C20391 VPWR.n2192 VGND 0.08393f
C20392 VPWR.n2193 VGND 0.08393f
C20393 VPWR.n2194 VGND 0.08393f
C20394 VPWR.n2195 VGND 0.08393f
C20395 VPWR.n2196 VGND 0.08393f
C20396 VPWR.n2197 VGND 0.08393f
C20397 VPWR.n2198 VGND 0.08393f
C20398 VPWR.n2199 VGND 0.08393f
C20399 VPWR.n2200 VGND 0.08393f
C20400 VPWR.n2201 VGND 0.08393f
C20401 VPWR.n2202 VGND 0.08393f
C20402 VPWR.n2203 VGND 0.08393f
C20403 VPWR.n2204 VGND 0.19469f
C20404 VPWR.n2205 VGND 1.02091f
C20405 VPWR.n2206 VGND 1.02091f
C20406 VPWR.n2207 VGND 0.19469f
C20407 VPWR.n2208 VGND 0.13984f
C20408 VPWR.n2209 VGND 0.01806f
C20409 VPWR.n2210 VGND 0.07657f
C20410 VPWR.t1292 VGND 0.13401f
C20411 VPWR.t1883 VGND 0.07889f
C20412 VPWR.t225 VGND 0.12017f
C20413 VPWR.n2211 VGND 0.10877f
C20414 VPWR.n2212 VGND 0.00732f
C20415 VPWR.n2213 VGND 0.01806f
C20416 VPWR.n2214 VGND 0.13984f
C20417 VPWR.n2215 VGND 0.08393f
C20418 VPWR.n2216 VGND 0.08393f
C20419 VPWR.n2217 VGND 0.13984f
C20420 VPWR.n2218 VGND 0.01806f
C20421 VPWR.n2219 VGND 0.00732f
C20422 VPWR.n2220 VGND 0.10877f
C20423 VPWR.t1054 VGND 0.09265f
C20424 VPWR.t1657 VGND 0.07889f
C20425 VPWR.t877 VGND 0.12017f
C20426 VPWR.n2221 VGND 0.10877f
C20427 VPWR.n2222 VGND 0.00732f
C20428 VPWR.n2223 VGND 0.01806f
C20429 VPWR.n2224 VGND 0.13984f
C20430 VPWR.n2225 VGND 0.08393f
C20431 VPWR.n2226 VGND 0.08393f
C20432 VPWR.n2227 VGND 0.13984f
C20433 VPWR.n2228 VGND 0.01806f
C20434 VPWR.n2229 VGND 0.00732f
C20435 VPWR.n2230 VGND 0.10877f
C20436 VPWR.t1003 VGND 0.09265f
C20437 VPWR.t1922 VGND 0.07889f
C20438 VPWR.t392 VGND 0.12017f
C20439 VPWR.n2231 VGND 0.10877f
C20440 VPWR.n2232 VGND 0.00732f
C20441 VPWR.n2233 VGND 0.01806f
C20442 VPWR.n2234 VGND 0.13984f
C20443 VPWR.n2235 VGND 0.08393f
C20444 VPWR.n2236 VGND 0.08393f
C20445 VPWR.n2237 VGND 0.13984f
C20446 VPWR.n2238 VGND 0.01806f
C20447 VPWR.n2239 VGND 0.00732f
C20448 VPWR.n2240 VGND 0.10877f
C20449 VPWR.t60 VGND 0.09265f
C20450 VPWR.t1661 VGND 0.07889f
C20451 VPWR.t139 VGND 0.12017f
C20452 VPWR.n2241 VGND 0.10877f
C20453 VPWR.n2242 VGND 0.00732f
C20454 VPWR.n2243 VGND 0.01806f
C20455 VPWR.n2244 VGND 0.13984f
C20456 VPWR.n2245 VGND 0.08393f
C20457 VPWR.n2246 VGND 0.08393f
C20458 VPWR.n2247 VGND 0.13984f
C20459 VPWR.n2248 VGND 0.01806f
C20460 VPWR.n2249 VGND 0.00732f
C20461 VPWR.n2250 VGND 0.10877f
C20462 VPWR.t161 VGND 0.09265f
C20463 VPWR.t1885 VGND 0.07889f
C20464 VPWR.t4 VGND 0.12017f
C20465 VPWR.n2251 VGND 0.10877f
C20466 VPWR.n2252 VGND 0.00732f
C20467 VPWR.n2253 VGND 0.01806f
C20468 VPWR.n2254 VGND 0.13984f
C20469 VPWR.n2255 VGND 0.08393f
C20470 VPWR.n2256 VGND 0.08393f
C20471 VPWR.n2257 VGND 0.13984f
C20472 VPWR.n2258 VGND 0.01806f
C20473 VPWR.n2259 VGND 0.00732f
C20474 VPWR.n2260 VGND 0.10877f
C20475 VPWR.t1761 VGND 0.09265f
C20476 VPWR.t1660 VGND 0.07889f
C20477 VPWR.t1874 VGND 0.12017f
C20478 VPWR.n2261 VGND 0.10877f
C20479 VPWR.n2262 VGND 0.00732f
C20480 VPWR.n2263 VGND 0.01806f
C20481 VPWR.n2264 VGND 0.13984f
C20482 VPWR.n2265 VGND 0.08393f
C20483 VPWR.n2266 VGND 0.08393f
C20484 VPWR.n2267 VGND 0.13984f
C20485 VPWR.n2268 VGND 0.01806f
C20486 VPWR.n2269 VGND 0.00732f
C20487 VPWR.n2270 VGND 0.10877f
C20488 VPWR.t1811 VGND 0.09265f
C20489 VPWR.t1654 VGND 0.07889f
C20490 VPWR.t1473 VGND 0.12017f
C20491 VPWR.n2271 VGND 0.10877f
C20492 VPWR.n2272 VGND 0.00732f
C20493 VPWR.n2273 VGND 0.01806f
C20494 VPWR.n2274 VGND 0.13984f
C20495 VPWR.n2275 VGND 0.08393f
C20496 VPWR.n2276 VGND 0.08393f
C20497 VPWR.n2277 VGND 0.13984f
C20498 VPWR.n2278 VGND 0.01806f
C20499 VPWR.n2279 VGND 0.00732f
C20500 VPWR.n2280 VGND 0.10877f
C20501 VPWR.t1586 VGND 0.09265f
C20502 VPWR.t1882 VGND 0.07889f
C20503 VPWR.t1557 VGND 0.12017f
C20504 VPWR.n2281 VGND 0.10877f
C20505 VPWR.n2282 VGND 0.00732f
C20506 VPWR.n2283 VGND 0.01806f
C20507 VPWR.n2284 VGND 0.13984f
C20508 VPWR.n2285 VGND 0.08393f
C20509 VPWR.n2286 VGND 1.01451f
C20510 VPWR.n2287 VGND 0.19469f
C20511 VPWR.n2288 VGND 0.08393f
C20512 VPWR.n2289 VGND 0.08393f
C20513 VPWR.n2290 VGND 0.08393f
C20514 VPWR.n2291 VGND 0.08393f
C20515 VPWR.n2292 VGND 0.08393f
C20516 VPWR.n2293 VGND 0.08393f
C20517 VPWR.n2294 VGND 0.08393f
C20518 VPWR.n2295 VGND 0.08393f
C20519 VPWR.n2296 VGND 0.08393f
C20520 VPWR.n2297 VGND 0.08393f
C20521 VPWR.n2298 VGND 0.08393f
C20522 VPWR.n2299 VGND 0.08393f
C20523 VPWR.n2300 VGND 0.08393f
C20524 VPWR.n2301 VGND 0.08393f
C20525 VPWR.n2302 VGND 0.08393f
C20526 VPWR.n2303 VGND 1.01451f
C20527 VPWR.n2304 VGND 1.01451f
C20528 VPWR.n2305 VGND 0.08393f
C20529 VPWR.n2306 VGND 0.13984f
C20530 VPWR.n2307 VGND 0.01806f
C20531 VPWR.n2308 VGND 0.00732f
C20532 VPWR.n2309 VGND 0.10877f
C20533 VPWR.t1842 VGND 0.12017f
C20534 VPWR.t1651 VGND 0.07889f
C20535 VPWR.t1836 VGND 0.09265f
C20536 VPWR.t1647 VGND 0.07889f
C20537 VPWR.t913 VGND 0.12017f
C20538 VPWR.n2310 VGND 0.10877f
C20539 VPWR.n2311 VGND 0.00732f
C20540 VPWR.n2312 VGND 0.01806f
C20541 VPWR.n2313 VGND 0.13984f
C20542 VPWR.n2314 VGND 0.08393f
C20543 VPWR.n2315 VGND 0.08393f
C20544 VPWR.n2316 VGND 0.13984f
C20545 VPWR.n2317 VGND 0.01806f
C20546 VPWR.n2318 VGND 0.00732f
C20547 VPWR.n2319 VGND 0.10877f
C20548 VPWR.t1519 VGND 0.12017f
C20549 VPWR.t1646 VGND 0.07889f
C20550 VPWR.t127 VGND 0.09265f
C20551 VPWR.t401 VGND 0.07889f
C20552 VPWR.t153 VGND 0.12017f
C20553 VPWR.n2320 VGND 0.10877f
C20554 VPWR.n2321 VGND 0.00732f
C20555 VPWR.n2322 VGND 0.01806f
C20556 VPWR.n2323 VGND 0.13984f
C20557 VPWR.n2324 VGND 0.08393f
C20558 VPWR.n2325 VGND 0.08393f
C20559 VPWR.n2326 VGND 0.13984f
C20560 VPWR.n2327 VGND 0.01806f
C20561 VPWR.n2328 VGND 0.00732f
C20562 VPWR.n2329 VGND 0.10877f
C20563 VPWR.t849 VGND 0.12017f
C20564 VPWR.t1866 VGND 0.07889f
C20565 VPWR.t948 VGND 0.09265f
C20566 VPWR.t1865 VGND 0.07889f
C20567 VPWR.t944 VGND 0.12017f
C20568 VPWR.n2330 VGND 0.10877f
C20569 VPWR.n2331 VGND 0.00732f
C20570 VPWR.n2332 VGND 0.01806f
C20571 VPWR.n2333 VGND 0.13984f
C20572 VPWR.n2334 VGND 0.08393f
C20573 VPWR.n2335 VGND 0.08393f
C20574 VPWR.n2336 VGND 0.13984f
C20575 VPWR.n2337 VGND 0.01806f
C20576 VPWR.n2338 VGND 0.00732f
C20577 VPWR.n2339 VGND 0.10877f
C20578 VPWR.t300 VGND 0.12017f
C20579 VPWR.t400 VGND 0.07889f
C20580 VPWR.t213 VGND 0.09265f
C20581 VPWR.t103 VGND 0.07889f
C20582 VPWR.t457 VGND 0.12017f
C20583 VPWR.n2340 VGND 0.10877f
C20584 VPWR.n2341 VGND 0.00732f
C20585 VPWR.n2342 VGND 0.01806f
C20586 VPWR.n2343 VGND 0.13984f
C20587 VPWR.n2344 VGND 0.08393f
C20588 VPWR.n2345 VGND 0.08393f
C20589 VPWR.n2346 VGND 0.13984f
C20590 VPWR.n2347 VGND 0.01806f
C20591 VPWR.n2348 VGND 0.00732f
C20592 VPWR.n2349 VGND 0.10877f
C20593 VPWR.t407 VGND 0.12017f
C20594 VPWR.t1867 VGND 0.07889f
C20595 VPWR.t72 VGND 0.09265f
C20596 VPWR.t1645 VGND 0.07889f
C20597 VPWR.t64 VGND 0.12017f
C20598 VPWR.n2350 VGND 0.10877f
C20599 VPWR.n2351 VGND 0.00732f
C20600 VPWR.n2352 VGND 0.01806f
C20601 VPWR.n2353 VGND 0.13984f
C20602 VPWR.n2354 VGND 0.08393f
C20603 VPWR.n2355 VGND 0.08393f
C20604 VPWR.n2356 VGND 0.13984f
C20605 VPWR.n2357 VGND 0.01806f
C20606 VPWR.n2358 VGND 0.00732f
C20607 VPWR.n2359 VGND 0.10877f
C20608 VPWR.t643 VGND 0.12017f
C20609 VPWR.t1644 VGND 0.07889f
C20610 VPWR.t209 VGND 0.09265f
C20611 VPWR.t1864 VGND 0.07889f
C20612 VPWR.t1007 VGND 0.12017f
C20613 VPWR.n2360 VGND 0.10877f
C20614 VPWR.n2361 VGND 0.00732f
C20615 VPWR.n2362 VGND 0.01806f
C20616 VPWR.n2363 VGND 0.13984f
C20617 VPWR.n2364 VGND 0.08393f
C20618 VPWR.n2365 VGND 0.08393f
C20619 VPWR.n2366 VGND 0.13984f
C20620 VPWR.n2367 VGND 0.01806f
C20621 VPWR.n2368 VGND 0.00732f
C20622 VPWR.n2369 VGND 0.10877f
C20623 VPWR.t98 VGND 0.12017f
C20624 VPWR.t1863 VGND 0.07889f
C20625 VPWR.t586 VGND 0.09265f
C20626 VPWR.t1862 VGND 0.07889f
C20627 VPWR.t1549 VGND 0.12017f
C20628 VPWR.n2370 VGND 0.10877f
C20629 VPWR.n2371 VGND 0.00732f
C20630 VPWR.n2372 VGND 0.01806f
C20631 VPWR.n2373 VGND 0.13984f
C20632 VPWR.n2374 VGND 0.08393f
C20633 VPWR.n2375 VGND 0.08393f
C20634 VPWR.n2376 VGND 0.13984f
C20635 VPWR.n2377 VGND 0.01806f
C20636 VPWR.n2378 VGND 0.00732f
C20637 VPWR.n2379 VGND 0.10877f
C20638 VPWR.t1058 VGND 0.12017f
C20639 VPWR.t1652 VGND 0.07889f
C20640 VPWR.t1225 VGND 0.13401f
C20641 VPWR.n2380 VGND 0.07657f
C20642 VPWR.n2381 VGND 0.01806f
C20643 VPWR.n2382 VGND 0.13984f
C20644 VPWR.n2383 VGND 0.19469f
C20645 VPWR.n2384 VGND 1.02091f
C20646 VPWR.n2385 VGND 0.08393f
C20647 VPWR.n2386 VGND 0.08393f
C20648 VPWR.n2387 VGND 0.08393f
C20649 VPWR.n2388 VGND 0.08393f
C20650 VPWR.n2389 VGND 0.08393f
C20651 VPWR.n2390 VGND 0.08393f
C20652 VPWR.n2391 VGND 0.08393f
C20653 VPWR.n2392 VGND 0.08393f
C20654 VPWR.n2393 VGND 0.08393f
C20655 VPWR.n2394 VGND 0.08393f
C20656 VPWR.n2395 VGND 0.08393f
C20657 VPWR.n2396 VGND 0.08393f
C20658 VPWR.n2397 VGND 0.08393f
C20659 VPWR.n2398 VGND 0.08393f
C20660 VPWR.n2399 VGND 0.08393f
C20661 VPWR.n2400 VGND 0.19469f
C20662 VPWR.n2401 VGND 1.02091f
C20663 VPWR.n2402 VGND 1.02091f
C20664 VPWR.n2403 VGND 0.19469f
C20665 VPWR.n2404 VGND 0.13984f
C20666 VPWR.n2405 VGND 0.01806f
C20667 VPWR.n2406 VGND 0.07657f
C20668 VPWR.t1395 VGND 0.13401f
C20669 VPWR.t345 VGND 0.07889f
C20670 VPWR.t167 VGND 0.12017f
C20671 VPWR.n2407 VGND 0.10877f
C20672 VPWR.n2408 VGND 0.00732f
C20673 VPWR.n2409 VGND 0.01806f
C20674 VPWR.n2410 VGND 0.13984f
C20675 VPWR.n2411 VGND 0.08393f
C20676 VPWR.n2412 VGND 0.08393f
C20677 VPWR.n2413 VGND 0.13984f
C20678 VPWR.n2414 VGND 0.01806f
C20679 VPWR.n2415 VGND 0.00732f
C20680 VPWR.n2416 VGND 0.10877f
C20681 VPWR.t1021 VGND 0.09265f
C20682 VPWR.t814 VGND 0.07889f
C20683 VPWR.t1797 VGND 0.12017f
C20684 VPWR.n2417 VGND 0.10877f
C20685 VPWR.n2418 VGND 0.00732f
C20686 VPWR.n2419 VGND 0.01806f
C20687 VPWR.n2420 VGND 0.13984f
C20688 VPWR.n2421 VGND 0.08393f
C20689 VPWR.n2422 VGND 0.08393f
C20690 VPWR.n2423 VGND 0.13984f
C20691 VPWR.n2424 VGND 0.01806f
C20692 VPWR.n2425 VGND 0.00732f
C20693 VPWR.n2426 VGND 0.10877f
C20694 VPWR.t993 VGND 0.09265f
C20695 VPWR.t932 VGND 0.07889f
C20696 VPWR.t1628 VGND 0.12017f
C20697 VPWR.n2427 VGND 0.10877f
C20698 VPWR.n2428 VGND 0.00732f
C20699 VPWR.n2429 VGND 0.01806f
C20700 VPWR.n2430 VGND 0.13984f
C20701 VPWR.n2431 VGND 0.08393f
C20702 VPWR.n2432 VGND 0.08393f
C20703 VPWR.n2433 VGND 0.13984f
C20704 VPWR.n2434 VGND 0.01806f
C20705 VPWR.n2435 VGND 0.00732f
C20706 VPWR.n2436 VGND 0.10877f
C20707 VPWR.t537 VGND 0.09265f
C20708 VPWR.t818 VGND 0.07889f
C20709 VPWR.t661 VGND 0.12017f
C20710 VPWR.n2437 VGND 0.10877f
C20711 VPWR.n2438 VGND 0.00732f
C20712 VPWR.n2439 VGND 0.01806f
C20713 VPWR.n2440 VGND 0.13984f
C20714 VPWR.n2441 VGND 0.08393f
C20715 VPWR.n2442 VGND 0.08393f
C20716 VPWR.n2443 VGND 0.13984f
C20717 VPWR.n2444 VGND 0.01806f
C20718 VPWR.n2445 VGND 0.00732f
C20719 VPWR.n2446 VGND 0.10877f
C20720 VPWR.t199 VGND 0.09265f
C20721 VPWR.t347 VGND 0.07889f
C20722 VPWR.t273 VGND 0.12017f
C20723 VPWR.n2447 VGND 0.10877f
C20724 VPWR.n2448 VGND 0.00732f
C20725 VPWR.n2449 VGND 0.01806f
C20726 VPWR.n2450 VGND 0.13984f
C20727 VPWR.n2451 VGND 0.08393f
C20728 VPWR.n2452 VGND 0.08393f
C20729 VPWR.n2453 VGND 0.13984f
C20730 VPWR.n2454 VGND 0.01806f
C20731 VPWR.n2455 VGND 0.00732f
C20732 VPWR.n2456 VGND 0.10877f
C20733 VPWR.t809 VGND 0.09265f
C20734 VPWR.t817 VGND 0.07889f
C20735 VPWR.t750 VGND 0.12017f
C20736 VPWR.n2457 VGND 0.10877f
C20737 VPWR.n2458 VGND 0.00732f
C20738 VPWR.n2459 VGND 0.01806f
C20739 VPWR.n2460 VGND 0.13984f
C20740 VPWR.n2461 VGND 0.08393f
C20741 VPWR.n2462 VGND 0.08393f
C20742 VPWR.n2463 VGND 0.13984f
C20743 VPWR.n2464 VGND 0.01806f
C20744 VPWR.n2465 VGND 0.00732f
C20745 VPWR.n2466 VGND 0.10877f
C20746 VPWR.t324 VGND 0.09265f
C20747 VPWR.t934 VGND 0.07889f
C20748 VPWR.t1485 VGND 0.12017f
C20749 VPWR.n2467 VGND 0.10877f
C20750 VPWR.n2468 VGND 0.00732f
C20751 VPWR.n2469 VGND 0.01806f
C20752 VPWR.n2470 VGND 0.13984f
C20753 VPWR.n2471 VGND 0.08393f
C20754 VPWR.n2472 VGND 0.08393f
C20755 VPWR.n2473 VGND 0.13984f
C20756 VPWR.n2474 VGND 0.01806f
C20757 VPWR.n2475 VGND 0.00732f
C20758 VPWR.n2476 VGND 0.10877f
C20759 VPWR.t707 VGND 0.09265f
C20760 VPWR.t344 VGND 0.07889f
C20761 VPWR.t1743 VGND 0.12017f
C20762 VPWR.n2477 VGND 0.10877f
C20763 VPWR.n2478 VGND 0.00732f
C20764 VPWR.n2479 VGND 0.01806f
C20765 VPWR.n2480 VGND 0.13984f
C20766 VPWR.n2481 VGND 0.08393f
C20767 VPWR.n2482 VGND 1.01451f
C20768 VPWR.n2483 VGND 0.19469f
C20769 VPWR.n2484 VGND 0.08393f
C20770 VPWR.n2485 VGND 0.08393f
C20771 VPWR.n2486 VGND 0.08393f
C20772 VPWR.n2487 VGND 0.08393f
C20773 VPWR.n2488 VGND 0.08393f
C20774 VPWR.n2489 VGND 0.08393f
C20775 VPWR.n2490 VGND 0.08393f
C20776 VPWR.n2491 VGND 0.08393f
C20777 VPWR.n2492 VGND 0.08393f
C20778 VPWR.n2493 VGND 0.08393f
C20779 VPWR.n2494 VGND 0.08393f
C20780 VPWR.n2495 VGND 0.08393f
C20781 VPWR.n2496 VGND 0.08393f
C20782 VPWR.n2497 VGND 0.08393f
C20783 VPWR.n2498 VGND 0.08393f
C20784 VPWR.n2499 VGND 1.01451f
C20785 VPWR.n2500 VGND 0.57419f
C20786 VPWR.n2501 VGND 0.08393f
C20787 VPWR.n2502 VGND 0.08698f
C20788 VPWR.n2503 VGND 0.00809f
C20789 VPWR.n2504 VGND 0.01723f
C20790 VPWR.n2505 VGND 0.00728f
C20791 VPWR.n2506 VGND 0.10877f
C20792 VPWR.t1274 VGND 0.12017f
C20793 VPWR.t1241 VGND 0.07889f
C20794 VPWR.t1365 VGND 0.09265f
C20795 VPWR.t1371 VGND 0.07889f
C20796 VPWR.t1386 VGND 0.12017f
C20797 VPWR.n2507 VGND 0.10877f
C20798 VPWR.n2508 VGND 0.00728f
C20799 VPWR.n2509 VGND 0.01723f
C20800 VPWR.n2510 VGND 0.00809f
C20801 VPWR.n2511 VGND 0.08698f
C20802 VPWR.n2512 VGND 0.08393f
C20803 VPWR.n2513 VGND 0.08393f
C20804 VPWR.n2514 VGND 0.08698f
C20805 VPWR.n2515 VGND 0.00809f
C20806 VPWR.n2516 VGND 0.01723f
C20807 VPWR.n2517 VGND 0.00728f
C20808 VPWR.n2518 VGND 0.10877f
C20809 VPWR.t1151 VGND 0.12017f
C20810 VPWR.t1411 VGND 0.07889f
C20811 VPWR.t1145 VGND 0.09265f
C20812 VPWR.t1135 VGND 0.07889f
C20813 VPWR.t1259 VGND 0.12017f
C20814 VPWR.n2519 VGND 0.10877f
C20815 VPWR.n2520 VGND 0.00728f
C20816 VPWR.n2521 VGND 0.01723f
C20817 VPWR.n2522 VGND 0.00809f
C20818 VPWR.n2523 VGND 0.08698f
C20819 VPWR.n2524 VGND 0.08393f
C20820 VPWR.n2525 VGND 0.08393f
C20821 VPWR.n2526 VGND 0.08698f
C20822 VPWR.n2527 VGND 0.00809f
C20823 VPWR.n2528 VGND 0.01723f
C20824 VPWR.n2529 VGND 0.00728f
C20825 VPWR.n2530 VGND 0.10877f
C20826 VPWR.t1271 VGND 0.12017f
C20827 VPWR.t1279 VGND 0.07889f
C20828 VPWR.t1408 VGND 0.09265f
C20829 VPWR.t1303 VGND 0.07889f
C20830 VPWR.t1427 VGND 0.12017f
C20831 VPWR.n2531 VGND 0.10877f
C20832 VPWR.n2532 VGND 0.00728f
C20833 VPWR.n2533 VGND 0.01723f
C20834 VPWR.n2534 VGND 0.00809f
C20835 VPWR.n2535 VGND 0.08698f
C20836 VPWR.n2536 VGND 0.08393f
C20837 VPWR.n2537 VGND 0.08393f
C20838 VPWR.n2538 VGND 0.08698f
C20839 VPWR.n2539 VGND 0.00809f
C20840 VPWR.n2540 VGND 0.01723f
C20841 VPWR.n2541 VGND 0.00728f
C20842 VPWR.n2542 VGND 0.10877f
C20843 VPWR.t1148 VGND 0.12017f
C20844 VPWR.t1140 VGND 0.07889f
C20845 VPWR.t1167 VGND 0.09265f
C20846 VPWR.t1175 VGND 0.07889f
C20847 VPWR.t1308 VGND 0.12017f
C20848 VPWR.n2543 VGND 0.10877f
C20849 VPWR.n2544 VGND 0.00728f
C20850 VPWR.n2545 VGND 0.01723f
C20851 VPWR.n2546 VGND 0.00809f
C20852 VPWR.n2547 VGND 0.08698f
C20853 VPWR.n2548 VGND 0.08393f
C20854 VPWR.n2549 VGND 0.08393f
C20855 VPWR.n2550 VGND 0.08698f
C20856 VPWR.n2551 VGND 0.00809f
C20857 VPWR.n2552 VGND 0.01723f
C20858 VPWR.n2553 VGND 0.00728f
C20859 VPWR.n2554 VGND 0.10877f
C20860 VPWR.t1324 VGND 0.12017f
C20861 VPWR.t1277 VGND 0.07889f
C20862 VPWR.t1405 VGND 0.09265f
C20863 VPWR.t1438 VGND 0.07889f
C20864 VPWR.t1454 VGND 0.12017f
C20865 VPWR.n2555 VGND 0.10877f
C20866 VPWR.n2556 VGND 0.00728f
C20867 VPWR.n2557 VGND 0.01723f
C20868 VPWR.n2558 VGND 0.00809f
C20869 VPWR.n2559 VGND 0.08698f
C20870 VPWR.n2560 VGND 0.08393f
C20871 VPWR.n2561 VGND 0.08393f
C20872 VPWR.n2562 VGND 0.08698f
C20873 VPWR.n2563 VGND 0.00809f
C20874 VPWR.n2564 VGND 0.01723f
C20875 VPWR.n2565 VGND 0.00728f
C20876 VPWR.n2566 VGND 0.10877f
C20877 VPWR.t1198 VGND 0.12017f
C20878 VPWR.t1457 VGND 0.07889f
C20879 VPWR.t1190 VGND 0.09265f
C20880 VPWR.t1311 VGND 0.07889f
C20881 VPWR.t1228 VGND 0.12017f
C20882 VPWR.n2567 VGND 0.10877f
C20883 VPWR.n2568 VGND 0.00728f
C20884 VPWR.n2569 VGND 0.01723f
C20885 VPWR.n2570 VGND 0.00809f
C20886 VPWR.n2571 VGND 0.08698f
C20887 VPWR.n2572 VGND 0.08393f
C20888 VPWR.n2573 VGND 0.08393f
C20889 VPWR.n2574 VGND 0.08698f
C20890 VPWR.n2575 VGND 0.00809f
C20891 VPWR.n2576 VGND 0.01723f
C20892 VPWR.n2577 VGND 0.00728f
C20893 VPWR.n2578 VGND 0.10877f
C20894 VPWR.t1078 VGND 0.12017f
C20895 VPWR.t1330 VGND 0.07889f
C20896 VPWR.t1451 VGND 0.09265f
C20897 VPWR.t1355 VGND 0.07889f
C20898 VPWR.t1097 VGND 0.12017f
C20899 VPWR.n2579 VGND 0.10877f
C20900 VPWR.n2580 VGND 0.00728f
C20901 VPWR.n2581 VGND 0.01723f
C20902 VPWR.n2582 VGND 0.00809f
C20903 VPWR.n2583 VGND 0.08698f
C20904 VPWR.n2584 VGND 0.08393f
C20905 VPWR.n2585 VGND 0.08393f
C20906 VPWR.n2586 VGND 0.08698f
C20907 VPWR.n2587 VGND 0.00809f
C20908 VPWR.n2588 VGND 0.01723f
C20909 VPWR.n2589 VGND 0.00728f
C20910 VPWR.n2590 VGND 0.10877f
C20911 VPWR.t1222 VGND 0.12017f
C20912 VPWR.t1206 VGND 0.07889f
C20913 VPWR.t1327 VGND 0.13401f
C20914 VPWR.n2591 VGND 0.07653f
C20915 VPWR.n2592 VGND 0.01707f
C20916 VPWR.n2593 VGND 0.00809f
C20917 VPWR.n2594 VGND 0.10908f
C20918 VPWR.n2595 VGND 0.19469f
C20919 VPWR.n2596 VGND 2.67612f
C20920 VPWR.n2597 VGND 1.08983f
C20921 VPWR.n2598 VGND 0.45664f
C20922 VPWR.t1899 VGND 0.05483f
C20923 VPWR.t1611 VGND 0.05483f
C20924 VPWR.n2599 VGND 0.09948f
C20925 VPWR.n2600 VGND 0.0471f
C20926 VPWR.t1898 VGND 0.0144f
C20927 VPWR.t1902 VGND 0.0144f
C20928 VPWR.n2601 VGND 0.03091f
C20929 VPWR.t1621 VGND 0.0144f
C20930 VPWR.t1609 VGND 0.0144f
C20931 VPWR.n2602 VGND 0.03091f
C20932 VPWR.n2603 VGND 0.0107f
C20933 VPWR.n2604 VGND 0.0471f
C20934 VPWR.t525 VGND 0.0144f
C20935 VPWR.t506 VGND 0.0144f
C20936 VPWR.n2605 VGND 0.03091f
C20937 VPWR.t489 VGND 0.0144f
C20938 VPWR.t495 VGND 0.0144f
C20939 VPWR.n2606 VGND 0.03091f
C20940 VPWR.t502 VGND 0.05743f
C20941 VPWR.t481 VGND 0.05743f
C20942 VPWR.n2607 VGND 0.13242f
C20943 VPWR.n2608 VGND 0.0425f
C20944 VPWR.n2609 VGND 0.01369f
C20945 VPWR.n2610 VGND 0.06214f
C20946 VPWR.n2611 VGND 0.00925f
C20947 VPWR.t483 VGND 0.0144f
C20948 VPWR.t1901 VGND 0.0144f
C20949 VPWR.n2612 VGND 0.03091f
C20950 VPWR.t501 VGND 0.0144f
C20951 VPWR.t1617 VGND 0.0144f
C20952 VPWR.n2613 VGND 0.03091f
C20953 VPWR.n2614 VGND 0.06214f
C20954 VPWR.n2615 VGND 0.01433f
C20955 VPWR.n2616 VGND 0.0471f
C20956 VPWR.n2617 VGND 0.0471f
C20957 VPWR.n2618 VGND 0.0471f
C20958 VPWR.n2619 VGND 0.01287f
C20959 VPWR.n2620 VGND 0.06214f
C20960 VPWR.n2621 VGND 0.01215f
C20961 VPWR.n2622 VGND 0.00988f
C20962 VPWR.n2623 VGND 0.0471f
C20963 VPWR.n2624 VGND 0.03533f
C20964 VPWR.n2625 VGND 0.00798f
C20965 VPWR.t480 VGND 0.17206f
C20966 VPWR.t488 VGND 0.25357f
C20967 VPWR.t494 VGND 0.25357f
C20968 VPWR.t482 VGND 0.25357f
C20969 VPWR.t1616 VGND 0.25357f
C20970 VPWR.t1620 VGND 0.25357f
C20971 VPWR.t1608 VGND 0.25357f
C20972 VPWR.t1610 VGND 0.56452f
C20973 VPWR.n2626 VGND 0.61616f
C20974 VPWR.n2627 VGND 0.01792f
C20975 VPWR.n2628 VGND 1.08075f
C20976 VPWR.n2629 VGND 0.0471f
C20977 VPWR.t478 VGND 0.17206f
C20978 VPWR.t491 VGND 0.25357f
C20979 VPWR.t465 VGND 0.25357f
C20980 VPWR.t517 VGND 0.25357f
C20981 VPWR.t1527 VGND 0.25357f
C20982 VPWR.t56 VGND 0.25357f
C20983 VPWR.t1525 VGND 0.25357f
C20984 VPWR.t54 VGND 0.41657f
C20985 VPWR.t237 VGND 0.44223f
C20986 VPWR.n2630 VGND 0.62407f
C20987 VPWR.n2631 VGND 0.17752f
C20988 VPWR.n2632 VGND 0.0471f
C20989 VPWR.t57 VGND 0.0144f
C20990 VPWR.t1526 VGND 0.0144f
C20991 VPWR.n2633 VGND 0.03091f
C20992 VPWR.t1780 VGND 0.0144f
C20993 VPWR.t1786 VGND 0.0144f
C20994 VPWR.n2634 VGND 0.03091f
C20995 VPWR.n2635 VGND 0.06214f
C20996 VPWR.n2636 VGND 0.0471f
C20997 VPWR.t528 VGND 0.0144f
C20998 VPWR.t1528 VGND 0.0144f
C20999 VPWR.n2637 VGND 0.03091f
C21000 VPWR.t518 VGND 0.0144f
C21001 VPWR.t1784 VGND 0.0144f
C21002 VPWR.n2638 VGND 0.03091f
C21003 VPWR.n2639 VGND 0.00925f
C21004 VPWR.t479 VGND 0.05743f
C21005 VPWR.t527 VGND 0.05743f
C21006 VPWR.n2640 VGND 0.13242f
C21007 VPWR.t510 VGND 0.0144f
C21008 VPWR.t485 VGND 0.0144f
C21009 VPWR.n2641 VGND 0.03091f
C21010 VPWR.t492 VGND 0.0144f
C21011 VPWR.t466 VGND 0.0144f
C21012 VPWR.n2642 VGND 0.03091f
C21013 VPWR.n2643 VGND 0.06214f
C21014 VPWR.n2644 VGND 0.01369f
C21015 VPWR.n2645 VGND 0.0425f
C21016 VPWR.n2646 VGND 0.0471f
C21017 VPWR.n2647 VGND 0.0471f
C21018 VPWR.n2648 VGND 0.01433f
C21019 VPWR.n2649 VGND 0.06214f
C21020 VPWR.n2650 VGND 0.0107f
C21021 VPWR.n2651 VGND 0.01287f
C21022 VPWR.n2652 VGND 0.0471f
C21023 VPWR.n2653 VGND 0.0471f
C21024 VPWR.n2654 VGND 0.01215f
C21025 VPWR.n2655 VGND 0.00988f
C21026 VPWR.t55 VGND 0.05483f
C21027 VPWR.t1782 VGND 0.05483f
C21028 VPWR.n2656 VGND 0.09948f
C21029 VPWR.n2657 VGND 0.00798f
C21030 VPWR.n2658 VGND 0.03533f
C21031 VPWR.n2659 VGND 0.01792f
C21032 VPWR.n2660 VGND 0.03533f
C21033 VPWR.n2661 VGND 0.01405f
C21034 VPWR.n2662 VGND 0.01088f
C21035 VPWR.t238 VGND 0.05737f
C21036 VPWR.t884 VGND 0.05737f
C21037 VPWR.n2663 VGND 0.11596f
C21038 VPWR.n2664 VGND 0.03277f
C21039 VPWR.n2665 VGND 1.64485f
C21040 VPWR.n2666 VGND 0.0471f
C21041 VPWR.t886 VGND 0.05631f
C21042 VPWR.t512 VGND 0.17206f
C21043 VPWR.t469 VGND 0.25357f
C21044 VPWR.t519 VGND 0.25357f
C21045 VPWR.t496 VGND 0.25357f
C21046 VPWR.t413 VGND 0.25357f
C21047 VPWR.t651 VGND 0.25357f
C21048 VPWR.t1018 VGND 0.25357f
C21049 VPWR.t143 VGND 0.41657f
C21050 VPWR.t398 VGND 0.15999f
C21051 VPWR.t885 VGND 0.12678f
C21052 VPWR.t615 VGND 0.28224f
C21053 VPWR.n2667 VGND 0.55313f
C21054 VPWR.n2668 VGND 0.17489f
C21055 VPWR.n2669 VGND 0.0471f
C21056 VPWR.t1014 VGND 0.0144f
C21057 VPWR.t1019 VGND 0.0144f
C21058 VPWR.n2670 VGND 0.03091f
C21059 VPWR.t652 VGND 0.0144f
C21060 VPWR.t1662 VGND 0.0144f
C21061 VPWR.n2671 VGND 0.03091f
C21062 VPWR.n2672 VGND 0.06214f
C21063 VPWR.n2673 VGND 0.0471f
C21064 VPWR.t514 VGND 0.0144f
C21065 VPWR.t1017 VGND 0.0144f
C21066 VPWR.n2674 VGND 0.03091f
C21067 VPWR.t497 VGND 0.0144f
C21068 VPWR.t414 VGND 0.0144f
C21069 VPWR.n2675 VGND 0.03091f
C21070 VPWR.n2676 VGND 0.00925f
C21071 VPWR.t526 VGND 0.05743f
C21072 VPWR.t513 VGND 0.05743f
C21073 VPWR.n2677 VGND 0.13242f
C21074 VPWR.t486 VGND 0.0144f
C21075 VPWR.t532 VGND 0.0144f
C21076 VPWR.n2678 VGND 0.03091f
C21077 VPWR.t470 VGND 0.0144f
C21078 VPWR.t520 VGND 0.0144f
C21079 VPWR.n2679 VGND 0.03091f
C21080 VPWR.n2680 VGND 0.06214f
C21081 VPWR.n2681 VGND 0.01369f
C21082 VPWR.n2682 VGND 0.0425f
C21083 VPWR.n2683 VGND 0.0471f
C21084 VPWR.n2684 VGND 0.0471f
C21085 VPWR.n2685 VGND 0.01433f
C21086 VPWR.n2686 VGND 0.06214f
C21087 VPWR.n2687 VGND 0.0107f
C21088 VPWR.n2688 VGND 0.01287f
C21089 VPWR.n2689 VGND 0.0471f
C21090 VPWR.n2690 VGND 0.0471f
C21091 VPWR.n2691 VGND 0.01215f
C21092 VPWR.n2692 VGND 0.00988f
C21093 VPWR.t1015 VGND 0.05483f
C21094 VPWR.t144 VGND 0.05483f
C21095 VPWR.n2693 VGND 0.09948f
C21096 VPWR.n2694 VGND 0.00798f
C21097 VPWR.n2695 VGND 0.03533f
C21098 VPWR.n2696 VGND 0.01792f
C21099 VPWR.n2697 VGND 0.03533f
C21100 VPWR.t616 VGND 0.05743f
C21101 VPWR.n2698 VGND 0.08004f
C21102 VPWR.n2699 VGND 0.0107f
C21103 VPWR.n2700 VGND 0.05857f
C21104 VPWR.t399 VGND 0.05646f
C21105 VPWR.n2701 VGND 0.07318f
C21106 VPWR.n2702 VGND 0.0279f
C21107 VPWR.n2703 VGND 1.64485f
C21108 VPWR.n2704 VGND 0.0471f
C21109 VPWR.t515 VGND 0.09758f
C21110 VPWR.t473 VGND 0.14381f
C21111 VPWR.t521 VGND 0.13981f
C21112 VPWR.t499 VGND 0.22359f
C21113 VPWR.t649 VGND 0.19017f
C21114 VPWR.t503 VGND 0.12678f
C21115 VPWR.t545 VGND 0.12678f
C21116 VPWR.t475 VGND 0.12678f
C21117 VPWR.t1066 VGND 0.12678f
C21118 VPWR.t507 VGND 0.12678f
C21119 VPWR.t292 VGND 0.12678f
C21120 VPWR.t530 VGND 0.17659f
C21121 VPWR.t1778 VGND 0.09962f
C21122 VPWR.t541 VGND 0.10867f
C21123 VPWR.t613 VGND 0.12678f
C21124 VPWR.t543 VGND 0.23545f
C21125 VPWR.n2705 VGND 0.37955f
C21126 VPWR.n2706 VGND 0.17507f
C21127 VPWR.t544 VGND 0.057f
C21128 VPWR.n2707 VGND 0.0471f
C21129 VPWR.t531 VGND 0.05635f
C21130 VPWR.t293 VGND 0.05425f
C21131 VPWR.t476 VGND 0.0144f
C21132 VPWR.t508 VGND 0.0144f
C21133 VPWR.n2708 VGND 0.03091f
C21134 VPWR.t546 VGND 0.0144f
C21135 VPWR.t1067 VGND 0.0144f
C21136 VPWR.n2709 VGND 0.03091f
C21137 VPWR.n2710 VGND 0.03524f
C21138 VPWR.n2711 VGND 0.0471f
C21139 VPWR.t500 VGND 0.0144f
C21140 VPWR.t650 VGND 0.0144f
C21141 VPWR.n2712 VGND 0.03091f
C21142 VPWR.n2713 VGND 0.00925f
C21143 VPWR.t516 VGND 0.05743f
C21144 VPWR.n2714 VGND 0.07237f
C21145 VPWR.t474 VGND 0.0144f
C21146 VPWR.t522 VGND 0.0144f
C21147 VPWR.n2715 VGND 0.03091f
C21148 VPWR.n2716 VGND 0.03524f
C21149 VPWR.n2717 VGND 0.01369f
C21150 VPWR.n2718 VGND 0.0425f
C21151 VPWR.n2719 VGND 0.0471f
C21152 VPWR.n2720 VGND 0.0471f
C21153 VPWR.n2721 VGND 0.01433f
C21154 VPWR.n2722 VGND 0.03443f
C21155 VPWR.t504 VGND 0.0504f
C21156 VPWR.n2723 VGND 0.04018f
C21157 VPWR.n2724 VGND 0.00988f
C21158 VPWR.n2725 VGND 0.0471f
C21159 VPWR.n2726 VGND 0.0471f
C21160 VPWR.n2727 VGND 0.03905f
C21161 VPWR.n2728 VGND 0.01215f
C21162 VPWR.n2729 VGND 0.05168f
C21163 VPWR.n2730 VGND 0.0681f
C21164 VPWR.n2731 VGND 0.00626f
C21165 VPWR.n2732 VGND 0.0279f
C21166 VPWR.n2733 VGND 0.01792f
C21167 VPWR.n2734 VGND 0.03533f
C21168 VPWR.t614 VGND 0.05749f
C21169 VPWR.n2735 VGND 0.1478f
C21170 VPWR.n2736 VGND 0.01088f
C21171 VPWR.t542 VGND 0.0574f
C21172 VPWR.n2737 VGND 0.06389f
C21173 VPWR.n2738 VGND 0.02765f
C21174 VPWR.n2739 VGND 1.64485f
C21175 VPWR.n2740 VGND 0.0425f
C21176 VPWR.t509 VGND 0.67014f
C21177 VPWR.t468 VGND 0.25357f
C21178 VPWR.t498 VGND 0.25357f
C21179 VPWR.t472 VGND 0.25357f
C21180 VPWR.t1614 VGND 0.25357f
C21181 VPWR.t1612 VGND 0.25357f
C21182 VPWR.t1618 VGND 0.25357f
C21183 VPWR.t1606 VGND 0.22942f
C21184 VPWR.t690 VGND 0.55543f
C21185 VPWR.t428 VGND 0.15395f
C21186 VPWR.n2741 VGND 0.33277f
C21187 VPWR.n2742 VGND 0.17752f
C21188 VPWR.t1903 VGND 0.0144f
C21189 VPWR.t1900 VGND 0.0144f
C21190 VPWR.n2743 VGND 0.03156f
C21191 VPWR.t1615 VGND 0.0144f
C21192 VPWR.t1613 VGND 0.0144f
C21193 VPWR.n2744 VGND 0.03156f
C21194 VPWR.n2745 VGND 0.1198f
C21195 VPWR.n2746 VGND 0.09713f
C21196 VPWR.t1904 VGND 0.0144f
C21197 VPWR.t1905 VGND 0.0144f
C21198 VPWR.n2747 VGND 0.03162f
C21199 VPWR.t1619 VGND 0.0144f
C21200 VPWR.t1607 VGND 0.0144f
C21201 VPWR.n2748 VGND 0.03162f
C21202 VPWR.n2749 VGND 0.13131f
C21203 VPWR.n2750 VGND 0.01124f
C21204 VPWR.n2751 VGND 0.37932f
C21205 VPWR.n2752 VGND 0.01792f
C21206 VPWR.n2753 VGND 0.01638f
C21207 VPWR.n2754 VGND 0.01405f
C21208 VPWR.n2755 VGND 0.01315f
C21209 VPWR.t1860 VGND 0.05749f
C21210 VPWR.t691 VGND 0.05749f
C21211 VPWR.n2756 VGND 0.16979f
C21212 VPWR.n2757 VGND 0.03533f
C21213 VPWR.n2758 VGND 1.64485f
C21214 VPWR.n2759 VGND 0.0425f
C21215 VPWR.t490 VGND 0.67014f
C21216 VPWR.t523 VGND 0.25357f
C21217 VPWR.t477 VGND 0.25357f
C21218 VPWR.t524 VGND 0.25357f
C21219 VPWR.t1523 VGND 0.25357f
C21220 VPWR.t52 VGND 0.25357f
C21221 VPWR.t48 VGND 0.25357f
C21222 VPWR.t46 VGND 0.22942f
C21223 VPWR.t1920 VGND 0.49355f
C21224 VPWR.t430 VGND 0.10867f
C21225 VPWR.t434 VGND 0.10716f
C21226 VPWR.n2760 VGND 0.33126f
C21227 VPWR.n2761 VGND 0.17752f
C21228 VPWR.t1524 VGND 0.0144f
C21229 VPWR.t53 VGND 0.0144f
C21230 VPWR.n2762 VGND 0.03156f
C21231 VPWR.t1779 VGND 0.0144f
C21232 VPWR.t1785 VGND 0.0144f
C21233 VPWR.n2763 VGND 0.03156f
C21234 VPWR.n2764 VGND 0.1198f
C21235 VPWR.n2765 VGND 0.09713f
C21236 VPWR.t49 VGND 0.0144f
C21237 VPWR.t47 VGND 0.0144f
C21238 VPWR.n2766 VGND 0.03162f
C21239 VPWR.t1781 VGND 0.0144f
C21240 VPWR.t1783 VGND 0.0144f
C21241 VPWR.n2767 VGND 0.03162f
C21242 VPWR.n2768 VGND 0.13131f
C21243 VPWR.n2769 VGND 0.01124f
C21244 VPWR.n2770 VGND 0.37932f
C21245 VPWR.n2771 VGND 0.01792f
C21246 VPWR.n2772 VGND 0.01613f
C21247 VPWR.n2773 VGND 0.00771f
C21248 VPWR.t431 VGND 0.05737f
C21249 VPWR.n2774 VGND 0.06132f
C21250 VPWR.n2775 VGND 0.00734f
C21251 VPWR.t1921 VGND 0.05749f
C21252 VPWR.n2776 VGND 0.09156f
C21253 VPWR.n2777 VGND 0.03533f
C21254 VPWR.n2778 VGND 1.64485f
C21255 VPWR.n2779 VGND 0.04301f
C21256 VPWR.t471 VGND 0.67014f
C21257 VPWR.t484 VGND 0.25357f
C21258 VPWR.t511 VGND 0.25357f
C21259 VPWR.t487 VGND 0.25357f
C21260 VPWR.t342 VGND 0.25357f
C21261 VPWR.t133 VGND 0.25357f
C21262 VPWR.t1011 VGND 0.25357f
C21263 VPWR.t548 VGND 0.22942f
C21264 VPWR.t688 VGND 0.52524f
C21265 VPWR.t426 VGND 0.18112f
C21266 VPWR.n2780 VGND 0.32975f
C21267 VPWR.n2781 VGND 0.17489f
C21268 VPWR.t429 VGND 0.05745f
C21269 VPWR.t1020 VGND 0.0144f
C21270 VPWR.t1016 VGND 0.0144f
C21271 VPWR.n2782 VGND 0.03156f
C21272 VPWR.t343 VGND 0.0144f
C21273 VPWR.t134 VGND 0.0144f
C21274 VPWR.n2783 VGND 0.03156f
C21275 VPWR.n2784 VGND 0.1198f
C21276 VPWR.n2785 VGND 0.09713f
C21277 VPWR.t1012 VGND 0.0144f
C21278 VPWR.t1013 VGND 0.0144f
C21279 VPWR.n2786 VGND 0.03162f
C21280 VPWR.t1559 VGND 0.0144f
C21281 VPWR.t549 VGND 0.0144f
C21282 VPWR.n2787 VGND 0.03162f
C21283 VPWR.n2788 VGND 0.13131f
C21284 VPWR.n2789 VGND 0.01124f
C21285 VPWR.n2790 VGND 0.37932f
C21286 VPWR.n2791 VGND 0.01792f
C21287 VPWR.n2792 VGND 0.01587f
C21288 VPWR.t427 VGND 0.05745f
C21289 VPWR.n2793 VGND 0.15135f
C21290 VPWR.n2794 VGND 0.01215f
C21291 VPWR.t1861 VGND 0.05743f
C21292 VPWR.t689 VGND 0.05743f
C21293 VPWR.n2795 VGND 0.13514f
C21294 VPWR.n2796 VGND 0.03533f
C21295 VPWR.n2797 VGND 1.64485f
C21296 VPWR.n2798 VGND 0.04301f
C21297 VPWR.t1919 VGND 0.05743f
C21298 VPWR.n2799 VGND 0.01587f
C21299 VPWR.t433 VGND 0.05745f
C21300 VPWR.n2800 VGND 0.01792f
C21301 VPWR.t505 VGND 0.38006f
C21302 VPWR.t529 VGND 0.14381f
C21303 VPWR.t493 VGND 0.14381f
C21304 VPWR.t467 VGND 0.14381f
C21305 VPWR.t290 VGND 0.14381f
C21306 VPWR.t50 VGND 0.14381f
C21307 VPWR.t1070 VGND 0.14381f
C21308 VPWR.t1912 VGND 0.13011f
C21309 VPWR.t1918 VGND 0.29789f
C21310 VPWR.t432 VGND 0.10272f
C21311 VPWR.n2801 VGND 0.18352f
C21312 VPWR.t1071 VGND 0.0144f
C21313 VPWR.t1913 VGND 0.0144f
C21314 VPWR.n2802 VGND 0.03162f
C21315 VPWR.n2803 VGND 0.07781f
C21316 VPWR.t291 VGND 0.0144f
C21317 VPWR.t51 VGND 0.0144f
C21318 VPWR.n2804 VGND 0.03291f
C21319 VPWR.n2805 VGND 0.17568f
C21320 VPWR.n2806 VGND 0.37932f
C21321 VPWR.n2807 VGND 0.01124f
C21322 VPWR.n2808 VGND 0.0971f
C21323 VPWR.n2809 VGND 0.08524f
C21324 VPWR.n2810 VGND 0.01215f
C21325 VPWR.n2811 VGND 0.07387f
C21326 VPWR.n2812 VGND 0.03533f
C21327 VPWR.n2813 VGND 2.39365f
C21328 VPWR.n2814 VGND 1.93855f
C21329 VPWR.t1561 VGND 0.0292f
C21330 VPWR.n2815 VGND 0.13089f
C21331 VPWR.n2816 VGND 0.28811f
C21332 VPWR.n2817 VGND 0.07598f
C21333 VPWR.n2818 VGND 0.03609f
C21334 VPWR.n2819 VGND 0.04406f
C21335 VPWR.n2820 VGND 0.08931f
C21336 VPWR.n2821 VGND 0.11642f
C21337 VPWR.n2822 VGND 0.08931f
C21338 VPWR.t556 VGND 2.8091f
C21339 VPWR.t1560 VGND 0.88722f
C21340 VPWR.n2823 VGND 0.11733f
C21341 VPWR.n2824 VGND 0.46422f
C21342 VPWR.t734 VGND 0.02919f
C21343 VPWR.n2825 VGND 0.17872f
C21344 VPWR.n2826 VGND 0.01804f
C21345 VPWR.n2827 VGND 0.09846f
C21346 VPWR.n2828 VGND 0.0884f
C21347 VPWR.n2829 VGND 0.11733f
C21348 VPWR.n2830 VGND 0.07389f
C21349 VPWR.t557 VGND 0.02919f
C21350 VPWR.n2831 VGND 0.17872f
C21351 VPWR.n2832 VGND 0.01804f
C21352 VPWR.n2833 VGND 0.11733f
C21353 VPWR.n2834 VGND 0.07678f
C21354 VPWR.n2835 VGND 0.08757f
C21355 VPWR.n2836 VGND 1.67873f
C21356 VPWR.n2837 VGND 0.08757f
C21357 VPWR.n2838 VGND 0.07678f
C21358 VPWR.n2839 VGND 0.11733f
C21359 VPWR.n2840 VGND 0.09837f
C21360 VPWR.n2841 VGND 0.08137f
C21361 VPWR.n2842 VGND 1.0091f
C21362 VPWR.n2843 VGND 0.06349f
C21363 VPWR.n2844 VGND 0.08881f
C21364 VPWR.n2845 VGND 0.06174f
C21365 VPWR.n2846 VGND 0.01804f
C21366 VPWR.n2847 VGND 0.06349f
C21367 VPWR.n2848 VGND 0.04875f
C21368 VPWR.n2849 VGND 0.17444f
C21369 VPWR.n2850 VGND 0.06872f
C21370 VPWR.n2851 VGND 0.04406f
C21371 VPWR.t447 VGND 0.34736f
C21372 VPWR.n2852 VGND 0.08137f
C21373 VPWR.n2853 VGND 0.09837f
C21374 VPWR.n2854 VGND 0.03609f
C21375 VPWR.n2855 VGND 2.0331f
C21376 VPWR.n2856 VGND 0.03609f
C21377 VPWR.n2857 VGND 0.03609f
C21378 VPWR.n2858 VGND 0.08967f
C21379 VPWR.n2859 VGND 0.04923f
C21380 VPWR.n2860 VGND 0.38128f
C21381 VPWR.n2861 VGND 0.31371f
C21382 VPWR.t448 VGND 0.02918f
C21383 VPWR.n2862 VGND 0.22078f
C21384 VPWR.n2863 VGND 3.49571f
C21385 XThR.Tn[2].t5 VGND 0.02313f
C21386 XThR.Tn[2].t2 VGND 0.02313f
C21387 XThR.Tn[2].n0 VGND 0.04668f
C21388 XThR.Tn[2].t4 VGND 0.02313f
C21389 XThR.Tn[2].t3 VGND 0.02313f
C21390 XThR.Tn[2].n1 VGND 0.05462f
C21391 XThR.Tn[2].n2 VGND 0.16384f
C21392 XThR.Tn[2].t7 VGND 0.01503f
C21393 XThR.Tn[2].t8 VGND 0.01503f
C21394 XThR.Tn[2].n3 VGND 0.03423f
C21395 XThR.Tn[2].t6 VGND 0.01503f
C21396 XThR.Tn[2].t1 VGND 0.01503f
C21397 XThR.Tn[2].n4 VGND 0.03423f
C21398 XThR.Tn[2].t9 VGND 0.01503f
C21399 XThR.Tn[2].t10 VGND 0.01503f
C21400 XThR.Tn[2].n5 VGND 0.05704f
C21401 XThR.Tn[2].t11 VGND 0.01503f
C21402 XThR.Tn[2].t0 VGND 0.01503f
C21403 XThR.Tn[2].n6 VGND 0.03423f
C21404 XThR.Tn[2].n7 VGND 0.16303f
C21405 XThR.Tn[2].n8 VGND 0.10078f
C21406 XThR.Tn[2].n9 VGND 0.11374f
C21407 XThR.Tn[2].t21 VGND 0.01808f
C21408 XThR.Tn[2].t14 VGND 0.01979f
C21409 XThR.Tn[2].n10 VGND 0.04833f
C21410 XThR.Tn[2].n11 VGND 0.09285f
C21411 XThR.Tn[2].t40 VGND 0.01808f
C21412 XThR.Tn[2].t31 VGND 0.01979f
C21413 XThR.Tn[2].n12 VGND 0.04833f
C21414 XThR.Tn[2].t55 VGND 0.01802f
C21415 XThR.Tn[2].t66 VGND 0.01973f
C21416 XThR.Tn[2].n13 VGND 0.05029f
C21417 XThR.Tn[2].n14 VGND 0.03533f
C21418 XThR.Tn[2].n15 VGND 0.00646f
C21419 XThR.Tn[2].n16 VGND 0.11337f
C21420 XThR.Tn[2].t15 VGND 0.01808f
C21421 XThR.Tn[2].t67 VGND 0.01979f
C21422 XThR.Tn[2].n17 VGND 0.04833f
C21423 XThR.Tn[2].t30 VGND 0.01802f
C21424 XThR.Tn[2].t43 VGND 0.01973f
C21425 XThR.Tn[2].n18 VGND 0.05029f
C21426 XThR.Tn[2].n19 VGND 0.03533f
C21427 XThR.Tn[2].n20 VGND 0.00646f
C21428 XThR.Tn[2].n21 VGND 0.11337f
C21429 XThR.Tn[2].t32 VGND 0.01808f
C21430 XThR.Tn[2].t23 VGND 0.01979f
C21431 XThR.Tn[2].n22 VGND 0.04833f
C21432 XThR.Tn[2].t47 VGND 0.01802f
C21433 XThR.Tn[2].t60 VGND 0.01973f
C21434 XThR.Tn[2].n23 VGND 0.05029f
C21435 XThR.Tn[2].n24 VGND 0.03533f
C21436 XThR.Tn[2].n25 VGND 0.00646f
C21437 XThR.Tn[2].n26 VGND 0.11337f
C21438 XThR.Tn[2].t58 VGND 0.01808f
C21439 XThR.Tn[2].t50 VGND 0.01979f
C21440 XThR.Tn[2].n27 VGND 0.04833f
C21441 XThR.Tn[2].t16 VGND 0.01802f
C21442 XThR.Tn[2].t28 VGND 0.01973f
C21443 XThR.Tn[2].n28 VGND 0.05029f
C21444 XThR.Tn[2].n29 VGND 0.03533f
C21445 XThR.Tn[2].n30 VGND 0.00646f
C21446 XThR.Tn[2].n31 VGND 0.11337f
C21447 XThR.Tn[2].t34 VGND 0.01808f
C21448 XThR.Tn[2].t25 VGND 0.01979f
C21449 XThR.Tn[2].n32 VGND 0.04833f
C21450 XThR.Tn[2].t48 VGND 0.01802f
C21451 XThR.Tn[2].t62 VGND 0.01973f
C21452 XThR.Tn[2].n33 VGND 0.05029f
C21453 XThR.Tn[2].n34 VGND 0.03533f
C21454 XThR.Tn[2].n35 VGND 0.00646f
C21455 XThR.Tn[2].n36 VGND 0.11337f
C21456 XThR.Tn[2].t70 VGND 0.01808f
C21457 XThR.Tn[2].t41 VGND 0.01979f
C21458 XThR.Tn[2].n37 VGND 0.04833f
C21459 XThR.Tn[2].t22 VGND 0.01802f
C21460 XThR.Tn[2].t20 VGND 0.01973f
C21461 XThR.Tn[2].n38 VGND 0.05029f
C21462 XThR.Tn[2].n39 VGND 0.03533f
C21463 XThR.Tn[2].n40 VGND 0.00646f
C21464 XThR.Tn[2].n41 VGND 0.11337f
C21465 XThR.Tn[2].t39 VGND 0.01808f
C21466 XThR.Tn[2].t35 VGND 0.01979f
C21467 XThR.Tn[2].n42 VGND 0.04833f
C21468 XThR.Tn[2].t54 VGND 0.01802f
C21469 XThR.Tn[2].t12 VGND 0.01973f
C21470 XThR.Tn[2].n43 VGND 0.05029f
C21471 XThR.Tn[2].n44 VGND 0.03533f
C21472 XThR.Tn[2].n45 VGND 0.00646f
C21473 XThR.Tn[2].n46 VGND 0.11337f
C21474 XThR.Tn[2].t44 VGND 0.01808f
C21475 XThR.Tn[2].t49 VGND 0.01979f
C21476 XThR.Tn[2].n47 VGND 0.04833f
C21477 XThR.Tn[2].t57 VGND 0.01802f
C21478 XThR.Tn[2].t27 VGND 0.01973f
C21479 XThR.Tn[2].n48 VGND 0.05029f
C21480 XThR.Tn[2].n49 VGND 0.03533f
C21481 XThR.Tn[2].n50 VGND 0.00646f
C21482 XThR.Tn[2].n51 VGND 0.11337f
C21483 XThR.Tn[2].t61 VGND 0.01808f
C21484 XThR.Tn[2].t69 VGND 0.01979f
C21485 XThR.Tn[2].n52 VGND 0.04833f
C21486 XThR.Tn[2].t18 VGND 0.01802f
C21487 XThR.Tn[2].t45 VGND 0.01973f
C21488 XThR.Tn[2].n53 VGND 0.05029f
C21489 XThR.Tn[2].n54 VGND 0.03533f
C21490 XThR.Tn[2].n55 VGND 0.00646f
C21491 XThR.Tn[2].n56 VGND 0.11337f
C21492 XThR.Tn[2].t52 VGND 0.01808f
C21493 XThR.Tn[2].t26 VGND 0.01979f
C21494 XThR.Tn[2].n57 VGND 0.04833f
C21495 XThR.Tn[2].t68 VGND 0.01802f
C21496 XThR.Tn[2].t63 VGND 0.01973f
C21497 XThR.Tn[2].n58 VGND 0.05029f
C21498 XThR.Tn[2].n59 VGND 0.03533f
C21499 XThR.Tn[2].n60 VGND 0.00646f
C21500 XThR.Tn[2].n61 VGND 0.11337f
C21501 XThR.Tn[2].t73 VGND 0.01808f
C21502 XThR.Tn[2].t64 VGND 0.01979f
C21503 XThR.Tn[2].n62 VGND 0.04833f
C21504 XThR.Tn[2].t24 VGND 0.01802f
C21505 XThR.Tn[2].t37 VGND 0.01973f
C21506 XThR.Tn[2].n63 VGND 0.05029f
C21507 XThR.Tn[2].n64 VGND 0.03533f
C21508 XThR.Tn[2].n65 VGND 0.00646f
C21509 XThR.Tn[2].n66 VGND 0.11337f
C21510 XThR.Tn[2].t42 VGND 0.01808f
C21511 XThR.Tn[2].t36 VGND 0.01979f
C21512 XThR.Tn[2].n67 VGND 0.04833f
C21513 XThR.Tn[2].t56 VGND 0.01802f
C21514 XThR.Tn[2].t13 VGND 0.01973f
C21515 XThR.Tn[2].n68 VGND 0.05029f
C21516 XThR.Tn[2].n69 VGND 0.03533f
C21517 XThR.Tn[2].n70 VGND 0.00646f
C21518 XThR.Tn[2].n71 VGND 0.11337f
C21519 XThR.Tn[2].t59 VGND 0.01808f
C21520 XThR.Tn[2].t51 VGND 0.01979f
C21521 XThR.Tn[2].n72 VGND 0.04833f
C21522 XThR.Tn[2].t17 VGND 0.01802f
C21523 XThR.Tn[2].t29 VGND 0.01973f
C21524 XThR.Tn[2].n73 VGND 0.05029f
C21525 XThR.Tn[2].n74 VGND 0.03533f
C21526 XThR.Tn[2].n75 VGND 0.00646f
C21527 XThR.Tn[2].n76 VGND 0.11337f
C21528 XThR.Tn[2].t19 VGND 0.01808f
C21529 XThR.Tn[2].t72 VGND 0.01979f
C21530 XThR.Tn[2].n77 VGND 0.04833f
C21531 XThR.Tn[2].t33 VGND 0.01802f
C21532 XThR.Tn[2].t46 VGND 0.01973f
C21533 XThR.Tn[2].n78 VGND 0.05029f
C21534 XThR.Tn[2].n79 VGND 0.03533f
C21535 XThR.Tn[2].n80 VGND 0.00646f
C21536 XThR.Tn[2].n81 VGND 0.11337f
C21537 XThR.Tn[2].t53 VGND 0.01808f
C21538 XThR.Tn[2].t65 VGND 0.01979f
C21539 XThR.Tn[2].n82 VGND 0.04833f
C21540 XThR.Tn[2].t71 VGND 0.01802f
C21541 XThR.Tn[2].t38 VGND 0.01973f
C21542 XThR.Tn[2].n83 VGND 0.05029f
C21543 XThR.Tn[2].n84 VGND 0.03533f
C21544 XThR.Tn[2].n85 VGND 0.00646f
C21545 XThR.Tn[2].n86 VGND 0.11337f
C21546 XThR.Tn[2].n87 VGND 0.10303f
C21547 XThR.Tn[2].n88 VGND 0.22327f
.ends

