** sch_path: /home/anton/projects/NEW-ttsky25b-analog-vga-dacs/xschem/vbias085.sch
.subckt vbias085 VPWR VGND bias[2] bias[1] bias[0] Vbias
*.PININFO VPWR:B VGND:B bias[2:0]:I Vbias:O
XM1 Vbias bias[2] VPWR VPWR sky130_fd_pr__pfet_01v8 L=0.5 W=0.85 nf=1 m=1
XM2 Vbias bias[1] VPWR VPWR sky130_fd_pr__pfet_01v8 L=1 W=0.85 nf=1 m=1
XM3 Vbias bias[0] VPWR VPWR sky130_fd_pr__pfet_01v8 L=2 W=0.85 nf=1 m=1
XM4 Vbias VGND VPWR VPWR sky130_fd_pr__pfet_01v8 L=2 W=0.85 nf=1 m=1
XMmirror Vbias Vbias VGND VGND sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2.6 nf=1 m=1
.ends
