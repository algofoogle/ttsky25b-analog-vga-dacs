* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1961 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t1541 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1540 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t234 VGND.t2415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1458 VPWR.t1460 VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t782 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t781 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t575 XThR.XTBN.Y.t4 a_n997_2667# VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t480 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t479 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t521 VPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t1988 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t3 XThC.XTBN.Y.t4 VGND.t512 VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1931 VGND.t497 VGND.t496 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t2577 VGND.t2576 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t513 XThC.XTBN.Y.t5 XThC.Tn[5].t3 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t162 VGND.t1682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t1990 VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t2438 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t2437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t219 VGND.t2333 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t53 VGND.t369 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t7 XThC.XTB5.Y VPWR.t683 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1932 VGND.t499 VGND.t498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t198 VGND.t1953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t835 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t3 VPWR.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1456 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1457 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t197 VGND.t1952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t225 VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t7 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t864 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1135 VGND.t1137 VGND.t1136 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t1310 VGND.t1309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t3 XThR.XTBN.Y.t5 a_n1049_5611# VPWR.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t1287 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t669 XThC.XTBN.Y.t8 XThC.Tn[2].t6 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t866 VGND.t865 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t222 VGND.t2338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t2263 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t2262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t1455 VPWR.t1453 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t501 VPWR.t1933 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t500 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t708 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t707 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t803 Vbias.t12 XA.XIR[14].XIC[11].icell.SM VGND.t802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t1748 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t2381 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t2380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t503 VPWR.t1934 XA.XIR[10].XIC_15.icell.PDM VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t766 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t765 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1450 VPWR.t1452 VPWR.t1451 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t7 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t805 Vbias.t13 XA.XIR[2].XIC[5].icell.SM VGND.t804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t450 VPWR.t449 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t7 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t641 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t640 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.XTB5.Y XThC.XTB7.B VGND.t965 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t7 XThC.XTBN.Y.t9 VPWR.t340 VPWR.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t2579 VGND.t2578 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t237 XThR.XTB7.Y XThR.Tn[6].t3 VGND.t236 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t1678 VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t282 XThR.XTBN.Y.t6 XThR.Tn[9].t11 VPWR.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t838 VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t710 VPWR.t709 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t712 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t711 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t1992 VGND.t1991 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t828 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t1539 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1538 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t2367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t482 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t481 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t1449 VPWR.t1447 XA.XIR[2].XIC_15.icell.PUM VPWR.t1448 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.XTB7.Y VPWR.t843 VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t1312 VGND.t1311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t7 XThR.XTBN.Y.t7 VPWR.t284 VPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t1522 VGND.t1521 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.XTBN.Y.t10 VGND.t671 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t807 Vbias.t14 XA.XIR[12].XIC[7].icell.SM VGND.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t601 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t132 VGND.t1512 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t182 VGND.t1841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t505 VPWR.t1935 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t504 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t577 XThR.XTBN.Y.t8 XThR.Tn[5].t7 VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t809 Vbias.t15 XA.XIR[15].XIC[8].icell.SM VGND.t808 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t811 Vbias.t16 XA.XIR[14].XIC[9].icell.SM VGND.t810 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t157 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t156 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t2440 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t2439 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t2340 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t2339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t1680 VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t649 XThR.XTB6.Y a_n1049_5611# VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t813 Vbias.t17 XA.XIR[9].XIC[7].icell.SM VGND.t812 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t2265 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t2264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t907 VPWR.t906 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1936 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t506 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 a_n1049_7787# XThR.XTB2.Y VPWR.t53 VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 VGND.t1685 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t1684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X96 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t2033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X97 VGND.t815 Vbias.t18 XA.XIR[2].XIC[0].icell.SM VGND.t814 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X98 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t452 VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X99 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t320 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X100 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1445 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1446 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 VGND.t817 Vbias.t19 XA.XIR[0].XIC[13].icell.SM VGND.t816 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X102 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t1524 VGND.t1523 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X103 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1682 VPWR.t1681 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X104 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t2035 VGND.t2034 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X105 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t2037 VGND.t2036 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t714 VPWR.t713 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X107 VGND.t2657 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X108 VPWR.t151 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X109 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t829 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X110 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t2268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 VPWR.t639 data[4].t0 a_n1335_4229# VPWR.t638 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X112 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1537 VPWR.t1536 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X113 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t254 VGND.t2615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X114 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X115 VGND.t579 XThR.XTBN.Y.t9 XThR.Tn[7].t3 VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X116 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t2279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X117 a_n1319_5317# XThR.XTB7.A VPWR.t456 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X118 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t2038 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X119 VPWR.t21 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X120 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X121 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t879 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X122 XThC.Tn[9].t7 XThC.XTB2.Y VPWR.t387 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 XA.XIR[15].XIC[4].icell.Ien VPWR.t1442 VPWR.t1444 VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X124 VGND.t819 Vbias.t20 XA.XIR[12].XIC[2].icell.SM VGND.t818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X125 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t100 VGND.t978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X126 VGND.t821 Vbias.t21 XA.XIR[11].XIC_15.icell.SM VGND.t820 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X127 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1439 VPWR.t1441 VPWR.t1440 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X128 XThC.Tn[5].t2 XThC.XTBN.Y.t11 VGND.t672 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t2295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X130 VGND.t823 Vbias.t22 XA.XIR[15].XIC[3].icell.SM VGND.t822 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X131 VGND.t825 Vbias.t23 XA.XIR[14].XIC[4].icell.SM VGND.t824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t603 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X133 VPWR.t1574 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t1573 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X134 VPWR.t1465 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t1464 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VGND.t1134 VGND.t1132 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X136 XThR.Tn[9].t3 XThR.XTB2.Y a_n997_3755# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X137 XThC.Tn[0].t2 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1937 VGND.t508 VGND.t507 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X139 XThC.Tn[5].t6 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X140 VGND.t1286 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X141 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t1736 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X142 VGND.t380 Vbias.t24 XA.XIR[9].XIC[2].icell.SM VGND.t379 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X143 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t3 VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X144 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X145 XThC.Tn[7].t3 XThC.XTBN.Y.t14 VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X146 XThC.Tn[2].t5 XThC.XTBN.Y.t15 VGND.t675 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 VGND.t784 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t783 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X148 a_n997_1579# XThR.XTBN.Y.t10 VGND.t581 VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X149 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t2270 VGND.t2269 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X150 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t2272 VGND.t2271 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1437 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t228 VGND.t2396 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X153 VGND.t643 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X154 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X155 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t105 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X156 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t868 VGND.t867 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t831 VGND.t830 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X159 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X160 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t1927 VGND.t1926 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t252 VGND.t2597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X162 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t154 VGND.t1658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t17 VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X164 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1922 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t1467 VPWR.t1466 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X166 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t139 VGND.t1577 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X167 XA.XIR[15].XIC[0].icell.Ien VPWR.t1434 VPWR.t1436 VPWR.t1435 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X168 VGND.t382 Vbias.t25 XA.XIR[8].XIC_15.icell.SM VGND.t381 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X169 VGND.t2505 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t2504 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X170 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1431 VPWR.t1433 VPWR.t1432 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X171 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t2280 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X172 VGND.t1662 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t1661 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X173 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t523 VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X174 VGND.t676 XThC.XTBN.Y.t16 XThC.Tn[1].t7 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VGND.t384 Vbias.t26 XA.XIR[1].XIC[5].icell.SM VGND.t383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X176 VPWR.t1469 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t1468 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X177 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t1765 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X178 XA.XIR[2].XIC_15.icell.PUM VPWR.t1429 XA.XIR[2].XIC_15.icell.Ien VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X180 VPWR.t1892 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t1891 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X181 VPWR.t1039 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t1038 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VGND.t386 Vbias.t27 XA.XIR[4].XIC[6].icell.SM VGND.t385 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X183 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1938 VGND.t510 VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X184 VPWR.t1428 VPWR.t1426 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1427 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X185 VPWR.t342 XThC.XTBN.Y.t17 XThC.Tn[10].t1 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VGND.t583 XThR.XTBN.Y.t11 XThR.Tn[3].t7 VGND.t582 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t2594 VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X188 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t458 VPWR.t457 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X189 XThR.Tn[0].t6 XThR.XTBN.Y.t12 a_n1049_8581# VPWR.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X191 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t85 VGND.t835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X192 VPWR.t622 VGND.t2689 XA.XIR[0].XIC[8].icell.PUM VPWR.t621 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X193 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t1494 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X194 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XThC.Tn[12].t6 XThC.XTB5.Y VPWR.t682 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X196 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t1809 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X197 XThR.Tn[11].t11 XThR.XTBN.Y.t13 VPWR.t287 VPWR.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t801 VPWR.t800 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X199 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t2592 VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X200 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t898 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t1929 VGND.t1928 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t1574 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X203 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t2499 VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X204 VGND.t2442 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t2441 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t440 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XThR.Tn[2].t2 XThR.XTBN.Y.t14 VGND.t585 VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VGND.t2444 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t2443 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X208 VGND.t1131 VGND.t1129 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X209 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t1471 VPWR.t1470 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X210 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1670 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X211 VPWR.t288 XThR.XTBN.Y.t15 XThR.Tn[12].t3 VPWR.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X212 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t833 VGND.t832 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X213 XThC.XTB7.A data[0].t0 VPWR.t233 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 VPWR.t1894 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t1893 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X215 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t1766 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X216 VGND.t388 Vbias.t28 XA.XIR[4].XIC[10].icell.SM VGND.t387 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X217 XA.XIR[0].XIC[13].icell.PDM VGND.t1126 VGND.t1128 VGND.t1127 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X218 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 VGND.t1322 VPWR.t1939 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t1321 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t2267 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t390 Vbias.t29 XA.XIR[11].XIC[8].icell.SM VGND.t389 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X222 XThC.Tn[9].t3 XThC.XTB2.Y a_7875_9569# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 VGND.t645 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X224 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t768 VPWR.t767 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X225 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1940 VGND.t1324 VGND.t1323 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X226 VGND.t2149 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t2148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t1760 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t1759 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t1326 VPWR.t1941 XA.XIR[3].XIC_15.icell.PDM VGND.t1325 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 a_n1319_5611# XThR.XTB6.A VPWR.t35 VPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X230 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X231 VGND.t587 XThR.XTBN.Y.t16 a_n997_3979# VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X232 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t72 VGND.t715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X233 VPWR.t344 XThC.XTBN.Y.t18 XThC.Tn[14].t3 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 VGND.t392 Vbias.t30 XA.XIR[1].XIC[0].icell.SM VGND.t391 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X235 VPWR.t1473 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t1472 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X236 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X237 VGND.t394 Vbias.t31 XA.XIR[4].XIC[1].icell.SM VGND.t393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X238 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t1642 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X239 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t1643 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t803 VPWR.t802 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X241 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t2590 VGND.t2589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X242 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t460 VPWR.t459 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X243 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t900 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X244 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t10 VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X245 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t454 VPWR.t453 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X246 VGND.t396 Vbias.t32 XA.XIR[2].XIC[14].icell.SM VGND.t395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X247 VGND.t2599 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t2598 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X248 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t2501 VGND.t2500 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 VPWR.t554 XThR.XTB4.Y a_n1049_6699# VPWR.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X250 VGND.t1328 VPWR.t1942 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t1327 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X251 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t174 VGND.t1816 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X252 VPWR.t620 VGND.t2690 XA.XIR[0].XIC[3].icell.PUM VPWR.t619 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X253 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t1898 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X254 VPWR.t991 XThC.XTB6.Y a_5949_9615# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VPWR.t968 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X256 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t2502 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X257 VPWR.t909 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t908 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X258 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t1690 VPWR.t1689 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X259 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t2581 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X260 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t30 VGND.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X261 VGND.t398 Vbias.t33 XA.XIR[5].XIC[7].icell.SM VGND.t397 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X262 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t325 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X263 VGND.t605 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t1239 XThR.XTB7.B a_n1335_8107# VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VPWR.t867 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t866 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X266 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X267 VPWR.t1425 VPWR.t1423 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X268 VGND.t607 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X269 VGND.t400 Vbias.t34 XA.XIR[8].XIC[8].icell.SM VGND.t399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X270 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t869 VPWR.t868 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X271 XThC.XTB4.Y.t1 XThC.XTB7.B VPWR.t561 VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X272 VGND.t1125 VGND.t1123 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X273 VGND.t159 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t158 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X274 VPWR.t1364 VPWR.t1362 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X275 XThR.Tn[2].t8 XThR.XTB3.Y VGND.t711 VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X276 VGND.t589 XThR.XTBN.Y.t17 a_n997_2891# VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 VPWR.t1896 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t1895 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X278 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t98 VGND.t974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X279 VPWR.t860 XThR.XTB5.Y XThR.Tn[12].t11 VPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t1919 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X281 VGND.t2631 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t2630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t402 Vbias.t35 XA.XIR[11].XIC[3].icell.SM VGND.t401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X283 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t901 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X284 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t75 VGND.t722 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X285 VGND.t591 XThR.XTBN.Y.t18 XThR.Tn[6].t11 VGND.t590 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t1705 VGND.t1704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X287 VPWR.t290 XThR.XTBN.Y.t19 XThR.Tn[9].t10 VPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t143 VGND.t1581 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X289 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X290 VGND.t1122 VGND.t1120 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X291 XA.XIR[14].XIC_15.icell.PUM VPWR.t1421 XA.XIR[14].XIC_15.icell.Ien VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X292 a_n997_715# XThR.XTBN.Y.t20 VGND.t2567 VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X293 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t1899 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X294 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XThC.Tn[1].t6 XThC.XTBN.Y.t19 VGND.t677 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 VPWR.t911 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t910 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X297 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X298 XThR.Tn[14].t7 XThR.XTB7.Y VPWR.t147 VPWR.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t195 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X300 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t179 VGND.t1822 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X301 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t87 VGND.t840 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[7].XIC_15.icell.PDM VPWR.t1943 VGND.t1330 VGND.t1329 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X303 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t204 VGND.t2028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X304 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t1899 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X305 VGND.t2157 Vbias.t36 XA.XIR[15].XIC[12].icell.SM VGND.t2156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X306 VGND.t2159 Vbias.t37 XA.XIR[14].XIC[13].icell.SM VGND.t2158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t2588 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X308 VPWR.t871 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t870 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X309 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t2132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X310 VPWR.t859 XThR.XTB5.Y a_n1049_6405# VPWR.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X311 VPWR.t1543 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1542 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X312 XThR.XTB7.B data[6].t0 VPWR.t259 VPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X313 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X314 VPWR.t226 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t58 VGND.t493 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X316 VGND.t2161 Vbias.t38 XA.XIR[5].XIC[2].icell.SM VGND.t2160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X317 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t1041 VPWR.t1040 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X318 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1359 VPWR.t1361 VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 VGND.t63 XThR.XTB2.Y XThR.Tn[1].t3 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t2289 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X321 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t1994 VGND.t1993 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X322 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t191 VGND.t1921 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X323 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t1245 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t226 VGND.t2393 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X325 VGND.t2163 Vbias.t39 XA.XIR[8].XIC[3].icell.SM VGND.t2162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X326 XA.XIR[15].XIC[13].icell.Ien VPWR.t1418 VPWR.t1420 VPWR.t1419 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X327 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t177 VGND.t1820 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X328 VPWR.t1848 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t1847 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X329 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1944 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t1331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X330 VPWR.t1043 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t1042 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X331 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t1645 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X332 a_n1049_7787# XThR.XTBN.Y.t21 XThR.Tn[1].t11 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X333 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t103 VGND.t1138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X334 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X335 VGND.t678 XThC.XTBN.Y.t20 XThC.Tn[4].t7 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X336 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X337 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t137 VGND.t1526 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X338 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t140 VGND.t1578 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1416 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1417 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X340 VGND.t1119 VGND.t1117 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X341 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t1799 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X342 VGND.t548 data[1].t1 a_8739_10571# VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 XA.XIR[0].XIC[1].icell.PDM VGND.t1114 VGND.t1116 VGND.t1115 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X344 VPWR.t51 XThR.XTB2.Y XThR.Tn[9].t7 VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND.t2569 XThR.XTBN.Y.t22 XThR.Tn[7].t2 VGND.t2568 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VGND.t2601 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t2600 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X347 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t251 VGND.t2596 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X348 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1945 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t1332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X349 XThR.Tn[13].t3 XThR.XTBN.Y.t23 VPWR.t1885 VPWR.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X350 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t1901 VGND.t1900 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X351 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t210 VGND.t2294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X352 VGND.t2165 Vbias.t40 XA.XIR[10].XIC[11].icell.SM VGND.t2164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X353 VGND.t1113 VGND.t1111 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t1045 VPWR.t1044 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X355 VPWR.t1535 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X356 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1413 VPWR.t1415 VPWR.t1414 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X357 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t1475 VPWR.t1474 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 VPWR.t462 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t461 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X359 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t926 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X360 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1365 VPWR.t1367 VPWR.t1366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X361 VPWR.t1850 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t1849 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X362 VGND.t2342 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t2341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X363 VGND.t1260 XThR.XTB6.Y XThR.Tn[5].t11 VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t296 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X365 XThR.Tn[9].t2 XThR.XTB2.Y a_n997_3755# VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 VGND.t2167 Vbias.t41 XA.XIR[1].XIC[14].icell.SM VGND.t2166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X367 XThR.XTB6.Y XThR.XTB6.A VGND.t52 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X368 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1946 VGND.t1334 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X369 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t20 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X370 a_n997_1579# XThR.XTBN.Y.t24 VGND.t2570 VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 VGND.t1687 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t1686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X372 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t6 VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X373 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t1313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X374 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t1314 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 VPWR.t525 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X376 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1411 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1412 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X377 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X378 VPWR.t11 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X379 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X380 XA.XIR[15].XIC[6].icell.Ien VPWR.t1408 VPWR.t1410 VPWR.t1409 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X381 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1947 VGND.t1336 VGND.t1335 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X382 VGND.t2169 Vbias.t42 XA.XIR[10].XIC[9].icell.SM VGND.t2168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X383 VPWR.t1477 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t1476 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X384 VPWR.t888 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t887 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 XA.XIR[15].XIC[9].icell.PDM VPWR.t1948 XA.XIR[15].XIC[9].icell.Ien VGND.t1337 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X386 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t716 VPWR.t715 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X387 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t1903 VGND.t1902 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X388 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t903 VGND.t902 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1949 VGND.t1339 VGND.t1338 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 VPWR.t1876 XThR.XTBN.A XThR.XTBN.Y.t3 VPWR.t1875 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X392 VPWR.t1852 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t1851 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X393 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t2281 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X394 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t323 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X395 VPWR.t527 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X396 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t113 VGND.t1281 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X397 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t1737 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X398 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1406 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1407 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 a_3523_10575# XThC.XTB7.B VGND.t964 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X401 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t883 VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X402 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t885 VGND.t884 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t1900 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t155 VGND.t1659 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X405 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t1860 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X406 VPWR.t949 XThC.XTBN.Y.t21 XThC.Tn[13].t3 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X408 VGND.t2171 Vbias.t43 XA.XIR[13].XIC[5].icell.SM VGND.t2170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X409 VGND.t338 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t337 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X410 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t1479 VPWR.t1478 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X411 XThC.Tn[5].t11 XThC.XTB6.Y VGND.t1858 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t1285 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t886 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X414 VGND.t1341 VPWR.t1950 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t1340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X415 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t1315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X416 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t529 VPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X417 VPWR.t531 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X418 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t1472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X419 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t11 VGND.t1258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 VPWR.t13 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X421 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X422 VPWR.t1898 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t1897 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X423 XA.XIR[15].XIC[1].icell.Ien VPWR.t1403 VPWR.t1405 VPWR.t1404 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X424 VGND.t2173 Vbias.t44 XA.XIR[11].XIC[12].icell.SM VGND.t2172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X425 VGND.t2175 Vbias.t45 XA.XIR[7].XIC_15.icell.SM VGND.t2174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1400 VPWR.t1402 VPWR.t1401 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X427 VGND.t2507 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t2506 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X428 VGND.t1465 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t1464 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t2 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 XThC.Tn[4].t6 XThC.XTBN.Y.t22 VGND.t1795 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VPWR.t1692 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t1691 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X432 a_n1049_5317# XThR.XTB7.Y VPWR.t145 VPWR.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X434 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t81 VGND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X435 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t905 VGND.t904 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X436 VGND.t2177 Vbias.t46 XA.XIR[10].XIC[4].icell.SM VGND.t2176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VGND.t1110 VGND.t1108 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VPWR.t890 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t889 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X439 VPWR.t499 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t498 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 XThC.XTB6.Y XThC.XTB7.B VGND.t963 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VPWR.t1399 VPWR.t1397 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X442 XA.XIR[15].XIC[4].icell.PDM VPWR.t1951 XA.XIR[15].XIC[4].icell.Ien VGND.t1342 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X443 VPWR.t718 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t717 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X444 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1952 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X445 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t1859 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X447 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t2135 VGND.t2134 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X448 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t1921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t16 VGND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X450 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t623 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X451 XThC.Tn[13].t11 XThC.XTB6.Y VPWR.t990 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X452 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t18 VGND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X453 VGND.t1796 XThC.XTBN.Y.t24 XThC.Tn[0].t7 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 XThR.Tn[3].t11 XThR.XTBN.Y.t25 a_n1049_6699# VPWR.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t887 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X456 VGND.t2344 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t2343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X457 VGND.t955 XThR.XTB4.Y XThR.Tn[3].t3 VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X459 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t2137 VGND.t2136 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X460 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t83 VGND.t826 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X462 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t196 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X463 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t889 VGND.t888 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t7 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X465 XA.XIR[0].XIC_15.icell.PDM VPWR.t1953 VGND.t1345 VGND.t1344 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X466 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t17 VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X467 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t2583 VGND.t2582 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X468 VGND.t2179 Vbias.t47 XA.XIR[13].XIC[0].icell.SM VGND.t2178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X469 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t184 VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X470 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t1901 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X471 VGND.t928 Vbias.t48 XA.XIR[8].XIC[12].icell.SM VGND.t927 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X472 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t15 VGND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X473 XThR.Tn[11].t3 XThR.XTB4.Y VPWR.t552 VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X474 VGND.t1467 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t1466 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X475 VGND.t2509 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t2508 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 XThC.Tn[14].t7 XThC.XTB7.Y a_10915_9569# VGND.t1596 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 VPWR.t1694 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X478 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t533 VPWR.t532 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X479 VGND.t420 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t419 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X480 VPWR.t501 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t500 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X481 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X482 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t297 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X483 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1954 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t1346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X484 VPWR.t1396 VPWR.t1394 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1395 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X485 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t562 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X486 VGND.t475 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VPWR.t386 XThC.XTB2.Y XThC.Tn[9].t6 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X488 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t1854 VPWR.t1853 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X489 VGND.t1762 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t1761 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X490 VGND.t930 Vbias.t49 XA.XIR[6].XIC[11].icell.SM VGND.t929 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X491 VGND.t1348 VPWR.t1955 XA.XIR[2].XIC_15.icell.PDM VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X492 VPWR.t858 XThR.XTB5.Y XThR.Tn[12].t10 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VGND.t1689 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t1688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X494 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t5 VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X495 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t355 VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X496 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t892 VPWR.t891 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t1960 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X498 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t843 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X499 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t844 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 VPWR.t143 XThR.XTB7.Y XThR.Tn[14].t6 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t2139 VGND.t2138 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X502 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X503 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t900 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X504 XThR.Tn[8].t8 XThR.XTB1.Y.t4 a_n997_3979# VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t442 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X506 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t2390 VGND.t2389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 VGND.t1647 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1956 VGND.t1350 VGND.t1349 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 VPWR.t720 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t719 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X510 VPWR.t779 data[2].t0 XThC.XTB7.B VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X511 VGND.t1107 VGND.t1105 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t1106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X512 VPWR.t1023 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t1022 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X513 VGND.t786 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X514 XThC.Tn[13].t6 XThC.XTB6.Y a_10051_9569# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X515 XThR.Tn[4].t3 XThR.XTBN.Y.t26 a_n1049_6405# VPWR.t1886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X517 VGND.t932 Vbias.t50 XA.XIR[4].XIC[7].icell.SM VGND.t931 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X518 XThC.Tn[8].t3 XThC.XTBN.Y.t25 VPWR.t951 VPWR.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X519 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t14 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X520 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t872 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t690 VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X523 VGND.t2151 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t2150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X524 VGND.t934 Vbias.t51 XA.XIR[7].XIC[8].icell.SM VGND.t933 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X525 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t464 VPWR.t463 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X526 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t1856 VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t406 VGND.t405 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X528 VGND.t968 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t967 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t936 Vbias.t52 XA.XIR[6].XIC[9].icell.SM VGND.t935 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X530 VGND.t938 Vbias.t53 XA.XIR[3].XIC[11].icell.SM VGND.t937 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 XThC.Tn[8].t6 XThC.XTB1.Y.t4 a_7651_9569# VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 XThC.Tn[13].t2 XThC.XTBN.Y.t26 VPWR.t952 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X533 VGND.t1764 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t1763 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X534 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t357 VPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X535 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t169 VGND.t1802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X536 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t170 VGND.t1803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 VPWR.t618 VGND.t2691 XA.XIR[0].XIC[9].icell.PUM VPWR.t617 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X538 VGND.t1857 XThC.XTB6.Y XThC.Tn[5].t10 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t1738 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X540 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1379 VPWR.t1381 VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X541 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t1943 VGND.t1942 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X542 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t1945 VGND.t1944 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t15 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X544 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t1641 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X545 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t298 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 VGND.t940 Vbias.t54 XA.XIR[12].XIC[5].icell.SM VGND.t939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X548 VGND.t340 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t339 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X549 a_n1049_5611# XThR.XTB6.Y VPWR.t648 VPWR.t144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 XA.XIR[13].XIC_15.icell.PUM VPWR.t1392 XA.XIR[13].XIC_15.icell.Ien VPWR.t1393 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X551 XThR.Tn[10].t3 XThR.XTB3.Y a_n997_2891# VGND.t709 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X552 VGND.t942 Vbias.t55 XA.XIR[15].XIC[6].icell.SM VGND.t941 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X553 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t2290 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X554 VGND.t647 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X555 VGND.t1691 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t1690 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VPWR.t954 XThC.XTBN.Y.t27 XThC.Tn[7].t6 VPWR.t953 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t845 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X558 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t2140 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 VPWR.t1025 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1024 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X560 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1390 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1391 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X561 VPWR.t49 XThR.XTB2.Y XThR.Tn[9].t6 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X563 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t327 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X564 VPWR.t1032 bias[1].t0 Vbias.t10 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.1275 pd=1.15 as=0.1955 ps=1.31 w=0.85 l=1
X565 VGND.t944 Vbias.t56 XA.XIR[9].XIC[5].icell.SM VGND.t943 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X566 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t894 VPWR.t893 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X567 VGND.t609 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X568 VPWR.t1063 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t1062 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X569 VPWR.t722 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t721 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X570 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t2291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X571 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1545 VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X572 VGND.t946 Vbias.t57 XA.XIR[3].XIC[9].icell.SM VGND.t945 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X573 VGND.t970 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t969 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X574 XA.XIR[15].XIC_15.icell.Ien VPWR.t1387 VPWR.t1389 VPWR.t1388 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X575 VPWR.t1027 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1026 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X576 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t1608 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X577 VPWR.t1858 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t1857 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X578 a_n1049_7493# XThR.XTBN.Y.t27 XThR.Tn[2].t11 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X579 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t1679 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X580 XThC.Tn[0].t6 XThC.XTBN.Y.t29 VGND.t1797 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X581 VGND.t948 Vbias.t58 XA.XIR[4].XIC[2].icell.SM VGND.t947 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X582 VPWR.t1386 VPWR.t1384 XA.XIR[9].XIC_15.icell.PUM VPWR.t1385 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X583 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t531 VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X584 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t533 VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X585 VGND.t950 Vbias.t59 XA.XIR[7].XIC[3].icell.SM VGND.t949 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X586 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t10 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X587 XThR.Tn[0].t1 XThR.XTB1.Y.t5 VGND.t473 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X588 VGND.t2571 XThR.XTBN.Y.t28 XThR.Tn[5].t6 VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t235 VGND.t2432 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X590 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t164 VPWR.t163 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X591 VGND.t1168 Vbias.t60 XA.XIR[6].XIC[4].icell.SM VGND.t1167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X592 XThR.Tn[14].t3 XThR.XTB7.Y a_n997_715# VGND.t235 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X593 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t408 VGND.t407 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X594 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t1318 VGND.t1317 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 VGND.t1170 Vbias.t61 XA.XIR[15].XIC[10].icell.SM VGND.t1169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X596 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t359 VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X597 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t1905 VGND.t1904 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X598 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t63 VGND.t599 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X599 VGND.t1352 VPWR.t1957 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t1351 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X600 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t846 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X601 VGND.t2572 XThR.XTBN.Y.t29 XThR.Tn[4].t7 VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X602 VPWR.t834 bias[1].t1 Vbias.t8 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.1275 pd=1.15 as=0.1955 ps=1.31 w=0.85 l=1
X603 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t1947 VGND.t1946 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t1739 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X605 VGND.t1354 VPWR.t1958 XA.XIR[14].XIC_15.icell.PDM VGND.t1353 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t6 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t1902 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 VGND.t1172 Vbias.t62 XA.XIR[12].XIC[0].icell.SM VGND.t1171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X609 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t157 VGND.t1663 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X610 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1382 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1383 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X611 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t1903 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t1174 Vbias.t63 XA.XIR[15].XIC[1].icell.SM VGND.t1173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X613 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X614 VGND.t342 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t341 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VGND.t1192 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t1191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X616 VGND.t1176 Vbias.t64 XA.XIR[10].XIC[13].icell.SM VGND.t1175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1547 VPWR.t1546 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X618 VGND.t422 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t421 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VPWR.t1065 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t1064 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X620 VGND.t1178 Vbias.t65 XA.XIR[13].XIC[14].icell.SM VGND.t1177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t186 VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X622 VGND.t1798 XThC.XTBN.Y.t31 a_8739_9569# VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 VGND.t2603 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t2602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X624 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1959 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t1355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X625 VGND.t1180 Vbias.t66 XA.XIR[9].XIC[0].icell.SM VGND.t1179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X626 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t1774 VPWR.t1773 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X627 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t896 VPWR.t895 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X628 VGND.t1182 Vbias.t67 XA.XIR[0].XIC_15.icell.SM VGND.t1181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X629 VGND.t1469 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X630 VGND.t2511 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t2510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1549 VPWR.t1548 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X632 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t1320 VGND.t1319 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X633 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t180 VGND.t1823 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X634 a_9827_9569# XThC.XTBN.Y.t32 VGND.t1799 VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X635 VGND.t1184 Vbias.t68 XA.XIR[3].XIC[4].icell.SM VGND.t1183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X636 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t229 VGND.t2410 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X637 VPWR.t1624 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X638 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t1680 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X639 VPWR.t251 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X640 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1960 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t1356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X641 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t194 VGND.t1924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X642 VPWR.t1776 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t1775 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X643 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t1995 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X644 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t1949 VGND.t1948 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X645 VPWR.t1378 VPWR.t1376 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1377 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X646 XA.XIR[15].XIC[13].icell.PDM VPWR.t1961 XA.XIR[15].XIC[13].icell.Ien VGND.t1357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X647 VGND.t2337 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X648 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t536 VGND.t535 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X649 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t73 VGND.t716 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X650 XThR.XTB7.A data[5].t1 VPWR.t1553 VPWR.t1552 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X651 VGND.t788 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t787 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X652 VPWR.t188 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X653 VGND.t764 XThC.XTBN.A XThC.XTBN.Y.t1 VGND.t763 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X655 VPWR.t636 XThR.XTB7.B XThR.XTB1.Y.t0 VPWR.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X656 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t10 VGND.t1257 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X657 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t899 VGND.t898 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X658 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t1778 VPWR.t1777 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X659 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t9 VGND.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X660 XA.XIR[14].XIC_15.icell.PDM VPWR.t1962 VGND.t1359 VGND.t1358 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X661 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1373 VPWR.t1375 VPWR.t1374 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X662 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t47 VGND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X663 VPWR.t938 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t937 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X664 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t299 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X665 XThC.Tn[7].t5 XThC.XTBN.Y.t33 VPWR.t956 VPWR.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X666 VGND.t1238 XThR.XTB7.B a_n1335_7243# VGND.t1237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X667 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X668 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t563 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t538 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1963 VGND.t1361 VGND.t1360 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[12].XIC_15.icell.PUM VPWR.t1371 XA.XIR[12].XIC_15.icell.Ien VPWR.t1372 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t2018 VGND.t2017 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X674 VGND.t1766 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t1765 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X675 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t741 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X676 VGND.t2217 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t2216 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t50 VGND.t353 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X678 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1533 VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X679 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t57 VGND.t492 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X680 XThC.Tn[11].t7 XThC.XTB4.Y.t6 VPWR.t1830 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 VGND.t2219 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t2218 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X682 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t61 VGND.t554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X683 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1368 VPWR.t1370 VPWR.t1369 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X684 a_n997_1803# XThR.XTBN.Y.t30 VGND.t2573 VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X685 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X686 XThR.Tn[3].t10 XThR.XTBN.Y.t31 a_n1049_6699# VPWR.t1887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X687 VPWR.t361 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t360 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X688 VGND.t2574 XThR.XTBN.Y.t32 XThR.Tn[3].t6 VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 VGND.t1186 Vbias.t69 XA.XIR[11].XIC[6].icell.SM VGND.t1185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X690 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t760 VPWR.t759 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X691 VGND.t1363 VPWR.t1964 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t1362 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X692 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1965 VGND.t1365 VGND.t1364 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X693 XThC.Tn[2].t9 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X694 VPWR.t253 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X695 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t17 VPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X696 VPWR.t1780 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t1779 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X697 VPWR.t190 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 XThR.Tn[11].t2 XThR.XTB4.Y VPWR.t550 VPWR.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 VPWR.t1358 VPWR.t1356 XA.XIR[8].XIC_15.icell.PUM VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X700 VPWR.t385 XThC.XTB2.Y a_3773_9615# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X701 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t1924 VPWR.t1923 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1354 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1355 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X703 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t897 VGND.t896 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X704 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 VGND.t1188 Vbias.t70 XA.XIR[0].XIC[8].icell.SM VGND.t1187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X706 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t1489 VGND.t1488 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X707 VGND.t972 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t971 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 VGND.t1104 VGND.t1102 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t1103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X709 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t361 VGND.t360 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X710 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t692 VGND.t691 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X711 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t25 VGND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X712 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1531 VPWR.t1530 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X713 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t125 VGND.t1497 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X714 VGND.t1367 VPWR.t1966 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t1366 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X715 VPWR.t67 XThC.XTB6.A a_5949_10571# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X716 VPWR.t940 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t939 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X717 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t154 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X718 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t1740 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 VGND.t708 XThR.XTB3.Y XThR.Tn[2].t7 VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 VPWR.t19 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X721 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1741 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X722 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t1642 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t1862 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t2020 VGND.t2019 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X725 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t209 VGND.t2293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X726 XThC.XTBN.Y.t3 XThC.XTBN.A VPWR.t418 VPWR.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X727 VGND.t1190 Vbias.t71 XA.XIR[5].XIC[5].icell.SM VGND.t1189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X728 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t927 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X729 VGND.t344 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t343 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 VGND.t1963 Vbias.t72 XA.XIR[11].XIC[10].icell.SM VGND.t1962 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X731 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t762 VPWR.t761 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X732 XThR.Tn[8].t2 XThR.XTB1.Y.t7 a_n997_3979# VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X733 XA.XIR[6].XIC_15.icell.PUM VPWR.t1352 XA.XIR[6].XIC_15.icell.Ien VPWR.t1353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X734 VGND.t2369 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t2368 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t1965 Vbias.t73 XA.XIR[12].XIC[14].icell.SM VGND.t1964 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X736 VGND.t346 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X737 VGND.t1967 Vbias.t74 XA.XIR[8].XIC[6].icell.SM VGND.t1966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X738 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t724 VPWR.t723 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X739 VGND.t1369 VPWR.t1967 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t1368 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X740 VGND.t649 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X741 VGND.t2605 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t2604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t1800 XThC.XTBN.Y.t35 a_9827_9569# VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X743 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t197 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X744 VPWR.t363 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X745 VPWR.t842 XThC.XTB7.Y XThC.Tn[14].t11 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X746 XThR.Tn[4].t2 XThR.XTBN.Y.t33 a_n1049_6405# VPWR.t1887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X747 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t906 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X748 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t907 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X749 VGND.t1969 Vbias.t75 XA.XIR[11].XIC[1].icell.SM VGND.t1968 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X750 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t764 VPWR.t763 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X751 VGND.t1971 Vbias.t76 XA.XIR[7].XIC[12].icell.SM VGND.t1970 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X752 VPWR.t548 XThR.XTB4.Y a_n1049_6699# VPWR.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X753 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t166 VPWR.t165 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X754 VGND.t1973 Vbias.t77 XA.XIR[6].XIC[13].icell.SM VGND.t1972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X755 VPWR.t484 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t483 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X756 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X757 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t365 VPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X758 VGND.t1975 Vbias.t78 XA.XIR[9].XIC[14].icell.SM VGND.t1974 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X759 VPWR.t1782 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t1781 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X760 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t156 VGND.t1660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X761 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t1570 VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X762 XA.XIR[15].XIC[1].icell.PDM VPWR.t1968 XA.XIR[15].XIC[1].icell.Ien VGND.t1370 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X763 VPWR.t1067 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t1066 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X764 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t1490 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X765 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1969 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t1371 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t486 VPWR.t485 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X767 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t624 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X768 VGND.t1977 Vbias.t79 XA.XIR[0].XIC[3].icell.SM VGND.t1976 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X769 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t115 VGND.t1300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X770 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t223 VGND.t2366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X771 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t363 VGND.t362 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X772 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1529 VPWR.t1528 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X773 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t2416 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X774 VGND.t1979 Vbias.t80 XA.XIR[8].XIC[10].icell.SM VGND.t1978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X775 VPWR.t1889 XThR.XTBN.Y.t34 XThR.Tn[8].t7 VPWR.t1888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X776 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t726 VPWR.t725 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X777 XThR.Tn[10].t2 XThR.XTB3.Y a_n997_2891# VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X778 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t535 VPWR.t534 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X779 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X780 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t560 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X781 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t246 VGND.t2564 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X782 VGND.t1981 Vbias.t81 XA.XIR[5].XIC[0].icell.SM VGND.t1980 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X783 VGND.t1101 VGND.t1099 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t1100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 VGND.t1983 Vbias.t82 XA.XIR[8].XIC[1].icell.SM VGND.t1982 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X785 VPWR.t65 XThC.XTB6.A XThC.XTB2.Y VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X786 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t1693 VGND.t1692 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X787 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t1695 VGND.t1694 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X788 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t188 VGND.t1907 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X789 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t1710 VPWR.t1709 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X790 VGND.t1985 Vbias.t83 XA.XIR[3].XIC[13].icell.SM VGND.t1984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X791 VGND.t1194 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t1193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X792 VGND.t424 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 XThR.XTB3.Y XThR.XTB7.A VPWR.t455 VPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X794 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t14 VGND.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X795 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X796 VGND.t2607 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t2606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X797 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X798 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1970 VGND.t1373 VGND.t1372 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X799 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t2 VGND.t234 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X800 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t908 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X801 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X802 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t942 VPWR.t941 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X803 VGND.t1204 Vbias.t84 XA.XIR[2].XIC[11].icell.SM VGND.t1203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X804 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t225 VGND.t2383 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X805 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t488 VPWR.t487 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X806 XThR.Tn[0].t10 XThR.XTBN.Y.t35 VGND.t2575 VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X807 VPWR.t857 XThR.XTB5.Y a_n1049_6405# VPWR.t547 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X808 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t1784 VPWR.t1783 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X809 VGND.t1206 Vbias.t85 XA.XIR[14].XIC_15.icell.SM VGND.t1205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X810 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t12 VGND.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X811 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X812 XThC.Tn[10].t0 XThC.XTB3.Y.t4 VPWR.t153 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t364 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X814 VPWR.t1890 XThR.XTBN.Y.t36 XThR.Tn[10].t11 VPWR.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t2006 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X816 VPWR.t903 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t902 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X817 VPWR.t1749 XThC.XTBN.Y.t36 XThC.Tn[13].t1 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X818 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t693 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X819 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t2021 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X820 a_3773_9615# XThC.XTB2.Y VPWR.t384 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X821 XThC.Tn[5].t9 XThC.XTB6.Y VGND.t1856 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t211 VGND.t2300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X823 XThC.Tn[2].t0 XThC.XTB3.Y.t5 VGND.t336 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X824 VPWR.t1069 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t1068 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X825 VPWR.t1527 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1526 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X826 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t412 VGND.t411 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X827 VGND.t790 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t789 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X828 VPWR.t466 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t465 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X829 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t133 VGND.t1513 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X830 VPWR.t168 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t167 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X831 VGND.t725 XThR.XTBN.Y.t37 a_n997_3755# VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X833 VPWR.t1731 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t1730 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t695 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X835 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1971 VGND.t1375 VGND.t1374 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X836 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t1884 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X837 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t944 VPWR.t943 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X838 VGND.t1208 Vbias.t86 XA.XIR[2].XIC[9].icell.SM VGND.t1207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X839 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X840 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t159 VGND.t1667 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X841 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t1697 VGND.t1696 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X842 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t128 VGND.t1507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X843 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t1227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t64 VGND.t638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t198 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X846 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t207 VGND.t2089 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X847 VGND.t1649 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t1648 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X848 XA.XIR[11].XIC_15.icell.PDM VPWR.t1972 VGND.t1377 VGND.t1376 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t147 VGND.t1597 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X850 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t365 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X851 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t2307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t21 VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X853 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X854 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t928 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X855 a_5155_9615# XThC.XTB5.Y VPWR.t681 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X856 XA.XIR[5].XIC_15.icell.PUM VPWR.t1350 XA.XIR[5].XIC_15.icell.Ien VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X857 VPWR.t905 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t904 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X858 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t848 VGND.t847 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X859 a_n1049_7493# XThR.XTB3.Y VPWR.t379 VPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X860 VGND.t2371 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t2370 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X861 XA.XIR[9].XIC_15.icell.PUM VPWR.t1348 XA.XIR[9].XIC_15.icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X862 VGND.t2153 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t2152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X863 VPWR.t1525 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X864 VPWR.t468 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t467 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X865 VGND.t1379 VPWR.t1973 XA.XIR[13].XIC_15.icell.PDM VGND.t1378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X866 XThC.Tn[8].t11 XThC.XTB1.Y.t7 VPWR.t1733 VPWR.t1732 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X867 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t1665 VPWR.t1664 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X868 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t1071 VPWR.t1070 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X869 VGND.t1628 XThR.XTB5.Y XThR.Tn[4].t11 VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X870 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t11 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X871 VGND.t1381 VPWR.t1974 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t1380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X872 VPWR.t1073 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t1072 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X873 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t416 VGND.t415 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t1523 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1522 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XThR.XTB5.Y XThR.XTB5.A VGND.t1801 VGND.t51 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X876 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t1699 VGND.t1698 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X877 VPWR.t470 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t469 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X878 VPWR.t946 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t945 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X879 VPWR.t170 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t169 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t444 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X881 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t1818 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X882 VPWR.t1322 VPWR.t1320 XA.XIR[1].XIC_15.icell.PUM VPWR.t1321 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X883 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t2256 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X884 VPWR.t1347 VPWR.t1345 XA.XIR[5].XIC_15.icell.PUM VPWR.t1346 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[15].XIC_15.icell.PDM VPWR.t1975 XA.XIR[15].XIC_15.icell.Ien VGND.t1382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X886 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t850 VGND.t849 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X887 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t948 VPWR.t947 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X888 VGND.t1210 Vbias.t87 XA.XIR[2].XIC[4].icell.SM VGND.t1209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X889 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t32 VGND.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X890 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t1478 VGND.t1477 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X891 VGND.t1212 Vbias.t88 XA.XIR[15].XIC[7].icell.SM VGND.t1211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X892 VGND.t1384 VPWR.t1976 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t1383 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t1214 Vbias.t89 XA.XIR[14].XIC[8].icell.SM VGND.t1213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X894 VGND.t611 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X895 VPWR.t1344 VPWR.t1342 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X896 XThC.Tn[14].t6 XThC.XTB7.Y a_10915_9569# VGND.t1595 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X897 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X898 a_n997_1803# XThR.XTBN.Y.t38 VGND.t727 VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t1904 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X900 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t1075 VPWR.t1074 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X901 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t1886 VGND.t1885 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t11 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X903 VGND.t2373 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2372 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t111 VGND.t1261 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X905 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t1888 VGND.t1887 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 VGND.t1216 Vbias.t90 XA.XIR[5].XIC[14].icell.SM VGND.t1215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X907 VGND.t2609 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t2608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X908 VPWR.t832 XThC.XTB5.A XThC.XTB1.Y.t2 VPWR.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X909 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1977 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X910 VGND.t131 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X911 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1978 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t1386 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t1794 VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t1700 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 VGND.t1218 Vbias.t91 XA.XIR[1].XIC[11].icell.SM VGND.t1217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X915 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t1667 VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X916 VGND.t1220 Vbias.t92 XA.XIR[0].XIC[12].icell.SM VGND.t1219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X917 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t1796 VPWR.t1795 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X918 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X919 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1340 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X920 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1521 VPWR.t1520 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X921 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t86 VGND.t839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X922 VGND.t1275 XThC.XTB3.Y.t6 XThC.Tn[2].t1 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t329 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X924 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t2 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X925 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t2022 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X926 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t2257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X927 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t2397 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X928 a_n1319_6405# XThR.XTB5.A VPWR.t960 VPWR.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X929 VPWR.t993 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t992 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X930 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t2478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X931 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t564 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X932 VPWR.t1339 VPWR.t1337 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X933 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t4 VGND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X934 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t1735 VPWR.t1734 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X935 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t490 VPWR.t489 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X936 VGND.t1222 Vbias.t93 XA.XIR[15].XIC[2].icell.SM VGND.t1221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X937 VGND.t1224 Vbias.t94 XA.XIR[14].XIC[3].icell.SM VGND.t1223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X938 XThR.Tn[12].t2 XThR.XTBN.Y.t39 VPWR.t388 VPWR.t286 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X939 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X940 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1334 VPWR.t1336 VPWR.t1335 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X941 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t253 VGND.t2614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X942 XThC.Tn[11].t3 XThC.XTBN.Y.t39 VPWR.t1750 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X943 VGND.t1247 data[4].t2 XThR.XTB5.A VGND.t1246 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X944 XThR.XTBN.Y.t1 XThR.XTBN.A VGND.t2529 VGND.t2528 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X945 VGND.t1499 data[3].t0 XThC.XTBN.A VGND.t1498 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X946 VGND.t1226 Vbias.t95 XA.XIR[1].XIC[9].icell.SM VGND.t1225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X947 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1979 VGND.t1388 VGND.t1387 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X948 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t2024 VGND.t2023 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X949 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t7 VGND.t1258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X950 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t1890 VGND.t1889 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t201 VGND.t1997 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X952 XA.XIR[10].XIC_15.icell.PDM VPWR.t1980 VGND.t1390 VGND.t1389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t192 VGND.t1922 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 a_n997_2667# XThR.XTBN.Y.t40 VGND.t728 VGND.t514 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1332 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X956 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t250 VGND.t2586 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X957 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t313 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X958 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t2142 VGND.t2141 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X959 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t2479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X960 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t874 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t565 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X962 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t2259 VGND.t2258 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 VPWR.t995 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t994 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X964 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t2026 VGND.t2025 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t743 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X966 VGND.t2221 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t2220 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X967 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t36 VGND.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X968 XThC.Tn[4].t10 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X969 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t2398 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X970 VGND.t1392 VPWR.t1981 XA.XIR[12].XIC_15.icell.PDM VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X971 VPWR.t192 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X972 VPWR.t390 XThR.XTBN.Y.t41 XThR.Tn[8].t6 VPWR.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X973 VGND.t2513 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t2512 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X974 VGND.t1471 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t1470 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X975 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t1643 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X977 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1329 VPWR.t1331 VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X978 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t5 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X979 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t1476 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X980 VGND.t1861 Vbias.t96 XA.XIR[4].XIC[5].icell.SM VGND.t1860 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X981 VPWR.t680 XThC.XTB5.Y XThC.Tn[12].t5 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1982 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t1393 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X983 VPWR.t1821 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t1820 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X984 VPWR.t1328 VPWR.t1326 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X985 VGND.t1863 Vbias.t97 XA.XIR[7].XIC[6].icell.SM VGND.t1862 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X986 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t472 VPWR.t471 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X987 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t172 VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X988 VGND.t651 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X989 VGND.t729 XThR.XTBN.Y.t42 XThR.Tn[1].t7 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X990 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t1892 VGND.t1891 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t2418 VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X992 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t367 VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X993 VPWR.t616 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t615 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X994 VPWR.t1325 VPWR.t1323 XA.XIR[4].XIC_15.icell.PUM VPWR.t1324 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X995 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t492 VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X996 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t23 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X997 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X998 VGND.t1865 Vbias.t98 XA.XIR[1].XIC[4].icell.SM VGND.t1864 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X999 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t1475 VGND.t1474 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1000 XThR.Tn[6].t2 XThR.XTB7.Y VGND.t233 VGND.t232 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1001 a_9827_9569# XThC.XTBN.Y.t41 VGND.t2351 VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1002 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t875 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1003 XThR.Tn[9].t9 XThR.XTBN.Y.t43 VPWR.t392 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1004 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t1278 VGND.t1277 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t2420 VGND.t2419 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1006 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t1658 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t1920 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1008 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t67 VGND.t698 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1009 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t871 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1010 XThC.Tn[1].t10 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1011 VGND.t1651 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t1650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1012 XThR.Tn[0].t9 XThR.XTBN.Y.t44 VGND.t730 VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 XThC.Tn[13].t5 XThC.XTB6.Y a_10051_9569# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1014 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1762 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1015 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t1473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1016 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1017 VPWR.t393 XThR.XTBN.Y.t45 XThR.Tn[10].t10 VPWR.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1018 VPWR.t369 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1019 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t929 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1020 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t2261 VGND.t2260 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1021 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1317 VPWR.t1319 VPWR.t1318 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1022 XA.XIR[0].XIC[12].icell.PDM VGND.t1096 VGND.t1098 VGND.t1097 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 VGND.t348 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1024 VGND.t2375 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2374 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1025 VGND.t1867 Vbias.t99 XA.XIR[11].XIC[7].icell.SM VGND.t1866 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1026 VGND.t1869 Vbias.t100 XA.XIR[7].XIC[10].icell.SM VGND.t1868 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1027 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t474 VPWR.t473 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1028 VPWR.t841 XThC.XTB7.Y a_6243_9615# VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1029 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t130 VGND.t1509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1030 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1983 VGND.t1395 VGND.t1394 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1031 VGND.t2377 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2376 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1032 VGND.t653 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1034 VGND.t2155 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t2154 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 VPWR.t614 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t613 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1036 VGND.t1768 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t1767 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t1492 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1038 VGND.t1397 VPWR.t1984 XA.XIR[6].XIC_15.icell.PDM VGND.t1396 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1039 VGND.t2352 XThC.XTBN.Y.t43 a_8963_9569# VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1040 VGND.t1871 Vbias.t101 XA.XIR[4].XIC[0].icell.SM VGND.t1870 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1041 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t155 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1042 VPWR.t1029 XThR.XTB1.Y.t8 XThR.Tn[8].t9 VPWR.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1043 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1315 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1044 VGND.t1873 Vbias.t102 XA.XIR[7].XIC[1].icell.SM VGND.t1872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1045 VGND.t1875 Vbias.t103 XA.XIR[2].XIC[13].icell.SM VGND.t1874 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1046 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t476 VPWR.t475 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1047 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t89 VGND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1048 VGND.t1196 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1049 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t1626 VPWR.t1625 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1050 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t1801 VPWR.t1800 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1051 VGND.t426 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1052 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t2422 VGND.t2421 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1053 XThR.XTBN.A data[7].t0 VPWR.t1568 VPWR.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1054 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t371 VPWR.t370 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1055 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t1669 VPWR.t1668 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1056 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t70 VGND.t713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1057 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1058 VPWR.t612 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t611 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1059 VPWR.t47 XThR.XTB2.Y a_n1049_7787# VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1060 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1061 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t851 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1062 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1063 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t25 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 VPWR.t1823 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t1822 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1065 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t1279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t90 VGND.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1067 XA.XIR[0].XIC[10].icell.PDM VGND.t1093 VGND.t1095 VGND.t1094 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1068 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t1599 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1069 VGND.t1877 Vbias.t104 XA.XIR[8].XIC[7].icell.SM VGND.t1876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1070 a_n1049_7493# XThR.XTBN.Y.t46 XThR.Tn[2].t9 VPWR.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t99 VGND.t975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1072 VGND.t625 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1073 XThC.Tn[8].t10 XThC.XTB1.Y.t10 VPWR.t693 VPWR.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1074 VPWR.t1009 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t1008 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1075 VPWR.t1314 VPWR.t1312 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1313 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1076 VGND.t1092 VGND.t1090 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t1091 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1077 VGND.t1616 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t1615 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1078 XThR.Tn[0].t2 XThR.XTB1.Y.t9 VGND.t842 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1079 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t2308 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1080 VGND.t1879 Vbias.t105 XA.XIR[11].XIC[2].icell.SM VGND.t1878 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1081 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t625 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1082 VPWR.t378 XThR.XTB3.Y XThR.Tn[10].t7 VPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1083 VGND.t792 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t791 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t2310 VGND.t2309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1085 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t2312 VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1086 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t71 VGND.t714 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1087 VPWR.t383 XThC.XTB2.Y a_3773_9615# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1088 VGND.t1198 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t1197 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1089 VGND.t732 XThR.XTBN.Y.t47 XThR.Tn[4].t6 VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1090 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1310 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1311 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t35 VGND.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1092 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t1864 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t1897 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1094 VPWR.t1751 XThC.XTBN.Y.t44 XThC.Tn[9].t11 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1985 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t1398 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1097 VGND.t2353 XThC.XTBN.Y.t45 XThC.Tn[5].t1 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1098 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t2400 VGND.t2399 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1099 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1100 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t216 VGND.t2318 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1101 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t144 VGND.t1582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1102 VGND.t734 XThR.XTBN.Y.t48 a_n997_1579# VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1103 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t199 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1104 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t51 VGND.t366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1105 VGND.t1881 Vbias.t106 XA.XIR[14].XIC[12].icell.SM VGND.t1880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1106 VGND.t1883 Vbias.t107 XA.XIR[10].XIC_15.icell.SM VGND.t1882 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1107 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t1 VPWR.t1752 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1108 VGND.t2515 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t2514 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1109 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1110 VGND.t919 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t2143 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VPWR.t1825 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t1824 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1113 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t850 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1114 XThC.Tn[12].t2 XThC.XTB5.Y a_9827_9569# VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1115 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1116 VPWR.t1011 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t1010 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1117 XThR.XTB6.A data[5].t2 VPWR.t182 VPWR.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1118 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t42 VGND.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1119 VPWR.t1309 VPWR.t1307 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1120 XThR.Tn[14].t1 XThR.XTB7.Y a_n997_715# VGND.t231 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1121 VPWR.t997 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t996 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1122 a_n1049_5317# XThR.XTBN.Y.t49 XThR.Tn[6].t7 VPWR.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1123 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1827 VPWR.t1826 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1124 VGND.t439 Vbias.t108 XA.XIR[8].XIC[2].icell.SM VGND.t438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1125 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t120 VGND.t1480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1126 XA.XIR[15].XIC[12].icell.Ien VPWR.t1304 VPWR.t1306 VPWR.t1305 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1127 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t206 VGND.t2030 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1128 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t24 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1129 VPWR.t1628 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t1627 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1130 VPWR.t667 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t666 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1131 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t1564 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1132 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1986 VGND.t1400 VGND.t1399 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1133 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t1601 VGND.t1600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1134 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t1659 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1135 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t1566 VGND.t1565 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t3 VGND.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1137 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t84 VGND.t827 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1138 XA.XIR[3].XIC_15.icell.PDM VPWR.t1987 VGND.t1402 VGND.t1401 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1139 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1140 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t121 VGND.t1481 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1141 a_6243_9615# XThC.XTB7.Y VPWR.t840 VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1142 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1302 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1303 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1143 VGND.t1089 VGND.t1087 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t1088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1144 XThC.Tn[10].t8 XThC.XTBN.Y.t47 VPWR.t1753 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1145 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t2144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1146 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t876 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1147 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t2402 VGND.t2401 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1148 VGND.t428 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t427 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XA.XIR[1].XIC_15.icell.PUM VPWR.t1300 XA.XIR[1].XIC_15.icell.Ien VPWR.t1301 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 XThC.Tn[10].t3 XThC.XTB3.Y.t8 a_8739_9569# VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1151 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t2146 VGND.t2145 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1152 VGND.t1594 XThC.XTB7.Y XThC.Tn[6].t11 VGND.t1593 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t145 VGND.t1583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1154 VGND.t1404 VPWR.t1988 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t1403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1155 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1989 VGND.t1406 VGND.t1405 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1156 XThR.Tn[11].t10 XThR.XTBN.Y.t50 VPWR.t396 VPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 VGND.t1630 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 VPWR.t1754 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 VGND.t1408 VPWR.t1990 XA.XIR[5].XIC_15.icell.PDM VGND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1160 XA.XIR[15].XIC[10].icell.Ien VPWR.t1297 VPWR.t1299 VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 VGND.t441 Vbias.t109 XA.XIR[13].XIC[11].icell.SM VGND.t440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1162 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t194 VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1163 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1829 VPWR.t1828 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1164 VGND.t1410 VPWR.t1991 XA.XIR[9].XIC_15.icell.PDM VGND.t1409 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1165 VPWR.t1803 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t1802 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1166 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t1645 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1167 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1294 VPWR.t1296 VPWR.t1295 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1168 VPWR.t669 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t668 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1169 VGND.t443 Vbias.t110 XA.XIR[1].XIC[13].icell.SM VGND.t442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1170 VGND.t445 Vbias.t111 XA.XIR[0].XIC[6].icell.SM VGND.t444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1171 VGND.t655 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1172 VGND.t447 Vbias.t112 XA.XIR[4].XIC[14].icell.SM VGND.t446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t2032 XThC.XTB7.A XThC.XTB7.Y VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1174 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t1568 VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1175 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1519 VPWR.t1518 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1176 VPWR.t1630 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t1629 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1177 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t6 VGND.t1257 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1178 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t97 VGND.t956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1179 a_n997_2667# XThR.XTBN.Y.t51 VGND.t735 VGND.t524 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 VPWR.t999 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t998 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1181 VPWR.t1906 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t1905 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1182 a_7875_9569# XThC.XTBN.Y.t49 VGND.t2354 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1183 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t1603 VGND.t1602 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1184 VGND.t794 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t793 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1185 VGND.t736 XThR.XTBN.Y.t52 a_n997_3979# VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1186 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t845 VPWR.t844 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1187 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t183 VGND.t1842 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1188 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1189 XThC.Tn[14].t2 XThC.XTBN.Y.t50 VPWR.t1755 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1190 a_n1049_6699# XThR.XTB4.Y VPWR.t546 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1191 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t7 VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1192 VGND.t449 Vbias.t113 XA.XIR[10].XIC[8].icell.SM VGND.t448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1193 VGND.t1618 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t1617 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1194 VGND.t451 Vbias.t114 XA.XIR[13].XIC[9].icell.SM VGND.t450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1195 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t1047 VPWR.t1046 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1196 XThC.Tn[2].t2 XThC.XTB3.Y.t9 VGND.t1276 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1197 XThC.Tn[9].t10 XThC.XTBN.Y.t52 VPWR.t228 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1198 XThC.Tn[5].t0 XThC.XTBN.Y.t53 VGND.t476 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1199 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 VGND.t453 Vbias.t115 XA.XIR[0].XIC[10].icell.SM VGND.t452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1201 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t2611 VGND.t2610 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1202 VGND.t133 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1203 XA.XIR[15].XIC[5].icell.Ien VPWR.t1291 VPWR.t1293 VPWR.t1292 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1204 VGND.t1086 VGND.t1084 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t1085 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1205 VPWR.t695 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1206 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1992 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t1411 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1207 XThC.Tn[0].t0 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1208 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 VPWR.t671 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t670 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1210 VPWR.t1908 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t1907 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1211 XThR.Tn[12].t9 XThR.XTB5.Y VPWR.t856 VPWR.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1212 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1213 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t200 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1214 VGND.t455 Vbias.t116 XA.XIR[0].XIC[1].icell.SM VGND.t454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1215 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1289 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1290 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t122 VGND.t1482 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1217 VGND.t1200 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t1199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1218 XThR.Tn[6].t10 XThR.XTBN.Y.t53 VGND.t738 VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1219 a_n1049_5611# XThR.XTBN.Y.t54 XThR.Tn[5].t2 VPWR.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1220 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1221 VGND.t1844 XThR.XTBN.Y.t55 a_n997_2891# VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1222 VGND.t1236 XThR.XTB7.B XThR.XTB7.Y VGND.t1235 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1223 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1517 VPWR.t1516 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1224 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t28 VGND.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1225 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t1751 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1226 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t2404 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1227 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t1001 VPWR.t1000 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1228 VPWR.t1003 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t1002 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1229 VGND.t1413 VPWR.t1993 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t1412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1230 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t536 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1231 VPWR.t1910 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t1909 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1232 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t7 VGND.t703 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1233 VPWR.t1288 VPWR.t1286 XA.XIR[12].XIC_15.icell.PUM VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t165 VGND.t1708 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1235 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t1013 VPWR.t1012 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1236 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1283 VPWR.t1285 VPWR.t1284 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1237 VGND.t457 Vbias.t117 XA.XIR[6].XIC_15.icell.SM VGND.t456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1238 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1239 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t96 VGND.t951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1240 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t2613 VGND.t2612 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1241 VGND.t459 Vbias.t118 XA.XIR[10].XIC[3].icell.SM VGND.t458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1242 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1280 VPWR.t1282 VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1243 VGND.t477 XThC.XTBN.Y.t55 XThC.Tn[1].t5 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 a_n1049_6405# XThR.XTB5.Y VPWR.t855 VPWR.t545 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1245 VGND.t461 Vbias.t119 XA.XIR[13].XIC[4].icell.SM VGND.t460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1246 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t1049 VPWR.t1048 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1247 VPWR.t805 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1248 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t1604 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1249 VGND.t1083 VGND.t1081 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t1082 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1250 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1994 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t1414 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t242 VPWR.t1995 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t241 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1252 VPWR.t1015 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t1014 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1253 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t1753 VGND.t1752 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t446 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1255 VPWR.t478 XThR.XTB1.Y.t10 XThR.Tn[8].t3 VPWR.t477 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1256 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t626 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1257 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t65 VGND.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1258 VPWR.t978 XThR.XTBN.Y.t56 XThR.Tn[7].t6 VPWR.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1259 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1278 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1260 VGND.t720 XThC.XTB2.Y XThC.Tn[1].t3 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1261 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1276 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1262 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t212 VGND.t2303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1263 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t2405 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1264 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t231 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t1501 VGND.t1500 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1266 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t1005 VPWR.t1004 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1267 VGND.t60 XThR.XTB2.Y XThR.Tn[1].t2 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1268 XThR.Tn[1].t10 XThR.XTBN.Y.t57 a_n1049_7787# VPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1269 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t1755 VGND.t1754 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1270 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t185 VGND.t1853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1271 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t201 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t1931 VGND.t1930 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1273 VGND.t1653 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t1652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t135 VGND.t1515 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1275 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t807 VPWR.t806 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1276 VGND.t2446 Vbias.t120 XA.XIR[3].XIC_15.icell.SM VGND.t2445 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1277 VGND.t2448 Vbias.t121 XA.XIR[12].XIC[11].icell.SM VGND.t2447 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1278 VGND.t1080 VGND.t1078 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t1079 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1279 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t1017 VPWR.t1016 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1280 VGND.t921 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t920 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1281 VGND.t2517 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t2516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1282 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t1007 VPWR.t1006 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1283 XThR.Tn[9].t5 XThR.XTB2.Y VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1284 XThR.Tn[7].t1 XThR.XTBN.Y.t58 VGND.t1846 VGND.t1845 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1285 VPWR.t769 data[1].t2 XThC.XTB6.A VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1286 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t861 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1287 VPWR.t809 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t808 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1288 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t314 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1289 VPWR.t1275 VPWR.t1273 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1274 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1290 VGND.t479 XThC.XTBN.Y.t57 a_7875_9569# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t1893 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1292 VPWR.t979 XThR.XTBN.Y.t59 XThR.Tn[13].t2 VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1293 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t771 VPWR.t770 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1294 VPWR.t1272 VPWR.t1270 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1295 VGND.t1832 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1296 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1297 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t218 VGND.t2332 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1298 VGND.t2450 Vbias.t122 XA.XIR[9].XIC[11].icell.SM VGND.t2449 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1299 VPWR.t377 XThR.XTB3.Y XThR.Tn[10].t6 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1300 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t673 VPWR.t672 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1301 VGND.t2223 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t2222 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1302 XThC.Tn[3].t6 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1303 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t2423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1304 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t2424 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1305 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t92 VPWR.t91 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1306 XThR.Tn[5].t10 XThR.XTB6.Y VGND.t1256 VGND.t1255 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1307 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1308 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1309 VPWR.t634 XThR.XTB7.B XThR.XTB4.Y VPWR.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1310 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t2587 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1311 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1312 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t1757 VGND.t1756 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1313 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t331 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1996 VGND.t244 VGND.t243 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t2305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1317 VGND.t2452 Vbias.t123 XA.XIR[12].XIC[9].icell.SM VGND.t2451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1318 VGND.t1655 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t1654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1319 VPWR.t1019 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t1018 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1320 VGND.t1077 VGND.t1075 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t1076 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1321 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t811 VPWR.t810 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1322 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t0 VGND.t230 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1323 VGND.t2379 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t2378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1324 VGND.t2454 Vbias.t124 XA.XIR[7].XIC[7].icell.SM VGND.t2453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1325 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t1805 VPWR.t1804 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1326 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t1933 VGND.t1932 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1327 VGND.t627 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1328 VGND.t2456 Vbias.t125 XA.XIR[6].XIC[8].icell.SM VGND.t2455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1329 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t125 VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1997 VGND.t246 VGND.t245 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1331 VGND.t1834 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t1833 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t264 VPWR.t263 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1333 VGND.t1632 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t1631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1335 VGND.t2458 Vbias.t126 XA.XIR[9].XIC[9].icell.SM VGND.t2457 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1336 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t675 VPWR.t674 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1337 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t80 VGND.t774 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1338 VPWR.t55 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t54 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1339 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1340 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1763 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1341 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t1894 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1342 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t109 VGND.t108 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t111 VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1344 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t773 VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1345 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t31 VGND.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1346 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1347 VGND.t2460 Vbias.t127 XA.XIR[15].XIC[5].icell.SM VGND.t2459 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1348 VGND.t2462 Vbias.t128 XA.XIR[14].XIC[6].icell.SM VGND.t2461 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1349 VGND.t1670 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t1669 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1350 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1351 VGND.t248 VPWR.t1998 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t247 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t2425 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1353 XThC.Tn[1].t4 XThC.XTBN.Y.t59 VGND.t480 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1354 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1356 VPWR.t1269 VPWR.t1267 XA.XIR[15].XIC_15.icell.PUM VPWR.t1268 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1357 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1358 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t1605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1359 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t94 VPWR.t93 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1360 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t1 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1361 VPWR.t1515 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1362 VGND.t2464 Vbias.t129 XA.XIR[3].XIC[8].icell.SM VGND.t2463 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1363 VGND.t629 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t628 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1364 XA.XIR[15].XIC[14].icell.Ien VPWR.t1264 VPWR.t1266 VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1365 VGND.t2466 Vbias.t130 XA.XIR[12].XIC[4].icell.SM VGND.t2465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1366 VPWR.t1021 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t1020 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1367 VGND.t1620 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t1619 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1368 VPWR.t69 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 VPWR.t1263 VPWR.t1261 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1262 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1370 XThR.Tn[13].t9 XThR.XTB6.Y a_n997_1579# VGND.t1254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1371 a_n1049_8581# XThR.XTBN.Y.t60 XThR.Tn[0].t5 VPWR.t980 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1372 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t973 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1373 VPWR.t657 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t656 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1374 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1375 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t2407 VGND.t2406 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1376 VGND.t2468 Vbias.t131 XA.XIR[7].XIC[2].icell.SM VGND.t2467 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1377 VGND.t1441 Vbias.t132 XA.XIR[6].XIC[3].icell.SM VGND.t1440 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1378 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t152 VGND.t1639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1379 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t128 VGND.t127 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1380 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t52 VGND.t368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1381 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t862 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 VGND.t1443 Vbias.t133 XA.XIR[9].XIC[4].icell.SM VGND.t1442 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1383 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t659 VPWR.t658 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1384 VGND.t1445 Vbias.t134 XA.XIR[14].XIC[10].icell.SM VGND.t1444 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1385 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t373 VGND.t372 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1386 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1387 VGND.t1280 data[2].t1 XThC.XTB7.B VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1388 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t752 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t1847 XThR.XTBN.Y.t61 XThR.Tn[2].t10 VGND.t582 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1390 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t2409 VGND.t2408 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1391 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t78 VGND.t766 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1392 a_n1049_5317# XThR.XTB7.Y VPWR.t141 VPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1393 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1394 VGND.t482 XThC.XTBN.Y.t60 XThC.Tn[4].t5 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1395 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t1913 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1396 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t115 VGND.t114 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1397 XA.XIR[2].XIC_15.icell.PDM VPWR.t1999 VGND.t250 VGND.t249 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t106 VGND.t1241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1399 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t149 VGND.t1624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1400 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1401 VGND.t1447 Vbias.t135 XA.XIR[15].XIC[0].icell.SM VGND.t1446 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1402 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t98 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 VGND.t1449 Vbias.t136 XA.XIR[14].XIC[1].icell.SM VGND.t1448 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 VGND.t1451 Vbias.t137 XA.XIR[10].XIC[12].icell.SM VGND.t1450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1405 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t221 VGND.t2335 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1406 XThR.Tn[3].t2 XThR.XTB4.Y VGND.t954 VGND.t701 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1407 VGND.t1453 Vbias.t138 XA.XIR[13].XIC[13].icell.SM VGND.t1452 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1408 VPWR.t1513 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1512 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1409 VGND.t2617 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t2616 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1410 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t1051 VPWR.t1050 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1411 VPWR.t71 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1412 VPWR.t839 XThC.XTB7.Y a_6243_9615# VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VPWR.t989 XThC.XTB6.Y XThC.Tn[13].t10 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1414 VPWR.t1260 VPWR.t1258 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1259 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1415 VGND.t2336 data[1].t3 XThC.XTB5.A VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1416 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t1607 VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1417 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t1798 VPWR.t1797 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1418 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t1271 VGND.t1270 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1419 Vbias.t11 bias[2].t0 VPWR.t1711 VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.1955 pd=1.31 as=0.2465 ps=2.28 w=0.85 l=0.5
X1420 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t96 VPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1421 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1255 VPWR.t1257 VPWR.t1256 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 VGND.t1455 Vbias.t139 XA.XIR[3].XIC[3].icell.SM VGND.t1454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1423 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t203 VGND.t2027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1424 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t244 VGND.t2562 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1425 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t174 VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1426 VPWR.t699 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t698 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1427 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t375 VGND.t374 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1428 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1429 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t230 VGND.t2411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1430 VGND.t484 XThC.XTBN.Y.t61 XThC.Tn[7].t2 VGND.t483 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1431 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1570 VGND.t1569 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1432 VPWR.t925 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t924 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1433 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1434 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t131 VGND.t1510 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1435 XA.XIR[15].XIC[12].icell.PDM VPWR.t2000 XA.XIR[15].XIC[12].icell.Ien VGND.t251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1436 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t1303 VGND.t1302 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1437 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t448 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XThR.Tn[12].t8 XThR.XTB5.Y VPWR.t854 VPWR.t549 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1439 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1440 a_10915_9569# XThC.XTBN.Y.t62 VGND.t486 VGND.t485 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1441 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t181 VGND.t1824 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1442 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1616 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1443 XThR.Tn[6].t9 XThR.XTBN.Y.t62 VGND.t1849 VGND.t1848 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1444 VPWR.t1053 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t1052 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1445 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t2481 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1446 XThC.Tn[9].t5 XThC.XTB2.Y VPWR.t382 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1447 VGND.t2091 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t2090 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1448 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t6 VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1449 VGND.t1657 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1450 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t1896 VGND.t1895 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t754 VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1452 VGND.t1457 Vbias.t140 XA.XIR[5].XIC[11].icell.SM VGND.t1456 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1453 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t813 VPWR.t812 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1454 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t43 VGND.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1455 VGND.t253 VPWR.t2001 XA.XIR[1].XIC_15.icell.PDM VGND.t252 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1456 VPWR.t775 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1457 VPWR.t701 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t700 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1458 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1459 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1252 VPWR.t1254 VPWR.t1253 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1460 VPWR.t1583 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t1582 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1461 XA.XIR[15].XIC[10].icell.PDM VPWR.t2002 XA.XIR[15].XIC[10].icell.Ien VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1462 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t86 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1463 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t315 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 VGND.t1234 XThR.XTB7.B a_n1335_8331# VGND.t1233 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1465 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t1305 VGND.t1304 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1466 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t1934 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1467 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t1273 VGND.t1272 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1468 VGND.t1836 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t1835 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 VPWR.t232 XThC.XTBN.Y.t63 XThC.Tn[9].t9 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1471 XA.XIR[15].XIC_15.icell.PUM VPWR.t1250 XA.XIR[15].XIC_15.icell.Ien VPWR.t1251 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1472 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t189 VGND.t1908 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1473 a_10051_9569# XThC.XTBN.Y.t64 VGND.t488 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1474 VGND.t2225 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t2224 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1475 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t134 VGND.t1514 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1476 VPWR.t982 XThR.XTBN.Y.t63 XThR.Tn[7].t5 VPWR.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1477 VPWR.t1055 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t1054 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1478 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1479 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1248 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1249 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1480 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t166 VGND.t1709 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1481 VPWR.t266 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t265 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1482 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t67 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1483 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1484 XThC.Tn[11].t8 XThC.XTB4.Y.t8 VPWR.t1831 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1485 VGND.t1850 XThR.XTBN.Y.t64 XThR.Tn[1].t6 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1486 XThR.Tn[1].t9 XThR.XTBN.Y.t65 a_n1049_7787# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1487 a_7651_9569# XThC.XTBN.Y.t65 VGND.t490 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1488 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1650 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1489 VGND.t1459 Vbias.t141 XA.XIR[11].XIC[5].icell.SM VGND.t1458 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1490 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t176 VPWR.t175 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1491 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1651 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1492 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t1912 VPWR.t1911 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1493 VGND.t1461 Vbias.t142 XA.XIR[5].XIC[9].icell.SM VGND.t1460 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1494 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2003 VGND.t256 VGND.t255 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1495 VPWR.t1057 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t1056 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1496 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t1986 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1497 VPWR.t59 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1498 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t1306 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1499 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t376 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XThR.Tn[6].t1 XThR.XTB7.Y VGND.t229 VGND.t228 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1501 a_n1049_5611# XThR.XTB6.Y VPWR.t647 VPWR.t140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 XThR.Tn[9].t4 XThR.XTB2.Y VPWR.t43 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 VPWR.t1247 VPWR.t1245 XA.XIR[11].XIC_15.icell.PUM VPWR.t1246 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1504 VGND.t1463 Vbias.t143 XA.XIR[0].XIC[7].icell.SM VGND.t1462 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1505 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t1935 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1506 Vbias.t9 bias[0].t0 VPWR.t882 VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.12325 pd=1.14 as=0.1275 ps=1.15 w=0.85 l=2
X1507 XThC.Tn[4].t4 XThC.XTBN.Y.t66 VGND.t1769 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1508 VGND.t631 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t630 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t756 VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1510 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t2321 VGND.t2320 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 VPWR.t983 XThR.XTBN.Y.t66 XThR.Tn[13].t1 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t560 VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1511 VPWR.t1510 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VGND.t1074 VGND.t1072 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t1073 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1516 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t1937 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t161 VGND.t1681 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1518 VPWR.t703 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t258 VPWR.t2004 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t257 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t1585 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t1584 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t268 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t267 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1764 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 VGND.t1641 XThR.XTB1.Y.t11 XThR.Tn[0].t11 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t164 VGND.t1707 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1526 XThR.Tn[5].t5 XThR.XTBN.Y.t67 VGND.t1851 VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t627 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t1069 VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t1066 VGND.t1068 VGND.t1067 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t1232 XThR.XTB7.B XThR.XTB6.Y VGND.t1230 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t973 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1532 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t87 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 VGND.t1770 XThC.XTBN.Y.t67 XThC.Tn[0].t5 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 VGND.t2659 Vbias.t144 XA.XIR[8].XIC[5].icell.SM VGND.t2658 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1536 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t1817 VPWR.t1816 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 VGND.t2661 Vbias.t145 XA.XIR[12].XIC[13].icell.SM VGND.t2660 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1538 VGND.t1672 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t1671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t260 VPWR.t2005 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t2619 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t2618 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t1771 XThC.XTBN.Y.t68 XThC.Tn[3].t3 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t2663 Vbias.t146 XA.XIR[15].XIC[14].icell.SM VGND.t2662 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1543 VGND.t2189 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t2188 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VGND.t135 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1545 VPWR.t270 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t269 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1546 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2006 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t261 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t75 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1549 XThC.Tn[7].t1 XThC.XTBN.Y.t69 VGND.t1773 VGND.t1772 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1550 VPWR.t930 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1551 VGND.t2665 Vbias.t147 XA.XIR[11].XIC[0].icell.SM VGND.t2664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t178 VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t73 VPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1554 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1242 VPWR.t1244 VPWR.t1243 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1555 VGND.t2667 Vbias.t148 XA.XIR[2].XIC_15.icell.SM VGND.t2666 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1556 VGND.t2669 Vbias.t149 XA.XIR[6].XIC[12].icell.SM VGND.t2668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1557 VGND.t923 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t922 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 VGND.t119 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VPWR.t41 XThR.XTB2.Y a_n1049_7787# VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1560 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t1819 VPWR.t1818 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1561 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t562 VGND.t561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1562 VGND.t2671 Vbias.t150 XA.XIR[5].XIC[4].icell.SM VGND.t2670 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1563 VGND.t2673 Vbias.t151 XA.XIR[9].XIC[13].icell.SM VGND.t2672 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1564 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t141 VGND.t1579 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1565 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t661 VPWR.t660 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 VGND.t1775 XThC.XTBN.Y.t71 a_10915_9569# VGND.t1774 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VPWR.t610 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t609 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 VPWR.t815 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t814 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1569 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t1509 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2007 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1572 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t231 VGND.t2412 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t1613 VPWR.t1612 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1574 XThC.Tn[11].t9 XThC.XTB4.Y.t9 a_8963_9569# VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t2472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1576 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2008 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1577 VPWR.t75 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1578 VGND.t2482 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t2675 Vbias.t152 XA.XIR[0].XIC[2].icell.SM VGND.t2674 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1580 XThR.Tn[14].t11 XThR.XTBN.Y.t68 VPWR.t400 VPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t628 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1240 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1241 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 a_7875_9569# XThC.XTBN.Y.t72 VGND.t1776 VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 VPWR.t646 XThR.XTB6.Y XThR.Tn[13].t7 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VGND.t2093 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t2092 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1586 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t1661 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t208 VGND.t2292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1589 XA.XIR[0].XIC[3].icell.PDM VGND.t1063 VGND.t1065 VGND.t1064 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1590 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1591 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1592 XThC.Tn[11].t10 XThC.XTB4.Y.t11 a_8963_9569# VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1593 VGND.t2677 Vbias.t153 XA.XIR[8].XIC[0].icell.SM VGND.t2676 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1594 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1595 VGND.t2679 Vbias.t154 XA.XIR[3].XIC[12].icell.SM VGND.t2678 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1596 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t77 VPWR.t76 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1597 VGND.t1062 VGND.t1060 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t1061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1598 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1238 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1239 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1599 XThC.Tn[0].t8 XThC.XTB1.Y.t12 VGND.t1298 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t102 VGND.t980 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1601 VGND.t1777 XThC.XTBN.Y.t73 a_10051_9569# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VGND.t1202 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t1201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1603 VPWR.t817 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t816 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 VGND.t2621 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t2620 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 XThR.XTB1.Y.t2 XThR.XTB5.A VPWR.t958 VPWR.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 VPWR.t608 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t607 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1607 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1608 XThR.Tn[13].t8 XThR.XTB6.Y a_n997_1579# VGND.t1253 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t2323 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1610 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t852 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2010 VGND.t266 VGND.t265 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1612 VGND.t1634 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1613 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t538 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1614 VGND.t1778 XThC.XTBN.Y.t74 a_7651_9569# VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1615 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t1587 VPWR.t1586 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t109 VGND.t1244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1617 XThC.XTBN.Y.t0 XThC.XTBN.A VGND.t762 VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t819 VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1619 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1235 VPWR.t1237 VPWR.t1236 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1620 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t1502 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1621 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t138 VGND.t1576 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1622 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t1503 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1852 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1624 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y VGND.t836 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t2473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t1274 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[0].XIC[7].icell.PDM VGND.t1057 VGND.t1059 VGND.t1058 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_n1049_5317# XThR.XTBN.Y.t69 XThR.Tn[6].t6 VPWR.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1630 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2011 VGND.t268 VGND.t267 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t664 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1632 VPWR.t932 XThC.XTBN.Y.t75 XThC.Tn[7].t4 VPWR.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1633 VPWR.t1507 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t2083 VGND.t2082 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1635 XA.XIR[15].XIC[8].icell.Ien VPWR.t1232 VPWR.t1234 VPWR.t1233 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 VPWR.t79 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t78 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1637 VGND.t745 XThR.XTBN.Y.t70 a_n997_1803# VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 VPWR.t408 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 XThR.Tn[3].t5 XThR.XTBN.Y.t71 VGND.t746 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1640 VGND.t2095 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t2094 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1641 VPWR.t663 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t662 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1642 VPWR.t1832 XThC.XTB4.Y.t12 XThC.Tn[11].t11 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 VGND.t2681 Vbias.t155 XA.XIR[2].XIC[8].icell.SM VGND.t2680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1646 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t1939 VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t777 VPWR.t776 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1648 VGND.t1622 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t1621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t2085 VGND.t2084 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t891 VGND.t890 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t1589 VPWR.t1588 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t116 VGND.t1301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 VGND.t270 VPWR.t2012 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1654 XThC.Tn[0].t4 XThC.XTBN.Y.t76 VGND.t1779 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t178 VGND.t1821 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 VPWR.t821 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1657 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t68 VGND.t699 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 XThC.Tn[3].t2 XThC.XTBN.Y.t77 VGND.t1780 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 VGND.t925 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t924 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 VGND.t121 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1663 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t88 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t863 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t89 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 XA.XIR[8].XIC_15.icell.PUM VPWR.t1230 XA.XIR[8].XIC_15.icell.Ien VPWR.t1231 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t1031 VPWR.t1030 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 VGND.t1784 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t182 VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1670 VPWR.t1229 VPWR.t1227 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1228 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1671 VGND.t2633 Vbias.t156 XA.XIR[10].XIC[6].icell.SM VGND.t2632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 VGND.t2191 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t2190 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1673 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t1808 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1674 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t1059 VPWR.t1058 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VPWR.t410 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1676 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 VGND.t2635 Vbias.t157 XA.XIR[1].XIC_15.icell.SM VGND.t2634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t99 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1679 XThC.XTB1.Y.t1 XThC.XTB5.A a_3299_10575# VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1680 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t823 VPWR.t822 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1681 VPWR.t1505 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1504 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1682 VGND.t705 XThR.XTB3.Y XThR.Tn[2].t6 VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 XA.XIR[15].XIC[3].icell.Ien VPWR.t1224 VPWR.t1226 VPWR.t1225 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1684 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t2087 VGND.t2086 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1685 VGND.t2637 Vbias.t158 XA.XIR[11].XIC[14].icell.SM VGND.t2636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t180 VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1687 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t1662 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1688 VPWR.t81 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t80 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t412 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t411 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1691 VPWR.t705 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t1571 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1693 VPWR.t1591 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t1590 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 VPWR.t121 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t120 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1695 VGND.t1782 XThC.XTBN.Y.t78 XThC.Tn[6].t2 VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VGND.t2639 Vbias.t159 XA.XIR[2].XIC[3].icell.SM VGND.t2638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1697 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t148 VGND.t1623 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 XThC.Tn[10].t4 XThC.XTB3.Y.t11 VPWR.t665 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t893 VGND.t892 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1700 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t72 VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1701 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t1593 VPWR.t1592 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 VGND.t1056 VGND.t1054 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t1055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 VGND.t2641 Vbias.t160 XA.XIR[14].XIC[7].icell.SM VGND.t2640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1704 VGND.t2643 Vbias.t161 XA.XIR[10].XIC[10].icell.SM VGND.t2642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1705 XThC.Tn[14].t10 XThC.XTB7.Y VPWR.t838 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t758 VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t272 VPWR.t2013 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t1299 XThC.XTB1.Y.t13 XThC.Tn[0].t9 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 VGND.t1636 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t1635 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t736 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t1915 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 VGND.t2645 Vbias.t162 XA.XIR[10].XIC[1].icell.SM VGND.t2644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1715 XThR.Tn[8].t5 XThR.XTBN.Y.t72 VPWR.t403 VPWR.t402 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t136 VGND.t1525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 VGND.t2647 Vbias.t163 XA.XIR[5].XIC[13].icell.SM VGND.t2646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1718 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t163 VGND.t1683 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1719 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t2475 VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t2477 VGND.t2476 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t1427 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t1426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 VGND.t2623 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t2622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t1061 VPWR.t1060 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1724 VGND.t2625 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t2624 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1725 VGND.t2649 Vbias.t164 XA.XIR[8].XIC[14].icell.SM VGND.t2648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t515 VPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t137 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2014 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y.t73 XThR.Tn[5].t1 VPWR.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t825 VPWR.t824 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t2072 VGND.t2071 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t30 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 VGND.t2651 Vbias.t165 XA.XIR[4].XIC[11].icell.SM VGND.t2650 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1734 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t82 VGND.t780 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1735 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t70 VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1736 XThR.XTBN.A data[7].t1 VGND.t1666 VGND.t1665 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1737 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1738 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1739 XThC.Tn[14].t9 XThC.XTB7.Y VPWR.t837 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1740 VPWR.t970 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t2088 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t316 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t606 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t605 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2015 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t274 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t873 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t872 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 XThC.XTB2.Y XThC.XTB7.B VPWR.t558 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t1617 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1749 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t205 VGND.t2029 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t789 VPWR.t788 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XThR.Tn[5].t4 XThR.XTBN.Y.t74 VGND.t747 VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VGND.t2227 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t2226 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1753 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t2326 VGND.t2325 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 VGND.t2653 Vbias.t166 XA.XIR[14].XIC[2].icell.SM VGND.t2652 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1755 VGND.t2097 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t2096 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t9 XThR.XTBN.Y.t75 VPWR.t404 VPWR.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t517 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t2099 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t2098 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# XThC.XTB6.Y VPWR.t988 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t2655 Vbias.t167 XA.XIR[1].XIC[8].icell.SM VGND.t2654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t2040 Vbias.t168 XA.XIR[4].XIC[9].icell.SM VGND.t2039 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t214 VGND.t2314 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1763 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t2328 VGND.t2327 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1764 VPWR.t780 XThC.XTB3.Y.t12 XThC.Tn[10].t5 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1765 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t1826 VGND.t1825 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1766 VGND.t1053 VGND.t1051 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t1052 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1767 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t56 VGND.t491 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t249 VGND.t2585 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XThC.Tn[13].t0 XThC.XTBN.Y.t79 VPWR.t917 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1770 XA.XIR[13].XIC_15.icell.PDM VPWR.t2016 VGND.t276 VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1771 a_n997_3755# XThR.XTBN.Y.t76 VGND.t748 VGND.t686 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1772 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t39 VGND.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1773 VPWR.t406 XThR.XTBN.Y.t77 XThR.Tn[14].t10 VPWR.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t220 VGND.t2334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1775 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t317 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t184 VGND.t183 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t355 VGND.t354 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t864 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2017 VGND.t278 VGND.t277 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1781 VPWR.t972 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t971 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1782 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t894 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1783 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t791 VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1784 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t171 VGND.t1804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1785 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t31 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1786 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t158 VGND.t1664 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1787 XThR.Tn[7].t0 XThR.XTBN.Y.t78 VGND.t750 VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t46 VGND.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1789 VPWR.t1223 VPWR.t1221 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1790 VGND.t2229 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t2228 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1791 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t1713 VPWR.t1712 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1792 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t933 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 VGND.t280 VPWR.t2018 XA.XIR[15].XIC_15.icell.PDM VGND.t279 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1794 XThC.XTB4.Y.t0 XThC.XTB7.B VGND.t962 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1795 VPWR.t645 XThR.XTB6.Y XThR.Tn[13].t6 VPWR.t142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t376 XThR.XTB3.Y a_n1049_7493# VPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1798 VPWR.t1615 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1614 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1799 VGND.t2042 Vbias.t169 XA.XIR[7].XIC[5].icell.SM VGND.t2041 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t85 VPWR.t84 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t414 VPWR.t413 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1802 VPWR.t641 data[4].t3 XThR.XTB7.A VPWR.t640 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1803 VGND.t1674 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t1673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 VGND.t2044 Vbias.t170 XA.XIR[6].XIC[6].icell.SM VGND.t2043 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VGND.t282 VPWR.t2019 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t281 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2020 VGND.t284 VGND.t283 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t2330 VGND.t2329 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 XThC.Tn[6].t1 XThC.XTBN.Y.t80 VGND.t1715 VGND.t1714 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1809 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t1828 VGND.t1827 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1810 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t272 VPWR.t271 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t123 VPWR.t122 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t604 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 VPWR.t827 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t826 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1814 XThR.Tn[5].t9 XThR.XTB6.Y VGND.t1252 VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1815 VPWR.t519 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1816 VPWR.t679 XThC.XTB5.Y a_5155_9615# VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 VPWR.t1220 VPWR.t1218 XA.XIR[3].XIC_15.icell.PUM VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1818 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t2483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1819 VPWR.t1217 VPWR.t1215 XA.XIR[7].XIC_15.icell.PUM VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1820 VGND.t2046 Vbias.t171 XA.XIR[1].XIC[3].icell.SM VGND.t2045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t684 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t10 XThR.XTB5.Y VGND.t1627 VGND.t1255 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1461 VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t5 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 VGND.t2048 Vbias.t172 XA.XIR[4].XIC[4].icell.SM VGND.t2047 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1826 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t760 VGND.t759 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 VGND.t286 VPWR.t2021 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1828 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t151 VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1829 VGND.t1716 XThC.XTBN.Y.t82 XThC.Tn[2].t4 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t288 VPWR.t2022 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t118 VGND.t1308 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1832 VPWR.t697 XThC.XTB1.Y.t14 XThC.Tn[8].t9 VPWR.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VGND.t1289 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t1288 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# XThC.XTBN.Y.t83 VGND.t1718 VGND.t1717 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t1715 VPWR.t1714 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t934 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t975 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1839 VPWR.t1605 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1604 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1840 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t793 VPWR.t792 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1841 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t865 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1842 VGND.t2050 Vbias.t173 XA.XIR[6].XIC[10].icell.SM VGND.t2049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t1878 VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1844 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t1987 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1845 VGND.t2052 Vbias.t174 XA.XIR[3].XIC[6].icell.SM VGND.t2051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 VGND.t1676 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t1675 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t1786 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 VGND.t2193 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t2192 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t274 VPWR.t273 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1850 VGND.t1838 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1837 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t1416 VGND.t1415 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1852 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t1829 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1853 XThR.Tn[3].t4 XThR.XTBN.Y.t79 VGND.t751 VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t101 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1855 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t1834 VPWR.t1833 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 VGND.t2054 Vbias.t175 XA.XIR[7].XIC[0].icell.SM VGND.t2053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 VGND.t2056 Vbias.t176 XA.XIR[2].XIC[12].icell.SM VGND.t2055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1858 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t1880 VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 VGND.t2058 Vbias.t177 XA.XIR[6].XIC[1].icell.SM VGND.t2057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1213 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1214 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t5 VGND.t1592 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t276 VPWR.t275 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1863 a_4387_10575# XThC.XTB7.B VGND.t961 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t158 VPWR.t157 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1865 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t224 VGND.t2382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t125 VPWR.t124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t602 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t729 VPWR.t728 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t463 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t76 VGND.t723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1871 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t2484 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2023 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t289 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t2554 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t1830 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1876 a_10051_9569# XThC.XTBN.Y.t84 VGND.t1719 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t2076 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1878 XThC.XTB1.Y.t0 XThC.XTB7.B VPWR.t556 VPWR.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1879 a_n1049_6699# XThR.XTBN.Y.t80 XThR.Tn[3].t9 VPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1880 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t37 VGND.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t49 VGND.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1882 VGND.t2060 Vbias.t178 XA.XIR[3].XIC[10].icell.SM VGND.t2059 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1210 VPWR.t1212 VPWR.t1211 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t2503 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1885 a_n1049_8581# XThR.XTBN.Y.t81 XThR.Tn[0].t4 VPWR.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_7651_9569# XThC.XTBN.Y.t85 VGND.t1720 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1887 VGND.t1050 VGND.t1048 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t1049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 VGND.t633 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t632 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1889 VPWR.t1572 XThC.XTB7.A a_6243_10571# VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1890 VPWR.t1209 VPWR.t1207 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1208 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1891 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t1518 VGND.t1517 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1892 VPWR.t1607 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1606 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1893 XThC.Tn[10].t6 XThC.XTB3.Y.t13 a_8739_9569# VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VGND.t2062 Vbias.t179 XA.XIR[3].XIC[1].icell.SM VGND.t2061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t199 VGND.t1954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1896 VGND.t1429 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t1428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 VGND.t680 XThR.XTBN.Y.t82 XThR.Tn[2].t3 VGND.t679 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1898 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t465 VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t467 VGND.t466 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t48 VGND.t351 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1901 XThR.XTB5.A data[5].t3 VGND.t977 VGND.t976 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t33 VGND.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1903 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1205 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1206 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t1418 VGND.t1417 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1905 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t895 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1907 XThR.Tn[12].t1 XThR.XTBN.Y.t83 VPWR.t347 VPWR.t346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1908 VGND.t291 VPWR.t2024 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t290 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 Vbias.t7 Vbias.t6 VGND.t1166 VGND.t1164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.754 pd=5.78 as=0.754 ps=5.78 w=2.6 l=0.5
X1910 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t2486 VGND.t2485 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1911 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t32 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1912 XThR.Tn[12].t5 XThR.XTB5.Y a_n997_1803# VGND.t1254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1913 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t233 VGND.t2414 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1914 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t33 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1915 XThR.Tn[3].t1 XThR.XTB4.Y VGND.t953 VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1916 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t227 VGND.t2394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1917 VGND.t681 XThR.XTBN.Y.t84 a_n997_2667# VGND.t588 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1918 XA.XIR[9].XIC_15.icell.PDM VPWR.t2025 VGND.t293 VGND.t292 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1919 Vbias.t3 bias[2].t1 VPWR.t799 VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.1955 pd=1.31 as=0.2465 ps=2.28 w=0.85 l=0.5
X1920 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t2555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1921 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t119 VGND.t1479 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1922 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t349 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1923 VGND.t2531 Vbias.t180 XA.XIR[13].XIC_15.icell.SM VGND.t2530 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1924 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1202 VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1925 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t318 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1926 VGND.t123 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1927 VGND.t35 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t34 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1928 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t612 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1929 Vbias.t0 bias[0].t1 VPWR.t223 VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.12325 pd=1.14 as=0.1275 ps=1.15 w=0.85 l=2
X1930 a_5155_9615# XThC.XTB5.Y VPWR.t678 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1931 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t356 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1932 VPWR.t677 XThC.XTB5.Y XThC.Tn[12].t4 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1933 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t1419 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1934 VPWR.t1717 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t1716 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1935 XA.XIR[7].XIC_15.icell.PUM VPWR.t1200 XA.XIR[7].XIC_15.icell.Ien VPWR.t1201 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1936 VPWR.t1632 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t1631 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1937 VPWR.t1199 VPWR.t1197 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1198 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1938 VGND.t2231 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t2230 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1939 XThC.Tn[5].t4 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t150 VGND.t1637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1941 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t1263 VGND.t1262 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1942 VGND.t1284 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1943 a_n1049_6405# XThR.XTBN.Y.t85 XThR.Tn[4].t1 VPWR.t348 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1944 VPWR.t962 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t961 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1945 VPWR.t795 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t794 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1946 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t184 VGND.t1843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1947 XThC.Tn[2].t3 XThC.XTBN.Y.t87 VGND.t1721 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1948 VPWR.t160 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t159 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1949 XA.XIR[15].XIC[14].icell.PDM VPWR.t2026 XA.XIR[15].XIC[14].icell.Ien VGND.t294 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1950 XA.XIR[15].XIC[8].icell.PDM VPWR.t2027 XA.XIR[15].XIC[8].icell.Ien VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1951 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t9 VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1952 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t1520 VGND.t1519 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1953 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t1265 VGND.t1264 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1954 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1955 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t129 VGND.t1508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1956 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1957 VPWR.t632 XThR.XTB7.B XThR.XTB2.Y VPWR.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1958 XThC.Tn[8].t4 XThC.XTB1.Y.t15 a_7651_9569# VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1959 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t469 VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t1291 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t1290 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1961 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t241 VGND.t2559 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1962 XA.XIR[6].XIC_15.icell.PDM VPWR.t2028 VGND.t297 VGND.t296 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1963 VGND.t1575 XThC.XTB5.A XThC.XTB5.Y VGND.t481 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1964 VGND.t1047 VGND.t1045 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t1046 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1965 VGND.t227 XThR.XTB7.Y XThR.Tn[6].t0 VGND.t226 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1966 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1967 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t90 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t102 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1969 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t2488 VGND.t2487 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1811 VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 VPWR.t1719 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t1718 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1972 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t103 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1973 XA.XIR[4].XIC_15.icell.PUM VPWR.t1195 XA.XIR[4].XIC_15.icell.Ien VPWR.t1196 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t359 VGND.t358 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1975 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t8 VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1976 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2029 VGND.t299 VGND.t298 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1977 XA.XIR[15].XIC[9].icell.Ien VPWR.t1192 VPWR.t1194 VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1978 VGND.t1840 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1839 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 XThR.Tn[9].t8 XThR.XTBN.Y.t86 VPWR.t349 VPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1980 VGND.t1722 XThC.XTBN.Y.t89 a_9827_9569# VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1981 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t935 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t964 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t963 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t145 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1984 VGND.t301 VPWR.t2030 XA.XIR[8].XIC_15.icell.PDM VGND.t300 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1985 VPWR.t127 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t126 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1986 VGND.t2533 Vbias.t181 XA.XIR[1].XIC[12].icell.SM VGND.t2532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1987 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t1721 VPWR.t1720 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1988 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1189 VPWR.t1191 VPWR.t1190 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1989 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t1940 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1990 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1187 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1188 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1991 XThC.Tn[0].t10 XThC.XTB1.Y.t16 VGND.t1516 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1992 VGND.t2535 Vbias.t182 XA.XIR[0].XIC[5].icell.SM VGND.t2534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1993 VGND.t2537 Vbias.t183 XA.XIR[4].XIC[13].icell.SM VGND.t2536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1994 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t1941 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1995 VGND.t1678 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t1677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1996 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t4 VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1997 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t1267 VGND.t1266 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1998 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1503 VPWR.t1502 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1999 VGND.t2539 Vbias.t184 XA.XIR[7].XIC[14].icell.SM VGND.t2538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2000 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t1836 VPWR.t1835 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2001 VPWR.t966 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t471 VGND.t470 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2003 VGND.t139 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2004 VPWR.t797 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t1598 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2006 XThR.Tn[14].t9 XThR.XTBN.Y.t87 VPWR.t351 VPWR.t350 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2007 VPWR.t162 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t161 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2008 VPWR.t1186 VPWR.t1184 XA.XIR[0].XIC_15.icell.PUM VPWR.t1185 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2009 VPWR.t1634 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t1633 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2010 XA.XIR[15].XIC[3].icell.PDM VPWR.t2031 XA.XIR[15].XIC[3].icell.Ien VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 a_n997_3755# XThR.XTBN.Y.t88 VGND.t682 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2012 XThR.Tn[8].t0 XThR.XTB1.Y.t13 VPWR.t29 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2013 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2014 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t1684 VPWR.t1683 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2015 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1813 VGND.t1812 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2016 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t146 VGND.t1584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t2541 Vbias.t185 XA.XIR[10].XIC[7].icell.SM VGND.t2540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2018 a_n1049_7787# XThR.XTB2.Y VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2019 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t55 VGND.t418 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2020 VGND.t635 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t634 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2021 VPWR.t203 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t202 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2022 a_n1331_2891# data[5].t4 VGND.t870 VGND.t869 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2023 VGND.t2543 Vbias.t186 XA.XIR[13].XIC[8].icell.SM VGND.t2542 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2024 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t205 VPWR.t204 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2025 VPWR.t1183 VPWR.t1181 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1182 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2026 VGND.t875 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t874 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2027 VPWR.t1723 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t1722 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2028 XThR.XTB7.B data[6].t1 VGND.t1910 VGND.t1909 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2029 XThR.Tn[2].t4 XThR.XTBN.Y.t89 a_n1049_7493# VPWR.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2030 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t614 VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2031 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t616 VGND.t615 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1501 VPWR.t1500 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2033 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t153 VGND.t1640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2034 VGND.t2627 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t2626 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2035 VGND.t141 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2036 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 XA.XIR[15].XIC[7].icell.PDM VPWR.t2033 XA.XIR[15].XIC[7].icell.Ien VGND.t304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2038 VGND.t2545 Vbias.t187 XA.XIR[0].XIC[0].icell.SM VGND.t2544 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2039 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t429 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 VPWR.t919 XThC.XTBN.Y.t90 XThC.Tn[8].t2 VPWR.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2041 XThR.Tn[10].t5 XThR.XTB3.Y VPWR.t375 VPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2042 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t1268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2043 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XThR.Tn[4].t5 XThR.XTBN.Y.t90 VGND.t684 VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2045 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2046 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1179 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2047 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1499 VPWR.t1498 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2048 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t27 VGND.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2049 VGND.t1231 XThR.XTB7.B XThR.XTB5.Y VGND.t1230 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2050 VGND.t2547 Vbias.t188 XA.XIR[12].XIC_15.icell.SM VGND.t2546 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2051 VGND.t565 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t564 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t1420 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2053 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t1725 VPWR.t1724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2054 VGND.t37 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2055 VPWR.t1636 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t1635 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t496 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2057 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 VPWR.t207 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t206 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2059 VPWR.t302 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t301 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2060 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t2489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2061 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t112 VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2062 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t2331 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2063 VPWR.t1609 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1608 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2064 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t1 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2065 XThC.Tn[4].t8 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2066 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t1638 VPWR.t1637 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2067 VGND.t2549 Vbias.t189 XA.XIR[10].XIC[2].icell.SM VGND.t2548 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2068 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t202 VGND.t2016 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2069 VGND.t2551 Vbias.t190 XA.XIR[9].XIC_15.icell.SM VGND.t2550 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2070 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t173 VGND.t1815 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2071 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1176 VPWR.t1178 VPWR.t1177 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2072 VGND.t2101 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t2100 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2073 VGND.t2553 Vbias.t191 XA.XIR[13].XIC[3].icell.SM VGND.t2552 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2074 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t2282 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2075 VPWR.t731 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t730 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2076 VGND.t685 XThR.XTBN.Y.t91 a_n997_1579# VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2077 VPWR.t221 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2078 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2034 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2081 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t1618 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2082 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t618 VGND.t617 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2083 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t0 VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2084 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t59 VGND.t495 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t1 VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2086 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t737 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2087 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t200 VGND.t1959 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2088 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1174 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1175 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t237 VGND.t2434 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2090 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2091 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t2297 VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[0].XIC[5].icell.PDM VGND.t1042 VGND.t1044 VGND.t1043 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2093 VPWR.t304 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t303 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2094 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t1422 VGND.t1421 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t215 VGND.t2317 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2096 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t2078 VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2097 VGND.t147 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2098 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t1727 VPWR.t1726 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 XThR.XTBN.Y.t2 XThR.XTBN.A VPWR.t1874 VPWR.t1873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2100 VGND.t198 Vbias.t192 XA.XIR[15].XIC[11].icell.SM VGND.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2101 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t1640 VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2102 VPWR.t651 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t650 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2103 VGND.t567 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2104 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t2283 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2105 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t976 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2106 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2107 VGND.t39 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1171 VPWR.t1173 VPWR.t1172 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2109 VPWR.t746 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t745 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2110 XA.XIR[0].XIC_15.icell.PUM VPWR.t1169 XA.XIR[0].XIC_15.icell.Ien VPWR.t1170 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2111 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t985 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2112 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t1926 VPWR.t1925 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2113 VGND.t200 Vbias.t193 XA.XIR[2].XIC[6].icell.SM VGND.t199 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2114 VGND.t1788 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t1787 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2115 VGND.t2195 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t2194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t353 XThR.XTBN.Y.t92 XThR.Tn[11].t9 VPWR.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2117 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t1696 VPWR.t1695 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2118 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t620 VGND.t619 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2119 VPWR.t727 data[1].t4 XThC.XTB7.A VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2120 VPWR.t733 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t732 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2121 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1611 VPWR.t1610 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2122 a_8739_9569# XThC.XTBN.Y.t92 VGND.t1723 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 VGND.t2527 XThR.XTBN.A XThR.XTBN.Y.t0 VGND.t2526 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2124 XThC.Tn[6].t10 XThC.XTB7.Y VGND.t1591 VGND.t1590 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2125 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2126 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2127 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1653 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2128 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t2285 VGND.t2284 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1034 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2130 XThR.Tn[12].t4 XThR.XTB5.Y a_n997_1803# VGND.t1253 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2131 VGND.t308 VPWR.t2035 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t202 Vbias.t194 XA.XIR[12].XIC[8].icell.SM VGND.t201 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 VGND.t1293 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t1292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2134 VGND.t877 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t876 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2135 VGND.t204 Vbias.t195 XA.XIR[15].XIC[9].icell.SM VGND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2136 a_n997_3979# XThR.XTBN.Y.t93 VGND.t687 VGND.t686 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2137 XThC.XTB7.Y XThC.XTB7.B VGND.t960 VGND.t959 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2138 XA.XIR[0].XIC[0].icell.PDM VGND.t1039 VGND.t1041 VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2139 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1166 VPWR.t1168 VPWR.t1167 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2140 VGND.t206 Vbias.t196 XA.XIR[6].XIC[7].icell.SM VGND.t205 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2141 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t1928 VPWR.t1927 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2142 VGND.t208 Vbias.t197 XA.XIR[2].XIC[10].icell.SM VGND.t207 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2143 XThC.Tn[8].t1 XThC.XTBN.Y.t93 VPWR.t921 VPWR.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2144 VGND.t1790 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t1789 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2145 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t2080 VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 VGND.t2274 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t2273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2147 VGND.t210 Vbias.t198 XA.XIR[9].XIC[8].icell.SM VGND.t209 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2148 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t420 VPWR.t419 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2150 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2036 VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2151 VGND.t149 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2152 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t2556 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2153 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1595 VPWR.t1594 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2154 a_n1049_6699# XThR.XTB4.Y VPWR.t544 VPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2155 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t175 VGND.t1817 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2156 VPWR.t593 VGND.t2700 Vbias.t2 VPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.2465 pd=2.28 as=0.12325 ps=1.14 w=0.85 l=2
X2157 VPWR.t748 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2158 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t621 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2159 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t846 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2160 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t1930 VPWR.t1929 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2161 VGND.t212 Vbias.t199 XA.XIR[2].XIC[1].icell.SM VGND.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2162 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1164 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1165 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2163 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t168 VGND.t1725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2164 VGND.t1431 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t1430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2165 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1162 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t1698 VPWR.t1697 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2167 VGND.t214 Vbias.t200 XA.XIR[0].XIC[14].icell.SM VGND.t213 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2168 VGND.t216 Vbias.t201 XA.XIR[14].XIC[5].icell.SM VGND.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2169 VGND.t143 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2170 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t2490 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2171 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2037 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t2682 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t313 VPWR.t2038 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t312 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2175 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2176 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2177 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t1423 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2178 VGND.t1505 data[1].t5 XThC.XTB6.A VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2179 VPWR.t577 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t576 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2180 VPWR.t1158 VPWR.t1156 XA.XIR[14].XIC_15.icell.PUM VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2181 a_n997_2891# XThR.XTBN.Y.t94 VGND.t515 VGND.t514 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2182 VGND.t218 Vbias.t202 XA.XIR[12].XIC[3].icell.SM VGND.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2183 VGND.t220 Vbias.t203 XA.XIR[3].XIC[7].icell.SM VGND.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2184 VGND.t637 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t636 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2185 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t686 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2186 VPWR.t1882 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2187 VPWR.t1161 VPWR.t1159 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1160 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VGND.t1727 Vbias.t204 XA.XIR[15].XIC[4].icell.SM VGND.t1726 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2189 VGND.t1038 VGND.t1036 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t1037 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2190 VGND.t879 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t878 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2191 VPWR.t1155 VPWR.t1153 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1154 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2192 VPWR.t209 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t208 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2193 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2039 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t314 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2194 XThR.Tn[11].t5 XThR.XTB4.Y a_n997_2667# VGND.t709 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2195 VGND.t1729 Vbias.t205 XA.XIR[6].XIC[2].icell.SM VGND.t1728 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2196 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t2492 VGND.t2491 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 VPWR.t676 XThC.XTB5.Y a_5155_9615# VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2198 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t738 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2199 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t62 VGND.t592 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2200 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t862 VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2201 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t860 VGND.t859 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2202 VGND.t1731 Vbias.t206 XA.XIR[9].XIC[3].icell.SM VGND.t1730 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2203 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2204 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t2558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2205 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1597 VPWR.t1596 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2206 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t1425 VGND.t1424 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2207 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t623 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2208 VGND.t2197 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t2196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2210 VGND.t517 XThR.XTBN.Y.t95 XThR.Tn[0].t8 VGND.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2211 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t2494 VGND.t2493 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2212 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t1646 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2213 a_n1049_6405# XThR.XTB5.Y VPWR.t853 VPWR.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2214 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t117 VGND.t1307 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2215 XThR.Tn[8].t10 XThR.XTB1.Y.t14 VPWR.t1729 VPWR.t1728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2216 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t22 VGND.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t1917 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t1733 Vbias.t207 XA.XIR[14].XIC[0].icell.SM VGND.t1732 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t987 VGND.t986 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t60 VGND.t553 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2221 XA.XIR[5].XIC_15.icell.PDM VPWR.t2040 VGND.t316 VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 VGND.t1735 Vbias.t208 XA.XIR[5].XIC_15.icell.SM VGND.t1734 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2223 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t128 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2224 VGND.t2181 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t2180 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2225 VGND.t569 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t2683 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2227 VGND.t1737 Vbias.t209 XA.XIR[13].XIC[12].icell.SM VGND.t1736 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2228 XThR.Tn[1].t1 XThR.XTB2.Y VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 VGND.t571 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2230 VGND.t2183 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t2182 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2231 VPWR.t1884 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t1883 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 VGND.t1724 XThC.XTBN.Y.t94 a_8739_9569# VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t579 VPWR.t578 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2234 VGND.t1739 Vbias.t210 XA.XIR[1].XIC[6].icell.SM VGND.t1738 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2235 VPWR.t1152 VPWR.t1150 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 XThC.Tn[1].t2 XThC.XTB2.Y VGND.t719 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2237 VGND.t1589 XThC.XTB7.Y XThC.Tn[6].t9 VGND.t1588 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2238 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2041 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2239 VPWR.t306 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2240 VPWR.t1149 VPWR.t1147 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1148 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2241 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t1741 Vbias.t211 XA.XIR[3].XIC[2].icell.SM VGND.t1740 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2243 VGND.t1743 Vbias.t212 XA.XIR[11].XIC[11].icell.SM VGND.t1742 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2244 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t750 VPWR.t749 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XThR.Tn[2].t0 XThR.XTBN.Y.t96 a_n1049_7493# VPWR.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2246 VGND.t319 VPWR.t2042 XA.XIR[7].XIC_15.icell.PDM VGND.t318 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t193 VGND.t1923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2248 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t115 VPWR.t114 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2249 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t239 VGND.t2436 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2250 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t2287 VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2251 XThR.Tn[13].t0 XThR.XTBN.Y.t97 VPWR.t236 VPWR.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2252 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t2496 VGND.t2495 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t1686 VPWR.t1685 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2255 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t79 VGND.t773 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2256 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1036 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2257 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t858 VGND.t857 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2258 XThR.Tn[10].t4 XThR.XTB3.Y VPWR.t374 VPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2259 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t1619 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2260 XThR.Tn[4].t4 XThR.XTBN.Y.t98 VGND.t519 VGND.t518 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2261 VPWR.t211 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t210 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2262 VGND.t1035 VGND.t1033 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t1034 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 VGND.t1250 XThR.XTB6.Y XThR.Tn[5].t8 VGND.t1249 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2264 VGND.t1433 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t104 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2266 VGND.t1745 Vbias.t213 XA.XIR[1].XIC[10].icell.SM VGND.t1744 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2267 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t5 VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2268 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t989 VGND.t988 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2269 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t2 VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2270 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t174 VGND.t173 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2271 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2043 VGND.t321 VGND.t320 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2272 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t0 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2273 VGND.t151 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t1747 Vbias.t214 XA.XIR[11].XIC[9].icell.SM VGND.t1746 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t752 VPWR.t751 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t108 VGND.t1243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2277 VGND.t153 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t152 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 VGND.t1749 Vbias.t215 XA.XIR[8].XIC[11].icell.SM VGND.t1748 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2279 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t653 VPWR.t652 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2280 VPWR.t1688 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t1687 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t323 VPWR.t2044 XA.XIR[4].XIC_15.icell.PDM VGND.t322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1144 VPWR.t1146 VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2283 VGND.t1140 Vbias.t216 XA.XIR[1].XIC[1].icell.SM VGND.t1139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2284 VPWR.t1700 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t1699 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2285 VGND.t1792 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t1791 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2286 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t319 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t277 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2288 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t856 VGND.t855 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t990 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2290 VGND.t325 VPWR.t2045 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2291 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t94 VGND.t917 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2292 VGND.t1913 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1912 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2293 VPWR.t373 XThR.XTB3.Y a_n1049_7493# VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2294 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t187 VGND.t1906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2295 VPWR.t308 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t307 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2296 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2297 VPWR.t1599 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2298 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t245 VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2299 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t117 VPWR.t116 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2301 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t77 VGND.t765 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2302 VGND.t1142 Vbias.t217 XA.XIR[5].XIC[8].icell.SM VGND.t1141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2303 VGND.t594 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VPWR.t213 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2305 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2306 VPWR.t1143 VPWR.t1141 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1142 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2307 VGND.t596 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t595 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2308 VGND.t1144 Vbias.t218 XA.XIR[8].XIC[9].icell.SM VGND.t1143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2309 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t655 VPWR.t654 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2310 XThR.Tn[4].t9 XThR.XTB5.Y VGND.t1626 VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2311 VPWR.t238 XThR.XTBN.Y.t99 XThR.Tn[14].t8 VPWR.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2312 VPWR.t754 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t753 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2313 XThC.Tn[13].t9 XThC.XTB6.Y VPWR.t987 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2314 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2315 VGND.t1855 XThC.XTB6.Y XThC.Tn[5].t8 VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2316 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t177 VGND.t176 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2317 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t126 VGND.t1504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2318 VPWR.t240 XThR.XTBN.Y.t100 XThR.Tn[11].t8 VPWR.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2319 VGND.t1146 Vbias.t219 XA.XIR[11].XIC[4].icell.SM VGND.t1145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2320 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t756 VPWR.t755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2321 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t432 VGND.t431 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2322 VGND.t1032 VGND.t1030 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t1031 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2323 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t2074 VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2324 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t127 VGND.t1506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2325 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2326 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2327 XThC.Tn[9].t0 XThC.XTB2.Y a_7875_9569# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[4].XIC_15.icell.PDM VPWR.t2046 VGND.t327 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t936 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2330 VGND.t78 XThC.XTB6.A XThC.XTB6.Y VGND.t77 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2331 VGND.t718 XThC.XTB2.Y XThC.Tn[1].t1 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2332 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t129 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2333 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t107 VGND.t1242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t1148 Vbias.t220 XA.XIR[12].XIC[12].icell.SM VGND.t1147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1139 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1140 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2336 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2337 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t238 VGND.t2435 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2338 VGND.t1150 Vbias.t221 XA.XIR[15].XIC[13].icell.SM VGND.t1149 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2339 VGND.t1152 Vbias.t222 XA.XIR[14].XIC[14].icell.SM VGND.t1151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2340 VGND.t2629 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t2628 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2341 VGND.t1610 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t853 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2343 VPWR.t139 XThR.XTB7.Y a_n1049_5317# VPWR.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2344 VPWR.t310 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t309 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2345 VGND.t329 VPWR.t2047 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2346 VPWR.t986 XThC.XTB6.Y XThC.Tn[13].t8 VPWR.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2347 VPWR.t1601 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1600 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2348 a_n997_3979# XThR.XTBN.Y.t101 VGND.t521 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2349 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t427 VPWR.t426 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t119 VPWR.t118 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2351 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t312 VPWR.t311 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2352 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t196 VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1136 VPWR.t1138 VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2354 VGND.t1154 Vbias.t223 XA.XIR[5].XIC[3].icell.SM VGND.t1153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2355 VGND.t1156 Vbias.t224 XA.XIR[9].XIC[12].icell.SM VGND.t1155 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2356 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t34 VGND.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2357 VGND.t952 XThR.XTB4.Y XThR.Tn[3].t0 VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2358 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t240 VGND.t2480 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2359 a_7331_10587# data[0].t2 VPWR.t829 VPWR.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2360 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t8 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2361 VPWR.t1497 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2362 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t434 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2363 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t242 VGND.t2560 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2364 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1603 VPWR.t1602 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2365 VGND.t1158 Vbias.t225 XA.XIR[8].XIC[4].icell.SM VGND.t1157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2366 VGND.t1029 VGND.t1027 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t1028 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2367 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t107 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2368 VPWR.t1838 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t1837 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2370 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t92 VGND.t910 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2371 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2048 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2372 VPWR.t429 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t428 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2373 a_n1049_6699# XThR.XTBN.Y.t102 XThR.Tn[3].t8 VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2374 VGND.t1165 Vbias.t4 Vbias.t5 VGND.t1164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.754 pd=5.78 as=0.754 ps=5.78 w=2.6 l=0.5
X2375 XA.XIR[0].XIC[11].icell.PDM VGND.t1024 VGND.t1026 VGND.t1025 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2376 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t739 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2377 XA.XIR[1].XIC_15.icell.PDM VPWR.t2049 VGND.t332 VGND.t331 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t101 VGND.t979 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2379 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t104 VGND.t1163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2380 XThC.Tn[3].t4 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2381 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t1 VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2382 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1134 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1135 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XThC.XTB5.A data[0].t3 VGND.t1573 VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2384 VGND.t2103 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t2102 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2385 VPWR.t542 XThR.XTB4.Y XThR.Tn[11].t1 VPWR.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2386 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t795 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2387 XA.XIR[0].XIC[2].icell.PDM VGND.t1021 VGND.t1023 VGND.t1022 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2388 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t45 VGND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2389 VGND.t1295 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t1294 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2390 VGND.t523 XThR.XTBN.Y.t103 a_n997_715# VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2391 a_n997_2891# XThR.XTBN.Y.t104 VGND.t525 VGND.t524 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2392 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t162 VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2393 VGND.t1020 VGND.t1018 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t1019 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2394 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t431 VPWR.t430 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2395 VPWR.t735 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t734 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2396 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t1555 VPWR.t1554 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2397 VPWR.t1495 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1494 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2398 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1131 VPWR.t1133 VPWR.t1132 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2399 VPWR.t1840 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2400 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t991 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2401 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2402 XThR.Tn[11].t4 XThR.XTB4.Y a_n997_2667# VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2403 VPWR.t1130 VPWR.t1128 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1129 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2404 VGND.t2276 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t2275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2405 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2406 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t95 VGND.t926 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2407 VPWR.t381 XThC.XTB2.Y XThC.Tn[9].t4 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2408 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t1786 VPWR.t1785 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2409 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t11 VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2410 VGND.t334 VPWR.t2050 XA.XIR[0].XIC_15.icell.PDM VGND.t333 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2411 VGND.t1915 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1914 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2412 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t123 VGND.t1485 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2413 VPWR.t923 XThC.XTBN.Y.t100 XThC.Tn[8].t0 VPWR.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2414 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t74 VGND.t721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2415 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2416 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t2299 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2417 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t494 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2418 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2419 VPWR.t581 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t580 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2420 XA.XIR[0].XIC[6].icell.PDM VGND.t1015 VGND.t1017 VGND.t1016 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2421 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t2075 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2422 a_n1049_6405# XThR.XTBN.Y.t105 XThR.Tn[4].t0 VPWR.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2423 XA.XIR[15].XIC[7].icell.Ien VPWR.t1125 VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2424 XThR.Tn[7].t4 XThR.XTBN.Y.t106 VPWR.t243 VPWR.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2425 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2051 VGND.t1528 VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2426 VPWR.t433 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t432 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2427 VGND.t1014 VGND.t1012 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t1013 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VPWR.t422 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t421 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2429 XThC.Tn[9].t8 XThC.XTBN.Y.t101 VPWR.t1868 VPWR.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2430 XThR.Tn[1].t5 XThR.XTBN.Y.t107 VGND.t657 VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2431 VPWR.t1124 VPWR.t1122 XA.XIR[13].XIC_15.icell.PUM VPWR.t1123 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2432 VGND.t1160 Vbias.t226 XA.XIR[2].XIC[7].icell.SM VGND.t1159 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2433 VGND.t740 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2434 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2435 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t2470 VGND.t2469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2436 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t164 VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2437 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2052 VGND.t1530 VGND.t1529 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t1702 VPWR.t1701 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2439 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t1788 VPWR.t1787 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2440 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t1487 VGND.t1486 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2441 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t26 VGND.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2442 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t993 VGND.t992 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2443 VPWR.t1869 XThC.XTBN.Y.t102 XThC.Tn[11].t2 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2444 VPWR.t1493 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1492 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2445 VPWR.t644 XThR.XTB6.Y a_n1049_5611# VPWR.t138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2446 VGND.t1532 VPWR.t2053 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1531 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2447 a_n997_2891# XThR.XTB3.Y XThR.Tn[10].t1 VGND.t703 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2448 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t2684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2449 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t44 VGND.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2450 VPWR.t1842 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2451 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t1756 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1120 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1121 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2453 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t186 VGND.t1854 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2454 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t2686 VGND.t2685 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t540 VGND.t539 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2456 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t1672 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2457 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t2471 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2458 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t772 VGND.t771 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t278 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 VGND.t1162 Vbias.t227 XA.XIR[10].XIC[5].icell.SM VGND.t1161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2461 XA.XIR[15].XIC[11].icell.Ien VPWR.t1117 VPWR.t1119 VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2462 VGND.t1612 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1611 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2463 VGND.t1534 VPWR.t2054 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1533 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 XA.XIR[11].XIC_15.icell.PUM VPWR.t1115 XA.XIR[11].XIC_15.icell.Ien VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2466 VGND.t2109 Vbias.t228 XA.XIR[13].XIC[6].icell.SM VGND.t2108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2467 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t215 VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2468 VGND.t2199 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2469 VGND.t1536 VPWR.t2055 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1535 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 XThC.Tn[2].t7 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2471 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t2345 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2472 VPWR.t567 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2473 VPWR.t583 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t582 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2474 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t1806 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2475 VGND.t1229 XThR.XTB7.B XThR.XTB4.Y VGND.t1228 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2476 VPWR.t1114 VPWR.t1112 XA.XIR[10].XIC_15.icell.PUM VPWR.t1113 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2477 VGND.t2111 Vbias.t229 XA.XIR[4].XIC_15.icell.SM VGND.t2110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2478 XA.XIR[15].XIC[2].icell.Ien VPWR.t1109 VPWR.t1111 VPWR.t1110 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2479 VGND.t2113 Vbias.t230 XA.XIR[11].XIC[13].icell.SM VGND.t2112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2480 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t758 VPWR.t757 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2481 VGND.t240 XThR.XTB1.Y.t16 XThR.Tn[0].t0 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2482 VPWR.t255 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2483 VPWR.t435 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t434 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2484 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t1551 VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2485 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t245 VGND.t2563 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2486 VPWR.t569 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2487 XA.XIR[15].XIC[5].icell.PDM VPWR.t2056 XA.XIR[15].XIC[5].icell.Ien VGND.t1537 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2488 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t2395 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2489 VGND.t1297 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t1296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 VGND.t2115 Vbias.t231 XA.XIR[2].XIC[2].icell.SM VGND.t2114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2491 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1106 VPWR.t1108 VPWR.t1107 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t29 VGND.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2493 a_8739_9569# XThC.XTBN.Y.t104 VGND.t2520 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2494 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t983 VGND.t982 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2495 XThC.Tn[6].t8 XThC.XTB7.Y VGND.t1587 VGND.t1586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2496 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t1790 VPWR.t1789 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2497 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t2064 VGND.t2063 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2498 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t776 VGND.t775 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2499 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2500 VGND.t2117 Vbias.t232 XA.XIR[13].XIC[10].icell.SM VGND.t2116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2501 VGND.t2522 XThC.XTBN.Y.t105 XThC.Tn[7].t0 VGND.t2521 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t1870 VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2503 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t217 VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2504 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t2346 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2505 VGND.t2278 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t2277 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 XThC.Tn[12].t0 XThC.XTB5.Y a_9827_9569# VGND.t1283 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t195 VGND.t1950 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2508 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t544 VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t1620 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2510 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t1807 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2511 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t4 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2512 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t124 VGND.t1496 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2513 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t130 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 VGND.t2119 Vbias.t233 XA.XIR[10].XIC[0].icell.SM VGND.t2118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2515 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1104 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1105 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2516 VGND.t2121 Vbias.t234 XA.XIR[5].XIC[12].icell.SM VGND.t2120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2517 VGND.t2185 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t2184 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 VGND.t573 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2519 XThR.Tn[13].t5 XThR.XTB6.Y VPWR.t643 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2520 VGND.t2123 Vbias.t235 XA.XIR[13].XIC[1].icell.SM VGND.t2122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2521 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2522 VGND.t1435 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t1434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2523 VGND.t2125 Vbias.t236 XA.XIR[8].XIC[13].icell.SM VGND.t2124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2524 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t109 VPWR.t108 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2525 VGND.t2427 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2526 VPWR.t257 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2527 VGND.t192 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2528 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t292 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2529 VGND.t2523 XThC.XTBN.Y.t107 a_7875_9569# VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2530 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t435 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2531 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2057 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1538 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2532 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2533 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1491 VPWR.t1490 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t994 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2535 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t114 VGND.t1282 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2536 VGND.t2127 Vbias.t237 XA.XIR[7].XIC[11].icell.SM VGND.t2126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2537 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t1844 VPWR.t1843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2538 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t437 VPWR.t436 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2539 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t243 VGND.t2561 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2540 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t1557 VPWR.t1556 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2541 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t778 VGND.t777 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2542 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2543 VPWR.t600 VGND.t2701 XA.XIR[0].XIC[12].icell.PUM VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2544 XA.XIR[15].XIC[0].icell.PDM VPWR.t2058 XA.XIR[15].XIC[0].icell.Ien VGND.t1539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2545 a_8963_9569# XThC.XTBN.Y.t108 VGND.t2524 VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2546 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t2065 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2547 VGND.t742 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t546 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2550 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t1999 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t1103 VPWR.t1101 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1102 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t1621 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t2001 VGND.t2000 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2554 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2555 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2556 VPWR.t111 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t110 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2557 VGND.t2105 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t2104 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2558 XThC.Tn[11].t1 XThC.XTBN.Y.t109 VPWR.t1871 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2559 VPWR.t1576 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2560 VGND.t2129 Vbias.t238 XA.XIR[1].XIC[7].icell.SM VGND.t2128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2561 XThR.Tn[6].t5 XThR.XTBN.Y.t108 a_n1049_5317# VPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2562 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1655 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 VPWR.t1462 XThC.XTB4.Y.t16 XThC.Tn[11].t5 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2564 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2565 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t688 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 VGND.t2131 Vbias.t239 XA.XIR[4].XIC[8].icell.SM VGND.t2130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2567 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t996 VGND.t995 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2568 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t2003 VGND.t2002 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2569 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t2008 VGND.t2007 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2570 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2059 VGND.t1541 VGND.t1540 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2571 VGND.t155 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t154 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2572 VGND.t2233 Vbias.t240 XA.XIR[7].XIC[9].icell.SM VGND.t2232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2573 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t1846 VPWR.t1845 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2574 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1489 VPWR.t1488 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2575 XA.XIR[12].XIC_15.icell.PDM VPWR.t2060 VGND.t1543 VGND.t1542 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2576 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t105 VGND.t1240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2577 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t232 VGND.t2413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2578 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t176 VGND.t1819 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2579 VPWR.t598 VGND.t2702 XA.XIR[0].XIC[10].icell.PUM VPWR.t597 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2580 VPWR.t781 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2581 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t398 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2582 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2583 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t1673 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2584 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2066 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2585 VGND.t659 XThR.XTBN.Y.t109 a_n997_1803# VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2586 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t165 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2587 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t247 VPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2588 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t424 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2589 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2590 XA.XIR[10].XIC_15.icell.PUM VPWR.t1099 XA.XIR[10].XIC_15.icell.Ien VPWR.t1100 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 a_3773_9615# XThC.XTB2.Y VPWR.t380 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2592 VPWR.t1098 VPWR.t1096 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1097 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2593 VGND.t2235 Vbias.t241 XA.XIR[12].XIC[6].icell.SM VGND.t2234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2594 VGND.t1917 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1916 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2595 VGND.t2201 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2596 VPWR.t113 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t112 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2597 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2598 VPWR.t540 XThR.XTB4.Y XThR.Tn[11].t0 VPWR.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2599 a_n997_715# XThR.XTBN.Y.t110 VGND.t661 VGND.t660 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2600 VGND.t2237 Vbias.t242 XA.XIR[6].XIC[5].icell.SM VGND.t2236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2601 VPWR.t149 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2602 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1656 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2603 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t439 VPWR.t438 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2604 XThR.Tn[14].t5 XThR.XTB7.Y VPWR.t137 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2605 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t2005 VGND.t2004 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2606 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t1559 VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2607 VGND.t2239 Vbias.t243 XA.XIR[9].XIC[6].icell.SM VGND.t2238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2608 VGND.t2525 XThC.XTBN.Y.t110 XThC.Tn[3].t1 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2609 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t571 VPWR.t570 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2610 VGND.t598 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2611 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2061 VGND.t1545 VGND.t1544 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2612 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2613 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t834 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2614 VPWR.t1 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2615 XThC.Tn[1].t0 XThC.XTB2.Y VGND.t717 VGND.t79 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2616 VPWR.t1487 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1486 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2617 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t1710 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2618 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1811 VPWR.t1810 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2619 VPWR.t416 XThC.XTBN.A XThC.XTBN.Y.t2 VPWR.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2620 VPWR.t1578 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2621 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t2009 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2622 VPWR.t1768 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t1767 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2623 VGND.t2241 Vbias.t244 XA.XIR[1].XIC[2].icell.SM VGND.t2240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2624 VPWR.t1095 VPWR.t1093 XA.XIR[6].XIC_15.icell.PUM VPWR.t1094 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2625 VGND.t2243 Vbias.t245 XA.XIR[4].XIC[3].icell.SM VGND.t2242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2626 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t3 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2627 XThR.Tn[2].t5 XThR.XTB3.Y VGND.t702 VGND.t701 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2628 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t2011 VGND.t2010 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2629 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2630 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t41 VGND.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2631 VGND.t2245 Vbias.t246 XA.XIR[7].XIC[4].icell.SM VGND.t2244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2632 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t1770 VPWR.t1769 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2633 VGND.t1011 VGND.t1009 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t1010 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2634 VGND.t2247 Vbias.t247 XA.XIR[12].XIC[10].icell.SM VGND.t2246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2635 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2636 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t1 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t91 VGND.t909 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2638 a_3299_10575# XThC.XTB7.B VGND.t958 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2639 VGND.t1547 VPWR.t2062 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2640 VGND.t663 XThR.XTBN.Y.t111 XThR.Tn[6].t8 VGND.t662 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2641 VPWR.t596 VGND.t2703 XA.XIR[0].XIC[5].icell.PUM VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2642 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t1757 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2643 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t740 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2644 VPWR.t1813 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1812 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2645 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1090 VPWR.t1092 VPWR.t1091 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2647 VGND.t2249 Vbias.t248 XA.XIR[12].XIC[1].icell.SM VGND.t2248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2648 VGND.t2251 Vbias.t249 XA.XIR[3].XIC[5].icell.SM VGND.t2250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2649 VGND.t1437 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t1436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2650 VPWR.t594 VGND.t2704 Vbias.t1 VPWR.t592 sky130_fd_pr__pfet_01v8 ad=0.2465 pd=2.28 as=0.12325 ps=1.14 w=0.85 l=2
X2651 VGND.t1614 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1613 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VGND.t2253 Vbias.t250 XA.XIR[9].XIC[10].icell.SM VGND.t2252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2653 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t573 VPWR.t572 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2654 VGND.t2356 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t2355 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2655 VGND.t2255 Vbias.t251 XA.XIR[10].XIC[14].icell.SM VGND.t2254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2656 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2657 VGND.t2211 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t2210 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2658 VPWR.t1872 XThC.XTBN.Y.t111 XThC.Tn[10].t11 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2659 VGND.t194 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2063 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t1548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2661 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t1808 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2662 VGND.t2359 XThC.XTBN.Y.t112 a_8963_9569# VGND.t670 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t913 VPWR.t912 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 VGND.t81 Vbias.t252 XA.XIR[6].XIC[0].icell.SM VGND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2665 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t2385 VGND.t2384 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2666 VPWR.t830 XThC.XTB5.A a_5155_10571# VPWR.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2667 VPWR.t836 XThC.XTB7.Y XThC.Tn[14].t8 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 XThR.Tn[1].t4 XThR.XTBN.Y.t112 VGND.t665 VGND.t664 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2669 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t503 VPWR.t502 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2670 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t1561 VPWR.t1560 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2671 VGND.t83 Vbias.t253 XA.XIR[9].XIC[1].icell.SM VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2672 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t575 VPWR.t574 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2673 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t1792 VPWR.t1791 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2674 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t255 VGND.t2687 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2675 VPWR.t1571 XThC.XTB7.A XThC.XTB3.Y.t2 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2676 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1815 VPWR.t1814 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2677 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t1711 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2678 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t190 VGND.t1911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2679 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t142 VGND.t1580 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2680 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t2301 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2681 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t2012 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2682 XThR.Tn[8].t4 XThR.XTBN.Y.t113 VPWR.t334 VPWR.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2683 VPWR.t505 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2684 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2064 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t1549 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2685 XThR.Tn[5].t0 XThR.XTBN.Y.t114 a_n1049_5611# VPWR.t332 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2686 a_n997_2891# XThR.XTB3.Y XThR.Tn[10].t0 VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2687 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t984 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2688 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2689 VPWR.t1089 VPWR.t1087 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1088 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2690 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t247 VGND.t2565 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2691 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t38 VGND.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2692 a_n1049_7787# XThR.XTBN.Y.t115 XThR.Tn[1].t8 VPWR.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2693 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t9 VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2694 VPWR.t630 XThR.XTB7.B XThR.XTB3.Y VPWR.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2065 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t1550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2696 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t1622 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2697 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t782 VPWR.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2698 VGND.t85 Vbias.t254 XA.XIR[3].XIC[0].icell.SM VGND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2699 VPWR.t783 XThC.XTB3.Y.t16 XThC.Tn[10].t7 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2700 VPWR.t1758 XThC.XTBN.Y.t114 XThC.Tn[14].t1 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2701 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t507 VPWR.t506 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2702 VGND.t1008 VGND.t1006 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t1007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2703 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t849 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2704 XA.XIR[15].XIC_15.icell.PDM VPWR.t2066 VGND.t1552 VGND.t1551 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2705 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t13 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2706 VGND.t1439 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t1438 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2707 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t66 VGND.t697 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2708 VGND.t667 XThR.XTBN.Y.t116 XThR.Tn[0].t7 VGND.t666 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2709 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t19 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2710 VGND.t1511 XThC.XTB3.Y.t17 XThC.Tn[2].t11 VGND.t335 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2711 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t294 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2712 XThR.Tn[10].t8 XThR.XTBN.Y.t117 VPWR.t337 VPWR.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2713 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t2387 VGND.t2386 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2714 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2067 VGND.t1554 VGND.t1553 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2715 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t1581 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2716 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t54 VGND.t378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2717 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t1648 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2718 VGND.t87 Vbias.t255 XA.XIR[0].XIC[11].icell.SM VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2719 VPWR.t985 XThC.XTB6.Y a_5949_9615# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2720 XThR.Tn[1].t0 XThR.XTB2.Y VGND.t54 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2721 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t69 VGND.t712 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2722 VGND.t668 XThR.XTBN.Y.t118 a_n997_3755# VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2723 VPWR.t423 data[3].t1 XThC.XTBN.A VPWR.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2724 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t217 VGND.t2319 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2725 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t785 VPWR.t784 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2726 XThC.Tn[3].t0 XThC.XTBN.Y.t115 VGND.t2360 VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2727 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1485 VPWR.t1484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2728 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t213 VGND.t2304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2729 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t2688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2730 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t2391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2731 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t279 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2732 VPWR.t1704 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t1703 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2733 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t40 VGND.t221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2734 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1580 VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2735 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2736 VPWR.t509 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t508 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2737 VPWR.t249 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2738 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2068 VGND.t2067 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t1076 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XThR.Tn[13].t4 XThR.XTB6.Y VPWR.t642 VPWR.t146 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2741 VPWR.t1743 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1742 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2742 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t88 VGND.t841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2743 a_n1049_7493# XThR.XTB3.Y VPWR.t372 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2744 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2745 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t690 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2746 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2747 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2748 VGND.t1005 VGND.t1003 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t1004 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2749 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t797 VGND.t796 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2750 VGND.t89 Vbias.t256 XA.XIR[0].XIC[9].icell.SM VGND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2751 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t2070 VGND.t2069 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2752 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t248 VGND.t2584 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2753 VPWR.t787 XThC.XTB1.Y.t18 XThC.Tn[8].t8 VPWR.t786 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2754 VGND.t371 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2755 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t11 VGND.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2756 VGND.t1625 XThR.XTB5.Y XThR.Tn[4].t8 VGND.t1249 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2757 XThC.Tn[10].t9 XThC.XTBN.Y.t116 VPWR.t1759 VPWR.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2758 VGND.t2362 XThC.XTBN.Y.t117 XThC.Tn[6].t0 VGND.t2361 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2759 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t2392 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2760 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t1675 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 VPWR.t585 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t584 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2762 VPWR.t1706 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t1705 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2763 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t1676 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t425 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 XA.XIR[3].XIC_15.icell.PUM VPWR.t1085 XA.XIR[3].XIC_15.icell.Ien VPWR.t1086 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t2348 VGND.t2347 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VGND.t91 Vbias.t257 XA.XIR[5].XIC[6].icell.SM VGND.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2769 VGND.t2358 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t2357 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2770 VGND.t1556 VPWR.t2068 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2771 VGND.t2213 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t2212 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2772 VGND.t1807 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t1806 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2773 VGND.t2215 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t2214 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2774 VPWR.t1565 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2775 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2776 VPWR.t1463 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2777 VPWR.t1745 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1744 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2778 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t587 VPWR.t586 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2779 XA.XIR[15].XIC[11].icell.PDM VPWR.t2069 XA.XIR[15].XIC[11].icell.Ien VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2780 VGND.t1559 VPWR.t2070 XA.XIR[11].XIC_15.icell.PDM VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2781 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t131 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2782 VGND.t93 Vbias.t258 XA.XIR[4].XIC[12].icell.SM VGND.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 XThR.Tn[6].t4 XThR.XTBN.Y.t119 a_n1049_5317# VPWR.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2784 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1083 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1084 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2785 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t4 VGND.t1585 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2786 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1483 VPWR.t1482 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2787 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1867 VPWR.t1866 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2788 VGND.t95 Vbias.t259 XA.XIR[7].XIC[13].icell.SM VGND.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2789 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t1772 VPWR.t1771 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2790 VGND.t2364 XThC.XTBN.Y.t118 a_10915_9569# VGND.t2363 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2791 VPWR.t511 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2792 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t915 VPWR.t914 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2793 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t2519 VGND.t2518 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2794 VGND.t2429 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t2428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2795 VGND.t97 Vbias.t260 XA.XIR[6].XIC[14].icell.SM VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2796 VPWR.t1567 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t1566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2797 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t1563 VPWR.t1562 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2798 VPWR.t1747 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1746 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2799 VPWR.t591 VGND.t2705 XA.XIR[0].XIC[14].icell.PUM VPWR.t590 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2800 XA.XIR[15].XIC[2].icell.PDM VPWR.t2071 XA.XIR[15].XIC[2].icell.Ien VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2801 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t801 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2802 XThC.Tn[1].t8 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2803 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t23 VGND.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2804 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t2302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2805 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t800 VGND.t799 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2806 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t2350 VGND.t2349 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2807 VGND.t99 Vbias.t261 XA.XIR[0].XIC[4].icell.SM VGND.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2808 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t93 VGND.t911 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2809 XThC.Tn[14].t0 XThC.XTBN.Y.t120 VPWR.t1760 VPWR.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2810 VGND.t101 Vbias.t262 XA.XIR[5].XIC[10].icell.SM VGND.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2811 VGND.t103 Vbias.t263 XA.XIR[13].XIC[7].icell.SM VGND.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2812 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2072 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t1561 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2813 VGND.t744 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t743 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2814 VGND.t550 XThR.XTBN.Y.t120 a_n997_715# VGND.t549 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2815 VPWR.t1082 VPWR.t1080 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1081 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2816 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t589 VPWR.t588 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2817 VPWR.t1708 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t1707 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2818 VPWR.t135 XThR.XTB7.Y XThR.Tn[14].t4 VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t437 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2820 VGND.t1002 VGND.t1000 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t1001 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2821 VGND.t2203 Vbias.t264 XA.XIR[5].XIC[1].icell.SM VGND.t2202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2822 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t167 VGND.t1713 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2823 XThR.XTB6.A data[5].t5 VGND.t2316 VGND.t2315 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2824 XThR.Tn[0].t3 XThR.XTBN.Y.t121 a_n1049_8581# VPWR.t260 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2825 VGND.t1956 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t1955 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t913 VGND.t912 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2827 a_5949_9615# XThC.XTB6.Y VPWR.t984 VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2828 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t915 VGND.t914 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2829 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t172 VGND.t1805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2830 VGND.t1958 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t1957 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 VGND.t2107 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t2106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2832 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2833 VGND.t2365 XThC.XTBN.Y.t121 a_10051_9569# VGND.t487 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2834 VGND.t2205 Vbias.t265 XA.XIR[3].XIC[14].icell.SM VGND.t2204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2835 VGND.t2431 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2836 VGND.t196 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t195 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2837 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2073 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t1562 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2838 XA.XIR[15].XIC[6].icell.PDM VPWR.t2074 XA.XIR[15].XIC[6].icell.Ien VGND.t1563 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2839 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t916 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2840 XA.XIR[0].XIC[9].icell.PDM VGND.t997 VGND.t999 VGND.t998 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2841 VPWR.t1761 XThC.XTBN.Y.t122 XThC.Tn[11].t0 VPWR.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2842 VGND.t688 XThC.XTBN.Y.t123 a_7651_9569# VGND.t489 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2843 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1481 VPWR.t1480 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2844 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t236 VGND.t2433 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2845 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t513 VPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2846 XThR.Tn[2].t1 XThR.XTBN.Y.t122 VGND.t552 VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2847 VPWR.t133 XThR.XTB7.Y a_n1049_5317# VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2848 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t367 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2849 VGND.t2207 Vbias.t266 XA.XIR[15].XIC_15.icell.SM VGND.t2206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2850 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t10 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2852 VGND.t1484 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t1483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2853 VGND.t2187 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t2186 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2854 VPWR.t262 XThR.XTBN.Y.t123 XThR.Tn[12].t0 VPWR.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2855 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t798 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2856 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t2388 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2857 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t1712 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2858 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t160 VGND.t1668 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2859 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t2013 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2860 VPWR.t1079 VPWR.t1077 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1078 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2861 VGND.t1919 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2862 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t110 VGND.t1248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2863 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t2015 VGND.t2014 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2864 VGND.t2209 Vbias.t267 XA.XIR[13].XIC[2].icell.SM VGND.t2208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2865 VPWR.t1794 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t1793 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n458 VGND.n298 1.04433e+06
R1 VGND.n2851 VGND.n458 74066.7
R2 VGND.n2869 VGND.n2868 21134.4
R3 VGND.n2922 VGND.n2921 13477
R4 VGND.n2923 VGND.n2922 11635.6
R5 VGND.n2874 VGND.n104 9309.26
R6 VGND.n2921 VGND.n2920 9223.7
R7 VGND.n2920 VGND.n2919 9223.7
R8 VGND.n2918 VGND.n2917 9223.7
R9 VGND.n2917 VGND.n103 9223.7
R10 VGND.n2869 VGND.n298 8212.42
R11 VGND.n3007 VGND.n103 7447.41
R12 VGND.n2226 VGND.n2225 7387.65
R13 VGND.n2227 VGND.n2226 7387.65
R14 VGND.n2850 VGND.n491 7387.65
R15 VGND.n2871 VGND.n2870 7387.65
R16 VGND.n2872 VGND.n2871 7387.65
R17 VGND.n2873 VGND.n2872 7387.65
R18 VGND.n2875 VGND.n2873 7387.65
R19 VGND.n2875 VGND.n2874 7387.65
R20 VGND.n2851 VGND.n2850 6977.14
R21 VGND.n1717 VGND.t1498 6324.96
R22 VGND.n2870 VGND.n2869 5925.11
R23 VGND.n2919 VGND.n2918 5231.11
R24 VGND.n1321 VGND.t277 5168.13
R25 VGND.n3006 VGND.n104 5074.71
R26 VGND.n1626 VGND.n1625 4539.15
R27 VGND VGND.n104 4240.58
R28 VGND.n2741 VGND.n560 4077.12
R29 VGND.n1319 VGND.n1318 3417.39
R30 VGND.n1318 VGND.n1051 3417.39
R31 VGND.n1719 VGND.n1718 3417.39
R32 VGND.n2157 VGND.n806 3417.39
R33 VGND.n687 VGND.n521 3417.39
R34 VGND.n2849 VGND.n2848 3417.39
R35 VGND.n2924 VGND.n297 3417.39
R36 VGND.n2742 VGND.n2741 3331.79
R37 VGND.n2743 VGND.n2742 3331.79
R38 VGND.n2744 VGND.n2743 3331.79
R39 VGND.n2745 VGND.n2744 3331.79
R40 VGND.n2746 VGND.n2745 3331.79
R41 VGND.n2747 VGND.n2746 3331.79
R42 VGND.n2748 VGND.n2747 3331.79
R43 VGND.n2749 VGND.n2748 3331.79
R44 VGND.n2750 VGND.n2749 3331.79
R45 VGND.n2751 VGND.n2750 3331.79
R46 VGND.n2752 VGND.n2751 3331.79
R47 VGND.n2753 VGND.n2752 3331.79
R48 VGND.n2754 VGND.n2753 3331.79
R49 VGND.n2754 VGND.n101 3331.79
R50 VGND.n3009 VGND.n101 3331.79
R51 VGND.n3009 VGND.n3008 3331.79
R52 VGND.n1626 VGND.n1051 3273.91
R53 VGND.n2158 VGND.n841 3265.22
R54 VGND.n2923 VGND.n298 3096.3
R55 VGND.n2848 VGND.n458 2756.52
R56 VGND.n2921 VGND.t582 2655.17
R57 VGND.n2920 VGND.t576 2655.17
R58 VGND.n3008 VGND.n3007 2602.7
R59 VGND.n2850 VGND.n2849 2517.39
R60 VGND.n1320 VGND.n1319 2173.91
R61 VGND.n2867 VGND.n453 2097.71
R62 VGND.n2867 VGND.n454 2097.71
R63 VGND.n2862 VGND.n454 2097.71
R64 VGND.n2862 VGND.n453 2097.71
R65 VGND.n2852 VGND.n452 2097.71
R66 VGND.n2853 VGND.n452 2097.71
R67 VGND.n2860 VGND.n2853 2097.71
R68 VGND.n2860 VGND.n2852 2097.71
R69 VGND.n2924 VGND.n2923 2082.61
R70 VGND.n2918 VGND 1997.7
R71 VGND.n2917 VGND 1997.7
R72 VGND VGND.n103 1997.7
R73 VGND.n2228 VGND.n491 1831.57
R74 VGND.n2919 VGND.t662 1807.04
R75 VGND.n126 VGND.t1665 1785.51
R76 VGND.n2227 VGND.n806 1691.3
R77 VGND.n2876 VGND.t64 1618.39
R78 VGND.t709 VGND.n2916 1618.39
R79 VGND.n127 VGND.t1254 1618.39
R80 VGND.n2922 VGND.t516 1517.24
R81 VGND.n2225 VGND.n842 1513.49
R82 VGND.n1717 VGND.n842 1370.36
R83 VGND.t998 VGND.n842 1270.28
R84 VGND.n1596 VGND.t487 1268.93
R85 VGND.n1596 VGND.t1283 1268.93
R86 VGND.n490 VGND.t474 1253.59
R87 VGND.t335 VGND.n490 1253.59
R88 VGND.n840 VGND.t77 1253.59
R89 VGND.t481 VGND.n840 1253.59
R90 VGND.n2224 VGND.t478 1253.59
R91 VGND.t489 VGND.n2224 1253.59
R92 VGND.n1716 VGND.t670 1253.59
R93 VGND.t547 VGND.n1716 1253.59
R94 VGND.n520 VGND.t79 1253.59
R95 VGND.t957 VGND.n520 1253.59
R96 VGND.n1321 VGND.n1320 1243.48
R97 VGND.t1043 VGND.n2228 1237.71
R98 VGND.n2876 VGND.t1246 1213.79
R99 VGND.n1625 VGND.n1624 1198.25
R100 VGND.n3006 VGND.n3005 1198.25
R101 VGND.n2734 VGND.n559 1180.79
R102 VGND.n2999 VGND.n102 1180.79
R103 VGND.n2827 VGND.n2826 1180.79
R104 VGND.n2756 VGND.n2755 1180.79
R105 VGND.n2639 VGND.n548 1180.79
R106 VGND.n2409 VGND.n549 1180.79
R107 VGND.n2404 VGND.n550 1180.79
R108 VGND.n2664 VGND.n551 1180.79
R109 VGND.n2127 VGND.n552 1180.79
R110 VGND.n2122 VGND.n553 1180.79
R111 VGND.n2689 VGND.n554 1180.79
R112 VGND.n1900 VGND.n555 1180.79
R113 VGND.n1895 VGND.n556 1180.79
R114 VGND.n2714 VGND.n557 1180.79
R115 VGND.n1288 VGND.n558 1180.79
R116 VGND.n3011 VGND.n3010 1180.79
R117 VGND.n1511 VGND.n560 1180.79
R118 VGND.n2740 VGND.n2739 1180.79
R119 VGND.n1330 VGND.n1329 1180.46
R120 VGND.n1397 VGND.n1396 1180.46
R121 VGND.n1395 VGND.n1394 1180.46
R122 VGND.n1390 VGND.n1389 1180.46
R123 VGND.n1385 VGND.n1384 1180.46
R124 VGND.n1380 VGND.n1379 1180.46
R125 VGND.n1375 VGND.n1374 1180.46
R126 VGND.n1370 VGND.n1369 1180.46
R127 VGND.n1365 VGND.n1364 1180.46
R128 VGND.n1360 VGND.n1359 1180.46
R129 VGND.n1355 VGND.n1354 1180.46
R130 VGND.n1350 VGND.n1349 1180.46
R131 VGND.n1345 VGND.n1344 1180.46
R132 VGND.n1340 VGND.n1339 1180.46
R133 VGND.n1335 VGND.n1334 1180.46
R134 VGND.n1508 VGND.n1507 1180.46
R135 VGND.n1506 VGND.n1505 1180.46
R136 VGND.n1489 VGND.n1488 1180.46
R137 VGND.n1487 VGND.n1486 1180.46
R138 VGND.n1476 VGND.n1475 1180.46
R139 VGND.n1474 VGND.n1473 1180.46
R140 VGND.n1457 VGND.n1456 1180.46
R141 VGND.n1455 VGND.n1454 1180.46
R142 VGND.n1444 VGND.n1443 1180.46
R143 VGND.n1442 VGND.n1441 1180.46
R144 VGND.n1425 VGND.n1424 1180.46
R145 VGND.n1423 VGND.n1422 1180.46
R146 VGND.n1411 VGND.n1064 1180.46
R147 VGND.n1566 VGND.n1565 1180.46
R148 VGND.n1568 VGND.n1567 1180.46
R149 VGND.n1145 VGND.n1144 1180.46
R150 VGND.n1150 VGND.n1149 1180.46
R151 VGND.n1202 VGND.n1201 1180.46
R152 VGND.n1200 VGND.n1199 1180.46
R153 VGND.n1195 VGND.n1194 1180.46
R154 VGND.n1190 VGND.n1189 1180.46
R155 VGND.n1185 VGND.n1184 1180.46
R156 VGND.n1180 VGND.n1179 1180.46
R157 VGND.n1175 VGND.n1174 1180.46
R158 VGND.n1170 VGND.n1169 1180.46
R159 VGND.n1165 VGND.n1164 1180.46
R160 VGND.n1160 VGND.n1159 1180.46
R161 VGND.n1155 VGND.n1154 1180.46
R162 VGND.n2729 VGND.n2728 1180.46
R163 VGND.n2731 VGND.n2730 1180.46
R164 VGND.n2926 VGND.n2925 1180.46
R165 VGND.n2934 VGND.n2933 1180.46
R166 VGND.n2936 VGND.n2935 1180.46
R167 VGND.n2944 VGND.n2943 1180.46
R168 VGND.n2946 VGND.n2945 1180.46
R169 VGND.n2954 VGND.n2953 1180.46
R170 VGND.n2956 VGND.n2955 1180.46
R171 VGND.n2964 VGND.n2963 1180.46
R172 VGND.n2966 VGND.n2965 1180.46
R173 VGND.n2974 VGND.n2973 1180.46
R174 VGND.n2976 VGND.n2975 1180.46
R175 VGND.n2984 VGND.n2983 1180.46
R176 VGND.n2986 VGND.n2985 1180.46
R177 VGND.n2994 VGND.n2993 1180.46
R178 VGND.n2996 VGND.n2995 1180.46
R179 VGND.n2847 VGND.n2846 1180.46
R180 VGND.n2760 VGND.n526 1180.46
R181 VGND.n2765 VGND.n2764 1180.46
R182 VGND.n2770 VGND.n2769 1180.46
R183 VGND.n2775 VGND.n2774 1180.46
R184 VGND.n2780 VGND.n2779 1180.46
R185 VGND.n2785 VGND.n2784 1180.46
R186 VGND.n2790 VGND.n2789 1180.46
R187 VGND.n2795 VGND.n2794 1180.46
R188 VGND.n2800 VGND.n2799 1180.46
R189 VGND.n2805 VGND.n2804 1180.46
R190 VGND.n2810 VGND.n2809 1180.46
R191 VGND.n2815 VGND.n2814 1180.46
R192 VGND.n2820 VGND.n2819 1180.46
R193 VGND.n2825 VGND.n2824 1180.46
R194 VGND.n2448 VGND.n2447 1180.46
R195 VGND.n2472 VGND.n2471 1180.46
R196 VGND.n2474 VGND.n2473 1180.46
R197 VGND.n2498 VGND.n2497 1180.46
R198 VGND.n2500 VGND.n2499 1180.46
R199 VGND.n2524 VGND.n2523 1180.46
R200 VGND.n2526 VGND.n2525 1180.46
R201 VGND.n2550 VGND.n2549 1180.46
R202 VGND.n2552 VGND.n2551 1180.46
R203 VGND.n2576 VGND.n2575 1180.46
R204 VGND.n2578 VGND.n2577 1180.46
R205 VGND.n2607 VGND.n2606 1180.46
R206 VGND.n2612 VGND.n2611 1180.46
R207 VGND.n2617 VGND.n2616 1180.46
R208 VGND.n2619 VGND.n2618 1180.46
R209 VGND.n2459 VGND.n2458 1180.46
R210 VGND.n2461 VGND.n2460 1180.46
R211 VGND.n2485 VGND.n2484 1180.46
R212 VGND.n2487 VGND.n2486 1180.46
R213 VGND.n2511 VGND.n2510 1180.46
R214 VGND.n2513 VGND.n2512 1180.46
R215 VGND.n2537 VGND.n2536 1180.46
R216 VGND.n2539 VGND.n2538 1180.46
R217 VGND.n2563 VGND.n2562 1180.46
R218 VGND.n2565 VGND.n2564 1180.46
R219 VGND.n2589 VGND.n2588 1180.46
R220 VGND.n2596 VGND.n2595 1180.46
R221 VGND.n2594 VGND.n2593 1180.46
R222 VGND.n2634 VGND.n2633 1180.46
R223 VGND.n2636 VGND.n2635 1180.46
R224 VGND.n692 VGND.n691 1180.46
R225 VGND.n697 VGND.n696 1180.46
R226 VGND.n702 VGND.n701 1180.46
R227 VGND.n707 VGND.n706 1180.46
R228 VGND.n712 VGND.n711 1180.46
R229 VGND.n717 VGND.n716 1180.46
R230 VGND.n722 VGND.n721 1180.46
R231 VGND.n727 VGND.n726 1180.46
R232 VGND.n732 VGND.n731 1180.46
R233 VGND.n737 VGND.n736 1180.46
R234 VGND.n742 VGND.n741 1180.46
R235 VGND.n747 VGND.n746 1180.46
R236 VGND.n2420 VGND.n2419 1180.46
R237 VGND.n2418 VGND.n2417 1180.46
R238 VGND.n2413 VGND.n2412 1180.46
R239 VGND.n2230 VGND.n2229 1180.46
R240 VGND.n2254 VGND.n2253 1180.46
R241 VGND.n2256 VGND.n2255 1180.46
R242 VGND.n2280 VGND.n2279 1180.46
R243 VGND.n2282 VGND.n2281 1180.46
R244 VGND.n2306 VGND.n2305 1180.46
R245 VGND.n2308 VGND.n2307 1180.46
R246 VGND.n2332 VGND.n2331 1180.46
R247 VGND.n2334 VGND.n2333 1180.46
R248 VGND.n2358 VGND.n2357 1180.46
R249 VGND.n2360 VGND.n2359 1180.46
R250 VGND.n2389 VGND.n2388 1180.46
R251 VGND.n2394 VGND.n2393 1180.46
R252 VGND.n2399 VGND.n2398 1180.46
R253 VGND.n2401 VGND.n2400 1180.46
R254 VGND.n2241 VGND.n2240 1180.46
R255 VGND.n2243 VGND.n2242 1180.46
R256 VGND.n2267 VGND.n2266 1180.46
R257 VGND.n2269 VGND.n2268 1180.46
R258 VGND.n2293 VGND.n2292 1180.46
R259 VGND.n2295 VGND.n2294 1180.46
R260 VGND.n2319 VGND.n2318 1180.46
R261 VGND.n2321 VGND.n2320 1180.46
R262 VGND.n2345 VGND.n2344 1180.46
R263 VGND.n2347 VGND.n2346 1180.46
R264 VGND.n2371 VGND.n2370 1180.46
R265 VGND.n2378 VGND.n2377 1180.46
R266 VGND.n2376 VGND.n2375 1180.46
R267 VGND.n2659 VGND.n2658 1180.46
R268 VGND.n2661 VGND.n2660 1180.46
R269 VGND.n2156 VGND.n2155 1180.46
R270 VGND.n869 VGND.n852 1180.46
R271 VGND.n874 VGND.n873 1180.46
R272 VGND.n879 VGND.n878 1180.46
R273 VGND.n884 VGND.n883 1180.46
R274 VGND.n889 VGND.n888 1180.46
R275 VGND.n894 VGND.n893 1180.46
R276 VGND.n899 VGND.n898 1180.46
R277 VGND.n904 VGND.n903 1180.46
R278 VGND.n909 VGND.n908 1180.46
R279 VGND.n914 VGND.n913 1180.46
R280 VGND.n919 VGND.n918 1180.46
R281 VGND.n2138 VGND.n2137 1180.46
R282 VGND.n2136 VGND.n2135 1180.46
R283 VGND.n2131 VGND.n2130 1180.46
R284 VGND.n1948 VGND.n1947 1180.46
R285 VGND.n1972 VGND.n1971 1180.46
R286 VGND.n1974 VGND.n1973 1180.46
R287 VGND.n1998 VGND.n1997 1180.46
R288 VGND.n2000 VGND.n1999 1180.46
R289 VGND.n2024 VGND.n2023 1180.46
R290 VGND.n2026 VGND.n2025 1180.46
R291 VGND.n2050 VGND.n2049 1180.46
R292 VGND.n2052 VGND.n2051 1180.46
R293 VGND.n2076 VGND.n2075 1180.46
R294 VGND.n2078 VGND.n2077 1180.46
R295 VGND.n2107 VGND.n2106 1180.46
R296 VGND.n2112 VGND.n2111 1180.46
R297 VGND.n2117 VGND.n2116 1180.46
R298 VGND.n2119 VGND.n2118 1180.46
R299 VGND.n1959 VGND.n1958 1180.46
R300 VGND.n1961 VGND.n1960 1180.46
R301 VGND.n1985 VGND.n1984 1180.46
R302 VGND.n1987 VGND.n1986 1180.46
R303 VGND.n2011 VGND.n2010 1180.46
R304 VGND.n2013 VGND.n2012 1180.46
R305 VGND.n2037 VGND.n2036 1180.46
R306 VGND.n2039 VGND.n2038 1180.46
R307 VGND.n2063 VGND.n2062 1180.46
R308 VGND.n2065 VGND.n2064 1180.46
R309 VGND.n2089 VGND.n2088 1180.46
R310 VGND.n2096 VGND.n2095 1180.46
R311 VGND.n2094 VGND.n2093 1180.46
R312 VGND.n2684 VGND.n2683 1180.46
R313 VGND.n2686 VGND.n2685 1180.46
R314 VGND.n1686 VGND.n1685 1180.46
R315 VGND.n1681 VGND.n1680 1180.46
R316 VGND.n1676 VGND.n1675 1180.46
R317 VGND.n1671 VGND.n1670 1180.46
R318 VGND.n1666 VGND.n1665 1180.46
R319 VGND.n1661 VGND.n1660 1180.46
R320 VGND.n1656 VGND.n1655 1180.46
R321 VGND.n1651 VGND.n1650 1180.46
R322 VGND.n1646 VGND.n1645 1180.46
R323 VGND.n1641 VGND.n1640 1180.46
R324 VGND.n1636 VGND.n1635 1180.46
R325 VGND.n1631 VGND.n1630 1180.46
R326 VGND.n1911 VGND.n1910 1180.46
R327 VGND.n1909 VGND.n1908 1180.46
R328 VGND.n1904 VGND.n1903 1180.46
R329 VGND.n1721 VGND.n1720 1180.46
R330 VGND.n1745 VGND.n1744 1180.46
R331 VGND.n1747 VGND.n1746 1180.46
R332 VGND.n1771 VGND.n1770 1180.46
R333 VGND.n1773 VGND.n1772 1180.46
R334 VGND.n1797 VGND.n1796 1180.46
R335 VGND.n1799 VGND.n1798 1180.46
R336 VGND.n1823 VGND.n1822 1180.46
R337 VGND.n1825 VGND.n1824 1180.46
R338 VGND.n1849 VGND.n1848 1180.46
R339 VGND.n1851 VGND.n1850 1180.46
R340 VGND.n1880 VGND.n1879 1180.46
R341 VGND.n1885 VGND.n1884 1180.46
R342 VGND.n1890 VGND.n1889 1180.46
R343 VGND.n1892 VGND.n1891 1180.46
R344 VGND.n1732 VGND.n1731 1180.46
R345 VGND.n1734 VGND.n1733 1180.46
R346 VGND.n1758 VGND.n1757 1180.46
R347 VGND.n1760 VGND.n1759 1180.46
R348 VGND.n1784 VGND.n1783 1180.46
R349 VGND.n1786 VGND.n1785 1180.46
R350 VGND.n1810 VGND.n1809 1180.46
R351 VGND.n1812 VGND.n1811 1180.46
R352 VGND.n1836 VGND.n1835 1180.46
R353 VGND.n1838 VGND.n1837 1180.46
R354 VGND.n1862 VGND.n1861 1180.46
R355 VGND.n1869 VGND.n1868 1180.46
R356 VGND.n1867 VGND.n1866 1180.46
R357 VGND.n2709 VGND.n2708 1180.46
R358 VGND.n2711 VGND.n2710 1180.46
R359 VGND.n1317 VGND.n1316 1180.46
R360 VGND.n1234 VGND.n1132 1180.46
R361 VGND.n1239 VGND.n1238 1180.46
R362 VGND.n1244 VGND.n1243 1180.46
R363 VGND.n1249 VGND.n1248 1180.46
R364 VGND.n1254 VGND.n1253 1180.46
R365 VGND.n1259 VGND.n1258 1180.46
R366 VGND.n1264 VGND.n1263 1180.46
R367 VGND.n1269 VGND.n1268 1180.46
R368 VGND.n1274 VGND.n1273 1180.46
R369 VGND.n1279 VGND.n1278 1180.46
R370 VGND.n1284 VGND.n1283 1180.46
R371 VGND.n1299 VGND.n1298 1180.46
R372 VGND.n1297 VGND.n1296 1180.46
R373 VGND.n1292 VGND.n1291 1180.46
R374 VGND.n296 VGND.n295 1180.46
R375 VGND.n291 VGND.n290 1180.46
R376 VGND.n286 VGND.n285 1180.46
R377 VGND.n281 VGND.n280 1180.46
R378 VGND.n276 VGND.n275 1180.46
R379 VGND.n271 VGND.n270 1180.46
R380 VGND.n266 VGND.n265 1180.46
R381 VGND.n261 VGND.n260 1180.46
R382 VGND.n256 VGND.n255 1180.46
R383 VGND.n251 VGND.n250 1180.46
R384 VGND.n246 VGND.n245 1180.46
R385 VGND.n241 VGND.n240 1180.46
R386 VGND.n236 VGND.n235 1180.46
R387 VGND.n231 VGND.n230 1180.46
R388 VGND.n226 VGND.n225 1180.46
R389 VGND.n2916 VGND.t1245 1180.08
R390 VGND.n1718 VGND.n1717 1169.57
R391 VGND.n2872 VGND.t51 1146.36
R392 VGND.n2870 VGND.t50 1112.64
R393 VGND.n2871 VGND.t836 1112.64
R394 VGND.n3007 VGND 1055.35
R395 VGND.n2228 VGND.n2227 1052.29
R396 VGND.n2861 VGND.t1164 1041.38
R397 VGND.n2868 VGND.t1164 1041.38
R398 VGND.t511 VGND.n2158 1032.59
R399 VGND.t532 VGND.n1145 988.926
R400 VGND.t539 VGND.n1150 988.926
R401 VGND.n1201 VGND.t859 988.926
R402 VGND.n1200 VGND.t1944 988.926
R403 VGND.n1195 VGND.t884 988.926
R404 VGND.n1190 VGND.t2269 988.926
R405 VGND.n1185 VGND.t108 988.926
R406 VGND.n1180 VGND.t2309 988.926
R407 VGND.n1175 VGND.t2034 988.926
R408 VGND.n1170 VGND.t613 988.926
R409 VGND.n1165 VGND.t464 988.926
R410 VGND.n1160 VGND.t1692 988.926
R411 VGND.n1155 VGND.t912 988.926
R412 VGND.t2476 VGND.n2729 988.926
R413 VGND.n2730 VGND.t1885 988.926
R414 VGND.n2925 VGND.t509 988.926
R415 VGND.t305 VGND.n2934 988.926
R416 VGND.n2935 VGND.t283 988.926
R417 VGND.t507 VGND.n2944 988.926
R418 VGND.n2945 VGND.t496 988.926
R419 VGND.t1544 VGND.n2954 988.926
R420 VGND.n2955 VGND.t1387 988.926
R421 VGND.t1364 VGND.n2964 988.926
R422 VGND.n2965 VGND.t1540 988.926
R423 VGND.t267 VGND.n2974 988.926
R424 VGND.n2975 VGND.t255 988.926
R425 VGND.t1335 VGND.n2984 988.926
R426 VGND.n2985 VGND.t1527 988.926
R427 VGND.t243 VGND.n2994 988.926
R428 VGND.n2995 VGND.t1349 988.926
R429 VGND.n2847 VGND.t2286 988.926
R430 VGND.t1500 VGND.n2760 988.926
R431 VGND.t1474 VGND.n2765 988.926
R432 VGND.t1424 VGND.n2770 988.926
R433 VGND.t2296 VGND.n2775 988.926
R434 VGND.t759 VGND.n2780 988.926
R435 VGND.t867 VGND.n2785 988.926
R436 VGND.t6 VGND.n2790 988.926
R437 VGND.t183 VGND.n2795 988.926
R438 VGND.t694 VGND.n2800 988.926
R439 VGND.t1488 VGND.n2805 988.926
R440 VGND.t2469 VGND.n2810 988.926
R441 VGND.t1938 VGND.n2815 988.926
R442 VGND.t13 VGND.n2820 988.926
R443 VGND.t995 VGND.n2825 988.926
R444 VGND.n2447 VGND.t1302 988.926
R445 VGND.t2136 VGND.n2472 988.926
R446 VGND.n2473 VGND.t2591 988.926
R447 VGND.t2408 VGND.n2498 988.926
R448 VGND.n2499 VGND.t1754 988.926
R449 VGND.t2419 VGND.n2524 988.926
R450 VGND.n2525 VGND.t2493 988.926
R451 VGND.t1264 VGND.n2550 988.926
R452 VGND.n2551 VGND.t2025 988.926
R453 VGND.t2576 VGND.n2576 988.926
R454 VGND.n2577 VGND.t2069 988.926
R455 VGND.t2084 VGND.n2607 988.926
R456 VGND.t413 VGND.n2612 988.926
R457 VGND.t2002 VGND.n2617 988.926
R458 VGND.n2618 VGND.t2327 988.926
R459 VGND.t535 VGND.n2459 988.926
R460 VGND.n2460 VGND.t543 988.926
R461 VGND.t857 VGND.n2485 988.926
R462 VGND.n2486 VGND.t1946 988.926
R463 VGND.t888 VGND.n2511 988.926
R464 VGND.n2512 VGND.t2498 988.926
R465 VGND.t114 VGND.n2537 988.926
R466 VGND.n2538 VGND.t1565 988.926
R467 VGND.t1926 VGND.n2563 988.926
R468 VGND.n2564 VGND.t617 988.926
R469 VGND.t468 VGND.n2589 988.926
R470 VGND.n2595 VGND.t1696 988.926
R471 VGND.n2594 VGND.t1989 988.926
R472 VGND.t1825 VGND.n2634 988.926
R473 VGND.n2635 VGND.t1889 988.926
R474 VGND.t1519 VGND.n692 988.926
R475 VGND.t2141 VGND.n697 988.926
R476 VGND.t896 VGND.n702 988.926
R477 VGND.t1417 VGND.n707 988.926
R478 VGND.t354 VGND.n712 988.926
R479 VGND.t755 VGND.n717 988.926
R480 VGND.t2386 VGND.n722 988.926
R481 VGND.t163 VGND.n727 988.926
R482 VGND.t1272 VGND.n732 988.926
R483 VGND.t689 VGND.n737 988.926
R484 VGND.t1902 VGND.n742 988.926
R485 VGND.t2079 VGND.n747 988.926
R486 VGND.n2419 VGND.t1932 988.926
R487 VGND.n2418 VGND.t8 988.926
R488 VGND.n2413 VGND.t988 988.926
R489 VGND.n2229 VGND.t1600 988.926
R490 VGND.t830 VGND.n2254 988.926
R491 VGND.n2255 VGND.t796 988.926
R492 VGND.t2399 VGND.n2280 988.926
R493 VGND.n2281 VGND.t2258 988.926
R494 VGND.t360 VGND.n2306 988.926
R495 VGND.n2307 VGND.t2485 988.926
R496 VGND.t890 VGND.n2332 988.926
R497 VGND.n2333 VGND.t2017 988.926
R498 VGND.t2007 VGND.n2358 988.926
R499 VGND.n2359 VGND.t1486 988.926
R500 VGND.t124 VGND.n2389 988.926
R501 VGND.t405 VGND.n2394 988.926
R502 VGND.t173 VGND.n2399 988.926
R503 VGND.n2400 VGND.t1895 988.926
R504 VGND.t1304 VGND.n2241 988.926
R505 VGND.n2242 VGND.t2138 988.926
R506 VGND.t2589 VGND.n2267 988.926
R507 VGND.n2268 VGND.t1569 988.926
R508 VGND.t1756 VGND.n2293 988.926
R509 VGND.n2294 VGND.t2421 988.926
R510 VGND.t2495 VGND.n2319 988.926
R511 VGND.n2320 VGND.t1266 988.926
R512 VGND.t1277 VGND.n2345 988.926
R513 VGND.n2346 VGND.t2578 988.926
R514 VGND.t2518 VGND.n2371 988.926
R515 VGND.n2377 VGND.t2086 988.926
R516 VGND.n2376 VGND.t415 988.926
R517 VGND.t2004 VGND.n2659 988.926
R518 VGND.n2660 VGND.t2329 988.926
R519 VGND.n2156 VGND.t537 988.926
R520 VGND.t545 VGND.n869 988.926
R521 VGND.t855 VGND.n874 988.926
R522 VGND.t1948 VGND.n879 988.926
R523 VGND.t2389 VGND.n884 988.926
R524 VGND.t2500 VGND.n889 988.926
R525 VGND.t116 VGND.n894 988.926
R526 VGND.t1567 VGND.n899 988.926
R527 VGND.t1928 VGND.n904 988.926
R528 VGND.t619 VGND.n909 988.926
R529 VGND.t470 VGND.n914 988.926
R530 VGND.t1698 VGND.n919 988.926
R531 VGND.n2137 VGND.t1991 988.926
R532 VGND.n2136 VGND.t1827 988.926
R533 VGND.n2131 VGND.t1891 988.926
R534 VGND.n1947 VGND.t530 988.926
R535 VGND.t2685 VGND.n1972 988.926
R536 VGND.n1973 VGND.t861 988.926
R537 VGND.t1942 VGND.n1998 988.926
R538 VGND.n1999 VGND.t882 988.926
R539 VGND.t2271 VGND.n2024 988.926
R540 VGND.n2025 VGND.t110 988.926
R541 VGND.t2311 VGND.n2050 988.926
R542 VGND.n2051 VGND.t2036 988.926
R543 VGND.t615 VGND.n2076 988.926
R544 VGND.n2077 VGND.t466 988.926
R545 VGND.t1694 VGND.n2107 988.926
R546 VGND.t914 VGND.n2112 988.926
R547 VGND.t2474 VGND.n2117 988.926
R548 VGND.n2118 VGND.t1887 988.926
R549 VGND.t1517 VGND.n1959 988.926
R550 VGND.n1960 VGND.t1793 988.926
R551 VGND.t898 VGND.n1985 988.926
R552 VGND.n1986 VGND.t1415 988.926
R553 VGND.t2071 VGND.n2011 988.926
R554 VGND.n2012 VGND.t753 988.926
R555 VGND.t2384 VGND.n2037 988.926
R556 VGND.n2038 VGND.t161 988.926
R557 VGND.t1270 VGND.n2063 988.926
R558 VGND.n2064 VGND.t2582 988.926
R559 VGND.t1900 VGND.n2089 988.926
R560 VGND.n2095 VGND.t2077 988.926
R561 VGND.n2094 VGND.t1930 988.926
R562 VGND.t16 VGND.n2684 988.926
R563 VGND.n2685 VGND.t986 988.926
R564 VGND.n1686 VGND.t1523 988.926
R565 VGND.n1681 VGND.t1812 988.926
R566 VGND.n1676 VGND.t69 988.926
R567 VGND.n1671 VGND.t1311 988.926
R568 VGND.n1666 VGND.t2349 988.926
R569 VGND.n1661 VGND.t777 988.926
R570 VGND.n1656 VGND.t849 988.926
R571 VGND.n1651 VGND.t1319 988.926
R572 VGND.n1646 VGND.t982 988.926
R573 VGND.n1641 VGND.t561 988.926
R574 VGND.n1636 VGND.t374 988.926
R575 VGND.n1631 VGND.t1993 988.926
R576 VGND.n1910 VGND.t433 988.926
R577 VGND.n1909 VGND.t2612 988.926
R578 VGND.n1904 VGND.t904 988.926
R579 VGND.n1720 VGND.t1606 988.926
R580 VGND.t2134 VGND.n1745 988.926
R581 VGND.n1746 VGND.t2593 988.926
R582 VGND.t2406 VGND.n1771 988.926
R583 VGND.n1772 VGND.t1752 988.926
R584 VGND.t2417 VGND.n1797 988.926
R585 VGND.n1798 VGND.t2491 988.926
R586 VGND.t1262 VGND.n1823 988.926
R587 VGND.n1824 VGND.t2023 988.926
R588 VGND.t2014 VGND.n1849 988.926
R589 VGND.n1850 VGND.t2067 988.926
R590 VGND.t2082 VGND.n1880 988.926
R591 VGND.t411 VGND.n1885 988.926
R592 VGND.t2000 VGND.n1890 988.926
R593 VGND.n1891 VGND.t2325 988.926
R594 VGND.t1521 VGND.n1732 988.926
R595 VGND.n1733 VGND.t1810 988.926
R596 VGND.t71 VGND.n1758 988.926
R597 VGND.n1759 VGND.t1309 988.926
R598 VGND.t2347 VGND.n1784 988.926
R599 VGND.n1785 VGND.t775 988.926
R600 VGND.t847 VGND.n1810 988.926
R601 VGND.n1811 VGND.t1317 988.926
R602 VGND.t771 VGND.n1836 988.926
R603 VGND.n1837 VGND.t559 988.926
R604 VGND.t372 VGND.n1862 988.926
R605 VGND.n1868 VGND.t1704 988.926
R606 VGND.n1867 VGND.t431 988.926
R607 VGND.t2610 VGND.n2709 988.926
R608 VGND.n2710 VGND.t902 988.926
R609 VGND.n1317 VGND.t2284 988.926
R610 VGND.t2145 VGND.n1234 988.926
R611 VGND.t1477 VGND.n1239 988.926
R612 VGND.t1421 VGND.n1244 988.926
R613 VGND.t358 VGND.n1249 988.926
R614 VGND.t757 VGND.n1254 988.926
R615 VGND.t865 VGND.n1259 988.926
R616 VGND.t4 VGND.n1264 988.926
R617 VGND.t181 VGND.n1269 988.926
R618 VGND.t691 VGND.n1274 988.926
R619 VGND.t1904 VGND.n1279 988.926
R620 VGND.t2073 VGND.n1284 988.926
R621 VGND.n1298 VGND.t1936 988.926
R622 VGND.n1297 VGND.t10 988.926
R623 VGND.n1292 VGND.t992 988.926
R624 VGND.n296 VGND.t1602 988.926
R625 VGND.n291 VGND.t832 988.926
R626 VGND.n286 VGND.t799 988.926
R627 VGND.n281 VGND.t2401 988.926
R628 VGND.n276 VGND.t2260 988.926
R629 VGND.n271 VGND.t362 988.926
R630 VGND.n266 VGND.t2487 988.926
R631 VGND.n261 VGND.t892 988.926
R632 VGND.n256 VGND.t2019 988.926
R633 VGND.n251 VGND.t2010 988.926
R634 VGND.n246 VGND.t2063 988.926
R635 VGND.n241 VGND.t127 988.926
R636 VGND.n236 VGND.t407 988.926
R637 VGND.n231 VGND.t176 988.926
R638 VGND.n226 VGND.t2320 988.926
R639 VGND.t331 VGND.n1330 988.926
R640 VGND.n1396 VGND.t249 988.926
R641 VGND.n1395 VGND.t1401 988.926
R642 VGND.n1390 VGND.t326 988.926
R643 VGND.n1385 VGND.t315 988.926
R644 VGND.n1380 VGND.t296 988.926
R645 VGND.n1375 VGND.t1329 988.926
R646 VGND.n1370 VGND.t498 988.926
R647 VGND.n1365 VGND.t292 988.926
R648 VGND.n1360 VGND.t1389 988.926
R649 VGND.n1355 VGND.t1376 988.926
R650 VGND.n1350 VGND.t1542 988.926
R651 VGND.n1345 VGND.t275 988.926
R652 VGND.n1340 VGND.t1358 988.926
R653 VGND.n1335 VGND.t1551 988.926
R654 VGND.n2225 VGND.n841 934.784
R655 VGND VGND.n391 927.203
R656 VGND VGND.n358 927.203
R657 VGND.n2159 VGND 918.774
R658 VGND VGND.n451 910.346
R659 VGND VGND.n422 910.346
R660 VGND.t235 VGND.n3006 909.365
R661 VGND.n2850 VGND.n521 900
R662 VGND.n1145 VGND.t1525 852.769
R663 VGND.n1150 VGND.t1663 852.769
R664 VGND.n1201 VGND.t40 852.769
R665 VGND.t1 VGND.n1200 852.769
R666 VGND.t2335 VGND.n1195 852.769
R667 VGND.t44 VGND.n1190 852.769
R668 VGND.t2435 VGND.n1185 852.769
R669 VGND.t2434 VGND.n1180 852.769
R670 VGND.t2303 VGND.n1175 852.769
R671 VGND.t2396 VGND.n1170 852.769
R672 VGND.t1952 VGND.n1165 852.769
R673 VGND.t167 VGND.n1160 852.769
R674 VGND.t2586 VGND.n1155 852.769
R675 VGND.n2729 VGND.t48 852.769
R676 VGND.n2730 VGND.t172 852.769
R677 VGND.t2334 VGND.n559 852.769
R678 VGND.n2925 VGND.t2305 852.769
R679 VGND.n2934 VGND.t1574 852.769
R680 VGND.n2935 VGND.t1814 852.769
R681 VGND.n2944 VGND.t1598 852.769
R682 VGND.n2945 VGND.t1920 852.769
R683 VGND.n2954 VGND.t2367 852.769
R684 VGND.n2955 VGND.t178 852.769
R685 VGND.n2964 VGND.t105 852.769
R686 VGND.n2965 VGND.t1818 852.769
R687 VGND.n2974 VGND.t834 852.769
R688 VGND.n2975 VGND.t2395 852.769
R689 VGND.n2984 VGND.t1227 852.769
R690 VGND.n2985 VGND.t1608 852.769
R691 VGND.n2994 VGND.t1859 852.769
R692 VGND.n2995 VGND.t1986 852.769
R693 VGND.t973 VGND.n102 852.769
R694 VGND.t2564 VGND.n2847 852.769
R695 VGND.n2760 VGND.t1950 852.769
R696 VGND.n2765 VGND.t238 852.769
R697 VGND.n2770 VGND.t1824 852.769
R698 VGND.n2775 VGND.t43 852.769
R699 VGND.n2780 VGND.t979 852.769
R700 VGND.n2785 VGND.t1241 852.769
R701 VGND.n2790 VGND.t1481 852.769
R702 VGND.n2795 VGND.t1526 852.769
R703 VGND.n2800 VGND.t495 852.769
R704 VGND.n2805 VGND.t2559 852.769
R705 VGND.n2810 VGND.t840 852.769
R706 VGND.n2815 VGND.t2333 852.769
R707 VGND.n2820 VGND.t30 852.769
R708 VGND.n2825 VGND.t1997 852.769
R709 VGND.n2826 VGND.t2089 852.769
R710 VGND.n2447 VGND.t223 852.769
R711 VGND.n2472 VGND.t1668 852.769
R712 VGND.n2473 VGND.t221 852.769
R713 VGND.n2498 VGND.t1804 852.769
R714 VGND.n2499 VGND.t2300 852.769
R715 VGND.n2524 VGND.t378 852.769
R716 VGND.n2525 VGND.t2029 852.769
R717 VGND.n2550 VGND.t1908 852.769
R718 VGND.n2551 VGND.t353 852.769
R719 VGND.n2576 VGND.t926 852.769
R720 VGND.n2577 VGND.t917 852.769
R721 VGND.n2607 VGND.t716 852.769
R722 VGND.n2612 VGND.t46 852.769
R723 VGND.n2617 VGND.t1816 852.769
R724 VGND.n2618 VGND.t2332 852.769
R725 VGND.n2755 VGND.t956 852.769
R726 VGND.n2459 VGND.t493 852.769
R727 VGND.n2460 VGND.t1269 852.769
R728 VGND.n2485 VGND.t1637 852.769
R729 VGND.n2486 VGND.t186 852.769
R730 VGND.n2511 VGND.t1248 852.769
R731 VGND.n2512 VGND.t2394 852.769
R732 VGND.n2537 VGND.t19 852.769
R733 VGND.n2538 VGND.t492 852.769
R734 VGND.n2563 VGND.t2319 852.769
R735 VGND.n2564 VGND.t1244 852.769
R736 VGND.n2589 VGND.t1514 852.769
R737 VGND.n2595 VGND.t188 852.769
R738 VGND.t1485 VGND.n2594 852.769
R739 VGND.n2634 VGND.t1906 852.769
R740 VGND.n2635 VGND.t20 852.769
R741 VGND.t21 VGND.n548 852.769
R742 VGND.n692 VGND.t1951 852.769
R743 VGND.n697 VGND.t1708 852.769
R744 VGND.n702 VGND.t1480 852.769
R745 VGND.n707 VGND.t1577 852.769
R746 VGND.n712 VGND.t2016 852.769
R747 VGND.n717 VGND.t366 852.769
R748 VGND.n722 VGND.t978 852.769
R749 VGND.n727 VGND.t2304 852.769
R750 VGND.n732 VGND.t1479 852.769
R751 VGND.n737 VGND.t31 852.769
R752 VGND.n742 VGND.t554 852.769
R753 VGND.n747 VGND.t352 852.769
R754 VGND.n2419 VGND.t1576 852.769
R755 VGND.t1709 VGND.n2418 852.769
R756 VGND.t2561 VGND.n2413 852.769
R757 VGND.t721 VGND.n549 852.769
R758 VGND.n2229 VGND.t1707 852.769
R759 VGND.n2254 VGND.t1281 852.769
R760 VGND.n2255 VGND.t1822 852.769
R761 VGND.n2280 VGND.t592 852.769
R762 VGND.n2281 VGND.t1482 852.769
R763 VGND.n2306 VGND.t974 852.769
R764 VGND.n2307 VGND.t1725 852.769
R765 VGND.n2332 VGND.t1954 852.769
R766 VGND.n2333 VGND.t714 852.769
R767 VGND.n2358 VGND.t1713 852.769
R768 VGND.n2359 VGND.t32 852.769
R769 VGND.n2389 VGND.t880 852.769
R770 VGND.n2394 VGND.t1907 852.769
R771 VGND.n2399 VGND.t350 852.769
R772 VGND.n2400 VGND.t1683 852.769
R773 VGND.t980 VGND.n550 852.769
R774 VGND.n2241 VGND.t2293 852.769
R775 VGND.n2242 VGND.t1854 852.769
R776 VGND.n2267 VGND.t1242 852.769
R777 VGND.n2268 VGND.t368 852.769
R778 VGND.n2293 VGND.t1659 852.769
R779 VGND.n2294 VGND.t1504 852.769
R780 VGND.n2319 VGND.t170 852.769
R781 VGND.n2320 VGND.t185 852.769
R782 VGND.n2345 VGND.t1581 852.769
R783 VGND.n2346 VGND.t1640 852.769
R784 VGND.n2371 VGND.t351 852.769
R785 VGND.n2377 VGND.t29 852.769
R786 VGND.t1805 VGND.n2376 852.769
R787 VGND.n2659 VGND.t45 852.769
R788 VGND.n2660 VGND.t1261 852.769
R789 VGND.t33 VGND.n551 852.769
R790 VGND.t881 VGND.n2156 852.769
R791 VGND.n869 VGND.t73 852.769
R792 VGND.n874 VGND.t2565 852.769
R793 VGND.n879 VGND.t780 852.769
R794 VGND.n884 VGND.t1300 852.769
R795 VGND.n889 VGND.t2687 852.769
R796 VGND.n894 VGND.t1623 852.769
R797 VGND.n899 VGND.t2027 852.769
R798 VGND.n904 VGND.t1823 852.769
R799 VGND.n909 VGND.t179 852.769
R800 VGND.n914 VGND.t1923 852.769
R801 VGND.n919 VGND.t2432 852.769
R802 VGND.n2137 VGND.t1921 852.769
R803 VGND.t835 VGND.n2136 852.769
R804 VGND.t951 VGND.n2131 852.769
R805 VGND.t74 VGND.n552 852.769
R806 VGND.n1947 VGND.t169 852.769
R807 VGND.n1972 VGND.t1584 852.769
R808 VGND.n1973 VGND.t187 852.769
R809 VGND.n1998 VGND.t839 852.769
R810 VGND.n1999 VGND.t911 852.769
R811 VGND.n2024 VGND.t2382 852.769
R812 VGND.n2025 VGND.t171 852.769
R813 VGND.n2050 VGND.t2410 852.769
R814 VGND.n2051 VGND.t1911 852.769
R815 VGND.n2076 VGND.t1579 852.769
R816 VGND.n2077 VGND.t2411 852.769
R817 VGND.n2107 VGND.t222 852.769
R818 VGND.n2112 VGND.t2560 852.769
R819 VGND.n2117 VGND.t2436 852.769
R820 VGND.n2118 VGND.t779 852.769
R821 VGND.t1820 VGND.n553 852.769
R822 VGND.n1959 VGND.t765 852.769
R823 VGND.n1960 VGND.t1842 852.769
R824 VGND.n1985 VGND.t975 852.769
R825 VGND.n1986 VGND.t2615 852.769
R826 VGND.n2011 VGND.t418 852.769
R827 VGND.n2012 VGND.t713 852.769
R828 VGND.n2037 VGND.t1512 852.769
R829 VGND.n2038 VGND.t1580 852.769
R830 VGND.n2063 VGND.t723 852.769
R831 VGND.n2064 VGND.t1660 852.769
R832 VGND.n2089 VGND.t1924 852.769
R833 VGND.n2095 VGND.t1638 852.769
R834 VGND.t2412 VGND.n2094 852.769
R835 VGND.n2684 VGND.t1510 852.769
R836 VGND.n2685 VGND.t2563 852.769
R837 VGND.t910 VGND.n554 852.769
R838 VGND.t2366 VGND.n1686 852.769
R839 VGND.t168 VGND.n1681 852.769
R840 VGND.t1163 VGND.n1676 852.769
R841 VGND.t2562 VGND.n1671 852.769
R842 VGND.t42 VGND.n1666 852.769
R843 VGND.t2480 VGND.n1661 852.769
R844 VGND.t1639 VGND.n1656 852.769
R845 VGND.t2030 VGND.n1651 852.769
R846 VGND.t2393 VGND.n1646 852.769
R847 VGND.t1815 VGND.n1641 852.769
R848 VGND.t1843 VGND.n1636 852.769
R849 VGND.t722 VGND.n1631 852.769
R850 VGND.n1910 VGND.t2415 852.769
R851 VGND.t841 VGND.n1909 852.769
R852 VGND.t2614 VGND.n1904 852.769
R853 VGND.t1513 VGND.n555 852.769
R854 VGND.n1720 VGND.t2 852.769
R855 VGND.n1745 VGND.t1583 852.769
R856 VGND.n1746 VGND.t1509 852.769
R857 VGND.n1771 VGND.t1841 852.769
R858 VGND.n1772 VGND.t27 852.769
R859 VGND.n1797 VGND.t698 852.769
R860 VGND.n1798 VGND.t2338 852.769
R861 VGND.n1823 VGND.t909 852.769
R862 VGND.n1824 VGND.t1308 852.769
R863 VGND.n1849 VGND.t104 852.769
R864 VGND.n1850 VGND.t599 852.769
R865 VGND.n1880 VGND.t1664 852.769
R866 VGND.n1885 VGND.t1681 852.769
R867 VGND.n1890 VGND.t766 852.769
R868 VGND.n1891 VGND.t160 852.769
R869 VGND.t1506 VGND.n556 852.769
R870 VGND.n1732 VGND.t22 852.769
R871 VGND.n1733 VGND.t49 852.769
R872 VGND.n1758 VGND.t2317 852.769
R873 VGND.n1759 VGND.t827 852.769
R874 VGND.n1784 VGND.t1658 852.769
R875 VGND.n1785 VGND.t0 852.769
R876 VGND.n1810 VGND.t1582 852.769
R877 VGND.n1811 VGND.t638 852.769
R878 VGND.n1836 VGND.t369 852.769
R879 VGND.n1837 VGND.t2585 852.769
R880 VGND.n1862 VGND.t1821 852.769
R881 VGND.n1868 VGND.t2433 852.769
R882 VGND.t1240 VGND.n1867 852.769
R883 VGND.n2709 VGND.t225 852.769
R884 VGND.n2710 VGND.t28 852.769
R885 VGND.t1803 VGND.n557 852.769
R886 VGND.t1496 VGND.n1317 852.769
R887 VGND.n1234 VGND.t1624 852.769
R888 VGND.n1239 VGND.t1515 852.769
R889 VGND.n1244 VGND.t1578 852.769
R890 VGND.n1249 VGND.t553 852.769
R891 VGND.n1254 VGND.t639 852.769
R892 VGND.n1259 VGND.t2028 852.769
R893 VGND.n1264 VGND.t1953 852.769
R894 VGND.n1269 VGND.t1959 852.769
R895 VGND.n1274 VGND.t1922 852.769
R896 VGND.n1279 VGND.t1597 852.769
R897 VGND.n1284 VGND.t166 852.769
R898 VGND.n1298 VGND.t190 852.769
R899 VGND.t699 VGND.n1297 852.769
R900 VGND.t697 VGND.n1292 852.769
R901 VGND.t1819 VGND.n558 852.769
R902 VGND.t2292 VGND.n296 852.769
R903 VGND.t826 VGND.n291 852.769
R904 VGND.t2596 VGND.n286 852.769
R905 VGND.t773 VGND.n281 852.769
R906 VGND.t1853 VGND.n276 852.769
R907 VGND.t1138 VGND.n271 852.769
R908 VGND.t1307 VGND.n266 852.769
R909 VGND.t1508 VGND.n261 852.769
R910 VGND.t18 VGND.n256 852.769
R911 VGND.t1682 VGND.n251 852.769
R912 VGND.t2584 VGND.n246 852.769
R913 VGND.t2318 VGND.n241 852.769
R914 VGND.t1667 VGND.n236 852.769
R915 VGND.t1497 VGND.n231 852.769
R916 VGND.t2314 VGND.n226 852.769
R917 VGND.n3010 VGND.t1301 852.769
R918 VGND.n1330 VGND.t2597 852.769
R919 VGND.n1396 VGND.t2414 852.769
R920 VGND.t239 VGND.n1395 852.769
R921 VGND.t1507 VGND.n1390 852.769
R922 VGND.t712 VGND.n1385 852.769
R923 VGND.t491 VGND.n1380 852.769
R924 VGND.t2383 VGND.n1375 852.769
R925 VGND.t1802 VGND.n1370 852.769
R926 VGND.t2413 VGND.n1365 852.769
R927 VGND.t224 VGND.n1360 852.769
R928 VGND.t774 VGND.n1355 852.769
R929 VGND.t1282 VGND.n1350 852.769
R930 VGND.t1243 VGND.n1345 852.769
R931 VGND.t1817 VGND.n1340 852.769
R932 VGND.t2294 VGND.n1335 852.769
R933 VGND.n2740 VGND.t715 852.769
R934 VGND.n2226 VGND 851.341
R935 VGND.n1319 VGND.t1067 809.773
R936 VGND.t1399 VGND.n2924 809.773
R937 VGND.n2848 VGND.t1115 809.773
R938 VGND.n2849 VGND.t1022 809.773
R939 VGND.t1064 VGND.n521 809.773
R940 VGND.t1136 VGND.n687 809.773
R941 VGND.n806 VGND.t1016 809.773
R942 VGND.n2157 VGND.t1058 809.773
R943 VGND.t1070 VGND.n841 809.773
R944 VGND.n1718 VGND.t1094 809.773
R945 VGND.t1025 VGND.n1719 809.773
R946 VGND.n1051 VGND.t1097 809.773
R947 VGND.n1318 VGND.t1127 809.773
R948 VGND.n297 VGND.t1040 809.773
R949 VGND.t1344 VGND.n1321 809.773
R950 VGND.t664 VGND.t516 708.047
R951 VGND.t666 VGND.t664 708.047
R952 VGND.t656 VGND.t666 708.047
R953 VGND.t59 VGND.t656 708.047
R954 VGND.t56 VGND.t59 708.047
R955 VGND.t62 VGND.t56 708.047
R956 VGND.t53 VGND.t62 708.047
R957 VGND.t50 VGND.t1233 708.047
R958 VGND.t584 VGND.t582 708.047
R959 VGND.t679 VGND.t584 708.047
R960 VGND.t551 VGND.t679 708.047
R961 VGND.t704 VGND.t551 708.047
R962 VGND.t701 VGND.t704 708.047
R963 VGND.t707 VGND.t701 708.047
R964 VGND.t710 VGND.t707 708.047
R965 VGND.t518 VGND.t576 708.047
R966 VGND.t731 VGND.t518 708.047
R967 VGND.t683 VGND.t731 708.047
R968 VGND.t1259 VGND.t683 708.047
R969 VGND.t1255 VGND.t1259 708.047
R970 VGND.t1249 VGND.t1255 708.047
R971 VGND.t1251 VGND.t1249 708.047
R972 VGND.t51 VGND.t1230 708.047
R973 VGND.t724 VGND.t520 708.047
R974 VGND.t686 VGND.t724 708.047
R975 VGND.t586 VGND.t686 708.047
R976 VGND.t55 VGND.t586 708.047
R977 VGND.t61 VGND.t55 708.047
R978 VGND.t58 VGND.t61 708.047
R979 VGND.t64 VGND.t58 708.047
R980 VGND.t524 VGND.t574 708.047
R981 VGND.t574 VGND.t514 708.047
R982 VGND.t514 VGND.t588 708.047
R983 VGND.t588 VGND.t700 708.047
R984 VGND.t700 VGND.t706 708.047
R985 VGND.t706 VGND.t703 708.047
R986 VGND.t703 VGND.t709 708.047
R987 VGND.t658 VGND.t726 708.047
R988 VGND.t580 VGND.t658 708.047
R989 VGND.t733 VGND.t580 708.047
R990 VGND.t1257 VGND.t733 708.047
R991 VGND.t1253 VGND.t1257 708.047
R992 VGND.t1258 VGND.t1253 708.047
R993 VGND.t1254 VGND.t1258 708.047
R994 VGND.n127 VGND.n126 708.047
R995 VGND.t761 VGND.t2031 691.188
R996 VGND.t837 VGND.t2526 691.188
R997 VGND.n458 VGND.n297 660.87
R998 VGND.t483 VGND.t1590 657.471
R999 VGND.t1772 VGND.t1588 657.471
R1000 VGND.t2521 VGND.t1586 657.471
R1001 VGND.t673 VGND.t1781 657.471
R1002 VGND.t2568 VGND.t737 657.471
R1003 VGND.t1845 VGND.t236 657.471
R1004 VGND.t578 VGND.t232 657.471
R1005 VGND.t749 VGND.t226 657.471
R1006 VGND.t1781 VGND.t1714 654.197
R1007 VGND.t737 VGND.t590 654.197
R1008 VGND.n2159 VGND 640.614
R1009 VGND.n451 VGND 640.614
R1010 VGND.n422 VGND 640.614
R1011 VGND.n391 VGND 640.614
R1012 VGND.n358 VGND 632.184
R1013 VGND.t527 VGND.t2510 630.62
R1014 VGND.t1502 VGND.t572 630.62
R1015 VGND.t66 VGND.t118 630.62
R1016 VGND.t2516 VGND.t1313 630.62
R1017 VGND.t2508 VGND.t2299 630.62
R1018 VGND.t568 VGND.t2424 630.62
R1019 VGND.t566 VGND.t843 630.62
R1020 VGND.t2506 VGND.t1642 630.62
R1021 VGND.t2504 VGND.t767 630.62
R1022 VGND.t570 VGND.t555 630.62
R1023 VGND.t2514 VGND.t1494 630.62
R1024 VGND.t2512 VGND.t1706 630.62
R1025 VGND.t564 VGND.t1940 630.62
R1026 VGND.t122 VGND.t23 630.62
R1027 VGND.t907 VGND.t120 630.62
R1028 VGND.t1483 VGND.t294 630.62
R1029 VGND.t311 VGND.t1321 630.62
R1030 VGND.t307 VGND.t1411 630.62
R1031 VGND.t1398 VGND.t1403 630.62
R1032 VGND.t1383 VGND.t1562 630.62
R1033 VGND.t303 VGND.t504 630.62
R1034 VGND.t285 VGND.t1385 630.62
R1035 VGND.t506 VGND.t271 630.62
R1036 VGND.t500 VGND.t1550 630.62
R1037 VGND.t273 VGND.t1546 630.62
R1038 VGND.t287 VGND.t1386 630.62
R1039 VGND.t1548 VGND.t1366 630.62
R1040 VGND.t1351 VGND.t1538 630.62
R1041 VGND.t264 VGND.t269 630.62
R1042 VGND.t257 VGND.t1355 630.62
R1043 VGND.t1332 VGND.t241 630.62
R1044 VGND.t1531 VGND.t261 630.62
R1045 VGND.t1791 VGND.t1605 630.62
R1046 VGND.t2133 VGND.t2378 630.62
R1047 VGND.t2588 VGND.t2341 630.62
R1048 VGND.t1420 VGND.t2339 630.62
R1049 VGND.t1751 VGND.t1789 630.62
R1050 VGND.t2268 VGND.t2374 630.62
R1051 VGND.t2490 VGND.t2372 630.62
R1052 VGND.t895 VGND.t1787 630.62
R1053 VGND.t2022 VGND.t1785 630.62
R1054 VGND.t2580 VGND.t2376 630.62
R1055 VGND.t463 VGND.t2357 630.62
R1056 VGND.t2088 VGND.t2355 630.62
R1057 VGND.t410 VGND.t2370 630.62
R1058 VGND.t2301 VGND.t2368 630.62
R1059 VGND.t991 VGND.t2343 630.62
R1060 VGND.t1370 VGND.t1783 630.62
R1061 VGND.t2291 VGND.t1835 630.62
R1062 VGND.t2150 VGND.t541 630.62
R1063 VGND.t853 VGND.t2275 630.62
R1064 VGND.t2273 VGND.t2404 630.62
R1065 VGND.t886 VGND.t1833 630.62
R1066 VGND.t2266 VGND.t2557 630.62
R1067 VGND.t112 VGND.t2264 630.62
R1068 VGND.t1831 VGND.t2313 630.62
R1069 VGND.t2038 VGND.t2154 630.62
R1070 VGND.t2148 VGND.t622 630.62
R1071 VGND.t1493 VGND.t1839 630.62
R1072 VGND.t1837 VGND.t2478 630.62
R1073 VGND.t916 VGND.t2262 630.62
R1074 VGND.t1830 VGND.t1806 630.62
R1075 VGND.t2323 VGND.t2277 630.62
R1076 VGND.t2152 VGND.t1560 630.62
R1077 VGND.t528 VGND.t1765 630.62
R1078 VGND.t1808 VGND.t154 630.62
R1079 VGND.t1633 VGND.t65 630.62
R1080 VGND.t1315 VGND.t1631 630.62
R1081 VGND.t1763 VGND.t2345 630.62
R1082 VGND.t2425 VGND.t150 630.62
R1083 VGND.t148 VGND.t845 630.62
R1084 VGND.t1644 VGND.t1761 630.62
R1085 VGND.t1759 VGND.t769 630.62
R1086 VGND.t557 VGND.t152 630.62
R1087 VGND.t1629 VGND.t1898 630.62
R1088 VGND.t1702 VGND.t1767 630.62
R1089 VGND.t146 VGND.t429 630.62
R1090 VGND.t144 VGND.t25 630.62
R1091 VGND.t908 VGND.t1635 630.62
R1092 VGND.t2380 VGND.t302 630.62
R1093 VGND.t1599 VGND.t1677 630.62
R1094 VGND.t829 VGND.t347 630.62
R1095 VGND.t798 VGND.t640 630.62
R1096 VGND.t1572 VGND.t1613 630.62
R1097 VGND.t2257 VGND.t1675 630.62
R1098 VGND.t1711 VGND.t343 630.62
R1099 VGND.t2484 VGND.t341 630.62
R1100 VGND.t76 VGND.t1673 630.62
R1101 VGND.t1680 VGND.t1671 630.62
R1102 VGND.t2012 VGND.t345 630.62
R1103 VGND.t377 VGND.t1611 630.62
R1104 VGND.t129 VGND.t1609 630.62
R1105 VGND.t404 VGND.t339 630.62
R1106 VGND.t337 VGND.t1998 630.62
R1107 VGND.t642 VGND.t985 630.62
R1108 VGND.t1669 VGND.t1342 630.62
R1109 VGND.t2288 VGND.t654 630.62
R1110 VGND.t644 VGND.t2682 630.62
R1111 VGND.t852 VGND.t2194 630.62
R1112 VGND.t2192 VGND.t2397 630.62
R1113 VGND.t2279 VGND.t652 630.62
R1114 VGND.t2212 VGND.t2554 630.62
R1115 VGND.t851 VGND.t2210 630.62
R1116 VGND.t650 VGND.t2306 630.62
R1117 VGND.t984 VGND.t648 630.62
R1118 VGND.t2214 VGND.t563 630.62
R1119 VGND.t1490 VGND.t2190 630.62
R1120 VGND.t2188 VGND.t1995 630.62
R1121 VGND.t435 VGND.t2200 630.62
R1122 VGND.t2472 VGND.t2198 630.62
R1123 VGND.t1893 VGND.t2196 630.62
R1124 VGND.t646 VGND.t1537 630.62
R1125 VGND.t630 VGND.t534 630.62
R1126 VGND.t542 VGND.t608 630.62
R1127 VGND.t739 VGND.t795 630.62
R1128 VGND.t2405 VGND.t636 630.62
R1129 VGND.t628 VGND.t887 630.62
R1130 VGND.t2558 VGND.t604 630.62
R1131 VGND.t602 VGND.t113 630.62
R1132 VGND.t1564 VGND.t626 630.62
R1133 VGND.t624 VGND.t1925 630.62
R1134 VGND.t623 VGND.t606 630.62
R1135 VGND.t634 VGND.t1897 630.62
R1136 VGND.t2479 VGND.t632 630.62
R1137 VGND.t600 VGND.t1988 630.62
R1138 VGND.t743 VGND.t2147 630.62
R1139 VGND.t2324 VGND.t741 630.62
R1140 VGND.t610 VGND.t1563 630.62
R1141 VGND.t971 VGND.t529 630.62
R1142 VGND.t1809 VGND.t597 630.62
R1143 VGND.t68 VGND.t1621 630.62
R1144 VGND.t1316 VGND.t1619 630.62
R1145 VGND.t2346 VGND.t969 630.62
R1146 VGND.t752 VGND.t593 630.62
R1147 VGND.t846 VGND.t878 630.62
R1148 VGND.t1645 VGND.t967 630.62
R1149 VGND.t770 VGND.t158 630.62
R1150 VGND.t558 VGND.t595 630.62
R1151 VGND.t1899 VGND.t1617 630.62
R1152 VGND.t1703 VGND.t1615 630.62
R1153 VGND.t430 VGND.t876 630.62
R1154 VGND.t874 VGND.t26 630.62
R1155 VGND.t872 VGND.t1884 630.62
R1156 VGND.t156 VGND.t304 630.62
R1157 VGND.t526 VGND.t1468 630.62
R1158 VGND.t2184 VGND.t1503 630.62
R1159 VGND.t67 VGND.t922 630.62
R1160 VGND.t920 VGND.t1314 630.62
R1161 VGND.t2298 VGND.t1466 630.62
R1162 VGND.t2180 VGND.t2423 630.62
R1163 VGND.t844 VGND.t38 630.62
R1164 VGND.t1464 VGND.t1643 630.62
R1165 VGND.t768 VGND.t1661 630.62
R1166 VGND.t2182 VGND.t556 630.62
R1167 VGND.t1495 VGND.t918 630.62
R1168 VGND.t1470 VGND.t1701 630.62
R1169 VGND.t1941 VGND.t36 630.62
R1170 VGND.t24 VGND.t34 630.62
R1171 VGND.t906 VGND.t924 630.62
R1172 VGND.t2186 VGND.t295 630.62
R1173 VGND.t871 VGND.t2230 630.62
R1174 VGND.t828 VGND.t2220 630.62
R1175 VGND.t1918 VGND.t801 630.62
R1176 VGND.t1571 VGND.t1916 630.62
R1177 VGND.t2228 VGND.t2256 630.62
R1178 VGND.t1710 VGND.t2216 630.62
R1179 VGND.t1690 VGND.t2483 630.62
R1180 VGND.t75 VGND.t2226 630.62
R1181 VGND.t2224 VGND.t1679 630.62
R1182 VGND.t2009 VGND.t2218 630.62
R1183 VGND.t1914 VGND.t376 630.62
R1184 VGND.t126 VGND.t1912 630.62
R1185 VGND.t1688 VGND.t403 630.62
R1186 VGND.t1686 VGND.t175 630.62
R1187 VGND.t2331 VGND.t1684 630.62
R1188 VGND.t2222 VGND.t1337 630.62
R1189 VGND.t783 VGND.t2283 630.62
R1190 VGND.t2100 VGND.t2144 630.62
R1191 VGND.t791 VGND.t1473 630.62
R1192 VGND.t789 VGND.t2392 630.62
R1193 VGND.t781 VGND.t357 630.62
R1194 VGND.t2096 VGND.t365 630.62
R1195 VGND.t2094 VGND.t864 630.62
R1196 VGND.t2106 VGND.t3 630.62
R1197 VGND.t2104 VGND.t180 630.62
R1198 VGND.t2098 VGND.t696 630.62
R1199 VGND.t787 VGND.t2066 630.62
R1200 VGND.t785 VGND.t2471 630.62
R1201 VGND.t2092 VGND.t1935 630.62
R1202 VGND.t2090 VGND.t15 630.62
R1203 VGND.t793 VGND.t901 630.62
R1204 VGND.t2102 VGND.t254 630.62
R1205 VGND.t2290 VGND.t1656 630.62
R1206 VGND.t1646 VGND.t2684 630.62
R1207 VGND.t854 VGND.t1294 630.62
R1208 VGND.t1292 VGND.t2403 630.62
R1209 VGND.t2281 VGND.t1654 630.62
R1210 VGND.t2441 VGND.t2556 630.62
R1211 VGND.t107 VGND.t2439 630.62
R1212 VGND.t1652 VGND.t2308 630.62
R1213 VGND.t2033 VGND.t1650 630.62
R1214 VGND.t2443 VGND.t621 630.62
R1215 VGND.t1492 VGND.t1290 630.62
R1216 VGND.t1288 VGND.t1700 630.62
R1217 VGND.t437 VGND.t2437 630.62
R1218 VGND.t1829 VGND.t370 630.62
R1219 VGND.t2322 VGND.t1296 630.62
R1220 VGND.t1648 VGND.t1557 630.62
R1221 VGND.t2656 VGND.t2282 630.62
R1222 VGND.t2143 VGND.t2626 630.62
R1223 VGND.t425 VGND.t1476 630.62
R1224 VGND.t2391 VGND.t423 630.62
R1225 VGND.t2430 VGND.t356 630.62
R1226 VGND.t364 VGND.t2622 630.62
R1227 VGND.t2620 VGND.t2388 630.62
R1228 VGND.t165 VGND.t2428 630.62
R1229 VGND.t2426 VGND.t1274 630.62
R1230 VGND.t693 VGND.t2624 630.62
R1231 VGND.t421 VGND.t2065 630.62
R1232 VGND.t2075 VGND.t419 630.62
R1233 VGND.t2618 VGND.t1934 630.62
R1234 VGND.t2616 VGND.t12 630.62
R1235 VGND.t900 VGND.t427 630.62
R1236 VGND.t2628 VGND.t251 630.62
R1237 VGND.t142 VGND.t1604 630.62
R1238 VGND.t2132 VGND.t132 630.62
R1239 VGND.t2595 VGND.t2598 630.62
R1240 VGND.t1419 VGND.t195 630.62
R1241 VGND.t1750 VGND.t140 630.62
R1242 VGND.t1712 VGND.t2608 630.62
R1243 VGND.t2489 VGND.t2606 630.62
R1244 VGND.t894 VGND.t138 630.62
R1245 VGND.t2021 VGND.t136 630.62
R1246 VGND.t2013 VGND.t130 630.62
R1247 VGND.t462 VGND.t193 630.62
R1248 VGND.t2081 VGND.t191 630.62
R1249 VGND.t409 VGND.t2604 630.62
R1250 VGND.t2602 VGND.t1999 630.62
R1251 VGND.t2600 VGND.t990 630.62
R1252 VGND.t134 VGND.t1357 630.62
R1253 VGND.t1199 VGND.t2289 630.62
R1254 VGND.t2630 VGND.t2683 630.62
R1255 VGND.t1430 VGND.t863 630.62
R1256 VGND.t1428 VGND.t2398 630.62
R1257 VGND.t1197 VGND.t2280 630.62
R1258 VGND.t1955 VGND.t2555 630.62
R1259 VGND.t1438 VGND.t106 630.62
R1260 VGND.t1195 VGND.t2307 630.62
R1261 VGND.t1193 VGND.t2688 630.62
R1262 VGND.t1957 VGND.t612 630.62
R1263 VGND.t1426 VGND.t1491 630.62
R1264 VGND.t1201 VGND.t1996 630.62
R1265 VGND.t1436 VGND.t436 630.62
R1266 VGND.t1434 VGND.t2473 630.62
R1267 VGND.t1432 VGND.t1894 630.62
R1268 VGND.t1191 VGND.t1539 630.62
R1269 VGND.t1306 VGND.t333 630.62
R1270 VGND.t2140 VGND.t252 630.62
R1271 VGND.t1347 VGND.t1472 630.62
R1272 VGND.t1325 VGND.t1423 630.62
R1273 VGND.t322 VGND.t1758 630.62
R1274 VGND.t1407 VGND.t2502 630.62
R1275 VGND.t1396 VGND.t2497 630.62
R1276 VGND.t318 VGND.t1268 630.62
R1277 VGND.t300 VGND.t1279 630.62
R1278 VGND.t1409 VGND.t2581 630.62
R1279 VGND.t502 VGND.t472 630.62
R1280 VGND.t1558 VGND.t2076 630.62
R1281 VGND.t1391 VGND.t417 630.62
R1282 VGND.t1378 VGND.t2302 630.62
R1283 VGND.t1353 VGND.t994 630.62
R1284 VGND.t279 VGND.t1382 630.62
R1285 VGND.n2187 VGND.n2159 599.125
R1286 VGND.n451 VGND.n450 599.125
R1287 VGND.n422 VGND.n421 599.125
R1288 VGND.n391 VGND.n390 599.125
R1289 VGND.n358 VGND.n357 599.125
R1290 VGND.n2877 VGND.n2876 599.125
R1291 VGND.n128 VGND.n127 599.125
R1292 VGND.n2916 VGND.n2915 599.125
R1293 VGND VGND.t869 581.61
R1294 VGND VGND.t53 573.181
R1295 VGND VGND.t710 573.181
R1296 VGND VGND.t1251 573.181
R1297 VGND VGND.t228 573.181
R1298 VGND VGND.t2528 564.751
R1299 VGND.n2873 VGND 564.751
R1300 VGND VGND.n2875 564.751
R1301 VGND.n2874 VGND 556.322
R1302 VGND VGND.t959 539.465
R1303 VGND.t976 VGND 539.465
R1304 VGND.n1626 VGND.t487 494.779
R1305 VGND.n2861 VGND.n2851 494.253
R1306 VGND.n1567 VGND.t1374 492.058
R1307 VGND.n1566 VGND.t1553 492.058
R1308 VGND.t1529 VGND.n1411 492.058
R1309 VGND.t1372 VGND.n1423 492.058
R1310 VGND.n1424 VGND.t1360 492.058
R1311 VGND.t1338 VGND.n1442 492.058
R1312 VGND.n1443 VGND.t265 492.058
R1313 VGND.t245 VGND.n1455 492.058
R1314 VGND.n1456 VGND.t1333 492.058
R1315 VGND.t320 VGND.n1474 492.058
R1316 VGND.n1475 VGND.t309 492.058
R1317 VGND.t1394 VGND.n1487 492.058
R1318 VGND.n1488 VGND.t1323 492.058
R1319 VGND.t298 VGND.n1506 492.058
R1320 VGND.n1507 VGND.t1405 492.058
R1321 VGND.t1714 VGND.t2361 481.877
R1322 VGND.t2361 VGND.t511 481.877
R1323 VGND.t1848 VGND.t662 481.877
R1324 VGND.t590 VGND.t1848 481.877
R1325 VGND.t1498 VGND 452.382
R1326 VGND.n1567 VGND.t966 424.312
R1327 VGND.t2295 VGND.n1566 424.312
R1328 VGND.n1411 VGND.t1961 424.312
R1329 VGND.n1423 VGND.t349 424.312
R1330 VGND.n1424 VGND.t41 424.312
R1331 VGND.n1442 VGND.t367 424.312
R1332 VGND.n1443 VGND.t2503 424.312
R1333 VGND.n1455 VGND.t1852 424.312
R1334 VGND.n1456 VGND.t2006 424.312
R1335 VGND.n1474 VGND.t189 424.312
R1336 VGND.n1475 VGND.t494 424.312
R1337 VGND.n1487 VGND.t2416 424.312
R1338 VGND.n1488 VGND.t1960 424.312
R1339 VGND.n1506 VGND.t47 424.312
R1340 VGND.n1507 VGND.t981 424.312
R1341 VGND.t2587 VGND.n560 424.312
R1342 VGND.t1283 VGND 419.68
R1343 VGND.n687 VGND.n491 413.043
R1344 VGND.t213 VGND.t1067 408.469
R1345 VGND.t2166 VGND.t532 408.469
R1346 VGND.t395 VGND.t539 408.469
R1347 VGND.t859 VGND.t2204 408.469
R1348 VGND.t1944 VGND.t446 408.469
R1349 VGND.t884 VGND.t1215 408.469
R1350 VGND.t2269 VGND.t96 408.469
R1351 VGND.t108 VGND.t2538 408.469
R1352 VGND.t2309 VGND.t2648 408.469
R1353 VGND.t2034 VGND.t1974 408.469
R1354 VGND.t613 VGND.t2254 408.469
R1355 VGND.t464 VGND.t2636 408.469
R1356 VGND.t1692 VGND.t1964 408.469
R1357 VGND.t912 VGND.t1177 408.469
R1358 VGND.t1151 VGND.t2476 408.469
R1359 VGND.t1885 VGND.t2662 408.469
R1360 VGND.t1052 VGND.t1399 408.469
R1361 VGND.t509 VGND.t1001 408.469
R1362 VGND.t1007 VGND.t305 408.469
R1363 VGND.t283 VGND.t1013 408.469
R1364 VGND.t1100 VGND.t507 408.469
R1365 VGND.t496 VGND.t1106 408.469
R1366 VGND.t1019 VGND.t1544 408.469
R1367 VGND.t1387 VGND.t1061 408.469
R1368 VGND.t1076 VGND.t1364 408.469
R1369 VGND.t1540 VGND.t1112 408.469
R1370 VGND.t1034 VGND.t267 408.469
R1371 VGND.t255 VGND.t1079 408.469
R1372 VGND.t1118 VGND.t1335 408.469
R1373 VGND.t1527 VGND.t1130 408.469
R1374 VGND.t1046 VGND.t243 408.469
R1375 VGND.t1349 VGND.t1088 408.469
R1376 VGND.t1115 VGND.t454 408.469
R1377 VGND.t1139 VGND.t2286 408.469
R1378 VGND.t211 VGND.t1500 408.469
R1379 VGND.t2061 VGND.t1474 408.469
R1380 VGND.t393 VGND.t1424 408.469
R1381 VGND.t2202 VGND.t2296 408.469
R1382 VGND.t2057 VGND.t759 408.469
R1383 VGND.t1872 VGND.t867 408.469
R1384 VGND.t1982 VGND.t6 408.469
R1385 VGND.t82 VGND.t183 408.469
R1386 VGND.t2644 VGND.t694 408.469
R1387 VGND.t1968 VGND.t1488 408.469
R1388 VGND.t2248 VGND.t2469 408.469
R1389 VGND.t2122 VGND.t1938 408.469
R1390 VGND.t1448 VGND.t13 408.469
R1391 VGND.t1173 VGND.t995 408.469
R1392 VGND.t2674 VGND.t1022 408.469
R1393 VGND.t1302 VGND.t2240 408.469
R1394 VGND.t2114 VGND.t2136 408.469
R1395 VGND.t2591 VGND.t1740 408.469
R1396 VGND.t947 VGND.t2408 408.469
R1397 VGND.t1754 VGND.t2160 408.469
R1398 VGND.t1728 VGND.t2419 408.469
R1399 VGND.t2493 VGND.t2467 408.469
R1400 VGND.t438 VGND.t1264 408.469
R1401 VGND.t2025 VGND.t379 408.469
R1402 VGND.t2548 VGND.t2576 408.469
R1403 VGND.t2069 VGND.t1878 408.469
R1404 VGND.t818 VGND.t2084 408.469
R1405 VGND.t2208 VGND.t413 408.469
R1406 VGND.t2652 VGND.t2002 408.469
R1407 VGND.t2327 VGND.t1221 408.469
R1408 VGND.t1976 VGND.t1064 408.469
R1409 VGND.t2045 VGND.t535 408.469
R1410 VGND.t543 VGND.t2638 408.469
R1411 VGND.t1454 VGND.t857 408.469
R1412 VGND.t1946 VGND.t2242 408.469
R1413 VGND.t1153 VGND.t888 408.469
R1414 VGND.t2498 VGND.t1440 408.469
R1415 VGND.t949 VGND.t114 408.469
R1416 VGND.t1565 VGND.t2162 408.469
R1417 VGND.t1730 VGND.t1926 408.469
R1418 VGND.t617 VGND.t458 408.469
R1419 VGND.t401 VGND.t468 408.469
R1420 VGND.t1696 VGND.t217 408.469
R1421 VGND.t1989 VGND.t2552 408.469
R1422 VGND.t1223 VGND.t1825 408.469
R1423 VGND.t1889 VGND.t822 408.469
R1424 VGND.t98 VGND.t1136 408.469
R1425 VGND.t1864 VGND.t1519 408.469
R1426 VGND.t1209 VGND.t2141 408.469
R1427 VGND.t1183 VGND.t896 408.469
R1428 VGND.t2047 VGND.t1417 408.469
R1429 VGND.t2670 VGND.t354 408.469
R1430 VGND.t1167 VGND.t755 408.469
R1431 VGND.t2244 VGND.t2386 408.469
R1432 VGND.t1157 VGND.t163 408.469
R1433 VGND.t1442 VGND.t1272 408.469
R1434 VGND.t2176 VGND.t689 408.469
R1435 VGND.t1145 VGND.t1902 408.469
R1436 VGND.t2465 VGND.t2079 408.469
R1437 VGND.t1932 VGND.t460 408.469
R1438 VGND.t8 VGND.t824 408.469
R1439 VGND.t988 VGND.t1726 408.469
R1440 VGND.t2534 VGND.t1043 408.469
R1441 VGND.t1600 VGND.t383 408.469
R1442 VGND.t804 VGND.t830 408.469
R1443 VGND.t796 VGND.t2250 408.469
R1444 VGND.t1860 VGND.t2399 408.469
R1445 VGND.t2258 VGND.t1189 408.469
R1446 VGND.t2236 VGND.t360 408.469
R1447 VGND.t2485 VGND.t2041 408.469
R1448 VGND.t2658 VGND.t890 408.469
R1449 VGND.t2017 VGND.t943 408.469
R1450 VGND.t1161 VGND.t2007 408.469
R1451 VGND.t1486 VGND.t1458 408.469
R1452 VGND.t939 VGND.t124 408.469
R1453 VGND.t2170 VGND.t405 408.469
R1454 VGND.t215 VGND.t173 408.469
R1455 VGND.t1895 VGND.t2459 408.469
R1456 VGND.t1016 VGND.t444 408.469
R1457 VGND.t1738 VGND.t1304 408.469
R1458 VGND.t2138 VGND.t199 408.469
R1459 VGND.t2051 VGND.t2589 408.469
R1460 VGND.t1569 VGND.t385 408.469
R1461 VGND.t90 VGND.t1756 408.469
R1462 VGND.t2421 VGND.t2043 408.469
R1463 VGND.t1862 VGND.t2495 408.469
R1464 VGND.t1266 VGND.t1966 408.469
R1465 VGND.t2238 VGND.t1277 408.469
R1466 VGND.t2578 VGND.t2632 408.469
R1467 VGND.t1185 VGND.t2518 408.469
R1468 VGND.t2086 VGND.t2234 408.469
R1469 VGND.t415 VGND.t2108 408.469
R1470 VGND.t2461 VGND.t2004 408.469
R1471 VGND.t2329 VGND.t941 408.469
R1472 VGND.t1058 VGND.t1462 408.469
R1473 VGND.t2128 VGND.t537 408.469
R1474 VGND.t1159 VGND.t545 408.469
R1475 VGND.t219 VGND.t855 408.469
R1476 VGND.t931 VGND.t1948 408.469
R1477 VGND.t397 VGND.t2389 408.469
R1478 VGND.t205 VGND.t2500 408.469
R1479 VGND.t2453 VGND.t116 408.469
R1480 VGND.t1876 VGND.t1567 408.469
R1481 VGND.t812 VGND.t1928 408.469
R1482 VGND.t2540 VGND.t619 408.469
R1483 VGND.t1866 VGND.t470 408.469
R1484 VGND.t806 VGND.t1698 408.469
R1485 VGND.t1991 VGND.t102 408.469
R1486 VGND.t1827 VGND.t2640 408.469
R1487 VGND.t1891 VGND.t1211 408.469
R1488 VGND.t1187 VGND.t1070 408.469
R1489 VGND.t530 VGND.t2654 408.469
R1490 VGND.t2680 VGND.t2685 408.469
R1491 VGND.t861 VGND.t2463 408.469
R1492 VGND.t2130 VGND.t1942 408.469
R1493 VGND.t882 VGND.t1141 408.469
R1494 VGND.t2455 VGND.t2271 408.469
R1495 VGND.t110 VGND.t933 408.469
R1496 VGND.t399 VGND.t2311 408.469
R1497 VGND.t2036 VGND.t209 408.469
R1498 VGND.t448 VGND.t615 408.469
R1499 VGND.t466 VGND.t389 408.469
R1500 VGND.t201 VGND.t1694 408.469
R1501 VGND.t2542 VGND.t914 408.469
R1502 VGND.t1213 VGND.t2474 408.469
R1503 VGND.t1887 VGND.t808 408.469
R1504 VGND.t88 VGND.t998 408.469
R1505 VGND.t1225 VGND.t1517 408.469
R1506 VGND.t1793 VGND.t1207 408.469
R1507 VGND.t945 VGND.t898 408.469
R1508 VGND.t1415 VGND.t2039 408.469
R1509 VGND.t1460 VGND.t2071 408.469
R1510 VGND.t753 VGND.t935 408.469
R1511 VGND.t2232 VGND.t2384 408.469
R1512 VGND.t161 VGND.t1143 408.469
R1513 VGND.t2457 VGND.t1270 408.469
R1514 VGND.t2582 VGND.t2168 408.469
R1515 VGND.t1746 VGND.t1900 408.469
R1516 VGND.t2077 VGND.t2451 408.469
R1517 VGND.t1930 VGND.t450 408.469
R1518 VGND.t810 VGND.t16 408.469
R1519 VGND.t986 VGND.t203 408.469
R1520 VGND.t1094 VGND.t452 408.469
R1521 VGND.t1523 VGND.t1744 408.469
R1522 VGND.t1812 VGND.t207 408.469
R1523 VGND.t69 VGND.t2059 408.469
R1524 VGND.t1311 VGND.t387 408.469
R1525 VGND.t2349 VGND.t100 408.469
R1526 VGND.t777 VGND.t2049 408.469
R1527 VGND.t849 VGND.t1868 408.469
R1528 VGND.t1319 VGND.t1978 408.469
R1529 VGND.t982 VGND.t2252 408.469
R1530 VGND.t561 VGND.t2642 408.469
R1531 VGND.t374 VGND.t1962 408.469
R1532 VGND.t1993 VGND.t2246 408.469
R1533 VGND.t433 VGND.t2116 408.469
R1534 VGND.t2612 VGND.t1444 408.469
R1535 VGND.t904 VGND.t1169 408.469
R1536 VGND.t86 VGND.t1025 408.469
R1537 VGND.t1606 VGND.t1217 408.469
R1538 VGND.t1203 VGND.t2134 408.469
R1539 VGND.t2593 VGND.t937 408.469
R1540 VGND.t2650 VGND.t2406 408.469
R1541 VGND.t1752 VGND.t1456 408.469
R1542 VGND.t929 VGND.t2417 408.469
R1543 VGND.t2491 VGND.t2126 408.469
R1544 VGND.t1748 VGND.t1262 408.469
R1545 VGND.t2023 VGND.t2449 408.469
R1546 VGND.t2164 VGND.t2014 408.469
R1547 VGND.t2067 VGND.t1742 408.469
R1548 VGND.t2447 VGND.t2082 408.469
R1549 VGND.t440 VGND.t411 408.469
R1550 VGND.t802 VGND.t2000 408.469
R1551 VGND.t2325 VGND.t197 408.469
R1552 VGND.t1097 VGND.t1219 408.469
R1553 VGND.t2532 VGND.t1521 408.469
R1554 VGND.t1810 VGND.t2055 408.469
R1555 VGND.t2678 VGND.t71 408.469
R1556 VGND.t1309 VGND.t92 408.469
R1557 VGND.t2120 VGND.t2347 408.469
R1558 VGND.t775 VGND.t2668 408.469
R1559 VGND.t1970 VGND.t847 408.469
R1560 VGND.t1317 VGND.t927 408.469
R1561 VGND.t1155 VGND.t771 408.469
R1562 VGND.t559 VGND.t1450 408.469
R1563 VGND.t2172 VGND.t372 408.469
R1564 VGND.t1704 VGND.t1147 408.469
R1565 VGND.t431 VGND.t1736 408.469
R1566 VGND.t1880 VGND.t2610 408.469
R1567 VGND.t902 VGND.t2156 408.469
R1568 VGND.t1127 VGND.t816 408.469
R1569 VGND.t442 VGND.t2284 408.469
R1570 VGND.t1874 VGND.t2145 408.469
R1571 VGND.t1984 VGND.t1477 408.469
R1572 VGND.t2536 VGND.t1421 408.469
R1573 VGND.t2646 VGND.t358 408.469
R1574 VGND.t1972 VGND.t757 408.469
R1575 VGND.t94 VGND.t865 408.469
R1576 VGND.t2124 VGND.t4 408.469
R1577 VGND.t2672 VGND.t181 408.469
R1578 VGND.t1175 VGND.t691 408.469
R1579 VGND.t2112 VGND.t1904 408.469
R1580 VGND.t2660 VGND.t2073 408.469
R1581 VGND.t1936 VGND.t1452 408.469
R1582 VGND.t10 VGND.t2158 408.469
R1583 VGND.t992 VGND.t1149 408.469
R1584 VGND.t1040 VGND.t2544 408.469
R1585 VGND.t1602 VGND.t391 408.469
R1586 VGND.t832 VGND.t814 408.469
R1587 VGND.t799 VGND.t84 408.469
R1588 VGND.t2401 VGND.t1870 408.469
R1589 VGND.t2260 VGND.t1980 408.469
R1590 VGND.t362 VGND.t80 408.469
R1591 VGND.t2487 VGND.t2053 408.469
R1592 VGND.t892 VGND.t2676 408.469
R1593 VGND.t2019 VGND.t1179 408.469
R1594 VGND.t2010 VGND.t2118 408.469
R1595 VGND.t2063 VGND.t2664 408.469
R1596 VGND.t127 VGND.t1171 408.469
R1597 VGND.t407 VGND.t2178 408.469
R1598 VGND.t176 VGND.t1732 408.469
R1599 VGND.t2320 VGND.t1446 408.469
R1600 VGND.t1181 VGND.t1344 408.469
R1601 VGND.t2634 VGND.t331 408.469
R1602 VGND.t249 VGND.t2666 408.469
R1603 VGND.t1401 VGND.t2445 408.469
R1604 VGND.t326 VGND.t2110 408.469
R1605 VGND.t315 VGND.t1734 408.469
R1606 VGND.t296 VGND.t456 408.469
R1607 VGND.t1329 VGND.t2174 408.469
R1608 VGND.t498 VGND.t381 408.469
R1609 VGND.t292 VGND.t2550 408.469
R1610 VGND.t1389 VGND.t1882 408.469
R1611 VGND.t1376 VGND.t820 408.469
R1612 VGND.t1542 VGND.t2546 408.469
R1613 VGND.t275 VGND.t2530 408.469
R1614 VGND.t1358 VGND.t1205 408.469
R1615 VGND.t1551 VGND.t2206 408.469
R1616 VGND.t2566 VGND.t549 397.848
R1617 VGND.t549 VGND.t660 397.848
R1618 VGND.t660 VGND.t522 397.848
R1619 VGND.t522 VGND.t230 397.848
R1620 VGND.t230 VGND.t231 397.848
R1621 VGND.t231 VGND.t234 397.848
R1622 VGND.t234 VGND.t235 397.848
R1623 VGND.t836 VGND.t1228 396.17
R1624 VGND.t1909 VGND.t1245 396.17
R1625 VGND.n2742 VGND.n559 394.137
R1626 VGND.n3008 VGND.n102 394.137
R1627 VGND.n2826 VGND.n101 394.137
R1628 VGND.n2755 VGND.n2754 394.137
R1629 VGND.n2753 VGND.n548 394.137
R1630 VGND.n2752 VGND.n549 394.137
R1631 VGND.n2751 VGND.n550 394.137
R1632 VGND.n2750 VGND.n551 394.137
R1633 VGND.n2749 VGND.n552 394.137
R1634 VGND.n2748 VGND.n553 394.137
R1635 VGND.n2747 VGND.n554 394.137
R1636 VGND.n2746 VGND.n555 394.137
R1637 VGND.n2745 VGND.n556 394.137
R1638 VGND.n2744 VGND.n557 394.137
R1639 VGND.n2743 VGND.n558 394.137
R1640 VGND.n3010 VGND.n3009 394.137
R1641 VGND.n2741 VGND.n2740 394.137
R1642 VGND.n491 VGND.t474 387.421
R1643 VGND.n2227 VGND.t77 387.421
R1644 VGND.n2225 VGND.t478 387.421
R1645 VGND.n1717 VGND.t670 387.421
R1646 VGND.n2850 VGND.t79 387.421
R1647 VGND.t1246 VGND.t2315 362.452
R1648 VGND.t2315 VGND.t976 345.594
R1649 VGND VGND.t335 328.616
R1650 VGND VGND.t481 328.616
R1651 VGND VGND.t489 328.616
R1652 VGND VGND.t547 328.616
R1653 VGND VGND.t957 328.616
R1654 VGND.t1380 VGND.t1561 313.776
R1655 VGND.t1555 VGND.t289 313.776
R1656 VGND.t274 VGND.t281 313.776
R1657 VGND.t1356 VGND.t259 313.776
R1658 VGND.t1549 VGND.t1368 313.776
R1659 VGND.t1533 VGND.t262 313.776
R1660 VGND.t1371 VGND.t328 313.776
R1661 VGND.t1362 VGND.t1346 313.776
R1662 VGND.t330 VGND.t1340 313.776
R1663 VGND.t1535 VGND.t263 313.776
R1664 VGND.t1343 VGND.t247 313.776
R1665 VGND.t1412 VGND.t1331 313.776
R1666 VGND.t317 VGND.t324 313.776
R1667 VGND.t312 VGND.t1414 313.776
R1668 VGND.t1393 VGND.t290 313.776
R1669 VGND.t1327 VGND.t314 313.776
R1670 VGND.t1228 VGND.t1237 311.877
R1671 VGND.t869 VGND.t1909 311.877
R1672 VGND.t1233 VGND 303.449
R1673 VGND.t1237 VGND 295.019
R1674 VGND.n333 VGND.t663 287.832
R1675 VGND VGND.t1593 286.591
R1676 VGND.n2161 VGND.t484 282.327
R1677 VGND.n346 VGND.t750 282.327
R1678 VGND.n2166 VGND.t674 281.13
R1679 VGND.n338 VGND.t2569 281.13
R1680 VGND.n470 VGND.t675 280.978
R1681 VGND.n470 VGND.t2360 280.978
R1682 VGND.n820 VGND.t1769 280.978
R1683 VGND.n820 VGND.t476 280.978
R1684 VGND.n2171 VGND.t512 280.978
R1685 VGND.n500 VGND.t1779 280.978
R1686 VGND.n500 VGND.t480 280.978
R1687 VGND.n434 VGND.t517 280.978
R1688 VGND.n434 VGND.t729 280.978
R1689 VGND.n403 VGND.t1847 280.978
R1690 VGND.n403 VGND.t583 280.978
R1691 VGND.n370 VGND.t2572 280.978
R1692 VGND.n370 VGND.t577 280.978
R1693 VGND.t763 VGND 278.161
R1694 VGND.n126 VGND 271.014
R1695 VGND.t1230 VGND 252.875
R1696 VGND.t1235 VGND 252.875
R1697 VGND.t520 VGND 252.875
R1698 VGND VGND.t524 252.875
R1699 VGND.t726 VGND 252.875
R1700 VGND.n2866 VGND.n455 244.329
R1701 VGND.n2864 VGND.n2863 244.329
R1702 VGND.n2859 VGND.n2854 244.329
R1703 VGND.n2857 VGND.n2856 244.329
R1704 VGND.n1323 VGND.t1182 241.393
R1705 VGND.n1135 VGND.t214 241.393
R1706 VGND.n220 VGND.t1053 241.393
R1707 VGND.n523 VGND.t455 241.393
R1708 VGND.n2443 VGND.t2675 241.393
R1709 VGND.n665 VGND.t1977 241.393
R1710 VGND.n671 VGND.t99 241.393
R1711 VGND.n802 VGND.t2535 241.393
R1712 VGND.n799 VGND.t445 241.393
R1713 VGND.n849 VGND.t1463 241.393
R1714 VGND.n1943 VGND.t1188 241.393
R1715 VGND.n971 VGND.t89 241.393
R1716 VGND.n977 VGND.t453 241.393
R1717 VGND.n1047 VGND.t87 241.393
R1718 VGND.n1044 VGND.t1220 241.393
R1719 VGND.n1129 VGND.t817 241.393
R1720 VGND.n55 VGND.t2545 241.393
R1721 VGND.n1058 VGND.t1056 241.393
R1722 VGND.n1328 VGND.t2635 241.284
R1723 VGND.n1127 VGND.t2667 241.284
R1724 VGND.n1393 VGND.t2446 241.284
R1725 VGND.n1388 VGND.t2111 241.284
R1726 VGND.n1383 VGND.t1735 241.284
R1727 VGND.n1378 VGND.t457 241.284
R1728 VGND.n1373 VGND.t2175 241.284
R1729 VGND.n1368 VGND.t382 241.284
R1730 VGND.n1363 VGND.t2551 241.284
R1731 VGND.n1358 VGND.t1883 241.284
R1732 VGND.n1353 VGND.t821 241.284
R1733 VGND.n1348 VGND.t2547 241.284
R1734 VGND.n1343 VGND.t2531 241.284
R1735 VGND.n1338 VGND.t1206 241.284
R1736 VGND.n1509 VGND.t1092 241.284
R1737 VGND.n1504 VGND.t1050 241.284
R1738 VGND.n1111 VGND.t1134 241.284
R1739 VGND.n1485 VGND.t1125 241.284
R1740 VGND.n1477 VGND.t1086 241.284
R1741 VGND.n1472 VGND.t1038 241.284
R1742 VGND.n1119 VGND.t1122 241.284
R1743 VGND.n1453 VGND.t1083 241.284
R1744 VGND.n1445 VGND.t1074 241.284
R1745 VGND.n1440 VGND.t1032 241.284
R1746 VGND.n1410 VGND.t1110 241.284
R1747 VGND.n1421 VGND.t1104 241.284
R1748 VGND.n1413 VGND.t1029 241.284
R1749 VGND.n1564 VGND.t1011 241.284
R1750 VGND.n1059 VGND.t1005 241.284
R1751 VGND.n1143 VGND.t2167 241.284
R1752 VGND.n1148 VGND.t396 241.284
R1753 VGND.n1140 VGND.t2205 241.284
R1754 VGND.n1198 VGND.t447 241.284
R1755 VGND.n1193 VGND.t1216 241.284
R1756 VGND.n1188 VGND.t97 241.284
R1757 VGND.n1183 VGND.t2539 241.284
R1758 VGND.n1178 VGND.t2649 241.284
R1759 VGND.n1173 VGND.t1975 241.284
R1760 VGND.n1168 VGND.t2255 241.284
R1761 VGND.n1163 VGND.t2637 241.284
R1762 VGND.n1158 VGND.t1965 241.284
R1763 VGND.n1153 VGND.t1178 241.284
R1764 VGND.n2727 VGND.t1152 241.284
R1765 VGND.n2732 VGND.t2663 241.284
R1766 VGND.n2927 VGND.t1002 241.284
R1767 VGND.n2932 VGND.t1008 241.284
R1768 VGND.n2937 VGND.t1014 241.284
R1769 VGND.n2942 VGND.t1101 241.284
R1770 VGND.n2947 VGND.t1107 241.284
R1771 VGND.n2952 VGND.t1020 241.284
R1772 VGND.n2957 VGND.t1062 241.284
R1773 VGND.n2962 VGND.t1077 241.284
R1774 VGND.n2967 VGND.t1113 241.284
R1775 VGND.n2972 VGND.t1035 241.284
R1776 VGND.n2977 VGND.t1080 241.284
R1777 VGND.n2982 VGND.t1119 241.284
R1778 VGND.n2987 VGND.t1131 241.284
R1779 VGND.n2992 VGND.t1047 241.284
R1780 VGND.n2997 VGND.t1089 241.284
R1781 VGND.n2845 VGND.t1140 241.284
R1782 VGND.n530 VGND.t212 241.284
R1783 VGND.n2763 VGND.t2062 241.284
R1784 VGND.n2768 VGND.t394 241.284
R1785 VGND.n2773 VGND.t2203 241.284
R1786 VGND.n2778 VGND.t2058 241.284
R1787 VGND.n2783 VGND.t1873 241.284
R1788 VGND.n2788 VGND.t1983 241.284
R1789 VGND.n2793 VGND.t83 241.284
R1790 VGND.n2798 VGND.t2645 241.284
R1791 VGND.n2803 VGND.t1969 241.284
R1792 VGND.n2808 VGND.t2249 241.284
R1793 VGND.n2813 VGND.t2123 241.284
R1794 VGND.n2818 VGND.t1449 241.284
R1795 VGND.n2823 VGND.t1174 241.284
R1796 VGND.n2446 VGND.t2241 241.284
R1797 VGND.n2470 VGND.t2115 241.284
R1798 VGND.n659 VGND.t1741 241.284
R1799 VGND.n2496 VGND.t948 241.284
R1800 VGND.n651 VGND.t2161 241.284
R1801 VGND.n2522 VGND.t1729 241.284
R1802 VGND.n643 VGND.t2468 241.284
R1803 VGND.n2548 VGND.t439 241.284
R1804 VGND.n635 VGND.t380 241.284
R1805 VGND.n2574 VGND.t2549 241.284
R1806 VGND.n627 VGND.t1879 241.284
R1807 VGND.n2605 VGND.t819 241.284
R1808 VGND.n2610 VGND.t2209 241.284
R1809 VGND.n2615 VGND.t2653 241.284
R1810 VGND.n619 VGND.t1222 241.284
R1811 VGND.n2457 VGND.t2046 241.284
R1812 VGND.n663 VGND.t2639 241.284
R1813 VGND.n2483 VGND.t1455 241.284
R1814 VGND.n655 VGND.t2243 241.284
R1815 VGND.n2509 VGND.t1154 241.284
R1816 VGND.n647 VGND.t1441 241.284
R1817 VGND.n2535 VGND.t950 241.284
R1818 VGND.n639 VGND.t2163 241.284
R1819 VGND.n2561 VGND.t1731 241.284
R1820 VGND.n631 VGND.t459 241.284
R1821 VGND.n2587 VGND.t402 241.284
R1822 VGND.n623 VGND.t218 241.284
R1823 VGND.n2592 VGND.t2553 241.284
R1824 VGND.n2632 VGND.t1224 241.284
R1825 VGND.n2637 VGND.t823 241.284
R1826 VGND.n690 VGND.t1865 241.284
R1827 VGND.n695 VGND.t1210 241.284
R1828 VGND.n700 VGND.t1184 241.284
R1829 VGND.n705 VGND.t2048 241.284
R1830 VGND.n710 VGND.t2671 241.284
R1831 VGND.n715 VGND.t1168 241.284
R1832 VGND.n720 VGND.t2245 241.284
R1833 VGND.n725 VGND.t1158 241.284
R1834 VGND.n730 VGND.t1443 241.284
R1835 VGND.n735 VGND.t2177 241.284
R1836 VGND.n740 VGND.t1146 241.284
R1837 VGND.n745 VGND.t2466 241.284
R1838 VGND.n686 VGND.t461 241.284
R1839 VGND.n2416 VGND.t825 241.284
R1840 VGND.n2411 VGND.t1727 241.284
R1841 VGND.n805 VGND.t384 241.284
R1842 VGND.n2252 VGND.t805 241.284
R1843 VGND.n793 VGND.t2251 241.284
R1844 VGND.n2278 VGND.t1861 241.284
R1845 VGND.n785 VGND.t1190 241.284
R1846 VGND.n2304 VGND.t2237 241.284
R1847 VGND.n777 VGND.t2042 241.284
R1848 VGND.n2330 VGND.t2659 241.284
R1849 VGND.n769 VGND.t944 241.284
R1850 VGND.n2356 VGND.t1162 241.284
R1851 VGND.n761 VGND.t1459 241.284
R1852 VGND.n2387 VGND.t940 241.284
R1853 VGND.n2392 VGND.t2171 241.284
R1854 VGND.n2397 VGND.t216 241.284
R1855 VGND.n2402 VGND.t2460 241.284
R1856 VGND.n2239 VGND.t1739 241.284
R1857 VGND.n797 VGND.t200 241.284
R1858 VGND.n2265 VGND.t2052 241.284
R1859 VGND.n789 VGND.t386 241.284
R1860 VGND.n2291 VGND.t91 241.284
R1861 VGND.n781 VGND.t2044 241.284
R1862 VGND.n2317 VGND.t1863 241.284
R1863 VGND.n773 VGND.t1967 241.284
R1864 VGND.n2343 VGND.t2239 241.284
R1865 VGND.n765 VGND.t2633 241.284
R1866 VGND.n2369 VGND.t1186 241.284
R1867 VGND.n757 VGND.t2235 241.284
R1868 VGND.n2374 VGND.t2109 241.284
R1869 VGND.n2657 VGND.t2462 241.284
R1870 VGND.n2662 VGND.t942 241.284
R1871 VGND.n2154 VGND.t2129 241.284
R1872 VGND.n854 VGND.t1160 241.284
R1873 VGND.n872 VGND.t220 241.284
R1874 VGND.n877 VGND.t932 241.284
R1875 VGND.n882 VGND.t398 241.284
R1876 VGND.n887 VGND.t206 241.284
R1877 VGND.n892 VGND.t2454 241.284
R1878 VGND.n897 VGND.t1877 241.284
R1879 VGND.n902 VGND.t813 241.284
R1880 VGND.n907 VGND.t2541 241.284
R1881 VGND.n912 VGND.t1867 241.284
R1882 VGND.n917 VGND.t807 241.284
R1883 VGND.n868 VGND.t103 241.284
R1884 VGND.n2134 VGND.t2641 241.284
R1885 VGND.n2129 VGND.t1212 241.284
R1886 VGND.n1946 VGND.t2655 241.284
R1887 VGND.n1970 VGND.t2681 241.284
R1888 VGND.n965 VGND.t2464 241.284
R1889 VGND.n1996 VGND.t2131 241.284
R1890 VGND.n957 VGND.t1142 241.284
R1891 VGND.n2022 VGND.t2456 241.284
R1892 VGND.n949 VGND.t934 241.284
R1893 VGND.n2048 VGND.t400 241.284
R1894 VGND.n941 VGND.t210 241.284
R1895 VGND.n2074 VGND.t449 241.284
R1896 VGND.n933 VGND.t390 241.284
R1897 VGND.n2105 VGND.t202 241.284
R1898 VGND.n2110 VGND.t2543 241.284
R1899 VGND.n2115 VGND.t1214 241.284
R1900 VGND.n2120 VGND.t809 241.284
R1901 VGND.n1957 VGND.t1226 241.284
R1902 VGND.n969 VGND.t1208 241.284
R1903 VGND.n1983 VGND.t946 241.284
R1904 VGND.n961 VGND.t2040 241.284
R1905 VGND.n2009 VGND.t1461 241.284
R1906 VGND.n953 VGND.t936 241.284
R1907 VGND.n2035 VGND.t2233 241.284
R1908 VGND.n945 VGND.t1144 241.284
R1909 VGND.n2061 VGND.t2458 241.284
R1910 VGND.n937 VGND.t2169 241.284
R1911 VGND.n2087 VGND.t1747 241.284
R1912 VGND.n929 VGND.t2452 241.284
R1913 VGND.n2092 VGND.t451 241.284
R1914 VGND.n2682 VGND.t811 241.284
R1915 VGND.n2687 VGND.t204 241.284
R1916 VGND.n1684 VGND.t1745 241.284
R1917 VGND.n1679 VGND.t208 241.284
R1918 VGND.n1674 VGND.t2060 241.284
R1919 VGND.n1669 VGND.t388 241.284
R1920 VGND.n1664 VGND.t101 241.284
R1921 VGND.n1659 VGND.t2050 241.284
R1922 VGND.n1654 VGND.t1869 241.284
R1923 VGND.n1649 VGND.t1979 241.284
R1924 VGND.n1644 VGND.t2253 241.284
R1925 VGND.n1639 VGND.t2643 241.284
R1926 VGND.n1634 VGND.t1963 241.284
R1927 VGND.n1629 VGND.t2247 241.284
R1928 VGND.n992 VGND.t2117 241.284
R1929 VGND.n1907 VGND.t1445 241.284
R1930 VGND.n1902 VGND.t1170 241.284
R1931 VGND.n1050 VGND.t1218 241.284
R1932 VGND.n1743 VGND.t1204 241.284
R1933 VGND.n1038 VGND.t938 241.284
R1934 VGND.n1769 VGND.t2651 241.284
R1935 VGND.n1030 VGND.t1457 241.284
R1936 VGND.n1795 VGND.t930 241.284
R1937 VGND.n1022 VGND.t2127 241.284
R1938 VGND.n1821 VGND.t1749 241.284
R1939 VGND.n1014 VGND.t2450 241.284
R1940 VGND.n1847 VGND.t2165 241.284
R1941 VGND.n1006 VGND.t1743 241.284
R1942 VGND.n1878 VGND.t2448 241.284
R1943 VGND.n1883 VGND.t441 241.284
R1944 VGND.n1888 VGND.t803 241.284
R1945 VGND.n1893 VGND.t198 241.284
R1946 VGND.n1730 VGND.t2533 241.284
R1947 VGND.n1042 VGND.t2056 241.284
R1948 VGND.n1756 VGND.t2679 241.284
R1949 VGND.n1034 VGND.t93 241.284
R1950 VGND.n1782 VGND.t2121 241.284
R1951 VGND.n1026 VGND.t2669 241.284
R1952 VGND.n1808 VGND.t1971 241.284
R1953 VGND.n1018 VGND.t928 241.284
R1954 VGND.n1834 VGND.t1156 241.284
R1955 VGND.n1010 VGND.t1451 241.284
R1956 VGND.n1860 VGND.t2173 241.284
R1957 VGND.n1002 VGND.t1148 241.284
R1958 VGND.n1865 VGND.t1737 241.284
R1959 VGND.n2707 VGND.t1881 241.284
R1960 VGND.n2712 VGND.t2157 241.284
R1961 VGND.n1315 VGND.t443 241.284
R1962 VGND.n1219 VGND.t1875 241.284
R1963 VGND.n1237 VGND.t1985 241.284
R1964 VGND.n1242 VGND.t2537 241.284
R1965 VGND.n1247 VGND.t2647 241.284
R1966 VGND.n1252 VGND.t1973 241.284
R1967 VGND.n1257 VGND.t95 241.284
R1968 VGND.n1262 VGND.t2125 241.284
R1969 VGND.n1267 VGND.t2673 241.284
R1970 VGND.n1272 VGND.t1176 241.284
R1971 VGND.n1277 VGND.t2113 241.284
R1972 VGND.n1282 VGND.t2661 241.284
R1973 VGND.n1233 VGND.t1453 241.284
R1974 VGND.n1295 VGND.t2159 241.284
R1975 VGND.n1290 VGND.t1150 241.284
R1976 VGND.n294 VGND.t392 241.284
R1977 VGND.n289 VGND.t815 241.284
R1978 VGND.n284 VGND.t85 241.284
R1979 VGND.n279 VGND.t1871 241.284
R1980 VGND.n274 VGND.t1981 241.284
R1981 VGND.n269 VGND.t81 241.284
R1982 VGND.n264 VGND.t2054 241.284
R1983 VGND.n259 VGND.t2677 241.284
R1984 VGND.n254 VGND.t1180 241.284
R1985 VGND.n249 VGND.t2119 241.284
R1986 VGND.n244 VGND.t2665 241.284
R1987 VGND.n239 VGND.t1172 241.284
R1988 VGND.n234 VGND.t2179 241.284
R1989 VGND.n229 VGND.t1733 241.284
R1990 VGND.n224 VGND.t1447 241.284
R1991 VGND.n1333 VGND.t2207 241.284
R1992 VGND.t2510 VGND.t213 222.15
R1993 VGND.t1525 VGND.t527 222.15
R1994 VGND.t572 VGND.t2166 222.15
R1995 VGND.t1663 VGND.t1502 222.15
R1996 VGND.t118 VGND.t395 222.15
R1997 VGND.t40 VGND.t66 222.15
R1998 VGND.t2204 VGND.t2516 222.15
R1999 VGND.t1313 VGND.t1 222.15
R2000 VGND.t446 VGND.t2508 222.15
R2001 VGND.t2299 VGND.t2335 222.15
R2002 VGND.t1215 VGND.t568 222.15
R2003 VGND.t2424 VGND.t44 222.15
R2004 VGND.t96 VGND.t566 222.15
R2005 VGND.t843 VGND.t2435 222.15
R2006 VGND.t2538 VGND.t2506 222.15
R2007 VGND.t1642 VGND.t2434 222.15
R2008 VGND.t2648 VGND.t2504 222.15
R2009 VGND.t767 VGND.t2303 222.15
R2010 VGND.t1974 VGND.t570 222.15
R2011 VGND.t555 VGND.t2396 222.15
R2012 VGND.t2254 VGND.t2514 222.15
R2013 VGND.t1494 VGND.t1952 222.15
R2014 VGND.t2636 VGND.t2512 222.15
R2015 VGND.t1706 VGND.t167 222.15
R2016 VGND.t1964 VGND.t564 222.15
R2017 VGND.t1940 VGND.t2586 222.15
R2018 VGND.t1177 VGND.t122 222.15
R2019 VGND.t23 VGND.t48 222.15
R2020 VGND.t120 VGND.t1151 222.15
R2021 VGND.t172 VGND.t907 222.15
R2022 VGND.t2662 VGND.t1483 222.15
R2023 VGND.t294 VGND.t2334 222.15
R2024 VGND.t1321 VGND.t1052 222.15
R2025 VGND.t2305 VGND.t311 222.15
R2026 VGND.t1001 VGND.t307 222.15
R2027 VGND.t1411 VGND.t1574 222.15
R2028 VGND.t1403 VGND.t1007 222.15
R2029 VGND.t1814 VGND.t1398 222.15
R2030 VGND.t1013 VGND.t1383 222.15
R2031 VGND.t1562 VGND.t1598 222.15
R2032 VGND.t504 VGND.t1100 222.15
R2033 VGND.t1920 VGND.t303 222.15
R2034 VGND.t1106 VGND.t285 222.15
R2035 VGND.t1385 VGND.t2367 222.15
R2036 VGND.t271 VGND.t1019 222.15
R2037 VGND.t178 VGND.t506 222.15
R2038 VGND.t1061 VGND.t500 222.15
R2039 VGND.t1550 VGND.t105 222.15
R2040 VGND.t1546 VGND.t1076 222.15
R2041 VGND.t1818 VGND.t273 222.15
R2042 VGND.t1112 VGND.t287 222.15
R2043 VGND.t1386 VGND.t834 222.15
R2044 VGND.t1366 VGND.t1034 222.15
R2045 VGND.t2395 VGND.t1548 222.15
R2046 VGND.t1079 VGND.t1351 222.15
R2047 VGND.t1538 VGND.t1227 222.15
R2048 VGND.t269 VGND.t1118 222.15
R2049 VGND.t1608 VGND.t264 222.15
R2050 VGND.t1130 VGND.t257 222.15
R2051 VGND.t1355 VGND.t1859 222.15
R2052 VGND.t241 VGND.t1046 222.15
R2053 VGND.t1986 VGND.t1332 222.15
R2054 VGND.t1088 VGND.t1531 222.15
R2055 VGND.t261 VGND.t973 222.15
R2056 VGND.t454 VGND.t1791 222.15
R2057 VGND.t1605 VGND.t2564 222.15
R2058 VGND.t2378 VGND.t1139 222.15
R2059 VGND.t1950 VGND.t2133 222.15
R2060 VGND.t2341 VGND.t211 222.15
R2061 VGND.t238 VGND.t2588 222.15
R2062 VGND.t2339 VGND.t2061 222.15
R2063 VGND.t1824 VGND.t1420 222.15
R2064 VGND.t1789 VGND.t393 222.15
R2065 VGND.t43 VGND.t1751 222.15
R2066 VGND.t2374 VGND.t2202 222.15
R2067 VGND.t979 VGND.t2268 222.15
R2068 VGND.t2372 VGND.t2057 222.15
R2069 VGND.t1241 VGND.t2490 222.15
R2070 VGND.t1787 VGND.t1872 222.15
R2071 VGND.t1481 VGND.t895 222.15
R2072 VGND.t1785 VGND.t1982 222.15
R2073 VGND.t1526 VGND.t2022 222.15
R2074 VGND.t2376 VGND.t82 222.15
R2075 VGND.t495 VGND.t2580 222.15
R2076 VGND.t2357 VGND.t2644 222.15
R2077 VGND.t2559 VGND.t463 222.15
R2078 VGND.t2355 VGND.t1968 222.15
R2079 VGND.t840 VGND.t2088 222.15
R2080 VGND.t2370 VGND.t2248 222.15
R2081 VGND.t2333 VGND.t410 222.15
R2082 VGND.t2368 VGND.t2122 222.15
R2083 VGND.t30 VGND.t2301 222.15
R2084 VGND.t2343 VGND.t1448 222.15
R2085 VGND.t1997 VGND.t991 222.15
R2086 VGND.t1783 VGND.t1173 222.15
R2087 VGND.t2089 VGND.t1370 222.15
R2088 VGND.t1835 VGND.t2674 222.15
R2089 VGND.t223 VGND.t2291 222.15
R2090 VGND.t2240 VGND.t2150 222.15
R2091 VGND.t541 VGND.t1668 222.15
R2092 VGND.t2275 VGND.t2114 222.15
R2093 VGND.t221 VGND.t853 222.15
R2094 VGND.t1740 VGND.t2273 222.15
R2095 VGND.t2404 VGND.t1804 222.15
R2096 VGND.t1833 VGND.t947 222.15
R2097 VGND.t2300 VGND.t886 222.15
R2098 VGND.t2160 VGND.t2266 222.15
R2099 VGND.t2557 VGND.t378 222.15
R2100 VGND.t2264 VGND.t1728 222.15
R2101 VGND.t2029 VGND.t112 222.15
R2102 VGND.t2467 VGND.t1831 222.15
R2103 VGND.t2313 VGND.t1908 222.15
R2104 VGND.t2154 VGND.t438 222.15
R2105 VGND.t353 VGND.t2038 222.15
R2106 VGND.t379 VGND.t2148 222.15
R2107 VGND.t622 VGND.t926 222.15
R2108 VGND.t1839 VGND.t2548 222.15
R2109 VGND.t917 VGND.t1493 222.15
R2110 VGND.t1878 VGND.t1837 222.15
R2111 VGND.t2478 VGND.t716 222.15
R2112 VGND.t2262 VGND.t818 222.15
R2113 VGND.t46 VGND.t916 222.15
R2114 VGND.t1806 VGND.t2208 222.15
R2115 VGND.t1816 VGND.t1830 222.15
R2116 VGND.t2277 VGND.t2652 222.15
R2117 VGND.t2332 VGND.t2323 222.15
R2118 VGND.t1221 VGND.t2152 222.15
R2119 VGND.t1560 VGND.t956 222.15
R2120 VGND.t1765 VGND.t1976 222.15
R2121 VGND.t493 VGND.t528 222.15
R2122 VGND.t154 VGND.t2045 222.15
R2123 VGND.t1269 VGND.t1808 222.15
R2124 VGND.t2638 VGND.t1633 222.15
R2125 VGND.t65 VGND.t1637 222.15
R2126 VGND.t1631 VGND.t1454 222.15
R2127 VGND.t186 VGND.t1315 222.15
R2128 VGND.t2242 VGND.t1763 222.15
R2129 VGND.t2345 VGND.t1248 222.15
R2130 VGND.t150 VGND.t1153 222.15
R2131 VGND.t2394 VGND.t2425 222.15
R2132 VGND.t1440 VGND.t148 222.15
R2133 VGND.t845 VGND.t19 222.15
R2134 VGND.t1761 VGND.t949 222.15
R2135 VGND.t492 VGND.t1644 222.15
R2136 VGND.t2162 VGND.t1759 222.15
R2137 VGND.t769 VGND.t2319 222.15
R2138 VGND.t152 VGND.t1730 222.15
R2139 VGND.t1244 VGND.t557 222.15
R2140 VGND.t458 VGND.t1629 222.15
R2141 VGND.t1898 VGND.t1514 222.15
R2142 VGND.t1767 VGND.t401 222.15
R2143 VGND.t188 VGND.t1702 222.15
R2144 VGND.t217 VGND.t146 222.15
R2145 VGND.t429 VGND.t1485 222.15
R2146 VGND.t2552 VGND.t144 222.15
R2147 VGND.t25 VGND.t1906 222.15
R2148 VGND.t1635 VGND.t1223 222.15
R2149 VGND.t20 VGND.t908 222.15
R2150 VGND.t822 VGND.t2380 222.15
R2151 VGND.t302 VGND.t21 222.15
R2152 VGND.t1677 VGND.t98 222.15
R2153 VGND.t1951 VGND.t1599 222.15
R2154 VGND.t347 VGND.t1864 222.15
R2155 VGND.t1708 VGND.t829 222.15
R2156 VGND.t640 VGND.t1209 222.15
R2157 VGND.t1480 VGND.t798 222.15
R2158 VGND.t1613 VGND.t1183 222.15
R2159 VGND.t1577 VGND.t1572 222.15
R2160 VGND.t1675 VGND.t2047 222.15
R2161 VGND.t2016 VGND.t2257 222.15
R2162 VGND.t343 VGND.t2670 222.15
R2163 VGND.t366 VGND.t1711 222.15
R2164 VGND.t341 VGND.t1167 222.15
R2165 VGND.t978 VGND.t2484 222.15
R2166 VGND.t1673 VGND.t2244 222.15
R2167 VGND.t2304 VGND.t76 222.15
R2168 VGND.t1671 VGND.t1157 222.15
R2169 VGND.t1479 VGND.t1680 222.15
R2170 VGND.t345 VGND.t1442 222.15
R2171 VGND.t31 VGND.t2012 222.15
R2172 VGND.t1611 VGND.t2176 222.15
R2173 VGND.t554 VGND.t377 222.15
R2174 VGND.t1609 VGND.t1145 222.15
R2175 VGND.t352 VGND.t129 222.15
R2176 VGND.t339 VGND.t2465 222.15
R2177 VGND.t1576 VGND.t404 222.15
R2178 VGND.t460 VGND.t337 222.15
R2179 VGND.t1998 VGND.t1709 222.15
R2180 VGND.t824 VGND.t642 222.15
R2181 VGND.t985 VGND.t2561 222.15
R2182 VGND.t1726 VGND.t1669 222.15
R2183 VGND.t1342 VGND.t721 222.15
R2184 VGND.t654 VGND.t2534 222.15
R2185 VGND.t1707 VGND.t2288 222.15
R2186 VGND.t383 VGND.t644 222.15
R2187 VGND.t2682 VGND.t1281 222.15
R2188 VGND.t2194 VGND.t804 222.15
R2189 VGND.t1822 VGND.t852 222.15
R2190 VGND.t2250 VGND.t2192 222.15
R2191 VGND.t2397 VGND.t592 222.15
R2192 VGND.t652 VGND.t1860 222.15
R2193 VGND.t1482 VGND.t2279 222.15
R2194 VGND.t1189 VGND.t2212 222.15
R2195 VGND.t2554 VGND.t974 222.15
R2196 VGND.t2210 VGND.t2236 222.15
R2197 VGND.t1725 VGND.t851 222.15
R2198 VGND.t2041 VGND.t650 222.15
R2199 VGND.t2306 VGND.t1954 222.15
R2200 VGND.t648 VGND.t2658 222.15
R2201 VGND.t714 VGND.t984 222.15
R2202 VGND.t943 VGND.t2214 222.15
R2203 VGND.t563 VGND.t1713 222.15
R2204 VGND.t2190 VGND.t1161 222.15
R2205 VGND.t32 VGND.t1490 222.15
R2206 VGND.t1458 VGND.t2188 222.15
R2207 VGND.t1995 VGND.t880 222.15
R2208 VGND.t2200 VGND.t939 222.15
R2209 VGND.t1907 VGND.t435 222.15
R2210 VGND.t2198 VGND.t2170 222.15
R2211 VGND.t350 VGND.t2472 222.15
R2212 VGND.t2196 VGND.t215 222.15
R2213 VGND.t1683 VGND.t1893 222.15
R2214 VGND.t2459 VGND.t646 222.15
R2215 VGND.t1537 VGND.t980 222.15
R2216 VGND.t444 VGND.t630 222.15
R2217 VGND.t534 VGND.t2293 222.15
R2218 VGND.t608 VGND.t1738 222.15
R2219 VGND.t1854 VGND.t542 222.15
R2220 VGND.t199 VGND.t739 222.15
R2221 VGND.t795 VGND.t1242 222.15
R2222 VGND.t636 VGND.t2051 222.15
R2223 VGND.t368 VGND.t2405 222.15
R2224 VGND.t385 VGND.t628 222.15
R2225 VGND.t887 VGND.t1659 222.15
R2226 VGND.t604 VGND.t90 222.15
R2227 VGND.t1504 VGND.t2558 222.15
R2228 VGND.t2043 VGND.t602 222.15
R2229 VGND.t113 VGND.t170 222.15
R2230 VGND.t626 VGND.t1862 222.15
R2231 VGND.t185 VGND.t1564 222.15
R2232 VGND.t1966 VGND.t624 222.15
R2233 VGND.t1925 VGND.t1581 222.15
R2234 VGND.t606 VGND.t2238 222.15
R2235 VGND.t1640 VGND.t623 222.15
R2236 VGND.t2632 VGND.t634 222.15
R2237 VGND.t1897 VGND.t351 222.15
R2238 VGND.t632 VGND.t1185 222.15
R2239 VGND.t29 VGND.t2479 222.15
R2240 VGND.t2234 VGND.t600 222.15
R2241 VGND.t1988 VGND.t1805 222.15
R2242 VGND.t2108 VGND.t743 222.15
R2243 VGND.t2147 VGND.t45 222.15
R2244 VGND.t741 VGND.t2461 222.15
R2245 VGND.t1261 VGND.t2324 222.15
R2246 VGND.t941 VGND.t610 222.15
R2247 VGND.t1563 VGND.t33 222.15
R2248 VGND.t1462 VGND.t971 222.15
R2249 VGND.t529 VGND.t881 222.15
R2250 VGND.t597 VGND.t2128 222.15
R2251 VGND.t73 VGND.t1809 222.15
R2252 VGND.t1621 VGND.t1159 222.15
R2253 VGND.t2565 VGND.t68 222.15
R2254 VGND.t1619 VGND.t219 222.15
R2255 VGND.t780 VGND.t1316 222.15
R2256 VGND.t969 VGND.t931 222.15
R2257 VGND.t1300 VGND.t2346 222.15
R2258 VGND.t593 VGND.t397 222.15
R2259 VGND.t2687 VGND.t752 222.15
R2260 VGND.t878 VGND.t205 222.15
R2261 VGND.t1623 VGND.t846 222.15
R2262 VGND.t967 VGND.t2453 222.15
R2263 VGND.t2027 VGND.t1645 222.15
R2264 VGND.t158 VGND.t1876 222.15
R2265 VGND.t1823 VGND.t770 222.15
R2266 VGND.t595 VGND.t812 222.15
R2267 VGND.t179 VGND.t558 222.15
R2268 VGND.t1617 VGND.t2540 222.15
R2269 VGND.t1923 VGND.t1899 222.15
R2270 VGND.t1615 VGND.t1866 222.15
R2271 VGND.t2432 VGND.t1703 222.15
R2272 VGND.t876 VGND.t806 222.15
R2273 VGND.t1921 VGND.t430 222.15
R2274 VGND.t102 VGND.t874 222.15
R2275 VGND.t26 VGND.t835 222.15
R2276 VGND.t2640 VGND.t872 222.15
R2277 VGND.t1884 VGND.t951 222.15
R2278 VGND.t1211 VGND.t156 222.15
R2279 VGND.t304 VGND.t74 222.15
R2280 VGND.t1468 VGND.t1187 222.15
R2281 VGND.t169 VGND.t526 222.15
R2282 VGND.t2654 VGND.t2184 222.15
R2283 VGND.t1503 VGND.t1584 222.15
R2284 VGND.t922 VGND.t2680 222.15
R2285 VGND.t187 VGND.t67 222.15
R2286 VGND.t2463 VGND.t920 222.15
R2287 VGND.t1314 VGND.t839 222.15
R2288 VGND.t1466 VGND.t2130 222.15
R2289 VGND.t911 VGND.t2298 222.15
R2290 VGND.t1141 VGND.t2180 222.15
R2291 VGND.t2423 VGND.t2382 222.15
R2292 VGND.t38 VGND.t2455 222.15
R2293 VGND.t171 VGND.t844 222.15
R2294 VGND.t933 VGND.t1464 222.15
R2295 VGND.t1643 VGND.t2410 222.15
R2296 VGND.t1661 VGND.t399 222.15
R2297 VGND.t1911 VGND.t768 222.15
R2298 VGND.t209 VGND.t2182 222.15
R2299 VGND.t556 VGND.t1579 222.15
R2300 VGND.t918 VGND.t448 222.15
R2301 VGND.t2411 VGND.t1495 222.15
R2302 VGND.t389 VGND.t1470 222.15
R2303 VGND.t1701 VGND.t222 222.15
R2304 VGND.t36 VGND.t201 222.15
R2305 VGND.t2560 VGND.t1941 222.15
R2306 VGND.t34 VGND.t2542 222.15
R2307 VGND.t2436 VGND.t24 222.15
R2308 VGND.t924 VGND.t1213 222.15
R2309 VGND.t779 VGND.t906 222.15
R2310 VGND.t808 VGND.t2186 222.15
R2311 VGND.t295 VGND.t1820 222.15
R2312 VGND.t2230 VGND.t88 222.15
R2313 VGND.t765 VGND.t871 222.15
R2314 VGND.t2220 VGND.t1225 222.15
R2315 VGND.t1842 VGND.t828 222.15
R2316 VGND.t1207 VGND.t1918 222.15
R2317 VGND.t801 VGND.t975 222.15
R2318 VGND.t1916 VGND.t945 222.15
R2319 VGND.t2615 VGND.t1571 222.15
R2320 VGND.t2039 VGND.t2228 222.15
R2321 VGND.t2256 VGND.t418 222.15
R2322 VGND.t2216 VGND.t1460 222.15
R2323 VGND.t713 VGND.t1710 222.15
R2324 VGND.t935 VGND.t1690 222.15
R2325 VGND.t2483 VGND.t1512 222.15
R2326 VGND.t2226 VGND.t2232 222.15
R2327 VGND.t1580 VGND.t75 222.15
R2328 VGND.t1143 VGND.t2224 222.15
R2329 VGND.t1679 VGND.t723 222.15
R2330 VGND.t2218 VGND.t2457 222.15
R2331 VGND.t1660 VGND.t2009 222.15
R2332 VGND.t2168 VGND.t1914 222.15
R2333 VGND.t376 VGND.t1924 222.15
R2334 VGND.t1912 VGND.t1746 222.15
R2335 VGND.t1638 VGND.t126 222.15
R2336 VGND.t2451 VGND.t1688 222.15
R2337 VGND.t403 VGND.t2412 222.15
R2338 VGND.t450 VGND.t1686 222.15
R2339 VGND.t175 VGND.t1510 222.15
R2340 VGND.t1684 VGND.t810 222.15
R2341 VGND.t2563 VGND.t2331 222.15
R2342 VGND.t203 VGND.t2222 222.15
R2343 VGND.t1337 VGND.t910 222.15
R2344 VGND.t452 VGND.t783 222.15
R2345 VGND.t2283 VGND.t2366 222.15
R2346 VGND.t1744 VGND.t2100 222.15
R2347 VGND.t2144 VGND.t168 222.15
R2348 VGND.t207 VGND.t791 222.15
R2349 VGND.t1473 VGND.t1163 222.15
R2350 VGND.t2059 VGND.t789 222.15
R2351 VGND.t2392 VGND.t2562 222.15
R2352 VGND.t387 VGND.t781 222.15
R2353 VGND.t357 VGND.t42 222.15
R2354 VGND.t100 VGND.t2096 222.15
R2355 VGND.t365 VGND.t2480 222.15
R2356 VGND.t2049 VGND.t2094 222.15
R2357 VGND.t864 VGND.t1639 222.15
R2358 VGND.t1868 VGND.t2106 222.15
R2359 VGND.t3 VGND.t2030 222.15
R2360 VGND.t1978 VGND.t2104 222.15
R2361 VGND.t180 VGND.t2393 222.15
R2362 VGND.t2252 VGND.t2098 222.15
R2363 VGND.t696 VGND.t1815 222.15
R2364 VGND.t2642 VGND.t787 222.15
R2365 VGND.t2066 VGND.t1843 222.15
R2366 VGND.t1962 VGND.t785 222.15
R2367 VGND.t2471 VGND.t722 222.15
R2368 VGND.t2246 VGND.t2092 222.15
R2369 VGND.t1935 VGND.t2415 222.15
R2370 VGND.t2116 VGND.t2090 222.15
R2371 VGND.t15 VGND.t841 222.15
R2372 VGND.t1444 VGND.t793 222.15
R2373 VGND.t901 VGND.t2614 222.15
R2374 VGND.t1169 VGND.t2102 222.15
R2375 VGND.t254 VGND.t1513 222.15
R2376 VGND.t1656 VGND.t86 222.15
R2377 VGND.t2 VGND.t2290 222.15
R2378 VGND.t1217 VGND.t1646 222.15
R2379 VGND.t2684 VGND.t1583 222.15
R2380 VGND.t1294 VGND.t1203 222.15
R2381 VGND.t1509 VGND.t854 222.15
R2382 VGND.t937 VGND.t1292 222.15
R2383 VGND.t2403 VGND.t1841 222.15
R2384 VGND.t1654 VGND.t2650 222.15
R2385 VGND.t27 VGND.t2281 222.15
R2386 VGND.t1456 VGND.t2441 222.15
R2387 VGND.t2556 VGND.t698 222.15
R2388 VGND.t2439 VGND.t929 222.15
R2389 VGND.t2338 VGND.t107 222.15
R2390 VGND.t2126 VGND.t1652 222.15
R2391 VGND.t2308 VGND.t909 222.15
R2392 VGND.t1650 VGND.t1748 222.15
R2393 VGND.t1308 VGND.t2033 222.15
R2394 VGND.t2449 VGND.t2443 222.15
R2395 VGND.t621 VGND.t104 222.15
R2396 VGND.t1290 VGND.t2164 222.15
R2397 VGND.t599 VGND.t1492 222.15
R2398 VGND.t1742 VGND.t1288 222.15
R2399 VGND.t1700 VGND.t1664 222.15
R2400 VGND.t2437 VGND.t2447 222.15
R2401 VGND.t1681 VGND.t437 222.15
R2402 VGND.t370 VGND.t440 222.15
R2403 VGND.t766 VGND.t1829 222.15
R2404 VGND.t1296 VGND.t802 222.15
R2405 VGND.t160 VGND.t2322 222.15
R2406 VGND.t197 VGND.t1648 222.15
R2407 VGND.t1557 VGND.t1506 222.15
R2408 VGND.t1219 VGND.t2656 222.15
R2409 VGND.t2282 VGND.t22 222.15
R2410 VGND.t2626 VGND.t2532 222.15
R2411 VGND.t49 VGND.t2143 222.15
R2412 VGND.t2055 VGND.t425 222.15
R2413 VGND.t1476 VGND.t2317 222.15
R2414 VGND.t423 VGND.t2678 222.15
R2415 VGND.t827 VGND.t2391 222.15
R2416 VGND.t92 VGND.t2430 222.15
R2417 VGND.t356 VGND.t1658 222.15
R2418 VGND.t2622 VGND.t2120 222.15
R2419 VGND.t0 VGND.t364 222.15
R2420 VGND.t2668 VGND.t2620 222.15
R2421 VGND.t2388 VGND.t1582 222.15
R2422 VGND.t2428 VGND.t1970 222.15
R2423 VGND.t638 VGND.t165 222.15
R2424 VGND.t927 VGND.t2426 222.15
R2425 VGND.t1274 VGND.t369 222.15
R2426 VGND.t2624 VGND.t1155 222.15
R2427 VGND.t2585 VGND.t693 222.15
R2428 VGND.t1450 VGND.t421 222.15
R2429 VGND.t2065 VGND.t1821 222.15
R2430 VGND.t419 VGND.t2172 222.15
R2431 VGND.t2433 VGND.t2075 222.15
R2432 VGND.t1147 VGND.t2618 222.15
R2433 VGND.t1934 VGND.t1240 222.15
R2434 VGND.t1736 VGND.t2616 222.15
R2435 VGND.t12 VGND.t225 222.15
R2436 VGND.t427 VGND.t1880 222.15
R2437 VGND.t28 VGND.t900 222.15
R2438 VGND.t2156 VGND.t2628 222.15
R2439 VGND.t251 VGND.t1803 222.15
R2440 VGND.t816 VGND.t142 222.15
R2441 VGND.t1604 VGND.t1496 222.15
R2442 VGND.t132 VGND.t442 222.15
R2443 VGND.t1624 VGND.t2132 222.15
R2444 VGND.t2598 VGND.t1874 222.15
R2445 VGND.t1515 VGND.t2595 222.15
R2446 VGND.t195 VGND.t1984 222.15
R2447 VGND.t1578 VGND.t1419 222.15
R2448 VGND.t140 VGND.t2536 222.15
R2449 VGND.t553 VGND.t1750 222.15
R2450 VGND.t2608 VGND.t2646 222.15
R2451 VGND.t639 VGND.t1712 222.15
R2452 VGND.t2606 VGND.t1972 222.15
R2453 VGND.t2028 VGND.t2489 222.15
R2454 VGND.t138 VGND.t94 222.15
R2455 VGND.t1953 VGND.t894 222.15
R2456 VGND.t136 VGND.t2124 222.15
R2457 VGND.t1959 VGND.t2021 222.15
R2458 VGND.t130 VGND.t2672 222.15
R2459 VGND.t1922 VGND.t2013 222.15
R2460 VGND.t193 VGND.t1175 222.15
R2461 VGND.t1597 VGND.t462 222.15
R2462 VGND.t191 VGND.t2112 222.15
R2463 VGND.t166 VGND.t2081 222.15
R2464 VGND.t2604 VGND.t2660 222.15
R2465 VGND.t190 VGND.t409 222.15
R2466 VGND.t1452 VGND.t2602 222.15
R2467 VGND.t1999 VGND.t699 222.15
R2468 VGND.t2158 VGND.t2600 222.15
R2469 VGND.t990 VGND.t697 222.15
R2470 VGND.t1149 VGND.t134 222.15
R2471 VGND.t1357 VGND.t1819 222.15
R2472 VGND.t2544 VGND.t1199 222.15
R2473 VGND.t2289 VGND.t2292 222.15
R2474 VGND.t391 VGND.t2630 222.15
R2475 VGND.t2683 VGND.t826 222.15
R2476 VGND.t814 VGND.t1430 222.15
R2477 VGND.t863 VGND.t2596 222.15
R2478 VGND.t84 VGND.t1428 222.15
R2479 VGND.t2398 VGND.t773 222.15
R2480 VGND.t1870 VGND.t1197 222.15
R2481 VGND.t2280 VGND.t1853 222.15
R2482 VGND.t1980 VGND.t1955 222.15
R2483 VGND.t2555 VGND.t1138 222.15
R2484 VGND.t80 VGND.t1438 222.15
R2485 VGND.t106 VGND.t1307 222.15
R2486 VGND.t2053 VGND.t1195 222.15
R2487 VGND.t2307 VGND.t1508 222.15
R2488 VGND.t2676 VGND.t1193 222.15
R2489 VGND.t2688 VGND.t18 222.15
R2490 VGND.t1179 VGND.t1957 222.15
R2491 VGND.t612 VGND.t1682 222.15
R2492 VGND.t2118 VGND.t1426 222.15
R2493 VGND.t1491 VGND.t2584 222.15
R2494 VGND.t2664 VGND.t1201 222.15
R2495 VGND.t1996 VGND.t2318 222.15
R2496 VGND.t1171 VGND.t1436 222.15
R2497 VGND.t436 VGND.t1667 222.15
R2498 VGND.t2178 VGND.t1434 222.15
R2499 VGND.t2473 VGND.t1497 222.15
R2500 VGND.t1732 VGND.t1432 222.15
R2501 VGND.t1894 VGND.t2314 222.15
R2502 VGND.t1446 VGND.t1191 222.15
R2503 VGND.t1539 VGND.t1301 222.15
R2504 VGND.t333 VGND.t1181 222.15
R2505 VGND.t2597 VGND.t1306 222.15
R2506 VGND.t252 VGND.t2634 222.15
R2507 VGND.t2414 VGND.t2140 222.15
R2508 VGND.t2666 VGND.t1347 222.15
R2509 VGND.t1472 VGND.t239 222.15
R2510 VGND.t2445 VGND.t1325 222.15
R2511 VGND.t1423 VGND.t1507 222.15
R2512 VGND.t2110 VGND.t322 222.15
R2513 VGND.t1758 VGND.t712 222.15
R2514 VGND.t1734 VGND.t1407 222.15
R2515 VGND.t2502 VGND.t491 222.15
R2516 VGND.t456 VGND.t1396 222.15
R2517 VGND.t2497 VGND.t2383 222.15
R2518 VGND.t2174 VGND.t318 222.15
R2519 VGND.t1268 VGND.t1802 222.15
R2520 VGND.t381 VGND.t300 222.15
R2521 VGND.t1279 VGND.t2413 222.15
R2522 VGND.t2550 VGND.t1409 222.15
R2523 VGND.t2581 VGND.t224 222.15
R2524 VGND.t1882 VGND.t502 222.15
R2525 VGND.t472 VGND.t774 222.15
R2526 VGND.t820 VGND.t1558 222.15
R2527 VGND.t2076 VGND.t1282 222.15
R2528 VGND.t2546 VGND.t1391 222.15
R2529 VGND.t417 VGND.t1243 222.15
R2530 VGND.t2530 VGND.t1378 222.15
R2531 VGND.t2302 VGND.t1817 222.15
R2532 VGND.t1205 VGND.t1353 222.15
R2533 VGND.t994 VGND.t2294 222.15
R2534 VGND.t2206 VGND.t279 222.15
R2535 VGND.t1382 VGND.t715 222.15
R2536 VGND.n477 VGND.n475 214.365
R2537 VGND.n477 VGND.n476 214.365
R2538 VGND.n467 VGND.n465 214.365
R2539 VGND.n467 VGND.n466 214.365
R2540 VGND.n485 VGND.n483 214.365
R2541 VGND.n485 VGND.n484 214.365
R2542 VGND.n827 VGND.n825 214.365
R2543 VGND.n827 VGND.n826 214.365
R2544 VGND.n817 VGND.n815 214.365
R2545 VGND.n817 VGND.n816 214.365
R2546 VGND.n835 VGND.n833 214.365
R2547 VGND.n835 VGND.n834 214.365
R2548 VGND.n2168 VGND.n2167 214.365
R2549 VGND.n507 VGND.n505 214.365
R2550 VGND.n507 VGND.n506 214.365
R2551 VGND.n497 VGND.n495 214.365
R2552 VGND.n497 VGND.n496 214.365
R2553 VGND.n515 VGND.n513 214.365
R2554 VGND.n515 VGND.n514 214.365
R2555 VGND.n1613 VGND.n1608 213.613
R2556 VGND.n1611 VGND.n1610 213.613
R2557 VGND.n1581 VGND.n1579 213.613
R2558 VGND.n1581 VGND.n1580 213.613
R2559 VGND.n1584 VGND.n1582 213.613
R2560 VGND.n1584 VGND.n1583 213.613
R2561 VGND.n2213 VGND.n2206 213.613
R2562 VGND.n2213 VGND.n2207 213.613
R2563 VGND.n2211 VGND.n2208 213.613
R2564 VGND.n2211 VGND.n2210 213.613
R2565 VGND.n1705 VGND.n1698 213.613
R2566 VGND.n1705 VGND.n1699 213.613
R2567 VGND.n1703 VGND.n1700 213.613
R2568 VGND.n1703 VGND.n1702 213.613
R2569 VGND.n2863 VGND.n457 212.329
R2570 VGND.n2859 VGND.n2858 212.329
R2571 VGND.n1625 VGND.t1585 211.359
R2572 VGND.n2165 VGND.n2164 207.965
R2573 VGND.n2182 VGND.n2162 207.965
R2574 VGND.n436 VGND.n432 207.965
R2575 VGND.n436 VGND.n433 207.965
R2576 VGND.n430 VGND.n428 207.965
R2577 VGND.n430 VGND.n429 207.965
R2578 VGND.n443 VGND.n426 207.965
R2579 VGND.n443 VGND.n427 207.965
R2580 VGND.n405 VGND.n401 207.965
R2581 VGND.n405 VGND.n402 207.965
R2582 VGND.n399 VGND.n397 207.965
R2583 VGND.n399 VGND.n398 207.965
R2584 VGND.n412 VGND.n395 207.965
R2585 VGND.n412 VGND.n396 207.965
R2586 VGND.n372 VGND.n368 207.965
R2587 VGND.n372 VGND.n369 207.965
R2588 VGND.n366 VGND.n364 207.965
R2589 VGND.n366 VGND.n365 207.965
R2590 VGND.n379 VGND.n362 207.965
R2591 VGND.n379 VGND.n363 207.965
R2592 VGND.n337 VGND.n336 207.965
R2593 VGND.n344 VGND.n328 207.965
R2594 VGND.n334 VGND.n332 207.965
R2595 VGND.n2181 VGND.n2163 207.213
R2596 VGND.n111 VGND.n110 207.213
R2597 VGND.n115 VGND.n109 207.213
R2598 VGND.n307 VGND.n305 207.213
R2599 VGND.n307 VGND.n306 207.213
R2600 VGND.n311 VGND.n303 207.213
R2601 VGND.n311 VGND.n304 207.213
R2602 VGND.n343 VGND.n329 207.213
R2603 VGND.n2886 VGND.n2884 207.213
R2604 VGND.n2886 VGND.n2885 207.213
R2605 VGND.n2890 VGND.n2881 207.213
R2606 VGND.n2890 VGND.n2882 207.213
R2607 VGND.n137 VGND.n135 207.213
R2608 VGND.n137 VGND.n136 207.213
R2609 VGND.n141 VGND.n132 207.213
R2610 VGND.n141 VGND.n133 207.213
R2611 VGND.t277 VGND.t1055 203.242
R2612 VGND.t1374 VGND.t1004 203.242
R2613 VGND.t1010 VGND.t1553 203.242
R2614 VGND.t1028 VGND.t1529 203.242
R2615 VGND.t1103 VGND.t1372 203.242
R2616 VGND.t1360 VGND.t1109 203.242
R2617 VGND.t1031 VGND.t1338 203.242
R2618 VGND.t265 VGND.t1073 203.242
R2619 VGND.t1082 VGND.t245 203.242
R2620 VGND.t1333 VGND.t1121 203.242
R2621 VGND.t1037 VGND.t320 203.242
R2622 VGND.t309 VGND.t1085 203.242
R2623 VGND.t1124 VGND.t1394 203.242
R2624 VGND.t1323 VGND.t1133 203.242
R2625 VGND.t1049 VGND.t298 203.242
R2626 VGND.t1405 VGND.t1091 203.242
R2627 VGND VGND.n204 194.419
R2628 VGND VGND.n2990 194.419
R2629 VGND VGND.n206 194.419
R2630 VGND VGND.n2980 194.419
R2631 VGND VGND.n208 194.419
R2632 VGND VGND.n2970 194.419
R2633 VGND VGND.n210 194.419
R2634 VGND VGND.n2960 194.419
R2635 VGND VGND.n212 194.419
R2636 VGND VGND.n2950 194.419
R2637 VGND VGND.n214 194.419
R2638 VGND VGND.n2940 194.419
R2639 VGND VGND.n216 194.419
R2640 VGND VGND.n2930 194.419
R2641 VGND VGND.n218 194.419
R2642 VGND.n1323 VGND.n1322 194.391
R2643 VGND.n1327 VGND.n1326 194.391
R2644 VGND.n1126 VGND.n1125 194.391
R2645 VGND.n1392 VGND.n1391 194.391
R2646 VGND.n1387 VGND.n1386 194.391
R2647 VGND.n1382 VGND.n1381 194.391
R2648 VGND.n1377 VGND.n1376 194.391
R2649 VGND.n1372 VGND.n1371 194.391
R2650 VGND.n1367 VGND.n1366 194.391
R2651 VGND.n1362 VGND.n1361 194.391
R2652 VGND.n1357 VGND.n1356 194.391
R2653 VGND.n1352 VGND.n1351 194.391
R2654 VGND.n1347 VGND.n1346 194.391
R2655 VGND.n1342 VGND.n1341 194.391
R2656 VGND.n1337 VGND.n1336 194.391
R2657 VGND.n1510 VGND.n1104 194.391
R2658 VGND.n1503 VGND.n1502 194.391
R2659 VGND.n1110 VGND.n1109 194.391
R2660 VGND.n1484 VGND.n1483 194.391
R2661 VGND.n1478 VGND.n1112 194.391
R2662 VGND.n1471 VGND.n1470 194.391
R2663 VGND.n1118 VGND.n1117 194.391
R2664 VGND.n1452 VGND.n1451 194.391
R2665 VGND.n1446 VGND.n1120 194.391
R2666 VGND.n1439 VGND.n1438 194.391
R2667 VGND.n1409 VGND.n1408 194.391
R2668 VGND.n1420 VGND.n1419 194.391
R2669 VGND.n1414 VGND.n1412 194.391
R2670 VGND.n1563 VGND.n1063 194.391
R2671 VGND.n1061 VGND.n1060 194.391
R2672 VGND.n1135 VGND.n1134 194.391
R2673 VGND.n1142 VGND.n1141 194.391
R2674 VGND.n1147 VGND.n1146 194.391
R2675 VGND.n1139 VGND.n1138 194.391
R2676 VGND.n1197 VGND.n1196 194.391
R2677 VGND.n1192 VGND.n1191 194.391
R2678 VGND.n1187 VGND.n1186 194.391
R2679 VGND.n1182 VGND.n1181 194.391
R2680 VGND.n1177 VGND.n1176 194.391
R2681 VGND.n1172 VGND.n1171 194.391
R2682 VGND.n1167 VGND.n1166 194.391
R2683 VGND.n1162 VGND.n1161 194.391
R2684 VGND.n1157 VGND.n1156 194.391
R2685 VGND.n1152 VGND.n1151 194.391
R2686 VGND.n2726 VGND.n2725 194.391
R2687 VGND.n2733 VGND.n565 194.391
R2688 VGND.n220 VGND.n219 194.391
R2689 VGND.n523 VGND.n522 194.391
R2690 VGND.n2844 VGND.n525 194.391
R2691 VGND.n531 VGND.n529 194.391
R2692 VGND.n2762 VGND.n2761 194.391
R2693 VGND.n2767 VGND.n2766 194.391
R2694 VGND.n2772 VGND.n2771 194.391
R2695 VGND.n2777 VGND.n2776 194.391
R2696 VGND.n2782 VGND.n2781 194.391
R2697 VGND.n2787 VGND.n2786 194.391
R2698 VGND.n2792 VGND.n2791 194.391
R2699 VGND.n2797 VGND.n2796 194.391
R2700 VGND.n2802 VGND.n2801 194.391
R2701 VGND.n2807 VGND.n2806 194.391
R2702 VGND.n2812 VGND.n2811 194.391
R2703 VGND.n2817 VGND.n2816 194.391
R2704 VGND.n2822 VGND.n2821 194.391
R2705 VGND.n2443 VGND.n2442 194.391
R2706 VGND.n2445 VGND.n2444 194.391
R2707 VGND.n2469 VGND.n2468 194.391
R2708 VGND.n658 VGND.n657 194.391
R2709 VGND.n2495 VGND.n2494 194.391
R2710 VGND.n650 VGND.n649 194.391
R2711 VGND.n2521 VGND.n2520 194.391
R2712 VGND.n642 VGND.n641 194.391
R2713 VGND.n2547 VGND.n2546 194.391
R2714 VGND.n634 VGND.n633 194.391
R2715 VGND.n2573 VGND.n2572 194.391
R2716 VGND.n626 VGND.n625 194.391
R2717 VGND.n2604 VGND.n2603 194.391
R2718 VGND.n2609 VGND.n2608 194.391
R2719 VGND.n2614 VGND.n2613 194.391
R2720 VGND.n618 VGND.n617 194.391
R2721 VGND.n665 VGND.n664 194.391
R2722 VGND.n2456 VGND.n2455 194.391
R2723 VGND.n662 VGND.n661 194.391
R2724 VGND.n2482 VGND.n2481 194.391
R2725 VGND.n654 VGND.n653 194.391
R2726 VGND.n2508 VGND.n2507 194.391
R2727 VGND.n646 VGND.n645 194.391
R2728 VGND.n2534 VGND.n2533 194.391
R2729 VGND.n638 VGND.n637 194.391
R2730 VGND.n2560 VGND.n2559 194.391
R2731 VGND.n630 VGND.n629 194.391
R2732 VGND.n2586 VGND.n2585 194.391
R2733 VGND.n622 VGND.n621 194.391
R2734 VGND.n2591 VGND.n2590 194.391
R2735 VGND.n2631 VGND.n2630 194.391
R2736 VGND.n2638 VGND.n613 194.391
R2737 VGND.n671 VGND.n670 194.391
R2738 VGND.n689 VGND.n688 194.391
R2739 VGND.n694 VGND.n693 194.391
R2740 VGND.n699 VGND.n698 194.391
R2741 VGND.n704 VGND.n703 194.391
R2742 VGND.n709 VGND.n708 194.391
R2743 VGND.n714 VGND.n713 194.391
R2744 VGND.n719 VGND.n718 194.391
R2745 VGND.n724 VGND.n723 194.391
R2746 VGND.n729 VGND.n728 194.391
R2747 VGND.n734 VGND.n733 194.391
R2748 VGND.n739 VGND.n738 194.391
R2749 VGND.n744 VGND.n743 194.391
R2750 VGND.n685 VGND.n684 194.391
R2751 VGND.n2415 VGND.n2414 194.391
R2752 VGND.n2410 VGND.n748 194.391
R2753 VGND.n802 VGND.n801 194.391
R2754 VGND.n804 VGND.n803 194.391
R2755 VGND.n2251 VGND.n2250 194.391
R2756 VGND.n792 VGND.n791 194.391
R2757 VGND.n2277 VGND.n2276 194.391
R2758 VGND.n784 VGND.n783 194.391
R2759 VGND.n2303 VGND.n2302 194.391
R2760 VGND.n776 VGND.n775 194.391
R2761 VGND.n2329 VGND.n2328 194.391
R2762 VGND.n768 VGND.n767 194.391
R2763 VGND.n2355 VGND.n2354 194.391
R2764 VGND.n760 VGND.n759 194.391
R2765 VGND.n2386 VGND.n2385 194.391
R2766 VGND.n2391 VGND.n2390 194.391
R2767 VGND.n2396 VGND.n2395 194.391
R2768 VGND.n2403 VGND.n751 194.391
R2769 VGND.n799 VGND.n798 194.391
R2770 VGND.n2238 VGND.n2237 194.391
R2771 VGND.n796 VGND.n795 194.391
R2772 VGND.n2264 VGND.n2263 194.391
R2773 VGND.n788 VGND.n787 194.391
R2774 VGND.n2290 VGND.n2289 194.391
R2775 VGND.n780 VGND.n779 194.391
R2776 VGND.n2316 VGND.n2315 194.391
R2777 VGND.n772 VGND.n771 194.391
R2778 VGND.n2342 VGND.n2341 194.391
R2779 VGND.n764 VGND.n763 194.391
R2780 VGND.n2368 VGND.n2367 194.391
R2781 VGND.n756 VGND.n755 194.391
R2782 VGND.n2373 VGND.n2372 194.391
R2783 VGND.n2656 VGND.n2655 194.391
R2784 VGND.n2663 VGND.n602 194.391
R2785 VGND.n849 VGND.n848 194.391
R2786 VGND.n2153 VGND.n851 194.391
R2787 VGND.n855 VGND.n853 194.391
R2788 VGND.n871 VGND.n870 194.391
R2789 VGND.n876 VGND.n875 194.391
R2790 VGND.n881 VGND.n880 194.391
R2791 VGND.n886 VGND.n885 194.391
R2792 VGND.n891 VGND.n890 194.391
R2793 VGND.n896 VGND.n895 194.391
R2794 VGND.n901 VGND.n900 194.391
R2795 VGND.n906 VGND.n905 194.391
R2796 VGND.n911 VGND.n910 194.391
R2797 VGND.n916 VGND.n915 194.391
R2798 VGND.n867 VGND.n866 194.391
R2799 VGND.n2133 VGND.n2132 194.391
R2800 VGND.n2128 VGND.n920 194.391
R2801 VGND.n1943 VGND.n1942 194.391
R2802 VGND.n1945 VGND.n1944 194.391
R2803 VGND.n1969 VGND.n1968 194.391
R2804 VGND.n964 VGND.n963 194.391
R2805 VGND.n1995 VGND.n1994 194.391
R2806 VGND.n956 VGND.n955 194.391
R2807 VGND.n2021 VGND.n2020 194.391
R2808 VGND.n948 VGND.n947 194.391
R2809 VGND.n2047 VGND.n2046 194.391
R2810 VGND.n940 VGND.n939 194.391
R2811 VGND.n2073 VGND.n2072 194.391
R2812 VGND.n932 VGND.n931 194.391
R2813 VGND.n2104 VGND.n2103 194.391
R2814 VGND.n2109 VGND.n2108 194.391
R2815 VGND.n2114 VGND.n2113 194.391
R2816 VGND.n2121 VGND.n923 194.391
R2817 VGND.n971 VGND.n970 194.391
R2818 VGND.n1956 VGND.n1955 194.391
R2819 VGND.n968 VGND.n967 194.391
R2820 VGND.n1982 VGND.n1981 194.391
R2821 VGND.n960 VGND.n959 194.391
R2822 VGND.n2008 VGND.n2007 194.391
R2823 VGND.n952 VGND.n951 194.391
R2824 VGND.n2034 VGND.n2033 194.391
R2825 VGND.n944 VGND.n943 194.391
R2826 VGND.n2060 VGND.n2059 194.391
R2827 VGND.n936 VGND.n935 194.391
R2828 VGND.n2086 VGND.n2085 194.391
R2829 VGND.n928 VGND.n927 194.391
R2830 VGND.n2091 VGND.n2090 194.391
R2831 VGND.n2681 VGND.n2680 194.391
R2832 VGND.n2688 VGND.n590 194.391
R2833 VGND.n977 VGND.n976 194.391
R2834 VGND.n1683 VGND.n1682 194.391
R2835 VGND.n1678 VGND.n1677 194.391
R2836 VGND.n1673 VGND.n1672 194.391
R2837 VGND.n1668 VGND.n1667 194.391
R2838 VGND.n1663 VGND.n1662 194.391
R2839 VGND.n1658 VGND.n1657 194.391
R2840 VGND.n1653 VGND.n1652 194.391
R2841 VGND.n1648 VGND.n1647 194.391
R2842 VGND.n1643 VGND.n1642 194.391
R2843 VGND.n1638 VGND.n1637 194.391
R2844 VGND.n1633 VGND.n1632 194.391
R2845 VGND.n1628 VGND.n1627 194.391
R2846 VGND.n991 VGND.n990 194.391
R2847 VGND.n1906 VGND.n1905 194.391
R2848 VGND.n1901 VGND.n993 194.391
R2849 VGND.n1047 VGND.n1046 194.391
R2850 VGND.n1049 VGND.n1048 194.391
R2851 VGND.n1742 VGND.n1741 194.391
R2852 VGND.n1037 VGND.n1036 194.391
R2853 VGND.n1768 VGND.n1767 194.391
R2854 VGND.n1029 VGND.n1028 194.391
R2855 VGND.n1794 VGND.n1793 194.391
R2856 VGND.n1021 VGND.n1020 194.391
R2857 VGND.n1820 VGND.n1819 194.391
R2858 VGND.n1013 VGND.n1012 194.391
R2859 VGND.n1846 VGND.n1845 194.391
R2860 VGND.n1005 VGND.n1004 194.391
R2861 VGND.n1877 VGND.n1876 194.391
R2862 VGND.n1882 VGND.n1881 194.391
R2863 VGND.n1887 VGND.n1886 194.391
R2864 VGND.n1894 VGND.n996 194.391
R2865 VGND.n1044 VGND.n1043 194.391
R2866 VGND.n1729 VGND.n1728 194.391
R2867 VGND.n1041 VGND.n1040 194.391
R2868 VGND.n1755 VGND.n1754 194.391
R2869 VGND.n1033 VGND.n1032 194.391
R2870 VGND.n1781 VGND.n1780 194.391
R2871 VGND.n1025 VGND.n1024 194.391
R2872 VGND.n1807 VGND.n1806 194.391
R2873 VGND.n1017 VGND.n1016 194.391
R2874 VGND.n1833 VGND.n1832 194.391
R2875 VGND.n1009 VGND.n1008 194.391
R2876 VGND.n1859 VGND.n1858 194.391
R2877 VGND.n1001 VGND.n1000 194.391
R2878 VGND.n1864 VGND.n1863 194.391
R2879 VGND.n2706 VGND.n2705 194.391
R2880 VGND.n2713 VGND.n577 194.391
R2881 VGND.n1129 VGND.n1128 194.391
R2882 VGND.n1314 VGND.n1131 194.391
R2883 VGND.n1220 VGND.n1218 194.391
R2884 VGND.n1236 VGND.n1235 194.391
R2885 VGND.n1241 VGND.n1240 194.391
R2886 VGND.n1246 VGND.n1245 194.391
R2887 VGND.n1251 VGND.n1250 194.391
R2888 VGND.n1256 VGND.n1255 194.391
R2889 VGND.n1261 VGND.n1260 194.391
R2890 VGND.n1266 VGND.n1265 194.391
R2891 VGND.n1271 VGND.n1270 194.391
R2892 VGND.n1276 VGND.n1275 194.391
R2893 VGND.n1281 VGND.n1280 194.391
R2894 VGND.n1232 VGND.n1231 194.391
R2895 VGND.n1294 VGND.n1293 194.391
R2896 VGND.n1289 VGND.n1285 194.391
R2897 VGND.n55 VGND.n54 194.391
R2898 VGND.n293 VGND.n292 194.391
R2899 VGND.n288 VGND.n287 194.391
R2900 VGND.n283 VGND.n282 194.391
R2901 VGND.n278 VGND.n277 194.391
R2902 VGND.n273 VGND.n272 194.391
R2903 VGND.n268 VGND.n267 194.391
R2904 VGND.n263 VGND.n262 194.391
R2905 VGND.n258 VGND.n257 194.391
R2906 VGND.n253 VGND.n252 194.391
R2907 VGND.n248 VGND.n247 194.391
R2908 VGND.n243 VGND.n242 194.391
R2909 VGND.n238 VGND.n237 194.391
R2910 VGND.n233 VGND.n232 194.391
R2911 VGND.n228 VGND.n227 194.391
R2912 VGND.n223 VGND.n222 194.391
R2913 VGND.n1058 VGND.n1057 194.391
R2914 VGND.n1332 VGND.n1331 194.391
R2915 VGND.n2865 VGND.n2864 176.941
R2916 VGND.n2855 VGND.n2854 176.941
R2917 VGND.n49 VGND.n48 161.308
R2918 VGND.n46 VGND.n45 161.308
R2919 VGND.n43 VGND.n42 161.308
R2920 VGND.n40 VGND.n39 161.308
R2921 VGND.n37 VGND.n36 161.308
R2922 VGND.n34 VGND.n33 161.308
R2923 VGND.n31 VGND.n30 161.308
R2924 VGND.n28 VGND.n27 161.308
R2925 VGND.n25 VGND.n24 161.308
R2926 VGND.n22 VGND.n21 161.308
R2927 VGND.n19 VGND.n18 161.308
R2928 VGND.n16 VGND.n15 161.308
R2929 VGND.n13 VGND.n12 161.308
R2930 VGND.n10 VGND.n9 161.308
R2931 VGND.n7 VGND.n6 161.308
R2932 VGND.n48 VGND.t2696 159.978
R2933 VGND.n45 VGND.t2699 159.978
R2934 VGND.n42 VGND.t2694 159.978
R2935 VGND.n39 VGND.t2690 159.978
R2936 VGND.n36 VGND.t2695 159.978
R2937 VGND.n33 VGND.t2703 159.978
R2938 VGND.n30 VGND.t2698 159.978
R2939 VGND.n27 VGND.t2692 159.978
R2940 VGND.n24 VGND.t2689 159.978
R2941 VGND.n21 VGND.t2691 159.978
R2942 VGND.n18 VGND.t2702 159.978
R2943 VGND.n15 VGND.t2693 159.978
R2944 VGND.n12 VGND.t2701 159.978
R2945 VGND.n9 VGND.t2697 159.978
R2946 VGND.n6 VGND.t2705 159.978
R2947 VGND.n2193 VGND.t764 159.315
R2948 VGND.n349 VGND.t2529 159.315
R2949 VGND.n1601 VGND.t1499 158.361
R2950 VGND.n155 VGND.t1666 158.361
R2951 VGND.n846 VGND.t762 157.291
R2952 VGND.n353 VGND.t2527 157.291
R2953 VGND.n808 VGND.t965 156.915
R2954 VGND.n360 VGND.t1231 156.915
R2955 VGND.n808 VGND.t963 156.915
R2956 VGND.n360 VGND.t1232 156.915
R2957 VGND.n810 VGND.t1575 154.131
R2958 VGND.n810 VGND.t78 154.131
R2959 VGND.n2193 VGND.t2032 154.131
R2960 VGND.n843 VGND.t1573 154.131
R2961 VGND.n385 VGND.t52 154.131
R2962 VGND.n385 VGND.t1801 154.131
R2963 VGND.n349 VGND.t838 154.131
R2964 VGND.n2902 VGND.t1247 154.131
R2965 VGND.n462 VGND.t962 153.631
R2966 VGND.n2199 VGND.t1505 153.631
R2967 VGND.n1691 VGND.t1280 153.631
R2968 VGND.n417 VGND.t1229 153.631
R2969 VGND.n2904 VGND.t2316 153.631
R2970 VGND.n2909 VGND.t1910 153.631
R2971 VGND.n2198 VGND.t2336 152.757
R2972 VGND.n2905 VGND.t977 152.757
R2973 VGND.n2188 VGND.t960 152.381
R2974 VGND.n326 VGND.t1236 152.381
R2975 VGND.n2158 VGND.n2157 152.174
R2976 VGND.n493 VGND.t964 150.922
R2977 VGND.n493 VGND.t958 150.922
R2978 VGND.n424 VGND.t1239 150.922
R2979 VGND.n424 VGND.t1234 150.922
R2980 VGND.n460 VGND.t475 150.922
R2981 VGND.n807 VGND.t1855 150.922
R2982 VGND.n492 VGND.t720 150.922
R2983 VGND.n423 VGND.t54 150.922
R2984 VGND.n392 VGND.t953 150.922
R2985 VGND.n359 VGND.t1252 150.922
R2986 VGND.n460 VGND.t1511 150.922
R2987 VGND.n807 VGND.t1284 150.922
R2988 VGND.n492 VGND.t2337 150.922
R2989 VGND.n423 VGND.t842 150.922
R2990 VGND.n392 VGND.t711 150.922
R2991 VGND.n359 VGND.t1626 150.922
R2992 VGND.n461 VGND.t961 147.411
R2993 VGND.n1690 VGND.t548 147.411
R2994 VGND.n416 VGND.t1238 147.411
R2995 VGND.n2910 VGND.t870 147.411
R2996 VGND.n847 VGND.t1594 146.964
R2997 VGND.n325 VGND.t229 146.964
R2998 VGND.n2860 VGND.n2859 146.25
R2999 VGND.n2861 VGND.n2860 146.25
R3000 VGND.n2856 VGND.n452 146.25
R3001 VGND.n2868 VGND.n452 146.25
R3002 VGND.n2863 VGND.n2862 146.25
R3003 VGND.n2862 VGND.n2861 146.25
R3004 VGND.n2867 VGND.n2866 146.25
R3005 VGND.n2868 VGND.n2867 146.25
R3006 VGND.n48 VGND.t1039 143.911
R3007 VGND.n45 VGND.t1114 143.911
R3008 VGND.n42 VGND.t1021 143.911
R3009 VGND.n39 VGND.t1063 143.911
R3010 VGND.n36 VGND.t1135 143.911
R3011 VGND.n33 VGND.t1042 143.911
R3012 VGND.n30 VGND.t1015 143.911
R3013 VGND.n27 VGND.t1057 143.911
R3014 VGND.n24 VGND.t1069 143.911
R3015 VGND.n21 VGND.t997 143.911
R3016 VGND.n18 VGND.t1093 143.911
R3017 VGND.n15 VGND.t1024 143.911
R3018 VGND.n12 VGND.t1096 143.911
R3019 VGND.n9 VGND.t1126 143.911
R3020 VGND.n6 VGND.t1066 143.911
R3021 VGND.n1719 VGND.n1626 143.478
R3022 VGND VGND.t2566 142.089
R3023 VGND.n1055 VGND.t1054 119.309
R3024 VGND.n1102 VGND.t1090 119.309
R3025 VGND.n202 VGND.t1087 119.309
R3026 VGND.n158 VGND.t1051 119.309
R3027 VGND.n160 VGND.t1000 119.309
R3028 VGND.n163 VGND.t1006 119.309
R3029 VGND.n166 VGND.t1012 119.309
R3030 VGND.n169 VGND.t1099 119.309
R3031 VGND.n172 VGND.t1105 119.309
R3032 VGND.n175 VGND.t1018 119.309
R3033 VGND.n178 VGND.t1060 119.309
R3034 VGND.n181 VGND.t1075 119.309
R3035 VGND.n184 VGND.t1111 119.309
R3036 VGND.n187 VGND.t1033 119.309
R3037 VGND.n190 VGND.t1078 119.309
R3038 VGND.n193 VGND.t1117 119.309
R3039 VGND.n196 VGND.t1129 119.309
R3040 VGND.n199 VGND.t1045 119.309
R3041 VGND.n1123 VGND.t1003 119.309
R3042 VGND.n1065 VGND.t1009 119.309
R3043 VGND.n1415 VGND.t1027 119.309
R3044 VGND.n1407 VGND.t1102 119.309
R3045 VGND.n1122 VGND.t1108 119.309
R3046 VGND.n1430 VGND.t1030 119.309
R3047 VGND.n1447 VGND.t1072 119.309
R3048 VGND.n1116 VGND.t1081 119.309
R3049 VGND.n1114 VGND.t1120 119.309
R3050 VGND.n1462 VGND.t1036 119.309
R3051 VGND.n1479 VGND.t1084 119.309
R3052 VGND.n1108 VGND.t1123 119.309
R3053 VGND.n1106 VGND.t1132 119.309
R3054 VGND.n1494 VGND.t1048 119.309
R3055 VGND.t1055 VGND.t1380 110.535
R3056 VGND.t1561 VGND.t966 110.535
R3057 VGND.t1004 VGND.t1555 110.535
R3058 VGND.t289 VGND.t2295 110.535
R3059 VGND.t281 VGND.t1010 110.535
R3060 VGND.t1961 VGND.t274 110.535
R3061 VGND.t259 VGND.t1028 110.535
R3062 VGND.t349 VGND.t1356 110.535
R3063 VGND.t1368 VGND.t1103 110.535
R3064 VGND.t41 VGND.t1549 110.535
R3065 VGND.t1109 VGND.t1533 110.535
R3066 VGND.t262 VGND.t367 110.535
R3067 VGND.t328 VGND.t1031 110.535
R3068 VGND.t2503 VGND.t1371 110.535
R3069 VGND.t1073 VGND.t1362 110.535
R3070 VGND.t1346 VGND.t1852 110.535
R3071 VGND.t1340 VGND.t1082 110.535
R3072 VGND.t2006 VGND.t330 110.535
R3073 VGND.t1121 VGND.t1535 110.535
R3074 VGND.t263 VGND.t189 110.535
R3075 VGND.t247 VGND.t1037 110.535
R3076 VGND.t494 VGND.t1343 110.535
R3077 VGND.t1085 VGND.t1412 110.535
R3078 VGND.t1331 VGND.t2416 110.535
R3079 VGND.t324 VGND.t1124 110.535
R3080 VGND.t1960 VGND.t317 110.535
R3081 VGND.t1133 VGND.t312 110.535
R3082 VGND.t1414 VGND.t47 110.535
R3083 VGND.t290 VGND.t1049 110.535
R3084 VGND.t981 VGND.t1393 110.535
R3085 VGND.t1091 VGND.t1327 110.535
R3086 VGND.t314 VGND.t2587 110.535
R3087 VGND.t1595 VGND.t1585 92.4699
R3088 VGND.t1592 VGND.t1595 92.4699
R3089 VGND.t1596 VGND.t1592 92.4699
R3090 VGND.t485 VGND.t1596 92.4699
R3091 VGND.t1774 VGND.t485 92.4699
R3092 VGND.t1717 VGND.t1774 92.4699
R3093 VGND.t2363 VGND.t1717 92.4699
R3094 VGND.n2865 VGND.t2700 88.3562
R3095 VGND.n2855 VGND.t2704 88.3562
R3096 VGND VGND.n1626 80.9529
R3097 VGND.n1626 VGND 75.1009
R3098 VGND.n1320 VGND 74.8566
R3099 VGND VGND.t2363 70.4533
R3100 VGND.n2866 VGND.n2865 67.3887
R3101 VGND.n2856 VGND.n2855 67.3887
R3102 VGND.n491 VGND 58.8055
R3103 VGND.n2227 VGND 58.8055
R3104 VGND.n2225 VGND 58.8055
R3105 VGND.n1717 VGND 58.8055
R3106 VGND.n2850 VGND 58.8055
R3107 VGND.n2854 VGND.n2852 53.1823
R3108 VGND.n2852 VGND.t1164 53.1823
R3109 VGND.n2857 VGND.n2853 53.1823
R3110 VGND.n2853 VGND.t1164 53.1823
R3111 VGND.n455 VGND.n453 53.1823
R3112 VGND.n453 VGND.t1164 53.1823
R3113 VGND.n2864 VGND.n454 53.1823
R3114 VGND.n454 VGND.t1164 53.1823
R3115 VGND.t1593 VGND.t483 50.5752
R3116 VGND.t1590 VGND.t1772 50.5752
R3117 VGND.t1588 VGND.t2521 50.5752
R3118 VGND.t1586 VGND.t673 50.5752
R3119 VGND.t236 VGND.t2568 50.5752
R3120 VGND.t232 VGND.t1845 50.5752
R3121 VGND.t226 VGND.t578 50.5752
R3122 VGND.t228 VGND.t749 50.5752
R3123 VGND VGND.n111 43.2063
R3124 VGND VGND.n307 43.2063
R3125 VGND VGND.n2886 43.2063
R3126 VGND VGND.n137 43.2063
R3127 VGND.n1322 VGND.t1345 34.8005
R3128 VGND.n1322 VGND.t334 34.8005
R3129 VGND.n1326 VGND.t332 34.8005
R3130 VGND.n1326 VGND.t253 34.8005
R3131 VGND.n1125 VGND.t250 34.8005
R3132 VGND.n1125 VGND.t1348 34.8005
R3133 VGND.n1391 VGND.t1402 34.8005
R3134 VGND.n1391 VGND.t1326 34.8005
R3135 VGND.n1386 VGND.t327 34.8005
R3136 VGND.n1386 VGND.t323 34.8005
R3137 VGND.n1381 VGND.t316 34.8005
R3138 VGND.n1381 VGND.t1408 34.8005
R3139 VGND.n1376 VGND.t297 34.8005
R3140 VGND.n1376 VGND.t1397 34.8005
R3141 VGND.n1371 VGND.t1330 34.8005
R3142 VGND.n1371 VGND.t319 34.8005
R3143 VGND.n1366 VGND.t499 34.8005
R3144 VGND.n1366 VGND.t301 34.8005
R3145 VGND.n1361 VGND.t293 34.8005
R3146 VGND.n1361 VGND.t1410 34.8005
R3147 VGND.n1356 VGND.t1390 34.8005
R3148 VGND.n1356 VGND.t503 34.8005
R3149 VGND.n1351 VGND.t1377 34.8005
R3150 VGND.n1351 VGND.t1559 34.8005
R3151 VGND.n1346 VGND.t1543 34.8005
R3152 VGND.n1346 VGND.t1392 34.8005
R3153 VGND.n1341 VGND.t276 34.8005
R3154 VGND.n1341 VGND.t1379 34.8005
R3155 VGND.n1336 VGND.t1359 34.8005
R3156 VGND.n1336 VGND.t1354 34.8005
R3157 VGND.n1104 VGND.t1406 34.8005
R3158 VGND.n1104 VGND.t1328 34.8005
R3159 VGND.n1502 VGND.t299 34.8005
R3160 VGND.n1502 VGND.t291 34.8005
R3161 VGND.n1109 VGND.t1324 34.8005
R3162 VGND.n1109 VGND.t313 34.8005
R3163 VGND.n1483 VGND.t1395 34.8005
R3164 VGND.n1483 VGND.t325 34.8005
R3165 VGND.n1112 VGND.t310 34.8005
R3166 VGND.n1112 VGND.t1413 34.8005
R3167 VGND.n1470 VGND.t321 34.8005
R3168 VGND.n1470 VGND.t248 34.8005
R3169 VGND.n1117 VGND.t1334 34.8005
R3170 VGND.n1117 VGND.t1536 34.8005
R3171 VGND.n1451 VGND.t246 34.8005
R3172 VGND.n1451 VGND.t1341 34.8005
R3173 VGND.n1120 VGND.t266 34.8005
R3174 VGND.n1120 VGND.t1363 34.8005
R3175 VGND.n1438 VGND.t1339 34.8005
R3176 VGND.n1438 VGND.t329 34.8005
R3177 VGND.n1408 VGND.t1361 34.8005
R3178 VGND.n1408 VGND.t1534 34.8005
R3179 VGND.n1419 VGND.t1373 34.8005
R3180 VGND.n1419 VGND.t1369 34.8005
R3181 VGND.n1412 VGND.t1530 34.8005
R3182 VGND.n1412 VGND.t260 34.8005
R3183 VGND.n1063 VGND.t1554 34.8005
R3184 VGND.n1063 VGND.t282 34.8005
R3185 VGND.n1060 VGND.t1375 34.8005
R3186 VGND.n1060 VGND.t1556 34.8005
R3187 VGND.n1134 VGND.t1068 34.8005
R3188 VGND.n1134 VGND.t2511 34.8005
R3189 VGND.n1141 VGND.t533 34.8005
R3190 VGND.n1141 VGND.t573 34.8005
R3191 VGND.n1146 VGND.t540 34.8005
R3192 VGND.n1146 VGND.t119 34.8005
R3193 VGND.n1138 VGND.t860 34.8005
R3194 VGND.n1138 VGND.t2517 34.8005
R3195 VGND.n1196 VGND.t1945 34.8005
R3196 VGND.n1196 VGND.t2509 34.8005
R3197 VGND.n1191 VGND.t885 34.8005
R3198 VGND.n1191 VGND.t569 34.8005
R3199 VGND.n1186 VGND.t2270 34.8005
R3200 VGND.n1186 VGND.t567 34.8005
R3201 VGND.n1181 VGND.t109 34.8005
R3202 VGND.n1181 VGND.t2507 34.8005
R3203 VGND.n1176 VGND.t2310 34.8005
R3204 VGND.n1176 VGND.t2505 34.8005
R3205 VGND.n1171 VGND.t2035 34.8005
R3206 VGND.n1171 VGND.t571 34.8005
R3207 VGND.n1166 VGND.t614 34.8005
R3208 VGND.n1166 VGND.t2515 34.8005
R3209 VGND.n1161 VGND.t465 34.8005
R3210 VGND.n1161 VGND.t2513 34.8005
R3211 VGND.n1156 VGND.t1693 34.8005
R3212 VGND.n1156 VGND.t565 34.8005
R3213 VGND.n1151 VGND.t913 34.8005
R3214 VGND.n1151 VGND.t123 34.8005
R3215 VGND.n2725 VGND.t2477 34.8005
R3216 VGND.n2725 VGND.t121 34.8005
R3217 VGND.n565 VGND.t1886 34.8005
R3218 VGND.n565 VGND.t1484 34.8005
R3219 VGND.n219 VGND.t1400 34.8005
R3220 VGND.n219 VGND.t1322 34.8005
R3221 VGND.n204 VGND.t1350 34.8005
R3222 VGND.n204 VGND.t1532 34.8005
R3223 VGND.n2990 VGND.t244 34.8005
R3224 VGND.n2990 VGND.t242 34.8005
R3225 VGND.n206 VGND.t1528 34.8005
R3226 VGND.n206 VGND.t258 34.8005
R3227 VGND.n2980 VGND.t1336 34.8005
R3228 VGND.n2980 VGND.t270 34.8005
R3229 VGND.n208 VGND.t256 34.8005
R3230 VGND.n208 VGND.t1352 34.8005
R3231 VGND.n2970 VGND.t268 34.8005
R3232 VGND.n2970 VGND.t1367 34.8005
R3233 VGND.n210 VGND.t1541 34.8005
R3234 VGND.n210 VGND.t288 34.8005
R3235 VGND.n2960 VGND.t1365 34.8005
R3236 VGND.n2960 VGND.t1547 34.8005
R3237 VGND.n212 VGND.t1388 34.8005
R3238 VGND.n212 VGND.t501 34.8005
R3239 VGND.n2950 VGND.t1545 34.8005
R3240 VGND.n2950 VGND.t272 34.8005
R3241 VGND.n214 VGND.t497 34.8005
R3242 VGND.n214 VGND.t286 34.8005
R3243 VGND.n2940 VGND.t508 34.8005
R3244 VGND.n2940 VGND.t505 34.8005
R3245 VGND.n216 VGND.t284 34.8005
R3246 VGND.n216 VGND.t1384 34.8005
R3247 VGND.n2930 VGND.t306 34.8005
R3248 VGND.n2930 VGND.t1404 34.8005
R3249 VGND.n218 VGND.t510 34.8005
R3250 VGND.n218 VGND.t308 34.8005
R3251 VGND.n522 VGND.t1116 34.8005
R3252 VGND.n522 VGND.t1792 34.8005
R3253 VGND.n525 VGND.t2287 34.8005
R3254 VGND.n525 VGND.t2379 34.8005
R3255 VGND.n529 VGND.t1501 34.8005
R3256 VGND.n529 VGND.t2342 34.8005
R3257 VGND.n2761 VGND.t1475 34.8005
R3258 VGND.n2761 VGND.t2340 34.8005
R3259 VGND.n2766 VGND.t1425 34.8005
R3260 VGND.n2766 VGND.t1790 34.8005
R3261 VGND.n2771 VGND.t2297 34.8005
R3262 VGND.n2771 VGND.t2375 34.8005
R3263 VGND.n2776 VGND.t760 34.8005
R3264 VGND.n2776 VGND.t2373 34.8005
R3265 VGND.n2781 VGND.t868 34.8005
R3266 VGND.n2781 VGND.t1788 34.8005
R3267 VGND.n2786 VGND.t7 34.8005
R3268 VGND.n2786 VGND.t1786 34.8005
R3269 VGND.n2791 VGND.t184 34.8005
R3270 VGND.n2791 VGND.t2377 34.8005
R3271 VGND.n2796 VGND.t695 34.8005
R3272 VGND.n2796 VGND.t2358 34.8005
R3273 VGND.n2801 VGND.t1489 34.8005
R3274 VGND.n2801 VGND.t2356 34.8005
R3275 VGND.n2806 VGND.t2470 34.8005
R3276 VGND.n2806 VGND.t2371 34.8005
R3277 VGND.n2811 VGND.t1939 34.8005
R3278 VGND.n2811 VGND.t2369 34.8005
R3279 VGND.n2816 VGND.t14 34.8005
R3280 VGND.n2816 VGND.t2344 34.8005
R3281 VGND.n2821 VGND.t996 34.8005
R3282 VGND.n2821 VGND.t1784 34.8005
R3283 VGND.n2442 VGND.t1023 34.8005
R3284 VGND.n2442 VGND.t1836 34.8005
R3285 VGND.n2444 VGND.t1303 34.8005
R3286 VGND.n2444 VGND.t2151 34.8005
R3287 VGND.n2468 VGND.t2137 34.8005
R3288 VGND.n2468 VGND.t2276 34.8005
R3289 VGND.n657 VGND.t2592 34.8005
R3290 VGND.n657 VGND.t2274 34.8005
R3291 VGND.n2494 VGND.t2409 34.8005
R3292 VGND.n2494 VGND.t1834 34.8005
R3293 VGND.n649 VGND.t1755 34.8005
R3294 VGND.n649 VGND.t2267 34.8005
R3295 VGND.n2520 VGND.t2420 34.8005
R3296 VGND.n2520 VGND.t2265 34.8005
R3297 VGND.n641 VGND.t2494 34.8005
R3298 VGND.n641 VGND.t1832 34.8005
R3299 VGND.n2546 VGND.t1265 34.8005
R3300 VGND.n2546 VGND.t2155 34.8005
R3301 VGND.n633 VGND.t2026 34.8005
R3302 VGND.n633 VGND.t2149 34.8005
R3303 VGND.n2572 VGND.t2577 34.8005
R3304 VGND.n2572 VGND.t1840 34.8005
R3305 VGND.n625 VGND.t2070 34.8005
R3306 VGND.n625 VGND.t1838 34.8005
R3307 VGND.n2603 VGND.t2085 34.8005
R3308 VGND.n2603 VGND.t2263 34.8005
R3309 VGND.n2608 VGND.t414 34.8005
R3310 VGND.n2608 VGND.t1807 34.8005
R3311 VGND.n2613 VGND.t2003 34.8005
R3312 VGND.n2613 VGND.t2278 34.8005
R3313 VGND.n617 VGND.t2328 34.8005
R3314 VGND.n617 VGND.t2153 34.8005
R3315 VGND.n664 VGND.t1065 34.8005
R3316 VGND.n664 VGND.t1766 34.8005
R3317 VGND.n2455 VGND.t536 34.8005
R3318 VGND.n2455 VGND.t155 34.8005
R3319 VGND.n661 VGND.t544 34.8005
R3320 VGND.n661 VGND.t1634 34.8005
R3321 VGND.n2481 VGND.t858 34.8005
R3322 VGND.n2481 VGND.t1632 34.8005
R3323 VGND.n653 VGND.t1947 34.8005
R3324 VGND.n653 VGND.t1764 34.8005
R3325 VGND.n2507 VGND.t889 34.8005
R3326 VGND.n2507 VGND.t151 34.8005
R3327 VGND.n645 VGND.t2499 34.8005
R3328 VGND.n645 VGND.t149 34.8005
R3329 VGND.n2533 VGND.t115 34.8005
R3330 VGND.n2533 VGND.t1762 34.8005
R3331 VGND.n637 VGND.t1566 34.8005
R3332 VGND.n637 VGND.t1760 34.8005
R3333 VGND.n2559 VGND.t1927 34.8005
R3334 VGND.n2559 VGND.t153 34.8005
R3335 VGND.n629 VGND.t618 34.8005
R3336 VGND.n629 VGND.t1630 34.8005
R3337 VGND.n2585 VGND.t469 34.8005
R3338 VGND.n2585 VGND.t1768 34.8005
R3339 VGND.n621 VGND.t1697 34.8005
R3340 VGND.n621 VGND.t147 34.8005
R3341 VGND.n2590 VGND.t1990 34.8005
R3342 VGND.n2590 VGND.t145 34.8005
R3343 VGND.n2630 VGND.t1826 34.8005
R3344 VGND.n2630 VGND.t1636 34.8005
R3345 VGND.n613 VGND.t1890 34.8005
R3346 VGND.n613 VGND.t2381 34.8005
R3347 VGND.n670 VGND.t1137 34.8005
R3348 VGND.n670 VGND.t1678 34.8005
R3349 VGND.n688 VGND.t1520 34.8005
R3350 VGND.n688 VGND.t348 34.8005
R3351 VGND.n693 VGND.t2142 34.8005
R3352 VGND.n693 VGND.t641 34.8005
R3353 VGND.n698 VGND.t897 34.8005
R3354 VGND.n698 VGND.t1614 34.8005
R3355 VGND.n703 VGND.t1418 34.8005
R3356 VGND.n703 VGND.t1676 34.8005
R3357 VGND.n708 VGND.t355 34.8005
R3358 VGND.n708 VGND.t344 34.8005
R3359 VGND.n713 VGND.t756 34.8005
R3360 VGND.n713 VGND.t342 34.8005
R3361 VGND.n718 VGND.t2387 34.8005
R3362 VGND.n718 VGND.t1674 34.8005
R3363 VGND.n723 VGND.t164 34.8005
R3364 VGND.n723 VGND.t1672 34.8005
R3365 VGND.n728 VGND.t1273 34.8005
R3366 VGND.n728 VGND.t346 34.8005
R3367 VGND.n733 VGND.t690 34.8005
R3368 VGND.n733 VGND.t1612 34.8005
R3369 VGND.n738 VGND.t1903 34.8005
R3370 VGND.n738 VGND.t1610 34.8005
R3371 VGND.n743 VGND.t2080 34.8005
R3372 VGND.n743 VGND.t340 34.8005
R3373 VGND.n684 VGND.t1933 34.8005
R3374 VGND.n684 VGND.t338 34.8005
R3375 VGND.n2414 VGND.t9 34.8005
R3376 VGND.n2414 VGND.t643 34.8005
R3377 VGND.n748 VGND.t989 34.8005
R3378 VGND.n748 VGND.t1670 34.8005
R3379 VGND.n801 VGND.t1044 34.8005
R3380 VGND.n801 VGND.t655 34.8005
R3381 VGND.n803 VGND.t1601 34.8005
R3382 VGND.n803 VGND.t645 34.8005
R3383 VGND.n2250 VGND.t831 34.8005
R3384 VGND.n2250 VGND.t2195 34.8005
R3385 VGND.n791 VGND.t797 34.8005
R3386 VGND.n791 VGND.t2193 34.8005
R3387 VGND.n2276 VGND.t2400 34.8005
R3388 VGND.n2276 VGND.t653 34.8005
R3389 VGND.n783 VGND.t2259 34.8005
R3390 VGND.n783 VGND.t2213 34.8005
R3391 VGND.n2302 VGND.t361 34.8005
R3392 VGND.n2302 VGND.t2211 34.8005
R3393 VGND.n775 VGND.t2486 34.8005
R3394 VGND.n775 VGND.t651 34.8005
R3395 VGND.n2328 VGND.t891 34.8005
R3396 VGND.n2328 VGND.t649 34.8005
R3397 VGND.n767 VGND.t2018 34.8005
R3398 VGND.n767 VGND.t2215 34.8005
R3399 VGND.n2354 VGND.t2008 34.8005
R3400 VGND.n2354 VGND.t2191 34.8005
R3401 VGND.n759 VGND.t1487 34.8005
R3402 VGND.n759 VGND.t2189 34.8005
R3403 VGND.n2385 VGND.t125 34.8005
R3404 VGND.n2385 VGND.t2201 34.8005
R3405 VGND.n2390 VGND.t406 34.8005
R3406 VGND.n2390 VGND.t2199 34.8005
R3407 VGND.n2395 VGND.t174 34.8005
R3408 VGND.n2395 VGND.t2197 34.8005
R3409 VGND.n751 VGND.t1896 34.8005
R3410 VGND.n751 VGND.t647 34.8005
R3411 VGND.n798 VGND.t1017 34.8005
R3412 VGND.n798 VGND.t631 34.8005
R3413 VGND.n2237 VGND.t1305 34.8005
R3414 VGND.n2237 VGND.t609 34.8005
R3415 VGND.n795 VGND.t2139 34.8005
R3416 VGND.n795 VGND.t740 34.8005
R3417 VGND.n2263 VGND.t2590 34.8005
R3418 VGND.n2263 VGND.t637 34.8005
R3419 VGND.n787 VGND.t1570 34.8005
R3420 VGND.n787 VGND.t629 34.8005
R3421 VGND.n2289 VGND.t1757 34.8005
R3422 VGND.n2289 VGND.t605 34.8005
R3423 VGND.n779 VGND.t2422 34.8005
R3424 VGND.n779 VGND.t603 34.8005
R3425 VGND.n2315 VGND.t2496 34.8005
R3426 VGND.n2315 VGND.t627 34.8005
R3427 VGND.n771 VGND.t1267 34.8005
R3428 VGND.n771 VGND.t625 34.8005
R3429 VGND.n2341 VGND.t1278 34.8005
R3430 VGND.n2341 VGND.t607 34.8005
R3431 VGND.n763 VGND.t2579 34.8005
R3432 VGND.n763 VGND.t635 34.8005
R3433 VGND.n2367 VGND.t2519 34.8005
R3434 VGND.n2367 VGND.t633 34.8005
R3435 VGND.n755 VGND.t2087 34.8005
R3436 VGND.n755 VGND.t601 34.8005
R3437 VGND.n2372 VGND.t416 34.8005
R3438 VGND.n2372 VGND.t744 34.8005
R3439 VGND.n2655 VGND.t2005 34.8005
R3440 VGND.n2655 VGND.t742 34.8005
R3441 VGND.n602 VGND.t2330 34.8005
R3442 VGND.n602 VGND.t611 34.8005
R3443 VGND.n848 VGND.t1059 34.8005
R3444 VGND.n848 VGND.t972 34.8005
R3445 VGND.n851 VGND.t538 34.8005
R3446 VGND.n851 VGND.t598 34.8005
R3447 VGND.n853 VGND.t546 34.8005
R3448 VGND.n853 VGND.t1622 34.8005
R3449 VGND.n870 VGND.t856 34.8005
R3450 VGND.n870 VGND.t1620 34.8005
R3451 VGND.n875 VGND.t1949 34.8005
R3452 VGND.n875 VGND.t970 34.8005
R3453 VGND.n880 VGND.t2390 34.8005
R3454 VGND.n880 VGND.t594 34.8005
R3455 VGND.n885 VGND.t2501 34.8005
R3456 VGND.n885 VGND.t879 34.8005
R3457 VGND.n890 VGND.t117 34.8005
R3458 VGND.n890 VGND.t968 34.8005
R3459 VGND.n895 VGND.t1568 34.8005
R3460 VGND.n895 VGND.t159 34.8005
R3461 VGND.n900 VGND.t1929 34.8005
R3462 VGND.n900 VGND.t596 34.8005
R3463 VGND.n905 VGND.t620 34.8005
R3464 VGND.n905 VGND.t1618 34.8005
R3465 VGND.n910 VGND.t471 34.8005
R3466 VGND.n910 VGND.t1616 34.8005
R3467 VGND.n915 VGND.t1699 34.8005
R3468 VGND.n915 VGND.t877 34.8005
R3469 VGND.n866 VGND.t1992 34.8005
R3470 VGND.n866 VGND.t875 34.8005
R3471 VGND.n2132 VGND.t1828 34.8005
R3472 VGND.n2132 VGND.t873 34.8005
R3473 VGND.n920 VGND.t1892 34.8005
R3474 VGND.n920 VGND.t157 34.8005
R3475 VGND.n1942 VGND.t1071 34.8005
R3476 VGND.n1942 VGND.t1469 34.8005
R3477 VGND.n1944 VGND.t531 34.8005
R3478 VGND.n1944 VGND.t2185 34.8005
R3479 VGND.n1968 VGND.t2686 34.8005
R3480 VGND.n1968 VGND.t923 34.8005
R3481 VGND.n963 VGND.t862 34.8005
R3482 VGND.n963 VGND.t921 34.8005
R3483 VGND.n1994 VGND.t1943 34.8005
R3484 VGND.n1994 VGND.t1467 34.8005
R3485 VGND.n955 VGND.t883 34.8005
R3486 VGND.n955 VGND.t2181 34.8005
R3487 VGND.n2020 VGND.t2272 34.8005
R3488 VGND.n2020 VGND.t39 34.8005
R3489 VGND.n947 VGND.t111 34.8005
R3490 VGND.n947 VGND.t1465 34.8005
R3491 VGND.n2046 VGND.t2312 34.8005
R3492 VGND.n2046 VGND.t1662 34.8005
R3493 VGND.n939 VGND.t2037 34.8005
R3494 VGND.n939 VGND.t2183 34.8005
R3495 VGND.n2072 VGND.t616 34.8005
R3496 VGND.n2072 VGND.t919 34.8005
R3497 VGND.n931 VGND.t467 34.8005
R3498 VGND.n931 VGND.t1471 34.8005
R3499 VGND.n2103 VGND.t1695 34.8005
R3500 VGND.n2103 VGND.t37 34.8005
R3501 VGND.n2108 VGND.t915 34.8005
R3502 VGND.n2108 VGND.t35 34.8005
R3503 VGND.n2113 VGND.t2475 34.8005
R3504 VGND.n2113 VGND.t925 34.8005
R3505 VGND.n923 VGND.t1888 34.8005
R3506 VGND.n923 VGND.t2187 34.8005
R3507 VGND.n970 VGND.t999 34.8005
R3508 VGND.n970 VGND.t2231 34.8005
R3509 VGND.n1955 VGND.t1518 34.8005
R3510 VGND.n1955 VGND.t2221 34.8005
R3511 VGND.n967 VGND.t1794 34.8005
R3512 VGND.n967 VGND.t1919 34.8005
R3513 VGND.n1981 VGND.t899 34.8005
R3514 VGND.n1981 VGND.t1917 34.8005
R3515 VGND.n959 VGND.t1416 34.8005
R3516 VGND.n959 VGND.t2229 34.8005
R3517 VGND.n2007 VGND.t2072 34.8005
R3518 VGND.n2007 VGND.t2217 34.8005
R3519 VGND.n951 VGND.t754 34.8005
R3520 VGND.n951 VGND.t1691 34.8005
R3521 VGND.n2033 VGND.t2385 34.8005
R3522 VGND.n2033 VGND.t2227 34.8005
R3523 VGND.n943 VGND.t162 34.8005
R3524 VGND.n943 VGND.t2225 34.8005
R3525 VGND.n2059 VGND.t1271 34.8005
R3526 VGND.n2059 VGND.t2219 34.8005
R3527 VGND.n935 VGND.t2583 34.8005
R3528 VGND.n935 VGND.t1915 34.8005
R3529 VGND.n2085 VGND.t1901 34.8005
R3530 VGND.n2085 VGND.t1913 34.8005
R3531 VGND.n927 VGND.t2078 34.8005
R3532 VGND.n927 VGND.t1689 34.8005
R3533 VGND.n2090 VGND.t1931 34.8005
R3534 VGND.n2090 VGND.t1687 34.8005
R3535 VGND.n2680 VGND.t17 34.8005
R3536 VGND.n2680 VGND.t1685 34.8005
R3537 VGND.n590 VGND.t987 34.8005
R3538 VGND.n590 VGND.t2223 34.8005
R3539 VGND.n976 VGND.t1095 34.8005
R3540 VGND.n976 VGND.t784 34.8005
R3541 VGND.n1682 VGND.t1524 34.8005
R3542 VGND.n1682 VGND.t2101 34.8005
R3543 VGND.n1677 VGND.t1813 34.8005
R3544 VGND.n1677 VGND.t792 34.8005
R3545 VGND.n1672 VGND.t70 34.8005
R3546 VGND.n1672 VGND.t790 34.8005
R3547 VGND.n1667 VGND.t1312 34.8005
R3548 VGND.n1667 VGND.t782 34.8005
R3549 VGND.n1662 VGND.t2350 34.8005
R3550 VGND.n1662 VGND.t2097 34.8005
R3551 VGND.n1657 VGND.t778 34.8005
R3552 VGND.n1657 VGND.t2095 34.8005
R3553 VGND.n1652 VGND.t850 34.8005
R3554 VGND.n1652 VGND.t2107 34.8005
R3555 VGND.n1647 VGND.t1320 34.8005
R3556 VGND.n1647 VGND.t2105 34.8005
R3557 VGND.n1642 VGND.t983 34.8005
R3558 VGND.n1642 VGND.t2099 34.8005
R3559 VGND.n1637 VGND.t562 34.8005
R3560 VGND.n1637 VGND.t788 34.8005
R3561 VGND.n1632 VGND.t375 34.8005
R3562 VGND.n1632 VGND.t786 34.8005
R3563 VGND.n1627 VGND.t1994 34.8005
R3564 VGND.n1627 VGND.t2093 34.8005
R3565 VGND.n990 VGND.t434 34.8005
R3566 VGND.n990 VGND.t2091 34.8005
R3567 VGND.n1905 VGND.t2613 34.8005
R3568 VGND.n1905 VGND.t794 34.8005
R3569 VGND.n993 VGND.t905 34.8005
R3570 VGND.n993 VGND.t2103 34.8005
R3571 VGND.n1046 VGND.t1026 34.8005
R3572 VGND.n1046 VGND.t1657 34.8005
R3573 VGND.n1048 VGND.t1607 34.8005
R3574 VGND.n1048 VGND.t1647 34.8005
R3575 VGND.n1741 VGND.t2135 34.8005
R3576 VGND.n1741 VGND.t1295 34.8005
R3577 VGND.n1036 VGND.t2594 34.8005
R3578 VGND.n1036 VGND.t1293 34.8005
R3579 VGND.n1767 VGND.t2407 34.8005
R3580 VGND.n1767 VGND.t1655 34.8005
R3581 VGND.n1028 VGND.t1753 34.8005
R3582 VGND.n1028 VGND.t2442 34.8005
R3583 VGND.n1793 VGND.t2418 34.8005
R3584 VGND.n1793 VGND.t2440 34.8005
R3585 VGND.n1020 VGND.t2492 34.8005
R3586 VGND.n1020 VGND.t1653 34.8005
R3587 VGND.n1819 VGND.t1263 34.8005
R3588 VGND.n1819 VGND.t1651 34.8005
R3589 VGND.n1012 VGND.t2024 34.8005
R3590 VGND.n1012 VGND.t2444 34.8005
R3591 VGND.n1845 VGND.t2015 34.8005
R3592 VGND.n1845 VGND.t1291 34.8005
R3593 VGND.n1004 VGND.t2068 34.8005
R3594 VGND.n1004 VGND.t1289 34.8005
R3595 VGND.n1876 VGND.t2083 34.8005
R3596 VGND.n1876 VGND.t2438 34.8005
R3597 VGND.n1881 VGND.t412 34.8005
R3598 VGND.n1881 VGND.t371 34.8005
R3599 VGND.n1886 VGND.t2001 34.8005
R3600 VGND.n1886 VGND.t1297 34.8005
R3601 VGND.n996 VGND.t2326 34.8005
R3602 VGND.n996 VGND.t1649 34.8005
R3603 VGND.n1043 VGND.t1098 34.8005
R3604 VGND.n1043 VGND.t2657 34.8005
R3605 VGND.n1728 VGND.t1522 34.8005
R3606 VGND.n1728 VGND.t2627 34.8005
R3607 VGND.n1040 VGND.t1811 34.8005
R3608 VGND.n1040 VGND.t426 34.8005
R3609 VGND.n1754 VGND.t72 34.8005
R3610 VGND.n1754 VGND.t424 34.8005
R3611 VGND.n1032 VGND.t1310 34.8005
R3612 VGND.n1032 VGND.t2431 34.8005
R3613 VGND.n1780 VGND.t2348 34.8005
R3614 VGND.n1780 VGND.t2623 34.8005
R3615 VGND.n1024 VGND.t776 34.8005
R3616 VGND.n1024 VGND.t2621 34.8005
R3617 VGND.n1806 VGND.t848 34.8005
R3618 VGND.n1806 VGND.t2429 34.8005
R3619 VGND.n1016 VGND.t1318 34.8005
R3620 VGND.n1016 VGND.t2427 34.8005
R3621 VGND.n1832 VGND.t772 34.8005
R3622 VGND.n1832 VGND.t2625 34.8005
R3623 VGND.n1008 VGND.t560 34.8005
R3624 VGND.n1008 VGND.t422 34.8005
R3625 VGND.n1858 VGND.t373 34.8005
R3626 VGND.n1858 VGND.t420 34.8005
R3627 VGND.n1000 VGND.t1705 34.8005
R3628 VGND.n1000 VGND.t2619 34.8005
R3629 VGND.n1863 VGND.t432 34.8005
R3630 VGND.n1863 VGND.t2617 34.8005
R3631 VGND.n2705 VGND.t2611 34.8005
R3632 VGND.n2705 VGND.t428 34.8005
R3633 VGND.n577 VGND.t903 34.8005
R3634 VGND.n577 VGND.t2629 34.8005
R3635 VGND.n1128 VGND.t1128 34.8005
R3636 VGND.n1128 VGND.t143 34.8005
R3637 VGND.n1131 VGND.t2285 34.8005
R3638 VGND.n1131 VGND.t133 34.8005
R3639 VGND.n1218 VGND.t2146 34.8005
R3640 VGND.n1218 VGND.t2599 34.8005
R3641 VGND.n1235 VGND.t1478 34.8005
R3642 VGND.n1235 VGND.t196 34.8005
R3643 VGND.n1240 VGND.t1422 34.8005
R3644 VGND.n1240 VGND.t141 34.8005
R3645 VGND.n1245 VGND.t359 34.8005
R3646 VGND.n1245 VGND.t2609 34.8005
R3647 VGND.n1250 VGND.t758 34.8005
R3648 VGND.n1250 VGND.t2607 34.8005
R3649 VGND.n1255 VGND.t866 34.8005
R3650 VGND.n1255 VGND.t139 34.8005
R3651 VGND.n1260 VGND.t5 34.8005
R3652 VGND.n1260 VGND.t137 34.8005
R3653 VGND.n1265 VGND.t182 34.8005
R3654 VGND.n1265 VGND.t131 34.8005
R3655 VGND.n1270 VGND.t692 34.8005
R3656 VGND.n1270 VGND.t194 34.8005
R3657 VGND.n1275 VGND.t1905 34.8005
R3658 VGND.n1275 VGND.t192 34.8005
R3659 VGND.n1280 VGND.t2074 34.8005
R3660 VGND.n1280 VGND.t2605 34.8005
R3661 VGND.n1231 VGND.t1937 34.8005
R3662 VGND.n1231 VGND.t2603 34.8005
R3663 VGND.n1293 VGND.t11 34.8005
R3664 VGND.n1293 VGND.t2601 34.8005
R3665 VGND.n1285 VGND.t993 34.8005
R3666 VGND.n1285 VGND.t135 34.8005
R3667 VGND.n54 VGND.t1041 34.8005
R3668 VGND.n54 VGND.t1200 34.8005
R3669 VGND.n292 VGND.t1603 34.8005
R3670 VGND.n292 VGND.t2631 34.8005
R3671 VGND.n287 VGND.t833 34.8005
R3672 VGND.n287 VGND.t1431 34.8005
R3673 VGND.n282 VGND.t800 34.8005
R3674 VGND.n282 VGND.t1429 34.8005
R3675 VGND.n277 VGND.t2402 34.8005
R3676 VGND.n277 VGND.t1198 34.8005
R3677 VGND.n272 VGND.t2261 34.8005
R3678 VGND.n272 VGND.t1956 34.8005
R3679 VGND.n267 VGND.t363 34.8005
R3680 VGND.n267 VGND.t1439 34.8005
R3681 VGND.n262 VGND.t2488 34.8005
R3682 VGND.n262 VGND.t1196 34.8005
R3683 VGND.n257 VGND.t893 34.8005
R3684 VGND.n257 VGND.t1194 34.8005
R3685 VGND.n252 VGND.t2020 34.8005
R3686 VGND.n252 VGND.t1958 34.8005
R3687 VGND.n247 VGND.t2011 34.8005
R3688 VGND.n247 VGND.t1427 34.8005
R3689 VGND.n242 VGND.t2064 34.8005
R3690 VGND.n242 VGND.t1202 34.8005
R3691 VGND.n237 VGND.t128 34.8005
R3692 VGND.n237 VGND.t1437 34.8005
R3693 VGND.n232 VGND.t408 34.8005
R3694 VGND.n232 VGND.t1435 34.8005
R3695 VGND.n227 VGND.t177 34.8005
R3696 VGND.n227 VGND.t1433 34.8005
R3697 VGND.n222 VGND.t2321 34.8005
R3698 VGND.n222 VGND.t1192 34.8005
R3699 VGND.n1057 VGND.t278 34.8005
R3700 VGND.n1057 VGND.t1381 34.8005
R3701 VGND.n1331 VGND.t1552 34.8005
R3702 VGND.n1331 VGND.t280 34.8005
R3703 VGND.n339 VGND.n335 34.6358
R3704 VGND.n1620 VGND.n1052 34.6358
R3705 VGND.n1620 VGND.n1619 34.6358
R3706 VGND.n1619 VGND.n1618 34.6358
R3707 VGND.n1618 VGND.n1606 34.6358
R3708 VGND.n1614 VGND.n1606 34.6358
R3709 VGND.n1600 VGND.n1574 34.6358
R3710 VGND.n1595 VGND.n1575 34.6358
R3711 VGND.n1591 VGND.n1575 34.6358
R3712 VGND.n1591 VGND.n1590 34.6358
R3713 VGND.n1590 VGND.n1589 34.6358
R3714 VGND.n1589 VGND.n1577 34.6358
R3715 VGND.n474 VGND.n469 34.6358
R3716 VGND.n479 VGND.n478 34.6358
R3717 VGND.n824 VGND.n819 34.6358
R3718 VGND.n829 VGND.n828 34.6358
R3719 VGND.n2173 VGND.n2172 34.6358
R3720 VGND.n2181 VGND.n2180 34.6358
R3721 VGND.n2177 VGND.n2176 34.6358
R3722 VGND.n2220 VGND.n844 34.6358
R3723 VGND.n2220 VGND.n2219 34.6358
R3724 VGND.n2219 VGND.n2218 34.6358
R3725 VGND.n2218 VGND.n2204 34.6358
R3726 VGND.n2214 VGND.n2204 34.6358
R3727 VGND.n1692 VGND.n1687 34.6358
R3728 VGND.n1712 VGND.n1688 34.6358
R3729 VGND.n1712 VGND.n1711 34.6358
R3730 VGND.n1711 VGND.n1710 34.6358
R3731 VGND.n1710 VGND.n1696 34.6358
R3732 VGND.n1706 VGND.n1696 34.6358
R3733 VGND.n504 VGND.n499 34.6358
R3734 VGND.n509 VGND.n508 34.6358
R3735 VGND.n114 VGND.n113 34.6358
R3736 VGND.n116 VGND.n107 34.6358
R3737 VGND.n120 VGND.n107 34.6358
R3738 VGND.n121 VGND.n120 34.6358
R3739 VGND.n122 VGND.n121 34.6358
R3740 VGND.n122 VGND.n105 34.6358
R3741 VGND.n310 VGND.n309 34.6358
R3742 VGND.n312 VGND.n301 34.6358
R3743 VGND.n316 VGND.n301 34.6358
R3744 VGND.n317 VGND.n316 34.6358
R3745 VGND.n318 VGND.n317 34.6358
R3746 VGND.n318 VGND.n299 34.6358
R3747 VGND.n438 VGND.n437 34.6358
R3748 VGND.n442 VGND.n441 34.6358
R3749 VGND.n407 VGND.n406 34.6358
R3750 VGND.n411 VGND.n410 34.6358
R3751 VGND.n374 VGND.n373 34.6358
R3752 VGND.n378 VGND.n377 34.6358
R3753 VGND.n343 VGND.n330 34.6358
R3754 VGND.n2889 VGND.n2883 34.6358
R3755 VGND.n2892 VGND.n2891 34.6358
R3756 VGND.n2892 VGND.n2879 34.6358
R3757 VGND.n2896 VGND.n2879 34.6358
R3758 VGND.n2897 VGND.n2896 34.6358
R3759 VGND.n2898 VGND.n2897 34.6358
R3760 VGND.n2914 VGND.n322 34.6358
R3761 VGND.n140 VGND.n134 34.6358
R3762 VGND.n143 VGND.n142 34.6358
R3763 VGND.n143 VGND.n130 34.6358
R3764 VGND.n147 VGND.n130 34.6358
R3765 VGND.n148 VGND.n147 34.6358
R3766 VGND.n149 VGND.n148 34.6358
R3767 VGND.n154 VGND.n153 34.6358
R3768 VGND.n456 VGND.t1165 34.1632
R3769 VGND.n2 VGND.t1166 34.1153
R3770 VGND.n2192 VGND.n846 33.1299
R3771 VGND.n353 VGND.n352 33.1299
R3772 VGND.n346 VGND.n345 32.377
R3773 VGND.n2183 VGND.n2182 32.377
R3774 VGND.n444 VGND.n443 32.377
R3775 VGND.n413 VGND.n412 32.377
R3776 VGND.n380 VGND.n379 32.377
R3777 VGND.n345 VGND.n344 32.377
R3778 VGND.n2183 VGND.n2161 32.0005
R3779 VGND.n457 VGND.n455 32.0005
R3780 VGND.n2858 VGND.n2857 32.0005
R3781 VGND.n485 VGND.n482 30.4946
R3782 VGND.n835 VGND.n832 30.4946
R3783 VGND.n515 VGND.n512 30.4946
R3784 VGND.n447 VGND.n424 29.8709
R3785 VGND.n1612 VGND.n1611 28.9887
R3786 VGND.n1585 VGND.n1584 28.9887
R3787 VGND.n2212 VGND.n2211 28.9887
R3788 VGND.n1704 VGND.n1703 28.9887
R3789 VGND.n115 VGND.n114 27.8593
R3790 VGND.n311 VGND.n310 27.8593
R3791 VGND.n2890 VGND.n2889 27.8593
R3792 VGND.n141 VGND.n140 27.8593
R3793 VGND.n463 VGND.n462 27.0003
R3794 VGND.n418 VGND.n417 26.8591
R3795 VGND.n2180 VGND.n2165 26.3534
R3796 VGND.n441 VGND.n430 26.3534
R3797 VGND.n410 VGND.n399 26.3534
R3798 VGND.n377 VGND.n366 26.3534
R3799 VGND.n337 VGND.n330 26.3534
R3800 VGND.n486 VGND.n485 25.977
R3801 VGND.n836 VGND.n835 25.977
R3802 VGND.n811 VGND.n808 25.977
R3803 VGND.n516 VGND.n515 25.977
R3804 VGND.n386 VGND.n360 25.977
R3805 VGND.n1608 VGND.t486 24.9236
R3806 VGND.n1608 VGND.t1775 24.9236
R3807 VGND.n1610 VGND.t1718 24.9236
R3808 VGND.n1610 VGND.t2364 24.9236
R3809 VGND.n1580 VGND.t1799 24.9236
R3810 VGND.n1580 VGND.t1800 24.9236
R3811 VGND.n1579 VGND.t488 24.9236
R3812 VGND.n1579 VGND.t1777 24.9236
R3813 VGND.n1583 VGND.t2351 24.9236
R3814 VGND.n1583 VGND.t1722 24.9236
R3815 VGND.n1582 VGND.t1719 24.9236
R3816 VGND.n1582 VGND.t2365 24.9236
R3817 VGND.n476 VGND.t1721 24.9236
R3818 VGND.n476 VGND.t669 24.9236
R3819 VGND.n475 VGND.t1780 24.9236
R3820 VGND.n475 VGND.t2525 24.9236
R3821 VGND.n466 VGND.t1276 24.9236
R3822 VGND.n466 VGND.t1716 24.9236
R3823 VGND.n465 VGND.t1987 24.9236
R3824 VGND.n465 VGND.t1771 24.9236
R3825 VGND.n484 VGND.t336 24.9236
R3826 VGND.n484 VGND.t1275 24.9236
R3827 VGND.n483 VGND.t2481 24.9236
R3828 VGND.n483 VGND.t2482 24.9236
R3829 VGND.n826 VGND.t1795 24.9236
R3830 VGND.n826 VGND.t482 24.9236
R3831 VGND.n825 VGND.t672 24.9236
R3832 VGND.n825 VGND.t2353 24.9236
R3833 VGND.n816 VGND.t1285 24.9236
R3834 VGND.n816 VGND.t678 24.9236
R3835 VGND.n815 VGND.t1856 24.9236
R3836 VGND.n815 VGND.t513 24.9236
R3837 VGND.n834 VGND.t1287 24.9236
R3838 VGND.n834 VGND.t1286 24.9236
R3839 VGND.n833 VGND.t1858 24.9236
R3840 VGND.n833 VGND.t1857 24.9236
R3841 VGND.n2163 VGND.t1773 24.9236
R3842 VGND.n2163 VGND.t2522 24.9236
R3843 VGND.n2164 VGND.t1587 24.9236
R3844 VGND.n2164 VGND.t1782 24.9236
R3845 VGND.n2162 VGND.t1591 24.9236
R3846 VGND.n2162 VGND.t1589 24.9236
R3847 VGND.n2167 VGND.t1715 24.9236
R3848 VGND.n2167 VGND.t2362 24.9236
R3849 VGND.n2207 VGND.t490 24.9236
R3850 VGND.n2207 VGND.t1778 24.9236
R3851 VGND.n2206 VGND.t2354 24.9236
R3852 VGND.n2206 VGND.t479 24.9236
R3853 VGND.n2210 VGND.t1720 24.9236
R3854 VGND.n2210 VGND.t688 24.9236
R3855 VGND.n2208 VGND.t1776 24.9236
R3856 VGND.n2208 VGND.t2523 24.9236
R3857 VGND.n1699 VGND.t1723 24.9236
R3858 VGND.n1699 VGND.t1724 24.9236
R3859 VGND.n1698 VGND.t2524 24.9236
R3860 VGND.n1698 VGND.t2359 24.9236
R3861 VGND.n1702 VGND.t2520 24.9236
R3862 VGND.n1702 VGND.t1798 24.9236
R3863 VGND.n1700 VGND.t671 24.9236
R3864 VGND.n1700 VGND.t2352 24.9236
R3865 VGND.n506 VGND.t1797 24.9236
R3866 VGND.n506 VGND.t1770 24.9236
R3867 VGND.n505 VGND.t677 24.9236
R3868 VGND.n505 VGND.t477 24.9236
R3869 VGND.n496 VGND.t1516 24.9236
R3870 VGND.n496 VGND.t1796 24.9236
R3871 VGND.n495 VGND.t717 24.9236
R3872 VGND.n495 VGND.t676 24.9236
R3873 VGND.n514 VGND.t1298 24.9236
R3874 VGND.n514 VGND.t1299 24.9236
R3875 VGND.n513 VGND.t719 24.9236
R3876 VGND.n513 VGND.t718 24.9236
R3877 VGND.n110 VGND.t2567 24.9236
R3878 VGND.n110 VGND.t550 24.9236
R3879 VGND.n109 VGND.t661 24.9236
R3880 VGND.n109 VGND.t523 24.9236
R3881 VGND.n306 VGND.t735 24.9236
R3882 VGND.n306 VGND.t575 24.9236
R3883 VGND.n305 VGND.t525 24.9236
R3884 VGND.n305 VGND.t1844 24.9236
R3885 VGND.n304 VGND.t728 24.9236
R3886 VGND.n304 VGND.t681 24.9236
R3887 VGND.n303 VGND.t515 24.9236
R3888 VGND.n303 VGND.t589 24.9236
R3889 VGND.n433 VGND.t665 24.9236
R3890 VGND.n433 VGND.t1850 24.9236
R3891 VGND.n432 VGND.t730 24.9236
R3892 VGND.n432 VGND.t667 24.9236
R3893 VGND.n429 VGND.t657 24.9236
R3894 VGND.n429 VGND.t60 24.9236
R3895 VGND.n428 VGND.t2575 24.9236
R3896 VGND.n428 VGND.t240 24.9236
R3897 VGND.n427 VGND.t57 24.9236
R3898 VGND.n427 VGND.t63 24.9236
R3899 VGND.n426 VGND.t473 24.9236
R3900 VGND.n426 VGND.t1641 24.9236
R3901 VGND.n402 VGND.t751 24.9236
R3902 VGND.n402 VGND.t2574 24.9236
R3903 VGND.n401 VGND.t585 24.9236
R3904 VGND.n401 VGND.t680 24.9236
R3905 VGND.n398 VGND.t746 24.9236
R3906 VGND.n398 VGND.t955 24.9236
R3907 VGND.n397 VGND.t552 24.9236
R3908 VGND.n397 VGND.t705 24.9236
R3909 VGND.n396 VGND.t954 24.9236
R3910 VGND.n396 VGND.t952 24.9236
R3911 VGND.n395 VGND.t702 24.9236
R3912 VGND.n395 VGND.t708 24.9236
R3913 VGND.n369 VGND.t747 24.9236
R3914 VGND.n369 VGND.t2571 24.9236
R3915 VGND.n368 VGND.t519 24.9236
R3916 VGND.n368 VGND.t732 24.9236
R3917 VGND.n365 VGND.t1851 24.9236
R3918 VGND.n365 VGND.t1260 24.9236
R3919 VGND.n364 VGND.t684 24.9236
R3920 VGND.n364 VGND.t1628 24.9236
R3921 VGND.n363 VGND.t1256 24.9236
R3922 VGND.n363 VGND.t1250 24.9236
R3923 VGND.n362 VGND.t1627 24.9236
R3924 VGND.n362 VGND.t1625 24.9236
R3925 VGND.n329 VGND.t1846 24.9236
R3926 VGND.n329 VGND.t579 24.9236
R3927 VGND.n336 VGND.t738 24.9236
R3928 VGND.n336 VGND.t237 24.9236
R3929 VGND.n328 VGND.t233 24.9236
R3930 VGND.n328 VGND.t227 24.9236
R3931 VGND.n332 VGND.t1849 24.9236
R3932 VGND.n332 VGND.t591 24.9236
R3933 VGND.n2885 VGND.t682 24.9236
R3934 VGND.n2885 VGND.t725 24.9236
R3935 VGND.n2884 VGND.t521 24.9236
R3936 VGND.n2884 VGND.t736 24.9236
R3937 VGND.n2882 VGND.t748 24.9236
R3938 VGND.n2882 VGND.t668 24.9236
R3939 VGND.n2881 VGND.t687 24.9236
R3940 VGND.n2881 VGND.t587 24.9236
R3941 VGND.n136 VGND.t2570 24.9236
R3942 VGND.n136 VGND.t685 24.9236
R3943 VGND.n135 VGND.t727 24.9236
R3944 VGND.n135 VGND.t659 24.9236
R3945 VGND.n133 VGND.t581 24.9236
R3946 VGND.n133 VGND.t734 24.9236
R3947 VGND.n132 VGND.t2573 24.9236
R3948 VGND.n132 VGND.t745 24.9236
R3949 VGND.n486 VGND.n460 24.4711
R3950 VGND.n836 VGND.n807 24.4711
R3951 VGND.n811 VGND.n810 24.4711
R3952 VGND.n2193 VGND.n2192 24.4711
R3953 VGND.n2200 VGND.n843 24.4711
R3954 VGND.n516 VGND.n492 24.4711
R3955 VGND.n444 VGND.n423 24.4711
R3956 VGND.n413 VGND.n392 24.4711
R3957 VGND.n380 VGND.n359 24.4711
R3958 VGND.n386 VGND.n385 24.4711
R3959 VGND.n352 VGND.n349 24.4711
R3960 VGND.n2903 VGND.n2902 24.4711
R3961 VGND.n421 VGND.n393 23.7181
R3962 VGND.n1624 VGND.n1052 23.7181
R3963 VGND.n1596 VGND.n1574 23.7181
R3964 VGND.n1596 VGND.n1595 23.7181
R3965 VGND.n490 VGND.n459 23.7181
R3966 VGND.n2187 VGND.n847 23.7181
R3967 VGND.n2224 VGND.n844 23.7181
R3968 VGND.n1716 VGND.n1687 23.7181
R3969 VGND.n1716 VGND.n1688 23.7181
R3970 VGND.n3005 VGND.n105 23.7181
R3971 VGND.n2915 VGND.n299 23.7181
R3972 VGND.n2898 VGND.n2877 23.7181
R3973 VGND.n2915 VGND.n2914 23.7181
R3974 VGND.n149 VGND.n128 23.7181
R3975 VGND.n153 VGND.n128 23.7181
R3976 VGND.n2188 VGND.n2187 23.3417
R3977 VGND.n357 VGND.n325 23.3417
R3978 VGND.n357 VGND.n326 23.3417
R3979 VGND.n1613 VGND.n1612 21.4593
R3980 VGND.n1585 VGND.n1581 21.4593
R3981 VGND.n2213 VGND.n2212 21.4593
R3982 VGND.n1705 VGND.n1704 21.4593
R3983 VGND.n436 VGND.n435 21.0905
R3984 VGND.n405 VGND.n404 21.0905
R3985 VGND.n372 VGND.n371 21.0905
R3986 VGND.n334 VGND.n333 21.0905
R3987 VGND.n437 VGND.n436 20.3299
R3988 VGND.n406 VGND.n405 20.3299
R3989 VGND.n373 VGND.n372 20.3299
R3990 VGND.n335 VGND.n334 20.3299
R3991 VGND.n482 VGND.n467 19.9534
R3992 VGND.n832 VGND.n817 19.9534
R3993 VGND.n512 VGND.n497 19.9534
R3994 VGND.n2200 VGND.n2199 19.2005
R3995 VGND.n1692 VGND.n1691 19.2005
R3996 VGND.n2904 VGND.n2903 19.2005
R3997 VGND.n2909 VGND.n322 19.2005
R3998 VGND.t2031 VGND.t763 16.8587
R3999 VGND.t959 VGND.t761 16.8587
R4000 VGND.t2526 VGND.t1235 16.8587
R4001 VGND.t2528 VGND.t837 16.8587
R4002 VGND.n1602 VGND.n1601 16.077
R4003 VGND.n156 VGND.n155 16.077
R4004 VGND.n2199 VGND.n2198 15.4358
R4005 VGND.n2905 VGND.n2904 15.4358
R4006 VGND.n462 VGND.n461 14.6829
R4007 VGND.n1691 VGND.n1690 14.6829
R4008 VGND.n417 VGND.n416 14.6829
R4009 VGND.n2910 VGND.n2909 14.6829
R4010 VGND.n471 VGND.n470 14.5711
R4011 VGND.n821 VGND.n820 14.5711
R4012 VGND.n2171 VGND.n2170 14.5711
R4013 VGND.n501 VGND.n500 14.5711
R4014 VGND.n840 VGND.n808 14.3064
R4015 VGND.n390 VGND.n360 14.3064
R4016 VGND.n478 VGND.n477 13.9299
R4017 VGND.n828 VGND.n827 13.9299
R4018 VGND.n2176 VGND.n2168 13.9299
R4019 VGND.n508 VGND.n507 13.9299
R4020 VGND.n2224 VGND.n843 13.5534
R4021 VGND.n2902 VGND.n2877 13.5534
R4022 VGND.n490 VGND.n460 13.177
R4023 VGND.n840 VGND.n807 13.177
R4024 VGND.n520 VGND.n492 13.177
R4025 VGND.n450 VGND.n423 13.177
R4026 VGND.n421 VGND.n392 13.177
R4027 VGND.n390 VGND.n359 13.177
R4028 VGND.n520 VGND.n493 12.8005
R4029 VGND.n450 VGND.n424 12.8005
R4030 VGND.n1601 VGND.n1600 10.5417
R4031 VGND.n155 VGND.n154 10.5417
R4032 VGND.n1690 VGND.n1689 10.0534
R4033 VGND.n2911 VGND.n2910 10.0534
R4034 VGND.n1612 VGND.n1607 9.3005
R4035 VGND.n1615 VGND.n1614 9.3005
R4036 VGND.n1616 VGND.n1606 9.3005
R4037 VGND.n1618 VGND.n1617 9.3005
R4038 VGND.n1619 VGND.n1605 9.3005
R4039 VGND.n1621 VGND.n1620 9.3005
R4040 VGND.n1622 VGND.n1052 9.3005
R4041 VGND.n1624 VGND.n1623 9.3005
R4042 VGND.n1586 VGND.n1585 9.3005
R4043 VGND.n1587 VGND.n1577 9.3005
R4044 VGND.n1589 VGND.n1588 9.3005
R4045 VGND.n1590 VGND.n1576 9.3005
R4046 VGND.n1592 VGND.n1591 9.3005
R4047 VGND.n1593 VGND.n1575 9.3005
R4048 VGND.n1595 VGND.n1594 9.3005
R4049 VGND.n1598 VGND.n1574 9.3005
R4050 VGND.n1600 VGND.n1599 9.3005
R4051 VGND.n1597 VGND.n1596 9.3005
R4052 VGND.n488 VGND.n460 9.3005
R4053 VGND.n472 VGND.n469 9.3005
R4054 VGND.n474 VGND.n473 9.3005
R4055 VGND.n478 VGND.n468 9.3005
R4056 VGND.n480 VGND.n479 9.3005
R4057 VGND.n482 VGND.n481 9.3005
R4058 VGND.n485 VGND.n464 9.3005
R4059 VGND.n487 VGND.n486 9.3005
R4060 VGND.n463 VGND.n459 9.3005
R4061 VGND.n490 VGND.n489 9.3005
R4062 VGND.n810 VGND.n809 9.3005
R4063 VGND.n813 VGND.n808 9.3005
R4064 VGND.n838 VGND.n807 9.3005
R4065 VGND.n822 VGND.n819 9.3005
R4066 VGND.n824 VGND.n823 9.3005
R4067 VGND.n828 VGND.n818 9.3005
R4068 VGND.n830 VGND.n829 9.3005
R4069 VGND.n832 VGND.n831 9.3005
R4070 VGND.n835 VGND.n814 9.3005
R4071 VGND.n837 VGND.n836 9.3005
R4072 VGND.n812 VGND.n811 9.3005
R4073 VGND.n840 VGND.n839 9.3005
R4074 VGND.n2194 VGND.n2193 9.3005
R4075 VGND.n2185 VGND.n847 9.3005
R4076 VGND.n2172 VGND.n2169 9.3005
R4077 VGND.n2174 VGND.n2173 9.3005
R4078 VGND.n2176 VGND.n2175 9.3005
R4079 VGND.n2178 VGND.n2177 9.3005
R4080 VGND.n2180 VGND.n2179 9.3005
R4081 VGND.n2181 VGND.n2160 9.3005
R4082 VGND.n2184 VGND.n2183 9.3005
R4083 VGND.n2190 VGND.n2189 9.3005
R4084 VGND.n2192 VGND.n2191 9.3005
R4085 VGND.n2187 VGND.n2186 9.3005
R4086 VGND.n2212 VGND.n2205 9.3005
R4087 VGND.n2215 VGND.n2214 9.3005
R4088 VGND.n2216 VGND.n2204 9.3005
R4089 VGND.n2218 VGND.n2217 9.3005
R4090 VGND.n2219 VGND.n2203 9.3005
R4091 VGND.n2221 VGND.n2220 9.3005
R4092 VGND.n2222 VGND.n844 9.3005
R4093 VGND.n2202 VGND.n843 9.3005
R4094 VGND.n2201 VGND.n2200 9.3005
R4095 VGND.n2198 VGND.n2197 9.3005
R4096 VGND.n2224 VGND.n2223 9.3005
R4097 VGND.n1704 VGND.n1697 9.3005
R4098 VGND.n1707 VGND.n1706 9.3005
R4099 VGND.n1708 VGND.n1696 9.3005
R4100 VGND.n1710 VGND.n1709 9.3005
R4101 VGND.n1711 VGND.n1695 9.3005
R4102 VGND.n1713 VGND.n1712 9.3005
R4103 VGND.n1714 VGND.n1688 9.3005
R4104 VGND.n1694 VGND.n1687 9.3005
R4105 VGND.n1693 VGND.n1692 9.3005
R4106 VGND.n1716 VGND.n1715 9.3005
R4107 VGND.n518 VGND.n492 9.3005
R4108 VGND.n502 VGND.n499 9.3005
R4109 VGND.n504 VGND.n503 9.3005
R4110 VGND.n508 VGND.n498 9.3005
R4111 VGND.n510 VGND.n509 9.3005
R4112 VGND.n512 VGND.n511 9.3005
R4113 VGND.n515 VGND.n494 9.3005
R4114 VGND.n517 VGND.n516 9.3005
R4115 VGND.n520 VGND.n519 9.3005
R4116 VGND.n3005 VGND.n3004 9.3005
R4117 VGND.n113 VGND.n112 9.3005
R4118 VGND.n114 VGND.n108 9.3005
R4119 VGND.n117 VGND.n116 9.3005
R4120 VGND.n118 VGND.n107 9.3005
R4121 VGND.n120 VGND.n119 9.3005
R4122 VGND.n121 VGND.n106 9.3005
R4123 VGND.n123 VGND.n122 9.3005
R4124 VGND.n124 VGND.n105 9.3005
R4125 VGND.n448 VGND.n424 9.3005
R4126 VGND.n437 VGND.n431 9.3005
R4127 VGND.n439 VGND.n438 9.3005
R4128 VGND.n441 VGND.n440 9.3005
R4129 VGND.n442 VGND.n425 9.3005
R4130 VGND.n445 VGND.n444 9.3005
R4131 VGND.n446 VGND.n423 9.3005
R4132 VGND.n450 VGND.n449 9.3005
R4133 VGND.n419 VGND.n393 9.3005
R4134 VGND.n406 VGND.n400 9.3005
R4135 VGND.n408 VGND.n407 9.3005
R4136 VGND.n410 VGND.n409 9.3005
R4137 VGND.n411 VGND.n394 9.3005
R4138 VGND.n414 VGND.n413 9.3005
R4139 VGND.n415 VGND.n392 9.3005
R4140 VGND.n421 VGND.n420 9.3005
R4141 VGND.n385 VGND.n384 9.3005
R4142 VGND.n373 VGND.n367 9.3005
R4143 VGND.n375 VGND.n374 9.3005
R4144 VGND.n377 VGND.n376 9.3005
R4145 VGND.n378 VGND.n361 9.3005
R4146 VGND.n381 VGND.n380 9.3005
R4147 VGND.n382 VGND.n359 9.3005
R4148 VGND.n388 VGND.n360 9.3005
R4149 VGND.n387 VGND.n386 9.3005
R4150 VGND.n390 VGND.n389 9.3005
R4151 VGND.n350 VGND.n349 9.3005
R4152 VGND.n335 VGND.n331 9.3005
R4153 VGND.n340 VGND.n339 9.3005
R4154 VGND.n341 VGND.n330 9.3005
R4155 VGND.n343 VGND.n342 9.3005
R4156 VGND.n345 VGND.n327 9.3005
R4157 VGND.n348 VGND.n347 9.3005
R4158 VGND.n355 VGND.n354 9.3005
R4159 VGND.n352 VGND.n351 9.3005
R4160 VGND.n357 VGND.n356 9.3005
R4161 VGND.n2906 VGND.n2905 9.3005
R4162 VGND.n2887 VGND.n2883 9.3005
R4163 VGND.n2889 VGND.n2888 9.3005
R4164 VGND.n2891 VGND.n2880 9.3005
R4165 VGND.n2893 VGND.n2892 9.3005
R4166 VGND.n2894 VGND.n2879 9.3005
R4167 VGND.n2896 VGND.n2895 9.3005
R4168 VGND.n2897 VGND.n2878 9.3005
R4169 VGND.n2899 VGND.n2898 9.3005
R4170 VGND.n2902 VGND.n2901 9.3005
R4171 VGND.n2903 VGND.n324 9.3005
R4172 VGND.n2900 VGND.n2877 9.3005
R4173 VGND.n309 VGND.n308 9.3005
R4174 VGND.n310 VGND.n302 9.3005
R4175 VGND.n313 VGND.n312 9.3005
R4176 VGND.n314 VGND.n301 9.3005
R4177 VGND.n316 VGND.n315 9.3005
R4178 VGND.n317 VGND.n300 9.3005
R4179 VGND.n319 VGND.n318 9.3005
R4180 VGND.n320 VGND.n299 9.3005
R4181 VGND.n2915 VGND.n321 9.3005
R4182 VGND.n2914 VGND.n2913 9.3005
R4183 VGND.n2912 VGND.n322 9.3005
R4184 VGND.n138 VGND.n134 9.3005
R4185 VGND.n140 VGND.n139 9.3005
R4186 VGND.n142 VGND.n131 9.3005
R4187 VGND.n144 VGND.n143 9.3005
R4188 VGND.n145 VGND.n130 9.3005
R4189 VGND.n147 VGND.n146 9.3005
R4190 VGND.n148 VGND.n129 9.3005
R4191 VGND.n150 VGND.n149 9.3005
R4192 VGND.n151 VGND.n128 9.3005
R4193 VGND.n153 VGND.n152 9.3005
R4194 VGND.n154 VGND.n125 9.3005
R4195 VGND.n438 VGND.n430 8.28285
R4196 VGND.n407 VGND.n399 8.28285
R4197 VGND.n374 VGND.n366 8.28285
R4198 VGND.n1207 VGND.n1136 7.9105
R4199 VGND.n528 VGND.n524 7.9105
R4200 VGND.n2843 VGND.n2842 7.9105
R4201 VGND.n2841 VGND.n532 7.9105
R4202 VGND.n2840 VGND.n533 7.9105
R4203 VGND.n2839 VGND.n534 7.9105
R4204 VGND.n2838 VGND.n535 7.9105
R4205 VGND.n2837 VGND.n536 7.9105
R4206 VGND.n2836 VGND.n537 7.9105
R4207 VGND.n2835 VGND.n538 7.9105
R4208 VGND.n2834 VGND.n539 7.9105
R4209 VGND.n2833 VGND.n540 7.9105
R4210 VGND.n2832 VGND.n541 7.9105
R4211 VGND.n2831 VGND.n542 7.9105
R4212 VGND.n2830 VGND.n543 7.9105
R4213 VGND.n2829 VGND.n544 7.9105
R4214 VGND.n2828 VGND.n2827 7.9105
R4215 VGND.n2450 VGND.n2449 7.9105
R4216 VGND.n2467 VGND.n2466 7.9105
R4217 VGND.n2476 VGND.n2475 7.9105
R4218 VGND.n2493 VGND.n2492 7.9105
R4219 VGND.n2502 VGND.n2501 7.9105
R4220 VGND.n2519 VGND.n2518 7.9105
R4221 VGND.n2528 VGND.n2527 7.9105
R4222 VGND.n2545 VGND.n2544 7.9105
R4223 VGND.n2554 VGND.n2553 7.9105
R4224 VGND.n2571 VGND.n2570 7.9105
R4225 VGND.n2580 VGND.n2579 7.9105
R4226 VGND.n2602 VGND.n2601 7.9105
R4227 VGND.n2624 VGND.n615 7.9105
R4228 VGND.n2623 VGND.n616 7.9105
R4229 VGND.n2621 VGND.n2620 7.9105
R4230 VGND.n2757 VGND.n2756 7.9105
R4231 VGND.n2454 VGND.n2453 7.9105
R4232 VGND.n2463 VGND.n2462 7.9105
R4233 VGND.n2480 VGND.n2479 7.9105
R4234 VGND.n2489 VGND.n2488 7.9105
R4235 VGND.n2506 VGND.n2505 7.9105
R4236 VGND.n2515 VGND.n2514 7.9105
R4237 VGND.n2532 VGND.n2531 7.9105
R4238 VGND.n2541 VGND.n2540 7.9105
R4239 VGND.n2558 VGND.n2557 7.9105
R4240 VGND.n2567 VGND.n2566 7.9105
R4241 VGND.n2584 VGND.n2583 7.9105
R4242 VGND.n2598 VGND.n2597 7.9105
R4243 VGND.n2627 VGND.n614 7.9105
R4244 VGND.n2629 VGND.n2628 7.9105
R4245 VGND.n2641 VGND.n611 7.9105
R4246 VGND.n2640 VGND.n2639 7.9105
R4247 VGND.n2434 VGND.n672 7.9105
R4248 VGND.n2433 VGND.n673 7.9105
R4249 VGND.n2432 VGND.n674 7.9105
R4250 VGND.n2431 VGND.n675 7.9105
R4251 VGND.n2430 VGND.n676 7.9105
R4252 VGND.n2429 VGND.n677 7.9105
R4253 VGND.n2428 VGND.n678 7.9105
R4254 VGND.n2427 VGND.n679 7.9105
R4255 VGND.n2426 VGND.n680 7.9105
R4256 VGND.n2425 VGND.n681 7.9105
R4257 VGND.n2424 VGND.n682 7.9105
R4258 VGND.n2423 VGND.n683 7.9105
R4259 VGND.n2422 VGND.n2421 7.9105
R4260 VGND.n2645 VGND.n608 7.9105
R4261 VGND.n2644 VGND.n609 7.9105
R4262 VGND.n2409 VGND.n2408 7.9105
R4263 VGND.n2232 VGND.n2231 7.9105
R4264 VGND.n2249 VGND.n2248 7.9105
R4265 VGND.n2258 VGND.n2257 7.9105
R4266 VGND.n2275 VGND.n2274 7.9105
R4267 VGND.n2284 VGND.n2283 7.9105
R4268 VGND.n2301 VGND.n2300 7.9105
R4269 VGND.n2310 VGND.n2309 7.9105
R4270 VGND.n2327 VGND.n2326 7.9105
R4271 VGND.n2336 VGND.n2335 7.9105
R4272 VGND.n2353 VGND.n2352 7.9105
R4273 VGND.n2362 VGND.n2361 7.9105
R4274 VGND.n2384 VGND.n2383 7.9105
R4275 VGND.n2649 VGND.n605 7.9105
R4276 VGND.n2648 VGND.n606 7.9105
R4277 VGND.n753 VGND.n752 7.9105
R4278 VGND.n2405 VGND.n2404 7.9105
R4279 VGND.n2236 VGND.n2235 7.9105
R4280 VGND.n2245 VGND.n2244 7.9105
R4281 VGND.n2262 VGND.n2261 7.9105
R4282 VGND.n2271 VGND.n2270 7.9105
R4283 VGND.n2288 VGND.n2287 7.9105
R4284 VGND.n2297 VGND.n2296 7.9105
R4285 VGND.n2314 VGND.n2313 7.9105
R4286 VGND.n2323 VGND.n2322 7.9105
R4287 VGND.n2340 VGND.n2339 7.9105
R4288 VGND.n2349 VGND.n2348 7.9105
R4289 VGND.n2366 VGND.n2365 7.9105
R4290 VGND.n2380 VGND.n2379 7.9105
R4291 VGND.n2652 VGND.n603 7.9105
R4292 VGND.n2654 VGND.n2653 7.9105
R4293 VGND.n2666 VGND.n599 7.9105
R4294 VGND.n2665 VGND.n2664 7.9105
R4295 VGND.n1937 VGND.n850 7.9105
R4296 VGND.n2152 VGND.n2151 7.9105
R4297 VGND.n2150 VGND.n856 7.9105
R4298 VGND.n2149 VGND.n857 7.9105
R4299 VGND.n2148 VGND.n858 7.9105
R4300 VGND.n2147 VGND.n859 7.9105
R4301 VGND.n2146 VGND.n860 7.9105
R4302 VGND.n2145 VGND.n861 7.9105
R4303 VGND.n2144 VGND.n862 7.9105
R4304 VGND.n2143 VGND.n863 7.9105
R4305 VGND.n2142 VGND.n864 7.9105
R4306 VGND.n2141 VGND.n865 7.9105
R4307 VGND.n2140 VGND.n2139 7.9105
R4308 VGND.n2670 VGND.n596 7.9105
R4309 VGND.n2669 VGND.n597 7.9105
R4310 VGND.n2127 VGND.n2126 7.9105
R4311 VGND.n1950 VGND.n1949 7.9105
R4312 VGND.n1967 VGND.n1966 7.9105
R4313 VGND.n1976 VGND.n1975 7.9105
R4314 VGND.n1993 VGND.n1992 7.9105
R4315 VGND.n2002 VGND.n2001 7.9105
R4316 VGND.n2019 VGND.n2018 7.9105
R4317 VGND.n2028 VGND.n2027 7.9105
R4318 VGND.n2045 VGND.n2044 7.9105
R4319 VGND.n2054 VGND.n2053 7.9105
R4320 VGND.n2071 VGND.n2070 7.9105
R4321 VGND.n2080 VGND.n2079 7.9105
R4322 VGND.n2102 VGND.n2101 7.9105
R4323 VGND.n2674 VGND.n593 7.9105
R4324 VGND.n2673 VGND.n594 7.9105
R4325 VGND.n925 VGND.n924 7.9105
R4326 VGND.n2123 VGND.n2122 7.9105
R4327 VGND.n1954 VGND.n1953 7.9105
R4328 VGND.n1963 VGND.n1962 7.9105
R4329 VGND.n1980 VGND.n1979 7.9105
R4330 VGND.n1989 VGND.n1988 7.9105
R4331 VGND.n2006 VGND.n2005 7.9105
R4332 VGND.n2015 VGND.n2014 7.9105
R4333 VGND.n2032 VGND.n2031 7.9105
R4334 VGND.n2041 VGND.n2040 7.9105
R4335 VGND.n2058 VGND.n2057 7.9105
R4336 VGND.n2067 VGND.n2066 7.9105
R4337 VGND.n2084 VGND.n2083 7.9105
R4338 VGND.n2098 VGND.n2097 7.9105
R4339 VGND.n2677 VGND.n591 7.9105
R4340 VGND.n2679 VGND.n2678 7.9105
R4341 VGND.n2691 VGND.n587 7.9105
R4342 VGND.n2690 VGND.n2689 7.9105
R4343 VGND.n1925 VGND.n978 7.9105
R4344 VGND.n1924 VGND.n979 7.9105
R4345 VGND.n1923 VGND.n980 7.9105
R4346 VGND.n1922 VGND.n981 7.9105
R4347 VGND.n1921 VGND.n982 7.9105
R4348 VGND.n1920 VGND.n983 7.9105
R4349 VGND.n1919 VGND.n984 7.9105
R4350 VGND.n1918 VGND.n985 7.9105
R4351 VGND.n1917 VGND.n986 7.9105
R4352 VGND.n1916 VGND.n987 7.9105
R4353 VGND.n1915 VGND.n988 7.9105
R4354 VGND.n1914 VGND.n989 7.9105
R4355 VGND.n1913 VGND.n1912 7.9105
R4356 VGND.n2695 VGND.n584 7.9105
R4357 VGND.n2694 VGND.n585 7.9105
R4358 VGND.n1900 VGND.n1899 7.9105
R4359 VGND.n1723 VGND.n1722 7.9105
R4360 VGND.n1740 VGND.n1739 7.9105
R4361 VGND.n1749 VGND.n1748 7.9105
R4362 VGND.n1766 VGND.n1765 7.9105
R4363 VGND.n1775 VGND.n1774 7.9105
R4364 VGND.n1792 VGND.n1791 7.9105
R4365 VGND.n1801 VGND.n1800 7.9105
R4366 VGND.n1818 VGND.n1817 7.9105
R4367 VGND.n1827 VGND.n1826 7.9105
R4368 VGND.n1844 VGND.n1843 7.9105
R4369 VGND.n1853 VGND.n1852 7.9105
R4370 VGND.n1875 VGND.n1874 7.9105
R4371 VGND.n2699 VGND.n581 7.9105
R4372 VGND.n2698 VGND.n582 7.9105
R4373 VGND.n998 VGND.n997 7.9105
R4374 VGND.n1896 VGND.n1895 7.9105
R4375 VGND.n1727 VGND.n1726 7.9105
R4376 VGND.n1736 VGND.n1735 7.9105
R4377 VGND.n1753 VGND.n1752 7.9105
R4378 VGND.n1762 VGND.n1761 7.9105
R4379 VGND.n1779 VGND.n1778 7.9105
R4380 VGND.n1788 VGND.n1787 7.9105
R4381 VGND.n1805 VGND.n1804 7.9105
R4382 VGND.n1814 VGND.n1813 7.9105
R4383 VGND.n1831 VGND.n1830 7.9105
R4384 VGND.n1840 VGND.n1839 7.9105
R4385 VGND.n1857 VGND.n1856 7.9105
R4386 VGND.n1871 VGND.n1870 7.9105
R4387 VGND.n2702 VGND.n578 7.9105
R4388 VGND.n2704 VGND.n2703 7.9105
R4389 VGND.n2716 VGND.n574 7.9105
R4390 VGND.n2715 VGND.n2714 7.9105
R4391 VGND.n1217 VGND.n1130 7.9105
R4392 VGND.n1313 VGND.n1312 7.9105
R4393 VGND.n1311 VGND.n1221 7.9105
R4394 VGND.n1310 VGND.n1222 7.9105
R4395 VGND.n1309 VGND.n1223 7.9105
R4396 VGND.n1308 VGND.n1224 7.9105
R4397 VGND.n1307 VGND.n1225 7.9105
R4398 VGND.n1306 VGND.n1226 7.9105
R4399 VGND.n1305 VGND.n1227 7.9105
R4400 VGND.n1304 VGND.n1228 7.9105
R4401 VGND.n1303 VGND.n1229 7.9105
R4402 VGND.n1302 VGND.n1230 7.9105
R4403 VGND.n1301 VGND.n1300 7.9105
R4404 VGND.n2720 VGND.n569 7.9105
R4405 VGND.n2719 VGND.n570 7.9105
R4406 VGND.n1288 VGND.n1287 7.9105
R4407 VGND.n3055 VGND.n56 7.9105
R4408 VGND.n3054 VGND.n57 7.9105
R4409 VGND.n3049 VGND.n62 7.9105
R4410 VGND.n3048 VGND.n63 7.9105
R4411 VGND.n3043 VGND.n68 7.9105
R4412 VGND.n3042 VGND.n69 7.9105
R4413 VGND.n3037 VGND.n74 7.9105
R4414 VGND.n3036 VGND.n75 7.9105
R4415 VGND.n3031 VGND.n80 7.9105
R4416 VGND.n3030 VGND.n81 7.9105
R4417 VGND.n3025 VGND.n86 7.9105
R4418 VGND.n3024 VGND.n87 7.9105
R4419 VGND.n3019 VGND.n92 7.9105
R4420 VGND.n3018 VGND.n93 7.9105
R4421 VGND.n3013 VGND.n98 7.9105
R4422 VGND.n3012 VGND.n3011 7.9105
R4423 VGND.n1205 VGND.n1137 7.9105
R4424 VGND.n1204 VGND.n1203 7.9105
R4425 VGND.n1554 VGND.n1071 7.9105
R4426 VGND.n1553 VGND.n1072 7.9105
R4427 VGND.n1546 VGND.n1077 7.9105
R4428 VGND.n1545 VGND.n1078 7.9105
R4429 VGND.n1538 VGND.n1083 7.9105
R4430 VGND.n1537 VGND.n1084 7.9105
R4431 VGND.n1530 VGND.n1089 7.9105
R4432 VGND.n1529 VGND.n1090 7.9105
R4433 VGND.n1522 VGND.n1095 7.9105
R4434 VGND.n1521 VGND.n1096 7.9105
R4435 VGND.n2724 VGND.n2723 7.9105
R4436 VGND.n571 VGND.n566 7.9105
R4437 VGND.n2735 VGND.n2734 7.9105
R4438 VGND.n1325 VGND.n1324 7.9105
R4439 VGND.n1399 VGND.n1398 7.9105
R4440 VGND.n1558 VGND.n1068 7.9105
R4441 VGND.n1557 VGND.n1069 7.9105
R4442 VGND.n1550 VGND.n1074 7.9105
R4443 VGND.n1549 VGND.n1075 7.9105
R4444 VGND.n1542 VGND.n1080 7.9105
R4445 VGND.n1541 VGND.n1081 7.9105
R4446 VGND.n1534 VGND.n1086 7.9105
R4447 VGND.n1533 VGND.n1087 7.9105
R4448 VGND.n1526 VGND.n1092 7.9105
R4449 VGND.n1525 VGND.n1093 7.9105
R4450 VGND.n1518 VGND.n1098 7.9105
R4451 VGND.n1517 VGND.n1099 7.9105
R4452 VGND.n1516 VGND.n1100 7.9105
R4453 VGND.n2739 VGND.n2738 7.9105
R4454 VGND.n477 VGND.n474 7.90638
R4455 VGND.n470 VGND.n469 7.90638
R4456 VGND.n827 VGND.n824 7.90638
R4457 VGND.n820 VGND.n819 7.90638
R4458 VGND.n2173 VGND.n2168 7.90638
R4459 VGND.n2172 VGND.n2171 7.90638
R4460 VGND.n507 VGND.n504 7.90638
R4461 VGND.n500 VGND.n499 7.90638
R4462 VGND.n1611 VGND.n1609 7.4049
R4463 VGND.n1584 VGND.n1578 7.4049
R4464 VGND.n2211 VGND.n2209 7.4049
R4465 VGND.n1703 VGND.n1701 7.4049
R4466 VGND VGND.n493 7.12482
R4467 VGND.n435 VGND.n434 6.85473
R4468 VGND.n404 VGND.n403 6.85473
R4469 VGND.n371 VGND.n370 6.85473
R4470 VGND.n116 VGND.n115 6.77697
R4471 VGND.n312 VGND.n311 6.77697
R4472 VGND.n2891 VGND.n2890 6.77697
R4473 VGND.n142 VGND.n141 6.77697
R4474 VGND.n2166 VGND.n2165 5.27109
R4475 VGND.n338 VGND.n337 5.27109
R4476 VGND.n161 VGND.n160 4.5005
R4477 VGND.n164 VGND.n163 4.5005
R4478 VGND.n167 VGND.n166 4.5005
R4479 VGND.n170 VGND.n169 4.5005
R4480 VGND.n173 VGND.n172 4.5005
R4481 VGND.n176 VGND.n175 4.5005
R4482 VGND.n179 VGND.n178 4.5005
R4483 VGND.n182 VGND.n181 4.5005
R4484 VGND.n185 VGND.n184 4.5005
R4485 VGND.n188 VGND.n187 4.5005
R4486 VGND.n191 VGND.n190 4.5005
R4487 VGND.n194 VGND.n193 4.5005
R4488 VGND.n197 VGND.n196 4.5005
R4489 VGND.n200 VGND.n199 4.5005
R4490 VGND.n205 VGND.n96 4.5005
R4491 VGND.n2989 VGND.n95 4.5005
R4492 VGND.n207 VGND.n90 4.5005
R4493 VGND.n2979 VGND.n89 4.5005
R4494 VGND.n209 VGND.n84 4.5005
R4495 VGND.n2969 VGND.n83 4.5005
R4496 VGND.n211 VGND.n78 4.5005
R4497 VGND.n2959 VGND.n77 4.5005
R4498 VGND.n213 VGND.n72 4.5005
R4499 VGND.n2949 VGND.n71 4.5005
R4500 VGND.n215 VGND.n66 4.5005
R4501 VGND.n2939 VGND.n65 4.5005
R4502 VGND.n217 VGND.n60 4.5005
R4503 VGND.n2929 VGND.n59 4.5005
R4504 VGND.n8 VGND.n7 4.5005
R4505 VGND.n11 VGND.n10 4.5005
R4506 VGND.n14 VGND.n13 4.5005
R4507 VGND.n17 VGND.n16 4.5005
R4508 VGND.n20 VGND.n19 4.5005
R4509 VGND.n23 VGND.n22 4.5005
R4510 VGND.n26 VGND.n25 4.5005
R4511 VGND.n29 VGND.n28 4.5005
R4512 VGND.n32 VGND.n31 4.5005
R4513 VGND.n35 VGND.n34 4.5005
R4514 VGND.n38 VGND.n37 4.5005
R4515 VGND.n41 VGND.n40 4.5005
R4516 VGND.n44 VGND.n43 4.5005
R4517 VGND.n47 VGND.n46 4.5005
R4518 VGND.n50 VGND.n49 4.5005
R4519 VGND.n221 VGND.n52 4.5005
R4520 VGND.n159 VGND.n158 4.5005
R4521 VGND.n203 VGND.n202 4.5005
R4522 VGND.n3000 VGND.n2999 4.5005
R4523 VGND.n1403 VGND.n1123 4.5005
R4524 VGND.n1066 VGND.n1065 4.5005
R4525 VGND.n1416 VGND.n1415 4.5005
R4526 VGND.n1428 VGND.n1407 4.5005
R4527 VGND.n1435 VGND.n1122 4.5005
R4528 VGND.n1432 VGND.n1430 4.5005
R4529 VGND.n1448 VGND.n1447 4.5005
R4530 VGND.n1460 VGND.n1116 4.5005
R4531 VGND.n1467 VGND.n1114 4.5005
R4532 VGND.n1464 VGND.n1462 4.5005
R4533 VGND.n1480 VGND.n1479 4.5005
R4534 VGND.n1492 VGND.n1108 4.5005
R4535 VGND.n1498 VGND.n1106 4.5005
R4536 VGND.n1495 VGND.n1494 4.5005
R4537 VGND.n1103 VGND.n1102 4.5005
R4538 VGND.n1056 VGND.n1055 4.5005
R4539 VGND.n1570 VGND.n1569 4.5005
R4540 VGND.n1402 VGND.n1062 4.5005
R4541 VGND.n1562 VGND.n1561 4.5005
R4542 VGND.n1418 VGND.n1417 4.5005
R4543 VGND.n1427 VGND.n1426 4.5005
R4544 VGND.n1437 VGND.n1436 4.5005
R4545 VGND.n1431 VGND.n1121 4.5005
R4546 VGND.n1450 VGND.n1449 4.5005
R4547 VGND.n1459 VGND.n1458 4.5005
R4548 VGND.n1469 VGND.n1468 4.5005
R4549 VGND.n1463 VGND.n1113 4.5005
R4550 VGND.n1482 VGND.n1481 4.5005
R4551 VGND.n1491 VGND.n1490 4.5005
R4552 VGND.n1501 VGND.n1500 4.5005
R4553 VGND.n1105 VGND.n1101 4.5005
R4554 VGND.n1512 VGND.n1511 4.5005
R4555 VGND.n1623 VGND.n1604 4.41365
R4556 VGND VGND.n3003 4.35375
R4557 VGND.n1603 VGND.n1602 4.05427
R4558 VGND.n809 VGND.n0 4.05427
R4559 VGND.n2195 VGND.n2194 4.05427
R4560 VGND.n2197 VGND.n2196 4.05427
R4561 VGND.n1689 VGND.n845 4.05427
R4562 VGND VGND.n383 3.99438
R4563 VGND VGND.n323 3.99438
R4564 VGND.n2907 VGND 3.99438
R4565 VGND VGND.n2908 3.99437
R4566 VGND.n157 VGND 3.99437
R4567 VGND.n1513 VGND.n561 3.77268
R4568 VGND.n3001 VGND.n99 3.77268
R4569 VGND.n1571 VGND.n1054 3.77268
R4570 VGND.n3057 VGND.n3056 3.77268
R4571 VGND.n1560 VGND.n1559 3.77268
R4572 VGND.n3051 VGND.n3050 3.77268
R4573 VGND.n1556 VGND.n1070 3.77268
R4574 VGND.n3047 VGND.n3046 3.77268
R4575 VGND.n1551 VGND.n1073 3.77268
R4576 VGND.n3045 VGND.n3044 3.77268
R4577 VGND.n1548 VGND.n1076 3.77268
R4578 VGND.n3041 VGND.n3040 3.77268
R4579 VGND.n1543 VGND.n1079 3.77268
R4580 VGND.n3039 VGND.n3038 3.77268
R4581 VGND.n1540 VGND.n1082 3.77268
R4582 VGND.n3035 VGND.n3034 3.77268
R4583 VGND.n1535 VGND.n1085 3.77268
R4584 VGND.n3033 VGND.n3032 3.77268
R4585 VGND.n1532 VGND.n1088 3.77268
R4586 VGND.n3029 VGND.n3028 3.77268
R4587 VGND.n1527 VGND.n1091 3.77268
R4588 VGND.n3027 VGND.n3026 3.77268
R4589 VGND.n1524 VGND.n1094 3.77268
R4590 VGND.n3023 VGND.n3022 3.77268
R4591 VGND.n1519 VGND.n1097 3.77268
R4592 VGND.n3021 VGND.n3020 3.77268
R4593 VGND.n1499 VGND.n567 3.77268
R4594 VGND.n3017 VGND.n3016 3.77268
R4595 VGND.n1515 VGND.n1514 3.77268
R4596 VGND.n3015 VGND.n3014 3.77268
R4597 VGND.n1401 VGND.n1400 3.77268
R4598 VGND.n3053 VGND.n3052 3.77268
R4599 VGND.n1208 VGND.n1133 3.76865
R4600 VGND.n162 VGND.n159 3.75914
R4601 VGND.n203 VGND.n201 3.75914
R4602 VGND.n1496 VGND.n1103 3.75914
R4603 VGND.n1404 VGND.n1056 3.75914
R4604 VGND.n527 VGND.n4 3.49421
R4605 VGND.n2441 VGND.n667 3.49421
R4606 VGND.n2438 VGND.n2437 3.49421
R4607 VGND.n2436 VGND.n2435 3.49421
R4608 VGND.n1931 VGND.n669 3.49421
R4609 VGND.n1935 VGND.n1934 3.49421
R4610 VGND.n1938 VGND.n1936 3.49421
R4611 VGND.n1941 VGND.n973 3.49421
R4612 VGND.n1929 VGND.n1928 3.49421
R4613 VGND.n1927 VGND.n1926 3.49421
R4614 VGND.n1210 VGND.n975 3.49421
R4615 VGND.n1213 VGND.n1212 3.49421
R4616 VGND.n1216 VGND.n1133 3.49421
R4617 VGND.n3061 VGND.n3060 3.49421
R4618 VGND.n162 VGND.n161 3.4105
R4619 VGND.n165 VGND.n164 3.4105
R4620 VGND.n168 VGND.n167 3.4105
R4621 VGND.n171 VGND.n170 3.4105
R4622 VGND.n174 VGND.n173 3.4105
R4623 VGND.n177 VGND.n176 3.4105
R4624 VGND.n180 VGND.n179 3.4105
R4625 VGND.n183 VGND.n182 3.4105
R4626 VGND.n186 VGND.n185 3.4105
R4627 VGND.n189 VGND.n188 3.4105
R4628 VGND.n192 VGND.n191 3.4105
R4629 VGND.n195 VGND.n194 3.4105
R4630 VGND.n198 VGND.n197 3.4105
R4631 VGND.n201 VGND.n200 3.4105
R4632 VGND.n3001 VGND.n3000 3.4105
R4633 VGND.n3015 VGND.n96 3.4105
R4634 VGND.n3016 VGND.n95 3.4105
R4635 VGND.n3021 VGND.n90 3.4105
R4636 VGND.n3022 VGND.n89 3.4105
R4637 VGND.n3027 VGND.n84 3.4105
R4638 VGND.n3028 VGND.n83 3.4105
R4639 VGND.n3033 VGND.n78 3.4105
R4640 VGND.n3034 VGND.n77 3.4105
R4641 VGND.n3039 VGND.n72 3.4105
R4642 VGND.n3040 VGND.n71 3.4105
R4643 VGND.n3045 VGND.n66 3.4105
R4644 VGND.n3046 VGND.n65 3.4105
R4645 VGND.n3051 VGND.n60 3.4105
R4646 VGND.n3052 VGND.n59 3.4105
R4647 VGND.n3057 VGND.n52 3.4105
R4648 VGND.n528 VGND.n53 3.4105
R4649 VGND.n2828 VGND.n545 3.4105
R4650 VGND.n2841 VGND.n61 3.4105
R4651 VGND.n2477 VGND.n2476 3.4105
R4652 VGND.n2451 VGND.n2450 3.4105
R4653 VGND.n2757 VGND.n547 3.4105
R4654 VGND.n2492 VGND.n2491 3.4105
R4655 VGND.n2840 VGND.n64 3.4105
R4656 VGND.n2490 VGND.n2489 3.4105
R4657 VGND.n2479 VGND.n2478 3.4105
R4658 VGND.n2453 VGND.n2452 3.4105
R4659 VGND.n2640 VGND.n612 3.4105
R4660 VGND.n2505 VGND.n2504 3.4105
R4661 VGND.n2503 VGND.n2502 3.4105
R4662 VGND.n2839 VGND.n67 3.4105
R4663 VGND.n2430 VGND.n648 3.4105
R4664 VGND.n2431 VGND.n652 3.4105
R4665 VGND.n2432 VGND.n656 3.4105
R4666 VGND.n2434 VGND.n666 3.4105
R4667 VGND.n2408 VGND.n749 3.4105
R4668 VGND.n2429 VGND.n644 3.4105
R4669 VGND.n2516 VGND.n2515 3.4105
R4670 VGND.n2518 VGND.n2517 3.4105
R4671 VGND.n2838 VGND.n70 3.4105
R4672 VGND.n2300 VGND.n2299 3.4105
R4673 VGND.n2285 VGND.n2284 3.4105
R4674 VGND.n2274 VGND.n2273 3.4105
R4675 VGND.n2259 VGND.n2258 3.4105
R4676 VGND.n2233 VGND.n2232 3.4105
R4677 VGND.n2405 VGND.n750 3.4105
R4678 VGND.n2311 VGND.n2310 3.4105
R4679 VGND.n2428 VGND.n640 3.4105
R4680 VGND.n2531 VGND.n2530 3.4105
R4681 VGND.n2529 VGND.n2528 3.4105
R4682 VGND.n2837 VGND.n73 3.4105
R4683 VGND.n2313 VGND.n2312 3.4105
R4684 VGND.n2298 VGND.n2297 3.4105
R4685 VGND.n2287 VGND.n2286 3.4105
R4686 VGND.n2272 VGND.n2271 3.4105
R4687 VGND.n2261 VGND.n2260 3.4105
R4688 VGND.n2235 VGND.n2234 3.4105
R4689 VGND.n2665 VGND.n600 3.4105
R4690 VGND.n2324 VGND.n2323 3.4105
R4691 VGND.n2326 VGND.n2325 3.4105
R4692 VGND.n2427 VGND.n636 3.4105
R4693 VGND.n2542 VGND.n2541 3.4105
R4694 VGND.n2544 VGND.n2543 3.4105
R4695 VGND.n2836 VGND.n76 3.4105
R4696 VGND.n2145 VGND.n770 3.4105
R4697 VGND.n2146 VGND.n774 3.4105
R4698 VGND.n2147 VGND.n778 3.4105
R4699 VGND.n2148 VGND.n782 3.4105
R4700 VGND.n2149 VGND.n786 3.4105
R4701 VGND.n2150 VGND.n790 3.4105
R4702 VGND.n1937 VGND.n800 3.4105
R4703 VGND.n2126 VGND.n921 3.4105
R4704 VGND.n2144 VGND.n766 3.4105
R4705 VGND.n2339 VGND.n2338 3.4105
R4706 VGND.n2337 VGND.n2336 3.4105
R4707 VGND.n2426 VGND.n632 3.4105
R4708 VGND.n2557 VGND.n2556 3.4105
R4709 VGND.n2555 VGND.n2554 3.4105
R4710 VGND.n2835 VGND.n79 3.4105
R4711 VGND.n2055 VGND.n2054 3.4105
R4712 VGND.n2044 VGND.n2043 3.4105
R4713 VGND.n2029 VGND.n2028 3.4105
R4714 VGND.n2018 VGND.n2017 3.4105
R4715 VGND.n2003 VGND.n2002 3.4105
R4716 VGND.n1992 VGND.n1991 3.4105
R4717 VGND.n1977 VGND.n1976 3.4105
R4718 VGND.n1951 VGND.n1950 3.4105
R4719 VGND.n2123 VGND.n922 3.4105
R4720 VGND.n2070 VGND.n2069 3.4105
R4721 VGND.n2143 VGND.n762 3.4105
R4722 VGND.n2350 VGND.n2349 3.4105
R4723 VGND.n2352 VGND.n2351 3.4105
R4724 VGND.n2425 VGND.n628 3.4105
R4725 VGND.n2568 VGND.n2567 3.4105
R4726 VGND.n2570 VGND.n2569 3.4105
R4727 VGND.n2834 VGND.n82 3.4105
R4728 VGND.n2068 VGND.n2067 3.4105
R4729 VGND.n2057 VGND.n2056 3.4105
R4730 VGND.n2042 VGND.n2041 3.4105
R4731 VGND.n2031 VGND.n2030 3.4105
R4732 VGND.n2016 VGND.n2015 3.4105
R4733 VGND.n2005 VGND.n2004 3.4105
R4734 VGND.n1990 VGND.n1989 3.4105
R4735 VGND.n1979 VGND.n1978 3.4105
R4736 VGND.n1953 VGND.n1952 3.4105
R4737 VGND.n2690 VGND.n588 3.4105
R4738 VGND.n2083 VGND.n2082 3.4105
R4739 VGND.n2081 VGND.n2080 3.4105
R4740 VGND.n2142 VGND.n758 3.4105
R4741 VGND.n2365 VGND.n2364 3.4105
R4742 VGND.n2363 VGND.n2362 3.4105
R4743 VGND.n2424 VGND.n624 3.4105
R4744 VGND.n2583 VGND.n2582 3.4105
R4745 VGND.n2581 VGND.n2580 3.4105
R4746 VGND.n2833 VGND.n85 3.4105
R4747 VGND.n1915 VGND.n930 3.4105
R4748 VGND.n1916 VGND.n934 3.4105
R4749 VGND.n1917 VGND.n938 3.4105
R4750 VGND.n1918 VGND.n942 3.4105
R4751 VGND.n1919 VGND.n946 3.4105
R4752 VGND.n1920 VGND.n950 3.4105
R4753 VGND.n1921 VGND.n954 3.4105
R4754 VGND.n1922 VGND.n958 3.4105
R4755 VGND.n1923 VGND.n962 3.4105
R4756 VGND.n1925 VGND.n972 3.4105
R4757 VGND.n1899 VGND.n994 3.4105
R4758 VGND.n1914 VGND.n926 3.4105
R4759 VGND.n2099 VGND.n2098 3.4105
R4760 VGND.n2101 VGND.n2100 3.4105
R4761 VGND.n2141 VGND.n754 3.4105
R4762 VGND.n2381 VGND.n2380 3.4105
R4763 VGND.n2383 VGND.n2382 3.4105
R4764 VGND.n2423 VGND.n620 3.4105
R4765 VGND.n2599 VGND.n2598 3.4105
R4766 VGND.n2601 VGND.n2600 3.4105
R4767 VGND.n2832 VGND.n88 3.4105
R4768 VGND.n1874 VGND.n1873 3.4105
R4769 VGND.n1854 VGND.n1853 3.4105
R4770 VGND.n1843 VGND.n1842 3.4105
R4771 VGND.n1828 VGND.n1827 3.4105
R4772 VGND.n1817 VGND.n1816 3.4105
R4773 VGND.n1802 VGND.n1801 3.4105
R4774 VGND.n1791 VGND.n1790 3.4105
R4775 VGND.n1776 VGND.n1775 3.4105
R4776 VGND.n1765 VGND.n1764 3.4105
R4777 VGND.n1750 VGND.n1749 3.4105
R4778 VGND.n1724 VGND.n1723 3.4105
R4779 VGND.n1896 VGND.n995 3.4105
R4780 VGND.n2700 VGND.n2699 3.4105
R4781 VGND.n1913 VGND.n580 3.4105
R4782 VGND.n2677 VGND.n2676 3.4105
R4783 VGND.n2675 VGND.n2674 3.4105
R4784 VGND.n2140 VGND.n592 3.4105
R4785 VGND.n2652 VGND.n2651 3.4105
R4786 VGND.n2650 VGND.n2649 3.4105
R4787 VGND.n2422 VGND.n604 3.4105
R4788 VGND.n2627 VGND.n2626 3.4105
R4789 VGND.n2625 VGND.n2624 3.4105
R4790 VGND.n2831 VGND.n91 3.4105
R4791 VGND.n2702 VGND.n2701 3.4105
R4792 VGND.n1872 VGND.n1871 3.4105
R4793 VGND.n1856 VGND.n1855 3.4105
R4794 VGND.n1841 VGND.n1840 3.4105
R4795 VGND.n1830 VGND.n1829 3.4105
R4796 VGND.n1815 VGND.n1814 3.4105
R4797 VGND.n1804 VGND.n1803 3.4105
R4798 VGND.n1789 VGND.n1788 3.4105
R4799 VGND.n1778 VGND.n1777 3.4105
R4800 VGND.n1763 VGND.n1762 3.4105
R4801 VGND.n1752 VGND.n1751 3.4105
R4802 VGND.n1726 VGND.n1725 3.4105
R4803 VGND.n2715 VGND.n575 3.4105
R4804 VGND.n2703 VGND.n568 3.4105
R4805 VGND.n2698 VGND.n2697 3.4105
R4806 VGND.n2696 VGND.n2695 3.4105
R4807 VGND.n2678 VGND.n583 3.4105
R4808 VGND.n2673 VGND.n2672 3.4105
R4809 VGND.n2671 VGND.n2670 3.4105
R4810 VGND.n2653 VGND.n595 3.4105
R4811 VGND.n2648 VGND.n2647 3.4105
R4812 VGND.n2646 VGND.n2645 3.4105
R4813 VGND.n2628 VGND.n607 3.4105
R4814 VGND.n2623 VGND.n2622 3.4105
R4815 VGND.n2830 VGND.n94 3.4105
R4816 VGND.n2721 VGND.n2720 3.4105
R4817 VGND.n1301 VGND.n579 3.4105
R4818 VGND.n1302 VGND.n999 3.4105
R4819 VGND.n1303 VGND.n1003 3.4105
R4820 VGND.n1304 VGND.n1007 3.4105
R4821 VGND.n1305 VGND.n1011 3.4105
R4822 VGND.n1306 VGND.n1015 3.4105
R4823 VGND.n1307 VGND.n1019 3.4105
R4824 VGND.n1308 VGND.n1023 3.4105
R4825 VGND.n1309 VGND.n1027 3.4105
R4826 VGND.n1310 VGND.n1031 3.4105
R4827 VGND.n1311 VGND.n1035 3.4105
R4828 VGND.n1217 VGND.n1045 3.4105
R4829 VGND.n1287 VGND.n1286 3.4105
R4830 VGND.n2719 VGND.n2718 3.4105
R4831 VGND.n2717 VGND.n2716 3.4105
R4832 VGND.n997 VGND.n573 3.4105
R4833 VGND.n2694 VGND.n2693 3.4105
R4834 VGND.n2692 VGND.n2691 3.4105
R4835 VGND.n924 VGND.n586 3.4105
R4836 VGND.n2669 VGND.n2668 3.4105
R4837 VGND.n2667 VGND.n2666 3.4105
R4838 VGND.n752 VGND.n598 3.4105
R4839 VGND.n2644 VGND.n2643 3.4105
R4840 VGND.n2642 VGND.n2641 3.4105
R4841 VGND.n2621 VGND.n610 3.4105
R4842 VGND.n2829 VGND.n97 3.4105
R4843 VGND.n3014 VGND.n3013 3.4105
R4844 VGND.n3018 VGND.n3017 3.4105
R4845 VGND.n3020 VGND.n3019 3.4105
R4846 VGND.n3024 VGND.n3023 3.4105
R4847 VGND.n3026 VGND.n3025 3.4105
R4848 VGND.n3030 VGND.n3029 3.4105
R4849 VGND.n3032 VGND.n3031 3.4105
R4850 VGND.n3036 VGND.n3035 3.4105
R4851 VGND.n3038 VGND.n3037 3.4105
R4852 VGND.n3042 VGND.n3041 3.4105
R4853 VGND.n3044 VGND.n3043 3.4105
R4854 VGND.n3048 VGND.n3047 3.4105
R4855 VGND.n3050 VGND.n3049 3.4105
R4856 VGND.n3056 VGND.n3055 3.4105
R4857 VGND.n3012 VGND.n99 3.4105
R4858 VGND.n572 VGND.n571 3.4105
R4859 VGND.n2723 VGND.n2722 3.4105
R4860 VGND.n1521 VGND.n1520 3.4105
R4861 VGND.n1523 VGND.n1522 3.4105
R4862 VGND.n1529 VGND.n1528 3.4105
R4863 VGND.n1531 VGND.n1530 3.4105
R4864 VGND.n1537 VGND.n1536 3.4105
R4865 VGND.n1539 VGND.n1538 3.4105
R4866 VGND.n1545 VGND.n1544 3.4105
R4867 VGND.n1547 VGND.n1546 3.4105
R4868 VGND.n1553 VGND.n1552 3.4105
R4869 VGND.n1555 VGND.n1554 3.4105
R4870 VGND.n1204 VGND.n1067 3.4105
R4871 VGND.n1207 VGND.n1206 3.4105
R4872 VGND.n2735 VGND.n564 3.4105
R4873 VGND.n1205 VGND.n1124 3.4105
R4874 VGND.n1312 VGND.n1039 3.4105
R4875 VGND.n1737 VGND.n1736 3.4105
R4876 VGND.n1739 VGND.n1738 3.4105
R4877 VGND.n1924 VGND.n966 3.4105
R4878 VGND.n1964 VGND.n1963 3.4105
R4879 VGND.n1966 VGND.n1965 3.4105
R4880 VGND.n2151 VGND.n794 3.4105
R4881 VGND.n2246 VGND.n2245 3.4105
R4882 VGND.n2248 VGND.n2247 3.4105
R4883 VGND.n2433 VGND.n660 3.4105
R4884 VGND.n2464 VGND.n2463 3.4105
R4885 VGND.n2466 VGND.n2465 3.4105
R4886 VGND.n2842 VGND.n58 3.4105
R4887 VGND.n3054 VGND.n3053 3.4105
R4888 VGND.n1514 VGND.n1101 3.4105
R4889 VGND.n1500 VGND.n1499 3.4105
R4890 VGND.n1491 VGND.n1097 3.4105
R4891 VGND.n1481 VGND.n1094 3.4105
R4892 VGND.n1463 VGND.n1091 3.4105
R4893 VGND.n1468 VGND.n1088 3.4105
R4894 VGND.n1459 VGND.n1085 3.4105
R4895 VGND.n1449 VGND.n1082 3.4105
R4896 VGND.n1431 VGND.n1079 3.4105
R4897 VGND.n1436 VGND.n1076 3.4105
R4898 VGND.n1427 VGND.n1073 3.4105
R4899 VGND.n1417 VGND.n1070 3.4105
R4900 VGND.n1561 VGND.n1560 3.4105
R4901 VGND.n1402 VGND.n1401 3.4105
R4902 VGND.n1513 VGND.n1512 3.4105
R4903 VGND.n1496 VGND.n1495 3.4105
R4904 VGND.n1498 VGND.n1497 3.4105
R4905 VGND.n1493 VGND.n1492 3.4105
R4906 VGND.n1480 VGND.n1107 3.4105
R4907 VGND.n1465 VGND.n1464 3.4105
R4908 VGND.n1467 VGND.n1466 3.4105
R4909 VGND.n1461 VGND.n1460 3.4105
R4910 VGND.n1448 VGND.n1115 3.4105
R4911 VGND.n1433 VGND.n1432 3.4105
R4912 VGND.n1435 VGND.n1434 3.4105
R4913 VGND.n1429 VGND.n1428 3.4105
R4914 VGND.n1416 VGND.n1406 3.4105
R4915 VGND.n1405 VGND.n1066 3.4105
R4916 VGND.n1404 VGND.n1403 3.4105
R4917 VGND.n1571 VGND.n1570 3.4105
R4918 VGND.n1516 VGND.n1515 3.4105
R4919 VGND.n1517 VGND.n567 3.4105
R4920 VGND.n1519 VGND.n1518 3.4105
R4921 VGND.n1525 VGND.n1524 3.4105
R4922 VGND.n1527 VGND.n1526 3.4105
R4923 VGND.n1533 VGND.n1532 3.4105
R4924 VGND.n1535 VGND.n1534 3.4105
R4925 VGND.n1541 VGND.n1540 3.4105
R4926 VGND.n1543 VGND.n1542 3.4105
R4927 VGND.n1549 VGND.n1548 3.4105
R4928 VGND.n1551 VGND.n1550 3.4105
R4929 VGND.n1557 VGND.n1556 3.4105
R4930 VGND.n1559 VGND.n1558 3.4105
R4931 VGND.n1400 VGND.n1399 3.4105
R4932 VGND.n1324 VGND.n1054 3.4105
R4933 VGND.n2738 VGND.n561 3.4105
R4934 VGND.n2177 VGND.n2166 3.01226
R4935 VGND.n339 VGND.n338 3.01226
R4936 VGND.n2161 VGND.n847 2.63579
R4937 VGND.n8 VGND 2.52282
R4938 VGND.n11 VGND 2.52282
R4939 VGND.n14 VGND 2.52282
R4940 VGND.n17 VGND 2.52282
R4941 VGND.n20 VGND 2.52282
R4942 VGND.n23 VGND 2.52282
R4943 VGND.n26 VGND 2.52282
R4944 VGND.n29 VGND 2.52282
R4945 VGND.n32 VGND 2.52282
R4946 VGND.n35 VGND 2.52282
R4947 VGND.n38 VGND 2.52282
R4948 VGND.n41 VGND 2.52282
R4949 VGND.n44 VGND 2.52282
R4950 VGND.n47 VGND 2.52282
R4951 VGND.n50 VGND 2.52282
R4952 VGND.n2182 VGND.n2181 2.25932
R4953 VGND.n443 VGND.n442 2.25932
R4954 VGND.n412 VGND.n411 2.25932
R4955 VGND.n379 VGND.n378 2.25932
R4956 VGND.n347 VGND.n346 2.25932
R4957 VGND.n344 VGND.n343 2.25932
R4958 VGND.n479 VGND.n467 1.88285
R4959 VGND.n829 VGND.n817 1.88285
R4960 VGND.n509 VGND.n497 1.88285
R4961 VGND.n457 VGND.n456 1.8605
R4962 VGND.n2858 VGND.n3 1.8605
R4963 VGND.n51 VGND 1.79514
R4964 VGND.n1573 VGND.n562 1.76378
R4965 VGND.n51 VGND 1.57193
R4966 VGND.n3002 VGND.n3001 1.54254
R4967 VGND.n2828 VGND.n2759 1.54254
R4968 VGND.n2758 VGND.n2757 1.54254
R4969 VGND.n2640 VGND.n546 1.54254
R4970 VGND.n2408 VGND.n2407 1.54254
R4971 VGND.n2406 VGND.n2405 1.54254
R4972 VGND.n2665 VGND.n601 1.54254
R4973 VGND.n2126 VGND.n2125 1.54254
R4974 VGND.n2124 VGND.n2123 1.54254
R4975 VGND.n2690 VGND.n589 1.54254
R4976 VGND.n1899 VGND.n1898 1.54254
R4977 VGND.n1897 VGND.n1896 1.54254
R4978 VGND.n2715 VGND.n576 1.54254
R4979 VGND.n1287 VGND.n563 1.54254
R4980 VGND.n3012 VGND.n100 1.54254
R4981 VGND.n2736 VGND.n2735 1.54254
R4982 VGND.n1513 VGND.n562 1.54254
R4983 VGND.n2738 VGND.n2737 1.54254
R4984 VGND.n2189 VGND.n846 1.50638
R4985 VGND.n354 VGND.n353 1.50638
R4986 VGND.n3058 VGND 1.3946
R4987 VGND.n1572 VGND 1.3946
R4988 VGND VGND.n1053 1.3946
R4989 VGND.n3063 VGND.n3062 1.36426
R4990 VGND.n1209 VGND.n1208 1.13717
R4991 VGND.n1216 VGND.n1215 1.13717
R4992 VGND.n1214 VGND.n1213 1.13717
R4993 VGND.n1211 VGND.n1210 1.13717
R4994 VGND.n1926 VGND.n974 1.13717
R4995 VGND.n1930 VGND.n1929 1.13717
R4996 VGND.n1941 VGND.n1940 1.13717
R4997 VGND.n1939 VGND.n1938 1.13717
R4998 VGND.n1934 VGND.n1933 1.13717
R4999 VGND.n1932 VGND.n1931 1.13717
R5000 VGND.n2435 VGND.n668 1.13717
R5001 VGND.n2439 VGND.n2438 1.13717
R5002 VGND.n2441 VGND.n2440 1.13717
R5003 VGND.n527 VGND.n5 1.13717
R5004 VGND.n3060 VGND.n3059 1.13717
R5005 VGND.n1604 VGND.n1573 1.04899
R5006 VGND.n161 VGND.n59 1.00149
R5007 VGND.n164 VGND.n60 1.00149
R5008 VGND.n167 VGND.n65 1.00149
R5009 VGND.n170 VGND.n66 1.00149
R5010 VGND.n173 VGND.n71 1.00149
R5011 VGND.n176 VGND.n72 1.00149
R5012 VGND.n179 VGND.n77 1.00149
R5013 VGND.n182 VGND.n78 1.00149
R5014 VGND.n185 VGND.n83 1.00149
R5015 VGND.n188 VGND.n84 1.00149
R5016 VGND.n191 VGND.n89 1.00149
R5017 VGND.n194 VGND.n90 1.00149
R5018 VGND.n197 VGND.n95 1.00149
R5019 VGND.n200 VGND.n96 1.00149
R5020 VGND.n3000 VGND.n203 1.00149
R5021 VGND.n1403 VGND.n1402 1.00149
R5022 VGND.n1561 VGND.n1066 1.00149
R5023 VGND.n1417 VGND.n1416 1.00149
R5024 VGND.n1428 VGND.n1427 1.00149
R5025 VGND.n1436 VGND.n1435 1.00149
R5026 VGND.n1432 VGND.n1431 1.00149
R5027 VGND.n1449 VGND.n1448 1.00149
R5028 VGND.n1460 VGND.n1459 1.00149
R5029 VGND.n1468 VGND.n1467 1.00149
R5030 VGND.n1464 VGND.n1463 1.00149
R5031 VGND.n1481 VGND.n1480 1.00149
R5032 VGND.n1492 VGND.n1491 1.00149
R5033 VGND.n1500 VGND.n1498 1.00149
R5034 VGND.n1495 VGND.n1101 1.00149
R5035 VGND.n1512 VGND.n1103 1.00149
R5036 VGND.n1570 VGND.n1056 1.00149
R5037 VGND.n159 VGND.n52 0.973133
R5038 VGND.n3062 VGND.n3 0.964047
R5039 VGND.n435 VGND.n431 0.929432
R5040 VGND.n404 VGND.n400 0.929432
R5041 VGND.n371 VGND.n367 0.929432
R5042 VGND.n333 VGND.n331 0.929432
R5043 VGND.n383 VGND.n1 0.916608
R5044 VGND VGND.n8 0.839786
R5045 VGND VGND.n11 0.839786
R5046 VGND VGND.n14 0.839786
R5047 VGND VGND.n17 0.839786
R5048 VGND VGND.n20 0.839786
R5049 VGND VGND.n23 0.839786
R5050 VGND VGND.n26 0.839786
R5051 VGND VGND.n29 0.839786
R5052 VGND VGND.n32 0.839786
R5053 VGND VGND.n35 0.839786
R5054 VGND VGND.n38 0.839786
R5055 VGND VGND.n41 0.839786
R5056 VGND VGND.n44 0.839786
R5057 VGND VGND.n47 0.839786
R5058 VGND VGND.n50 0.839786
R5059 VGND.n461 VGND.n459 0.753441
R5060 VGND.n113 VGND.n111 0.753441
R5061 VGND.n309 VGND.n307 0.753441
R5062 VGND.n416 VGND.n393 0.753441
R5063 VGND.n2886 VGND.n2883 0.753441
R5064 VGND.n137 VGND.n134 0.753441
R5065 VGND.n3064 VGND.n3063 0.669548
R5066 VGND VGND.n0 0.542567
R5067 VGND.n3064 VGND.n1 0.507317
R5068 VGND.n3003 VGND.n3002 0.404308
R5069 VGND.n1614 VGND.n1613 0.376971
R5070 VGND.n1581 VGND.n1577 0.376971
R5071 VGND.n2189 VGND.n2188 0.376971
R5072 VGND.n2214 VGND.n2213 0.376971
R5073 VGND.n1706 VGND.n1705 0.376971
R5074 VGND.n347 VGND.n325 0.376971
R5075 VGND.n354 VGND.n326 0.376971
R5076 VGND VGND.n3064 0.37415
R5077 VGND.n564 VGND.n561 0.362676
R5078 VGND.n1286 VGND.n564 0.362676
R5079 VGND.n1286 VGND.n575 0.362676
R5080 VGND.n995 VGND.n575 0.362676
R5081 VGND.n995 VGND.n994 0.362676
R5082 VGND.n994 VGND.n588 0.362676
R5083 VGND.n922 VGND.n588 0.362676
R5084 VGND.n922 VGND.n921 0.362676
R5085 VGND.n921 VGND.n600 0.362676
R5086 VGND.n750 VGND.n600 0.362676
R5087 VGND.n750 VGND.n749 0.362676
R5088 VGND.n749 VGND.n612 0.362676
R5089 VGND.n612 VGND.n547 0.362676
R5090 VGND.n547 VGND.n545 0.362676
R5091 VGND.n545 VGND.n99 0.362676
R5092 VGND.n1206 VGND.n1054 0.362676
R5093 VGND.n1206 VGND.n1045 0.362676
R5094 VGND.n1725 VGND.n1045 0.362676
R5095 VGND.n1725 VGND.n1724 0.362676
R5096 VGND.n1724 VGND.n972 0.362676
R5097 VGND.n1952 VGND.n972 0.362676
R5098 VGND.n1952 VGND.n1951 0.362676
R5099 VGND.n1951 VGND.n800 0.362676
R5100 VGND.n2234 VGND.n800 0.362676
R5101 VGND.n2234 VGND.n2233 0.362676
R5102 VGND.n2233 VGND.n666 0.362676
R5103 VGND.n2452 VGND.n666 0.362676
R5104 VGND.n2452 VGND.n2451 0.362676
R5105 VGND.n2451 VGND.n53 0.362676
R5106 VGND.n3056 VGND.n53 0.362676
R5107 VGND.n1559 VGND.n1067 0.362676
R5108 VGND.n1067 VGND.n1035 0.362676
R5109 VGND.n1751 VGND.n1035 0.362676
R5110 VGND.n1751 VGND.n1750 0.362676
R5111 VGND.n1750 VGND.n962 0.362676
R5112 VGND.n1978 VGND.n962 0.362676
R5113 VGND.n1978 VGND.n1977 0.362676
R5114 VGND.n1977 VGND.n790 0.362676
R5115 VGND.n2260 VGND.n790 0.362676
R5116 VGND.n2260 VGND.n2259 0.362676
R5117 VGND.n2259 VGND.n656 0.362676
R5118 VGND.n2478 VGND.n656 0.362676
R5119 VGND.n2478 VGND.n2477 0.362676
R5120 VGND.n2477 VGND.n61 0.362676
R5121 VGND.n3050 VGND.n61 0.362676
R5122 VGND.n1556 VGND.n1555 0.362676
R5123 VGND.n1555 VGND.n1031 0.362676
R5124 VGND.n1763 VGND.n1031 0.362676
R5125 VGND.n1764 VGND.n1763 0.362676
R5126 VGND.n1764 VGND.n958 0.362676
R5127 VGND.n1990 VGND.n958 0.362676
R5128 VGND.n1991 VGND.n1990 0.362676
R5129 VGND.n1991 VGND.n786 0.362676
R5130 VGND.n2272 VGND.n786 0.362676
R5131 VGND.n2273 VGND.n2272 0.362676
R5132 VGND.n2273 VGND.n652 0.362676
R5133 VGND.n2490 VGND.n652 0.362676
R5134 VGND.n2491 VGND.n2490 0.362676
R5135 VGND.n2491 VGND.n64 0.362676
R5136 VGND.n3047 VGND.n64 0.362676
R5137 VGND.n1552 VGND.n1551 0.362676
R5138 VGND.n1552 VGND.n1027 0.362676
R5139 VGND.n1777 VGND.n1027 0.362676
R5140 VGND.n1777 VGND.n1776 0.362676
R5141 VGND.n1776 VGND.n954 0.362676
R5142 VGND.n2004 VGND.n954 0.362676
R5143 VGND.n2004 VGND.n2003 0.362676
R5144 VGND.n2003 VGND.n782 0.362676
R5145 VGND.n2286 VGND.n782 0.362676
R5146 VGND.n2286 VGND.n2285 0.362676
R5147 VGND.n2285 VGND.n648 0.362676
R5148 VGND.n2504 VGND.n648 0.362676
R5149 VGND.n2504 VGND.n2503 0.362676
R5150 VGND.n2503 VGND.n67 0.362676
R5151 VGND.n3044 VGND.n67 0.362676
R5152 VGND.n1548 VGND.n1547 0.362676
R5153 VGND.n1547 VGND.n1023 0.362676
R5154 VGND.n1789 VGND.n1023 0.362676
R5155 VGND.n1790 VGND.n1789 0.362676
R5156 VGND.n1790 VGND.n950 0.362676
R5157 VGND.n2016 VGND.n950 0.362676
R5158 VGND.n2017 VGND.n2016 0.362676
R5159 VGND.n2017 VGND.n778 0.362676
R5160 VGND.n2298 VGND.n778 0.362676
R5161 VGND.n2299 VGND.n2298 0.362676
R5162 VGND.n2299 VGND.n644 0.362676
R5163 VGND.n2516 VGND.n644 0.362676
R5164 VGND.n2517 VGND.n2516 0.362676
R5165 VGND.n2517 VGND.n70 0.362676
R5166 VGND.n3041 VGND.n70 0.362676
R5167 VGND.n1544 VGND.n1543 0.362676
R5168 VGND.n1544 VGND.n1019 0.362676
R5169 VGND.n1803 VGND.n1019 0.362676
R5170 VGND.n1803 VGND.n1802 0.362676
R5171 VGND.n1802 VGND.n946 0.362676
R5172 VGND.n2030 VGND.n946 0.362676
R5173 VGND.n2030 VGND.n2029 0.362676
R5174 VGND.n2029 VGND.n774 0.362676
R5175 VGND.n2312 VGND.n774 0.362676
R5176 VGND.n2312 VGND.n2311 0.362676
R5177 VGND.n2311 VGND.n640 0.362676
R5178 VGND.n2530 VGND.n640 0.362676
R5179 VGND.n2530 VGND.n2529 0.362676
R5180 VGND.n2529 VGND.n73 0.362676
R5181 VGND.n3038 VGND.n73 0.362676
R5182 VGND.n1540 VGND.n1539 0.362676
R5183 VGND.n1539 VGND.n1015 0.362676
R5184 VGND.n1815 VGND.n1015 0.362676
R5185 VGND.n1816 VGND.n1815 0.362676
R5186 VGND.n1816 VGND.n942 0.362676
R5187 VGND.n2042 VGND.n942 0.362676
R5188 VGND.n2043 VGND.n2042 0.362676
R5189 VGND.n2043 VGND.n770 0.362676
R5190 VGND.n2324 VGND.n770 0.362676
R5191 VGND.n2325 VGND.n2324 0.362676
R5192 VGND.n2325 VGND.n636 0.362676
R5193 VGND.n2542 VGND.n636 0.362676
R5194 VGND.n2543 VGND.n2542 0.362676
R5195 VGND.n2543 VGND.n76 0.362676
R5196 VGND.n3035 VGND.n76 0.362676
R5197 VGND.n1536 VGND.n1535 0.362676
R5198 VGND.n1536 VGND.n1011 0.362676
R5199 VGND.n1829 VGND.n1011 0.362676
R5200 VGND.n1829 VGND.n1828 0.362676
R5201 VGND.n1828 VGND.n938 0.362676
R5202 VGND.n2056 VGND.n938 0.362676
R5203 VGND.n2056 VGND.n2055 0.362676
R5204 VGND.n2055 VGND.n766 0.362676
R5205 VGND.n2338 VGND.n766 0.362676
R5206 VGND.n2338 VGND.n2337 0.362676
R5207 VGND.n2337 VGND.n632 0.362676
R5208 VGND.n2556 VGND.n632 0.362676
R5209 VGND.n2556 VGND.n2555 0.362676
R5210 VGND.n2555 VGND.n79 0.362676
R5211 VGND.n3032 VGND.n79 0.362676
R5212 VGND.n1532 VGND.n1531 0.362676
R5213 VGND.n1531 VGND.n1007 0.362676
R5214 VGND.n1841 VGND.n1007 0.362676
R5215 VGND.n1842 VGND.n1841 0.362676
R5216 VGND.n1842 VGND.n934 0.362676
R5217 VGND.n2068 VGND.n934 0.362676
R5218 VGND.n2069 VGND.n2068 0.362676
R5219 VGND.n2069 VGND.n762 0.362676
R5220 VGND.n2350 VGND.n762 0.362676
R5221 VGND.n2351 VGND.n2350 0.362676
R5222 VGND.n2351 VGND.n628 0.362676
R5223 VGND.n2568 VGND.n628 0.362676
R5224 VGND.n2569 VGND.n2568 0.362676
R5225 VGND.n2569 VGND.n82 0.362676
R5226 VGND.n3029 VGND.n82 0.362676
R5227 VGND.n1528 VGND.n1527 0.362676
R5228 VGND.n1528 VGND.n1003 0.362676
R5229 VGND.n1855 VGND.n1003 0.362676
R5230 VGND.n1855 VGND.n1854 0.362676
R5231 VGND.n1854 VGND.n930 0.362676
R5232 VGND.n2082 VGND.n930 0.362676
R5233 VGND.n2082 VGND.n2081 0.362676
R5234 VGND.n2081 VGND.n758 0.362676
R5235 VGND.n2364 VGND.n758 0.362676
R5236 VGND.n2364 VGND.n2363 0.362676
R5237 VGND.n2363 VGND.n624 0.362676
R5238 VGND.n2582 VGND.n624 0.362676
R5239 VGND.n2582 VGND.n2581 0.362676
R5240 VGND.n2581 VGND.n85 0.362676
R5241 VGND.n3026 VGND.n85 0.362676
R5242 VGND.n1524 VGND.n1523 0.362676
R5243 VGND.n1523 VGND.n999 0.362676
R5244 VGND.n1872 VGND.n999 0.362676
R5245 VGND.n1873 VGND.n1872 0.362676
R5246 VGND.n1873 VGND.n926 0.362676
R5247 VGND.n2099 VGND.n926 0.362676
R5248 VGND.n2100 VGND.n2099 0.362676
R5249 VGND.n2100 VGND.n754 0.362676
R5250 VGND.n2381 VGND.n754 0.362676
R5251 VGND.n2382 VGND.n2381 0.362676
R5252 VGND.n2382 VGND.n620 0.362676
R5253 VGND.n2599 VGND.n620 0.362676
R5254 VGND.n2600 VGND.n2599 0.362676
R5255 VGND.n2600 VGND.n88 0.362676
R5256 VGND.n3023 VGND.n88 0.362676
R5257 VGND.n1520 VGND.n1519 0.362676
R5258 VGND.n1520 VGND.n579 0.362676
R5259 VGND.n2701 VGND.n579 0.362676
R5260 VGND.n2701 VGND.n2700 0.362676
R5261 VGND.n2700 VGND.n580 0.362676
R5262 VGND.n2676 VGND.n580 0.362676
R5263 VGND.n2676 VGND.n2675 0.362676
R5264 VGND.n2675 VGND.n592 0.362676
R5265 VGND.n2651 VGND.n592 0.362676
R5266 VGND.n2651 VGND.n2650 0.362676
R5267 VGND.n2650 VGND.n604 0.362676
R5268 VGND.n2626 VGND.n604 0.362676
R5269 VGND.n2626 VGND.n2625 0.362676
R5270 VGND.n2625 VGND.n91 0.362676
R5271 VGND.n3020 VGND.n91 0.362676
R5272 VGND.n2722 VGND.n567 0.362676
R5273 VGND.n2722 VGND.n2721 0.362676
R5274 VGND.n2721 VGND.n568 0.362676
R5275 VGND.n2697 VGND.n568 0.362676
R5276 VGND.n2697 VGND.n2696 0.362676
R5277 VGND.n2696 VGND.n583 0.362676
R5278 VGND.n2672 VGND.n583 0.362676
R5279 VGND.n2672 VGND.n2671 0.362676
R5280 VGND.n2671 VGND.n595 0.362676
R5281 VGND.n2647 VGND.n595 0.362676
R5282 VGND.n2647 VGND.n2646 0.362676
R5283 VGND.n2646 VGND.n607 0.362676
R5284 VGND.n2622 VGND.n607 0.362676
R5285 VGND.n2622 VGND.n94 0.362676
R5286 VGND.n3017 VGND.n94 0.362676
R5287 VGND.n1515 VGND.n572 0.362676
R5288 VGND.n2718 VGND.n572 0.362676
R5289 VGND.n2718 VGND.n2717 0.362676
R5290 VGND.n2717 VGND.n573 0.362676
R5291 VGND.n2693 VGND.n573 0.362676
R5292 VGND.n2693 VGND.n2692 0.362676
R5293 VGND.n2692 VGND.n586 0.362676
R5294 VGND.n2668 VGND.n586 0.362676
R5295 VGND.n2668 VGND.n2667 0.362676
R5296 VGND.n2667 VGND.n598 0.362676
R5297 VGND.n2643 VGND.n598 0.362676
R5298 VGND.n2643 VGND.n2642 0.362676
R5299 VGND.n2642 VGND.n610 0.362676
R5300 VGND.n610 VGND.n97 0.362676
R5301 VGND.n3014 VGND.n97 0.362676
R5302 VGND.n1400 VGND.n1124 0.362676
R5303 VGND.n1124 VGND.n1039 0.362676
R5304 VGND.n1737 VGND.n1039 0.362676
R5305 VGND.n1738 VGND.n1737 0.362676
R5306 VGND.n1738 VGND.n966 0.362676
R5307 VGND.n1964 VGND.n966 0.362676
R5308 VGND.n1965 VGND.n1964 0.362676
R5309 VGND.n1965 VGND.n794 0.362676
R5310 VGND.n2246 VGND.n794 0.362676
R5311 VGND.n2247 VGND.n2246 0.362676
R5312 VGND.n2247 VGND.n660 0.362676
R5313 VGND.n2464 VGND.n660 0.362676
R5314 VGND.n2465 VGND.n2464 0.362676
R5315 VGND.n2465 VGND.n58 0.362676
R5316 VGND.n3053 VGND.n58 0.362676
R5317 VGND.n165 VGND.n162 0.349144
R5318 VGND.n168 VGND.n165 0.349144
R5319 VGND.n171 VGND.n168 0.349144
R5320 VGND.n174 VGND.n171 0.349144
R5321 VGND.n177 VGND.n174 0.349144
R5322 VGND.n180 VGND.n177 0.349144
R5323 VGND.n183 VGND.n180 0.349144
R5324 VGND.n186 VGND.n183 0.349144
R5325 VGND.n189 VGND.n186 0.349144
R5326 VGND.n192 VGND.n189 0.349144
R5327 VGND.n195 VGND.n192 0.349144
R5328 VGND.n198 VGND.n195 0.349144
R5329 VGND.n201 VGND.n198 0.349144
R5330 VGND.n1497 VGND.n1496 0.349144
R5331 VGND.n1497 VGND.n1493 0.349144
R5332 VGND.n1493 VGND.n1107 0.349144
R5333 VGND.n1465 VGND.n1107 0.349144
R5334 VGND.n1466 VGND.n1465 0.349144
R5335 VGND.n1466 VGND.n1461 0.349144
R5336 VGND.n1461 VGND.n1115 0.349144
R5337 VGND.n1433 VGND.n1115 0.349144
R5338 VGND.n1434 VGND.n1433 0.349144
R5339 VGND.n1434 VGND.n1429 0.349144
R5340 VGND.n1429 VGND.n1406 0.349144
R5341 VGND.n1406 VGND.n1405 0.349144
R5342 VGND.n1405 VGND.n1404 0.349144
R5343 VGND.n2731 VGND.n566 0.327628
R5344 VGND.n2728 VGND.n2724 0.327628
R5345 VGND.n1154 VGND.n1096 0.327628
R5346 VGND.n1159 VGND.n1095 0.327628
R5347 VGND.n1164 VGND.n1090 0.327628
R5348 VGND.n1169 VGND.n1089 0.327628
R5349 VGND.n1174 VGND.n1084 0.327628
R5350 VGND.n1179 VGND.n1083 0.327628
R5351 VGND.n1184 VGND.n1078 0.327628
R5352 VGND.n1189 VGND.n1077 0.327628
R5353 VGND.n1194 VGND.n1072 0.327628
R5354 VGND.n1199 VGND.n1071 0.327628
R5355 VGND.n1203 VGND.n1202 0.327628
R5356 VGND.n1149 VGND.n1137 0.327628
R5357 VGND.n1144 VGND.n1136 0.327628
R5358 VGND.n2996 VGND.n205 0.327628
R5359 VGND.n2993 VGND.n2989 0.327628
R5360 VGND.n2986 VGND.n207 0.327628
R5361 VGND.n2983 VGND.n2979 0.327628
R5362 VGND.n2976 VGND.n209 0.327628
R5363 VGND.n2973 VGND.n2969 0.327628
R5364 VGND.n2966 VGND.n211 0.327628
R5365 VGND.n2963 VGND.n2959 0.327628
R5366 VGND.n2956 VGND.n213 0.327628
R5367 VGND.n2953 VGND.n2949 0.327628
R5368 VGND.n2946 VGND.n215 0.327628
R5369 VGND.n2943 VGND.n2939 0.327628
R5370 VGND.n2936 VGND.n217 0.327628
R5371 VGND.n2933 VGND.n2929 0.327628
R5372 VGND.n2926 VGND.n221 0.327628
R5373 VGND.n2824 VGND.n544 0.327628
R5374 VGND.n2819 VGND.n543 0.327628
R5375 VGND.n2814 VGND.n542 0.327628
R5376 VGND.n2809 VGND.n541 0.327628
R5377 VGND.n2804 VGND.n540 0.327628
R5378 VGND.n2799 VGND.n539 0.327628
R5379 VGND.n2794 VGND.n538 0.327628
R5380 VGND.n2789 VGND.n537 0.327628
R5381 VGND.n2784 VGND.n536 0.327628
R5382 VGND.n2779 VGND.n535 0.327628
R5383 VGND.n2774 VGND.n534 0.327628
R5384 VGND.n2769 VGND.n533 0.327628
R5385 VGND.n2764 VGND.n532 0.327628
R5386 VGND.n2843 VGND.n526 0.327628
R5387 VGND.n2846 VGND.n524 0.327628
R5388 VGND.n2620 VGND.n2619 0.327628
R5389 VGND.n2616 VGND.n616 0.327628
R5390 VGND.n2611 VGND.n615 0.327628
R5391 VGND.n2606 VGND.n2602 0.327628
R5392 VGND.n2579 VGND.n2578 0.327628
R5393 VGND.n2575 VGND.n2571 0.327628
R5394 VGND.n2553 VGND.n2552 0.327628
R5395 VGND.n2549 VGND.n2545 0.327628
R5396 VGND.n2527 VGND.n2526 0.327628
R5397 VGND.n2523 VGND.n2519 0.327628
R5398 VGND.n2501 VGND.n2500 0.327628
R5399 VGND.n2497 VGND.n2493 0.327628
R5400 VGND.n2475 VGND.n2474 0.327628
R5401 VGND.n2471 VGND.n2467 0.327628
R5402 VGND.n2449 VGND.n2448 0.327628
R5403 VGND.n2636 VGND.n611 0.327628
R5404 VGND.n2633 VGND.n2629 0.327628
R5405 VGND.n2593 VGND.n614 0.327628
R5406 VGND.n2597 VGND.n2596 0.327628
R5407 VGND.n2588 VGND.n2584 0.327628
R5408 VGND.n2566 VGND.n2565 0.327628
R5409 VGND.n2562 VGND.n2558 0.327628
R5410 VGND.n2540 VGND.n2539 0.327628
R5411 VGND.n2536 VGND.n2532 0.327628
R5412 VGND.n2514 VGND.n2513 0.327628
R5413 VGND.n2510 VGND.n2506 0.327628
R5414 VGND.n2488 VGND.n2487 0.327628
R5415 VGND.n2484 VGND.n2480 0.327628
R5416 VGND.n2462 VGND.n2461 0.327628
R5417 VGND.n2458 VGND.n2454 0.327628
R5418 VGND.n2412 VGND.n609 0.327628
R5419 VGND.n2417 VGND.n608 0.327628
R5420 VGND.n2421 VGND.n2420 0.327628
R5421 VGND.n746 VGND.n683 0.327628
R5422 VGND.n741 VGND.n682 0.327628
R5423 VGND.n736 VGND.n681 0.327628
R5424 VGND.n731 VGND.n680 0.327628
R5425 VGND.n726 VGND.n679 0.327628
R5426 VGND.n721 VGND.n678 0.327628
R5427 VGND.n716 VGND.n677 0.327628
R5428 VGND.n711 VGND.n676 0.327628
R5429 VGND.n706 VGND.n675 0.327628
R5430 VGND.n701 VGND.n674 0.327628
R5431 VGND.n696 VGND.n673 0.327628
R5432 VGND.n691 VGND.n672 0.327628
R5433 VGND.n2401 VGND.n753 0.327628
R5434 VGND.n2398 VGND.n606 0.327628
R5435 VGND.n2393 VGND.n605 0.327628
R5436 VGND.n2388 VGND.n2384 0.327628
R5437 VGND.n2361 VGND.n2360 0.327628
R5438 VGND.n2357 VGND.n2353 0.327628
R5439 VGND.n2335 VGND.n2334 0.327628
R5440 VGND.n2331 VGND.n2327 0.327628
R5441 VGND.n2309 VGND.n2308 0.327628
R5442 VGND.n2305 VGND.n2301 0.327628
R5443 VGND.n2283 VGND.n2282 0.327628
R5444 VGND.n2279 VGND.n2275 0.327628
R5445 VGND.n2257 VGND.n2256 0.327628
R5446 VGND.n2253 VGND.n2249 0.327628
R5447 VGND.n2231 VGND.n2230 0.327628
R5448 VGND.n2661 VGND.n599 0.327628
R5449 VGND.n2658 VGND.n2654 0.327628
R5450 VGND.n2375 VGND.n603 0.327628
R5451 VGND.n2379 VGND.n2378 0.327628
R5452 VGND.n2370 VGND.n2366 0.327628
R5453 VGND.n2348 VGND.n2347 0.327628
R5454 VGND.n2344 VGND.n2340 0.327628
R5455 VGND.n2322 VGND.n2321 0.327628
R5456 VGND.n2318 VGND.n2314 0.327628
R5457 VGND.n2296 VGND.n2295 0.327628
R5458 VGND.n2292 VGND.n2288 0.327628
R5459 VGND.n2270 VGND.n2269 0.327628
R5460 VGND.n2266 VGND.n2262 0.327628
R5461 VGND.n2244 VGND.n2243 0.327628
R5462 VGND.n2240 VGND.n2236 0.327628
R5463 VGND.n2130 VGND.n597 0.327628
R5464 VGND.n2135 VGND.n596 0.327628
R5465 VGND.n2139 VGND.n2138 0.327628
R5466 VGND.n918 VGND.n865 0.327628
R5467 VGND.n913 VGND.n864 0.327628
R5468 VGND.n908 VGND.n863 0.327628
R5469 VGND.n903 VGND.n862 0.327628
R5470 VGND.n898 VGND.n861 0.327628
R5471 VGND.n893 VGND.n860 0.327628
R5472 VGND.n888 VGND.n859 0.327628
R5473 VGND.n883 VGND.n858 0.327628
R5474 VGND.n878 VGND.n857 0.327628
R5475 VGND.n873 VGND.n856 0.327628
R5476 VGND.n2152 VGND.n852 0.327628
R5477 VGND.n2155 VGND.n850 0.327628
R5478 VGND.n2119 VGND.n925 0.327628
R5479 VGND.n2116 VGND.n594 0.327628
R5480 VGND.n2111 VGND.n593 0.327628
R5481 VGND.n2106 VGND.n2102 0.327628
R5482 VGND.n2079 VGND.n2078 0.327628
R5483 VGND.n2075 VGND.n2071 0.327628
R5484 VGND.n2053 VGND.n2052 0.327628
R5485 VGND.n2049 VGND.n2045 0.327628
R5486 VGND.n2027 VGND.n2026 0.327628
R5487 VGND.n2023 VGND.n2019 0.327628
R5488 VGND.n2001 VGND.n2000 0.327628
R5489 VGND.n1997 VGND.n1993 0.327628
R5490 VGND.n1975 VGND.n1974 0.327628
R5491 VGND.n1971 VGND.n1967 0.327628
R5492 VGND.n1949 VGND.n1948 0.327628
R5493 VGND.n2686 VGND.n587 0.327628
R5494 VGND.n2683 VGND.n2679 0.327628
R5495 VGND.n2093 VGND.n591 0.327628
R5496 VGND.n2097 VGND.n2096 0.327628
R5497 VGND.n2088 VGND.n2084 0.327628
R5498 VGND.n2066 VGND.n2065 0.327628
R5499 VGND.n2062 VGND.n2058 0.327628
R5500 VGND.n2040 VGND.n2039 0.327628
R5501 VGND.n2036 VGND.n2032 0.327628
R5502 VGND.n2014 VGND.n2013 0.327628
R5503 VGND.n2010 VGND.n2006 0.327628
R5504 VGND.n1988 VGND.n1987 0.327628
R5505 VGND.n1984 VGND.n1980 0.327628
R5506 VGND.n1962 VGND.n1961 0.327628
R5507 VGND.n1958 VGND.n1954 0.327628
R5508 VGND.n1903 VGND.n585 0.327628
R5509 VGND.n1908 VGND.n584 0.327628
R5510 VGND.n1912 VGND.n1911 0.327628
R5511 VGND.n1630 VGND.n989 0.327628
R5512 VGND.n1635 VGND.n988 0.327628
R5513 VGND.n1640 VGND.n987 0.327628
R5514 VGND.n1645 VGND.n986 0.327628
R5515 VGND.n1650 VGND.n985 0.327628
R5516 VGND.n1655 VGND.n984 0.327628
R5517 VGND.n1660 VGND.n983 0.327628
R5518 VGND.n1665 VGND.n982 0.327628
R5519 VGND.n1670 VGND.n981 0.327628
R5520 VGND.n1675 VGND.n980 0.327628
R5521 VGND.n1680 VGND.n979 0.327628
R5522 VGND.n1685 VGND.n978 0.327628
R5523 VGND.n1892 VGND.n998 0.327628
R5524 VGND.n1889 VGND.n582 0.327628
R5525 VGND.n1884 VGND.n581 0.327628
R5526 VGND.n1879 VGND.n1875 0.327628
R5527 VGND.n1852 VGND.n1851 0.327628
R5528 VGND.n1848 VGND.n1844 0.327628
R5529 VGND.n1826 VGND.n1825 0.327628
R5530 VGND.n1822 VGND.n1818 0.327628
R5531 VGND.n1800 VGND.n1799 0.327628
R5532 VGND.n1796 VGND.n1792 0.327628
R5533 VGND.n1774 VGND.n1773 0.327628
R5534 VGND.n1770 VGND.n1766 0.327628
R5535 VGND.n1748 VGND.n1747 0.327628
R5536 VGND.n1744 VGND.n1740 0.327628
R5537 VGND.n1722 VGND.n1721 0.327628
R5538 VGND.n2711 VGND.n574 0.327628
R5539 VGND.n2708 VGND.n2704 0.327628
R5540 VGND.n1866 VGND.n578 0.327628
R5541 VGND.n1870 VGND.n1869 0.327628
R5542 VGND.n1861 VGND.n1857 0.327628
R5543 VGND.n1839 VGND.n1838 0.327628
R5544 VGND.n1835 VGND.n1831 0.327628
R5545 VGND.n1813 VGND.n1812 0.327628
R5546 VGND.n1809 VGND.n1805 0.327628
R5547 VGND.n1787 VGND.n1786 0.327628
R5548 VGND.n1783 VGND.n1779 0.327628
R5549 VGND.n1761 VGND.n1760 0.327628
R5550 VGND.n1757 VGND.n1753 0.327628
R5551 VGND.n1735 VGND.n1734 0.327628
R5552 VGND.n1731 VGND.n1727 0.327628
R5553 VGND.n1291 VGND.n570 0.327628
R5554 VGND.n1296 VGND.n569 0.327628
R5555 VGND.n1300 VGND.n1299 0.327628
R5556 VGND.n1283 VGND.n1230 0.327628
R5557 VGND.n1278 VGND.n1229 0.327628
R5558 VGND.n1273 VGND.n1228 0.327628
R5559 VGND.n1268 VGND.n1227 0.327628
R5560 VGND.n1263 VGND.n1226 0.327628
R5561 VGND.n1258 VGND.n1225 0.327628
R5562 VGND.n1253 VGND.n1224 0.327628
R5563 VGND.n1248 VGND.n1223 0.327628
R5564 VGND.n1243 VGND.n1222 0.327628
R5565 VGND.n1238 VGND.n1221 0.327628
R5566 VGND.n1313 VGND.n1132 0.327628
R5567 VGND.n1316 VGND.n1130 0.327628
R5568 VGND.n225 VGND.n98 0.327628
R5569 VGND.n230 VGND.n93 0.327628
R5570 VGND.n235 VGND.n92 0.327628
R5571 VGND.n240 VGND.n87 0.327628
R5572 VGND.n245 VGND.n86 0.327628
R5573 VGND.n250 VGND.n81 0.327628
R5574 VGND.n255 VGND.n80 0.327628
R5575 VGND.n260 VGND.n75 0.327628
R5576 VGND.n265 VGND.n74 0.327628
R5577 VGND.n270 VGND.n69 0.327628
R5578 VGND.n275 VGND.n68 0.327628
R5579 VGND.n280 VGND.n63 0.327628
R5580 VGND.n285 VGND.n62 0.327628
R5581 VGND.n290 VGND.n57 0.327628
R5582 VGND.n295 VGND.n56 0.327628
R5583 VGND.n1569 VGND.n1568 0.327628
R5584 VGND.n1565 VGND.n1062 0.327628
R5585 VGND.n1562 VGND.n1064 0.327628
R5586 VGND.n1422 VGND.n1418 0.327628
R5587 VGND.n1426 VGND.n1425 0.327628
R5588 VGND.n1441 VGND.n1437 0.327628
R5589 VGND.n1444 VGND.n1121 0.327628
R5590 VGND.n1454 VGND.n1450 0.327628
R5591 VGND.n1458 VGND.n1457 0.327628
R5592 VGND.n1473 VGND.n1469 0.327628
R5593 VGND.n1476 VGND.n1113 0.327628
R5594 VGND.n1486 VGND.n1482 0.327628
R5595 VGND.n1490 VGND.n1489 0.327628
R5596 VGND.n1505 VGND.n1501 0.327628
R5597 VGND.n1508 VGND.n1105 0.327628
R5598 VGND.n1334 VGND.n1100 0.327628
R5599 VGND.n1339 VGND.n1099 0.327628
R5600 VGND.n1344 VGND.n1098 0.327628
R5601 VGND.n1349 VGND.n1093 0.327628
R5602 VGND.n1354 VGND.n1092 0.327628
R5603 VGND.n1359 VGND.n1087 0.327628
R5604 VGND.n1364 VGND.n1086 0.327628
R5605 VGND.n1369 VGND.n1081 0.327628
R5606 VGND.n1374 VGND.n1080 0.327628
R5607 VGND.n1379 VGND.n1075 0.327628
R5608 VGND.n1384 VGND.n1074 0.327628
R5609 VGND.n1389 VGND.n1069 0.327628
R5610 VGND.n1394 VGND.n1068 0.327628
R5611 VGND.n1398 VGND.n1397 0.327628
R5612 VGND.n1329 VGND.n1325 0.327628
R5613 VGND.n1212 VGND.n1133 0.274941
R5614 VGND.n1212 VGND.n975 0.274941
R5615 VGND.n1927 VGND.n975 0.274941
R5616 VGND.n1928 VGND.n1927 0.274941
R5617 VGND.n1928 VGND.n973 0.274941
R5618 VGND.n1936 VGND.n973 0.274941
R5619 VGND.n1936 VGND.n1935 0.274941
R5620 VGND.n1935 VGND.n669 0.274941
R5621 VGND.n2436 VGND.n669 0.274941
R5622 VGND.n2437 VGND.n2436 0.274941
R5623 VGND.n2437 VGND.n667 0.274941
R5624 VGND.n667 VGND.n4 0.2218
R5625 VGND VGND.n527 0.218797
R5626 VGND VGND.n2441 0.218797
R5627 VGND.n2438 VGND 0.218797
R5628 VGND.n2435 VGND 0.218797
R5629 VGND.n1931 VGND 0.218797
R5630 VGND.n1934 VGND 0.218797
R5631 VGND.n1938 VGND 0.218797
R5632 VGND VGND.n1941 0.218797
R5633 VGND.n1929 VGND 0.218797
R5634 VGND.n1926 VGND 0.218797
R5635 VGND.n1210 VGND 0.218797
R5636 VGND.n1213 VGND 0.218797
R5637 VGND VGND.n1216 0.218797
R5638 VGND.n3060 VGND 0.218797
R5639 VGND.n1208 VGND 0.218797
R5640 VGND.n383 VGND.n323 0.213567
R5641 VGND.n2907 VGND.n323 0.213567
R5642 VGND.n2908 VGND.n2907 0.213567
R5643 VGND.n2908 VGND.n157 0.213567
R5644 VGND.n1604 VGND.n1603 0.213567
R5645 VGND.n1603 VGND.n845 0.213567
R5646 VGND.n2196 VGND.n845 0.213567
R5647 VGND.n2196 VGND.n2195 0.213567
R5648 VGND.n2195 VGND.n0 0.213567
R5649 VGND.n3003 VGND.n157 0.2073
R5650 VGND.n1573 VGND.n1572 0.175967
R5651 VGND.n3057 VGND 0.169807
R5652 VGND.n3052 VGND 0.169807
R5653 VGND.n3051 VGND 0.169807
R5654 VGND.n3046 VGND 0.169807
R5655 VGND.n3045 VGND 0.169807
R5656 VGND.n3040 VGND 0.169807
R5657 VGND.n3039 VGND 0.169807
R5658 VGND.n3034 VGND 0.169807
R5659 VGND.n3033 VGND 0.169807
R5660 VGND.n3028 VGND 0.169807
R5661 VGND.n3027 VGND 0.169807
R5662 VGND.n3022 VGND 0.169807
R5663 VGND.n3021 VGND 0.169807
R5664 VGND.n3016 VGND 0.169807
R5665 VGND.n3015 VGND 0.169807
R5666 VGND VGND.n528 0.169807
R5667 VGND.n2842 VGND 0.169807
R5668 VGND.n2841 VGND 0.169807
R5669 VGND.n2840 VGND 0.169807
R5670 VGND.n2839 VGND 0.169807
R5671 VGND.n2838 VGND 0.169807
R5672 VGND.n2837 VGND 0.169807
R5673 VGND.n2836 VGND 0.169807
R5674 VGND.n2835 VGND 0.169807
R5675 VGND.n2834 VGND 0.169807
R5676 VGND.n2833 VGND 0.169807
R5677 VGND.n2832 VGND 0.169807
R5678 VGND.n2831 VGND 0.169807
R5679 VGND.n2830 VGND 0.169807
R5680 VGND.n2829 VGND 0.169807
R5681 VGND.n2450 VGND 0.169807
R5682 VGND.n2466 VGND 0.169807
R5683 VGND.n2476 VGND 0.169807
R5684 VGND.n2492 VGND 0.169807
R5685 VGND.n2502 VGND 0.169807
R5686 VGND.n2518 VGND 0.169807
R5687 VGND.n2528 VGND 0.169807
R5688 VGND.n2544 VGND 0.169807
R5689 VGND.n2554 VGND 0.169807
R5690 VGND.n2570 VGND 0.169807
R5691 VGND.n2580 VGND 0.169807
R5692 VGND.n2601 VGND 0.169807
R5693 VGND.n2624 VGND 0.169807
R5694 VGND.n2623 VGND 0.169807
R5695 VGND.n2621 VGND 0.169807
R5696 VGND.n2453 VGND 0.169807
R5697 VGND.n2463 VGND 0.169807
R5698 VGND.n2479 VGND 0.169807
R5699 VGND.n2489 VGND 0.169807
R5700 VGND.n2505 VGND 0.169807
R5701 VGND.n2515 VGND 0.169807
R5702 VGND.n2531 VGND 0.169807
R5703 VGND.n2541 VGND 0.169807
R5704 VGND.n2557 VGND 0.169807
R5705 VGND.n2567 VGND 0.169807
R5706 VGND.n2583 VGND 0.169807
R5707 VGND.n2598 VGND 0.169807
R5708 VGND VGND.n2627 0.169807
R5709 VGND.n2628 VGND 0.169807
R5710 VGND.n2641 VGND 0.169807
R5711 VGND.n2434 VGND 0.169807
R5712 VGND.n2433 VGND 0.169807
R5713 VGND.n2432 VGND 0.169807
R5714 VGND.n2431 VGND 0.169807
R5715 VGND.n2430 VGND 0.169807
R5716 VGND.n2429 VGND 0.169807
R5717 VGND.n2428 VGND 0.169807
R5718 VGND.n2427 VGND 0.169807
R5719 VGND.n2426 VGND 0.169807
R5720 VGND.n2425 VGND 0.169807
R5721 VGND.n2424 VGND 0.169807
R5722 VGND.n2423 VGND 0.169807
R5723 VGND.n2422 VGND 0.169807
R5724 VGND.n2645 VGND 0.169807
R5725 VGND.n2644 VGND 0.169807
R5726 VGND.n2232 VGND 0.169807
R5727 VGND.n2248 VGND 0.169807
R5728 VGND.n2258 VGND 0.169807
R5729 VGND.n2274 VGND 0.169807
R5730 VGND.n2284 VGND 0.169807
R5731 VGND.n2300 VGND 0.169807
R5732 VGND.n2310 VGND 0.169807
R5733 VGND.n2326 VGND 0.169807
R5734 VGND.n2336 VGND 0.169807
R5735 VGND.n2352 VGND 0.169807
R5736 VGND.n2362 VGND 0.169807
R5737 VGND.n2383 VGND 0.169807
R5738 VGND.n2649 VGND 0.169807
R5739 VGND.n2648 VGND 0.169807
R5740 VGND.n752 VGND 0.169807
R5741 VGND.n2235 VGND 0.169807
R5742 VGND.n2245 VGND 0.169807
R5743 VGND.n2261 VGND 0.169807
R5744 VGND.n2271 VGND 0.169807
R5745 VGND.n2287 VGND 0.169807
R5746 VGND.n2297 VGND 0.169807
R5747 VGND.n2313 VGND 0.169807
R5748 VGND.n2323 VGND 0.169807
R5749 VGND.n2339 VGND 0.169807
R5750 VGND.n2349 VGND 0.169807
R5751 VGND.n2365 VGND 0.169807
R5752 VGND.n2380 VGND 0.169807
R5753 VGND VGND.n2652 0.169807
R5754 VGND.n2653 VGND 0.169807
R5755 VGND.n2666 VGND 0.169807
R5756 VGND.n1937 VGND 0.169807
R5757 VGND.n2151 VGND 0.169807
R5758 VGND.n2150 VGND 0.169807
R5759 VGND.n2149 VGND 0.169807
R5760 VGND.n2148 VGND 0.169807
R5761 VGND.n2147 VGND 0.169807
R5762 VGND.n2146 VGND 0.169807
R5763 VGND.n2145 VGND 0.169807
R5764 VGND.n2144 VGND 0.169807
R5765 VGND.n2143 VGND 0.169807
R5766 VGND.n2142 VGND 0.169807
R5767 VGND.n2141 VGND 0.169807
R5768 VGND.n2140 VGND 0.169807
R5769 VGND.n2670 VGND 0.169807
R5770 VGND.n2669 VGND 0.169807
R5771 VGND.n1950 VGND 0.169807
R5772 VGND.n1966 VGND 0.169807
R5773 VGND.n1976 VGND 0.169807
R5774 VGND.n1992 VGND 0.169807
R5775 VGND.n2002 VGND 0.169807
R5776 VGND.n2018 VGND 0.169807
R5777 VGND.n2028 VGND 0.169807
R5778 VGND.n2044 VGND 0.169807
R5779 VGND.n2054 VGND 0.169807
R5780 VGND.n2070 VGND 0.169807
R5781 VGND.n2080 VGND 0.169807
R5782 VGND.n2101 VGND 0.169807
R5783 VGND.n2674 VGND 0.169807
R5784 VGND.n2673 VGND 0.169807
R5785 VGND.n924 VGND 0.169807
R5786 VGND.n1953 VGND 0.169807
R5787 VGND.n1963 VGND 0.169807
R5788 VGND.n1979 VGND 0.169807
R5789 VGND.n1989 VGND 0.169807
R5790 VGND.n2005 VGND 0.169807
R5791 VGND.n2015 VGND 0.169807
R5792 VGND.n2031 VGND 0.169807
R5793 VGND.n2041 VGND 0.169807
R5794 VGND.n2057 VGND 0.169807
R5795 VGND.n2067 VGND 0.169807
R5796 VGND.n2083 VGND 0.169807
R5797 VGND.n2098 VGND 0.169807
R5798 VGND VGND.n2677 0.169807
R5799 VGND.n2678 VGND 0.169807
R5800 VGND.n2691 VGND 0.169807
R5801 VGND.n1925 VGND 0.169807
R5802 VGND.n1924 VGND 0.169807
R5803 VGND.n1923 VGND 0.169807
R5804 VGND.n1922 VGND 0.169807
R5805 VGND.n1921 VGND 0.169807
R5806 VGND.n1920 VGND 0.169807
R5807 VGND.n1919 VGND 0.169807
R5808 VGND.n1918 VGND 0.169807
R5809 VGND.n1917 VGND 0.169807
R5810 VGND.n1916 VGND 0.169807
R5811 VGND.n1915 VGND 0.169807
R5812 VGND.n1914 VGND 0.169807
R5813 VGND.n1913 VGND 0.169807
R5814 VGND.n2695 VGND 0.169807
R5815 VGND.n2694 VGND 0.169807
R5816 VGND.n1723 VGND 0.169807
R5817 VGND.n1739 VGND 0.169807
R5818 VGND.n1749 VGND 0.169807
R5819 VGND.n1765 VGND 0.169807
R5820 VGND.n1775 VGND 0.169807
R5821 VGND.n1791 VGND 0.169807
R5822 VGND.n1801 VGND 0.169807
R5823 VGND.n1817 VGND 0.169807
R5824 VGND.n1827 VGND 0.169807
R5825 VGND.n1843 VGND 0.169807
R5826 VGND.n1853 VGND 0.169807
R5827 VGND.n1874 VGND 0.169807
R5828 VGND.n2699 VGND 0.169807
R5829 VGND.n2698 VGND 0.169807
R5830 VGND.n997 VGND 0.169807
R5831 VGND.n1726 VGND 0.169807
R5832 VGND.n1736 VGND 0.169807
R5833 VGND.n1752 VGND 0.169807
R5834 VGND.n1762 VGND 0.169807
R5835 VGND.n1778 VGND 0.169807
R5836 VGND.n1788 VGND 0.169807
R5837 VGND.n1804 VGND 0.169807
R5838 VGND.n1814 VGND 0.169807
R5839 VGND.n1830 VGND 0.169807
R5840 VGND.n1840 VGND 0.169807
R5841 VGND.n1856 VGND 0.169807
R5842 VGND.n1871 VGND 0.169807
R5843 VGND VGND.n2702 0.169807
R5844 VGND.n2703 VGND 0.169807
R5845 VGND.n2716 VGND 0.169807
R5846 VGND VGND.n1217 0.169807
R5847 VGND.n1312 VGND 0.169807
R5848 VGND.n1311 VGND 0.169807
R5849 VGND.n1310 VGND 0.169807
R5850 VGND.n1309 VGND 0.169807
R5851 VGND.n1308 VGND 0.169807
R5852 VGND.n1307 VGND 0.169807
R5853 VGND.n1306 VGND 0.169807
R5854 VGND.n1305 VGND 0.169807
R5855 VGND.n1304 VGND 0.169807
R5856 VGND.n1303 VGND 0.169807
R5857 VGND.n1302 VGND 0.169807
R5858 VGND.n1301 VGND 0.169807
R5859 VGND.n2720 VGND 0.169807
R5860 VGND.n2719 VGND 0.169807
R5861 VGND.n3055 VGND 0.169807
R5862 VGND.n3054 VGND 0.169807
R5863 VGND.n3049 VGND 0.169807
R5864 VGND.n3048 VGND 0.169807
R5865 VGND.n3043 VGND 0.169807
R5866 VGND.n3042 VGND 0.169807
R5867 VGND.n3037 VGND 0.169807
R5868 VGND.n3036 VGND 0.169807
R5869 VGND.n3031 VGND 0.169807
R5870 VGND.n3030 VGND 0.169807
R5871 VGND.n3025 VGND 0.169807
R5872 VGND.n3024 VGND 0.169807
R5873 VGND.n3019 VGND 0.169807
R5874 VGND.n3018 VGND 0.169807
R5875 VGND.n3013 VGND 0.169807
R5876 VGND.n1207 VGND 0.169807
R5877 VGND.n1205 VGND 0.169807
R5878 VGND.n1204 VGND 0.169807
R5879 VGND.n1554 VGND 0.169807
R5880 VGND.n1553 VGND 0.169807
R5881 VGND.n1546 VGND 0.169807
R5882 VGND.n1545 VGND 0.169807
R5883 VGND.n1538 VGND 0.169807
R5884 VGND.n1537 VGND 0.169807
R5885 VGND.n1530 VGND 0.169807
R5886 VGND.n1529 VGND 0.169807
R5887 VGND.n1522 VGND 0.169807
R5888 VGND.n1521 VGND 0.169807
R5889 VGND.n2723 VGND 0.169807
R5890 VGND.n571 VGND 0.169807
R5891 VGND.n1571 VGND 0.169807
R5892 VGND.n1401 VGND 0.169807
R5893 VGND.n1560 VGND 0.169807
R5894 VGND VGND.n1070 0.169807
R5895 VGND VGND.n1073 0.169807
R5896 VGND VGND.n1076 0.169807
R5897 VGND VGND.n1079 0.169807
R5898 VGND VGND.n1082 0.169807
R5899 VGND VGND.n1085 0.169807
R5900 VGND VGND.n1088 0.169807
R5901 VGND VGND.n1091 0.169807
R5902 VGND VGND.n1094 0.169807
R5903 VGND VGND.n1097 0.169807
R5904 VGND.n1499 VGND 0.169807
R5905 VGND.n1514 VGND 0.169807
R5906 VGND.n1324 VGND 0.169807
R5907 VGND.n1399 VGND 0.169807
R5908 VGND.n1558 VGND 0.169807
R5909 VGND.n1557 VGND 0.169807
R5910 VGND.n1550 VGND 0.169807
R5911 VGND.n1549 VGND 0.169807
R5912 VGND.n1542 VGND 0.169807
R5913 VGND.n1541 VGND 0.169807
R5914 VGND.n1534 VGND 0.169807
R5915 VGND.n1533 VGND 0.169807
R5916 VGND.n1526 VGND 0.169807
R5917 VGND.n1525 VGND 0.169807
R5918 VGND.n1518 VGND 0.169807
R5919 VGND.n1517 VGND 0.169807
R5920 VGND.n1516 VGND 0.169807
R5921 VGND.n447 VGND 0.159538
R5922 VGND.n418 VGND 0.159538
R5923 VGND.n3061 VGND.n4 0.156949
R5924 VGND.n2737 VGND.n562 0.154425
R5925 VGND.n2737 VGND.n2736 0.154425
R5926 VGND.n2736 VGND.n563 0.154425
R5927 VGND.n576 VGND.n563 0.154425
R5928 VGND.n1897 VGND.n576 0.154425
R5929 VGND.n1898 VGND.n1897 0.154425
R5930 VGND.n1898 VGND.n589 0.154425
R5931 VGND.n2124 VGND.n589 0.154425
R5932 VGND.n2125 VGND.n2124 0.154425
R5933 VGND.n2125 VGND.n601 0.154425
R5934 VGND.n2406 VGND.n601 0.154425
R5935 VGND.n2407 VGND.n2406 0.154425
R5936 VGND.n2407 VGND.n546 0.154425
R5937 VGND.n2758 VGND.n546 0.154425
R5938 VGND.n2759 VGND.n2758 0.154425
R5939 VGND.n2759 VGND.n100 0.154425
R5940 VGND.n3002 VGND.n100 0.154425
R5941 VGND.n1572 VGND.n1053 0.154425
R5942 VGND.n1209 VGND.n1053 0.154425
R5943 VGND.n1215 VGND.n1209 0.154425
R5944 VGND.n1215 VGND.n1214 0.154425
R5945 VGND.n1214 VGND.n1211 0.154425
R5946 VGND.n1211 VGND.n974 0.154425
R5947 VGND.n1930 VGND.n974 0.154425
R5948 VGND.n1940 VGND.n1930 0.154425
R5949 VGND.n1940 VGND.n1939 0.154425
R5950 VGND.n1939 VGND.n1933 0.154425
R5951 VGND.n1933 VGND.n1932 0.154425
R5952 VGND.n1932 VGND.n668 0.154425
R5953 VGND.n2439 VGND.n668 0.154425
R5954 VGND.n2440 VGND.n2439 0.154425
R5955 VGND.n2440 VGND.n5 0.154425
R5956 VGND.n3059 VGND.n5 0.154425
R5957 VGND.n3059 VGND.n3058 0.154425
R5958 VGND.n1609 VGND.n1607 0.144904
R5959 VGND.n1586 VGND.n1578 0.144904
R5960 VGND.n2209 VGND.n2205 0.144904
R5961 VGND.n1701 VGND.n1697 0.144904
R5962 VGND.n52 VGND.n51 0.138284
R5963 VGND.n2732 VGND.n2731 0.13638
R5964 VGND.n2728 VGND.n2727 0.13638
R5965 VGND.n1154 VGND.n1153 0.13638
R5966 VGND.n1159 VGND.n1158 0.13638
R5967 VGND.n1164 VGND.n1163 0.13638
R5968 VGND.n1169 VGND.n1168 0.13638
R5969 VGND.n1174 VGND.n1173 0.13638
R5970 VGND.n1179 VGND.n1178 0.13638
R5971 VGND.n1184 VGND.n1183 0.13638
R5972 VGND.n1189 VGND.n1188 0.13638
R5973 VGND.n1194 VGND.n1193 0.13638
R5974 VGND.n1199 VGND.n1198 0.13638
R5975 VGND.n1202 VGND.n1140 0.13638
R5976 VGND.n1149 VGND.n1148 0.13638
R5977 VGND.n1144 VGND.n1143 0.13638
R5978 VGND.n2997 VGND.n2996 0.13638
R5979 VGND.n2993 VGND.n2992 0.13638
R5980 VGND.n2987 VGND.n2986 0.13638
R5981 VGND.n2983 VGND.n2982 0.13638
R5982 VGND.n2977 VGND.n2976 0.13638
R5983 VGND.n2973 VGND.n2972 0.13638
R5984 VGND.n2967 VGND.n2966 0.13638
R5985 VGND.n2963 VGND.n2962 0.13638
R5986 VGND.n2957 VGND.n2956 0.13638
R5987 VGND.n2953 VGND.n2952 0.13638
R5988 VGND.n2947 VGND.n2946 0.13638
R5989 VGND.n2943 VGND.n2942 0.13638
R5990 VGND.n2937 VGND.n2936 0.13638
R5991 VGND.n2933 VGND.n2932 0.13638
R5992 VGND.n2927 VGND.n2926 0.13638
R5993 VGND.n2824 VGND.n2823 0.13638
R5994 VGND.n2819 VGND.n2818 0.13638
R5995 VGND.n2814 VGND.n2813 0.13638
R5996 VGND.n2809 VGND.n2808 0.13638
R5997 VGND.n2804 VGND.n2803 0.13638
R5998 VGND.n2799 VGND.n2798 0.13638
R5999 VGND.n2794 VGND.n2793 0.13638
R6000 VGND.n2789 VGND.n2788 0.13638
R6001 VGND.n2784 VGND.n2783 0.13638
R6002 VGND.n2779 VGND.n2778 0.13638
R6003 VGND.n2774 VGND.n2773 0.13638
R6004 VGND.n2769 VGND.n2768 0.13638
R6005 VGND.n2764 VGND.n2763 0.13638
R6006 VGND.n530 VGND.n526 0.13638
R6007 VGND.n2846 VGND.n2845 0.13638
R6008 VGND.n2619 VGND.n619 0.13638
R6009 VGND.n2616 VGND.n2615 0.13638
R6010 VGND.n2611 VGND.n2610 0.13638
R6011 VGND.n2606 VGND.n2605 0.13638
R6012 VGND.n2578 VGND.n627 0.13638
R6013 VGND.n2575 VGND.n2574 0.13638
R6014 VGND.n2552 VGND.n635 0.13638
R6015 VGND.n2549 VGND.n2548 0.13638
R6016 VGND.n2526 VGND.n643 0.13638
R6017 VGND.n2523 VGND.n2522 0.13638
R6018 VGND.n2500 VGND.n651 0.13638
R6019 VGND.n2497 VGND.n2496 0.13638
R6020 VGND.n2474 VGND.n659 0.13638
R6021 VGND.n2471 VGND.n2470 0.13638
R6022 VGND.n2448 VGND.n2446 0.13638
R6023 VGND.n2637 VGND.n2636 0.13638
R6024 VGND.n2633 VGND.n2632 0.13638
R6025 VGND.n2593 VGND.n2592 0.13638
R6026 VGND.n2596 VGND.n623 0.13638
R6027 VGND.n2588 VGND.n2587 0.13638
R6028 VGND.n2565 VGND.n631 0.13638
R6029 VGND.n2562 VGND.n2561 0.13638
R6030 VGND.n2539 VGND.n639 0.13638
R6031 VGND.n2536 VGND.n2535 0.13638
R6032 VGND.n2513 VGND.n647 0.13638
R6033 VGND.n2510 VGND.n2509 0.13638
R6034 VGND.n2487 VGND.n655 0.13638
R6035 VGND.n2484 VGND.n2483 0.13638
R6036 VGND.n2461 VGND.n663 0.13638
R6037 VGND.n2458 VGND.n2457 0.13638
R6038 VGND.n2412 VGND.n2411 0.13638
R6039 VGND.n2417 VGND.n2416 0.13638
R6040 VGND.n2420 VGND.n686 0.13638
R6041 VGND.n746 VGND.n745 0.13638
R6042 VGND.n741 VGND.n740 0.13638
R6043 VGND.n736 VGND.n735 0.13638
R6044 VGND.n731 VGND.n730 0.13638
R6045 VGND.n726 VGND.n725 0.13638
R6046 VGND.n721 VGND.n720 0.13638
R6047 VGND.n716 VGND.n715 0.13638
R6048 VGND.n711 VGND.n710 0.13638
R6049 VGND.n706 VGND.n705 0.13638
R6050 VGND.n701 VGND.n700 0.13638
R6051 VGND.n696 VGND.n695 0.13638
R6052 VGND.n691 VGND.n690 0.13638
R6053 VGND.n2402 VGND.n2401 0.13638
R6054 VGND.n2398 VGND.n2397 0.13638
R6055 VGND.n2393 VGND.n2392 0.13638
R6056 VGND.n2388 VGND.n2387 0.13638
R6057 VGND.n2360 VGND.n761 0.13638
R6058 VGND.n2357 VGND.n2356 0.13638
R6059 VGND.n2334 VGND.n769 0.13638
R6060 VGND.n2331 VGND.n2330 0.13638
R6061 VGND.n2308 VGND.n777 0.13638
R6062 VGND.n2305 VGND.n2304 0.13638
R6063 VGND.n2282 VGND.n785 0.13638
R6064 VGND.n2279 VGND.n2278 0.13638
R6065 VGND.n2256 VGND.n793 0.13638
R6066 VGND.n2253 VGND.n2252 0.13638
R6067 VGND.n2230 VGND.n805 0.13638
R6068 VGND.n2662 VGND.n2661 0.13638
R6069 VGND.n2658 VGND.n2657 0.13638
R6070 VGND.n2375 VGND.n2374 0.13638
R6071 VGND.n2378 VGND.n757 0.13638
R6072 VGND.n2370 VGND.n2369 0.13638
R6073 VGND.n2347 VGND.n765 0.13638
R6074 VGND.n2344 VGND.n2343 0.13638
R6075 VGND.n2321 VGND.n773 0.13638
R6076 VGND.n2318 VGND.n2317 0.13638
R6077 VGND.n2295 VGND.n781 0.13638
R6078 VGND.n2292 VGND.n2291 0.13638
R6079 VGND.n2269 VGND.n789 0.13638
R6080 VGND.n2266 VGND.n2265 0.13638
R6081 VGND.n2243 VGND.n797 0.13638
R6082 VGND.n2240 VGND.n2239 0.13638
R6083 VGND.n2130 VGND.n2129 0.13638
R6084 VGND.n2135 VGND.n2134 0.13638
R6085 VGND.n2138 VGND.n868 0.13638
R6086 VGND.n918 VGND.n917 0.13638
R6087 VGND.n913 VGND.n912 0.13638
R6088 VGND.n908 VGND.n907 0.13638
R6089 VGND.n903 VGND.n902 0.13638
R6090 VGND.n898 VGND.n897 0.13638
R6091 VGND.n893 VGND.n892 0.13638
R6092 VGND.n888 VGND.n887 0.13638
R6093 VGND.n883 VGND.n882 0.13638
R6094 VGND.n878 VGND.n877 0.13638
R6095 VGND.n873 VGND.n872 0.13638
R6096 VGND.n854 VGND.n852 0.13638
R6097 VGND.n2155 VGND.n2154 0.13638
R6098 VGND.n2120 VGND.n2119 0.13638
R6099 VGND.n2116 VGND.n2115 0.13638
R6100 VGND.n2111 VGND.n2110 0.13638
R6101 VGND.n2106 VGND.n2105 0.13638
R6102 VGND.n2078 VGND.n933 0.13638
R6103 VGND.n2075 VGND.n2074 0.13638
R6104 VGND.n2052 VGND.n941 0.13638
R6105 VGND.n2049 VGND.n2048 0.13638
R6106 VGND.n2026 VGND.n949 0.13638
R6107 VGND.n2023 VGND.n2022 0.13638
R6108 VGND.n2000 VGND.n957 0.13638
R6109 VGND.n1997 VGND.n1996 0.13638
R6110 VGND.n1974 VGND.n965 0.13638
R6111 VGND.n1971 VGND.n1970 0.13638
R6112 VGND.n1948 VGND.n1946 0.13638
R6113 VGND.n2687 VGND.n2686 0.13638
R6114 VGND.n2683 VGND.n2682 0.13638
R6115 VGND.n2093 VGND.n2092 0.13638
R6116 VGND.n2096 VGND.n929 0.13638
R6117 VGND.n2088 VGND.n2087 0.13638
R6118 VGND.n2065 VGND.n937 0.13638
R6119 VGND.n2062 VGND.n2061 0.13638
R6120 VGND.n2039 VGND.n945 0.13638
R6121 VGND.n2036 VGND.n2035 0.13638
R6122 VGND.n2013 VGND.n953 0.13638
R6123 VGND.n2010 VGND.n2009 0.13638
R6124 VGND.n1987 VGND.n961 0.13638
R6125 VGND.n1984 VGND.n1983 0.13638
R6126 VGND.n1961 VGND.n969 0.13638
R6127 VGND.n1958 VGND.n1957 0.13638
R6128 VGND.n1903 VGND.n1902 0.13638
R6129 VGND.n1908 VGND.n1907 0.13638
R6130 VGND.n1911 VGND.n992 0.13638
R6131 VGND.n1630 VGND.n1629 0.13638
R6132 VGND.n1635 VGND.n1634 0.13638
R6133 VGND.n1640 VGND.n1639 0.13638
R6134 VGND.n1645 VGND.n1644 0.13638
R6135 VGND.n1650 VGND.n1649 0.13638
R6136 VGND.n1655 VGND.n1654 0.13638
R6137 VGND.n1660 VGND.n1659 0.13638
R6138 VGND.n1665 VGND.n1664 0.13638
R6139 VGND.n1670 VGND.n1669 0.13638
R6140 VGND.n1675 VGND.n1674 0.13638
R6141 VGND.n1680 VGND.n1679 0.13638
R6142 VGND.n1685 VGND.n1684 0.13638
R6143 VGND.n1893 VGND.n1892 0.13638
R6144 VGND.n1889 VGND.n1888 0.13638
R6145 VGND.n1884 VGND.n1883 0.13638
R6146 VGND.n1879 VGND.n1878 0.13638
R6147 VGND.n1851 VGND.n1006 0.13638
R6148 VGND.n1848 VGND.n1847 0.13638
R6149 VGND.n1825 VGND.n1014 0.13638
R6150 VGND.n1822 VGND.n1821 0.13638
R6151 VGND.n1799 VGND.n1022 0.13638
R6152 VGND.n1796 VGND.n1795 0.13638
R6153 VGND.n1773 VGND.n1030 0.13638
R6154 VGND.n1770 VGND.n1769 0.13638
R6155 VGND.n1747 VGND.n1038 0.13638
R6156 VGND.n1744 VGND.n1743 0.13638
R6157 VGND.n1721 VGND.n1050 0.13638
R6158 VGND.n2712 VGND.n2711 0.13638
R6159 VGND.n2708 VGND.n2707 0.13638
R6160 VGND.n1866 VGND.n1865 0.13638
R6161 VGND.n1869 VGND.n1002 0.13638
R6162 VGND.n1861 VGND.n1860 0.13638
R6163 VGND.n1838 VGND.n1010 0.13638
R6164 VGND.n1835 VGND.n1834 0.13638
R6165 VGND.n1812 VGND.n1018 0.13638
R6166 VGND.n1809 VGND.n1808 0.13638
R6167 VGND.n1786 VGND.n1026 0.13638
R6168 VGND.n1783 VGND.n1782 0.13638
R6169 VGND.n1760 VGND.n1034 0.13638
R6170 VGND.n1757 VGND.n1756 0.13638
R6171 VGND.n1734 VGND.n1042 0.13638
R6172 VGND.n1731 VGND.n1730 0.13638
R6173 VGND.n1291 VGND.n1290 0.13638
R6174 VGND.n1296 VGND.n1295 0.13638
R6175 VGND.n1299 VGND.n1233 0.13638
R6176 VGND.n1283 VGND.n1282 0.13638
R6177 VGND.n1278 VGND.n1277 0.13638
R6178 VGND.n1273 VGND.n1272 0.13638
R6179 VGND.n1268 VGND.n1267 0.13638
R6180 VGND.n1263 VGND.n1262 0.13638
R6181 VGND.n1258 VGND.n1257 0.13638
R6182 VGND.n1253 VGND.n1252 0.13638
R6183 VGND.n1248 VGND.n1247 0.13638
R6184 VGND.n1243 VGND.n1242 0.13638
R6185 VGND.n1238 VGND.n1237 0.13638
R6186 VGND.n1219 VGND.n1132 0.13638
R6187 VGND.n1316 VGND.n1315 0.13638
R6188 VGND.n225 VGND.n224 0.13638
R6189 VGND.n230 VGND.n229 0.13638
R6190 VGND.n235 VGND.n234 0.13638
R6191 VGND.n240 VGND.n239 0.13638
R6192 VGND.n245 VGND.n244 0.13638
R6193 VGND.n250 VGND.n249 0.13638
R6194 VGND.n255 VGND.n254 0.13638
R6195 VGND.n260 VGND.n259 0.13638
R6196 VGND.n265 VGND.n264 0.13638
R6197 VGND.n270 VGND.n269 0.13638
R6198 VGND.n275 VGND.n274 0.13638
R6199 VGND.n280 VGND.n279 0.13638
R6200 VGND.n285 VGND.n284 0.13638
R6201 VGND.n290 VGND.n289 0.13638
R6202 VGND.n295 VGND.n294 0.13638
R6203 VGND.n1568 VGND.n1059 0.13638
R6204 VGND.n1565 VGND.n1564 0.13638
R6205 VGND.n1413 VGND.n1064 0.13638
R6206 VGND.n1422 VGND.n1421 0.13638
R6207 VGND.n1425 VGND.n1410 0.13638
R6208 VGND.n1441 VGND.n1440 0.13638
R6209 VGND.n1445 VGND.n1444 0.13638
R6210 VGND.n1454 VGND.n1453 0.13638
R6211 VGND.n1457 VGND.n1119 0.13638
R6212 VGND.n1473 VGND.n1472 0.13638
R6213 VGND.n1477 VGND.n1476 0.13638
R6214 VGND.n1486 VGND.n1485 0.13638
R6215 VGND.n1489 VGND.n1111 0.13638
R6216 VGND.n1505 VGND.n1504 0.13638
R6217 VGND.n1509 VGND.n1508 0.13638
R6218 VGND.n1334 VGND.n1333 0.13638
R6219 VGND.n1339 VGND.n1338 0.13638
R6220 VGND.n1344 VGND.n1343 0.13638
R6221 VGND.n1349 VGND.n1348 0.13638
R6222 VGND.n1354 VGND.n1353 0.13638
R6223 VGND.n1359 VGND.n1358 0.13638
R6224 VGND.n1364 VGND.n1363 0.13638
R6225 VGND.n1369 VGND.n1368 0.13638
R6226 VGND.n1374 VGND.n1373 0.13638
R6227 VGND.n1379 VGND.n1378 0.13638
R6228 VGND.n1384 VGND.n1383 0.13638
R6229 VGND.n1389 VGND.n1388 0.13638
R6230 VGND.n1394 VGND.n1393 0.13638
R6231 VGND.n1397 VGND.n1127 0.13638
R6232 VGND.n1329 VGND.n1328 0.13638
R6233 VGND VGND.n447 0.120838
R6234 VGND.n1622 VGND.n1621 0.120292
R6235 VGND.n1621 VGND.n1605 0.120292
R6236 VGND.n1617 VGND.n1605 0.120292
R6237 VGND.n1617 VGND.n1616 0.120292
R6238 VGND.n1616 VGND.n1615 0.120292
R6239 VGND.n1615 VGND.n1607 0.120292
R6240 VGND.n1599 VGND.n1598 0.120292
R6241 VGND.n1594 VGND.n1593 0.120292
R6242 VGND.n1593 VGND.n1592 0.120292
R6243 VGND.n1592 VGND.n1576 0.120292
R6244 VGND.n1588 VGND.n1576 0.120292
R6245 VGND.n1588 VGND.n1587 0.120292
R6246 VGND.n1587 VGND.n1586 0.120292
R6247 VGND.n487 VGND.n464 0.120292
R6248 VGND.n481 VGND.n464 0.120292
R6249 VGND.n481 VGND.n480 0.120292
R6250 VGND.n480 VGND.n468 0.120292
R6251 VGND.n473 VGND.n468 0.120292
R6252 VGND.n473 VGND.n472 0.120292
R6253 VGND.n472 VGND.n471 0.120292
R6254 VGND.n812 VGND.n809 0.120292
R6255 VGND.n813 VGND.n812 0.120292
R6256 VGND.n837 VGND.n814 0.120292
R6257 VGND.n831 VGND.n814 0.120292
R6258 VGND.n831 VGND.n830 0.120292
R6259 VGND.n830 VGND.n818 0.120292
R6260 VGND.n823 VGND.n818 0.120292
R6261 VGND.n823 VGND.n822 0.120292
R6262 VGND.n822 VGND.n821 0.120292
R6263 VGND.n2191 VGND.n2190 0.120292
R6264 VGND.n2184 VGND.n2160 0.120292
R6265 VGND.n2179 VGND.n2160 0.120292
R6266 VGND.n2179 VGND.n2178 0.120292
R6267 VGND.n2175 VGND.n2174 0.120292
R6268 VGND.n2174 VGND.n2169 0.120292
R6269 VGND.n2170 VGND.n2169 0.120292
R6270 VGND.n2202 VGND.n2201 0.120292
R6271 VGND.n2222 VGND.n2221 0.120292
R6272 VGND.n2221 VGND.n2203 0.120292
R6273 VGND.n2217 VGND.n2203 0.120292
R6274 VGND.n2217 VGND.n2216 0.120292
R6275 VGND.n2216 VGND.n2215 0.120292
R6276 VGND.n2215 VGND.n2205 0.120292
R6277 VGND.n1694 VGND.n1693 0.120292
R6278 VGND.n1714 VGND.n1713 0.120292
R6279 VGND.n1713 VGND.n1695 0.120292
R6280 VGND.n1709 VGND.n1695 0.120292
R6281 VGND.n1709 VGND.n1708 0.120292
R6282 VGND.n1708 VGND.n1707 0.120292
R6283 VGND.n1707 VGND.n1697 0.120292
R6284 VGND.n517 VGND.n494 0.120292
R6285 VGND.n511 VGND.n494 0.120292
R6286 VGND.n511 VGND.n510 0.120292
R6287 VGND.n510 VGND.n498 0.120292
R6288 VGND.n503 VGND.n498 0.120292
R6289 VGND.n503 VGND.n502 0.120292
R6290 VGND.n502 VGND.n501 0.120292
R6291 VGND.n112 VGND.n108 0.120292
R6292 VGND.n117 VGND.n108 0.120292
R6293 VGND.n118 VGND.n117 0.120292
R6294 VGND.n119 VGND.n118 0.120292
R6295 VGND.n119 VGND.n106 0.120292
R6296 VGND.n123 VGND.n106 0.120292
R6297 VGND.n124 VGND.n123 0.120292
R6298 VGND.n439 VGND.n431 0.120292
R6299 VGND.n440 VGND.n439 0.120292
R6300 VGND.n440 VGND.n425 0.120292
R6301 VGND.n445 VGND.n425 0.120292
R6302 VGND.n446 VGND.n445 0.120292
R6303 VGND.n408 VGND.n400 0.120292
R6304 VGND.n409 VGND.n408 0.120292
R6305 VGND.n409 VGND.n394 0.120292
R6306 VGND.n414 VGND.n394 0.120292
R6307 VGND.n415 VGND.n414 0.120292
R6308 VGND.n375 VGND.n367 0.120292
R6309 VGND.n376 VGND.n375 0.120292
R6310 VGND.n376 VGND.n361 0.120292
R6311 VGND.n381 VGND.n361 0.120292
R6312 VGND.n382 VGND.n381 0.120292
R6313 VGND.n387 VGND.n384 0.120292
R6314 VGND.n340 VGND.n331 0.120292
R6315 VGND.n341 VGND.n340 0.120292
R6316 VGND.n342 VGND.n341 0.120292
R6317 VGND.n342 VGND.n327 0.120292
R6318 VGND.n348 VGND.n327 0.120292
R6319 VGND.n351 VGND.n350 0.120292
R6320 VGND.n2888 VGND.n2887 0.120292
R6321 VGND.n2888 VGND.n2880 0.120292
R6322 VGND.n2893 VGND.n2880 0.120292
R6323 VGND.n2894 VGND.n2893 0.120292
R6324 VGND.n2895 VGND.n2894 0.120292
R6325 VGND.n2895 VGND.n2878 0.120292
R6326 VGND.n2899 VGND.n2878 0.120292
R6327 VGND.n2901 VGND.n324 0.120292
R6328 VGND.n2906 VGND.n324 0.120292
R6329 VGND.n308 VGND.n302 0.120292
R6330 VGND.n313 VGND.n302 0.120292
R6331 VGND.n314 VGND.n313 0.120292
R6332 VGND.n315 VGND.n314 0.120292
R6333 VGND.n315 VGND.n300 0.120292
R6334 VGND.n319 VGND.n300 0.120292
R6335 VGND.n320 VGND.n319 0.120292
R6336 VGND.n2913 VGND.n2912 0.120292
R6337 VGND.n2912 VGND.n2911 0.120292
R6338 VGND.n139 VGND.n138 0.120292
R6339 VGND.n139 VGND.n131 0.120292
R6340 VGND.n144 VGND.n131 0.120292
R6341 VGND.n145 VGND.n144 0.120292
R6342 VGND.n146 VGND.n145 0.120292
R6343 VGND.n146 VGND.n129 0.120292
R6344 VGND.n150 VGND.n129 0.120292
R6345 VGND.n152 VGND.n125 0.120292
R6346 VGND.n156 VGND.n125 0.120292
R6347 VGND VGND.n418 0.119536
R6348 VGND.n1609 VGND 0.117202
R6349 VGND.n1578 VGND 0.117202
R6350 VGND.n2209 VGND 0.117202
R6351 VGND.n1701 VGND 0.117202
R6352 VGND.n2733 VGND.n2732 0.110872
R6353 VGND.n2727 VGND.n2726 0.110872
R6354 VGND.n1153 VGND.n1152 0.110872
R6355 VGND.n1158 VGND.n1157 0.110872
R6356 VGND.n1163 VGND.n1162 0.110872
R6357 VGND.n1168 VGND.n1167 0.110872
R6358 VGND.n1173 VGND.n1172 0.110872
R6359 VGND.n1178 VGND.n1177 0.110872
R6360 VGND.n1183 VGND.n1182 0.110872
R6361 VGND.n1188 VGND.n1187 0.110872
R6362 VGND.n1193 VGND.n1192 0.110872
R6363 VGND.n1198 VGND.n1197 0.110872
R6364 VGND.n1140 VGND.n1139 0.110872
R6365 VGND.n1148 VGND.n1147 0.110872
R6366 VGND.n1143 VGND.n1142 0.110872
R6367 VGND.n2823 VGND.n2822 0.110872
R6368 VGND.n2818 VGND.n2817 0.110872
R6369 VGND.n2813 VGND.n2812 0.110872
R6370 VGND.n2808 VGND.n2807 0.110872
R6371 VGND.n2803 VGND.n2802 0.110872
R6372 VGND.n2798 VGND.n2797 0.110872
R6373 VGND.n2793 VGND.n2792 0.110872
R6374 VGND.n2788 VGND.n2787 0.110872
R6375 VGND.n2783 VGND.n2782 0.110872
R6376 VGND.n2778 VGND.n2777 0.110872
R6377 VGND.n2773 VGND.n2772 0.110872
R6378 VGND.n2768 VGND.n2767 0.110872
R6379 VGND.n2763 VGND.n2762 0.110872
R6380 VGND.n531 VGND.n530 0.110872
R6381 VGND.n2845 VGND.n2844 0.110872
R6382 VGND.n619 VGND.n618 0.110872
R6383 VGND.n2615 VGND.n2614 0.110872
R6384 VGND.n2610 VGND.n2609 0.110872
R6385 VGND.n2605 VGND.n2604 0.110872
R6386 VGND.n627 VGND.n626 0.110872
R6387 VGND.n2574 VGND.n2573 0.110872
R6388 VGND.n635 VGND.n634 0.110872
R6389 VGND.n2548 VGND.n2547 0.110872
R6390 VGND.n643 VGND.n642 0.110872
R6391 VGND.n2522 VGND.n2521 0.110872
R6392 VGND.n651 VGND.n650 0.110872
R6393 VGND.n2496 VGND.n2495 0.110872
R6394 VGND.n659 VGND.n658 0.110872
R6395 VGND.n2470 VGND.n2469 0.110872
R6396 VGND.n2446 VGND.n2445 0.110872
R6397 VGND.n2638 VGND.n2637 0.110872
R6398 VGND.n2632 VGND.n2631 0.110872
R6399 VGND.n2592 VGND.n2591 0.110872
R6400 VGND.n623 VGND.n622 0.110872
R6401 VGND.n2587 VGND.n2586 0.110872
R6402 VGND.n631 VGND.n630 0.110872
R6403 VGND.n2561 VGND.n2560 0.110872
R6404 VGND.n639 VGND.n638 0.110872
R6405 VGND.n2535 VGND.n2534 0.110872
R6406 VGND.n647 VGND.n646 0.110872
R6407 VGND.n2509 VGND.n2508 0.110872
R6408 VGND.n655 VGND.n654 0.110872
R6409 VGND.n2483 VGND.n2482 0.110872
R6410 VGND.n663 VGND.n662 0.110872
R6411 VGND.n2457 VGND.n2456 0.110872
R6412 VGND.n2411 VGND.n2410 0.110872
R6413 VGND.n2416 VGND.n2415 0.110872
R6414 VGND.n686 VGND.n685 0.110872
R6415 VGND.n745 VGND.n744 0.110872
R6416 VGND.n740 VGND.n739 0.110872
R6417 VGND.n735 VGND.n734 0.110872
R6418 VGND.n730 VGND.n729 0.110872
R6419 VGND.n725 VGND.n724 0.110872
R6420 VGND.n720 VGND.n719 0.110872
R6421 VGND.n715 VGND.n714 0.110872
R6422 VGND.n710 VGND.n709 0.110872
R6423 VGND.n705 VGND.n704 0.110872
R6424 VGND.n700 VGND.n699 0.110872
R6425 VGND.n695 VGND.n694 0.110872
R6426 VGND.n690 VGND.n689 0.110872
R6427 VGND.n2403 VGND.n2402 0.110872
R6428 VGND.n2397 VGND.n2396 0.110872
R6429 VGND.n2392 VGND.n2391 0.110872
R6430 VGND.n2387 VGND.n2386 0.110872
R6431 VGND.n761 VGND.n760 0.110872
R6432 VGND.n2356 VGND.n2355 0.110872
R6433 VGND.n769 VGND.n768 0.110872
R6434 VGND.n2330 VGND.n2329 0.110872
R6435 VGND.n777 VGND.n776 0.110872
R6436 VGND.n2304 VGND.n2303 0.110872
R6437 VGND.n785 VGND.n784 0.110872
R6438 VGND.n2278 VGND.n2277 0.110872
R6439 VGND.n793 VGND.n792 0.110872
R6440 VGND.n2252 VGND.n2251 0.110872
R6441 VGND.n805 VGND.n804 0.110872
R6442 VGND.n2663 VGND.n2662 0.110872
R6443 VGND.n2657 VGND.n2656 0.110872
R6444 VGND.n2374 VGND.n2373 0.110872
R6445 VGND.n757 VGND.n756 0.110872
R6446 VGND.n2369 VGND.n2368 0.110872
R6447 VGND.n765 VGND.n764 0.110872
R6448 VGND.n2343 VGND.n2342 0.110872
R6449 VGND.n773 VGND.n772 0.110872
R6450 VGND.n2317 VGND.n2316 0.110872
R6451 VGND.n781 VGND.n780 0.110872
R6452 VGND.n2291 VGND.n2290 0.110872
R6453 VGND.n789 VGND.n788 0.110872
R6454 VGND.n2265 VGND.n2264 0.110872
R6455 VGND.n797 VGND.n796 0.110872
R6456 VGND.n2239 VGND.n2238 0.110872
R6457 VGND.n2129 VGND.n2128 0.110872
R6458 VGND.n2134 VGND.n2133 0.110872
R6459 VGND.n868 VGND.n867 0.110872
R6460 VGND.n917 VGND.n916 0.110872
R6461 VGND.n912 VGND.n911 0.110872
R6462 VGND.n907 VGND.n906 0.110872
R6463 VGND.n902 VGND.n901 0.110872
R6464 VGND.n897 VGND.n896 0.110872
R6465 VGND.n892 VGND.n891 0.110872
R6466 VGND.n887 VGND.n886 0.110872
R6467 VGND.n882 VGND.n881 0.110872
R6468 VGND.n877 VGND.n876 0.110872
R6469 VGND.n872 VGND.n871 0.110872
R6470 VGND.n855 VGND.n854 0.110872
R6471 VGND.n2154 VGND.n2153 0.110872
R6472 VGND.n2121 VGND.n2120 0.110872
R6473 VGND.n2115 VGND.n2114 0.110872
R6474 VGND.n2110 VGND.n2109 0.110872
R6475 VGND.n2105 VGND.n2104 0.110872
R6476 VGND.n933 VGND.n932 0.110872
R6477 VGND.n2074 VGND.n2073 0.110872
R6478 VGND.n941 VGND.n940 0.110872
R6479 VGND.n2048 VGND.n2047 0.110872
R6480 VGND.n949 VGND.n948 0.110872
R6481 VGND.n2022 VGND.n2021 0.110872
R6482 VGND.n957 VGND.n956 0.110872
R6483 VGND.n1996 VGND.n1995 0.110872
R6484 VGND.n965 VGND.n964 0.110872
R6485 VGND.n1970 VGND.n1969 0.110872
R6486 VGND.n1946 VGND.n1945 0.110872
R6487 VGND.n2688 VGND.n2687 0.110872
R6488 VGND.n2682 VGND.n2681 0.110872
R6489 VGND.n2092 VGND.n2091 0.110872
R6490 VGND.n929 VGND.n928 0.110872
R6491 VGND.n2087 VGND.n2086 0.110872
R6492 VGND.n937 VGND.n936 0.110872
R6493 VGND.n2061 VGND.n2060 0.110872
R6494 VGND.n945 VGND.n944 0.110872
R6495 VGND.n2035 VGND.n2034 0.110872
R6496 VGND.n953 VGND.n952 0.110872
R6497 VGND.n2009 VGND.n2008 0.110872
R6498 VGND.n961 VGND.n960 0.110872
R6499 VGND.n1983 VGND.n1982 0.110872
R6500 VGND.n969 VGND.n968 0.110872
R6501 VGND.n1957 VGND.n1956 0.110872
R6502 VGND.n1902 VGND.n1901 0.110872
R6503 VGND.n1907 VGND.n1906 0.110872
R6504 VGND.n992 VGND.n991 0.110872
R6505 VGND.n1629 VGND.n1628 0.110872
R6506 VGND.n1634 VGND.n1633 0.110872
R6507 VGND.n1639 VGND.n1638 0.110872
R6508 VGND.n1644 VGND.n1643 0.110872
R6509 VGND.n1649 VGND.n1648 0.110872
R6510 VGND.n1654 VGND.n1653 0.110872
R6511 VGND.n1659 VGND.n1658 0.110872
R6512 VGND.n1664 VGND.n1663 0.110872
R6513 VGND.n1669 VGND.n1668 0.110872
R6514 VGND.n1674 VGND.n1673 0.110872
R6515 VGND.n1679 VGND.n1678 0.110872
R6516 VGND.n1684 VGND.n1683 0.110872
R6517 VGND.n1894 VGND.n1893 0.110872
R6518 VGND.n1888 VGND.n1887 0.110872
R6519 VGND.n1883 VGND.n1882 0.110872
R6520 VGND.n1878 VGND.n1877 0.110872
R6521 VGND.n1006 VGND.n1005 0.110872
R6522 VGND.n1847 VGND.n1846 0.110872
R6523 VGND.n1014 VGND.n1013 0.110872
R6524 VGND.n1821 VGND.n1820 0.110872
R6525 VGND.n1022 VGND.n1021 0.110872
R6526 VGND.n1795 VGND.n1794 0.110872
R6527 VGND.n1030 VGND.n1029 0.110872
R6528 VGND.n1769 VGND.n1768 0.110872
R6529 VGND.n1038 VGND.n1037 0.110872
R6530 VGND.n1743 VGND.n1742 0.110872
R6531 VGND.n1050 VGND.n1049 0.110872
R6532 VGND.n2713 VGND.n2712 0.110872
R6533 VGND.n2707 VGND.n2706 0.110872
R6534 VGND.n1865 VGND.n1864 0.110872
R6535 VGND.n1002 VGND.n1001 0.110872
R6536 VGND.n1860 VGND.n1859 0.110872
R6537 VGND.n1010 VGND.n1009 0.110872
R6538 VGND.n1834 VGND.n1833 0.110872
R6539 VGND.n1018 VGND.n1017 0.110872
R6540 VGND.n1808 VGND.n1807 0.110872
R6541 VGND.n1026 VGND.n1025 0.110872
R6542 VGND.n1782 VGND.n1781 0.110872
R6543 VGND.n1034 VGND.n1033 0.110872
R6544 VGND.n1756 VGND.n1755 0.110872
R6545 VGND.n1042 VGND.n1041 0.110872
R6546 VGND.n1730 VGND.n1729 0.110872
R6547 VGND.n1290 VGND.n1289 0.110872
R6548 VGND.n1295 VGND.n1294 0.110872
R6549 VGND.n1233 VGND.n1232 0.110872
R6550 VGND.n1282 VGND.n1281 0.110872
R6551 VGND.n1277 VGND.n1276 0.110872
R6552 VGND.n1272 VGND.n1271 0.110872
R6553 VGND.n1267 VGND.n1266 0.110872
R6554 VGND.n1262 VGND.n1261 0.110872
R6555 VGND.n1257 VGND.n1256 0.110872
R6556 VGND.n1252 VGND.n1251 0.110872
R6557 VGND.n1247 VGND.n1246 0.110872
R6558 VGND.n1242 VGND.n1241 0.110872
R6559 VGND.n1237 VGND.n1236 0.110872
R6560 VGND.n1220 VGND.n1219 0.110872
R6561 VGND.n1315 VGND.n1314 0.110872
R6562 VGND.n224 VGND.n223 0.110872
R6563 VGND.n229 VGND.n228 0.110872
R6564 VGND.n234 VGND.n233 0.110872
R6565 VGND.n239 VGND.n238 0.110872
R6566 VGND.n244 VGND.n243 0.110872
R6567 VGND.n249 VGND.n248 0.110872
R6568 VGND.n254 VGND.n253 0.110872
R6569 VGND.n259 VGND.n258 0.110872
R6570 VGND.n264 VGND.n263 0.110872
R6571 VGND.n269 VGND.n268 0.110872
R6572 VGND.n274 VGND.n273 0.110872
R6573 VGND.n279 VGND.n278 0.110872
R6574 VGND.n284 VGND.n283 0.110872
R6575 VGND.n289 VGND.n288 0.110872
R6576 VGND.n294 VGND.n293 0.110872
R6577 VGND.n1061 VGND.n1059 0.110872
R6578 VGND.n1564 VGND.n1563 0.110872
R6579 VGND.n1414 VGND.n1413 0.110872
R6580 VGND.n1421 VGND.n1420 0.110872
R6581 VGND.n1410 VGND.n1409 0.110872
R6582 VGND.n1440 VGND.n1439 0.110872
R6583 VGND.n1446 VGND.n1445 0.110872
R6584 VGND.n1453 VGND.n1452 0.110872
R6585 VGND.n1119 VGND.n1118 0.110872
R6586 VGND.n1472 VGND.n1471 0.110872
R6587 VGND.n1478 VGND.n1477 0.110872
R6588 VGND.n1485 VGND.n1484 0.110872
R6589 VGND.n1111 VGND.n1110 0.110872
R6590 VGND.n1504 VGND.n1503 0.110872
R6591 VGND.n1510 VGND.n1509 0.110872
R6592 VGND.n1333 VGND.n1332 0.110872
R6593 VGND.n1338 VGND.n1337 0.110872
R6594 VGND.n1343 VGND.n1342 0.110872
R6595 VGND.n1348 VGND.n1347 0.110872
R6596 VGND.n1353 VGND.n1352 0.110872
R6597 VGND.n1358 VGND.n1357 0.110872
R6598 VGND.n1363 VGND.n1362 0.110872
R6599 VGND.n1368 VGND.n1367 0.110872
R6600 VGND.n1373 VGND.n1372 0.110872
R6601 VGND.n1378 VGND.n1377 0.110872
R6602 VGND.n1383 VGND.n1382 0.110872
R6603 VGND.n1388 VGND.n1387 0.110872
R6604 VGND.n1393 VGND.n1392 0.110872
R6605 VGND.n1127 VGND.n1126 0.110872
R6606 VGND.n1328 VGND.n1327 0.110872
R6607 VGND.n1599 VGND 0.0981562
R6608 VGND.n2191 VGND 0.0981562
R6609 VGND.n1693 VGND 0.0981562
R6610 VGND VGND.n487 0.0968542
R6611 VGND VGND.n837 0.0968542
R6612 VGND VGND.n2184 0.0968542
R6613 VGND.n2201 VGND 0.0968542
R6614 VGND VGND.n517 0.0968542
R6615 VGND.n112 VGND 0.0968542
R6616 VGND VGND.n387 0.0968542
R6617 VGND.n351 VGND 0.0968542
R6618 VGND.n2887 VGND 0.0968542
R6619 VGND.n308 VGND 0.0968542
R6620 VGND.n138 VGND 0.0968542
R6621 VGND.n3058 VGND 0.088625
R6622 VGND VGND.n3057 0.0790114
R6623 VGND.n3052 VGND 0.0790114
R6624 VGND VGND.n3051 0.0790114
R6625 VGND.n3046 VGND 0.0790114
R6626 VGND VGND.n3045 0.0790114
R6627 VGND.n3040 VGND 0.0790114
R6628 VGND VGND.n3039 0.0790114
R6629 VGND.n3034 VGND 0.0790114
R6630 VGND VGND.n3033 0.0790114
R6631 VGND.n3028 VGND 0.0790114
R6632 VGND VGND.n3027 0.0790114
R6633 VGND.n3022 VGND 0.0790114
R6634 VGND VGND.n3021 0.0790114
R6635 VGND.n3016 VGND 0.0790114
R6636 VGND VGND.n3015 0.0790114
R6637 VGND.n3001 VGND 0.0790114
R6638 VGND.n528 VGND 0.0790114
R6639 VGND.n2842 VGND 0.0790114
R6640 VGND VGND.n2841 0.0790114
R6641 VGND VGND.n2840 0.0790114
R6642 VGND VGND.n2839 0.0790114
R6643 VGND VGND.n2838 0.0790114
R6644 VGND VGND.n2837 0.0790114
R6645 VGND VGND.n2836 0.0790114
R6646 VGND VGND.n2835 0.0790114
R6647 VGND VGND.n2834 0.0790114
R6648 VGND VGND.n2833 0.0790114
R6649 VGND VGND.n2832 0.0790114
R6650 VGND VGND.n2831 0.0790114
R6651 VGND VGND.n2830 0.0790114
R6652 VGND VGND.n2829 0.0790114
R6653 VGND VGND.n2828 0.0790114
R6654 VGND.n2450 VGND 0.0790114
R6655 VGND.n2466 VGND 0.0790114
R6656 VGND.n2476 VGND 0.0790114
R6657 VGND.n2492 VGND 0.0790114
R6658 VGND.n2502 VGND 0.0790114
R6659 VGND.n2518 VGND 0.0790114
R6660 VGND.n2528 VGND 0.0790114
R6661 VGND.n2544 VGND 0.0790114
R6662 VGND.n2554 VGND 0.0790114
R6663 VGND.n2570 VGND 0.0790114
R6664 VGND.n2580 VGND 0.0790114
R6665 VGND.n2601 VGND 0.0790114
R6666 VGND.n2624 VGND 0.0790114
R6667 VGND VGND.n2623 0.0790114
R6668 VGND VGND.n2621 0.0790114
R6669 VGND.n2757 VGND 0.0790114
R6670 VGND.n2453 VGND 0.0790114
R6671 VGND.n2463 VGND 0.0790114
R6672 VGND.n2479 VGND 0.0790114
R6673 VGND.n2489 VGND 0.0790114
R6674 VGND.n2505 VGND 0.0790114
R6675 VGND.n2515 VGND 0.0790114
R6676 VGND.n2531 VGND 0.0790114
R6677 VGND.n2541 VGND 0.0790114
R6678 VGND.n2557 VGND 0.0790114
R6679 VGND.n2567 VGND 0.0790114
R6680 VGND.n2583 VGND 0.0790114
R6681 VGND.n2598 VGND 0.0790114
R6682 VGND.n2627 VGND 0.0790114
R6683 VGND.n2628 VGND 0.0790114
R6684 VGND.n2641 VGND 0.0790114
R6685 VGND VGND.n2640 0.0790114
R6686 VGND VGND.n2434 0.0790114
R6687 VGND VGND.n2433 0.0790114
R6688 VGND VGND.n2432 0.0790114
R6689 VGND VGND.n2431 0.0790114
R6690 VGND VGND.n2430 0.0790114
R6691 VGND VGND.n2429 0.0790114
R6692 VGND VGND.n2428 0.0790114
R6693 VGND VGND.n2427 0.0790114
R6694 VGND VGND.n2426 0.0790114
R6695 VGND VGND.n2425 0.0790114
R6696 VGND VGND.n2424 0.0790114
R6697 VGND VGND.n2423 0.0790114
R6698 VGND VGND.n2422 0.0790114
R6699 VGND.n2645 VGND 0.0790114
R6700 VGND VGND.n2644 0.0790114
R6701 VGND.n2408 VGND 0.0790114
R6702 VGND.n2232 VGND 0.0790114
R6703 VGND.n2248 VGND 0.0790114
R6704 VGND.n2258 VGND 0.0790114
R6705 VGND.n2274 VGND 0.0790114
R6706 VGND.n2284 VGND 0.0790114
R6707 VGND.n2300 VGND 0.0790114
R6708 VGND.n2310 VGND 0.0790114
R6709 VGND.n2326 VGND 0.0790114
R6710 VGND.n2336 VGND 0.0790114
R6711 VGND.n2352 VGND 0.0790114
R6712 VGND.n2362 VGND 0.0790114
R6713 VGND.n2383 VGND 0.0790114
R6714 VGND.n2649 VGND 0.0790114
R6715 VGND VGND.n2648 0.0790114
R6716 VGND.n752 VGND 0.0790114
R6717 VGND.n2405 VGND 0.0790114
R6718 VGND.n2235 VGND 0.0790114
R6719 VGND.n2245 VGND 0.0790114
R6720 VGND.n2261 VGND 0.0790114
R6721 VGND.n2271 VGND 0.0790114
R6722 VGND.n2287 VGND 0.0790114
R6723 VGND.n2297 VGND 0.0790114
R6724 VGND.n2313 VGND 0.0790114
R6725 VGND.n2323 VGND 0.0790114
R6726 VGND.n2339 VGND 0.0790114
R6727 VGND.n2349 VGND 0.0790114
R6728 VGND.n2365 VGND 0.0790114
R6729 VGND.n2380 VGND 0.0790114
R6730 VGND.n2652 VGND 0.0790114
R6731 VGND.n2653 VGND 0.0790114
R6732 VGND.n2666 VGND 0.0790114
R6733 VGND VGND.n2665 0.0790114
R6734 VGND VGND.n1937 0.0790114
R6735 VGND.n2151 VGND 0.0790114
R6736 VGND VGND.n2150 0.0790114
R6737 VGND VGND.n2149 0.0790114
R6738 VGND VGND.n2148 0.0790114
R6739 VGND VGND.n2147 0.0790114
R6740 VGND VGND.n2146 0.0790114
R6741 VGND VGND.n2145 0.0790114
R6742 VGND VGND.n2144 0.0790114
R6743 VGND VGND.n2143 0.0790114
R6744 VGND VGND.n2142 0.0790114
R6745 VGND VGND.n2141 0.0790114
R6746 VGND VGND.n2140 0.0790114
R6747 VGND.n2670 VGND 0.0790114
R6748 VGND VGND.n2669 0.0790114
R6749 VGND.n2126 VGND 0.0790114
R6750 VGND.n1950 VGND 0.0790114
R6751 VGND.n1966 VGND 0.0790114
R6752 VGND.n1976 VGND 0.0790114
R6753 VGND.n1992 VGND 0.0790114
R6754 VGND.n2002 VGND 0.0790114
R6755 VGND.n2018 VGND 0.0790114
R6756 VGND.n2028 VGND 0.0790114
R6757 VGND.n2044 VGND 0.0790114
R6758 VGND.n2054 VGND 0.0790114
R6759 VGND.n2070 VGND 0.0790114
R6760 VGND.n2080 VGND 0.0790114
R6761 VGND.n2101 VGND 0.0790114
R6762 VGND.n2674 VGND 0.0790114
R6763 VGND VGND.n2673 0.0790114
R6764 VGND.n924 VGND 0.0790114
R6765 VGND.n2123 VGND 0.0790114
R6766 VGND.n1953 VGND 0.0790114
R6767 VGND.n1963 VGND 0.0790114
R6768 VGND.n1979 VGND 0.0790114
R6769 VGND.n1989 VGND 0.0790114
R6770 VGND.n2005 VGND 0.0790114
R6771 VGND.n2015 VGND 0.0790114
R6772 VGND.n2031 VGND 0.0790114
R6773 VGND.n2041 VGND 0.0790114
R6774 VGND.n2057 VGND 0.0790114
R6775 VGND.n2067 VGND 0.0790114
R6776 VGND.n2083 VGND 0.0790114
R6777 VGND.n2098 VGND 0.0790114
R6778 VGND.n2677 VGND 0.0790114
R6779 VGND.n2678 VGND 0.0790114
R6780 VGND.n2691 VGND 0.0790114
R6781 VGND VGND.n2690 0.0790114
R6782 VGND VGND.n1925 0.0790114
R6783 VGND VGND.n1924 0.0790114
R6784 VGND VGND.n1923 0.0790114
R6785 VGND VGND.n1922 0.0790114
R6786 VGND VGND.n1921 0.0790114
R6787 VGND VGND.n1920 0.0790114
R6788 VGND VGND.n1919 0.0790114
R6789 VGND VGND.n1918 0.0790114
R6790 VGND VGND.n1917 0.0790114
R6791 VGND VGND.n1916 0.0790114
R6792 VGND VGND.n1915 0.0790114
R6793 VGND VGND.n1914 0.0790114
R6794 VGND VGND.n1913 0.0790114
R6795 VGND.n2695 VGND 0.0790114
R6796 VGND VGND.n2694 0.0790114
R6797 VGND.n1899 VGND 0.0790114
R6798 VGND.n1723 VGND 0.0790114
R6799 VGND.n1739 VGND 0.0790114
R6800 VGND.n1749 VGND 0.0790114
R6801 VGND.n1765 VGND 0.0790114
R6802 VGND.n1775 VGND 0.0790114
R6803 VGND.n1791 VGND 0.0790114
R6804 VGND.n1801 VGND 0.0790114
R6805 VGND.n1817 VGND 0.0790114
R6806 VGND.n1827 VGND 0.0790114
R6807 VGND.n1843 VGND 0.0790114
R6808 VGND.n1853 VGND 0.0790114
R6809 VGND.n1874 VGND 0.0790114
R6810 VGND.n2699 VGND 0.0790114
R6811 VGND VGND.n2698 0.0790114
R6812 VGND.n997 VGND 0.0790114
R6813 VGND.n1896 VGND 0.0790114
R6814 VGND.n1726 VGND 0.0790114
R6815 VGND.n1736 VGND 0.0790114
R6816 VGND.n1752 VGND 0.0790114
R6817 VGND.n1762 VGND 0.0790114
R6818 VGND.n1778 VGND 0.0790114
R6819 VGND.n1788 VGND 0.0790114
R6820 VGND.n1804 VGND 0.0790114
R6821 VGND.n1814 VGND 0.0790114
R6822 VGND.n1830 VGND 0.0790114
R6823 VGND.n1840 VGND 0.0790114
R6824 VGND.n1856 VGND 0.0790114
R6825 VGND.n1871 VGND 0.0790114
R6826 VGND.n2702 VGND 0.0790114
R6827 VGND.n2703 VGND 0.0790114
R6828 VGND.n2716 VGND 0.0790114
R6829 VGND VGND.n2715 0.0790114
R6830 VGND.n1217 VGND 0.0790114
R6831 VGND.n1312 VGND 0.0790114
R6832 VGND VGND.n1311 0.0790114
R6833 VGND VGND.n1310 0.0790114
R6834 VGND VGND.n1309 0.0790114
R6835 VGND VGND.n1308 0.0790114
R6836 VGND VGND.n1307 0.0790114
R6837 VGND VGND.n1306 0.0790114
R6838 VGND VGND.n1305 0.0790114
R6839 VGND VGND.n1304 0.0790114
R6840 VGND VGND.n1303 0.0790114
R6841 VGND VGND.n1302 0.0790114
R6842 VGND VGND.n1301 0.0790114
R6843 VGND.n2720 VGND 0.0790114
R6844 VGND VGND.n2719 0.0790114
R6845 VGND.n1287 VGND 0.0790114
R6846 VGND.n3055 VGND 0.0790114
R6847 VGND VGND.n3054 0.0790114
R6848 VGND.n3049 VGND 0.0790114
R6849 VGND VGND.n3048 0.0790114
R6850 VGND.n3043 VGND 0.0790114
R6851 VGND VGND.n3042 0.0790114
R6852 VGND.n3037 VGND 0.0790114
R6853 VGND VGND.n3036 0.0790114
R6854 VGND.n3031 VGND 0.0790114
R6855 VGND VGND.n3030 0.0790114
R6856 VGND.n3025 VGND 0.0790114
R6857 VGND VGND.n3024 0.0790114
R6858 VGND.n3019 VGND 0.0790114
R6859 VGND VGND.n3018 0.0790114
R6860 VGND.n3013 VGND 0.0790114
R6861 VGND VGND.n3012 0.0790114
R6862 VGND VGND.n1207 0.0790114
R6863 VGND VGND.n1205 0.0790114
R6864 VGND VGND.n1204 0.0790114
R6865 VGND.n1554 VGND 0.0790114
R6866 VGND VGND.n1553 0.0790114
R6867 VGND.n1546 VGND 0.0790114
R6868 VGND VGND.n1545 0.0790114
R6869 VGND.n1538 VGND 0.0790114
R6870 VGND VGND.n1537 0.0790114
R6871 VGND.n1530 VGND 0.0790114
R6872 VGND VGND.n1529 0.0790114
R6873 VGND.n1522 VGND 0.0790114
R6874 VGND VGND.n1521 0.0790114
R6875 VGND.n2723 VGND 0.0790114
R6876 VGND.n571 VGND 0.0790114
R6877 VGND.n2735 VGND 0.0790114
R6878 VGND VGND.n1571 0.0790114
R6879 VGND.n1401 VGND 0.0790114
R6880 VGND.n1560 VGND 0.0790114
R6881 VGND.n1070 VGND 0.0790114
R6882 VGND.n1073 VGND 0.0790114
R6883 VGND.n1076 VGND 0.0790114
R6884 VGND.n1079 VGND 0.0790114
R6885 VGND.n1082 VGND 0.0790114
R6886 VGND.n1085 VGND 0.0790114
R6887 VGND.n1088 VGND 0.0790114
R6888 VGND.n1091 VGND 0.0790114
R6889 VGND.n1094 VGND 0.0790114
R6890 VGND.n1097 VGND 0.0790114
R6891 VGND.n1499 VGND 0.0790114
R6892 VGND.n1514 VGND 0.0790114
R6893 VGND VGND.n1513 0.0790114
R6894 VGND.n1324 VGND 0.0790114
R6895 VGND.n1399 VGND 0.0790114
R6896 VGND.n1558 VGND 0.0790114
R6897 VGND VGND.n1557 0.0790114
R6898 VGND.n1550 VGND 0.0790114
R6899 VGND VGND.n1549 0.0790114
R6900 VGND.n1542 VGND 0.0790114
R6901 VGND VGND.n1541 0.0790114
R6902 VGND.n1534 VGND 0.0790114
R6903 VGND VGND.n1533 0.0790114
R6904 VGND.n1526 VGND 0.0790114
R6905 VGND VGND.n1525 0.0790114
R6906 VGND.n1518 VGND 0.0790114
R6907 VGND VGND.n1517 0.0790114
R6908 VGND VGND.n1516 0.0790114
R6909 VGND.n2738 VGND 0.0790114
R6910 VGND.n2998 VGND.n2997 0.0656596
R6911 VGND.n2992 VGND.n2991 0.0656596
R6912 VGND.n2988 VGND.n2987 0.0656596
R6913 VGND.n2982 VGND.n2981 0.0656596
R6914 VGND.n2978 VGND.n2977 0.0656596
R6915 VGND.n2972 VGND.n2971 0.0656596
R6916 VGND.n2968 VGND.n2967 0.0656596
R6917 VGND.n2962 VGND.n2961 0.0656596
R6918 VGND.n2958 VGND.n2957 0.0656596
R6919 VGND.n2952 VGND.n2951 0.0656596
R6920 VGND.n2948 VGND.n2947 0.0656596
R6921 VGND.n2942 VGND.n2941 0.0656596
R6922 VGND.n2938 VGND.n2937 0.0656596
R6923 VGND.n2932 VGND.n2931 0.0656596
R6924 VGND.n2928 VGND.n2927 0.0656596
R6925 VGND.n49 VGND 0.063
R6926 VGND.n46 VGND 0.063
R6927 VGND.n43 VGND 0.063
R6928 VGND.n40 VGND 0.063
R6929 VGND.n37 VGND 0.063
R6930 VGND.n34 VGND 0.063
R6931 VGND.n31 VGND 0.063
R6932 VGND.n28 VGND 0.063
R6933 VGND.n25 VGND 0.063
R6934 VGND.n22 VGND 0.063
R6935 VGND.n19 VGND 0.063
R6936 VGND.n16 VGND 0.063
R6937 VGND.n13 VGND 0.063
R6938 VGND.n10 VGND 0.063
R6939 VGND.n7 VGND 0.063
R6940 VGND VGND.n1622 0.0603958
R6941 VGND.n1598 VGND 0.0603958
R6942 VGND VGND.n1597 0.0603958
R6943 VGND.n1594 VGND 0.0603958
R6944 VGND.n489 VGND 0.0603958
R6945 VGND VGND.n488 0.0603958
R6946 VGND.n471 VGND 0.0603958
R6947 VGND.n839 VGND 0.0603958
R6948 VGND VGND.n838 0.0603958
R6949 VGND.n821 VGND 0.0603958
R6950 VGND.n2186 VGND 0.0603958
R6951 VGND VGND.n2185 0.0603958
R6952 VGND.n2178 VGND 0.0603958
R6953 VGND.n2175 VGND 0.0603958
R6954 VGND.n2170 VGND 0.0603958
R6955 VGND VGND.n2202 0.0603958
R6956 VGND.n2223 VGND 0.0603958
R6957 VGND VGND.n2222 0.0603958
R6958 VGND VGND.n1694 0.0603958
R6959 VGND.n1715 VGND 0.0603958
R6960 VGND VGND.n1714 0.0603958
R6961 VGND.n519 VGND 0.0603958
R6962 VGND VGND.n518 0.0603958
R6963 VGND.n501 VGND 0.0603958
R6964 VGND VGND.n124 0.0603958
R6965 VGND.n3004 VGND 0.0603958
R6966 VGND.n449 VGND 0.0603958
R6967 VGND VGND.n448 0.0603958
R6968 VGND.n420 VGND 0.0603958
R6969 VGND VGND.n419 0.0603958
R6970 VGND.n389 VGND 0.0603958
R6971 VGND VGND.n388 0.0603958
R6972 VGND.n384 VGND 0.0603958
R6973 VGND.n356 VGND 0.0603958
R6974 VGND VGND.n355 0.0603958
R6975 VGND VGND.n2899 0.0603958
R6976 VGND.n2900 VGND 0.0603958
R6977 VGND.n2901 VGND 0.0603958
R6978 VGND VGND.n320 0.0603958
R6979 VGND.n321 VGND 0.0603958
R6980 VGND.n2913 VGND 0.0603958
R6981 VGND VGND.n150 0.0603958
R6982 VGND.n151 VGND 0.0603958
R6983 VGND.n152 VGND 0.0603958
R6984 VGND.n2998 VGND 0.0574853
R6985 VGND.n2991 VGND 0.0574853
R6986 VGND.n2988 VGND 0.0574853
R6987 VGND.n2981 VGND 0.0574853
R6988 VGND.n2978 VGND 0.0574853
R6989 VGND.n2971 VGND 0.0574853
R6990 VGND.n2968 VGND 0.0574853
R6991 VGND.n2961 VGND 0.0574853
R6992 VGND.n2958 VGND 0.0574853
R6993 VGND.n2951 VGND 0.0574853
R6994 VGND.n2948 VGND 0.0574853
R6995 VGND.n2941 VGND 0.0574853
R6996 VGND.n2938 VGND 0.0574853
R6997 VGND.n2931 VGND 0.0574853
R6998 VGND.n2928 VGND 0.0574853
R6999 VGND.n1055 VGND 0.0489375
R7000 VGND.n1102 VGND 0.0489375
R7001 VGND.n202 VGND 0.0489375
R7002 VGND.n158 VGND 0.0489375
R7003 VGND.n160 VGND 0.0489375
R7004 VGND.n163 VGND 0.0489375
R7005 VGND.n166 VGND 0.0489375
R7006 VGND.n169 VGND 0.0489375
R7007 VGND.n172 VGND 0.0489375
R7008 VGND.n175 VGND 0.0489375
R7009 VGND.n178 VGND 0.0489375
R7010 VGND.n181 VGND 0.0489375
R7011 VGND.n184 VGND 0.0489375
R7012 VGND.n187 VGND 0.0489375
R7013 VGND.n190 VGND 0.0489375
R7014 VGND.n193 VGND 0.0489375
R7015 VGND.n196 VGND 0.0489375
R7016 VGND.n199 VGND 0.0489375
R7017 VGND.n1123 VGND 0.0489375
R7018 VGND.n1065 VGND 0.0489375
R7019 VGND.n1415 VGND 0.0489375
R7020 VGND.n1407 VGND 0.0489375
R7021 VGND.n1122 VGND 0.0489375
R7022 VGND.n1430 VGND 0.0489375
R7023 VGND.n1447 VGND 0.0489375
R7024 VGND.n1116 VGND 0.0489375
R7025 VGND.n1114 VGND 0.0489375
R7026 VGND.n1462 VGND 0.0489375
R7027 VGND.n1479 VGND 0.0489375
R7028 VGND.n1108 VGND 0.0489375
R7029 VGND.n1106 VGND 0.0489375
R7030 VGND.n1494 VGND 0.0489375
R7031 VGND.n2 VGND 0.0445
R7032 VGND.n3 VGND.n2 0.043
R7033 VGND VGND.n2733 0.037734
R7034 VGND.n2726 VGND 0.037734
R7035 VGND.n1152 VGND 0.037734
R7036 VGND.n1157 VGND 0.037734
R7037 VGND.n1162 VGND 0.037734
R7038 VGND.n1167 VGND 0.037734
R7039 VGND.n1172 VGND 0.037734
R7040 VGND.n1177 VGND 0.037734
R7041 VGND.n1182 VGND 0.037734
R7042 VGND.n1187 VGND 0.037734
R7043 VGND.n1192 VGND 0.037734
R7044 VGND.n1197 VGND 0.037734
R7045 VGND.n1139 VGND 0.037734
R7046 VGND.n1147 VGND 0.037734
R7047 VGND.n1142 VGND 0.037734
R7048 VGND VGND.n1135 0.037734
R7049 VGND VGND.n220 0.037734
R7050 VGND.n2822 VGND 0.037734
R7051 VGND.n2817 VGND 0.037734
R7052 VGND.n2812 VGND 0.037734
R7053 VGND.n2807 VGND 0.037734
R7054 VGND.n2802 VGND 0.037734
R7055 VGND.n2797 VGND 0.037734
R7056 VGND.n2792 VGND 0.037734
R7057 VGND.n2787 VGND 0.037734
R7058 VGND.n2782 VGND 0.037734
R7059 VGND.n2777 VGND 0.037734
R7060 VGND.n2772 VGND 0.037734
R7061 VGND.n2767 VGND 0.037734
R7062 VGND.n2762 VGND 0.037734
R7063 VGND VGND.n531 0.037734
R7064 VGND.n2844 VGND 0.037734
R7065 VGND VGND.n523 0.037734
R7066 VGND.n618 VGND 0.037734
R7067 VGND.n2614 VGND 0.037734
R7068 VGND.n2609 VGND 0.037734
R7069 VGND.n2604 VGND 0.037734
R7070 VGND.n626 VGND 0.037734
R7071 VGND.n2573 VGND 0.037734
R7072 VGND.n634 VGND 0.037734
R7073 VGND.n2547 VGND 0.037734
R7074 VGND.n642 VGND 0.037734
R7075 VGND.n2521 VGND 0.037734
R7076 VGND.n650 VGND 0.037734
R7077 VGND.n2495 VGND 0.037734
R7078 VGND.n658 VGND 0.037734
R7079 VGND.n2469 VGND 0.037734
R7080 VGND.n2445 VGND 0.037734
R7081 VGND VGND.n2443 0.037734
R7082 VGND VGND.n2638 0.037734
R7083 VGND.n2631 VGND 0.037734
R7084 VGND.n2591 VGND 0.037734
R7085 VGND.n622 VGND 0.037734
R7086 VGND.n2586 VGND 0.037734
R7087 VGND.n630 VGND 0.037734
R7088 VGND.n2560 VGND 0.037734
R7089 VGND.n638 VGND 0.037734
R7090 VGND.n2534 VGND 0.037734
R7091 VGND.n646 VGND 0.037734
R7092 VGND.n2508 VGND 0.037734
R7093 VGND.n654 VGND 0.037734
R7094 VGND.n2482 VGND 0.037734
R7095 VGND.n662 VGND 0.037734
R7096 VGND.n2456 VGND 0.037734
R7097 VGND VGND.n665 0.037734
R7098 VGND.n2410 VGND 0.037734
R7099 VGND.n2415 VGND 0.037734
R7100 VGND.n685 VGND 0.037734
R7101 VGND.n744 VGND 0.037734
R7102 VGND.n739 VGND 0.037734
R7103 VGND.n734 VGND 0.037734
R7104 VGND.n729 VGND 0.037734
R7105 VGND.n724 VGND 0.037734
R7106 VGND.n719 VGND 0.037734
R7107 VGND.n714 VGND 0.037734
R7108 VGND.n709 VGND 0.037734
R7109 VGND.n704 VGND 0.037734
R7110 VGND.n699 VGND 0.037734
R7111 VGND.n694 VGND 0.037734
R7112 VGND.n689 VGND 0.037734
R7113 VGND VGND.n671 0.037734
R7114 VGND VGND.n2403 0.037734
R7115 VGND.n2396 VGND 0.037734
R7116 VGND.n2391 VGND 0.037734
R7117 VGND.n2386 VGND 0.037734
R7118 VGND.n760 VGND 0.037734
R7119 VGND.n2355 VGND 0.037734
R7120 VGND.n768 VGND 0.037734
R7121 VGND.n2329 VGND 0.037734
R7122 VGND.n776 VGND 0.037734
R7123 VGND.n2303 VGND 0.037734
R7124 VGND.n784 VGND 0.037734
R7125 VGND.n2277 VGND 0.037734
R7126 VGND.n792 VGND 0.037734
R7127 VGND.n2251 VGND 0.037734
R7128 VGND.n804 VGND 0.037734
R7129 VGND VGND.n802 0.037734
R7130 VGND VGND.n2663 0.037734
R7131 VGND.n2656 VGND 0.037734
R7132 VGND.n2373 VGND 0.037734
R7133 VGND.n756 VGND 0.037734
R7134 VGND.n2368 VGND 0.037734
R7135 VGND.n764 VGND 0.037734
R7136 VGND.n2342 VGND 0.037734
R7137 VGND.n772 VGND 0.037734
R7138 VGND.n2316 VGND 0.037734
R7139 VGND.n780 VGND 0.037734
R7140 VGND.n2290 VGND 0.037734
R7141 VGND.n788 VGND 0.037734
R7142 VGND.n2264 VGND 0.037734
R7143 VGND.n796 VGND 0.037734
R7144 VGND.n2238 VGND 0.037734
R7145 VGND VGND.n799 0.037734
R7146 VGND.n2128 VGND 0.037734
R7147 VGND.n2133 VGND 0.037734
R7148 VGND.n867 VGND 0.037734
R7149 VGND.n916 VGND 0.037734
R7150 VGND.n911 VGND 0.037734
R7151 VGND.n906 VGND 0.037734
R7152 VGND.n901 VGND 0.037734
R7153 VGND.n896 VGND 0.037734
R7154 VGND.n891 VGND 0.037734
R7155 VGND.n886 VGND 0.037734
R7156 VGND.n881 VGND 0.037734
R7157 VGND.n876 VGND 0.037734
R7158 VGND.n871 VGND 0.037734
R7159 VGND VGND.n855 0.037734
R7160 VGND.n2153 VGND 0.037734
R7161 VGND VGND.n849 0.037734
R7162 VGND VGND.n2121 0.037734
R7163 VGND.n2114 VGND 0.037734
R7164 VGND.n2109 VGND 0.037734
R7165 VGND.n2104 VGND 0.037734
R7166 VGND.n932 VGND 0.037734
R7167 VGND.n2073 VGND 0.037734
R7168 VGND.n940 VGND 0.037734
R7169 VGND.n2047 VGND 0.037734
R7170 VGND.n948 VGND 0.037734
R7171 VGND.n2021 VGND 0.037734
R7172 VGND.n956 VGND 0.037734
R7173 VGND.n1995 VGND 0.037734
R7174 VGND.n964 VGND 0.037734
R7175 VGND.n1969 VGND 0.037734
R7176 VGND.n1945 VGND 0.037734
R7177 VGND VGND.n1943 0.037734
R7178 VGND VGND.n2688 0.037734
R7179 VGND.n2681 VGND 0.037734
R7180 VGND.n2091 VGND 0.037734
R7181 VGND.n928 VGND 0.037734
R7182 VGND.n2086 VGND 0.037734
R7183 VGND.n936 VGND 0.037734
R7184 VGND.n2060 VGND 0.037734
R7185 VGND.n944 VGND 0.037734
R7186 VGND.n2034 VGND 0.037734
R7187 VGND.n952 VGND 0.037734
R7188 VGND.n2008 VGND 0.037734
R7189 VGND.n960 VGND 0.037734
R7190 VGND.n1982 VGND 0.037734
R7191 VGND.n968 VGND 0.037734
R7192 VGND.n1956 VGND 0.037734
R7193 VGND VGND.n971 0.037734
R7194 VGND.n1901 VGND 0.037734
R7195 VGND.n1906 VGND 0.037734
R7196 VGND.n991 VGND 0.037734
R7197 VGND.n1628 VGND 0.037734
R7198 VGND.n1633 VGND 0.037734
R7199 VGND.n1638 VGND 0.037734
R7200 VGND.n1643 VGND 0.037734
R7201 VGND.n1648 VGND 0.037734
R7202 VGND.n1653 VGND 0.037734
R7203 VGND.n1658 VGND 0.037734
R7204 VGND.n1663 VGND 0.037734
R7205 VGND.n1668 VGND 0.037734
R7206 VGND.n1673 VGND 0.037734
R7207 VGND.n1678 VGND 0.037734
R7208 VGND.n1683 VGND 0.037734
R7209 VGND VGND.n977 0.037734
R7210 VGND VGND.n1894 0.037734
R7211 VGND.n1887 VGND 0.037734
R7212 VGND.n1882 VGND 0.037734
R7213 VGND.n1877 VGND 0.037734
R7214 VGND.n1005 VGND 0.037734
R7215 VGND.n1846 VGND 0.037734
R7216 VGND.n1013 VGND 0.037734
R7217 VGND.n1820 VGND 0.037734
R7218 VGND.n1021 VGND 0.037734
R7219 VGND.n1794 VGND 0.037734
R7220 VGND.n1029 VGND 0.037734
R7221 VGND.n1768 VGND 0.037734
R7222 VGND.n1037 VGND 0.037734
R7223 VGND.n1742 VGND 0.037734
R7224 VGND.n1049 VGND 0.037734
R7225 VGND VGND.n1047 0.037734
R7226 VGND VGND.n2713 0.037734
R7227 VGND.n2706 VGND 0.037734
R7228 VGND.n1864 VGND 0.037734
R7229 VGND.n1001 VGND 0.037734
R7230 VGND.n1859 VGND 0.037734
R7231 VGND.n1009 VGND 0.037734
R7232 VGND.n1833 VGND 0.037734
R7233 VGND.n1017 VGND 0.037734
R7234 VGND.n1807 VGND 0.037734
R7235 VGND.n1025 VGND 0.037734
R7236 VGND.n1781 VGND 0.037734
R7237 VGND.n1033 VGND 0.037734
R7238 VGND.n1755 VGND 0.037734
R7239 VGND.n1041 VGND 0.037734
R7240 VGND.n1729 VGND 0.037734
R7241 VGND VGND.n1044 0.037734
R7242 VGND.n1289 VGND 0.037734
R7243 VGND.n1294 VGND 0.037734
R7244 VGND.n1232 VGND 0.037734
R7245 VGND.n1281 VGND 0.037734
R7246 VGND.n1276 VGND 0.037734
R7247 VGND.n1271 VGND 0.037734
R7248 VGND.n1266 VGND 0.037734
R7249 VGND.n1261 VGND 0.037734
R7250 VGND.n1256 VGND 0.037734
R7251 VGND.n1251 VGND 0.037734
R7252 VGND.n1246 VGND 0.037734
R7253 VGND.n1241 VGND 0.037734
R7254 VGND.n1236 VGND 0.037734
R7255 VGND VGND.n1220 0.037734
R7256 VGND.n1314 VGND 0.037734
R7257 VGND VGND.n1129 0.037734
R7258 VGND.n223 VGND 0.037734
R7259 VGND.n228 VGND 0.037734
R7260 VGND.n233 VGND 0.037734
R7261 VGND.n238 VGND 0.037734
R7262 VGND.n243 VGND 0.037734
R7263 VGND.n248 VGND 0.037734
R7264 VGND.n253 VGND 0.037734
R7265 VGND.n258 VGND 0.037734
R7266 VGND.n263 VGND 0.037734
R7267 VGND.n268 VGND 0.037734
R7268 VGND.n273 VGND 0.037734
R7269 VGND.n278 VGND 0.037734
R7270 VGND.n283 VGND 0.037734
R7271 VGND.n288 VGND 0.037734
R7272 VGND.n293 VGND 0.037734
R7273 VGND VGND.n55 0.037734
R7274 VGND VGND.n1058 0.037734
R7275 VGND VGND.n1061 0.037734
R7276 VGND.n1563 VGND 0.037734
R7277 VGND VGND.n1414 0.037734
R7278 VGND.n1420 VGND 0.037734
R7279 VGND.n1409 VGND 0.037734
R7280 VGND.n1439 VGND 0.037734
R7281 VGND VGND.n1446 0.037734
R7282 VGND.n1452 VGND 0.037734
R7283 VGND.n1118 VGND 0.037734
R7284 VGND.n1471 VGND 0.037734
R7285 VGND VGND.n1478 0.037734
R7286 VGND.n1484 VGND 0.037734
R7287 VGND.n1110 VGND 0.037734
R7288 VGND.n1503 VGND 0.037734
R7289 VGND VGND.n1510 0.037734
R7290 VGND.n1332 VGND 0.037734
R7291 VGND.n1337 VGND 0.037734
R7292 VGND.n1342 VGND 0.037734
R7293 VGND.n1347 VGND 0.037734
R7294 VGND.n1352 VGND 0.037734
R7295 VGND.n1357 VGND 0.037734
R7296 VGND.n1362 VGND 0.037734
R7297 VGND.n1367 VGND 0.037734
R7298 VGND.n1372 VGND 0.037734
R7299 VGND.n1377 VGND 0.037734
R7300 VGND.n1382 VGND 0.037734
R7301 VGND.n1387 VGND 0.037734
R7302 VGND.n1392 VGND 0.037734
R7303 VGND.n1126 VGND 0.037734
R7304 VGND.n1327 VGND 0.037734
R7305 VGND VGND.n1323 0.037734
R7306 VGND.n1623 VGND 0.0343542
R7307 VGND.n1597 VGND 0.0343542
R7308 VGND.n489 VGND 0.0343542
R7309 VGND.n839 VGND 0.0343542
R7310 VGND.n2186 VGND 0.0343542
R7311 VGND.n2223 VGND 0.0343542
R7312 VGND.n1715 VGND 0.0343542
R7313 VGND.n519 VGND 0.0343542
R7314 VGND.n3004 VGND 0.0330521
R7315 VGND.n449 VGND 0.0330521
R7316 VGND.n420 VGND 0.0330521
R7317 VGND.n389 VGND 0.0330521
R7318 VGND.n356 VGND 0.0330521
R7319 VGND VGND.n2900 0.0330521
R7320 VGND VGND.n321 0.0330521
R7321 VGND VGND.n151 0.0330521
R7322 VGND.n3003 VGND 0.024
R7323 VGND.n1 VGND 0.024
R7324 VGND.n488 VGND 0.0239375
R7325 VGND.n838 VGND 0.0239375
R7326 VGND.n518 VGND 0.0239375
R7327 VGND.n388 VGND 0.0239375
R7328 VGND.n355 VGND 0.0239375
R7329 VGND.n1602 VGND 0.0226354
R7330 VGND VGND.n463 0.0226354
R7331 VGND.n2194 VGND 0.0226354
R7332 VGND.n2185 VGND 0.0226354
R7333 VGND.n2197 VGND 0.0226354
R7334 VGND.n350 VGND 0.0226354
R7335 VGND.n2911 VGND 0.0226354
R7336 VGND VGND.n156 0.0226354
R7337 VGND VGND.n813 0.0213333
R7338 VGND.n2190 VGND 0.0213333
R7339 VGND.n1689 VGND 0.0213333
R7340 VGND VGND.n446 0.0213333
R7341 VGND.n448 VGND 0.0213333
R7342 VGND VGND.n415 0.0213333
R7343 VGND.n419 VGND 0.0213333
R7344 VGND VGND.n382 0.0213333
R7345 VGND VGND.n348 0.0213333
R7346 VGND VGND.n2906 0.0213333
R7347 VGND.n3003 VGND 0.0161667
R7348 VGND.n456 VGND 0.0144286
R7349 VGND.n3062 VGND.n3061 0.0105664
R7350 VGND.n2734 VGND 0.00980851
R7351 VGND VGND.n566 0.00980851
R7352 VGND.n2724 VGND 0.00980851
R7353 VGND VGND.n1096 0.00980851
R7354 VGND VGND.n1095 0.00980851
R7355 VGND VGND.n1090 0.00980851
R7356 VGND VGND.n1089 0.00980851
R7357 VGND VGND.n1084 0.00980851
R7358 VGND VGND.n1083 0.00980851
R7359 VGND VGND.n1078 0.00980851
R7360 VGND VGND.n1077 0.00980851
R7361 VGND VGND.n1072 0.00980851
R7362 VGND VGND.n1071 0.00980851
R7363 VGND.n1203 VGND 0.00980851
R7364 VGND VGND.n1137 0.00980851
R7365 VGND.n1136 VGND 0.00980851
R7366 VGND.n221 VGND 0.00980851
R7367 VGND.n2827 VGND 0.00980851
R7368 VGND VGND.n544 0.00980851
R7369 VGND VGND.n543 0.00980851
R7370 VGND VGND.n542 0.00980851
R7371 VGND VGND.n541 0.00980851
R7372 VGND VGND.n540 0.00980851
R7373 VGND VGND.n539 0.00980851
R7374 VGND VGND.n538 0.00980851
R7375 VGND VGND.n537 0.00980851
R7376 VGND VGND.n536 0.00980851
R7377 VGND VGND.n535 0.00980851
R7378 VGND VGND.n534 0.00980851
R7379 VGND VGND.n533 0.00980851
R7380 VGND.n532 VGND 0.00980851
R7381 VGND VGND.n2843 0.00980851
R7382 VGND.n524 VGND 0.00980851
R7383 VGND.n2756 VGND 0.00980851
R7384 VGND.n2620 VGND 0.00980851
R7385 VGND VGND.n616 0.00980851
R7386 VGND VGND.n615 0.00980851
R7387 VGND.n2602 VGND 0.00980851
R7388 VGND.n2579 VGND 0.00980851
R7389 VGND.n2571 VGND 0.00980851
R7390 VGND.n2553 VGND 0.00980851
R7391 VGND.n2545 VGND 0.00980851
R7392 VGND.n2527 VGND 0.00980851
R7393 VGND.n2519 VGND 0.00980851
R7394 VGND.n2501 VGND 0.00980851
R7395 VGND.n2493 VGND 0.00980851
R7396 VGND.n2475 VGND 0.00980851
R7397 VGND.n2467 VGND 0.00980851
R7398 VGND.n2449 VGND 0.00980851
R7399 VGND.n2639 VGND 0.00980851
R7400 VGND VGND.n611 0.00980851
R7401 VGND.n2629 VGND 0.00980851
R7402 VGND VGND.n614 0.00980851
R7403 VGND.n2597 VGND 0.00980851
R7404 VGND.n2584 VGND 0.00980851
R7405 VGND.n2566 VGND 0.00980851
R7406 VGND.n2558 VGND 0.00980851
R7407 VGND.n2540 VGND 0.00980851
R7408 VGND.n2532 VGND 0.00980851
R7409 VGND.n2514 VGND 0.00980851
R7410 VGND.n2506 VGND 0.00980851
R7411 VGND.n2488 VGND 0.00980851
R7412 VGND.n2480 VGND 0.00980851
R7413 VGND.n2462 VGND 0.00980851
R7414 VGND.n2454 VGND 0.00980851
R7415 VGND VGND.n2409 0.00980851
R7416 VGND VGND.n609 0.00980851
R7417 VGND VGND.n608 0.00980851
R7418 VGND.n2421 VGND 0.00980851
R7419 VGND VGND.n683 0.00980851
R7420 VGND VGND.n682 0.00980851
R7421 VGND VGND.n681 0.00980851
R7422 VGND VGND.n680 0.00980851
R7423 VGND VGND.n679 0.00980851
R7424 VGND VGND.n678 0.00980851
R7425 VGND VGND.n677 0.00980851
R7426 VGND VGND.n676 0.00980851
R7427 VGND VGND.n675 0.00980851
R7428 VGND VGND.n674 0.00980851
R7429 VGND VGND.n673 0.00980851
R7430 VGND.n672 VGND 0.00980851
R7431 VGND.n2404 VGND 0.00980851
R7432 VGND VGND.n753 0.00980851
R7433 VGND VGND.n606 0.00980851
R7434 VGND VGND.n605 0.00980851
R7435 VGND.n2384 VGND 0.00980851
R7436 VGND.n2361 VGND 0.00980851
R7437 VGND.n2353 VGND 0.00980851
R7438 VGND.n2335 VGND 0.00980851
R7439 VGND.n2327 VGND 0.00980851
R7440 VGND.n2309 VGND 0.00980851
R7441 VGND.n2301 VGND 0.00980851
R7442 VGND.n2283 VGND 0.00980851
R7443 VGND.n2275 VGND 0.00980851
R7444 VGND.n2257 VGND 0.00980851
R7445 VGND.n2249 VGND 0.00980851
R7446 VGND.n2231 VGND 0.00980851
R7447 VGND.n2664 VGND 0.00980851
R7448 VGND VGND.n599 0.00980851
R7449 VGND.n2654 VGND 0.00980851
R7450 VGND VGND.n603 0.00980851
R7451 VGND.n2379 VGND 0.00980851
R7452 VGND.n2366 VGND 0.00980851
R7453 VGND.n2348 VGND 0.00980851
R7454 VGND.n2340 VGND 0.00980851
R7455 VGND.n2322 VGND 0.00980851
R7456 VGND.n2314 VGND 0.00980851
R7457 VGND.n2296 VGND 0.00980851
R7458 VGND.n2288 VGND 0.00980851
R7459 VGND.n2270 VGND 0.00980851
R7460 VGND.n2262 VGND 0.00980851
R7461 VGND.n2244 VGND 0.00980851
R7462 VGND.n2236 VGND 0.00980851
R7463 VGND VGND.n2127 0.00980851
R7464 VGND VGND.n597 0.00980851
R7465 VGND VGND.n596 0.00980851
R7466 VGND.n2139 VGND 0.00980851
R7467 VGND VGND.n865 0.00980851
R7468 VGND VGND.n864 0.00980851
R7469 VGND VGND.n863 0.00980851
R7470 VGND VGND.n862 0.00980851
R7471 VGND VGND.n861 0.00980851
R7472 VGND VGND.n860 0.00980851
R7473 VGND VGND.n859 0.00980851
R7474 VGND VGND.n858 0.00980851
R7475 VGND VGND.n857 0.00980851
R7476 VGND.n856 VGND 0.00980851
R7477 VGND VGND.n2152 0.00980851
R7478 VGND.n850 VGND 0.00980851
R7479 VGND.n2122 VGND 0.00980851
R7480 VGND VGND.n925 0.00980851
R7481 VGND VGND.n594 0.00980851
R7482 VGND VGND.n593 0.00980851
R7483 VGND.n2102 VGND 0.00980851
R7484 VGND.n2079 VGND 0.00980851
R7485 VGND.n2071 VGND 0.00980851
R7486 VGND.n2053 VGND 0.00980851
R7487 VGND.n2045 VGND 0.00980851
R7488 VGND.n2027 VGND 0.00980851
R7489 VGND.n2019 VGND 0.00980851
R7490 VGND.n2001 VGND 0.00980851
R7491 VGND.n1993 VGND 0.00980851
R7492 VGND.n1975 VGND 0.00980851
R7493 VGND.n1967 VGND 0.00980851
R7494 VGND.n1949 VGND 0.00980851
R7495 VGND.n2689 VGND 0.00980851
R7496 VGND VGND.n587 0.00980851
R7497 VGND.n2679 VGND 0.00980851
R7498 VGND VGND.n591 0.00980851
R7499 VGND.n2097 VGND 0.00980851
R7500 VGND.n2084 VGND 0.00980851
R7501 VGND.n2066 VGND 0.00980851
R7502 VGND.n2058 VGND 0.00980851
R7503 VGND.n2040 VGND 0.00980851
R7504 VGND.n2032 VGND 0.00980851
R7505 VGND.n2014 VGND 0.00980851
R7506 VGND.n2006 VGND 0.00980851
R7507 VGND.n1988 VGND 0.00980851
R7508 VGND.n1980 VGND 0.00980851
R7509 VGND.n1962 VGND 0.00980851
R7510 VGND.n1954 VGND 0.00980851
R7511 VGND VGND.n1900 0.00980851
R7512 VGND VGND.n585 0.00980851
R7513 VGND VGND.n584 0.00980851
R7514 VGND.n1912 VGND 0.00980851
R7515 VGND VGND.n989 0.00980851
R7516 VGND VGND.n988 0.00980851
R7517 VGND VGND.n987 0.00980851
R7518 VGND VGND.n986 0.00980851
R7519 VGND VGND.n985 0.00980851
R7520 VGND VGND.n984 0.00980851
R7521 VGND VGND.n983 0.00980851
R7522 VGND VGND.n982 0.00980851
R7523 VGND VGND.n981 0.00980851
R7524 VGND VGND.n980 0.00980851
R7525 VGND VGND.n979 0.00980851
R7526 VGND.n978 VGND 0.00980851
R7527 VGND.n1895 VGND 0.00980851
R7528 VGND VGND.n998 0.00980851
R7529 VGND VGND.n582 0.00980851
R7530 VGND VGND.n581 0.00980851
R7531 VGND.n1875 VGND 0.00980851
R7532 VGND.n1852 VGND 0.00980851
R7533 VGND.n1844 VGND 0.00980851
R7534 VGND.n1826 VGND 0.00980851
R7535 VGND.n1818 VGND 0.00980851
R7536 VGND.n1800 VGND 0.00980851
R7537 VGND.n1792 VGND 0.00980851
R7538 VGND.n1774 VGND 0.00980851
R7539 VGND.n1766 VGND 0.00980851
R7540 VGND.n1748 VGND 0.00980851
R7541 VGND.n1740 VGND 0.00980851
R7542 VGND.n1722 VGND 0.00980851
R7543 VGND.n2714 VGND 0.00980851
R7544 VGND VGND.n574 0.00980851
R7545 VGND.n2704 VGND 0.00980851
R7546 VGND VGND.n578 0.00980851
R7547 VGND.n1870 VGND 0.00980851
R7548 VGND.n1857 VGND 0.00980851
R7549 VGND.n1839 VGND 0.00980851
R7550 VGND.n1831 VGND 0.00980851
R7551 VGND.n1813 VGND 0.00980851
R7552 VGND.n1805 VGND 0.00980851
R7553 VGND.n1787 VGND 0.00980851
R7554 VGND.n1779 VGND 0.00980851
R7555 VGND.n1761 VGND 0.00980851
R7556 VGND.n1753 VGND 0.00980851
R7557 VGND.n1735 VGND 0.00980851
R7558 VGND.n1727 VGND 0.00980851
R7559 VGND VGND.n1288 0.00980851
R7560 VGND VGND.n570 0.00980851
R7561 VGND VGND.n569 0.00980851
R7562 VGND.n1300 VGND 0.00980851
R7563 VGND VGND.n1230 0.00980851
R7564 VGND VGND.n1229 0.00980851
R7565 VGND VGND.n1228 0.00980851
R7566 VGND VGND.n1227 0.00980851
R7567 VGND VGND.n1226 0.00980851
R7568 VGND VGND.n1225 0.00980851
R7569 VGND VGND.n1224 0.00980851
R7570 VGND VGND.n1223 0.00980851
R7571 VGND VGND.n1222 0.00980851
R7572 VGND.n1221 VGND 0.00980851
R7573 VGND VGND.n1313 0.00980851
R7574 VGND.n1130 VGND 0.00980851
R7575 VGND.n3011 VGND 0.00980851
R7576 VGND VGND.n98 0.00980851
R7577 VGND VGND.n93 0.00980851
R7578 VGND VGND.n92 0.00980851
R7579 VGND VGND.n87 0.00980851
R7580 VGND VGND.n86 0.00980851
R7581 VGND VGND.n81 0.00980851
R7582 VGND VGND.n80 0.00980851
R7583 VGND VGND.n75 0.00980851
R7584 VGND VGND.n74 0.00980851
R7585 VGND VGND.n69 0.00980851
R7586 VGND VGND.n68 0.00980851
R7587 VGND VGND.n63 0.00980851
R7588 VGND VGND.n62 0.00980851
R7589 VGND VGND.n57 0.00980851
R7590 VGND.n56 VGND 0.00980851
R7591 VGND.n1569 VGND 0.00980851
R7592 VGND.n1062 VGND 0.00980851
R7593 VGND VGND.n1562 0.00980851
R7594 VGND.n1418 VGND 0.00980851
R7595 VGND.n1426 VGND 0.00980851
R7596 VGND.n1437 VGND 0.00980851
R7597 VGND VGND.n1121 0.00980851
R7598 VGND.n1450 VGND 0.00980851
R7599 VGND.n1458 VGND 0.00980851
R7600 VGND.n1469 VGND 0.00980851
R7601 VGND VGND.n1113 0.00980851
R7602 VGND.n1482 VGND 0.00980851
R7603 VGND.n1490 VGND 0.00980851
R7604 VGND.n1501 VGND 0.00980851
R7605 VGND VGND.n1105 0.00980851
R7606 VGND.n1511 VGND 0.00980851
R7607 VGND.n2739 VGND 0.00980851
R7608 VGND VGND.n1100 0.00980851
R7609 VGND VGND.n1099 0.00980851
R7610 VGND VGND.n1098 0.00980851
R7611 VGND VGND.n1093 0.00980851
R7612 VGND VGND.n1092 0.00980851
R7613 VGND VGND.n1087 0.00980851
R7614 VGND VGND.n1086 0.00980851
R7615 VGND VGND.n1081 0.00980851
R7616 VGND VGND.n1080 0.00980851
R7617 VGND VGND.n1075 0.00980851
R7618 VGND VGND.n1074 0.00980851
R7619 VGND VGND.n1069 0.00980851
R7620 VGND VGND.n1068 0.00980851
R7621 VGND.n1398 VGND 0.00980851
R7622 VGND.n1325 VGND 0.00980851
R7623 VGND.n3063 VGND 0.00835714
R7624 VGND.n2999 VGND.n2998 0.00182979
R7625 VGND.n2991 VGND.n205 0.00182979
R7626 VGND.n2989 VGND.n2988 0.00182979
R7627 VGND.n2981 VGND.n207 0.00182979
R7628 VGND.n2979 VGND.n2978 0.00182979
R7629 VGND.n2971 VGND.n209 0.00182979
R7630 VGND.n2969 VGND.n2968 0.00182979
R7631 VGND.n2961 VGND.n211 0.00182979
R7632 VGND.n2959 VGND.n2958 0.00182979
R7633 VGND.n2951 VGND.n213 0.00182979
R7634 VGND.n2949 VGND.n2948 0.00182979
R7635 VGND.n2941 VGND.n215 0.00182979
R7636 VGND.n2939 VGND.n2938 0.00182979
R7637 VGND.n2931 VGND.n217 0.00182979
R7638 VGND.n2929 VGND.n2928 0.00182979
R7639 XThR.Tn[2].n2 XThR.Tn[2].n0 332.332
R7640 XThR.Tn[2].n2 XThR.Tn[2].n1 296.493
R7641 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7642 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7643 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7644 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7645 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7646 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7647 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7648 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7649 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7650 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7651 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7652 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7653 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7654 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7655 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7656 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7657 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7658 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7659 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7660 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7661 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7662 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7663 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7664 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7665 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7666 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7667 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7668 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7669 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7670 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7671 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7672 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7673 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7674 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7675 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7676 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7677 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7678 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7679 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7680 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7681 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7682 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7683 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7684 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7685 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7686 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7687 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7688 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7689 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7690 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7691 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7692 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7693 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7694 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7695 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7696 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7697 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7698 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7699 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7700 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7701 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7702 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7703 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7704 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7705 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7706 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7707 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7708 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7709 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7710 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7711 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7712 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7713 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7714 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7715 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7716 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7717 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7718 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7719 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7720 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7721 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7722 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7723 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7724 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7725 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7726 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7727 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7728 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7729 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7730 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7731 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7732 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7733 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7734 XThR.Tn[2].n5 XThR.Tn[2].n3 135.249
R7735 XThR.Tn[2].n5 XThR.Tn[2].n4 98.982
R7736 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R7737 XThR.Tn[2].n9 XThR.Tn[2].n8 98.982
R7738 XThR.Tn[2].n7 XThR.Tn[2].n5 36.2672
R7739 XThR.Tn[2].n9 XThR.Tn[2].n7 36.2672
R7740 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7741 XThR.Tn[2].n0 XThR.Tn[2].t9 26.5955
R7742 XThR.Tn[2].n0 XThR.Tn[2].t4 26.5955
R7743 XThR.Tn[2].n1 XThR.Tn[2].t11 26.5955
R7744 XThR.Tn[2].n1 XThR.Tn[2].t0 26.5955
R7745 XThR.Tn[2].n3 XThR.Tn[2].t7 24.9236
R7746 XThR.Tn[2].n3 XThR.Tn[2].t8 24.9236
R7747 XThR.Tn[2].n4 XThR.Tn[2].t6 24.9236
R7748 XThR.Tn[2].n4 XThR.Tn[2].t5 24.9236
R7749 XThR.Tn[2].n6 XThR.Tn[2].t3 24.9236
R7750 XThR.Tn[2].n6 XThR.Tn[2].t1 24.9236
R7751 XThR.Tn[2].n8 XThR.Tn[2].t10 24.9236
R7752 XThR.Tn[2].n8 XThR.Tn[2].t2 24.9236
R7753 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7754 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7755 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7756 XThR.Tn[2] XThR.Tn[2].n11 5.4407
R7757 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7758 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7759 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7760 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7761 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7762 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7763 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7764 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7765 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7766 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7767 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7768 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7769 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7770 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7771 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7772 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7773 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7774 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7775 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7776 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7777 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7778 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7779 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7780 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7781 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7782 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7783 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7784 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7785 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7786 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7787 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7788 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7789 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7790 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7791 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7792 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7793 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7794 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7795 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7796 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7797 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7798 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7799 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7800 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7801 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7802 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7803 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7804 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7805 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7806 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7807 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7808 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7809 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7810 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7811 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7812 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7813 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7814 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7815 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7816 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7817 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7818 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7819 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7820 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7821 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7822 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7823 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7824 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7825 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7826 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7827 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7828 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7829 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7830 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7831 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7832 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7833 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7834 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7835 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7836 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7837 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7838 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7839 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7840 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7841 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7842 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7843 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7844 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7845 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7846 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7847 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7848 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7849 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7850 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7851 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7852 VPWR.n3110 VPWR.n29 3532.94
R7853 VPWR.n3110 VPWR.n30 3532.94
R7854 VPWR.n3119 VPWR.n29 3532.94
R7855 VPWR.n3119 VPWR.n30 3532.94
R7856 VPWR.n3108 VPWR.n27 3532.94
R7857 VPWR.n3108 VPWR.n28 3532.94
R7858 VPWR.n3121 VPWR.n27 3532.94
R7859 VPWR.n3121 VPWR.n28 3532.94
R7860 VPWR.n2662 VPWR.t1225 1005.7
R7861 VPWR.n2493 VPWR.t1443 1005.7
R7862 VPWR.n537 VPWR.t1292 1005.7
R7863 VPWR.n2353 VPWR.t1409 1005.7
R7864 VPWR.t1126 VPWR.n2258 1005.7
R7865 VPWR.t1233 VPWR.n2238 1005.7
R7866 VPWR.n2226 VPWR.t1193 1005.7
R7867 VPWR.t1298 VPWR.n2025 1005.7
R7868 VPWR.t1118 VPWR.n1995 1005.7
R7869 VPWR.t1305 VPWR.n834 1005.7
R7870 VPWR.t1110 VPWR.n2603 1005.7
R7871 VPWR.n1858 VPWR.t1419 1005.7
R7872 VPWR.n2673 VPWR.t1404 1005.7
R7873 VPWR.n1722 VPWR.t1265 1005.7
R7874 VPWR.n1712 VPWR.t1388 1005.7
R7875 VPWR.n317 VPWR.t1435 1005.7
R7876 VPWR.t1211 VPWR.n1587 1005.7
R7877 VPWR.n2847 VPWR.t1330 1005.7
R7878 VPWR.t796 VPWR.n492 983.14
R7879 VPWR.n496 VPWR.t1629 983.14
R7880 VPWR.n495 VPWR.t1538 983.14
R7881 VPWR.n2541 VPWR.t732 983.14
R7882 VPWR.n2540 VPWR.t161 983.14
R7883 VPWR.n2534 VPWR.t169 983.14
R7884 VPWR.n2533 VPWR.t481 983.14
R7885 VPWR.t518 VPWR.n2513 983.14
R7886 VPWR.t120 VPWR.n2516 983.14
R7887 VPWR.n2521 VPWR.t362 983.14
R7888 VPWR.n2520 VPWR.t1577 983.14
R7889 VPWR.t1600 VPWR.n2646 983.14
R7890 VPWR.n2647 VPWR.t189 983.14
R7891 VPWR.t12 VPWR.n2658 983.14
R7892 VPWR.t582 VPWR.n2661 983.14
R7893 VPWR.n486 VPWR.t1691 983.14
R7894 VPWR.t254 VPWR.n2426 983.14
R7895 VPWR.n2427 VPWR.t1514 983.14
R7896 VPWR.t1062 VPWR.n2433 983.14
R7897 VPWR.t498 VPWR.n2436 983.14
R7898 VPWR.n2442 VPWR.t1881 983.14
R7899 VPWR.n2441 VPWR.t68 983.14
R7900 VPWR.t866 VPWR.n2464 983.14
R7901 VPWR.n2465 VPWR.t1573 983.14
R7902 VPWR.t301 VPWR.n2471 983.14
R7903 VPWR.t1008 VPWR.n2476 983.14
R7904 VPWR.n2477 VPWR.t902 983.14
R7905 VPWR.t202 VPWR.n2484 983.14
R7906 VPWR.n2485 VPWR.t969 983.14
R7907 VPWR.t992 VPWR.n2492 983.14
R7908 VPWR.t702 VPWR.n509 983.14
R7909 VPWR.t939 VPWR.n512 983.14
R7910 VPWR.n2407 VPWR.t1492 983.14
R7911 VPWR.n2406 VPWR.t820 983.14
R7912 VPWR.n2400 VPWR.t1584 983.14
R7913 VPWR.n2399 VPWR.t1851 983.14
R7914 VPWR.n2393 VPWR.t1841 983.14
R7915 VPWR.n2392 VPWR.t54 983.14
R7916 VPWR.n2386 VPWR.t670 983.14
R7917 VPWR.n2385 VPWR.t1895 983.14
R7918 VPWR.n2379 VPWR.t747 983.14
R7919 VPWR.n2378 VPWR.t1606 983.14
R7920 VPWR.t1472 VPWR.n533 983.14
R7921 VPWR.n2367 VPWR.t1707 983.14
R7922 VPWR.n2366 VPWR.t1722 983.14
R7923 VPWR.t252 VPWR.n688 983.14
R7924 VPWR.n696 VPWR.t508 983.14
R7925 VPWR.n695 VPWR.t1506 983.14
R7926 VPWR.n691 VPWR.t1068 983.14
R7927 VPWR.n2288 VPWR.t1779 983.14
R7928 VPWR.n2287 VPWR.t432 983.14
R7929 VPWR.n571 VPWR.t78 983.14
R7930 VPWR.n570 VPWR.t719 983.14
R7931 VPWR.t887 VPWR.n2311 983.14
R7932 VPWR.t307 VPWR.n2314 983.14
R7933 VPWR.n2328 VPWR.t1018 983.14
R7934 VPWR.n2327 VPWR.t1822 983.14
R7935 VPWR.n2321 VPWR.t210 983.14
R7936 VPWR.n2320 VPWR.t1633 983.14
R7937 VPWR.t998 VPWR.n2352 983.14
R7938 VPWR.t248 VPWR.n632 983.14
R7939 VPWR.n680 VPWR.t961 983.14
R7940 VPWR.n679 VPWR.t1526 983.14
R7941 VPWR.n673 VPWR.t1793 983.14
R7942 VPWR.n672 VPWR.t1742 983.14
R7943 VPWR.n668 VPWR.t407 983.14
R7944 VPWR.n662 VPWR.t465 983.14
R7945 VPWR.n661 VPWR.t110 983.14
R7946 VPWR.n655 VPWR.t421 983.14
R7947 VPWR.n654 VPWR.t265 983.14
R7948 VPWR.n648 VPWR.t1022 983.14
R7949 VPWR.n647 VPWR.t908 983.14
R7950 VPWR.n2266 VPWR.t1052 983.14
R7951 VPWR.n2265 VPWR.t1905 983.14
R7952 VPWR.n2259 VPWR.t524 983.14
R7953 VPWR.n625 VPWR.t794 983.14
R7954 VPWR.t1627 VPWR.n2139 983.14
R7955 VPWR.n2143 VPWR.t1540 983.14
R7956 VPWR.n2142 VPWR.t730 983.14
R7957 VPWR.t159 VPWR.n2156 983.14
R7958 VPWR.n2157 VPWR.t167 983.14
R7959 VPWR.t479 VPWR.n2168 983.14
R7960 VPWR.n2169 VPWR.t516 983.14
R7961 VPWR.t662 VPWR.n2180 983.14
R7962 VPWR.t360 VPWR.n2183 983.14
R7963 VPWR.n2196 VPWR.t1575 983.14
R7964 VPWR.n2195 VPWR.t1598 983.14
R7965 VPWR.n2189 VPWR.t187 983.14
R7966 VPWR.n2188 VPWR.t10 983.14
R7967 VPWR.n2239 VPWR.t580 983.14
R7968 VPWR.n2072 VPWR.t1687 983.14
R7969 VPWR.t774 VPWR.n2078 983.14
R7970 VPWR.n2079 VPWR.t1534 983.14
R7971 VPWR.t734 VPWR.n2086 983.14
R7972 VPWR.t1699 VPWR.n2089 983.14
R7973 VPWR.n2114 VPWR.t1802 983.14
R7974 VPWR.n2113 VPWR.t461 983.14
R7975 VPWR.n2107 VPWR.t650 983.14
R7976 VPWR.n2106 VPWR.t126 983.14
R7977 VPWR.n2100 VPWR.t368 983.14
R7978 VPWR.n2099 VPWR.t765 983.14
R7979 VPWR.t1812 VPWR.n2214 983.14
R7980 VPWR.n2215 VPWR.t191 983.14
R7981 VPWR.t18 VPWR.n2222 983.14
R7982 VPWR.t584 VPWR.n2225 983.14
R7983 VPWR.n1923 VPWR.t700 983.14
R7984 VPWR.t937 VPWR.n1933 983.14
R7985 VPWR.t1494 VPWR.n1936 983.14
R7986 VPWR.n1944 VPWR.t816 983.14
R7987 VPWR.n1943 VPWR.t1582 983.14
R7988 VPWR.n1939 VPWR.t1849 983.14
R7989 VPWR.n2057 VPWR.t1839 983.14
R7990 VPWR.n2056 VPWR.t808 983.14
R7991 VPWR.t668 VPWR.n723 983.14
R7992 VPWR.n2045 VPWR.t1893 983.14
R7993 VPWR.n2044 VPWR.t745 983.14
R7994 VPWR.n2038 VPWR.t1604 983.14
R7995 VPWR.n2037 VPWR.t1468 983.14
R7996 VPWR.t1705 VPWR.n735 983.14
R7997 VPWR.n2026 VPWR.t1718 983.14
R7998 VPWR.t1564 VPWR.n770 983.14
R7999 VPWR.n790 VPWR.t963 983.14
R8000 VPWR.n789 VPWR.t1524 983.14
R8001 VPWR.n783 VPWR.t707 983.14
R8002 VPWR.n782 VPWR.t1744 983.14
R8003 VPWR.n776 VPWR.t409 983.14
R8004 VPWR.t467 VPWR.n1963 983.14
R8005 VPWR.n1964 VPWR.t112 983.14
R8006 VPWR.t566 VPWR.n1971 983.14
R8007 VPWR.n1972 VPWR.t267 983.14
R8008 VPWR.t1024 VPWR.n1987 983.14
R8009 VPWR.t910 VPWR.n1990 983.14
R8010 VPWR.n2003 VPWR.t1054 983.14
R8011 VPWR.n2002 VPWR.t1907 983.14
R8012 VPWR.n1996 VPWR.t526 983.14
R8013 VPWR.t698 VPWR.n802 983.14
R8014 VPWR.t1623 VPWR.n805 983.14
R8015 VPWR.n1909 VPWR.t1496 983.14
R8016 VPWR.n1908 VPWR.t814 983.14
R8017 VPWR.n1902 VPWR.t924 983.14
R8018 VPWR.n1901 VPWR.t1847 983.14
R8019 VPWR.t1837 VPWR.n819 983.14
R8020 VPWR.t804 VPWR.n822 983.14
R8021 VPWR.n1889 VPWR.t666 983.14
R8022 VPWR.n1888 VPWR.t1891 983.14
R8023 VPWR.n1882 VPWR.t220 983.14
R8024 VPWR.n1881 VPWR.t1614 983.14
R8025 VPWR.n1875 VPWR.t1464 983.14
R8026 VPWR.n1874 VPWR.t1703 983.14
R8027 VPWR.n835 VPWR.t1716 983.14
R8028 VPWR.t1566 VPWR.n2555 983.14
R8029 VPWR.t965 VPWR.n2558 983.14
R8030 VPWR.n2564 VPWR.t1522 983.14
R8031 VPWR.n2563 VPWR.t711 983.14
R8032 VPWR.t1746 VPWR.n2581 983.14
R8033 VPWR.n2582 VPWR.t411 983.14
R8034 VPWR.t469 VPWR.n2589 983.14
R8035 VPWR.t0 VPWR.n2592 983.14
R8036 VPWR.n2625 VPWR.t568 983.14
R8037 VPWR.n2624 VPWR.t269 983.14
R8038 VPWR.n2618 VPWR.t1026 983.14
R8039 VPWR.n2617 VPWR.t1542 983.14
R8040 VPWR.n2611 VPWR.t1056 983.14
R8041 VPWR.n2610 VPWR.t1909 983.14
R8042 VPWR.n2604 VPWR.t530 983.14
R8043 VPWR.t250 VPWR.n1780 983.14
R8044 VPWR.n1781 VPWR.t504 983.14
R8045 VPWR.t1508 VPWR.n1787 983.14
R8046 VPWR.t1066 VPWR.n1790 983.14
R8047 VPWR.n1799 VPWR.t1775 983.14
R8048 VPWR.n1798 VPWR.t428 983.14
R8049 VPWR.n1793 VPWR.t74 983.14
R8050 VPWR.t717 VPWR.n1822 983.14
R8051 VPWR.n1823 VPWR.t1042 983.14
R8052 VPWR.t305 VPWR.n1834 983.14
R8053 VPWR.n1838 VPWR.t1014 983.14
R8054 VPWR.n1837 VPWR.t1820 983.14
R8055 VPWR.t208 VPWR.n1849 983.14
R8056 VPWR.n1850 VPWR.t1631 983.14
R8057 VPWR.t996 VPWR.n1857 983.14
R8058 VPWR.t483 VPWR.n376 983.14
R8059 VPWR.n2732 VPWR.t510 983.14
R8060 VPWR.n2731 VPWR.t1504 983.14
R8061 VPWR.t1072 VPWR.n385 983.14
R8062 VPWR.n2720 VPWR.t1781 983.14
R8063 VPWR.n2719 VPWR.t434 983.14
R8064 VPWR.t80 VPWR.n394 983.14
R8065 VPWR.n2708 VPWR.t721 983.14
R8066 VPWR.n2707 VPWR.t889 983.14
R8067 VPWR.t309 VPWR.n403 983.14
R8068 VPWR.n2696 VPWR.t1020 983.14
R8069 VPWR.n2695 VPWR.t1824 983.14
R8070 VPWR.t212 VPWR.n412 983.14
R8071 VPWR.n2684 VPWR.t1635 983.14
R8072 VPWR.n2683 VPWR.t1002 983.14
R8073 VPWR.t704 VPWR.n880 983.14
R8074 VPWR.t945 VPWR.n883 983.14
R8075 VPWR.n1767 VPWR.t1486 983.14
R8076 VPWR.n1766 VPWR.t826 983.14
R8077 VPWR.n1760 VPWR.t1590 983.14
R8078 VPWR.n1759 VPWR.t1857 983.14
R8079 VPWR.t1767 VPWR.n900 983.14
R8080 VPWR.t58 VPWR.n903 983.14
R8081 VPWR.n1747 VPWR.t656 983.14
R8082 VPWR.n1746 VPWR.t1897 983.14
R8083 VPWR.n1740 VPWR.t753 983.14
R8084 VPWR.n1739 VPWR.t1608 983.14
R8085 VPWR.n1733 VPWR.t1476 983.14
R8086 VPWR.n1732 VPWR.t20 983.14
R8087 VPWR.t576 VPWR.n1721 983.14
R8088 VPWR.t1321 VPWR.n1191 983.14
R8089 VPWR.n1192 VPWR.t1448 983.14
R8090 VPWR.t1219 VPWR.n1199 983.14
R8091 VPWR.t1324 VPWR.n1205 983.14
R8092 VPWR.n1659 VPWR.t1346 983.14
R8093 VPWR.n1658 VPWR.t1094 983.14
R8094 VPWR.n1652 VPWR.t1216 983.14
R8095 VPWR.n1651 VPWR.t1357 983.14
R8096 VPWR.n1645 VPWR.t1385 983.14
R8097 VPWR.n1644 VPWR.t1113 983.14
R8098 VPWR.t1246 VPWR.n1625 983.14
R8099 VPWR.n1632 VPWR.t1287 983.14
R8100 VPWR.n1631 VPWR.t1123 983.14
R8101 VPWR.t1157 VPWR.n1705 983.14
R8102 VPWR.t1268 VPWR.n1711 983.14
R8103 VPWR.t1693 VPWR.n295 983.14
R8104 VPWR.n365 VPWR.t256 983.14
R8105 VPWR.n364 VPWR.t1512 983.14
R8106 VPWR.n358 VPWR.t1064 983.14
R8107 VPWR.n357 VPWR.t500 983.14
R8108 VPWR.n351 VPWR.t1883 983.14
R8109 VPWR.n350 VPWR.t70 983.14
R8110 VPWR.n344 VPWR.t870 983.14
R8111 VPWR.n343 VPWR.t1038 983.14
R8112 VPWR.n337 VPWR.t303 983.14
R8113 VPWR.n336 VPWR.t1010 983.14
R8114 VPWR.n330 VPWR.t904 983.14
R8115 VPWR.n329 VPWR.t206 983.14
R8116 VPWR.n323 VPWR.t971 983.14
R8117 VPWR.n322 VPWR.t994 983.14
R8118 VPWR.t1160 VPWR.n1163 983.14
R8119 VPWR.n1672 VPWR.t1262 983.14
R8120 VPWR.n1671 VPWR.t1424 983.14
R8121 VPWR.n1278 VPWR.t1142 983.14
R8122 VPWR.t1154 VPWR.n1488 983.14
R8123 VPWR.n1489 VPWR.t1313 983.14
R8124 VPWR.t1363 VPWR.n1500 983.14
R8125 VPWR.n1501 VPWR.t1182 983.14
R8126 VPWR.t1208 VPWR.n1514 983.14
R8127 VPWR.n1515 VPWR.t1338 983.14
R8128 VPWR.t1081 VPWR.n1523 983.14
R8129 VPWR.n1532 VPWR.t1102 983.14
R8130 VPWR.n1531 VPWR.t1343 983.14
R8131 VPWR.n1526 VPWR.t1377 983.14
R8132 VPWR.n1588 VPWR.t1088 983.14
R8133 VPWR.t1274 VPWR.n2762 983.14
R8134 VPWR.n2763 VPWR.t1395 983.14
R8135 VPWR.t1151 VPWR.n2774 983.14
R8136 VPWR.n2775 VPWR.t1259 983.14
R8137 VPWR.t1271 VPWR.n2786 983.14
R8138 VPWR.n2787 VPWR.t1427 983.14
R8139 VPWR.t1148 VPWR.n2798 983.14
R8140 VPWR.n2799 VPWR.t1308 983.14
R8141 VPWR.t1327 VPWR.n2810 983.14
R8142 VPWR.n2811 VPWR.t1454 983.14
R8143 VPWR.t1198 VPWR.n2822 983.14
R8144 VPWR.n2823 VPWR.t1228 983.14
R8145 VPWR.t1078 VPWR.n2834 983.14
R8146 VPWR.n2835 VPWR.t1097 983.14
R8147 VPWR.t1222 VPWR.n2846 983.14
R8148 VPWR.n1016 VPWR.t340 877.144
R8149 VPWR.n3012 VPWR.t982 877.144
R8150 VPWR.n906 VPWR.t1898 738.074
R8151 VPWR.n904 VPWR.t657 738.074
R8152 VPWR.n895 VPWR.t59 738.074
R8153 VPWR.n901 VPWR.t1768 738.074
R8154 VPWR.n896 VPWR.t1858 738.074
R8155 VPWR.n887 VPWR.t1591 738.074
R8156 VPWR.n858 VPWR.t718 738.074
R8157 VPWR.n859 VPWR.t75 738.074
R8158 VPWR.n459 VPWR.t170 738.074
R8159 VPWR.n458 VPWR.t162 738.074
R8160 VPWR.n456 VPWR.t733 738.074
R8161 VPWR.n455 VPWR.t1539 738.074
R8162 VPWR.n493 VPWR.t1630 738.074
R8163 VPWR.n491 VPWR.t797 738.074
R8164 VPWR.n489 VPWR.t620 738.074
R8165 VPWR.n2509 VPWR.t482 738.074
R8166 VPWR.n2514 VPWR.t519 738.074
R8167 VPWR.n2508 VPWR.t121 738.074
R8168 VPWR.n2517 VPWR.t363 738.074
R8169 VPWR.n430 VPWR.t1578 738.074
R8170 VPWR.n429 VPWR.t1601 738.074
R8171 VPWR.n423 VPWR.t190 738.074
R8172 VPWR.n2659 VPWR.t13 738.074
R8173 VPWR.n422 VPWR.t583 738.074
R8174 VPWR.n2437 VPWR.t1882 738.074
R8175 VPWR.n481 VPWR.t499 738.074
R8176 VPWR.n2434 VPWR.t1063 738.074
R8177 VPWR.n482 VPWR.t1515 738.074
R8178 VPWR.n483 VPWR.t255 738.074
R8179 VPWR.n484 VPWR.t1692 738.074
R8180 VPWR.n485 VPWR.t610 738.074
R8181 VPWR.n473 VPWR.t69 738.074
R8182 VPWR.n472 VPWR.t867 738.074
R8183 VPWR.n471 VPWR.t1574 738.074
R8184 VPWR.n2472 VPWR.t302 738.074
R8185 VPWR.n470 VPWR.t1009 738.074
R8186 VPWR.n469 VPWR.t903 738.074
R8187 VPWR.n468 VPWR.t203 738.074
R8188 VPWR.n467 VPWR.t970 738.074
R8189 VPWR.n466 VPWR.t993 738.074
R8190 VPWR.n518 VPWR.t1852 738.074
R8191 VPWR.n516 VPWR.t1585 738.074
R8192 VPWR.n515 VPWR.t821 738.074
R8193 VPWR.n513 VPWR.t1493 738.074
R8194 VPWR.n505 VPWR.t940 738.074
R8195 VPWR.n510 VPWR.t703 738.074
R8196 VPWR.n506 VPWR.t596 738.074
R8197 VPWR.n519 VPWR.t1842 738.074
R8198 VPWR.n521 VPWR.t55 738.074
R8199 VPWR.n522 VPWR.t671 738.074
R8200 VPWR.n524 VPWR.t1896 738.074
R8201 VPWR.n525 VPWR.t748 738.074
R8202 VPWR.n531 VPWR.t1607 738.074
R8203 VPWR.n530 VPWR.t1473 738.074
R8204 VPWR.n534 VPWR.t1708 738.074
R8205 VPWR.n536 VPWR.t1723 738.074
R8206 VPWR.n567 VPWR.t433 738.074
R8207 VPWR.n566 VPWR.t1780 738.074
R8208 VPWR.n565 VPWR.t1069 738.074
R8209 VPWR.n689 VPWR.t1507 738.074
R8210 VPWR.n692 VPWR.t509 738.074
R8211 VPWR.n687 VPWR.t253 738.074
R8212 VPWR.n684 VPWR.t604 738.074
R8213 VPWR.n568 VPWR.t79 738.074
R8214 VPWR.n555 VPWR.t720 738.074
R8215 VPWR.n2312 VPWR.t888 738.074
R8216 VPWR.n554 VPWR.t308 738.074
R8217 VPWR.n2315 VPWR.t1019 738.074
R8218 VPWR.n2317 VPWR.t1823 738.074
R8219 VPWR.n2318 VPWR.t211 738.074
R8220 VPWR.n543 VPWR.t1634 738.074
R8221 VPWR.n542 VPWR.t999 738.074
R8222 VPWR.n638 VPWR.t408 738.074
R8223 VPWR.n636 VPWR.t1743 738.074
R8224 VPWR.n669 VPWR.t1794 738.074
R8225 VPWR.n635 VPWR.t1527 738.074
R8226 VPWR.n633 VPWR.t962 738.074
R8227 VPWR.n631 VPWR.t249 738.074
R8228 VPWR.n628 VPWR.t616 738.074
R8229 VPWR.n639 VPWR.t466 738.074
R8230 VPWR.n641 VPWR.t111 738.074
R8231 VPWR.n642 VPWR.t422 738.074
R8232 VPWR.n644 VPWR.t266 738.074
R8233 VPWR.n645 VPWR.t1023 738.074
R8234 VPWR.n580 VPWR.t909 738.074
R8235 VPWR.n581 VPWR.t1053 738.074
R8236 VPWR.n2254 VPWR.t1906 738.074
R8237 VPWR.n2255 VPWR.t525 738.074
R8238 VPWR.n611 VPWR.t168 738.074
R8239 VPWR.n614 VPWR.t160 738.074
R8240 VPWR.n615 VPWR.t731 738.074
R8241 VPWR.n2140 VPWR.t1541 738.074
R8242 VPWR.n619 VPWR.t1628 738.074
R8243 VPWR.n620 VPWR.t795 738.074
R8244 VPWR.n624 VPWR.t622 738.074
R8245 VPWR.n610 VPWR.t480 738.074
R8246 VPWR.n607 VPWR.t517 738.074
R8247 VPWR.n2181 VPWR.t663 738.074
R8248 VPWR.n606 VPWR.t361 738.074
R8249 VPWR.n2184 VPWR.t1576 738.074
R8250 VPWR.n2185 VPWR.t1599 738.074
R8251 VPWR.n2186 VPWR.t188 738.074
R8252 VPWR.n588 VPWR.t11 738.074
R8253 VPWR.n589 VPWR.t581 738.074
R8254 VPWR.n2090 VPWR.t1803 738.074
R8255 VPWR.n2067 VPWR.t1700 738.074
R8256 VPWR.n2087 VPWR.t735 738.074
R8257 VPWR.n2068 VPWR.t1535 738.074
R8258 VPWR.n2069 VPWR.t775 738.074
R8259 VPWR.n2070 VPWR.t1688 738.074
R8260 VPWR.n2071 VPWR.t618 738.074
R8261 VPWR.n2092 VPWR.t462 738.074
R8262 VPWR.n2093 VPWR.t651 738.074
R8263 VPWR.n2095 VPWR.t127 738.074
R8264 VPWR.n2096 VPWR.t369 738.074
R8265 VPWR.n599 VPWR.t766 738.074
R8266 VPWR.n598 VPWR.t1813 738.074
R8267 VPWR.n597 VPWR.t192 738.074
R8268 VPWR.n2223 VPWR.t19 738.074
R8269 VPWR.n596 VPWR.t585 738.074
R8270 VPWR.n714 VPWR.t1850 738.074
R8271 VPWR.n1937 VPWR.t1583 738.074
R8272 VPWR.n1940 VPWR.t817 738.074
R8273 VPWR.n762 VPWR.t1495 738.074
R8274 VPWR.n1934 VPWR.t938 738.074
R8275 VPWR.n763 VPWR.t701 738.074
R8276 VPWR.n1922 VPWR.t598 738.074
R8277 VPWR.n715 VPWR.t1840 738.074
R8278 VPWR.n721 VPWR.t809 738.074
R8279 VPWR.n720 VPWR.t669 738.074
R8280 VPWR.n724 VPWR.t1894 738.074
R8281 VPWR.n726 VPWR.t746 738.074
R8282 VPWR.n727 VPWR.t1605 738.074
R8283 VPWR.n733 VPWR.t1469 738.074
R8284 VPWR.n732 VPWR.t1706 738.074
R8285 VPWR.n736 VPWR.t1719 738.074
R8286 VPWR.n753 VPWR.t410 738.074
R8287 VPWR.n775 VPWR.t1745 738.074
R8288 VPWR.n773 VPWR.t708 738.074
R8289 VPWR.n772 VPWR.t1525 738.074
R8290 VPWR.n771 VPWR.t964 738.074
R8291 VPWR.n769 VPWR.t1565 738.074
R8292 VPWR.n766 VPWR.t614 738.074
R8293 VPWR.n752 VPWR.t468 738.074
R8294 VPWR.n751 VPWR.t113 738.074
R8295 VPWR.n750 VPWR.t567 738.074
R8296 VPWR.n747 VPWR.t268 738.074
R8297 VPWR.n1988 VPWR.t1025 738.074
R8298 VPWR.n746 VPWR.t911 738.074
R8299 VPWR.n1991 VPWR.t1055 738.074
R8300 VPWR.n1992 VPWR.t1908 738.074
R8301 VPWR.n1993 VPWR.t527 738.074
R8302 VPWR.n815 VPWR.t1848 738.074
R8303 VPWR.n809 VPWR.t925 738.074
R8304 VPWR.n808 VPWR.t815 738.074
R8305 VPWR.n806 VPWR.t1497 738.074
R8306 VPWR.n798 VPWR.t1624 738.074
R8307 VPWR.n803 VPWR.t699 738.074
R8308 VPWR.n799 VPWR.t600 738.074
R8309 VPWR.n820 VPWR.t1838 738.074
R8310 VPWR.n814 VPWR.t805 738.074
R8311 VPWR.n823 VPWR.t667 738.074
R8312 VPWR.n825 VPWR.t1892 738.074
R8313 VPWR.n826 VPWR.t221 738.074
R8314 VPWR.n828 VPWR.t1615 738.074
R8315 VPWR.n829 VPWR.t1465 738.074
R8316 VPWR.n830 VPWR.t1704 738.074
R8317 VPWR.n831 VPWR.t1717 738.074
R8318 VPWR.n445 VPWR.t712 738.074
R8319 VPWR.n2559 VPWR.t1523 738.074
R8320 VPWR.n2551 VPWR.t966 738.074
R8321 VPWR.n2556 VPWR.t1567 738.074
R8322 VPWR.n2552 VPWR.t612 738.074
R8323 VPWR.n444 VPWR.t1747 738.074
R8324 VPWR.n443 VPWR.t412 738.074
R8325 VPWR.n2590 VPWR.t470 738.074
R8326 VPWR.n442 VPWR.t1 738.074
R8327 VPWR.n2593 VPWR.t569 738.074
R8328 VPWR.n2594 VPWR.t270 738.074
R8329 VPWR.n2595 VPWR.t1027 738.074
R8330 VPWR.n2597 VPWR.t1543 738.074
R8331 VPWR.n2598 VPWR.t1057 738.074
R8332 VPWR.n2600 VPWR.t1910 738.074
R8333 VPWR.n2601 VPWR.t531 738.074
R8334 VPWR.n1791 VPWR.t429 738.074
R8335 VPWR.n1794 VPWR.t1776 738.074
R8336 VPWR.n868 VPWR.t1067 738.074
R8337 VPWR.n1788 VPWR.t1509 738.074
R8338 VPWR.n869 VPWR.t505 738.074
R8339 VPWR.n870 VPWR.t251 738.074
R8340 VPWR.n871 VPWR.t606 738.074
R8341 VPWR.n850 VPWR.t1043 738.074
R8342 VPWR.n849 VPWR.t306 738.074
R8343 VPWR.n1835 VPWR.t1015 738.074
R8344 VPWR.n845 VPWR.t1821 738.074
R8345 VPWR.n844 VPWR.t209 738.074
R8346 VPWR.n843 VPWR.t1632 738.074
R8347 VPWR.n842 VPWR.t997 738.074
R8348 VPWR.n377 VPWR.t511 738.074
R8349 VPWR.n375 VPWR.t484 738.074
R8350 VPWR.n372 VPWR.t602 738.074
R8351 VPWR.n383 VPWR.t1505 738.074
R8352 VPWR.n382 VPWR.t1073 738.074
R8353 VPWR.n386 VPWR.t1782 738.074
R8354 VPWR.n392 VPWR.t435 738.074
R8355 VPWR.n391 VPWR.t81 738.074
R8356 VPWR.n395 VPWR.t722 738.074
R8357 VPWR.n401 VPWR.t890 738.074
R8358 VPWR.n400 VPWR.t310 738.074
R8359 VPWR.n404 VPWR.t1021 738.074
R8360 VPWR.n410 VPWR.t1825 738.074
R8361 VPWR.n409 VPWR.t213 738.074
R8362 VPWR.n413 VPWR.t1636 738.074
R8363 VPWR.n2672 VPWR.t1003 738.074
R8364 VPWR.n886 VPWR.t827 738.074
R8365 VPWR.n884 VPWR.t1487 738.074
R8366 VPWR.n877 VPWR.t946 738.074
R8367 VPWR.n881 VPWR.t705 738.074
R8368 VPWR.n878 VPWR.t591 738.074
R8369 VPWR.n907 VPWR.t754 738.074
R8370 VPWR.n909 VPWR.t1609 738.074
R8371 VPWR.n910 VPWR.t1477 738.074
R8372 VPWR.n1719 VPWR.t21 738.074
R8373 VPWR.n1718 VPWR.t577 738.074
R8374 VPWR.n291 VPWR.t608 738.074
R8375 VPWR.n294 VPWR.t1694 738.074
R8376 VPWR.n296 VPWR.t257 738.074
R8377 VPWR.n298 VPWR.t1513 738.074
R8378 VPWR.n299 VPWR.t1065 738.074
R8379 VPWR.n301 VPWR.t501 738.074
R8380 VPWR.n302 VPWR.t1884 738.074
R8381 VPWR.n304 VPWR.t71 738.074
R8382 VPWR.n305 VPWR.t871 738.074
R8383 VPWR.n307 VPWR.t1039 738.074
R8384 VPWR.n308 VPWR.t304 738.074
R8385 VPWR.n310 VPWR.t1011 738.074
R8386 VPWR.n311 VPWR.t905 738.074
R8387 VPWR.n313 VPWR.t207 738.074
R8388 VPWR.n314 VPWR.t972 738.074
R8389 VPWR.n316 VPWR.t995 738.074
R8390 VPWR.n1161 VPWR.t1399 738.074
R8391 VPWR.n1160 VPWR.t1161 738.074
R8392 VPWR.n1164 VPWR.t1263 738.074
R8393 VPWR.n1277 VPWR.t1425 738.074
R8394 VPWR.n1271 VPWR.t1143 738.074
R8395 VPWR.n1270 VPWR.t1155 738.074
R8396 VPWR.n1266 VPWR.t1314 738.074
R8397 VPWR.n1265 VPWR.t1364 738.074
R8398 VPWR.n1261 VPWR.t1183 738.074
R8399 VPWR.n1260 VPWR.t1209 738.074
R8400 VPWR.n1254 VPWR.t1339 738.074
R8401 VPWR.n1253 VPWR.t1082 738.074
R8402 VPWR.n1527 VPWR.t1103 738.074
R8403 VPWR.n1524 VPWR.t1344 738.074
R8404 VPWR.n1238 VPWR.t1378 738.074
R8405 VPWR.n1239 VPWR.t1089 738.074
R8406 VPWR.n85 VPWR.t1275 738.074
R8407 VPWR.n80 VPWR.t1396 738.074
R8408 VPWR.n79 VPWR.t1152 738.074
R8409 VPWR.n74 VPWR.t1260 738.074
R8410 VPWR.n73 VPWR.t1272 738.074
R8411 VPWR.n68 VPWR.t1428 738.074
R8412 VPWR.n67 VPWR.t1149 738.074
R8413 VPWR.n62 VPWR.t1309 738.074
R8414 VPWR.n61 VPWR.t1328 738.074
R8415 VPWR.n56 VPWR.t1455 738.074
R8416 VPWR.n55 VPWR.t1199 738.074
R8417 VPWR.n50 VPWR.t1229 738.074
R8418 VPWR.n49 VPWR.t1079 738.074
R8419 VPWR.n44 VPWR.t1098 738.074
R8420 VPWR.n43 VPWR.t1223 738.074
R8421 VPWR.n86 VPWR.t1130 738.074
R8422 VPWR.n924 VPWR.t1389 646.071
R8423 VPWR.n1619 VPWR.t1613 646.071
R8424 VPWR.n1623 VPWR.t180 646.071
R8425 VPWR.n1227 VPWR.t1563 646.071
R8426 VPWR.n1223 VPWR.t1570 646.071
R8427 VPWR.n1218 VPWR.t515 646.071
R8428 VPWR.n1214 VPWR.t1836 646.071
R8429 VPWR.n1209 VPWR.t915 646.071
R8430 VPWR.n1176 VPWR.t1669 646.071
R8431 VPWR.n1718 VPWR.t1266 646.071
R8432 VPWR.n907 VPWR.t1603 646.071
R8433 VPWR.n906 VPWR.t758 646.071
R8434 VPWR.n904 VPWR.t365 646.071
R8435 VPWR.n895 VPWR.t661 646.071
R8436 VPWR.n901 VPWR.t109 646.071
R8437 VPWR.n896 VPWR.t1772 646.071
R8438 VPWR.n887 VPWR.t166 646.071
R8439 VPWR.n842 VPWR.t1420 646.071
R8440 VPWR.n850 VPWR.t1557 646.071
R8441 VPWR.n858 VPWR.t892 646.071
R8442 VPWR.n859 VPWR.t57 646.071
R8443 VPWR.n422 VPWR.t1226 646.071
R8444 VPWR.n2509 VPWR.t5 646.071
R8445 VPWR.n459 VPWR.t460 646.071
R8446 VPWR.n458 VPWR.t1801 646.071
R8447 VPWR.n456 VPWR.t1698 646.071
R8448 VPWR.n455 VPWR.t714 646.071
R8449 VPWR.n493 VPWR.t1517 646.071
R8450 VPWR.n491 VPWR.t773 646.071
R8451 VPWR.n489 VPWR.t245 646.071
R8452 VPWR.n2514 VPWR.t125 646.071
R8453 VPWR.n2508 VPWR.t371 646.071
R8454 VPWR.n2517 VPWR.t1867 646.071
R8455 VPWR.n430 VPWR.t1815 646.071
R8456 VPWR.n429 VPWR.t1061 646.071
R8457 VPWR.n423 VPWR.t25 646.071
R8458 VPWR.n2659 VPWR.t533 646.071
R8459 VPWR.n466 VPWR.t1444 646.071
R8460 VPWR.n473 VPWR.t807 646.071
R8461 VPWR.n2437 VPWR.t73 646.071
R8462 VPWR.n481 VPWR.t427 646.071
R8463 VPWR.n2434 VPWR.t1774 646.071
R8464 VPWR.n482 VPWR.t1798 646.071
R8465 VPWR.n483 VPWR.t1491 646.071
R8466 VPWR.n484 VPWR.t503 646.071
R8467 VPWR.n485 VPWR.t486 646.071
R8468 VPWR.n472 VPWR.t1041 646.071
R8469 VPWR.n471 VPWR.t312 646.071
R8470 VPWR.n2472 VPWR.t1013 646.071
R8471 VPWR.n470 VPWR.t1827 646.071
R8472 VPWR.n469 VPWR.t1467 646.071
R8473 VPWR.n468 VPWR.t1638 646.071
R8474 VPWR.n467 VPWR.t1713 646.071
R8475 VPWR.n536 VPWR.t1293 646.071
R8476 VPWR.n519 VPWR.t107 646.071
R8477 VPWR.n518 VPWR.t1770 646.071
R8478 VPWR.n516 VPWR.t164 646.071
R8479 VPWR.n515 VPWR.t1593 646.071
R8480 VPWR.n513 VPWR.t1790 646.071
R8481 VPWR.n505 VPWR.t1529 646.071
R8482 VPWR.n510 VPWR.t948 646.071
R8483 VPWR.n506 VPWR.t793 646.071
R8484 VPWR.n521 VPWR.t659 646.071
R8485 VPWR.n522 VPWR.t359 646.071
R8486 VPWR.n524 VPWR.t756 646.071
R8487 VPWR.n525 VPWR.t1597 646.071
R8488 VPWR.n531 VPWR.t1049 646.071
R8489 VPWR.n530 VPWR.t9 646.071
R8490 VPWR.n534 VPWR.t521 646.071
R8491 VPWR.n542 VPWR.t1410 646.071
R8492 VPWR.n568 VPWR.t61 646.071
R8493 VPWR.n567 VPWR.t85 646.071
R8494 VPWR.n566 VPWR.t439 646.071
R8495 VPWR.n565 VPWR.t1665 646.071
R8496 VPWR.n689 VPWR.t823 646.071
R8497 VPWR.n692 VPWR.t1483 646.071
R8498 VPWR.n687 VPWR.t450 646.071
R8499 VPWR.n684 VPWR.t492 646.071
R8500 VPWR.n555 VPWR.t894 646.071
R8501 VPWR.n2312 VPWR.t1559 646.071
R8502 VPWR.n554 VPWR.t176 646.071
R8503 VPWR.n2315 VPWR.t94 646.071
R8504 VPWR.n2317 VPWR.t1479 646.071
R8505 VPWR.n2318 VPWR.t117 646.071
R8506 VPWR.n543 VPWR.t1725 646.071
R8507 VPWR.n2255 VPWR.t1127 646.071
R8508 VPWR.n639 VPWR.t724 646.071
R8509 VPWR.n638 VPWR.t472 646.071
R8510 VPWR.n636 VPWR.t414 646.071
R8511 VPWR.n669 VPWR.t1678 646.071
R8512 VPWR.n635 VPWR.t1071 646.071
R8513 VPWR.n633 VPWR.t1503 646.071
R8514 VPWR.n631 VPWR.t1926 646.071
R8515 VPWR.n628 VPWR.t801 646.071
R8516 VPWR.n641 VPWR.t571 646.071
R8517 VPWR.n642 VPWR.t272 646.071
R8518 VPWR.n644 VPWR.t760 646.071
R8519 VPWR.n645 VPWR.t1545 646.071
R8520 VPWR.n580 VPWR.t215 646.071
R8521 VPWR.n581 VPWR.t1912 646.071
R8522 VPWR.n2254 VPWR.t1001 646.071
R8523 VPWR.n589 VPWR.t1234 646.071
R8524 VPWR.n610 VPWR.t3 646.071
R8525 VPWR.n611 VPWR.t458 646.071
R8526 VPWR.n614 VPWR.t172 646.071
R8527 VPWR.n615 VPWR.t1696 646.071
R8528 VPWR.n2140 VPWR.t710 646.071
R8529 VPWR.n619 VPWR.t1519 646.071
R8530 VPWR.n620 VPWR.t771 646.071
R8531 VPWR.n624 VPWR.t1686 646.071
R8532 VPWR.n607 VPWR.t123 646.071
R8533 VPWR.n2181 VPWR.t367 646.071
R8534 VPWR.n606 VPWR.t1580 646.071
R8535 VPWR.n2184 VPWR.t1811 646.071
R8536 VPWR.n2185 VPWR.t1059 646.071
R8537 VPWR.n2186 VPWR.t17 646.071
R8538 VPWR.n588 VPWR.t529 646.071
R8539 VPWR.n596 VPWR.t1194 646.071
R8540 VPWR.n2092 VPWR.t869 646.071
R8541 VPWR.n2090 VPWR.t464 646.071
R8542 VPWR.n2067 VPWR.t1805 646.071
R8543 VPWR.n2087 VPWR.t1702 646.071
R8544 VPWR.n2068 VPWR.t716 646.071
R8545 VPWR.n2069 VPWR.t1511 646.071
R8546 VPWR.n2070 VPWR.t777 646.071
R8547 VPWR.n2071 VPWR.t247 646.071
R8548 VPWR.n2093 VPWR.t420 646.071
R8549 VPWR.n2095 VPWR.t264 646.071
R8550 VPWR.n2096 VPWR.t768 646.071
R8551 VPWR.n599 VPWR.t907 646.071
R8552 VPWR.n598 VPWR.t205 646.071
R8553 VPWR.n597 VPWR.t27 646.071
R8554 VPWR.n2223 VPWR.t535 646.071
R8555 VPWR.n736 VPWR.t1299 646.071
R8556 VPWR.n715 VPWR.t655 646.071
R8557 VPWR.n714 VPWR.t1846 646.071
R8558 VPWR.n1937 VPWR.t1856 646.071
R8559 VPWR.n1940 VPWR.t1589 646.071
R8560 VPWR.n762 VPWR.t1788 646.071
R8561 VPWR.n1934 VPWR.t1531 646.071
R8562 VPWR.n763 VPWR.t944 646.071
R8563 VPWR.n1922 VPWR.t791 646.071
R8564 VPWR.n721 VPWR.t675 646.071
R8565 VPWR.n720 VPWR.t357 646.071
R8566 VPWR.n724 VPWR.t752 646.071
R8567 VPWR.n726 VPWR.t1595 646.071
R8568 VPWR.n727 VPWR.t1047 646.071
R8569 VPWR.n733 VPWR.t7 646.071
R8570 VPWR.n732 VPWR.t589 646.071
R8571 VPWR.n1993 VPWR.t1119 646.071
R8572 VPWR.n752 VPWR.t726 646.071
R8573 VPWR.n753 VPWR.t474 646.071
R8574 VPWR.n775 VPWR.t1878 646.071
R8575 VPWR.n773 VPWR.t1680 646.071
R8576 VPWR.n772 VPWR.t1075 646.071
R8577 VPWR.n771 VPWR.t1501 646.071
R8578 VPWR.n769 VPWR.t1928 646.071
R8579 VPWR.n766 VPWR.t803 646.071
R8580 VPWR.n751 VPWR.t573 646.071
R8581 VPWR.n750 VPWR.t274 646.071
R8582 VPWR.n747 VPWR.t762 646.071
R8583 VPWR.n1988 VPWR.t1547 646.071
R8584 VPWR.n746 VPWR.t217 646.071
R8585 VPWR.n1991 VPWR.t1817 646.071
R8586 VPWR.n1992 VPWR.t1005 646.071
R8587 VPWR.n831 VPWR.t1306 646.071
R8588 VPWR.n820 VPWR.t653 646.071
R8589 VPWR.n815 VPWR.t1844 646.071
R8590 VPWR.n809 VPWR.t1854 646.071
R8591 VPWR.n808 VPWR.t1587 646.071
R8592 VPWR.n806 VPWR.t1786 646.071
R8593 VPWR.n798 VPWR.t1533 646.071
R8594 VPWR.n803 VPWR.t942 646.071
R8595 VPWR.n799 VPWR.t789 646.071
R8596 VPWR.n814 VPWR.t673 646.071
R8597 VPWR.n823 VPWR.t355 646.071
R8598 VPWR.n825 VPWR.t750 646.071
R8599 VPWR.n826 VPWR.t1611 646.071
R8600 VPWR.n828 VPWR.t194 646.071
R8601 VPWR.n829 VPWR.t23 646.071
R8602 VPWR.n830 VPWR.t587 646.071
R8603 VPWR.n2601 VPWR.t1111 646.071
R8604 VPWR.n444 VPWR.t1880 646.071
R8605 VPWR.n445 VPWR.t1682 646.071
R8606 VPWR.n2559 VPWR.t1796 646.071
R8607 VPWR.n2551 VPWR.t1499 646.071
R8608 VPWR.n2556 VPWR.t1930 646.071
R8609 VPWR.n2552 VPWR.t1690 646.071
R8610 VPWR.n443 VPWR.t476 646.071
R8611 VPWR.n2590 VPWR.t1710 646.071
R8612 VPWR.n442 VPWR.t575 646.071
R8613 VPWR.n2593 VPWR.t276 646.071
R8614 VPWR.n2594 VPWR.t764 646.071
R8615 VPWR.n2595 VPWR.t1549 646.071
R8616 VPWR.n2597 VPWR.t219 646.071
R8617 VPWR.n2598 VPWR.t1819 646.071
R8618 VPWR.n2600 VPWR.t1007 646.071
R8619 VPWR.n1791 VPWR.t83 646.071
R8620 VPWR.n1794 VPWR.t437 646.071
R8621 VPWR.n868 VPWR.t1784 646.071
R8622 VPWR.n1788 VPWR.t819 646.071
R8623 VPWR.n869 VPWR.t1485 646.071
R8624 VPWR.n870 VPWR.t513 646.071
R8625 VPWR.n871 VPWR.t490 646.071
R8626 VPWR.n849 VPWR.t174 646.071
R8627 VPWR.n1835 VPWR.t92 646.071
R8628 VPWR.n845 VPWR.t1475 646.071
R8629 VPWR.n844 VPWR.t115 646.071
R8630 VPWR.n843 VPWR.t1721 646.071
R8631 VPWR.n2672 VPWR.t1405 646.071
R8632 VPWR.n383 VPWR.t825 646.071
R8633 VPWR.n377 VPWR.t1481 646.071
R8634 VPWR.n375 VPWR.t452 646.071
R8635 VPWR.n372 VPWR.t494 646.071
R8636 VPWR.n382 VPWR.t1667 646.071
R8637 VPWR.n386 VPWR.t913 646.071
R8638 VPWR.n392 VPWR.t1834 646.071
R8639 VPWR.n391 VPWR.t63 646.071
R8640 VPWR.n395 VPWR.t896 646.071
R8641 VPWR.n401 VPWR.t1561 646.071
R8642 VPWR.n400 VPWR.t178 646.071
R8643 VPWR.n404 VPWR.t96 646.071
R8644 VPWR.n410 VPWR.t184 646.071
R8645 VPWR.n409 VPWR.t119 646.071
R8646 VPWR.n413 VPWR.t1727 646.071
R8647 VPWR.n886 VPWR.t158 646.071
R8648 VPWR.n884 VPWR.t1792 646.071
R8649 VPWR.n877 VPWR.t1521 646.071
R8650 VPWR.n881 VPWR.t1626 646.071
R8651 VPWR.n878 VPWR.t1684 646.071
R8652 VPWR.n909 VPWR.t1051 646.071
R8653 VPWR.n910 VPWR.t15 646.071
R8654 VPWR.n1719 VPWR.t523 646.071
R8655 VPWR.n1203 VPWR.t729 646.071
R8656 VPWR.n1180 VPWR.t1537 646.071
R8657 VPWR.n1184 VPWR.t454 646.071
R8658 VPWR.n1188 VPWR.t845 646.071
R8659 VPWR.n1629 VPWR.t186 646.071
R8660 VPWR.n928 VPWR.t1551 646.071
R8661 VPWR.n1709 VPWR.t579 646.071
R8662 VPWR.n316 VPWR.t1436 646.071
R8663 VPWR.n294 VPWR.t507 646.071
R8664 VPWR.n291 VPWR.t488 646.071
R8665 VPWR.n296 VPWR.t1489 646.071
R8666 VPWR.n298 VPWR.t813 646.071
R8667 VPWR.n299 VPWR.t1778 646.071
R8668 VPWR.n301 VPWR.t431 646.071
R8669 VPWR.n302 VPWR.t77 646.071
R8670 VPWR.n304 VPWR.t811 646.071
R8671 VPWR.n305 VPWR.t1045 646.071
R8672 VPWR.n307 VPWR.t1555 646.071
R8673 VPWR.n308 VPWR.t1017 646.071
R8674 VPWR.n310 VPWR.t1829 646.071
R8675 VPWR.n311 VPWR.t1471 646.071
R8676 VPWR.n313 VPWR.t1640 646.071
R8677 VPWR.n314 VPWR.t1715 646.071
R8678 VPWR.n1239 VPWR.t1212 646.071
R8679 VPWR.n1161 VPWR.t1108 646.071
R8680 VPWR.n1160 VPWR.t1244 646.071
R8681 VPWR.n1164 VPWR.t1257 646.071
R8682 VPWR.n1277 VPWR.t1361 646.071
R8683 VPWR.n1271 VPWR.t1138 646.071
R8684 VPWR.n1270 VPWR.t1285 646.071
R8685 VPWR.n1266 VPWR.t1402 646.071
R8686 VPWR.n1265 VPWR.t1433 646.071
R8687 VPWR.n1261 VPWR.t1178 646.071
R8688 VPWR.n1260 VPWR.t1282 646.071
R8689 VPWR.n1254 VPWR.t1441 646.071
R8690 VPWR.n1253 VPWR.t1460 646.071
R8691 VPWR.n1527 VPWR.t1204 646.071
R8692 VPWR.n1524 VPWR.t1336 646.071
R8693 VPWR.n1238 VPWR.t1370 646.071
R8694 VPWR.n86 VPWR.t1237 646.071
R8695 VPWR.n85 VPWR.t1375 646.071
R8696 VPWR.n80 VPWR.t1381 646.071
R8697 VPWR.n79 VPWR.t1146 646.071
R8698 VPWR.n74 VPWR.t1254 646.071
R8699 VPWR.n73 VPWR.t1415 646.071
R8700 VPWR.n68 VPWR.t1133 646.071
R8701 VPWR.n67 VPWR.t1168 646.071
R8702 VPWR.n62 VPWR.t1296 646.071
R8703 VPWR.n61 VPWR.t1367 646.071
R8704 VPWR.n56 VPWR.t1173 646.071
R8705 VPWR.n55 VPWR.t1191 646.071
R8706 VPWR.n50 VPWR.t1319 646.071
R8707 VPWR.n49 VPWR.t1452 646.071
R8708 VPWR.n44 VPWR.t1092 646.071
R8709 VPWR.n43 VPWR.t1331 646.071
R8710 VPWR.n1618 VPWR.t1247 642.13
R8711 VPWR.n1622 VPWR.t1114 642.13
R8712 VPWR.n1226 VPWR.t1386 642.13
R8713 VPWR.n1222 VPWR.t1358 642.13
R8714 VPWR.n1217 VPWR.t1217 642.13
R8715 VPWR.n1213 VPWR.t1095 642.13
R8716 VPWR.n1208 VPWR.t1347 642.13
R8717 VPWR.n1175 VPWR.t1325 642.13
R8718 VPWR.n1202 VPWR.t1220 642.13
R8719 VPWR.n1179 VPWR.t1449 642.13
R8720 VPWR.n1183 VPWR.t1322 642.13
R8721 VPWR.n1187 VPWR.t1186 642.13
R8722 VPWR.n1628 VPWR.t1288 642.13
R8723 VPWR.n927 VPWR.t1124 642.13
R8724 VPWR.n1708 VPWR.t1158 642.13
R8725 VPWR.n923 VPWR.t1269 642.13
R8726 VPWR.n492 VPWR.t244 629.652
R8727 VPWR.n496 VPWR.t772 629.652
R8728 VPWR.t1516 VPWR.n495 629.652
R8729 VPWR.n2541 VPWR.t713 629.652
R8730 VPWR.t1697 VPWR.n2540 629.652
R8731 VPWR.n2534 VPWR.t1800 629.652
R8732 VPWR.t459 VPWR.n2533 629.652
R8733 VPWR.n2513 VPWR.t4 629.652
R8734 VPWR.n2516 VPWR.t124 629.652
R8735 VPWR.n2521 VPWR.t370 629.652
R8736 VPWR.t1866 VPWR.n2520 629.652
R8737 VPWR.n2646 VPWR.t1814 629.652
R8738 VPWR.n2647 VPWR.t1060 629.652
R8739 VPWR.n2658 VPWR.t24 629.652
R8740 VPWR.n2661 VPWR.t532 629.652
R8741 VPWR.n486 VPWR.t485 629.652
R8742 VPWR.n2426 VPWR.t502 629.652
R8743 VPWR.n2427 VPWR.t1490 629.652
R8744 VPWR.n2433 VPWR.t1797 629.652
R8745 VPWR.n2436 VPWR.t1773 629.652
R8746 VPWR.n2442 VPWR.t426 629.652
R8747 VPWR.t72 VPWR.n2441 629.652
R8748 VPWR.n2464 VPWR.t806 629.652
R8749 VPWR.n2465 VPWR.t1040 629.652
R8750 VPWR.n2471 VPWR.t311 629.652
R8751 VPWR.n2476 VPWR.t1012 629.652
R8752 VPWR.n2477 VPWR.t1826 629.652
R8753 VPWR.n2484 VPWR.t1466 629.652
R8754 VPWR.n2485 VPWR.t1637 629.652
R8755 VPWR.n2492 VPWR.t1712 629.652
R8756 VPWR.n509 VPWR.t792 629.652
R8757 VPWR.n512 VPWR.t947 629.652
R8758 VPWR.n2407 VPWR.t1528 629.652
R8759 VPWR.t1789 VPWR.n2406 629.652
R8760 VPWR.n2400 VPWR.t1592 629.652
R8761 VPWR.t163 VPWR.n2399 629.652
R8762 VPWR.n2393 VPWR.t1769 629.652
R8763 VPWR.t106 VPWR.n2392 629.652
R8764 VPWR.n2386 VPWR.t658 629.652
R8765 VPWR.t358 VPWR.n2385 629.652
R8766 VPWR.n2379 VPWR.t755 629.652
R8767 VPWR.t1596 VPWR.n2378 629.652
R8768 VPWR.n533 VPWR.t1048 629.652
R8769 VPWR.n2367 VPWR.t8 629.652
R8770 VPWR.t520 VPWR.n2366 629.652
R8771 VPWR.n688 VPWR.t491 629.652
R8772 VPWR.n696 VPWR.t449 629.652
R8773 VPWR.t1482 VPWR.n695 629.652
R8774 VPWR.t822 VPWR.n691 629.652
R8775 VPWR.n2288 VPWR.t1664 629.652
R8776 VPWR.t438 VPWR.n2287 629.652
R8777 VPWR.n571 VPWR.t84 629.652
R8778 VPWR.t60 VPWR.n570 629.652
R8779 VPWR.n2311 VPWR.t893 629.652
R8780 VPWR.n2314 VPWR.t1558 629.652
R8781 VPWR.n2328 VPWR.t175 629.652
R8782 VPWR.t93 VPWR.n2327 629.652
R8783 VPWR.n2321 VPWR.t1478 629.652
R8784 VPWR.t116 VPWR.n2320 629.652
R8785 VPWR.n2352 VPWR.t1724 629.652
R8786 VPWR.n632 VPWR.t800 629.652
R8787 VPWR.n680 VPWR.t1925 629.652
R8788 VPWR.t1502 VPWR.n679 629.652
R8789 VPWR.n673 VPWR.t1070 629.652
R8790 VPWR.t1677 VPWR.n672 629.652
R8791 VPWR.t413 VPWR.n668 629.652
R8792 VPWR.n662 VPWR.t471 629.652
R8793 VPWR.t723 VPWR.n661 629.652
R8794 VPWR.n655 VPWR.t570 629.652
R8795 VPWR.t271 VPWR.n654 629.652
R8796 VPWR.n648 VPWR.t759 629.652
R8797 VPWR.t1544 VPWR.n647 629.652
R8798 VPWR.n2266 VPWR.t214 629.652
R8799 VPWR.t1911 VPWR.n2265 629.652
R8800 VPWR.n2259 VPWR.t1000 629.652
R8801 VPWR.n625 VPWR.t1685 629.652
R8802 VPWR.n2139 VPWR.t770 629.652
R8803 VPWR.n2143 VPWR.t1518 629.652
R8804 VPWR.t709 VPWR.n2142 629.652
R8805 VPWR.n2156 VPWR.t1695 629.652
R8806 VPWR.n2157 VPWR.t171 629.652
R8807 VPWR.n2168 VPWR.t457 629.652
R8808 VPWR.n2169 VPWR.t2 629.652
R8809 VPWR.n2180 VPWR.t122 629.652
R8810 VPWR.n2183 VPWR.t366 629.652
R8811 VPWR.n2196 VPWR.t1579 629.652
R8812 VPWR.t1810 VPWR.n2195 629.652
R8813 VPWR.n2189 VPWR.t1058 629.652
R8814 VPWR.t16 VPWR.n2188 629.652
R8815 VPWR.n2239 VPWR.t528 629.652
R8816 VPWR.n2072 VPWR.t246 629.652
R8817 VPWR.n2078 VPWR.t776 629.652
R8818 VPWR.n2079 VPWR.t1510 629.652
R8819 VPWR.n2086 VPWR.t715 629.652
R8820 VPWR.n2089 VPWR.t1701 629.652
R8821 VPWR.n2114 VPWR.t1804 629.652
R8822 VPWR.t463 VPWR.n2113 629.652
R8823 VPWR.n2107 VPWR.t868 629.652
R8824 VPWR.t419 VPWR.n2106 629.652
R8825 VPWR.n2100 VPWR.t263 629.652
R8826 VPWR.t767 VPWR.n2099 629.652
R8827 VPWR.n2214 VPWR.t906 629.652
R8828 VPWR.n2215 VPWR.t204 629.652
R8829 VPWR.n2222 VPWR.t26 629.652
R8830 VPWR.n2225 VPWR.t534 629.652
R8831 VPWR.n1923 VPWR.t790 629.652
R8832 VPWR.n1933 VPWR.t943 629.652
R8833 VPWR.n1936 VPWR.t1530 629.652
R8834 VPWR.n1944 VPWR.t1787 629.652
R8835 VPWR.t1588 VPWR.n1943 629.652
R8836 VPWR.t1855 VPWR.n1939 629.652
R8837 VPWR.n2057 VPWR.t1845 629.652
R8838 VPWR.t654 VPWR.n2056 629.652
R8839 VPWR.n723 VPWR.t674 629.652
R8840 VPWR.n2045 VPWR.t356 629.652
R8841 VPWR.t751 VPWR.n2044 629.652
R8842 VPWR.n2038 VPWR.t1594 629.652
R8843 VPWR.t1046 VPWR.n2037 629.652
R8844 VPWR.n735 VPWR.t6 629.652
R8845 VPWR.n2026 VPWR.t588 629.652
R8846 VPWR.n770 VPWR.t802 629.652
R8847 VPWR.n790 VPWR.t1927 629.652
R8848 VPWR.t1500 VPWR.n789 629.652
R8849 VPWR.n783 VPWR.t1074 629.652
R8850 VPWR.t1679 VPWR.n782 629.652
R8851 VPWR.n776 VPWR.t1877 629.652
R8852 VPWR.n1963 VPWR.t473 629.652
R8853 VPWR.n1964 VPWR.t725 629.652
R8854 VPWR.n1971 VPWR.t572 629.652
R8855 VPWR.n1972 VPWR.t273 629.652
R8856 VPWR.n1987 VPWR.t761 629.652
R8857 VPWR.n1990 VPWR.t1546 629.652
R8858 VPWR.n2003 VPWR.t216 629.652
R8859 VPWR.t1816 VPWR.n2002 629.652
R8860 VPWR.n1996 VPWR.t1004 629.652
R8861 VPWR.n802 VPWR.t788 629.652
R8862 VPWR.n805 VPWR.t941 629.652
R8863 VPWR.n1909 VPWR.t1532 629.652
R8864 VPWR.t1785 VPWR.n1908 629.652
R8865 VPWR.n1902 VPWR.t1586 629.652
R8866 VPWR.t1853 VPWR.n1901 629.652
R8867 VPWR.n819 VPWR.t1843 629.652
R8868 VPWR.n822 VPWR.t652 629.652
R8869 VPWR.n1889 VPWR.t672 629.652
R8870 VPWR.t354 VPWR.n1888 629.652
R8871 VPWR.n1882 VPWR.t749 629.652
R8872 VPWR.t1610 VPWR.n1881 629.652
R8873 VPWR.n1875 VPWR.t193 629.652
R8874 VPWR.t22 VPWR.n1874 629.652
R8875 VPWR.n835 VPWR.t586 629.652
R8876 VPWR.n2555 VPWR.t1689 629.652
R8877 VPWR.n2558 VPWR.t1929 629.652
R8878 VPWR.n2564 VPWR.t1498 629.652
R8879 VPWR.t1795 VPWR.n2563 629.652
R8880 VPWR.n2581 VPWR.t1681 629.652
R8881 VPWR.n2582 VPWR.t1879 629.652
R8882 VPWR.n2589 VPWR.t475 629.652
R8883 VPWR.n2592 VPWR.t1709 629.652
R8884 VPWR.n2625 VPWR.t574 629.652
R8885 VPWR.t275 VPWR.n2624 629.652
R8886 VPWR.n2618 VPWR.t763 629.652
R8887 VPWR.t1548 VPWR.n2617 629.652
R8888 VPWR.n2611 VPWR.t218 629.652
R8889 VPWR.t1818 VPWR.n2610 629.652
R8890 VPWR.n2604 VPWR.t1006 629.652
R8891 VPWR.n1780 VPWR.t489 629.652
R8892 VPWR.n1781 VPWR.t512 629.652
R8893 VPWR.n1787 VPWR.t1484 629.652
R8894 VPWR.n1790 VPWR.t818 629.652
R8895 VPWR.n1799 VPWR.t1783 629.652
R8896 VPWR.t436 VPWR.n1798 629.652
R8897 VPWR.t82 VPWR.n1793 629.652
R8898 VPWR.n1822 VPWR.t56 629.652
R8899 VPWR.n1823 VPWR.t891 629.652
R8900 VPWR.n1834 VPWR.t1556 629.652
R8901 VPWR.n1838 VPWR.t173 629.652
R8902 VPWR.t91 VPWR.n1837 629.652
R8903 VPWR.n1849 VPWR.t1474 629.652
R8904 VPWR.n1850 VPWR.t114 629.652
R8905 VPWR.n1857 VPWR.t1720 629.652
R8906 VPWR.n376 VPWR.t493 629.652
R8907 VPWR.n2732 VPWR.t451 629.652
R8908 VPWR.t1480 VPWR.n2731 629.652
R8909 VPWR.n385 VPWR.t824 629.652
R8910 VPWR.n2720 VPWR.t1666 629.652
R8911 VPWR.t912 VPWR.n2719 629.652
R8912 VPWR.n394 VPWR.t1833 629.652
R8913 VPWR.n2708 VPWR.t62 629.652
R8914 VPWR.t895 VPWR.n2707 629.652
R8915 VPWR.n403 VPWR.t1560 629.652
R8916 VPWR.n2696 VPWR.t177 629.652
R8917 VPWR.t95 VPWR.n2695 629.652
R8918 VPWR.n412 VPWR.t183 629.652
R8919 VPWR.n2684 VPWR.t118 629.652
R8920 VPWR.t1726 VPWR.n2683 629.652
R8921 VPWR.n880 VPWR.t1683 629.652
R8922 VPWR.n883 VPWR.t1625 629.652
R8923 VPWR.n1767 VPWR.t1520 629.652
R8924 VPWR.t1791 VPWR.n1766 629.652
R8925 VPWR.n1760 VPWR.t157 629.652
R8926 VPWR.t165 VPWR.n1759 629.652
R8927 VPWR.n900 VPWR.t1771 629.652
R8928 VPWR.n903 VPWR.t108 629.652
R8929 VPWR.n1747 VPWR.t660 629.652
R8930 VPWR.t364 VPWR.n1746 629.652
R8931 VPWR.n1740 VPWR.t757 629.652
R8932 VPWR.t1602 VPWR.n1739 629.652
R8933 VPWR.n1733 VPWR.t1050 629.652
R8934 VPWR.t14 VPWR.n1732 629.652
R8935 VPWR.n1721 VPWR.t522 629.652
R8936 VPWR.n1191 VPWR.t844 629.652
R8937 VPWR.n1192 VPWR.t453 629.652
R8938 VPWR.n1199 VPWR.t1536 629.652
R8939 VPWR.n1205 VPWR.t728 629.652
R8940 VPWR.n1659 VPWR.t1668 629.652
R8941 VPWR.t914 VPWR.n1658 629.652
R8942 VPWR.n1652 VPWR.t1835 629.652
R8943 VPWR.t514 VPWR.n1651 629.652
R8944 VPWR.n1645 VPWR.t1569 629.652
R8945 VPWR.t1562 VPWR.n1644 629.652
R8946 VPWR.n1625 VPWR.t179 629.652
R8947 VPWR.n1632 VPWR.t1612 629.652
R8948 VPWR.t185 VPWR.n1631 629.652
R8949 VPWR.n1705 VPWR.t1550 629.652
R8950 VPWR.n1711 VPWR.t578 629.652
R8951 VPWR.n295 VPWR.t487 629.652
R8952 VPWR.n365 VPWR.t506 629.652
R8953 VPWR.t1488 VPWR.n364 629.652
R8954 VPWR.n358 VPWR.t812 629.652
R8955 VPWR.t1777 VPWR.n357 629.652
R8956 VPWR.n351 VPWR.t430 629.652
R8957 VPWR.t76 VPWR.n350 629.652
R8958 VPWR.n344 VPWR.t810 629.652
R8959 VPWR.t1044 VPWR.n343 629.652
R8960 VPWR.n337 VPWR.t1554 629.652
R8961 VPWR.t1016 VPWR.n336 629.652
R8962 VPWR.n330 VPWR.t1828 629.652
R8963 VPWR.t1470 VPWR.n329 629.652
R8964 VPWR.n323 VPWR.t1639 629.652
R8965 VPWR.t1714 VPWR.n322 629.652
R8966 VPWR.n1163 VPWR.t1107 629.652
R8967 VPWR.n1672 VPWR.t1243 629.652
R8968 VPWR.t1256 VPWR.n1671 629.652
R8969 VPWR.n1278 VPWR.t1360 629.652
R8970 VPWR.n1488 VPWR.t1137 629.652
R8971 VPWR.n1489 VPWR.t1284 629.652
R8972 VPWR.n1500 VPWR.t1401 629.652
R8973 VPWR.n1501 VPWR.t1432 629.652
R8974 VPWR.n1514 VPWR.t1177 629.652
R8975 VPWR.n1515 VPWR.t1281 629.652
R8976 VPWR.n1523 VPWR.t1440 629.652
R8977 VPWR.n1532 VPWR.t1459 629.652
R8978 VPWR.t1203 VPWR.n1531 629.652
R8979 VPWR.t1335 VPWR.n1526 629.652
R8980 VPWR.n1588 VPWR.t1369 629.652
R8981 VPWR.n2762 VPWR.t1236 629.652
R8982 VPWR.n2763 VPWR.t1374 629.652
R8983 VPWR.n2774 VPWR.t1380 629.652
R8984 VPWR.n2775 VPWR.t1145 629.652
R8985 VPWR.n2786 VPWR.t1253 629.652
R8986 VPWR.n2787 VPWR.t1414 629.652
R8987 VPWR.n2798 VPWR.t1132 629.652
R8988 VPWR.n2799 VPWR.t1167 629.652
R8989 VPWR.n2810 VPWR.t1295 629.652
R8990 VPWR.n2811 VPWR.t1366 629.652
R8991 VPWR.n2822 VPWR.t1172 629.652
R8992 VPWR.n2823 VPWR.t1190 629.652
R8993 VPWR.n2834 VPWR.t1318 629.652
R8994 VPWR.n2835 VPWR.t1451 629.652
R8995 VPWR.n2846 VPWR.t1091 629.652
R8996 VPWR.t244 VPWR.t926 486.048
R8997 VPWR.t772 VPWR.t104 486.048
R8998 VPWR.t861 VPWR.t1516 486.048
R8999 VPWR.t929 VPWR.t713 486.048
R9000 VPWR.t1766 VPWR.t1697 486.048
R9001 VPWR.t1800 VPWR.t102 486.048
R9002 VPWR.t865 VPWR.t459 486.048
R9003 VPWR.t4 VPWR.t1765 486.048
R9004 VPWR.t124 VPWR.t425 486.048
R9005 VPWR.t370 VPWR.t103 486.048
R9006 VPWR.t928 VPWR.t1866 486.048
R9007 VPWR.t927 VPWR.t1814 486.048
R9008 VPWR.t1060 VPWR.t864 486.048
R9009 VPWR.t863 VPWR.t24 486.048
R9010 VPWR.t532 VPWR.t862 486.048
R9011 VPWR.t1225 VPWR.t424 486.048
R9012 VPWR.t485 VPWR.t885 486.048
R9013 VPWR.t154 VPWR.t502 486.048
R9014 VPWR.t1490 VPWR.t848 486.048
R9015 VPWR.t847 VPWR.t1797 486.048
R9016 VPWR.t1773 VPWR.t884 486.048
R9017 VPWR.t426 VPWR.t323 486.048
R9018 VPWR.t322 VPWR.t72 486.048
R9019 VPWR.t883 VPWR.t806 486.048
R9020 VPWR.t1040 VPWR.t156 486.048
R9021 VPWR.t324 VPWR.t311 486.048
R9022 VPWR.t1012 VPWR.t846 486.048
R9023 VPWR.t1826 VPWR.t886 486.048
R9024 VPWR.t321 VPWR.t1466 486.048
R9025 VPWR.t1637 VPWR.t320 486.048
R9026 VPWR.t849 VPWR.t1712 486.048
R9027 VPWR.t1443 VPWR.t155 486.048
R9028 VPWR.t792 VPWR.t1657 486.048
R9029 VPWR.t947 VPWR.t1652 486.048
R9030 VPWR.t1528 VPWR.t328 486.048
R9031 VPWR.t327 VPWR.t1789 486.048
R9032 VPWR.t1592 VPWR.t1656 486.048
R9033 VPWR.t1650 VPWR.t163 486.048
R9034 VPWR.t1769 VPWR.t1649 486.048
R9035 VPWR.t1655 VPWR.t106 486.048
R9036 VPWR.t658 VPWR.t1654 486.048
R9037 VPWR.t1651 VPWR.t358 486.048
R9038 VPWR.t755 VPWR.t326 486.048
R9039 VPWR.t325 VPWR.t1596 486.048
R9040 VPWR.t1048 VPWR.t331 486.048
R9041 VPWR.t8 VPWR.t330 486.048
R9042 VPWR.t329 VPWR.t520 486.048
R9043 VPWR.t1292 VPWR.t1653 486.048
R9044 VPWR.t491 VPWR.t318 486.048
R9045 VPWR.t449 VPWR.t313 486.048
R9046 VPWR.t399 VPWR.t1482 486.048
R9047 VPWR.t398 VPWR.t822 486.048
R9048 VPWR.t317 VPWR.t1664 486.048
R9049 VPWR.t299 VPWR.t438 486.048
R9050 VPWR.t84 VPWR.t298 486.048
R9051 VPWR.t316 VPWR.t60 486.048
R9052 VPWR.t315 VPWR.t893 486.048
R9053 VPWR.t1558 VPWR.t300 486.048
R9054 VPWR.t175 VPWR.t397 486.048
R9055 VPWR.t319 VPWR.t93 486.048
R9056 VPWR.t1478 VPWR.t297 486.048
R9057 VPWR.t296 VPWR.t116 486.048
R9058 VPWR.t295 VPWR.t1724 486.048
R9059 VPWR.t1409 VPWR.t314 486.048
R9060 VPWR.t800 VPWR.t850 486.048
R9061 VPWR.t1925 VPWR.t105 486.048
R9062 VPWR.t496 VPWR.t1502 486.048
R9063 VPWR.t1070 VPWR.t495 486.048
R9064 VPWR.t565 VPWR.t1677 486.048
R9065 VPWR.t294 VPWR.t413 486.048
R9066 VPWR.t471 VPWR.t293 486.048
R9067 VPWR.t564 VPWR.t723 486.048
R9068 VPWR.t570 VPWR.t563 486.048
R9069 VPWR.t1581 VPWR.t271 486.048
R9070 VPWR.t759 VPWR.t852 486.048
R9071 VPWR.t851 VPWR.t1544 486.048
R9072 VPWR.t292 VPWR.t214 486.048
R9073 VPWR.t291 VPWR.t1911 486.048
R9074 VPWR.t1000 VPWR.t497 486.048
R9075 VPWR.t562 VPWR.t1126 486.048
R9076 VPWR.t1685 VPWR.t881 486.048
R9077 VPWR.t1646 VPWR.t770 486.048
R9078 VPWR.t1518 VPWR.t536 486.048
R9079 VPWR.t743 VPWR.t709 486.048
R9080 VPWR.t880 VPWR.t1695 486.048
R9081 VPWR.t171 VPWR.t32 486.048
R9082 VPWR.t31 VPWR.t457 486.048
R9083 VPWR.t2 VPWR.t879 486.048
R9084 VPWR.t1648 VPWR.t122 486.048
R9085 VPWR.t366 VPWR.t33 486.048
R9086 VPWR.t1579 VPWR.t742 486.048
R9087 VPWR.t741 VPWR.t1810 486.048
R9088 VPWR.t1058 VPWR.t30 486.048
R9089 VPWR.t538 VPWR.t16 486.048
R9090 VPWR.t537 VPWR.t528 486.048
R9091 VPWR.t1647 VPWR.t1233 486.048
R9092 VPWR.t246 VPWR.t901 486.048
R9093 VPWR.t1037 VPWR.t776 486.048
R9094 VPWR.t1510 VPWR.t1661 486.048
R9095 VPWR.t1660 VPWR.t715 486.048
R9096 VPWR.t1701 VPWR.t900 486.048
R9097 VPWR.t1804 VPWR.t1035 486.048
R9098 VPWR.t1034 VPWR.t463 486.048
R9099 VPWR.t868 VPWR.t899 486.048
R9100 VPWR.t898 VPWR.t419 486.048
R9101 VPWR.t263 VPWR.t1036 486.048
R9102 VPWR.t1659 VPWR.t767 486.048
R9103 VPWR.t1658 VPWR.t906 486.048
R9104 VPWR.t204 VPWR.t1033 486.048
R9105 VPWR.t1663 VPWR.t26 486.048
R9106 VPWR.t534 VPWR.t1662 486.048
R9107 VPWR.t1193 VPWR.t897 486.048
R9108 VPWR.t790 VPWR.t1622 486.048
R9109 VPWR.t1617 VPWR.t943 486.048
R9110 VPWR.t1530 VPWR.t443 486.048
R9111 VPWR.t1787 VPWR.t442 486.048
R9112 VPWR.t1621 VPWR.t1588 486.048
R9113 VPWR.t448 VPWR.t1855 486.048
R9114 VPWR.t447 VPWR.t1845 486.048
R9115 VPWR.t1620 VPWR.t654 486.048
R9116 VPWR.t674 VPWR.t1619 486.048
R9117 VPWR.t356 VPWR.t1616 486.048
R9118 VPWR.t441 VPWR.t751 486.048
R9119 VPWR.t1594 VPWR.t440 486.048
R9120 VPWR.t446 VPWR.t1046 486.048
R9121 VPWR.t6 VPWR.t445 486.048
R9122 VPWR.t588 VPWR.t444 486.048
R9123 VPWR.t1618 VPWR.t1298 486.048
R9124 VPWR.t802 VPWR.t876 486.048
R9125 VPWR.t1927 VPWR.t1809 486.048
R9126 VPWR.t685 VPWR.t1500 486.048
R9127 VPWR.t1074 VPWR.t684 486.048
R9128 VPWR.t875 VPWR.t1679 486.048
R9129 VPWR.t1877 VPWR.t690 486.048
R9130 VPWR.t689 VPWR.t473 486.048
R9131 VPWR.t725 VPWR.t874 486.048
R9132 VPWR.t873 VPWR.t572 486.048
R9133 VPWR.t273 VPWR.t691 486.048
R9134 VPWR.t878 VPWR.t761 486.048
R9135 VPWR.t1546 VPWR.t877 486.048
R9136 VPWR.t216 VPWR.t688 486.048
R9137 VPWR.t687 VPWR.t1816 486.048
R9138 VPWR.t1004 VPWR.t686 486.048
R9139 VPWR.t872 VPWR.t1118 486.048
R9140 VPWR.t788 VPWR.t1808 486.048
R9141 VPWR.t941 VPWR.t1915 486.048
R9142 VPWR.t1532 VPWR.t197 486.048
R9143 VPWR.t196 VPWR.t1785 486.048
R9144 VPWR.t1586 VPWR.t1807 486.048
R9145 VPWR.t1913 VPWR.t1853 486.048
R9146 VPWR.t1843 VPWR.t201 486.048
R9147 VPWR.t652 VPWR.t1806 486.048
R9148 VPWR.t672 VPWR.t1917 486.048
R9149 VPWR.t1914 VPWR.t354 486.048
R9150 VPWR.t749 VPWR.t195 486.048
R9151 VPWR.t1922 VPWR.t1610 486.048
R9152 VPWR.t193 VPWR.t200 486.048
R9153 VPWR.t199 VPWR.t22 486.048
R9154 VPWR.t586 VPWR.t198 486.048
R9155 VPWR.t1916 VPWR.t1305 486.048
R9156 VPWR.t1689 VPWR.t1645 486.048
R9157 VPWR.t1929 VPWR.t1670 486.048
R9158 VPWR.t1498 VPWR.t976 486.048
R9159 VPWR.t975 VPWR.t1795 486.048
R9160 VPWR.t1644 VPWR.t1681 486.048
R9161 VPWR.t1879 VPWR.t1675 486.048
R9162 VPWR.t1674 VPWR.t475 486.048
R9163 VPWR.t1709 VPWR.t1643 486.048
R9164 VPWR.t574 VPWR.t1642 486.048
R9165 VPWR.t1676 VPWR.t275 486.048
R9166 VPWR.t763 VPWR.t974 486.048
R9167 VPWR.t973 VPWR.t1548 486.048
R9168 VPWR.t218 VPWR.t1673 486.048
R9169 VPWR.t1672 VPWR.t1818 486.048
R9170 VPWR.t1006 VPWR.t1671 486.048
R9171 VPWR.t1641 VPWR.t1110 486.048
R9172 VPWR.t489 VPWR.t101 486.048
R9173 VPWR.t512 VPWR.t1904 486.048
R9174 VPWR.t131 VPWR.t1484 486.048
R9175 VPWR.t818 VPWR.t130 486.048
R9176 VPWR.t1783 VPWR.t100 486.048
R9177 VPWR.t1902 VPWR.t436 486.048
R9178 VPWR.t1901 VPWR.t82 486.048
R9179 VPWR.t99 VPWR.t56 486.048
R9180 VPWR.t891 VPWR.t98 486.048
R9181 VPWR.t1903 VPWR.t1556 486.048
R9182 VPWR.t173 VPWR.t129 486.048
R9183 VPWR.t128 VPWR.t91 486.048
R9184 VPWR.t1900 VPWR.t1474 486.048
R9185 VPWR.t114 VPWR.t1899 486.048
R9186 VPWR.t835 VPWR.t1720 486.048
R9187 VPWR.t1419 VPWR.t97 486.048
R9188 VPWR.t493 VPWR.t935 486.048
R9189 VPWR.t451 VPWR.t1762 486.048
R9190 VPWR.t1748 VPWR.t1480 486.048
R9191 VPWR.t824 VPWR.t1757 486.048
R9192 VPWR.t1666 VPWR.t934 486.048
R9193 VPWR.t1740 VPWR.t912 486.048
R9194 VPWR.t1833 VPWR.t1739 486.048
R9195 VPWR.t62 VPWR.t933 486.048
R9196 VPWR.t1764 VPWR.t895 486.048
R9197 VPWR.t1560 VPWR.t1741 486.048
R9198 VPWR.t177 VPWR.t1756 486.048
R9199 VPWR.t936 VPWR.t95 486.048
R9200 VPWR.t183 VPWR.t1738 486.048
R9201 VPWR.t118 VPWR.t1737 486.048
R9202 VPWR.t1736 VPWR.t1726 486.048
R9203 VPWR.t1404 VPWR.t1763 486.048
R9204 VPWR.t1683 VPWR.t1859 486.048
R9205 VPWR.t1625 VPWR.t90 486.048
R9206 VPWR.t1520 VPWR.t1863 486.048
R9207 VPWR.t1862 VPWR.t1791 486.048
R9208 VPWR.t157 VPWR.t744 486.048
R9209 VPWR.t88 VPWR.t165 486.048
R9210 VPWR.t1771 VPWR.t87 486.048
R9211 VPWR.t108 VPWR.t279 486.048
R9212 VPWR.t660 VPWR.t278 486.048
R9213 VPWR.t89 VPWR.t364 486.048
R9214 VPWR.t757 VPWR.t1861 486.048
R9215 VPWR.t1860 VPWR.t1602 486.048
R9216 VPWR.t1050 VPWR.t86 486.048
R9217 VPWR.t1865 VPWR.t14 486.048
R9218 VPWR.t522 VPWR.t1864 486.048
R9219 VPWR.t1265 VPWR.t277 486.048
R9220 VPWR.t844 VPWR.t1170 486.048
R9221 VPWR.t453 VPWR.t1301 486.048
R9222 VPWR.t1430 VPWR.t1536 486.048
R9223 VPWR.t728 VPWR.t1086 486.048
R9224 VPWR.t1668 VPWR.t1196 486.048
R9225 VPWR.t1351 VPWR.t914 486.048
R9226 VPWR.t1835 VPWR.t1353 486.048
R9227 VPWR.t1201 VPWR.t514 486.048
R9228 VPWR.t1569 VPWR.t1231 486.048
R9229 VPWR.t1349 VPWR.t1562 486.048
R9230 VPWR.t179 VPWR.t1100 486.048
R9231 VPWR.t1612 VPWR.t1116 486.048
R9232 VPWR.t1372 VPWR.t185 486.048
R9233 VPWR.t1393 VPWR.t1550 486.048
R9234 VPWR.t578 VPWR.t1422 486.048
R9235 VPWR.t1388 VPWR.t1251 486.048
R9236 VPWR.t487 VPWR.t736 486.048
R9237 VPWR.t506 VPWR.t624 486.048
R9238 VPWR.t740 VPWR.t1488 486.048
R9239 VPWR.t812 VPWR.t739 486.048
R9240 VPWR.t628 VPWR.t1777 486.048
R9241 VPWR.t430 VPWR.t1921 486.048
R9242 VPWR.t1920 VPWR.t76 486.048
R9243 VPWR.t810 VPWR.t627 486.048
R9244 VPWR.t626 VPWR.t1044 486.048
R9245 VPWR.t1554 VPWR.t623 486.048
R9246 VPWR.t738 VPWR.t1016 486.048
R9247 VPWR.t1828 VPWR.t737 486.048
R9248 VPWR.t1919 VPWR.t1470 486.048
R9249 VPWR.t1639 VPWR.t1918 486.048
R9250 VPWR.t1076 VPWR.t1714 486.048
R9251 VPWR.t1435 VPWR.t625 486.048
R9252 VPWR.t1107 VPWR.t1391 486.048
R9253 VPWR.t1243 VPWR.t1121 486.048
R9254 VPWR.t1249 VPWR.t1256 486.048
R9255 VPWR.t1360 VPWR.t1290 486.048
R9256 VPWR.t1407 VPWR.t1137 486.048
R9257 VPWR.t1284 VPWR.t1165 486.048
R9258 VPWR.t1180 VPWR.t1401 486.048
R9259 VPWR.t1432 VPWR.t1412 486.048
R9260 VPWR.t1446 VPWR.t1177 486.048
R9261 VPWR.t1281 VPWR.t1163 486.048
R9262 VPWR.t1316 VPWR.t1440 486.048
R9263 VPWR.t1459 VPWR.t1341 486.048
R9264 VPWR.t1188 VPWR.t1203 486.048
R9265 VPWR.t1214 VPWR.t1335 486.048
R9266 VPWR.t1239 VPWR.t1369 486.048
R9267 VPWR.t1084 VPWR.t1211 486.048
R9268 VPWR.t1236 VPWR.t1105 486.048
R9269 VPWR.t1374 VPWR.t1241 486.048
R9270 VPWR.t1383 VPWR.t1380 486.048
R9271 VPWR.t1145 VPWR.t1417 486.048
R9272 VPWR.t1135 VPWR.t1253 486.048
R9273 VPWR.t1414 VPWR.t1279 486.048
R9274 VPWR.t1303 VPWR.t1132 486.048
R9275 VPWR.t1167 VPWR.t1140 486.048
R9276 VPWR.t1175 VPWR.t1295 486.048
R9277 VPWR.t1366 VPWR.t1277 486.048
R9278 VPWR.t1438 VPWR.t1172 486.048
R9279 VPWR.t1190 VPWR.t1457 486.048
R9280 VPWR.t1311 VPWR.t1318 486.048
R9281 VPWR.t1451 VPWR.t1333 486.048
R9282 VPWR.t1355 VPWR.t1091 486.048
R9283 VPWR.t1330 VPWR.t1206 486.048
R9284 VPWR.t926 VPWR.t619 463.954
R9285 VPWR.t104 VPWR.t796 463.954
R9286 VPWR.t1629 VPWR.t861 463.954
R9287 VPWR.t1538 VPWR.t929 463.954
R9288 VPWR.t732 VPWR.t1766 463.954
R9289 VPWR.t102 VPWR.t161 463.954
R9290 VPWR.t169 VPWR.t865 463.954
R9291 VPWR.t1765 VPWR.t481 463.954
R9292 VPWR.t425 VPWR.t518 463.954
R9293 VPWR.t103 VPWR.t120 463.954
R9294 VPWR.t362 VPWR.t928 463.954
R9295 VPWR.t1577 VPWR.t927 463.954
R9296 VPWR.t864 VPWR.t1600 463.954
R9297 VPWR.t189 VPWR.t863 463.954
R9298 VPWR.t862 VPWR.t12 463.954
R9299 VPWR.t424 VPWR.t582 463.954
R9300 VPWR.t885 VPWR.t609 463.954
R9301 VPWR.t1691 VPWR.t154 463.954
R9302 VPWR.t848 VPWR.t254 463.954
R9303 VPWR.t1514 VPWR.t847 463.954
R9304 VPWR.t884 VPWR.t1062 463.954
R9305 VPWR.t323 VPWR.t498 463.954
R9306 VPWR.t1881 VPWR.t322 463.954
R9307 VPWR.t68 VPWR.t883 463.954
R9308 VPWR.t156 VPWR.t866 463.954
R9309 VPWR.t1573 VPWR.t324 463.954
R9310 VPWR.t846 VPWR.t301 463.954
R9311 VPWR.t886 VPWR.t1008 463.954
R9312 VPWR.t902 VPWR.t321 463.954
R9313 VPWR.t320 VPWR.t202 463.954
R9314 VPWR.t969 VPWR.t849 463.954
R9315 VPWR.t155 VPWR.t992 463.954
R9316 VPWR.t1657 VPWR.t595 463.954
R9317 VPWR.t1652 VPWR.t702 463.954
R9318 VPWR.t328 VPWR.t939 463.954
R9319 VPWR.t1492 VPWR.t327 463.954
R9320 VPWR.t1656 VPWR.t820 463.954
R9321 VPWR.t1584 VPWR.t1650 463.954
R9322 VPWR.t1649 VPWR.t1851 463.954
R9323 VPWR.t1841 VPWR.t1655 463.954
R9324 VPWR.t1654 VPWR.t54 463.954
R9325 VPWR.t670 VPWR.t1651 463.954
R9326 VPWR.t326 VPWR.t1895 463.954
R9327 VPWR.t747 VPWR.t325 463.954
R9328 VPWR.t331 VPWR.t1606 463.954
R9329 VPWR.t330 VPWR.t1472 463.954
R9330 VPWR.t1707 VPWR.t329 463.954
R9331 VPWR.t1653 VPWR.t1722 463.954
R9332 VPWR.t318 VPWR.t603 463.954
R9333 VPWR.t313 VPWR.t252 463.954
R9334 VPWR.t508 VPWR.t399 463.954
R9335 VPWR.t1506 VPWR.t398 463.954
R9336 VPWR.t1068 VPWR.t317 463.954
R9337 VPWR.t1779 VPWR.t299 463.954
R9338 VPWR.t298 VPWR.t432 463.954
R9339 VPWR.t78 VPWR.t316 463.954
R9340 VPWR.t719 VPWR.t315 463.954
R9341 VPWR.t300 VPWR.t887 463.954
R9342 VPWR.t397 VPWR.t307 463.954
R9343 VPWR.t1018 VPWR.t319 463.954
R9344 VPWR.t297 VPWR.t1822 463.954
R9345 VPWR.t210 VPWR.t296 463.954
R9346 VPWR.t1633 VPWR.t295 463.954
R9347 VPWR.t314 VPWR.t998 463.954
R9348 VPWR.t850 VPWR.t615 463.954
R9349 VPWR.t105 VPWR.t248 463.954
R9350 VPWR.t961 VPWR.t496 463.954
R9351 VPWR.t495 VPWR.t1526 463.954
R9352 VPWR.t1793 VPWR.t565 463.954
R9353 VPWR.t1742 VPWR.t294 463.954
R9354 VPWR.t293 VPWR.t407 463.954
R9355 VPWR.t465 VPWR.t564 463.954
R9356 VPWR.t563 VPWR.t110 463.954
R9357 VPWR.t421 VPWR.t1581 463.954
R9358 VPWR.t852 VPWR.t265 463.954
R9359 VPWR.t1022 VPWR.t851 463.954
R9360 VPWR.t908 VPWR.t292 463.954
R9361 VPWR.t1052 VPWR.t291 463.954
R9362 VPWR.t497 VPWR.t1905 463.954
R9363 VPWR.t524 VPWR.t562 463.954
R9364 VPWR.t881 VPWR.t621 463.954
R9365 VPWR.t794 VPWR.t1646 463.954
R9366 VPWR.t536 VPWR.t1627 463.954
R9367 VPWR.t1540 VPWR.t743 463.954
R9368 VPWR.t730 VPWR.t880 463.954
R9369 VPWR.t32 VPWR.t159 463.954
R9370 VPWR.t167 VPWR.t31 463.954
R9371 VPWR.t879 VPWR.t479 463.954
R9372 VPWR.t516 VPWR.t1648 463.954
R9373 VPWR.t33 VPWR.t662 463.954
R9374 VPWR.t742 VPWR.t360 463.954
R9375 VPWR.t1575 VPWR.t741 463.954
R9376 VPWR.t30 VPWR.t1598 463.954
R9377 VPWR.t187 VPWR.t538 463.954
R9378 VPWR.t10 VPWR.t537 463.954
R9379 VPWR.t580 VPWR.t1647 463.954
R9380 VPWR.t901 VPWR.t617 463.954
R9381 VPWR.t1687 VPWR.t1037 463.954
R9382 VPWR.t1661 VPWR.t774 463.954
R9383 VPWR.t1534 VPWR.t1660 463.954
R9384 VPWR.t900 VPWR.t734 463.954
R9385 VPWR.t1035 VPWR.t1699 463.954
R9386 VPWR.t1802 VPWR.t1034 463.954
R9387 VPWR.t899 VPWR.t461 463.954
R9388 VPWR.t650 VPWR.t898 463.954
R9389 VPWR.t1036 VPWR.t126 463.954
R9390 VPWR.t368 VPWR.t1659 463.954
R9391 VPWR.t765 VPWR.t1658 463.954
R9392 VPWR.t1033 VPWR.t1812 463.954
R9393 VPWR.t191 VPWR.t1663 463.954
R9394 VPWR.t1662 VPWR.t18 463.954
R9395 VPWR.t897 VPWR.t584 463.954
R9396 VPWR.t1622 VPWR.t597 463.954
R9397 VPWR.t700 VPWR.t1617 463.954
R9398 VPWR.t443 VPWR.t937 463.954
R9399 VPWR.t442 VPWR.t1494 463.954
R9400 VPWR.t816 VPWR.t1621 463.954
R9401 VPWR.t1582 VPWR.t448 463.954
R9402 VPWR.t1849 VPWR.t447 463.954
R9403 VPWR.t1839 VPWR.t1620 463.954
R9404 VPWR.t1619 VPWR.t808 463.954
R9405 VPWR.t1616 VPWR.t668 463.954
R9406 VPWR.t1893 VPWR.t441 463.954
R9407 VPWR.t440 VPWR.t745 463.954
R9408 VPWR.t1604 VPWR.t446 463.954
R9409 VPWR.t445 VPWR.t1468 463.954
R9410 VPWR.t444 VPWR.t1705 463.954
R9411 VPWR.t1718 VPWR.t1618 463.954
R9412 VPWR.t876 VPWR.t613 463.954
R9413 VPWR.t1809 VPWR.t1564 463.954
R9414 VPWR.t963 VPWR.t685 463.954
R9415 VPWR.t684 VPWR.t1524 463.954
R9416 VPWR.t707 VPWR.t875 463.954
R9417 VPWR.t690 VPWR.t1744 463.954
R9418 VPWR.t409 VPWR.t689 463.954
R9419 VPWR.t874 VPWR.t467 463.954
R9420 VPWR.t112 VPWR.t873 463.954
R9421 VPWR.t691 VPWR.t566 463.954
R9422 VPWR.t267 VPWR.t878 463.954
R9423 VPWR.t877 VPWR.t1024 463.954
R9424 VPWR.t688 VPWR.t910 463.954
R9425 VPWR.t1054 VPWR.t687 463.954
R9426 VPWR.t686 VPWR.t1907 463.954
R9427 VPWR.t526 VPWR.t872 463.954
R9428 VPWR.t1808 VPWR.t599 463.954
R9429 VPWR.t1915 VPWR.t698 463.954
R9430 VPWR.t197 VPWR.t1623 463.954
R9431 VPWR.t1496 VPWR.t196 463.954
R9432 VPWR.t1807 VPWR.t814 463.954
R9433 VPWR.t924 VPWR.t1913 463.954
R9434 VPWR.t201 VPWR.t1847 463.954
R9435 VPWR.t1806 VPWR.t1837 463.954
R9436 VPWR.t1917 VPWR.t804 463.954
R9437 VPWR.t666 VPWR.t1914 463.954
R9438 VPWR.t195 VPWR.t1891 463.954
R9439 VPWR.t220 VPWR.t1922 463.954
R9440 VPWR.t200 VPWR.t1614 463.954
R9441 VPWR.t1464 VPWR.t199 463.954
R9442 VPWR.t198 VPWR.t1703 463.954
R9443 VPWR.t1716 VPWR.t1916 463.954
R9444 VPWR.t1645 VPWR.t611 463.954
R9445 VPWR.t1670 VPWR.t1566 463.954
R9446 VPWR.t976 VPWR.t965 463.954
R9447 VPWR.t1522 VPWR.t975 463.954
R9448 VPWR.t711 VPWR.t1644 463.954
R9449 VPWR.t1675 VPWR.t1746 463.954
R9450 VPWR.t411 VPWR.t1674 463.954
R9451 VPWR.t1643 VPWR.t469 463.954
R9452 VPWR.t1642 VPWR.t0 463.954
R9453 VPWR.t568 VPWR.t1676 463.954
R9454 VPWR.t974 VPWR.t269 463.954
R9455 VPWR.t1026 VPWR.t973 463.954
R9456 VPWR.t1673 VPWR.t1542 463.954
R9457 VPWR.t1056 VPWR.t1672 463.954
R9458 VPWR.t1671 VPWR.t1909 463.954
R9459 VPWR.t530 VPWR.t1641 463.954
R9460 VPWR.t101 VPWR.t605 463.954
R9461 VPWR.t1904 VPWR.t250 463.954
R9462 VPWR.t504 VPWR.t131 463.954
R9463 VPWR.t130 VPWR.t1508 463.954
R9464 VPWR.t100 VPWR.t1066 463.954
R9465 VPWR.t1775 VPWR.t1902 463.954
R9466 VPWR.t428 VPWR.t1901 463.954
R9467 VPWR.t74 VPWR.t99 463.954
R9468 VPWR.t98 VPWR.t717 463.954
R9469 VPWR.t1042 VPWR.t1903 463.954
R9470 VPWR.t129 VPWR.t305 463.954
R9471 VPWR.t1014 VPWR.t128 463.954
R9472 VPWR.t1820 VPWR.t1900 463.954
R9473 VPWR.t1899 VPWR.t208 463.954
R9474 VPWR.t1631 VPWR.t835 463.954
R9475 VPWR.t97 VPWR.t996 463.954
R9476 VPWR.t935 VPWR.t601 463.954
R9477 VPWR.t1762 VPWR.t483 463.954
R9478 VPWR.t510 VPWR.t1748 463.954
R9479 VPWR.t1757 VPWR.t1504 463.954
R9480 VPWR.t934 VPWR.t1072 463.954
R9481 VPWR.t1781 VPWR.t1740 463.954
R9482 VPWR.t1739 VPWR.t434 463.954
R9483 VPWR.t933 VPWR.t80 463.954
R9484 VPWR.t721 VPWR.t1764 463.954
R9485 VPWR.t1741 VPWR.t889 463.954
R9486 VPWR.t1756 VPWR.t309 463.954
R9487 VPWR.t1020 VPWR.t936 463.954
R9488 VPWR.t1738 VPWR.t1824 463.954
R9489 VPWR.t1737 VPWR.t212 463.954
R9490 VPWR.t1635 VPWR.t1736 463.954
R9491 VPWR.t1763 VPWR.t1002 463.954
R9492 VPWR.t1859 VPWR.t590 463.954
R9493 VPWR.t90 VPWR.t704 463.954
R9494 VPWR.t1863 VPWR.t945 463.954
R9495 VPWR.t1486 VPWR.t1862 463.954
R9496 VPWR.t744 VPWR.t826 463.954
R9497 VPWR.t1590 VPWR.t88 463.954
R9498 VPWR.t87 VPWR.t1857 463.954
R9499 VPWR.t279 VPWR.t1767 463.954
R9500 VPWR.t278 VPWR.t58 463.954
R9501 VPWR.t656 VPWR.t89 463.954
R9502 VPWR.t1861 VPWR.t1897 463.954
R9503 VPWR.t753 VPWR.t1860 463.954
R9504 VPWR.t86 VPWR.t1608 463.954
R9505 VPWR.t1476 VPWR.t1865 463.954
R9506 VPWR.t1864 VPWR.t20 463.954
R9507 VPWR.t277 VPWR.t576 463.954
R9508 VPWR.t1170 VPWR.t1185 463.954
R9509 VPWR.t1301 VPWR.t1321 463.954
R9510 VPWR.t1448 VPWR.t1430 463.954
R9511 VPWR.t1086 VPWR.t1219 463.954
R9512 VPWR.t1196 VPWR.t1324 463.954
R9513 VPWR.t1346 VPWR.t1351 463.954
R9514 VPWR.t1353 VPWR.t1094 463.954
R9515 VPWR.t1216 VPWR.t1201 463.954
R9516 VPWR.t1231 VPWR.t1357 463.954
R9517 VPWR.t1385 VPWR.t1349 463.954
R9518 VPWR.t1100 VPWR.t1113 463.954
R9519 VPWR.t1116 VPWR.t1246 463.954
R9520 VPWR.t1287 VPWR.t1372 463.954
R9521 VPWR.t1123 VPWR.t1393 463.954
R9522 VPWR.t1422 VPWR.t1157 463.954
R9523 VPWR.t1251 VPWR.t1268 463.954
R9524 VPWR.t736 VPWR.t607 463.954
R9525 VPWR.t624 VPWR.t1693 463.954
R9526 VPWR.t256 VPWR.t740 463.954
R9527 VPWR.t739 VPWR.t1512 463.954
R9528 VPWR.t1064 VPWR.t628 463.954
R9529 VPWR.t1921 VPWR.t500 463.954
R9530 VPWR.t1883 VPWR.t1920 463.954
R9531 VPWR.t627 VPWR.t70 463.954
R9532 VPWR.t870 VPWR.t626 463.954
R9533 VPWR.t623 VPWR.t1038 463.954
R9534 VPWR.t303 VPWR.t738 463.954
R9535 VPWR.t737 VPWR.t1010 463.954
R9536 VPWR.t904 VPWR.t1919 463.954
R9537 VPWR.t1918 VPWR.t206 463.954
R9538 VPWR.t971 VPWR.t1076 463.954
R9539 VPWR.t625 VPWR.t994 463.954
R9540 VPWR.t1391 VPWR.t1398 463.954
R9541 VPWR.t1121 VPWR.t1160 463.954
R9542 VPWR.t1262 VPWR.t1249 463.954
R9543 VPWR.t1290 VPWR.t1424 463.954
R9544 VPWR.t1142 VPWR.t1407 463.954
R9545 VPWR.t1165 VPWR.t1154 463.954
R9546 VPWR.t1313 VPWR.t1180 463.954
R9547 VPWR.t1412 VPWR.t1363 463.954
R9548 VPWR.t1182 VPWR.t1446 463.954
R9549 VPWR.t1163 VPWR.t1208 463.954
R9550 VPWR.t1338 VPWR.t1316 463.954
R9551 VPWR.t1341 VPWR.t1081 463.954
R9552 VPWR.t1102 VPWR.t1188 463.954
R9553 VPWR.t1343 VPWR.t1214 463.954
R9554 VPWR.t1377 VPWR.t1239 463.954
R9555 VPWR.t1088 VPWR.t1084 463.954
R9556 VPWR.t1105 VPWR.t1129 463.954
R9557 VPWR.t1241 VPWR.t1274 463.954
R9558 VPWR.t1395 VPWR.t1383 463.954
R9559 VPWR.t1417 VPWR.t1151 463.954
R9560 VPWR.t1259 VPWR.t1135 463.954
R9561 VPWR.t1279 VPWR.t1271 463.954
R9562 VPWR.t1427 VPWR.t1303 463.954
R9563 VPWR.t1140 VPWR.t1148 463.954
R9564 VPWR.t1308 VPWR.t1175 463.954
R9565 VPWR.t1277 VPWR.t1327 463.954
R9566 VPWR.t1454 VPWR.t1438 463.954
R9567 VPWR.t1457 VPWR.t1198 463.954
R9568 VPWR.t1228 VPWR.t1311 463.954
R9569 VPWR.t1333 VPWR.t1078 463.954
R9570 VPWR.t1097 VPWR.t1355 463.954
R9571 VPWR.t1206 VPWR.t1222 463.954
R9572 VPWR.n2915 VPWR.t136 428.822
R9573 VPWR.t592 VPWR.n3105 376.524
R9574 VPWR.n1633 VPWR.n1632 376.045
R9575 VPWR.n1625 VPWR.n1624 376.045
R9576 VPWR.n1644 VPWR.n1643 376.045
R9577 VPWR.n1646 VPWR.n1645 376.045
R9578 VPWR.n1651 VPWR.n1650 376.045
R9579 VPWR.n1653 VPWR.n1652 376.045
R9580 VPWR.n1658 VPWR.n1657 376.045
R9581 VPWR.n1660 VPWR.n1659 376.045
R9582 VPWR.n1741 VPWR.n1740 376.045
R9583 VPWR.n1746 VPWR.n1745 376.045
R9584 VPWR.n1748 VPWR.n1747 376.045
R9585 VPWR.n903 VPWR.n902 376.045
R9586 VPWR.n900 VPWR.n899 376.045
R9587 VPWR.n1759 VPWR.n1758 376.045
R9588 VPWR.n1824 VPWR.n1823 376.045
R9589 VPWR.n1822 VPWR.n1821 376.045
R9590 VPWR.n2533 VPWR.n2532 376.045
R9591 VPWR.n2535 VPWR.n2534 376.045
R9592 VPWR.n2540 VPWR.n2539 376.045
R9593 VPWR.n2542 VPWR.n2541 376.045
R9594 VPWR.n495 VPWR.n494 376.045
R9595 VPWR.n497 VPWR.n496 376.045
R9596 VPWR.n492 VPWR.n490 376.045
R9597 VPWR.n2513 VPWR.n2512 376.045
R9598 VPWR.n2516 VPWR.n2515 376.045
R9599 VPWR.n2522 VPWR.n2521 376.045
R9600 VPWR.n2520 VPWR.n2519 376.045
R9601 VPWR.n2646 VPWR.n2645 376.045
R9602 VPWR.n2648 VPWR.n2647 376.045
R9603 VPWR.n2658 VPWR.n2657 376.045
R9604 VPWR.n2661 VPWR.n2660 376.045
R9605 VPWR.n2441 VPWR.n2440 376.045
R9606 VPWR.n2443 VPWR.n2442 376.045
R9607 VPWR.n2436 VPWR.n2435 376.045
R9608 VPWR.n2433 VPWR.n2432 376.045
R9609 VPWR.n2428 VPWR.n2427 376.045
R9610 VPWR.n2426 VPWR.n2425 376.045
R9611 VPWR.n487 VPWR.n486 376.045
R9612 VPWR.n2464 VPWR.n2463 376.045
R9613 VPWR.n2466 VPWR.n2465 376.045
R9614 VPWR.n2471 VPWR.n2470 376.045
R9615 VPWR.n2476 VPWR.n2475 376.045
R9616 VPWR.n2478 VPWR.n2477 376.045
R9617 VPWR.n2484 VPWR.n2483 376.045
R9618 VPWR.n2486 VPWR.n2485 376.045
R9619 VPWR.n2492 VPWR.n2491 376.045
R9620 VPWR.n2394 VPWR.n2393 376.045
R9621 VPWR.n2399 VPWR.n2398 376.045
R9622 VPWR.n2401 VPWR.n2400 376.045
R9623 VPWR.n2406 VPWR.n2405 376.045
R9624 VPWR.n2408 VPWR.n2407 376.045
R9625 VPWR.n512 VPWR.n511 376.045
R9626 VPWR.n509 VPWR.n508 376.045
R9627 VPWR.n2392 VPWR.n2391 376.045
R9628 VPWR.n2387 VPWR.n2386 376.045
R9629 VPWR.n2385 VPWR.n2384 376.045
R9630 VPWR.n2380 VPWR.n2379 376.045
R9631 VPWR.n2378 VPWR.n2377 376.045
R9632 VPWR.n533 VPWR.n532 376.045
R9633 VPWR.n2368 VPWR.n2367 376.045
R9634 VPWR.n2366 VPWR.n2365 376.045
R9635 VPWR.n572 VPWR.n571 376.045
R9636 VPWR.n2287 VPWR.n2286 376.045
R9637 VPWR.n2289 VPWR.n2288 376.045
R9638 VPWR.n691 VPWR.n690 376.045
R9639 VPWR.n695 VPWR.n694 376.045
R9640 VPWR.n697 VPWR.n696 376.045
R9641 VPWR.n688 VPWR.n685 376.045
R9642 VPWR.n570 VPWR.n569 376.045
R9643 VPWR.n2311 VPWR.n2310 376.045
R9644 VPWR.n2314 VPWR.n2313 376.045
R9645 VPWR.n2329 VPWR.n2328 376.045
R9646 VPWR.n2327 VPWR.n2326 376.045
R9647 VPWR.n2322 VPWR.n2321 376.045
R9648 VPWR.n2320 VPWR.n2319 376.045
R9649 VPWR.n2352 VPWR.n2351 376.045
R9650 VPWR.n663 VPWR.n662 376.045
R9651 VPWR.n668 VPWR.n667 376.045
R9652 VPWR.n672 VPWR.n671 376.045
R9653 VPWR.n674 VPWR.n673 376.045
R9654 VPWR.n679 VPWR.n678 376.045
R9655 VPWR.n681 VPWR.n680 376.045
R9656 VPWR.n632 VPWR.n629 376.045
R9657 VPWR.n661 VPWR.n660 376.045
R9658 VPWR.n656 VPWR.n655 376.045
R9659 VPWR.n654 VPWR.n653 376.045
R9660 VPWR.n649 VPWR.n648 376.045
R9661 VPWR.n647 VPWR.n646 376.045
R9662 VPWR.n2267 VPWR.n2266 376.045
R9663 VPWR.n2265 VPWR.n2264 376.045
R9664 VPWR.n2260 VPWR.n2259 376.045
R9665 VPWR.n2168 VPWR.n2167 376.045
R9666 VPWR.n2158 VPWR.n2157 376.045
R9667 VPWR.n2156 VPWR.n2155 376.045
R9668 VPWR.n2142 VPWR.n2141 376.045
R9669 VPWR.n2144 VPWR.n2143 376.045
R9670 VPWR.n2139 VPWR.n2138 376.045
R9671 VPWR.n626 VPWR.n625 376.045
R9672 VPWR.n2170 VPWR.n2169 376.045
R9673 VPWR.n2180 VPWR.n2179 376.045
R9674 VPWR.n2183 VPWR.n2182 376.045
R9675 VPWR.n2197 VPWR.n2196 376.045
R9676 VPWR.n2195 VPWR.n2194 376.045
R9677 VPWR.n2190 VPWR.n2189 376.045
R9678 VPWR.n2188 VPWR.n2187 376.045
R9679 VPWR.n2240 VPWR.n2239 376.045
R9680 VPWR.n2113 VPWR.n2112 376.045
R9681 VPWR.n2115 VPWR.n2114 376.045
R9682 VPWR.n2089 VPWR.n2088 376.045
R9683 VPWR.n2086 VPWR.n2085 376.045
R9684 VPWR.n2080 VPWR.n2079 376.045
R9685 VPWR.n2078 VPWR.n2077 376.045
R9686 VPWR.n2073 VPWR.n2072 376.045
R9687 VPWR.n2108 VPWR.n2107 376.045
R9688 VPWR.n2106 VPWR.n2105 376.045
R9689 VPWR.n2101 VPWR.n2100 376.045
R9690 VPWR.n2099 VPWR.n2098 376.045
R9691 VPWR.n2214 VPWR.n2213 376.045
R9692 VPWR.n2216 VPWR.n2215 376.045
R9693 VPWR.n2222 VPWR.n2221 376.045
R9694 VPWR.n2225 VPWR.n2224 376.045
R9695 VPWR.n2058 VPWR.n2057 376.045
R9696 VPWR.n1939 VPWR.n1938 376.045
R9697 VPWR.n1943 VPWR.n1942 376.045
R9698 VPWR.n1945 VPWR.n1944 376.045
R9699 VPWR.n1936 VPWR.n1935 376.045
R9700 VPWR.n1933 VPWR.n1932 376.045
R9701 VPWR.n1924 VPWR.n1923 376.045
R9702 VPWR.n2056 VPWR.n2055 376.045
R9703 VPWR.n723 VPWR.n722 376.045
R9704 VPWR.n2046 VPWR.n2045 376.045
R9705 VPWR.n2044 VPWR.n2043 376.045
R9706 VPWR.n2039 VPWR.n2038 376.045
R9707 VPWR.n2037 VPWR.n2036 376.045
R9708 VPWR.n735 VPWR.n734 376.045
R9709 VPWR.n2027 VPWR.n2026 376.045
R9710 VPWR.n1963 VPWR.n1962 376.045
R9711 VPWR.n777 VPWR.n776 376.045
R9712 VPWR.n782 VPWR.n781 376.045
R9713 VPWR.n784 VPWR.n783 376.045
R9714 VPWR.n789 VPWR.n788 376.045
R9715 VPWR.n791 VPWR.n790 376.045
R9716 VPWR.n770 VPWR.n767 376.045
R9717 VPWR.n1965 VPWR.n1964 376.045
R9718 VPWR.n1971 VPWR.n1970 376.045
R9719 VPWR.n1973 VPWR.n1972 376.045
R9720 VPWR.n1987 VPWR.n1986 376.045
R9721 VPWR.n1990 VPWR.n1989 376.045
R9722 VPWR.n2004 VPWR.n2003 376.045
R9723 VPWR.n2002 VPWR.n2001 376.045
R9724 VPWR.n1997 VPWR.n1996 376.045
R9725 VPWR.n819 VPWR.n818 376.045
R9726 VPWR.n1901 VPWR.n1900 376.045
R9727 VPWR.n1903 VPWR.n1902 376.045
R9728 VPWR.n1908 VPWR.n1907 376.045
R9729 VPWR.n1910 VPWR.n1909 376.045
R9730 VPWR.n805 VPWR.n804 376.045
R9731 VPWR.n802 VPWR.n801 376.045
R9732 VPWR.n822 VPWR.n821 376.045
R9733 VPWR.n1890 VPWR.n1889 376.045
R9734 VPWR.n1888 VPWR.n1887 376.045
R9735 VPWR.n1883 VPWR.n1882 376.045
R9736 VPWR.n1881 VPWR.n1880 376.045
R9737 VPWR.n1876 VPWR.n1875 376.045
R9738 VPWR.n1874 VPWR.n1873 376.045
R9739 VPWR.n836 VPWR.n835 376.045
R9740 VPWR.n2581 VPWR.n2580 376.045
R9741 VPWR.n2563 VPWR.n2562 376.045
R9742 VPWR.n2565 VPWR.n2564 376.045
R9743 VPWR.n2558 VPWR.n2557 376.045
R9744 VPWR.n2555 VPWR.n2554 376.045
R9745 VPWR.n2583 VPWR.n2582 376.045
R9746 VPWR.n2589 VPWR.n2588 376.045
R9747 VPWR.n2592 VPWR.n2591 376.045
R9748 VPWR.n2626 VPWR.n2625 376.045
R9749 VPWR.n2624 VPWR.n2623 376.045
R9750 VPWR.n2619 VPWR.n2618 376.045
R9751 VPWR.n2617 VPWR.n2616 376.045
R9752 VPWR.n2612 VPWR.n2611 376.045
R9753 VPWR.n2610 VPWR.n2609 376.045
R9754 VPWR.n2605 VPWR.n2604 376.045
R9755 VPWR.n1793 VPWR.n1792 376.045
R9756 VPWR.n1798 VPWR.n1797 376.045
R9757 VPWR.n1800 VPWR.n1799 376.045
R9758 VPWR.n1790 VPWR.n1789 376.045
R9759 VPWR.n1787 VPWR.n1786 376.045
R9760 VPWR.n1782 VPWR.n1781 376.045
R9761 VPWR.n1780 VPWR.n1779 376.045
R9762 VPWR.n1834 VPWR.n1833 376.045
R9763 VPWR.n1839 VPWR.n1838 376.045
R9764 VPWR.n1837 VPWR.n1836 376.045
R9765 VPWR.n1849 VPWR.n1848 376.045
R9766 VPWR.n1851 VPWR.n1850 376.045
R9767 VPWR.n1857 VPWR.n1856 376.045
R9768 VPWR.n2731 VPWR.n2730 376.045
R9769 VPWR.n2733 VPWR.n2732 376.045
R9770 VPWR.n376 VPWR.n373 376.045
R9771 VPWR.n385 VPWR.n384 376.045
R9772 VPWR.n2721 VPWR.n2720 376.045
R9773 VPWR.n2719 VPWR.n2718 376.045
R9774 VPWR.n394 VPWR.n393 376.045
R9775 VPWR.n2709 VPWR.n2708 376.045
R9776 VPWR.n2707 VPWR.n2706 376.045
R9777 VPWR.n403 VPWR.n402 376.045
R9778 VPWR.n2697 VPWR.n2696 376.045
R9779 VPWR.n2695 VPWR.n2694 376.045
R9780 VPWR.n412 VPWR.n411 376.045
R9781 VPWR.n2685 VPWR.n2684 376.045
R9782 VPWR.n2683 VPWR.n2682 376.045
R9783 VPWR.n1761 VPWR.n1760 376.045
R9784 VPWR.n1766 VPWR.n1765 376.045
R9785 VPWR.n1768 VPWR.n1767 376.045
R9786 VPWR.n883 VPWR.n882 376.045
R9787 VPWR.n880 VPWR.n879 376.045
R9788 VPWR.n1739 VPWR.n1738 376.045
R9789 VPWR.n1734 VPWR.n1733 376.045
R9790 VPWR.n1732 VPWR.n1731 376.045
R9791 VPWR.n1721 VPWR.n1720 376.045
R9792 VPWR.n1205 VPWR.n1204 376.045
R9793 VPWR.n1199 VPWR.n1198 376.045
R9794 VPWR.n1193 VPWR.n1192 376.045
R9795 VPWR.n1191 VPWR.n1190 376.045
R9796 VPWR.n1631 VPWR.n1630 376.045
R9797 VPWR.n1705 VPWR.n1704 376.045
R9798 VPWR.n1711 VPWR.n1710 376.045
R9799 VPWR.n295 VPWR.n292 376.045
R9800 VPWR.n366 VPWR.n365 376.045
R9801 VPWR.n364 VPWR.n363 376.045
R9802 VPWR.n359 VPWR.n358 376.045
R9803 VPWR.n357 VPWR.n356 376.045
R9804 VPWR.n352 VPWR.n351 376.045
R9805 VPWR.n350 VPWR.n349 376.045
R9806 VPWR.n345 VPWR.n344 376.045
R9807 VPWR.n343 VPWR.n342 376.045
R9808 VPWR.n338 VPWR.n337 376.045
R9809 VPWR.n336 VPWR.n335 376.045
R9810 VPWR.n331 VPWR.n330 376.045
R9811 VPWR.n329 VPWR.n328 376.045
R9812 VPWR.n324 VPWR.n323 376.045
R9813 VPWR.n322 VPWR.n321 376.045
R9814 VPWR.n1163 VPWR.n1162 376.045
R9815 VPWR.n1673 VPWR.n1672 376.045
R9816 VPWR.n1671 VPWR.n1670 376.045
R9817 VPWR.n1279 VPWR.n1278 376.045
R9818 VPWR.n1488 VPWR.n1487 376.045
R9819 VPWR.n1490 VPWR.n1489 376.045
R9820 VPWR.n1500 VPWR.n1499 376.045
R9821 VPWR.n1502 VPWR.n1501 376.045
R9822 VPWR.n1514 VPWR.n1513 376.045
R9823 VPWR.n1516 VPWR.n1515 376.045
R9824 VPWR.n1523 VPWR.n1522 376.045
R9825 VPWR.n1533 VPWR.n1532 376.045
R9826 VPWR.n1531 VPWR.n1530 376.045
R9827 VPWR.n1526 VPWR.n1525 376.045
R9828 VPWR.n1589 VPWR.n1588 376.045
R9829 VPWR.n2764 VPWR.n2763 376.045
R9830 VPWR.n2774 VPWR.n2773 376.045
R9831 VPWR.n2776 VPWR.n2775 376.045
R9832 VPWR.n2786 VPWR.n2785 376.045
R9833 VPWR.n2788 VPWR.n2787 376.045
R9834 VPWR.n2798 VPWR.n2797 376.045
R9835 VPWR.n2800 VPWR.n2799 376.045
R9836 VPWR.n2810 VPWR.n2809 376.045
R9837 VPWR.n2812 VPWR.n2811 376.045
R9838 VPWR.n2822 VPWR.n2821 376.045
R9839 VPWR.n2824 VPWR.n2823 376.045
R9840 VPWR.n2834 VPWR.n2833 376.045
R9841 VPWR.n2836 VPWR.n2835 376.045
R9842 VPWR.n2846 VPWR.n2845 376.045
R9843 VPWR.n2762 VPWR.n2761 376.045
R9844 VPWR.n3112 VPWR.n3104 350.719
R9845 VPWR.n3112 VPWR.n3111 350.719
R9846 VPWR.n3107 VPWR.n25 350.719
R9847 VPWR.n3107 VPWR.n3106 350.719
R9848 VPWR.n1047 VPWR.t783 342.841
R9849 VPWR.n1086 VPWR.t677 342.841
R9850 VPWR.n1123 VPWR.t842 342.841
R9851 VPWR.n2982 VPWR.t375 342.841
R9852 VPWR.n2945 VPWR.t856 342.841
R9853 VPWR.n2888 VPWR.t137 342.841
R9854 VPWR.n1047 VPWR.t386 342.839
R9855 VPWR.n1086 VPWR.t1462 342.839
R9856 VPWR.n1123 VPWR.t986 342.839
R9857 VPWR.n2982 VPWR.t45 342.839
R9858 VPWR.n2945 VPWR.t552 342.839
R9859 VPWR.n2888 VPWR.t643 342.839
R9860 VPWR.n1014 VPWR.t787 338.488
R9861 VPWR.n3018 VPWR.t29 338.488
R9862 VPWR.n1023 VPWR.n1022 327.377
R9863 VPWR.n1016 VPWR.n1015 327.377
R9864 VPWR.n1030 VPWR.n1029 327.377
R9865 VPWR.n1060 VPWR.n1058 327.377
R9866 VPWR.n1053 VPWR.n1051 327.377
R9867 VPWR.n1068 VPWR.n1066 327.377
R9868 VPWR.n1099 VPWR.n1097 327.377
R9869 VPWR.n1092 VPWR.n1090 327.377
R9870 VPWR.n1107 VPWR.n1105 327.377
R9871 VPWR.n1136 VPWR.n1134 327.377
R9872 VPWR.n1129 VPWR.n1127 327.377
R9873 VPWR.n1144 VPWR.n1142 327.377
R9874 VPWR.n1032 VPWR.n1031 327.375
R9875 VPWR.n1060 VPWR.n1059 327.375
R9876 VPWR.n1053 VPWR.n1052 327.375
R9877 VPWR.n1068 VPWR.n1067 327.375
R9878 VPWR.n1099 VPWR.n1098 327.375
R9879 VPWR.n1092 VPWR.n1091 327.375
R9880 VPWR.n1107 VPWR.n1106 327.375
R9881 VPWR.n1136 VPWR.n1135 327.375
R9882 VPWR.n1129 VPWR.n1128 327.375
R9883 VPWR.n1144 VPWR.n1143 327.375
R9884 VPWR.n3118 VPWR.t1711 326.106
R9885 VPWR.n3122 VPWR.t799 326.106
R9886 VPWR.n3107 VPWR.t593 326.106
R9887 VPWR.n3112 VPWR.t594 326.106
R9888 VPWR.n1 VPWR 325.546
R9889 VPWR.n2956 VPWR.t44 322.262
R9890 VPWR.n2919 VPWR.t551 322.262
R9891 VPWR.n3094 VPWR.n3093 321.642
R9892 VPWR.n3011 VPWR.n3001 320.976
R9893 VPWR.n3005 VPWR.n3004 320.976
R9894 VPWR.n2999 VPWR.n2998 320.976
R9895 VPWR.n2969 VPWR.n2968 320.976
R9896 VPWR.n2975 VPWR.n2964 320.976
R9897 VPWR.n2961 VPWR.n2960 320.976
R9898 VPWR.n2932 VPWR.n2931 320.976
R9899 VPWR.n2938 VPWR.n2927 320.976
R9900 VPWR.n2924 VPWR.n2923 320.976
R9901 VPWR.n2899 VPWR.n2895 320.976
R9902 VPWR.n2903 VPWR.n2902 320.976
R9903 VPWR.n2909 VPWR.n2891 320.976
R9904 VPWR.n3016 VPWR.n2997 320.976
R9905 VPWR.n2969 VPWR.n2967 320.976
R9906 VPWR.n2975 VPWR.n2963 320.976
R9907 VPWR.n2961 VPWR.n2959 320.976
R9908 VPWR.n2932 VPWR.n2930 320.976
R9909 VPWR.n2938 VPWR.n2926 320.976
R9910 VPWR.n2924 VPWR.n2922 320.976
R9911 VPWR.n2899 VPWR.n2894 320.976
R9912 VPWR.n2903 VPWR.n2901 320.976
R9913 VPWR.n2909 VPWR.n2890 320.976
R9914 VPWR.n3090 VPWR 319.627
R9915 VPWR.n6 VPWR.n5 316.245
R9916 VPWR.n949 VPWR.n947 316.245
R9917 VPWR.n972 VPWR.n970 316.245
R9918 VPWR.n996 VPWR.n994 316.245
R9919 VPWR.n3073 VPWR.n3072 316.245
R9920 VPWR.n3053 VPWR.n3052 316.245
R9921 VPWR.n3034 VPWR.n3033 316.245
R9922 VPWR.n949 VPWR.n948 316.245
R9923 VPWR.n972 VPWR.n971 316.245
R9924 VPWR.n996 VPWR.n995 316.245
R9925 VPWR.n3073 VPWR.n3071 316.245
R9926 VPWR.n3053 VPWR.n3051 316.245
R9927 VPWR.n3034 VPWR.n3032 316.245
R9928 VPWR.n2919 VPWR.t258 313.87
R9929 VPWR.n10 VPWR.n4 310.502
R9930 VPWR.n954 VPWR.n946 310.502
R9931 VPWR.n977 VPWR.n969 310.502
R9932 VPWR.n1001 VPWR.n993 310.502
R9933 VPWR.n3092 VPWR.n3091 310.502
R9934 VPWR.n3077 VPWR.n3076 310.502
R9935 VPWR.n3057 VPWR.n3056 310.502
R9936 VPWR.n3038 VPWR.n3037 310.502
R9937 VPWR.n954 VPWR.n953 310.5
R9938 VPWR.n977 VPWR.n976 310.5
R9939 VPWR.n1001 VPWR.n1000 310.5
R9940 VPWR.n3077 VPWR.n3075 310.5
R9941 VPWR.n3057 VPWR.n3055 310.5
R9942 VPWR.n3038 VPWR.n3036 310.5
R9943 VPWR.t222 VPWR.t833 297.909
R9944 VPWR.n3125 VPWR.n3124 292.5
R9945 VPWR.n33 VPWR.n32 292.5
R9946 VPWR.n3109 VPWR.t592 272.257
R9947 VPWR.n3123 VPWR.n3122 256.226
R9948 VPWR.n3118 VPWR.n31 256.226
R9949 VPWR.n1120 VPWR.t423 255.905
R9950 VPWR.n2952 VPWR.t1568 255.905
R9951 VPWR.n983 VPWR.t561 255.904
R9952 VPWR.n1120 VPWR.t779 255.904
R9953 VPWR.n3063 VPWR.t634 255.904
R9954 VPWR.n2952 VPWR.t259 255.904
R9955 VPWR.n26 VPWR.n24 255.653
R9956 VPWR.n3117 VPWR.n35 255.653
R9957 VPWR.n1011 VPWR.t418 254.019
R9958 VPWR.n3024 VPWR.t1876 254.019
R9959 VPWR.n1043 VPWR.t416 252.948
R9960 VPWR.n3026 VPWR.t1874 252.948
R9961 VPWR.n1081 VPWR.t769 250.722
R9962 VPWR.n2989 VPWR.t182 250.722
R9963 VPWR.n1018 VPWR.t951 249.901
R9964 VPWR.n1054 VPWR.t1753 249.901
R9965 VPWR.n1093 VPWR.t1870 249.901
R9966 VPWR.n1130 VPWR.t1755 249.901
R9967 VPWR.n3003 VPWR.t390 249.901
R9968 VPWR.n2966 VPWR.t393 249.901
R9969 VPWR.n2929 VPWR.t288 249.901
R9970 VPWR.n2896 VPWR.t238 249.901
R9971 VPWR.n1054 VPWR.t1868 249.901
R9972 VPWR.n1093 VPWR.t1750 249.901
R9973 VPWR.n1130 VPWR.t917 249.901
R9974 VPWR.n2966 VPWR.t290 249.901
R9975 VPWR.n2929 VPWR.t240 249.901
R9976 VPWR.n2896 VPWR.t983 249.901
R9977 VPWR.n961 VPWR.t1571 249.363
R9978 VPWR.n1046 VPWR.t233 249.363
R9979 VPWR.n3100 VPWR.t958 249.363
R9980 VPWR.n3084 VPWR.t455 249.363
R9981 VPWR.n2987 VPWR.t641 249.363
R9982 VPWR.n17 VPWR.t832 249.362
R9983 VPWR.n961 VPWR.t65 249.362
R9984 VPWR.n3084 VPWR.t37 249.362
R9985 VPWR.t555 VPWR.t831 248.599
R9986 VPWR.t784 VPWR.t1730 248.599
R9987 VPWR.t1730 VPWR.t1734 248.599
R9988 VPWR.t1734 VPWR.t694 248.599
R9989 VPWR.t694 VPWR.t338 248.599
R9990 VPWR.t338 VPWR.t341 248.599
R9991 VPWR.t341 VPWR.t1752 248.599
R9992 VPWR.t1752 VPWR.t229 248.599
R9993 VPWR.t920 VPWR.t922 248.599
R9994 VPWR.t922 VPWR.t950 248.599
R9995 VPWR.t285 VPWR.t980 248.599
R9996 VPWR.t345 VPWR.t285 248.599
R9997 VPWR.t260 VPWR.t345 248.599
R9998 VPWR.t1030 VPWR.t260 248.599
R9999 VPWR.t148 VPWR.t1030 248.599
R10000 VPWR.t1923 VPWR.t148 248.599
R10001 VPWR.t967 VPWR.t1923 248.599
R10002 VPWR.t635 VPWR.t957 248.599
R10003 VPWR.t333 VPWR.t389 248.599
R10004 VPWR.t1888 VPWR.t333 248.599
R10005 VPWR.n15 VPWR.t556 247.394
R10006 VPWR.n959 VPWR.t560 247.394
R10007 VPWR.n3098 VPWR.t636 247.394
R10008 VPWR.n3082 VPWR.t630 247.394
R10009 VPWR.n959 VPWR.t558 247.394
R10010 VPWR.n3082 VPWR.t632 247.394
R10011 VPWR.n1012 VPWR.t954 244.737
R10012 VPWR.n3019 VPWR.t284 244.737
R10013 VPWR.n1082 VPWR.t727 243.886
R10014 VPWR.n2990 VPWR.t1553 243.886
R10015 VPWR.n985 VPWR.t830 243.512
R10016 VPWR.n1008 VPWR.t1572 243.512
R10017 VPWR.n1011 VPWR.t829 243.512
R10018 VPWR.n3065 VPWR.t960 243.512
R10019 VPWR.n3045 VPWR.t456 243.512
R10020 VPWR.n3024 VPWR.t639 243.512
R10021 VPWR.n1008 VPWR.t67 243.512
R10022 VPWR.n3045 VPWR.t35 243.512
R10023 VPWR.n1037 VPWR.t417 238.339
R10024 VPWR.n2994 VPWR.t1875 238.339
R10025 VPWR.n2956 VPWR.t640 234.982
R10026 VPWR.t918 VPWR.t920 228.101
R10027 VPWR.t402 VPWR.t1888 228.101
R10028 VPWR.n3090 VPWR 224.923
R10029 VPWR.n1 VPWR 219.004
R10030 VPWR.n1152 VPWR.n1151 214.613
R10031 VPWR.n1152 VPWR.n1150 214.613
R10032 VPWR.n944 VPWR.n943 214.326
R10033 VPWR.n967 VPWR.n966 214.326
R10034 VPWR.n991 VPWR.n990 214.326
R10035 VPWR.n1076 VPWR.n1075 214.326
R10036 VPWR.n1115 VPWR.n1114 214.326
R10037 VPWR.n944 VPWR.n942 214.326
R10038 VPWR.n967 VPWR.n965 214.326
R10039 VPWR.n991 VPWR.n989 214.326
R10040 VPWR.n1076 VPWR.n1074 214.326
R10041 VPWR.n1115 VPWR.n1113 214.326
R10042 VPWR.n2 VPWR.n1 213.119
R10043 VPWR.n3097 VPWR.n3090 213.119
R10044 VPWR VPWR.t555 207.166
R10045 VPWR VPWR.t967 201.246
R10046 VPWR.t833 VPWR.t798 200.262
R10047 VPWR.t950 VPWR 189.409
R10048 VPWR.n3030 VPWR 184.63
R10049 VPWR.n1037 VPWR 182.952
R10050 VPWR.n3049 VPWR 182.952
R10051 VPWR.n3069 VPWR 181.273
R10052 VPWR.t258 VPWR 177.916
R10053 VPWR.n1436 VPWR.n1434 161.365
R10054 VPWR.n1420 VPWR.n1418 161.365
R10055 VPWR.n1426 VPWR.n1424 161.365
R10056 VPWR.n1441 VPWR.n1439 161.365
R10057 VPWR.n1446 VPWR.n1444 161.365
R10058 VPWR.n1451 VPWR.n1449 161.365
R10059 VPWR.n1456 VPWR.n1454 161.365
R10060 VPWR.n1461 VPWR.n1459 161.365
R10061 VPWR.n1470 VPWR.n1468 161.365
R10062 VPWR.n1465 VPWR.n1463 161.365
R10063 VPWR.n1600 VPWR.n1598 161.365
R10064 VPWR.n1609 VPWR.n1607 161.365
R10065 VPWR.n1604 VPWR.n1602 161.365
R10066 VPWR.n935 VPWR.n933 161.365
R10067 VPWR.n1693 VPWR.n1691 161.365
R10068 VPWR.n1689 VPWR.n1687 161.365
R10069 VPWR VPWR.n2880 161.363
R10070 VPWR VPWR.n2878 161.363
R10071 VPWR VPWR.n2876 161.363
R10072 VPWR VPWR.n2874 161.363
R10073 VPWR VPWR.n2872 161.363
R10074 VPWR VPWR.n2870 161.363
R10075 VPWR VPWR.n2868 161.363
R10076 VPWR VPWR.n2866 161.363
R10077 VPWR VPWR.n2864 161.363
R10078 VPWR VPWR.n2862 161.363
R10079 VPWR VPWR.n2860 161.363
R10080 VPWR VPWR.n2858 161.363
R10081 VPWR VPWR.n2856 161.363
R10082 VPWR VPWR.n2854 161.363
R10083 VPWR VPWR.n2852 161.363
R10084 VPWR VPWR.n2850 161.363
R10085 VPWR.n1289 VPWR.n1288 161.303
R10086 VPWR.n94 VPWR.n93 161.303
R10087 VPWR.n1584 VPWR.n1583 161.3
R10088 VPWR.n1244 VPWR.n1243 161.3
R10089 VPWR.n1241 VPWR.n1240 161.3
R10090 VPWR.n1573 VPWR.n1572 161.3
R10091 VPWR.n1571 VPWR.n1570 161.3
R10092 VPWR.n1568 VPWR.n1567 161.3
R10093 VPWR.n1565 VPWR.n1564 161.3
R10094 VPWR.n1559 VPWR.n1558 161.3
R10095 VPWR.n1556 VPWR.n1555 161.3
R10096 VPWR.n1553 VPWR.n1552 161.3
R10097 VPWR.n1249 VPWR.n1248 161.3
R10098 VPWR.n1538 VPWR.n1537 161.3
R10099 VPWR.n1541 VPWR.n1540 161.3
R10100 VPWR.n1252 VPWR.n1251 161.3
R10101 VPWR.n1257 VPWR.n1256 161.3
R10102 VPWR.n1350 VPWR.n1349 161.3
R10103 VPWR.n1355 VPWR.n1354 161.3
R10104 VPWR.n1358 VPWR.n1357 161.3
R10105 VPWR.n1361 VPWR.n1360 161.3
R10106 VPWR.n1366 VPWR.n1365 161.3
R10107 VPWR.n1369 VPWR.n1368 161.3
R10108 VPWR.n1372 VPWR.n1371 161.3
R10109 VPWR.n1377 VPWR.n1376 161.3
R10110 VPWR.n1380 VPWR.n1379 161.3
R10111 VPWR.n1383 VPWR.n1382 161.3
R10112 VPWR.n1388 VPWR.n1387 161.3
R10113 VPWR.n1391 VPWR.n1390 161.3
R10114 VPWR.n1394 VPWR.n1393 161.3
R10115 VPWR.n1399 VPWR.n1398 161.3
R10116 VPWR.n1402 VPWR.n1401 161.3
R10117 VPWR.n1405 VPWR.n1404 161.3
R10118 VPWR.n1410 VPWR.n1409 161.3
R10119 VPWR.n1413 VPWR.n1412 161.3
R10120 VPWR.n1336 VPWR.n1335 161.3
R10121 VPWR.n1334 VPWR.n1333 161.3
R10122 VPWR.n1331 VPWR.n1330 161.3
R10123 VPWR.n1328 VPWR.n1327 161.3
R10124 VPWR.n1322 VPWR.n1321 161.3
R10125 VPWR.n1319 VPWR.n1318 161.3
R10126 VPWR.n1316 VPWR.n1315 161.3
R10127 VPWR.n1286 VPWR.n1285 161.3
R10128 VPWR.n1283 VPWR.n1282 161.3
R10129 VPWR.n1304 VPWR.n1303 161.3
R10130 VPWR.n1302 VPWR.n1301 161.3
R10131 VPWR.n1299 VPWR.n1298 161.3
R10132 VPWR.n1296 VPWR.n1295 161.3
R10133 VPWR.n1291 VPWR.n1290 161.3
R10134 VPWR.n92 VPWR.n91 161.3
R10135 VPWR.n289 VPWR.n288 161.3
R10136 VPWR.n286 VPWR.n285 161.3
R10137 VPWR.n88 VPWR.n87 161.3
R10138 VPWR.n273 VPWR.n272 161.3
R10139 VPWR.n276 VPWR.n275 161.3
R10140 VPWR.n270 VPWR.n269 161.3
R10141 VPWR.n267 VPWR.n266 161.3
R10142 VPWR.n264 VPWR.n263 161.3
R10143 VPWR.n258 VPWR.n257 161.3
R10144 VPWR.n255 VPWR.n254 161.3
R10145 VPWR.n252 VPWR.n251 161.3
R10146 VPWR.n103 VPWR.n102 161.3
R10147 VPWR.n239 VPWR.n238 161.3
R10148 VPWR.n242 VPWR.n241 161.3
R10149 VPWR.n236 VPWR.n235 161.3
R10150 VPWR.n233 VPWR.n232 161.3
R10151 VPWR.n230 VPWR.n229 161.3
R10152 VPWR.n224 VPWR.n223 161.3
R10153 VPWR.n221 VPWR.n220 161.3
R10154 VPWR.n218 VPWR.n217 161.3
R10155 VPWR.n108 VPWR.n107 161.3
R10156 VPWR.n205 VPWR.n204 161.3
R10157 VPWR.n208 VPWR.n207 161.3
R10158 VPWR.n202 VPWR.n201 161.3
R10159 VPWR.n199 VPWR.n198 161.3
R10160 VPWR.n196 VPWR.n195 161.3
R10161 VPWR.n190 VPWR.n189 161.3
R10162 VPWR.n187 VPWR.n186 161.3
R10163 VPWR.n184 VPWR.n183 161.3
R10164 VPWR.n113 VPWR.n112 161.3
R10165 VPWR.n171 VPWR.n170 161.3
R10166 VPWR.n174 VPWR.n173 161.3
R10167 VPWR.n168 VPWR.n167 161.3
R10168 VPWR.n165 VPWR.n164 161.3
R10169 VPWR.n162 VPWR.n161 161.3
R10170 VPWR.n156 VPWR.n155 161.3
R10171 VPWR.n153 VPWR.n152 161.3
R10172 VPWR.n150 VPWR.n149 161.3
R10173 VPWR.n118 VPWR.n117 161.3
R10174 VPWR.n137 VPWR.n136 161.3
R10175 VPWR.n140 VPWR.n139 161.3
R10176 VPWR.n134 VPWR.n133 161.3
R10177 VPWR.n131 VPWR.n130 161.3
R10178 VPWR.n96 VPWR.n95 161.3
R10179 VPWR.n128 VPWR.n127 161.3
R10180 VPWR.n123 VPWR.n122 161.3
R10181 VPWR.n1434 VPWR.t1429 161.202
R10182 VPWR.n1418 VPWR.t1300 161.202
R10183 VPWR.n1424 VPWR.t1169 161.202
R10184 VPWR.n1439 VPWR.t1085 161.202
R10185 VPWR.n1444 VPWR.t1195 161.202
R10186 VPWR.n1449 VPWR.t1350 161.202
R10187 VPWR.n1454 VPWR.t1352 161.202
R10188 VPWR.n1459 VPWR.t1200 161.202
R10189 VPWR.n1468 VPWR.t1230 161.202
R10190 VPWR.n1463 VPWR.t1348 161.202
R10191 VPWR.n1598 VPWR.t1099 161.202
R10192 VPWR.n1607 VPWR.t1115 161.202
R10193 VPWR.n1602 VPWR.t1371 161.202
R10194 VPWR.n933 VPWR.t1392 161.202
R10195 VPWR.n1691 VPWR.t1421 161.202
R10196 VPWR.n1687 VPWR.t1250 161.202
R10197 VPWR.n1243 VPWR.t1083 161.202
R10198 VPWR.n1570 VPWR.t1238 161.202
R10199 VPWR.n1558 VPWR.t1213 161.202
R10200 VPWR.n1248 VPWR.t1187 161.202
R10201 VPWR.n1251 VPWR.t1340 161.202
R10202 VPWR.n1354 VPWR.t1315 161.202
R10203 VPWR.n1365 VPWR.t1162 161.202
R10204 VPWR.n1376 VPWR.t1445 161.202
R10205 VPWR.n1387 VPWR.t1411 161.202
R10206 VPWR.n1398 VPWR.t1179 161.202
R10207 VPWR.n1409 VPWR.t1164 161.202
R10208 VPWR.n1333 VPWR.t1406 161.202
R10209 VPWR.n1321 VPWR.t1289 161.202
R10210 VPWR.n1285 VPWR.t1248 161.202
R10211 VPWR.n1301 VPWR.t1120 161.202
R10212 VPWR.n1290 VPWR.t1390 161.202
R10213 VPWR.n285 VPWR.t1240 161.202
R10214 VPWR.n275 VPWR.t1382 161.202
R10215 VPWR.n263 VPWR.t1416 161.202
R10216 VPWR.n251 VPWR.t1134 161.202
R10217 VPWR.n241 VPWR.t1278 161.202
R10218 VPWR.n229 VPWR.t1302 161.202
R10219 VPWR.n217 VPWR.t1139 161.202
R10220 VPWR.n207 VPWR.t1174 161.202
R10221 VPWR.n195 VPWR.t1276 161.202
R10222 VPWR.n183 VPWR.t1437 161.202
R10223 VPWR.n173 VPWR.t1456 161.202
R10224 VPWR.n161 VPWR.t1310 161.202
R10225 VPWR.n149 VPWR.t1332 161.202
R10226 VPWR.n139 VPWR.t1354 161.202
R10227 VPWR.n95 VPWR.t1104 161.202
R10228 VPWR.n127 VPWR.t1205 161.202
R10229 VPWR.n1583 VPWR.t1210 161.106
R10230 VPWR.n1572 VPWR.t1368 161.106
R10231 VPWR.n1564 VPWR.t1334 161.106
R10232 VPWR.n1552 VPWR.t1202 161.106
R10233 VPWR.n1540 VPWR.t1458 161.106
R10234 VPWR.n1349 VPWR.t1439 161.106
R10235 VPWR.n1360 VPWR.t1280 161.106
R10236 VPWR.n1371 VPWR.t1176 161.106
R10237 VPWR.n1382 VPWR.t1431 161.106
R10238 VPWR.n1393 VPWR.t1400 161.106
R10239 VPWR.n1404 VPWR.t1283 161.106
R10240 VPWR.n1335 VPWR.t1136 161.106
R10241 VPWR.n1327 VPWR.t1359 161.106
R10242 VPWR.n1315 VPWR.t1255 161.106
R10243 VPWR.n1303 VPWR.t1242 161.106
R10244 VPWR.n1295 VPWR.t1106 161.106
R10245 VPWR.n91 VPWR.t1235 161.106
R10246 VPWR.n87 VPWR.t1373 161.106
R10247 VPWR.n269 VPWR.t1379 161.106
R10248 VPWR.n257 VPWR.t1144 161.106
R10249 VPWR.n102 VPWR.t1252 161.106
R10250 VPWR.n235 VPWR.t1413 161.106
R10251 VPWR.n223 VPWR.t1131 161.106
R10252 VPWR.n107 VPWR.t1166 161.106
R10253 VPWR.n201 VPWR.t1294 161.106
R10254 VPWR.n189 VPWR.t1365 161.106
R10255 VPWR.n112 VPWR.t1171 161.106
R10256 VPWR.n167 VPWR.t1189 161.106
R10257 VPWR.n155 VPWR.t1317 161.106
R10258 VPWR.n117 VPWR.t1450 161.106
R10259 VPWR.n133 VPWR.t1090 161.106
R10260 VPWR.n122 VPWR.t1329 161.106
R10261 VPWR.n2880 VPWR.t1434 161.106
R10262 VPWR.n2878 VPWR.t1403 161.106
R10263 VPWR.n2876 VPWR.t1109 161.106
R10264 VPWR.n2874 VPWR.t1224 161.106
R10265 VPWR.n2872 VPWR.t1442 161.106
R10266 VPWR.n2870 VPWR.t1291 161.106
R10267 VPWR.n2868 VPWR.t1408 161.106
R10268 VPWR.n2866 VPWR.t1125 161.106
R10269 VPWR.n2864 VPWR.t1232 161.106
R10270 VPWR.n2862 VPWR.t1192 161.106
R10271 VPWR.n2860 VPWR.t1297 161.106
R10272 VPWR.n2858 VPWR.t1117 161.106
R10273 VPWR.n2856 VPWR.t1304 161.106
R10274 VPWR.n2854 VPWR.t1418 161.106
R10275 VPWR.n2852 VPWR.t1264 161.106
R10276 VPWR.n2850 VPWR.t1387 161.106
R10277 VPWR.n1616 VPWR.t1245 159.978
R10278 VPWR.n1620 VPWR.t1112 159.978
R10279 VPWR.n1224 VPWR.t1384 159.978
R10280 VPWR.n1220 VPWR.t1356 159.978
R10281 VPWR.n1215 VPWR.t1215 159.978
R10282 VPWR.n1211 VPWR.t1093 159.978
R10283 VPWR.n1206 VPWR.t1345 159.978
R10284 VPWR.n1173 VPWR.t1323 159.978
R10285 VPWR.n1200 VPWR.t1218 159.978
R10286 VPWR.n1177 VPWR.t1447 159.978
R10287 VPWR.n1181 VPWR.t1320 159.978
R10288 VPWR.n1185 VPWR.t1184 159.978
R10289 VPWR.n1626 VPWR.t1286 159.978
R10290 VPWR.n925 VPWR.t1122 159.978
R10291 VPWR.n1706 VPWR.t1156 159.978
R10292 VPWR.n921 VPWR.t1267 159.978
R10293 VPWR.n1240 VPWR.t1087 159.978
R10294 VPWR.n1567 VPWR.t1376 159.978
R10295 VPWR.n1555 VPWR.t1342 159.978
R10296 VPWR.n1537 VPWR.t1101 159.978
R10297 VPWR.n1256 VPWR.t1080 159.978
R10298 VPWR.n1357 VPWR.t1337 159.978
R10299 VPWR.n1368 VPWR.t1207 159.978
R10300 VPWR.n1379 VPWR.t1181 159.978
R10301 VPWR.n1390 VPWR.t1362 159.978
R10302 VPWR.n1401 VPWR.t1312 159.978
R10303 VPWR.n1412 VPWR.t1153 159.978
R10304 VPWR.n1330 VPWR.t1141 159.978
R10305 VPWR.n1318 VPWR.t1423 159.978
R10306 VPWR.n1282 VPWR.t1261 159.978
R10307 VPWR.n1298 VPWR.t1159 159.978
R10308 VPWR.n1288 VPWR.t1397 159.978
R10309 VPWR.n288 VPWR.t1273 159.978
R10310 VPWR.n272 VPWR.t1394 159.978
R10311 VPWR.n266 VPWR.t1150 159.978
R10312 VPWR.n254 VPWR.t1258 159.978
R10313 VPWR.n238 VPWR.t1270 159.978
R10314 VPWR.n232 VPWR.t1426 159.978
R10315 VPWR.n220 VPWR.t1147 159.978
R10316 VPWR.n204 VPWR.t1307 159.978
R10317 VPWR.n198 VPWR.t1326 159.978
R10318 VPWR.n186 VPWR.t1453 159.978
R10319 VPWR.n170 VPWR.t1197 159.978
R10320 VPWR.n164 VPWR.t1227 159.978
R10321 VPWR.n152 VPWR.t1077 159.978
R10322 VPWR.n136 VPWR.t1096 159.978
R10323 VPWR.n130 VPWR.t1221 159.978
R10324 VPWR.n93 VPWR.t1128 159.978
R10325 VPWR.n1617 VPWR.n1616 152
R10326 VPWR.n1621 VPWR.n1620 152
R10327 VPWR.n1225 VPWR.n1224 152
R10328 VPWR.n1221 VPWR.n1220 152
R10329 VPWR.n1216 VPWR.n1215 152
R10330 VPWR.n1212 VPWR.n1211 152
R10331 VPWR.n1207 VPWR.n1206 152
R10332 VPWR.n1174 VPWR.n1173 152
R10333 VPWR.n1201 VPWR.n1200 152
R10334 VPWR.n1178 VPWR.n1177 152
R10335 VPWR.n1182 VPWR.n1181 152
R10336 VPWR.n1186 VPWR.n1185 152
R10337 VPWR.n1627 VPWR.n1626 152
R10338 VPWR.n926 VPWR.n925 152
R10339 VPWR.n1707 VPWR.n1706 152
R10340 VPWR.n922 VPWR.n921 152
R10341 VPWR.n3120 VPWR.t798 148.127
R10342 VPWR.n1434 VPWR.t1955 145.137
R10343 VPWR.n1418 VPWR.t2001 145.137
R10344 VPWR.n1424 VPWR.t2050 145.137
R10345 VPWR.n1439 VPWR.t1941 145.137
R10346 VPWR.n1444 VPWR.t2044 145.137
R10347 VPWR.n1449 VPWR.t1990 145.137
R10348 VPWR.n1454 VPWR.t1984 145.137
R10349 VPWR.n1459 VPWR.t2042 145.137
R10350 VPWR.n1468 VPWR.t2030 145.137
R10351 VPWR.n1463 VPWR.t1991 145.137
R10352 VPWR.n1598 VPWR.t1934 145.137
R10353 VPWR.n1607 VPWR.t2070 145.137
R10354 VPWR.n1602 VPWR.t1981 145.137
R10355 VPWR.n933 VPWR.t1973 145.137
R10356 VPWR.n1691 VPWR.t1958 145.137
R10357 VPWR.n1687 VPWR.t2018 145.137
R10358 VPWR.n1243 VPWR.t1942 145.137
R10359 VPWR.n1570 VPWR.t2024 145.137
R10360 VPWR.n1558 VPWR.t2038 145.137
R10361 VPWR.n1248 VPWR.t2045 145.137
R10362 VPWR.n1251 VPWR.t1993 145.137
R10363 VPWR.n1354 VPWR.t1998 145.137
R10364 VPWR.n1365 VPWR.t2055 145.137
R10365 VPWR.n1376 VPWR.t1950 145.137
R10366 VPWR.n1387 VPWR.t1964 145.137
R10367 VPWR.n1398 VPWR.t2047 145.137
R10368 VPWR.n1409 VPWR.t2054 145.137
R10369 VPWR.n1333 VPWR.t1967 145.137
R10370 VPWR.n1321 VPWR.t2005 145.137
R10371 VPWR.n1285 VPWR.t2019 145.137
R10372 VPWR.n1301 VPWR.t2068 145.137
R10373 VPWR.n1290 VPWR.t1974 145.137
R10374 VPWR.n285 VPWR.t2035 145.137
R10375 VPWR.n275 VPWR.t1988 145.137
R10376 VPWR.n263 VPWR.t1976 145.137
R10377 VPWR.n251 VPWR.t1935 145.137
R10378 VPWR.n241 VPWR.t2021 145.137
R10379 VPWR.n229 VPWR.t2013 145.137
R10380 VPWR.n217 VPWR.t1933 145.137
R10381 VPWR.n207 VPWR.t2062 145.137
R10382 VPWR.n195 VPWR.t2022 145.137
R10383 VPWR.n183 VPWR.t1966 145.137
R10384 VPWR.n173 VPWR.t1957 145.137
R10385 VPWR.n161 VPWR.t2012 145.137
R10386 VPWR.n149 VPWR.t2004 145.137
R10387 VPWR.n139 VPWR.t1995 145.137
R10388 VPWR.n95 VPWR.t1939 145.137
R10389 VPWR.n127 VPWR.t2053 145.137
R10390 VPWR.n1583 VPWR.t2039 145.038
R10391 VPWR.n1572 VPWR.t1982 145.038
R10392 VPWR.n1564 VPWR.t1994 145.038
R10393 VPWR.n1552 VPWR.t2041 145.038
R10394 VPWR.n1540 VPWR.t1944 145.038
R10395 VPWR.n1349 VPWR.t1952 145.038
R10396 VPWR.n1360 VPWR.t2008 145.038
R10397 VPWR.n1371 VPWR.t2048 145.038
R10398 VPWR.n1382 VPWR.t1954 145.038
R10399 VPWR.n1393 VPWR.t1969 145.038
R10400 VPWR.n1404 VPWR.t2007 145.038
R10401 VPWR.n1335 VPWR.t2064 145.038
R10402 VPWR.n1327 VPWR.t1960 145.038
R10403 VPWR.n1315 VPWR.t2015 145.038
R10404 VPWR.n1303 VPWR.t2023 145.038
R10405 VPWR.n1295 VPWR.t2072 145.038
R10406 VPWR.n91 VPWR.t2037 145.038
R10407 VPWR.n87 VPWR.t1992 145.038
R10408 VPWR.n269 VPWR.t1985 145.038
R10409 VPWR.n257 VPWR.t2073 145.038
R10410 VPWR.n102 VPWR.t2032 145.038
R10411 VPWR.n235 VPWR.t1977 145.038
R10412 VPWR.n223 VPWR.t1936 145.038
R10413 VPWR.n107 VPWR.t2065 145.038
R10414 VPWR.n201 VPWR.t2014 145.038
R10415 VPWR.n189 VPWR.t1978 145.038
R10416 VPWR.n112 VPWR.t2063 145.038
R10417 VPWR.n167 VPWR.t2057 145.038
R10418 VPWR.n155 VPWR.t2009 145.038
R10419 VPWR.n117 VPWR.t1959 145.038
R10420 VPWR.n133 VPWR.t1945 145.038
R10421 VPWR.n122 VPWR.t2006 145.038
R10422 VPWR.n2880 VPWR.t2058 145.038
R10423 VPWR.n2878 VPWR.t1968 145.038
R10424 VPWR.n2876 VPWR.t2071 145.038
R10425 VPWR.n2874 VPWR.t2031 145.038
R10426 VPWR.n2872 VPWR.t1951 145.038
R10427 VPWR.n2870 VPWR.t2056 145.038
R10428 VPWR.n2868 VPWR.t2074 145.038
R10429 VPWR.n2866 VPWR.t2033 145.038
R10430 VPWR.n2864 VPWR.t2027 145.038
R10431 VPWR.n2862 VPWR.t1948 145.038
R10432 VPWR.n2860 VPWR.t2002 145.038
R10433 VPWR.n2858 VPWR.t2069 145.038
R10434 VPWR.n2856 VPWR.t2000 145.038
R10435 VPWR.n2854 VPWR.t1961 145.038
R10436 VPWR.n2852 VPWR.t2026 145.038
R10437 VPWR.n2850 VPWR.t1975 145.038
R10438 VPWR.n1616 VPWR.t1972 143.911
R10439 VPWR.n1620 VPWR.t1980 143.911
R10440 VPWR.n1224 VPWR.t2025 143.911
R10441 VPWR.n1220 VPWR.t1932 143.911
R10442 VPWR.n1215 VPWR.t1943 143.911
R10443 VPWR.n1211 VPWR.t2028 143.911
R10444 VPWR.n1206 VPWR.t2040 143.911
R10445 VPWR.n1173 VPWR.t2046 143.911
R10446 VPWR.n1200 VPWR.t1987 143.911
R10447 VPWR.n1177 VPWR.t1999 143.911
R10448 VPWR.n1181 VPWR.t2049 143.911
R10449 VPWR.n1185 VPWR.t1953 143.911
R10450 VPWR.n1626 VPWR.t2060 143.911
R10451 VPWR.n925 VPWR.t2016 143.911
R10452 VPWR.n1706 VPWR.t1962 143.911
R10453 VPWR.n921 VPWR.t2066 143.911
R10454 VPWR.n1240 VPWR.t1989 143.911
R10455 VPWR.n1567 VPWR.t2029 143.911
R10456 VPWR.n1555 VPWR.t1940 143.911
R10457 VPWR.n1537 VPWR.t1983 143.911
R10458 VPWR.n1256 VPWR.t2036 143.911
R10459 VPWR.n1357 VPWR.t2043 143.911
R10460 VPWR.n1368 VPWR.t1946 143.911
R10461 VPWR.n1379 VPWR.t1997 143.911
R10462 VPWR.n1390 VPWR.t2010 143.911
R10463 VPWR.n1401 VPWR.t1949 143.911
R10464 VPWR.n1412 VPWR.t1963 143.911
R10465 VPWR.n1330 VPWR.t1970 143.911
R10466 VPWR.n1318 VPWR.t2052 143.911
R10467 VPWR.n1282 VPWR.t2067 143.911
R10468 VPWR.n1298 VPWR.t1971 143.911
R10469 VPWR.n1288 VPWR.t2017 143.911
R10470 VPWR.n288 VPWR.t1938 143.911
R10471 VPWR.n272 VPWR.t2034 143.911
R10472 VPWR.n266 VPWR.t2020 143.911
R10473 VPWR.n254 VPWR.t1937 143.911
R10474 VPWR.n238 VPWR.t1931 143.911
R10475 VPWR.n232 VPWR.t2061 143.911
R10476 VPWR.n220 VPWR.t1979 143.911
R10477 VPWR.n204 VPWR.t1965 143.911
R10478 VPWR.n198 VPWR.t2059 143.911
R10479 VPWR.n186 VPWR.t2011 143.911
R10480 VPWR.n170 VPWR.t2003 143.911
R10481 VPWR.n164 VPWR.t1947 143.911
R10482 VPWR.n152 VPWR.t2051 143.911
R10483 VPWR.n136 VPWR.t1996 143.911
R10484 VPWR.n130 VPWR.t1956 143.911
R10485 VPWR.n93 VPWR.t1986 143.911
R10486 VPWR.t692 VPWR.t918 140.989
R10487 VPWR.t234 VPWR.t335 140.989
R10488 VPWR.t394 VPWR.t234 140.989
R10489 VPWR.t352 VPWR.t394 140.989
R10490 VPWR.t52 VPWR.t352 140.989
R10491 VPWR.t46 VPWR.t52 140.989
R10492 VPWR.t38 VPWR.t46 140.989
R10493 VPWR.t40 VPWR.t38 140.989
R10494 VPWR.t629 VPWR.t36 140.989
R10495 VPWR.t1887 VPWR.t348 140.989
R10496 VPWR.t241 VPWR.t1887 140.989
R10497 VPWR.t1886 VPWR.t241 140.989
R10498 VPWR.t543 VPWR.t1886 140.989
R10499 VPWR.t553 VPWR.t543 140.989
R10500 VPWR.t545 VPWR.t553 140.989
R10501 VPWR.t547 VPWR.t545 140.989
R10502 VPWR.t280 VPWR.t395 140.989
R10503 VPWR.t401 VPWR.t280 140.989
R10504 VPWR.t332 VPWR.t401 140.989
R10505 VPWR.t140 VPWR.t332 140.989
R10506 VPWR.t138 VPWR.t140 140.989
R10507 VPWR.t144 VPWR.t138 140.989
R10508 VPWR.t132 VPWR.t144 140.989
R10509 VPWR.t477 VPWR.t402 140.989
R10510 VPWR.t336 VPWR.t289 140.989
R10511 VPWR.t281 VPWR.t336 140.989
R10512 VPWR.t391 VPWR.t281 140.989
R10513 VPWR.t48 VPWR.t391 140.989
R10514 VPWR.t42 VPWR.t48 140.989
R10515 VPWR.t50 VPWR.t42 140.989
R10516 VPWR.t44 VPWR.t50 140.989
R10517 VPWR.t346 VPWR.t239 140.989
R10518 VPWR.t261 VPWR.t346 140.989
R10519 VPWR.t286 VPWR.t261 140.989
R10520 VPWR.t539 VPWR.t286 140.989
R10521 VPWR.t549 VPWR.t539 140.989
R10522 VPWR.t541 VPWR.t549 140.989
R10523 VPWR.t551 VPWR.t541 140.989
R10524 VPWR.t350 VPWR.t237 140.989
R10525 VPWR.t405 VPWR.t350 140.989
R10526 VPWR.t235 VPWR.t405 140.989
R10527 VPWR.t142 VPWR.t235 140.989
R10528 VPWR.t146 VPWR.t142 140.989
R10529 VPWR.t134 VPWR.t146 140.989
R10530 VPWR.t136 VPWR.t134 140.989
R10531 VPWR VPWR.n1150 133.312
R10532 VPWR.n3069 VPWR 127.562
R10533 VPWR.n3049 VPWR 127.562
R10534 VPWR.n3030 VPWR 127.562
R10535 VPWR VPWR.t283 125.883
R10536 VPWR.n2994 VPWR 125.883
R10537 VPWR.t631 VPWR.t34 120.849
R10538 VPWR.t828 VPWR.t415 117.492
R10539 VPWR.t638 VPWR.t1873 117.492
R10540 VPWR.t1552 VPWR 115.814
R10541 VPWR VPWR.t40 114.135
R10542 VPWR VPWR.t547 114.135
R10543 VPWR VPWR.t132 114.135
R10544 VPWR.t706 VPWR 107.421
R10545 VPWR.n1038 VPWR.n1037 106.561
R10546 VPWR.n3070 VPWR.n3069 106.561
R10547 VPWR.n3050 VPWR.n3049 106.561
R10548 VPWR.n3031 VPWR.n3030 106.561
R10549 VPWR.n2995 VPWR.n2994 106.561
R10550 VPWR.n2957 VPWR.n2956 106.561
R10551 VPWR.n2920 VPWR.n2919 106.561
R10552 VPWR VPWR.t635 106.543
R10553 VPWR VPWR.n942 104.8
R10554 VPWR VPWR.n965 104.8
R10555 VPWR VPWR.n989 104.8
R10556 VPWR VPWR.n1074 104.8
R10557 VPWR VPWR.n1113 104.8
R10558 VPWR.n1151 VPWR 100.883
R10559 VPWR VPWR.t784 100.624
R10560 VPWR.n1619 VPWR.n1618 91.8492
R10561 VPWR.n1623 VPWR.n1622 91.8492
R10562 VPWR.n1227 VPWR.n1226 91.8492
R10563 VPWR.n1223 VPWR.n1222 91.8492
R10564 VPWR.n1218 VPWR.n1217 91.8492
R10565 VPWR.n1214 VPWR.n1213 91.8492
R10566 VPWR.n1209 VPWR.n1208 91.8492
R10567 VPWR.n1176 VPWR.n1175 91.8492
R10568 VPWR.n1203 VPWR.n1202 91.8492
R10569 VPWR.n1180 VPWR.n1179 91.8492
R10570 VPWR.n1184 VPWR.n1183 91.8492
R10571 VPWR.n1188 VPWR.n1187 91.8492
R10572 VPWR.n1629 VPWR.n1628 91.8492
R10573 VPWR.n928 VPWR.n927 91.8492
R10574 VPWR.n1709 VPWR.n1708 91.8492
R10575 VPWR.n924 VPWR.n923 91.8492
R10576 VPWR.t389 VPWR 88.7855
R10577 VPWR.n3125 VPWR.n3123 83.2005
R10578 VPWR.n33 VPWR.n31 83.2005
R10579 VPWR.n3126 VPWR.n24 82.4894
R10580 VPWR.n35 VPWR.n34 82.4894
R10581 VPWR.n3111 VPWR.n35 80.9417
R10582 VPWR.n3123 VPWR.n25 80.9417
R10583 VPWR.n3106 VPWR.n24 80.9417
R10584 VPWR.n3104 VPWR.n31 80.9417
R10585 VPWR.n943 VPWR 79.407
R10586 VPWR.n966 VPWR 79.407
R10587 VPWR.n990 VPWR 79.407
R10588 VPWR.n1075 VPWR 79.407
R10589 VPWR.n1114 VPWR 79.407
R10590 VPWR.t640 VPWR.t181 78.8874
R10591 VPWR.t953 VPWR.t786 70.4952
R10592 VPWR.t786 VPWR.t955 70.4952
R10593 VPWR.t955 VPWR.t1732 70.4952
R10594 VPWR.t1732 VPWR.t931 70.4952
R10595 VPWR.t931 VPWR.t696 70.4952
R10596 VPWR.t696 VPWR.t339 70.4952
R10597 VPWR.t339 VPWR.t692 70.4952
R10598 VPWR.t981 VPWR.t477 70.4952
R10599 VPWR.t1728 VPWR.t981 70.4952
R10600 VPWR.t242 VPWR.t1728 70.4952
R10601 VPWR.t1028 VPWR.t242 70.4952
R10602 VPWR.t977 VPWR.t1028 70.4952
R10603 VPWR.t28 VPWR.t977 70.4952
R10604 VPWR.t283 VPWR.t28 70.4952
R10605 VPWR VPWR.t953 68.8168
R10606 VPWR.t637 VPWR.t633 68.8168
R10607 VPWR.t181 VPWR.t1552 62.103
R10608 VPWR VPWR.t629 60.4245
R10609 VPWR.t633 VPWR.t959 52.0323
R10610 VPWR.t1799 VPWR 50.3539
R10611 VPWR VPWR.t637 50.3539
R10612 VPWR VPWR.t631 50.3539
R10613 VPWR.t289 VPWR 50.3539
R10614 VPWR.t239 VPWR 50.3539
R10615 VPWR.t237 VPWR 50.3539
R10616 VPWR.n3112 VPWR.n3110 37.0005
R10617 VPWR.n3110 VPWR.n3109 37.0005
R10618 VPWR.n3108 VPWR.n3107 37.0005
R10619 VPWR.n3109 VPWR.n3108 37.0005
R10620 VPWR.n3122 VPWR.n3121 37.0005
R10621 VPWR.n3121 VPWR.n3120 37.0005
R10622 VPWR.n3119 VPWR.n3118 37.0005
R10623 VPWR.n3120 VPWR.n3119 37.0005
R10624 VPWR.n32 VPWR.t223 34.7652
R10625 VPWR.n32 VPWR.t1032 34.7652
R10626 VPWR.n3124 VPWR.t882 34.7652
R10627 VPWR.n3124 VPWR.t834 34.7652
R10628 VPWR.n1618 VPWR.n1617 34.7473
R10629 VPWR.n1622 VPWR.n1621 34.7473
R10630 VPWR.n1226 VPWR.n1225 34.7473
R10631 VPWR.n1222 VPWR.n1221 34.7473
R10632 VPWR.n1217 VPWR.n1216 34.7473
R10633 VPWR.n1213 VPWR.n1212 34.7473
R10634 VPWR.n1208 VPWR.n1207 34.7473
R10635 VPWR.n1175 VPWR.n1174 34.7473
R10636 VPWR.n1202 VPWR.n1201 34.7473
R10637 VPWR.n1179 VPWR.n1178 34.7473
R10638 VPWR.n1183 VPWR.n1182 34.7473
R10639 VPWR.n1187 VPWR.n1186 34.7473
R10640 VPWR.n1628 VPWR.n1627 34.7473
R10641 VPWR.n927 VPWR.n926 34.7473
R10642 VPWR.n1708 VPWR.n1707 34.7473
R10643 VPWR.n923 VPWR.n922 34.7473
R10644 VPWR.n1007 VPWR.n1006 34.6358
R10645 VPWR.n1065 VPWR.n1049 34.6358
R10646 VPWR.n1070 VPWR.n1069 34.6358
R10647 VPWR.n1104 VPWR.n1088 34.6358
R10648 VPWR.n1109 VPWR.n1108 34.6358
R10649 VPWR.n1119 VPWR.n1085 34.6358
R10650 VPWR.n1141 VPWR.n1125 34.6358
R10651 VPWR.n1146 VPWR.n1145 34.6358
R10652 VPWR.n3044 VPWR.n3043 34.6358
R10653 VPWR.n3010 VPWR.n3002 34.6358
R10654 VPWR.n3017 VPWR.n3016 34.6358
R10655 VPWR.n2974 VPWR.n2965 34.6358
R10656 VPWR.n2977 VPWR.n2976 34.6358
R10657 VPWR.n2981 VPWR.n2980 34.6358
R10658 VPWR.n2937 VPWR.n2928 34.6358
R10659 VPWR.n2940 VPWR.n2939 34.6358
R10660 VPWR.n2944 VPWR.n2943 34.6358
R10661 VPWR.n2951 VPWR.n2950 34.6358
R10662 VPWR.n2904 VPWR.n2900 34.6358
R10663 VPWR.n2908 VPWR.n2892 34.6358
R10664 VPWR.n2911 VPWR.n2910 34.6358
R10665 VPWR.n1024 VPWR.n1023 32.0005
R10666 VPWR.n1061 VPWR.n1060 32.0005
R10667 VPWR.n1100 VPWR.n1099 32.0005
R10668 VPWR.n1137 VPWR.n1136 32.0005
R10669 VPWR.n3006 VPWR.n3005 30.8711
R10670 VPWR.n2970 VPWR.n2969 30.8711
R10671 VPWR.n2933 VPWR.n2932 30.8711
R10672 VPWR.n2899 VPWR.n2898 30.8711
R10673 VPWR.n1033 VPWR.n1032 28.2358
R10674 VPWR.n5 VPWR.t1735 26.5955
R10675 VPWR.n5 VPWR.t695 26.5955
R10676 VPWR.n4 VPWR.t785 26.5955
R10677 VPWR.n4 VPWR.t1731 26.5955
R10678 VPWR.n948 VPWR.t384 26.5955
R10679 VPWR.n948 VPWR.t383 26.5955
R10680 VPWR.n947 VPWR.t782 26.5955
R10681 VPWR.n947 VPWR.t151 26.5955
R10682 VPWR.n953 VPWR.t380 26.5955
R10683 VPWR.n953 VPWR.t385 26.5955
R10684 VPWR.n946 VPWR.t664 26.5955
R10685 VPWR.n946 VPWR.t781 26.5955
R10686 VPWR.n971 VPWR.t225 26.5955
R10687 VPWR.n971 VPWR.t226 26.5955
R10688 VPWR.n970 VPWR.t678 26.5955
R10689 VPWR.n970 VPWR.t676 26.5955
R10690 VPWR.n976 VPWR.t1461 26.5955
R10691 VPWR.n976 VPWR.t1463 26.5955
R10692 VPWR.n969 VPWR.t681 26.5955
R10693 VPWR.n969 VPWR.t679 26.5955
R10694 VPWR.n995 VPWR.t984 26.5955
R10695 VPWR.n995 VPWR.t991 26.5955
R10696 VPWR.n994 VPWR.t840 26.5955
R10697 VPWR.n994 VPWR.t839 26.5955
R10698 VPWR.n1000 VPWR.t988 26.5955
R10699 VPWR.n1000 VPWR.t985 26.5955
R10700 VPWR.n993 VPWR.t843 26.5955
R10701 VPWR.n993 VPWR.t841 26.5955
R10702 VPWR.n1022 VPWR.t921 26.5955
R10703 VPWR.n1022 VPWR.t923 26.5955
R10704 VPWR.n1015 VPWR.t693 26.5955
R10705 VPWR.n1015 VPWR.t919 26.5955
R10706 VPWR.n1029 VPWR.t1733 26.5955
R10707 VPWR.n1029 VPWR.t697 26.5955
R10708 VPWR.n1031 VPWR.t956 26.5955
R10709 VPWR.n1031 VPWR.t932 26.5955
R10710 VPWR.n1059 VPWR.t228 26.5955
R10711 VPWR.n1059 VPWR.t232 26.5955
R10712 VPWR.n1058 VPWR.t1759 26.5955
R10713 VPWR.n1058 VPWR.t342 26.5955
R10714 VPWR.n1052 VPWR.t387 26.5955
R10715 VPWR.n1052 VPWR.t1751 26.5955
R10716 VPWR.n1051 VPWR.t665 26.5955
R10717 VPWR.n1051 VPWR.t1872 26.5955
R10718 VPWR.n1067 VPWR.t382 26.5955
R10719 VPWR.n1067 VPWR.t381 26.5955
R10720 VPWR.n1066 VPWR.t153 26.5955
R10721 VPWR.n1066 VPWR.t780 26.5955
R10722 VPWR.n1098 VPWR.t1871 26.5955
R10723 VPWR.n1098 VPWR.t1761 26.5955
R10724 VPWR.n1097 VPWR.t231 26.5955
R10725 VPWR.n1097 VPWR.t930 26.5955
R10726 VPWR.n1091 VPWR.t1831 26.5955
R10727 VPWR.n1091 VPWR.t1869 26.5955
R10728 VPWR.n1090 VPWR.t682 26.5955
R10729 VPWR.n1090 VPWR.t1754 26.5955
R10730 VPWR.n1106 VPWR.t1830 26.5955
R10731 VPWR.n1106 VPWR.t1832 26.5955
R10732 VPWR.n1105 VPWR.t683 26.5955
R10733 VPWR.n1105 VPWR.t680 26.5955
R10734 VPWR.n1135 VPWR.t952 26.5955
R10735 VPWR.n1135 VPWR.t1749 26.5955
R10736 VPWR.n1134 VPWR.t1760 26.5955
R10737 VPWR.n1134 VPWR.t344 26.5955
R10738 VPWR.n1128 VPWR.t987 26.5955
R10739 VPWR.n1128 VPWR.t949 26.5955
R10740 VPWR.n1127 VPWR.t837 26.5955
R10741 VPWR.n1127 VPWR.t1758 26.5955
R10742 VPWR.n1143 VPWR.t990 26.5955
R10743 VPWR.n1143 VPWR.t989 26.5955
R10744 VPWR.n1142 VPWR.t838 26.5955
R10745 VPWR.n1142 VPWR.t836 26.5955
R10746 VPWR.n3091 VPWR.t1924 26.5955
R10747 VPWR.n3091 VPWR.t968 26.5955
R10748 VPWR.n3093 VPWR.t1031 26.5955
R10749 VPWR.n3093 VPWR.t149 26.5955
R10750 VPWR.n3071 VPWR.t53 26.5955
R10751 VPWR.n3071 VPWR.t47 26.5955
R10752 VPWR.n3072 VPWR.t379 26.5955
R10753 VPWR.n3072 VPWR.t376 26.5955
R10754 VPWR.n3075 VPWR.t39 26.5955
R10755 VPWR.n3075 VPWR.t41 26.5955
R10756 VPWR.n3076 VPWR.t372 26.5955
R10757 VPWR.n3076 VPWR.t373 26.5955
R10758 VPWR.n3051 VPWR.t544 26.5955
R10759 VPWR.n3051 VPWR.t554 26.5955
R10760 VPWR.n3052 VPWR.t853 26.5955
R10761 VPWR.n3052 VPWR.t859 26.5955
R10762 VPWR.n3055 VPWR.t546 26.5955
R10763 VPWR.n3055 VPWR.t548 26.5955
R10764 VPWR.n3056 VPWR.t855 26.5955
R10765 VPWR.n3056 VPWR.t857 26.5955
R10766 VPWR.n3032 VPWR.t647 26.5955
R10767 VPWR.n3032 VPWR.t644 26.5955
R10768 VPWR.n3033 VPWR.t141 26.5955
R10769 VPWR.n3033 VPWR.t139 26.5955
R10770 VPWR.n3036 VPWR.t648 26.5955
R10771 VPWR.n3036 VPWR.t649 26.5955
R10772 VPWR.n3037 VPWR.t145 26.5955
R10773 VPWR.n3037 VPWR.t133 26.5955
R10774 VPWR.n2997 VPWR.t243 26.5955
R10775 VPWR.n2997 VPWR.t978 26.5955
R10776 VPWR.n3001 VPWR.t403 26.5955
R10777 VPWR.n3001 VPWR.t478 26.5955
R10778 VPWR.n3004 VPWR.t334 26.5955
R10779 VPWR.n3004 VPWR.t1889 26.5955
R10780 VPWR.n2998 VPWR.t1729 26.5955
R10781 VPWR.n2998 VPWR.t1029 26.5955
R10782 VPWR.n2968 VPWR.t337 26.5955
R10783 VPWR.n2968 VPWR.t1890 26.5955
R10784 VPWR.n2967 VPWR.t349 26.5955
R10785 VPWR.n2967 VPWR.t282 26.5955
R10786 VPWR.n2964 VPWR.t404 26.5955
R10787 VPWR.n2964 VPWR.t377 26.5955
R10788 VPWR.n2963 VPWR.t392 26.5955
R10789 VPWR.n2963 VPWR.t49 26.5955
R10790 VPWR.n2960 VPWR.t374 26.5955
R10791 VPWR.n2960 VPWR.t378 26.5955
R10792 VPWR.n2959 VPWR.t43 26.5955
R10793 VPWR.n2959 VPWR.t51 26.5955
R10794 VPWR.n2931 VPWR.t347 26.5955
R10795 VPWR.n2931 VPWR.t262 26.5955
R10796 VPWR.n2930 VPWR.t396 26.5955
R10797 VPWR.n2930 VPWR.t353 26.5955
R10798 VPWR.n2927 VPWR.t388 26.5955
R10799 VPWR.n2927 VPWR.t858 26.5955
R10800 VPWR.n2926 VPWR.t287 26.5955
R10801 VPWR.n2926 VPWR.t540 26.5955
R10802 VPWR.n2923 VPWR.t854 26.5955
R10803 VPWR.n2923 VPWR.t860 26.5955
R10804 VPWR.n2922 VPWR.t550 26.5955
R10805 VPWR.n2922 VPWR.t542 26.5955
R10806 VPWR.n2895 VPWR.t351 26.5955
R10807 VPWR.n2895 VPWR.t406 26.5955
R10808 VPWR.n2894 VPWR.t1885 26.5955
R10809 VPWR.n2894 VPWR.t979 26.5955
R10810 VPWR.n2902 VPWR.t400 26.5955
R10811 VPWR.n2902 VPWR.t143 26.5955
R10812 VPWR.n2901 VPWR.t236 26.5955
R10813 VPWR.n2901 VPWR.t645 26.5955
R10814 VPWR.n2891 VPWR.t147 26.5955
R10815 VPWR.n2891 VPWR.t135 26.5955
R10816 VPWR.n2890 VPWR.t642 26.5955
R10817 VPWR.n2890 VPWR.t646 26.5955
R10818 VPWR.n17 VPWR.n16 25.977
R10819 VPWR.n961 VPWR.n960 25.977
R10820 VPWR.n1021 VPWR.n1018 25.977
R10821 VPWR.n1057 VPWR.n1054 25.977
R10822 VPWR.n1080 VPWR.n1046 25.977
R10823 VPWR.n1096 VPWR.n1093 25.977
R10824 VPWR.n1133 VPWR.n1130 25.977
R10825 VPWR.n3100 VPWR.n3099 25.977
R10826 VPWR.n3084 VPWR.n3083 25.977
R10827 VPWR.n3006 VPWR.n3003 25.977
R10828 VPWR.n2970 VPWR.n2966 25.977
R10829 VPWR.n2988 VPWR.n2987 25.977
R10830 VPWR.n2933 VPWR.n2929 25.977
R10831 VPWR.n2898 VPWR.n2896 25.977
R10832 VPWR.n1043 VPWR.n1042 25.224
R10833 VPWR.n3026 VPWR.n3025 25.224
R10834 VPWR.n3011 VPWR.n3010 24.8476
R10835 VPWR.n2975 VPWR.n2974 24.8476
R10836 VPWR.n2938 VPWR.n2937 24.8476
R10837 VPWR.n2904 VPWR.n2903 24.8476
R10838 VPWR.n16 VPWR.n15 24.4711
R10839 VPWR.n960 VPWR.n959 24.4711
R10840 VPWR.n1023 VPWR.n1021 24.4711
R10841 VPWR.n1060 VPWR.n1057 24.4711
R10842 VPWR.n1099 VPWR.n1096 24.4711
R10843 VPWR.n1136 VPWR.n1133 24.4711
R10844 VPWR.n3099 VPWR.n3098 24.4711
R10845 VPWR.n3083 VPWR.n3082 24.4711
R10846 VPWR.n11 VPWR.n2 23.7181
R10847 VPWR.n955 VPWR.n944 23.7181
R10848 VPWR.n978 VPWR.n967 23.7181
R10849 VPWR.n982 VPWR.n967 23.7181
R10850 VPWR.n1002 VPWR.n991 23.7181
R10851 VPWR.n1006 VPWR.n991 23.7181
R10852 VPWR.n1038 VPWR.n1036 23.7181
R10853 VPWR.n1076 VPWR.n1073 23.7181
R10854 VPWR.n1115 VPWR.n1112 23.7181
R10855 VPWR.n1115 VPWR.n1085 23.7181
R10856 VPWR.n1152 VPWR.n1149 23.7181
R10857 VPWR.n3097 VPWR.n3096 23.7181
R10858 VPWR.n3078 VPWR.n3070 23.7181
R10859 VPWR.n3058 VPWR.n3050 23.7181
R10860 VPWR.n3062 VPWR.n3050 23.7181
R10861 VPWR.n3039 VPWR.n3031 23.7181
R10862 VPWR.n3043 VPWR.n3031 23.7181
R10863 VPWR.n3020 VPWR.n2995 23.7181
R10864 VPWR.n2983 VPWR.n2957 23.7181
R10865 VPWR.n2946 VPWR.n2920 23.7181
R10866 VPWR.n2950 VPWR.n2920 23.7181
R10867 VPWR.n2915 VPWR.n2914 23.7181
R10868 VPWR.t417 VPWR.t828 23.4987
R10869 VPWR.t1875 VPWR.t638 23.4987
R10870 VPWR.n11 VPWR.n10 22.9652
R10871 VPWR.n955 VPWR.n954 22.9652
R10872 VPWR.n978 VPWR.n977 22.9652
R10873 VPWR.n1002 VPWR.n1001 22.9652
R10874 VPWR.n3096 VPWR.n3092 22.9652
R10875 VPWR.n3078 VPWR.n3077 22.9652
R10876 VPWR.n3058 VPWR.n3057 22.9652
R10877 VPWR.n3039 VPWR.n3038 22.9652
R10878 VPWR.n1028 VPWR.n1016 22.2123
R10879 VPWR.n3013 VPWR.n3012 22.2123
R10880 VPWR.n10 VPWR.n3 21.4593
R10881 VPWR.n954 VPWR.n945 21.4593
R10882 VPWR.n977 VPWR.n968 21.4593
R10883 VPWR.n1001 VPWR.n992 21.4593
R10884 VPWR.n1150 VPWR.t343 20.5957
R10885 VPWR.n1151 VPWR.t916 20.5957
R10886 VPWR.n985 VPWR.n984 19.9534
R10887 VPWR.n1008 VPWR.n1007 19.9534
R10888 VPWR.n1042 VPWR.n1011 19.9534
R10889 VPWR.n3065 VPWR.n3064 19.9534
R10890 VPWR.n3045 VPWR.n3044 19.9534
R10891 VPWR.n3025 VPWR.n3024 19.9534
R10892 VPWR.n3013 VPWR.n2999 18.824
R10893 VPWR.n2977 VPWR.n2961 18.824
R10894 VPWR.n2940 VPWR.n2924 18.824
R10895 VPWR.n2909 VPWR.n2908 18.824
R10896 VPWR.n1024 VPWR.n1016 18.4476
R10897 VPWR.n1061 VPWR.n1053 18.4476
R10898 VPWR.n1081 VPWR.n1080 18.4476
R10899 VPWR.n1100 VPWR.n1092 18.4476
R10900 VPWR.n1137 VPWR.n1129 18.4476
R10901 VPWR.n2989 VPWR.n2988 18.4476
R10902 VPWR.n1121 VPWR.n1120 17.5829
R10903 VPWR.n2953 VPWR.n2952 17.5829
R10904 VPWR.n6 VPWR.n3 16.9417
R10905 VPWR.n949 VPWR.n945 16.9417
R10906 VPWR.n972 VPWR.n968 16.9417
R10907 VPWR.n996 VPWR.n992 16.9417
R10908 VPWR.n3019 VPWR.n3018 16.5652
R10909 VPWR.n1014 VPWR.n1012 16.1887
R10910 VPWR.n1082 VPWR.n1081 16.1887
R10911 VPWR.n2990 VPWR.n2989 16.1887
R10912 VPWR.n943 VPWR.t64 16.0935
R10913 VPWR.n966 VPWR.t224 16.0935
R10914 VPWR.n990 VPWR.t66 16.0935
R10915 VPWR.n1075 VPWR.t227 16.0935
R10916 VPWR.n1114 VPWR.t778 16.0935
R10917 VPWR.n942 VPWR.t150 16.0935
R10918 VPWR.n965 VPWR.t557 16.0935
R10919 VPWR.n989 VPWR.t559 16.0935
R10920 VPWR.n1074 VPWR.t152 16.0935
R10921 VPWR.n1113 VPWR.t230 16.0935
R10922 VPWR.n1033 VPWR.n1014 15.8123
R10923 VPWR.n3016 VPWR.n2999 15.8123
R10924 VPWR.n3018 VPWR.n3017 15.8123
R10925 VPWR.n2980 VPWR.n2961 15.8123
R10926 VPWR.n2943 VPWR.n2924 15.8123
R10927 VPWR.n2910 VPWR.n2909 15.8123
R10928 VPWR.n1038 VPWR.n1011 13.5534
R10929 VPWR.n3024 VPWR.n2995 13.5534
R10930 VPWR.n15 VPWR.n2 12.8005
R10931 VPWR.n959 VPWR.n944 12.8005
R10932 VPWR.n1076 VPWR.n1046 12.8005
R10933 VPWR.n3098 VPWR.n3097 12.8005
R10934 VPWR.n3082 VPWR.n3070 12.8005
R10935 VPWR.n2987 VPWR.n2957 12.8005
R10936 VPWR.n1030 VPWR.n1028 12.424
R10937 VPWR.n1068 VPWR.n1065 12.424
R10938 VPWR.n1107 VPWR.n1104 12.424
R10939 VPWR.n1144 VPWR.n1141 12.424
R10940 VPWR.n984 VPWR.n983 10.5417
R10941 VPWR.n1120 VPWR.n1119 10.5417
R10942 VPWR.n3064 VPWR.n3063 10.5417
R10943 VPWR.n2952 VPWR.n2951 10.5417
R10944 VPWR.n2976 VPWR.n2975 9.78874
R10945 VPWR.n2939 VPWR.n2938 9.78874
R10946 VPWR.n2903 VPWR.n2892 9.78874
R10947 VPWR.n1069 VPWR.n1068 9.41227
R10948 VPWR.n1073 VPWR.n1047 9.41227
R10949 VPWR.n1108 VPWR.n1107 9.41227
R10950 VPWR.n1112 VPWR.n1086 9.41227
R10951 VPWR.n1145 VPWR.n1144 9.41227
R10952 VPWR.n1149 VPWR.n1123 9.41227
R10953 VPWR.n2983 VPWR.n2982 9.41227
R10954 VPWR.n2946 VPWR.n2945 9.41227
R10955 VPWR.n2914 VPWR.n2888 9.41227
R10956 VPWR.n1617 VPWR 9.37021
R10957 VPWR.n1621 VPWR 9.37021
R10958 VPWR.n1225 VPWR 9.37021
R10959 VPWR.n1221 VPWR 9.37021
R10960 VPWR.n1216 VPWR 9.37021
R10961 VPWR.n1212 VPWR 9.37021
R10962 VPWR.n1207 VPWR 9.37021
R10963 VPWR.n1174 VPWR 9.37021
R10964 VPWR.n1201 VPWR 9.37021
R10965 VPWR.n1178 VPWR 9.37021
R10966 VPWR.n1182 VPWR 9.37021
R10967 VPWR.n1186 VPWR 9.37021
R10968 VPWR.n1627 VPWR 9.37021
R10969 VPWR.n926 VPWR 9.37021
R10970 VPWR.n1707 VPWR 9.37021
R10971 VPWR.n922 VPWR 9.37021
R10972 VPWR.n3003 VPWR 9.32394
R10973 VPWR.n2966 VPWR 9.32394
R10974 VPWR.n2929 VPWR 9.32394
R10975 VPWR VPWR.n2896 9.32394
R10976 VPWR.n499 VPWR.n490 9.30691
R10977 VPWR.n2422 VPWR.n487 9.30691
R10978 VPWR.n508 VPWR.n507 9.30691
R10979 VPWR.n699 VPWR.n685 9.30691
R10980 VPWR.n683 VPWR.n629 9.30691
R10981 VPWR.n627 VPWR.n626 9.30691
R10982 VPWR.n2074 VPWR.n2073 9.30691
R10983 VPWR.n1925 VPWR.n1924 9.30691
R10984 VPWR.n793 VPWR.n767 9.30691
R10985 VPWR.n801 VPWR.n800 9.30691
R10986 VPWR.n2554 VPWR.n2553 9.30691
R10987 VPWR.n1779 VPWR.n1778 9.30691
R10988 VPWR.n2735 VPWR.n373 9.30691
R10989 VPWR.n879 VPWR.n873 9.30691
R10990 VPWR.n1190 VPWR.n1189 9.30691
R10991 VPWR.n368 VPWR.n292 9.30691
R10992 VPWR.n18 VPWR.n17 9.3005
R10993 VPWR.n15 VPWR.n14 9.3005
R10994 VPWR.n13 VPWR.n2 9.3005
R10995 VPWR.n10 VPWR.n9 9.3005
R10996 VPWR.n8 VPWR.n3 9.3005
R10997 VPWR.n12 VPWR.n11 9.3005
R10998 VPWR.n16 VPWR.n0 9.3005
R10999 VPWR.n962 VPWR.n961 9.3005
R11000 VPWR.n959 VPWR.n958 9.3005
R11001 VPWR.n957 VPWR.n944 9.3005
R11002 VPWR.n954 VPWR.n952 9.3005
R11003 VPWR.n951 VPWR.n945 9.3005
R11004 VPWR.n956 VPWR.n955 9.3005
R11005 VPWR.n960 VPWR.n941 9.3005
R11006 VPWR.n986 VPWR.n985 9.3005
R11007 VPWR.n980 VPWR.n967 9.3005
R11008 VPWR.n977 VPWR.n975 9.3005
R11009 VPWR.n974 VPWR.n968 9.3005
R11010 VPWR.n979 VPWR.n978 9.3005
R11011 VPWR.n982 VPWR.n981 9.3005
R11012 VPWR.n984 VPWR.n964 9.3005
R11013 VPWR.n1009 VPWR.n1008 9.3005
R11014 VPWR.n1004 VPWR.n991 9.3005
R11015 VPWR.n1001 VPWR.n999 9.3005
R11016 VPWR.n998 VPWR.n992 9.3005
R11017 VPWR.n1003 VPWR.n1002 9.3005
R11018 VPWR.n1006 VPWR.n1005 9.3005
R11019 VPWR.n1007 VPWR.n988 9.3005
R11020 VPWR.n1040 VPWR.n1011 9.3005
R11021 VPWR.n1039 VPWR.n1038 9.3005
R11022 VPWR.n1019 VPWR.n1018 9.3005
R11023 VPWR.n1021 VPWR.n1020 9.3005
R11024 VPWR.n1023 VPWR.n1017 9.3005
R11025 VPWR.n1025 VPWR.n1024 9.3005
R11026 VPWR.n1026 VPWR.n1016 9.3005
R11027 VPWR.n1028 VPWR.n1027 9.3005
R11028 VPWR.n1032 VPWR.n1013 9.3005
R11029 VPWR.n1034 VPWR.n1033 9.3005
R11030 VPWR.n1036 VPWR.n1035 9.3005
R11031 VPWR.n1042 VPWR.n1041 9.3005
R11032 VPWR.n1044 VPWR.n1043 9.3005
R11033 VPWR.n1083 VPWR.n1082 9.3005
R11034 VPWR.n1078 VPWR.n1046 9.3005
R11035 VPWR.n1077 VPWR.n1076 9.3005
R11036 VPWR.n1055 VPWR.n1054 9.3005
R11037 VPWR.n1057 VPWR.n1056 9.3005
R11038 VPWR.n1060 VPWR.n1050 9.3005
R11039 VPWR.n1062 VPWR.n1061 9.3005
R11040 VPWR.n1063 VPWR.n1049 9.3005
R11041 VPWR.n1065 VPWR.n1064 9.3005
R11042 VPWR.n1069 VPWR.n1048 9.3005
R11043 VPWR.n1071 VPWR.n1070 9.3005
R11044 VPWR.n1073 VPWR.n1072 9.3005
R11045 VPWR.n1080 VPWR.n1079 9.3005
R11046 VPWR.n1116 VPWR.n1115 9.3005
R11047 VPWR.n1094 VPWR.n1093 9.3005
R11048 VPWR.n1096 VPWR.n1095 9.3005
R11049 VPWR.n1099 VPWR.n1089 9.3005
R11050 VPWR.n1101 VPWR.n1100 9.3005
R11051 VPWR.n1102 VPWR.n1088 9.3005
R11052 VPWR.n1104 VPWR.n1103 9.3005
R11053 VPWR.n1108 VPWR.n1087 9.3005
R11054 VPWR.n1110 VPWR.n1109 9.3005
R11055 VPWR.n1112 VPWR.n1111 9.3005
R11056 VPWR.n1117 VPWR.n1085 9.3005
R11057 VPWR.n1119 VPWR.n1118 9.3005
R11058 VPWR.n1153 VPWR.n1152 9.3005
R11059 VPWR.n1131 VPWR.n1130 9.3005
R11060 VPWR.n1133 VPWR.n1132 9.3005
R11061 VPWR.n1136 VPWR.n1126 9.3005
R11062 VPWR.n1138 VPWR.n1137 9.3005
R11063 VPWR.n1139 VPWR.n1125 9.3005
R11064 VPWR.n1141 VPWR.n1140 9.3005
R11065 VPWR.n1145 VPWR.n1124 9.3005
R11066 VPWR.n1147 VPWR.n1146 9.3005
R11067 VPWR.n1149 VPWR.n1148 9.3005
R11068 VPWR.n3096 VPWR.n3095 9.3005
R11069 VPWR.n3097 VPWR.n3089 9.3005
R11070 VPWR.n3098 VPWR.n3088 9.3005
R11071 VPWR.n3099 VPWR.n3087 9.3005
R11072 VPWR.n3101 VPWR.n3100 9.3005
R11073 VPWR.n3085 VPWR.n3084 9.3005
R11074 VPWR.n3079 VPWR.n3078 9.3005
R11075 VPWR.n3080 VPWR.n3070 9.3005
R11076 VPWR.n3082 VPWR.n3081 9.3005
R11077 VPWR.n3083 VPWR.n3068 9.3005
R11078 VPWR.n3066 VPWR.n3065 9.3005
R11079 VPWR.n3064 VPWR.n3048 9.3005
R11080 VPWR.n3059 VPWR.n3058 9.3005
R11081 VPWR.n3060 VPWR.n3050 9.3005
R11082 VPWR.n3062 VPWR.n3061 9.3005
R11083 VPWR.n3046 VPWR.n3045 9.3005
R11084 VPWR.n3040 VPWR.n3039 9.3005
R11085 VPWR.n3041 VPWR.n3031 9.3005
R11086 VPWR.n3043 VPWR.n3042 9.3005
R11087 VPWR.n3044 VPWR.n3029 9.3005
R11088 VPWR.n3027 VPWR.n3026 9.3005
R11089 VPWR.n3007 VPWR.n3006 9.3005
R11090 VPWR.n3008 VPWR.n3002 9.3005
R11091 VPWR.n3010 VPWR.n3009 9.3005
R11092 VPWR.n3012 VPWR.n3000 9.3005
R11093 VPWR.n3014 VPWR.n3013 9.3005
R11094 VPWR.n3016 VPWR.n3015 9.3005
R11095 VPWR.n3017 VPWR.n2996 9.3005
R11096 VPWR.n3021 VPWR.n3020 9.3005
R11097 VPWR.n3022 VPWR.n2995 9.3005
R11098 VPWR.n3024 VPWR.n3023 9.3005
R11099 VPWR.n3025 VPWR.n2993 9.3005
R11100 VPWR.n2991 VPWR.n2990 9.3005
R11101 VPWR.n2971 VPWR.n2970 9.3005
R11102 VPWR.n2972 VPWR.n2965 9.3005
R11103 VPWR.n2974 VPWR.n2973 9.3005
R11104 VPWR.n2976 VPWR.n2962 9.3005
R11105 VPWR.n2978 VPWR.n2977 9.3005
R11106 VPWR.n2980 VPWR.n2979 9.3005
R11107 VPWR.n2981 VPWR.n2958 9.3005
R11108 VPWR.n2984 VPWR.n2983 9.3005
R11109 VPWR.n2985 VPWR.n2957 9.3005
R11110 VPWR.n2987 VPWR.n2986 9.3005
R11111 VPWR.n2988 VPWR.n2955 9.3005
R11112 VPWR.n2934 VPWR.n2933 9.3005
R11113 VPWR.n2935 VPWR.n2928 9.3005
R11114 VPWR.n2937 VPWR.n2936 9.3005
R11115 VPWR.n2939 VPWR.n2925 9.3005
R11116 VPWR.n2941 VPWR.n2940 9.3005
R11117 VPWR.n2943 VPWR.n2942 9.3005
R11118 VPWR.n2944 VPWR.n2921 9.3005
R11119 VPWR.n2947 VPWR.n2946 9.3005
R11120 VPWR.n2948 VPWR.n2920 9.3005
R11121 VPWR.n2950 VPWR.n2949 9.3005
R11122 VPWR.n2951 VPWR.n2918 9.3005
R11123 VPWR.n2916 VPWR.n2915 9.3005
R11124 VPWR.n2898 VPWR.n2897 9.3005
R11125 VPWR.n2900 VPWR.n2893 9.3005
R11126 VPWR.n2905 VPWR.n2904 9.3005
R11127 VPWR.n2906 VPWR.n2892 9.3005
R11128 VPWR.n2908 VPWR.n2907 9.3005
R11129 VPWR.n2910 VPWR.n2889 9.3005
R11130 VPWR.n2912 VPWR.n2911 9.3005
R11131 VPWR.n2914 VPWR.n2913 9.3005
R11132 VPWR.n498 VPWR.n497 9.3005
R11133 VPWR.n494 VPWR.n453 9.3005
R11134 VPWR.n2543 VPWR.n2542 9.3005
R11135 VPWR.n2539 VPWR.n2538 9.3005
R11136 VPWR.n2536 VPWR.n2535 9.3005
R11137 VPWR.n2532 VPWR.n2531 9.3005
R11138 VPWR.n2512 VPWR.n2511 9.3005
R11139 VPWR.n2663 VPWR.n2662 9.3005
R11140 VPWR.n2660 VPWR.n420 9.3005
R11141 VPWR.n2657 VPWR.n2656 9.3005
R11142 VPWR.n2649 VPWR.n2648 9.3005
R11143 VPWR.n2645 VPWR.n2644 9.3005
R11144 VPWR.n2519 VPWR.n2518 9.3005
R11145 VPWR.n2523 VPWR.n2522 9.3005
R11146 VPWR.n2515 VPWR.n462 9.3005
R11147 VPWR.n2425 VPWR.n2424 9.3005
R11148 VPWR.n2429 VPWR.n2428 9.3005
R11149 VPWR.n2432 VPWR.n2431 9.3005
R11150 VPWR.n2435 VPWR.n480 9.3005
R11151 VPWR.n2444 VPWR.n2443 9.3005
R11152 VPWR.n2440 VPWR.n2439 9.3005
R11153 VPWR.n2463 VPWR.n2462 9.3005
R11154 VPWR.n2494 VPWR.n2493 9.3005
R11155 VPWR.n2491 VPWR.n2490 9.3005
R11156 VPWR.n2487 VPWR.n2486 9.3005
R11157 VPWR.n2483 VPWR.n2482 9.3005
R11158 VPWR.n2479 VPWR.n2478 9.3005
R11159 VPWR.n2475 VPWR.n2474 9.3005
R11160 VPWR.n2470 VPWR.n2469 9.3005
R11161 VPWR.n2467 VPWR.n2466 9.3005
R11162 VPWR.n511 VPWR.n503 9.3005
R11163 VPWR.n2409 VPWR.n2408 9.3005
R11164 VPWR.n2405 VPWR.n2404 9.3005
R11165 VPWR.n2402 VPWR.n2401 9.3005
R11166 VPWR.n2398 VPWR.n2397 9.3005
R11167 VPWR.n2395 VPWR.n2394 9.3005
R11168 VPWR.n2391 VPWR.n2390 9.3005
R11169 VPWR.n538 VPWR.n537 9.3005
R11170 VPWR.n2365 VPWR.n2364 9.3005
R11171 VPWR.n2369 VPWR.n2368 9.3005
R11172 VPWR.n532 VPWR.n528 9.3005
R11173 VPWR.n2377 VPWR.n2376 9.3005
R11174 VPWR.n2381 VPWR.n2380 9.3005
R11175 VPWR.n2384 VPWR.n2383 9.3005
R11176 VPWR.n2388 VPWR.n2387 9.3005
R11177 VPWR.n698 VPWR.n697 9.3005
R11178 VPWR.n694 VPWR.n693 9.3005
R11179 VPWR.n690 VPWR.n563 9.3005
R11180 VPWR.n2290 VPWR.n2289 9.3005
R11181 VPWR.n2286 VPWR.n2285 9.3005
R11182 VPWR.n573 VPWR.n572 9.3005
R11183 VPWR.n569 VPWR.n556 9.3005
R11184 VPWR.n2354 VPWR.n2353 9.3005
R11185 VPWR.n2351 VPWR.n2350 9.3005
R11186 VPWR.n2319 VPWR.n544 9.3005
R11187 VPWR.n2323 VPWR.n2322 9.3005
R11188 VPWR.n2326 VPWR.n2325 9.3005
R11189 VPWR.n2330 VPWR.n2329 9.3005
R11190 VPWR.n2313 VPWR.n553 9.3005
R11191 VPWR.n2310 VPWR.n2309 9.3005
R11192 VPWR.n682 VPWR.n681 9.3005
R11193 VPWR.n678 VPWR.n677 9.3005
R11194 VPWR.n675 VPWR.n674 9.3005
R11195 VPWR.n671 VPWR.n670 9.3005
R11196 VPWR.n667 VPWR.n666 9.3005
R11197 VPWR.n664 VPWR.n663 9.3005
R11198 VPWR.n660 VPWR.n659 9.3005
R11199 VPWR.n2258 VPWR.n2257 9.3005
R11200 VPWR.n2261 VPWR.n2260 9.3005
R11201 VPWR.n2264 VPWR.n2263 9.3005
R11202 VPWR.n2268 VPWR.n2267 9.3005
R11203 VPWR.n646 VPWR.n578 9.3005
R11204 VPWR.n650 VPWR.n649 9.3005
R11205 VPWR.n653 VPWR.n652 9.3005
R11206 VPWR.n657 VPWR.n656 9.3005
R11207 VPWR.n2138 VPWR.n2137 9.3005
R11208 VPWR.n2145 VPWR.n2144 9.3005
R11209 VPWR.n2141 VPWR.n616 9.3005
R11210 VPWR.n2155 VPWR.n2154 9.3005
R11211 VPWR.n2159 VPWR.n2158 9.3005
R11212 VPWR.n2167 VPWR.n2166 9.3005
R11213 VPWR.n2171 VPWR.n2170 9.3005
R11214 VPWR.n2238 VPWR.n2237 9.3005
R11215 VPWR.n2241 VPWR.n2240 9.3005
R11216 VPWR.n2187 VPWR.n586 9.3005
R11217 VPWR.n2191 VPWR.n2190 9.3005
R11218 VPWR.n2194 VPWR.n2193 9.3005
R11219 VPWR.n2198 VPWR.n2197 9.3005
R11220 VPWR.n2182 VPWR.n605 9.3005
R11221 VPWR.n2179 VPWR.n2178 9.3005
R11222 VPWR.n2077 VPWR.n2076 9.3005
R11223 VPWR.n2081 VPWR.n2080 9.3005
R11224 VPWR.n2085 VPWR.n2084 9.3005
R11225 VPWR.n2088 VPWR.n2065 9.3005
R11226 VPWR.n2116 VPWR.n2115 9.3005
R11227 VPWR.n2112 VPWR.n2111 9.3005
R11228 VPWR.n2109 VPWR.n2108 9.3005
R11229 VPWR.n2227 VPWR.n2226 9.3005
R11230 VPWR.n2224 VPWR.n594 9.3005
R11231 VPWR.n2221 VPWR.n2220 9.3005
R11232 VPWR.n2217 VPWR.n2216 9.3005
R11233 VPWR.n2213 VPWR.n2212 9.3005
R11234 VPWR.n2098 VPWR.n2097 9.3005
R11235 VPWR.n2102 VPWR.n2101 9.3005
R11236 VPWR.n2105 VPWR.n2104 9.3005
R11237 VPWR.n1932 VPWR.n1931 9.3005
R11238 VPWR.n1935 VPWR.n761 9.3005
R11239 VPWR.n1946 VPWR.n1945 9.3005
R11240 VPWR.n1942 VPWR.n1941 9.3005
R11241 VPWR.n1938 VPWR.n712 9.3005
R11242 VPWR.n2059 VPWR.n2058 9.3005
R11243 VPWR.n2055 VPWR.n2054 9.3005
R11244 VPWR.n2025 VPWR.n2024 9.3005
R11245 VPWR.n2028 VPWR.n2027 9.3005
R11246 VPWR.n734 VPWR.n730 9.3005
R11247 VPWR.n2036 VPWR.n2035 9.3005
R11248 VPWR.n2040 VPWR.n2039 9.3005
R11249 VPWR.n2043 VPWR.n2042 9.3005
R11250 VPWR.n2047 VPWR.n2046 9.3005
R11251 VPWR.n722 VPWR.n718 9.3005
R11252 VPWR.n792 VPWR.n791 9.3005
R11253 VPWR.n788 VPWR.n787 9.3005
R11254 VPWR.n785 VPWR.n784 9.3005
R11255 VPWR.n781 VPWR.n780 9.3005
R11256 VPWR.n778 VPWR.n777 9.3005
R11257 VPWR.n1962 VPWR.n1961 9.3005
R11258 VPWR.n1966 VPWR.n1965 9.3005
R11259 VPWR.n1995 VPWR.n1994 9.3005
R11260 VPWR.n1998 VPWR.n1997 9.3005
R11261 VPWR.n2001 VPWR.n2000 9.3005
R11262 VPWR.n2005 VPWR.n2004 9.3005
R11263 VPWR.n1989 VPWR.n744 9.3005
R11264 VPWR.n1986 VPWR.n1985 9.3005
R11265 VPWR.n1974 VPWR.n1973 9.3005
R11266 VPWR.n1970 VPWR.n1969 9.3005
R11267 VPWR.n804 VPWR.n796 9.3005
R11268 VPWR.n1911 VPWR.n1910 9.3005
R11269 VPWR.n1907 VPWR.n1906 9.3005
R11270 VPWR.n1904 VPWR.n1903 9.3005
R11271 VPWR.n1900 VPWR.n1899 9.3005
R11272 VPWR.n818 VPWR.n817 9.3005
R11273 VPWR.n821 VPWR.n812 9.3005
R11274 VPWR.n834 VPWR.n833 9.3005
R11275 VPWR.n837 VPWR.n836 9.3005
R11276 VPWR.n1873 VPWR.n1872 9.3005
R11277 VPWR.n1877 VPWR.n1876 9.3005
R11278 VPWR.n1880 VPWR.n1879 9.3005
R11279 VPWR.n1884 VPWR.n1883 9.3005
R11280 VPWR.n1887 VPWR.n1886 9.3005
R11281 VPWR.n1891 VPWR.n1890 9.3005
R11282 VPWR.n2557 VPWR.n2549 9.3005
R11283 VPWR.n2566 VPWR.n2565 9.3005
R11284 VPWR.n2562 VPWR.n2561 9.3005
R11285 VPWR.n2580 VPWR.n2579 9.3005
R11286 VPWR.n2584 VPWR.n2583 9.3005
R11287 VPWR.n2603 VPWR.n2602 9.3005
R11288 VPWR.n2606 VPWR.n2605 9.3005
R11289 VPWR.n2609 VPWR.n2608 9.3005
R11290 VPWR.n2613 VPWR.n2612 9.3005
R11291 VPWR.n2616 VPWR.n2615 9.3005
R11292 VPWR.n2620 VPWR.n2619 9.3005
R11293 VPWR.n2623 VPWR.n2622 9.3005
R11294 VPWR.n2627 VPWR.n2626 9.3005
R11295 VPWR.n2591 VPWR.n440 9.3005
R11296 VPWR.n2588 VPWR.n2587 9.3005
R11297 VPWR.n1783 VPWR.n1782 9.3005
R11298 VPWR.n1786 VPWR.n1785 9.3005
R11299 VPWR.n1789 VPWR.n867 9.3005
R11300 VPWR.n1801 VPWR.n1800 9.3005
R11301 VPWR.n1797 VPWR.n1796 9.3005
R11302 VPWR.n1792 VPWR.n860 9.3005
R11303 VPWR.n1821 VPWR.n1820 9.3005
R11304 VPWR.n1825 VPWR.n1824 9.3005
R11305 VPWR.n1833 VPWR.n1832 9.3005
R11306 VPWR.n1859 VPWR.n1858 9.3005
R11307 VPWR.n1856 VPWR.n1855 9.3005
R11308 VPWR.n1852 VPWR.n1851 9.3005
R11309 VPWR.n1848 VPWR.n1847 9.3005
R11310 VPWR.n1836 VPWR.n846 9.3005
R11311 VPWR.n1840 VPWR.n1839 9.3005
R11312 VPWR.n2734 VPWR.n2733 9.3005
R11313 VPWR.n2730 VPWR.n2729 9.3005
R11314 VPWR.n384 VPWR.n380 9.3005
R11315 VPWR.n2674 VPWR.n2673 9.3005
R11316 VPWR.n2682 VPWR.n2681 9.3005
R11317 VPWR.n2686 VPWR.n2685 9.3005
R11318 VPWR.n411 VPWR.n407 9.3005
R11319 VPWR.n2694 VPWR.n2693 9.3005
R11320 VPWR.n2698 VPWR.n2697 9.3005
R11321 VPWR.n402 VPWR.n398 9.3005
R11322 VPWR.n2706 VPWR.n2705 9.3005
R11323 VPWR.n2710 VPWR.n2709 9.3005
R11324 VPWR.n393 VPWR.n389 9.3005
R11325 VPWR.n2718 VPWR.n2717 9.3005
R11326 VPWR.n2722 VPWR.n2721 9.3005
R11327 VPWR.n882 VPWR.n875 9.3005
R11328 VPWR.n1769 VPWR.n1768 9.3005
R11329 VPWR.n1765 VPWR.n1764 9.3005
R11330 VPWR.n1762 VPWR.n1761 9.3005
R11331 VPWR.n1758 VPWR.n1757 9.3005
R11332 VPWR.n899 VPWR.n898 9.3005
R11333 VPWR.n902 VPWR.n893 9.3005
R11334 VPWR.n1749 VPWR.n1748 9.3005
R11335 VPWR.n1745 VPWR.n1744 9.3005
R11336 VPWR.n1742 VPWR.n1741 9.3005
R11337 VPWR.n1738 VPWR.n1737 9.3005
R11338 VPWR.n1723 VPWR.n1722 9.3005
R11339 VPWR.n1720 VPWR.n1716 9.3005
R11340 VPWR.n1731 VPWR.n1730 9.3005
R11341 VPWR.n1735 VPWR.n1734 9.3005
R11342 VPWR.n1194 VPWR.n1193 9.3005
R11343 VPWR.n1198 VPWR.n1197 9.3005
R11344 VPWR.n1204 VPWR.n1171 9.3005
R11345 VPWR.n1661 VPWR.n1660 9.3005
R11346 VPWR.n1657 VPWR.n1656 9.3005
R11347 VPWR.n1654 VPWR.n1653 9.3005
R11348 VPWR.n1650 VPWR.n1649 9.3005
R11349 VPWR.n1647 VPWR.n1646 9.3005
R11350 VPWR.n1643 VPWR.n1642 9.3005
R11351 VPWR.n1624 VPWR.n1232 9.3005
R11352 VPWR.n1634 VPWR.n1633 9.3005
R11353 VPWR.n1630 VPWR.n929 9.3005
R11354 VPWR.n1713 VPWR.n1712 9.3005
R11355 VPWR.n1710 VPWR.n919 9.3005
R11356 VPWR.n1704 VPWR.n1703 9.3005
R11357 VPWR.n367 VPWR.n366 9.3005
R11358 VPWR.n318 VPWR.n317 9.3005
R11359 VPWR.n321 VPWR.n320 9.3005
R11360 VPWR.n325 VPWR.n324 9.3005
R11361 VPWR.n328 VPWR.n327 9.3005
R11362 VPWR.n332 VPWR.n331 9.3005
R11363 VPWR.n335 VPWR.n334 9.3005
R11364 VPWR.n339 VPWR.n338 9.3005
R11365 VPWR.n342 VPWR.n341 9.3005
R11366 VPWR.n346 VPWR.n345 9.3005
R11367 VPWR.n349 VPWR.n348 9.3005
R11368 VPWR.n353 VPWR.n352 9.3005
R11369 VPWR.n356 VPWR.n355 9.3005
R11370 VPWR.n360 VPWR.n359 9.3005
R11371 VPWR.n363 VPWR.n362 9.3005
R11372 VPWR.n1587 VPWR.n1586 9.3005
R11373 VPWR.n1590 VPWR.n1589 9.3005
R11374 VPWR.n1525 VPWR.n1235 9.3005
R11375 VPWR.n1530 VPWR.n1529 9.3005
R11376 VPWR.n1534 VPWR.n1533 9.3005
R11377 VPWR.n1522 VPWR.n1521 9.3005
R11378 VPWR.n1517 VPWR.n1516 9.3005
R11379 VPWR.n1513 VPWR.n1512 9.3005
R11380 VPWR.n1503 VPWR.n1502 9.3005
R11381 VPWR.n1499 VPWR.n1498 9.3005
R11382 VPWR.n1491 VPWR.n1490 9.3005
R11383 VPWR.n1487 VPWR.n1486 9.3005
R11384 VPWR.n1280 VPWR.n1279 9.3005
R11385 VPWR.n1670 VPWR.n1669 9.3005
R11386 VPWR.n1674 VPWR.n1673 9.3005
R11387 VPWR.n1162 VPWR.n1157 9.3005
R11388 VPWR.n2761 VPWR.n2760 9.3005
R11389 VPWR.n2765 VPWR.n2764 9.3005
R11390 VPWR.n2773 VPWR.n2772 9.3005
R11391 VPWR.n2777 VPWR.n2776 9.3005
R11392 VPWR.n2785 VPWR.n2784 9.3005
R11393 VPWR.n2789 VPWR.n2788 9.3005
R11394 VPWR.n2797 VPWR.n2796 9.3005
R11395 VPWR.n2801 VPWR.n2800 9.3005
R11396 VPWR.n2809 VPWR.n2808 9.3005
R11397 VPWR.n2813 VPWR.n2812 9.3005
R11398 VPWR.n2821 VPWR.n2820 9.3005
R11399 VPWR.n2825 VPWR.n2824 9.3005
R11400 VPWR.n2833 VPWR.n2832 9.3005
R11401 VPWR.n2837 VPWR.n2836 9.3005
R11402 VPWR.n2845 VPWR.n2844 9.3005
R11403 VPWR.n2848 VPWR.n2847 9.3005
R11404 VPWR.n3111 VPWR.n30 8.40959
R11405 VPWR.n3105 VPWR.n30 8.40959
R11406 VPWR.n28 VPWR.n25 8.40959
R11407 VPWR.n3105 VPWR.n28 8.40959
R11408 VPWR.n3106 VPWR.n27 8.40959
R11409 VPWR.n3105 VPWR.n27 8.40959
R11410 VPWR.n3104 VPWR.n29 8.40959
R11411 VPWR.n3105 VPWR.n29 8.40959
R11412 VPWR.n983 VPWR.n982 8.28285
R11413 VPWR.n3063 VPWR.n3062 8.28285
R11414 VPWR.n1309 VPWR.n1287 8.25914
R11415 VPWR.n1579 VPWR.n1578 8.25914
R11416 VPWR.n282 VPWR.n100 8.25914
R11417 VPWR.n145 VPWR.n121 8.25914
R11418 VPWR.n2853 VPWR.n2851 7.96303
R11419 VPWR.n1690 VPWR.n1689 7.91351
R11420 VPWR.n1437 VPWR.n1436 7.9105
R11421 VPWR.n1421 VPWR.n1420 7.9105
R11422 VPWR.n1427 VPWR.n1426 7.9105
R11423 VPWR.n1442 VPWR.n1441 7.9105
R11424 VPWR.n1447 VPWR.n1446 7.9105
R11425 VPWR.n1452 VPWR.n1451 7.9105
R11426 VPWR.n1457 VPWR.n1456 7.9105
R11427 VPWR.n1462 VPWR.n1461 7.9105
R11428 VPWR.n1471 VPWR.n1470 7.9105
R11429 VPWR.n1466 VPWR.n1465 7.9105
R11430 VPWR.n1601 VPWR.n1600 7.9105
R11431 VPWR.n1610 VPWR.n1609 7.9105
R11432 VPWR.n1605 VPWR.n1604 7.9105
R11433 VPWR.n936 VPWR.n935 7.9105
R11434 VPWR.n1694 VPWR.n1693 7.9105
R11435 VPWR.n1309 VPWR.n1308 7.9105
R11436 VPWR.n1311 VPWR.n1310 7.9105
R11437 VPWR.n1323 VPWR.n1276 7.9105
R11438 VPWR.n1341 VPWR.n1340 7.9105
R11439 VPWR.n1342 VPWR.n1272 7.9105
R11440 VPWR.n1343 VPWR.n1273 7.9105
R11441 VPWR.n1344 VPWR.n1274 7.9105
R11442 VPWR.n1345 VPWR.n1275 7.9105
R11443 VPWR.n1347 VPWR.n1346 7.9105
R11444 VPWR.n1348 VPWR.n1250 7.9105
R11445 VPWR.n1546 VPWR.n1545 7.9105
R11446 VPWR.n1548 VPWR.n1547 7.9105
R11447 VPWR.n1560 VPWR.n1245 7.9105
R11448 VPWR.n1578 VPWR.n1577 7.9105
R11449 VPWR.n145 VPWR.n144 7.9105
R11450 VPWR.n147 VPWR.n146 7.9105
R11451 VPWR.n159 VPWR.n116 7.9105
R11452 VPWR.n179 VPWR.n178 7.9105
R11453 VPWR.n181 VPWR.n180 7.9105
R11454 VPWR.n193 VPWR.n111 7.9105
R11455 VPWR.n213 VPWR.n212 7.9105
R11456 VPWR.n215 VPWR.n214 7.9105
R11457 VPWR.n227 VPWR.n106 7.9105
R11458 VPWR.n247 VPWR.n246 7.9105
R11459 VPWR.n249 VPWR.n248 7.9105
R11460 VPWR.n261 VPWR.n101 7.9105
R11461 VPWR.n281 VPWR.n280 7.9105
R11462 VPWR.n283 VPWR.n282 7.9105
R11463 VPWR.n7 VPWR.n6 7.56315
R11464 VPWR.n950 VPWR.n949 7.56315
R11465 VPWR.n973 VPWR.n972 7.56315
R11466 VPWR.n997 VPWR.n996 7.56315
R11467 VPWR.n3114 VPWR.n3113 7.0697
R11468 VPWR.n3130 VPWR.n3129 6.57193
R11469 VPWR.n3094 VPWR.n3092 6.4511
R11470 VPWR.n3077 VPWR.n3074 6.4511
R11471 VPWR.n3057 VPWR.n3054 6.4511
R11472 VPWR.n3038 VPWR.n3035 6.4511
R11473 VPWR.n1070 VPWR.n1047 6.4005
R11474 VPWR.n1109 VPWR.n1086 6.4005
R11475 VPWR.n1146 VPWR.n1123 6.4005
R11476 VPWR.n3012 VPWR.n3011 6.4005
R11477 VPWR.n2982 VPWR.n2981 6.4005
R11478 VPWR.n2945 VPWR.n2944 6.4005
R11479 VPWR.n2911 VPWR.n2888 6.4005
R11480 VPWR.n1633 VPWR.n1619 6.04494
R11481 VPWR.n1624 VPWR.n1623 6.04494
R11482 VPWR.n1643 VPWR.n1227 6.04494
R11483 VPWR.n1646 VPWR.n1223 6.04494
R11484 VPWR.n1650 VPWR.n1218 6.04494
R11485 VPWR.n1653 VPWR.n1214 6.04494
R11486 VPWR.n1657 VPWR.n1209 6.04494
R11487 VPWR.n1660 VPWR.n1176 6.04494
R11488 VPWR.n1741 VPWR.n906 6.04494
R11489 VPWR.n1745 VPWR.n904 6.04494
R11490 VPWR.n1748 VPWR.n895 6.04494
R11491 VPWR.n902 VPWR.n901 6.04494
R11492 VPWR.n899 VPWR.n896 6.04494
R11493 VPWR.n1758 VPWR.n887 6.04494
R11494 VPWR.n1824 VPWR.n858 6.04494
R11495 VPWR.n1821 VPWR.n859 6.04494
R11496 VPWR.n2532 VPWR.n459 6.04494
R11497 VPWR.n2535 VPWR.n458 6.04494
R11498 VPWR.n2539 VPWR.n456 6.04494
R11499 VPWR.n2542 VPWR.n455 6.04494
R11500 VPWR.n494 VPWR.n493 6.04494
R11501 VPWR.n497 VPWR.n491 6.04494
R11502 VPWR.n490 VPWR.n489 6.04494
R11503 VPWR.n2512 VPWR.n2509 6.04494
R11504 VPWR.n2515 VPWR.n2514 6.04494
R11505 VPWR.n2522 VPWR.n2508 6.04494
R11506 VPWR.n2519 VPWR.n2517 6.04494
R11507 VPWR.n2645 VPWR.n430 6.04494
R11508 VPWR.n2648 VPWR.n429 6.04494
R11509 VPWR.n2657 VPWR.n423 6.04494
R11510 VPWR.n2660 VPWR.n2659 6.04494
R11511 VPWR.n2662 VPWR.n422 6.04494
R11512 VPWR.n2440 VPWR.n2437 6.04494
R11513 VPWR.n2443 VPWR.n481 6.04494
R11514 VPWR.n2435 VPWR.n2434 6.04494
R11515 VPWR.n2432 VPWR.n482 6.04494
R11516 VPWR.n2428 VPWR.n483 6.04494
R11517 VPWR.n2425 VPWR.n484 6.04494
R11518 VPWR.n487 VPWR.n485 6.04494
R11519 VPWR.n2463 VPWR.n473 6.04494
R11520 VPWR.n2466 VPWR.n472 6.04494
R11521 VPWR.n2470 VPWR.n471 6.04494
R11522 VPWR.n2475 VPWR.n2472 6.04494
R11523 VPWR.n2478 VPWR.n470 6.04494
R11524 VPWR.n2483 VPWR.n469 6.04494
R11525 VPWR.n2486 VPWR.n468 6.04494
R11526 VPWR.n2491 VPWR.n467 6.04494
R11527 VPWR.n2493 VPWR.n466 6.04494
R11528 VPWR.n2394 VPWR.n518 6.04494
R11529 VPWR.n2398 VPWR.n516 6.04494
R11530 VPWR.n2401 VPWR.n515 6.04494
R11531 VPWR.n2405 VPWR.n513 6.04494
R11532 VPWR.n2408 VPWR.n505 6.04494
R11533 VPWR.n511 VPWR.n510 6.04494
R11534 VPWR.n508 VPWR.n506 6.04494
R11535 VPWR.n2391 VPWR.n519 6.04494
R11536 VPWR.n2387 VPWR.n521 6.04494
R11537 VPWR.n2384 VPWR.n522 6.04494
R11538 VPWR.n2380 VPWR.n524 6.04494
R11539 VPWR.n2377 VPWR.n525 6.04494
R11540 VPWR.n532 VPWR.n531 6.04494
R11541 VPWR.n2368 VPWR.n530 6.04494
R11542 VPWR.n2365 VPWR.n534 6.04494
R11543 VPWR.n537 VPWR.n536 6.04494
R11544 VPWR.n572 VPWR.n567 6.04494
R11545 VPWR.n2286 VPWR.n566 6.04494
R11546 VPWR.n2289 VPWR.n565 6.04494
R11547 VPWR.n690 VPWR.n689 6.04494
R11548 VPWR.n694 VPWR.n692 6.04494
R11549 VPWR.n697 VPWR.n687 6.04494
R11550 VPWR.n685 VPWR.n684 6.04494
R11551 VPWR.n569 VPWR.n568 6.04494
R11552 VPWR.n2310 VPWR.n555 6.04494
R11553 VPWR.n2313 VPWR.n2312 6.04494
R11554 VPWR.n2329 VPWR.n554 6.04494
R11555 VPWR.n2326 VPWR.n2315 6.04494
R11556 VPWR.n2322 VPWR.n2317 6.04494
R11557 VPWR.n2319 VPWR.n2318 6.04494
R11558 VPWR.n2351 VPWR.n543 6.04494
R11559 VPWR.n2353 VPWR.n542 6.04494
R11560 VPWR.n663 VPWR.n638 6.04494
R11561 VPWR.n667 VPWR.n636 6.04494
R11562 VPWR.n671 VPWR.n669 6.04494
R11563 VPWR.n674 VPWR.n635 6.04494
R11564 VPWR.n678 VPWR.n633 6.04494
R11565 VPWR.n681 VPWR.n631 6.04494
R11566 VPWR.n629 VPWR.n628 6.04494
R11567 VPWR.n660 VPWR.n639 6.04494
R11568 VPWR.n656 VPWR.n641 6.04494
R11569 VPWR.n653 VPWR.n642 6.04494
R11570 VPWR.n649 VPWR.n644 6.04494
R11571 VPWR.n646 VPWR.n645 6.04494
R11572 VPWR.n2267 VPWR.n580 6.04494
R11573 VPWR.n2264 VPWR.n581 6.04494
R11574 VPWR.n2260 VPWR.n2254 6.04494
R11575 VPWR.n2258 VPWR.n2255 6.04494
R11576 VPWR.n2167 VPWR.n611 6.04494
R11577 VPWR.n2158 VPWR.n614 6.04494
R11578 VPWR.n2155 VPWR.n615 6.04494
R11579 VPWR.n2141 VPWR.n2140 6.04494
R11580 VPWR.n2144 VPWR.n619 6.04494
R11581 VPWR.n2138 VPWR.n620 6.04494
R11582 VPWR.n626 VPWR.n624 6.04494
R11583 VPWR.n2170 VPWR.n610 6.04494
R11584 VPWR.n2179 VPWR.n607 6.04494
R11585 VPWR.n2182 VPWR.n2181 6.04494
R11586 VPWR.n2197 VPWR.n606 6.04494
R11587 VPWR.n2194 VPWR.n2184 6.04494
R11588 VPWR.n2190 VPWR.n2185 6.04494
R11589 VPWR.n2187 VPWR.n2186 6.04494
R11590 VPWR.n2240 VPWR.n588 6.04494
R11591 VPWR.n2238 VPWR.n589 6.04494
R11592 VPWR.n2112 VPWR.n2090 6.04494
R11593 VPWR.n2115 VPWR.n2067 6.04494
R11594 VPWR.n2088 VPWR.n2087 6.04494
R11595 VPWR.n2085 VPWR.n2068 6.04494
R11596 VPWR.n2080 VPWR.n2069 6.04494
R11597 VPWR.n2077 VPWR.n2070 6.04494
R11598 VPWR.n2073 VPWR.n2071 6.04494
R11599 VPWR.n2108 VPWR.n2092 6.04494
R11600 VPWR.n2105 VPWR.n2093 6.04494
R11601 VPWR.n2101 VPWR.n2095 6.04494
R11602 VPWR.n2098 VPWR.n2096 6.04494
R11603 VPWR.n2213 VPWR.n599 6.04494
R11604 VPWR.n2216 VPWR.n598 6.04494
R11605 VPWR.n2221 VPWR.n597 6.04494
R11606 VPWR.n2224 VPWR.n2223 6.04494
R11607 VPWR.n2226 VPWR.n596 6.04494
R11608 VPWR.n2058 VPWR.n714 6.04494
R11609 VPWR.n1938 VPWR.n1937 6.04494
R11610 VPWR.n1942 VPWR.n1940 6.04494
R11611 VPWR.n1945 VPWR.n762 6.04494
R11612 VPWR.n1935 VPWR.n1934 6.04494
R11613 VPWR.n1932 VPWR.n763 6.04494
R11614 VPWR.n1924 VPWR.n1922 6.04494
R11615 VPWR.n2055 VPWR.n715 6.04494
R11616 VPWR.n722 VPWR.n721 6.04494
R11617 VPWR.n2046 VPWR.n720 6.04494
R11618 VPWR.n2043 VPWR.n724 6.04494
R11619 VPWR.n2039 VPWR.n726 6.04494
R11620 VPWR.n2036 VPWR.n727 6.04494
R11621 VPWR.n734 VPWR.n733 6.04494
R11622 VPWR.n2027 VPWR.n732 6.04494
R11623 VPWR.n2025 VPWR.n736 6.04494
R11624 VPWR.n1962 VPWR.n753 6.04494
R11625 VPWR.n777 VPWR.n775 6.04494
R11626 VPWR.n781 VPWR.n773 6.04494
R11627 VPWR.n784 VPWR.n772 6.04494
R11628 VPWR.n788 VPWR.n771 6.04494
R11629 VPWR.n791 VPWR.n769 6.04494
R11630 VPWR.n767 VPWR.n766 6.04494
R11631 VPWR.n1965 VPWR.n752 6.04494
R11632 VPWR.n1970 VPWR.n751 6.04494
R11633 VPWR.n1973 VPWR.n750 6.04494
R11634 VPWR.n1986 VPWR.n747 6.04494
R11635 VPWR.n1989 VPWR.n1988 6.04494
R11636 VPWR.n2004 VPWR.n746 6.04494
R11637 VPWR.n2001 VPWR.n1991 6.04494
R11638 VPWR.n1997 VPWR.n1992 6.04494
R11639 VPWR.n1995 VPWR.n1993 6.04494
R11640 VPWR.n818 VPWR.n815 6.04494
R11641 VPWR.n1900 VPWR.n809 6.04494
R11642 VPWR.n1903 VPWR.n808 6.04494
R11643 VPWR.n1907 VPWR.n806 6.04494
R11644 VPWR.n1910 VPWR.n798 6.04494
R11645 VPWR.n804 VPWR.n803 6.04494
R11646 VPWR.n801 VPWR.n799 6.04494
R11647 VPWR.n821 VPWR.n820 6.04494
R11648 VPWR.n1890 VPWR.n814 6.04494
R11649 VPWR.n1887 VPWR.n823 6.04494
R11650 VPWR.n1883 VPWR.n825 6.04494
R11651 VPWR.n1880 VPWR.n826 6.04494
R11652 VPWR.n1876 VPWR.n828 6.04494
R11653 VPWR.n1873 VPWR.n829 6.04494
R11654 VPWR.n836 VPWR.n830 6.04494
R11655 VPWR.n834 VPWR.n831 6.04494
R11656 VPWR.n2580 VPWR.n445 6.04494
R11657 VPWR.n2562 VPWR.n2559 6.04494
R11658 VPWR.n2565 VPWR.n2551 6.04494
R11659 VPWR.n2557 VPWR.n2556 6.04494
R11660 VPWR.n2554 VPWR.n2552 6.04494
R11661 VPWR.n2583 VPWR.n444 6.04494
R11662 VPWR.n2588 VPWR.n443 6.04494
R11663 VPWR.n2591 VPWR.n2590 6.04494
R11664 VPWR.n2626 VPWR.n442 6.04494
R11665 VPWR.n2623 VPWR.n2593 6.04494
R11666 VPWR.n2619 VPWR.n2594 6.04494
R11667 VPWR.n2616 VPWR.n2595 6.04494
R11668 VPWR.n2612 VPWR.n2597 6.04494
R11669 VPWR.n2609 VPWR.n2598 6.04494
R11670 VPWR.n2605 VPWR.n2600 6.04494
R11671 VPWR.n2603 VPWR.n2601 6.04494
R11672 VPWR.n1792 VPWR.n1791 6.04494
R11673 VPWR.n1797 VPWR.n1794 6.04494
R11674 VPWR.n1800 VPWR.n868 6.04494
R11675 VPWR.n1789 VPWR.n1788 6.04494
R11676 VPWR.n1786 VPWR.n869 6.04494
R11677 VPWR.n1782 VPWR.n870 6.04494
R11678 VPWR.n1779 VPWR.n871 6.04494
R11679 VPWR.n1833 VPWR.n850 6.04494
R11680 VPWR.n1839 VPWR.n849 6.04494
R11681 VPWR.n1836 VPWR.n1835 6.04494
R11682 VPWR.n1848 VPWR.n845 6.04494
R11683 VPWR.n1851 VPWR.n844 6.04494
R11684 VPWR.n1856 VPWR.n843 6.04494
R11685 VPWR.n1858 VPWR.n842 6.04494
R11686 VPWR.n2730 VPWR.n377 6.04494
R11687 VPWR.n2733 VPWR.n375 6.04494
R11688 VPWR.n373 VPWR.n372 6.04494
R11689 VPWR.n384 VPWR.n383 6.04494
R11690 VPWR.n2721 VPWR.n382 6.04494
R11691 VPWR.n2718 VPWR.n386 6.04494
R11692 VPWR.n393 VPWR.n392 6.04494
R11693 VPWR.n2709 VPWR.n391 6.04494
R11694 VPWR.n2706 VPWR.n395 6.04494
R11695 VPWR.n402 VPWR.n401 6.04494
R11696 VPWR.n2697 VPWR.n400 6.04494
R11697 VPWR.n2694 VPWR.n404 6.04494
R11698 VPWR.n411 VPWR.n410 6.04494
R11699 VPWR.n2685 VPWR.n409 6.04494
R11700 VPWR.n2682 VPWR.n413 6.04494
R11701 VPWR.n2673 VPWR.n2672 6.04494
R11702 VPWR.n1761 VPWR.n886 6.04494
R11703 VPWR.n1765 VPWR.n884 6.04494
R11704 VPWR.n1768 VPWR.n877 6.04494
R11705 VPWR.n882 VPWR.n881 6.04494
R11706 VPWR.n879 VPWR.n878 6.04494
R11707 VPWR.n1738 VPWR.n907 6.04494
R11708 VPWR.n1734 VPWR.n909 6.04494
R11709 VPWR.n1731 VPWR.n910 6.04494
R11710 VPWR.n1720 VPWR.n1719 6.04494
R11711 VPWR.n1722 VPWR.n1718 6.04494
R11712 VPWR.n1204 VPWR.n1203 6.04494
R11713 VPWR.n1198 VPWR.n1180 6.04494
R11714 VPWR.n1193 VPWR.n1184 6.04494
R11715 VPWR.n1190 VPWR.n1188 6.04494
R11716 VPWR.n1630 VPWR.n1629 6.04494
R11717 VPWR.n1704 VPWR.n928 6.04494
R11718 VPWR.n1710 VPWR.n1709 6.04494
R11719 VPWR.n1712 VPWR.n924 6.04494
R11720 VPWR.n292 VPWR.n291 6.04494
R11721 VPWR.n366 VPWR.n294 6.04494
R11722 VPWR.n363 VPWR.n296 6.04494
R11723 VPWR.n359 VPWR.n298 6.04494
R11724 VPWR.n356 VPWR.n299 6.04494
R11725 VPWR.n352 VPWR.n301 6.04494
R11726 VPWR.n349 VPWR.n302 6.04494
R11727 VPWR.n345 VPWR.n304 6.04494
R11728 VPWR.n342 VPWR.n305 6.04494
R11729 VPWR.n338 VPWR.n307 6.04494
R11730 VPWR.n335 VPWR.n308 6.04494
R11731 VPWR.n331 VPWR.n310 6.04494
R11732 VPWR.n328 VPWR.n311 6.04494
R11733 VPWR.n324 VPWR.n313 6.04494
R11734 VPWR.n321 VPWR.n314 6.04494
R11735 VPWR.n317 VPWR.n316 6.04494
R11736 VPWR.n1162 VPWR.n1161 6.04494
R11737 VPWR.n1673 VPWR.n1160 6.04494
R11738 VPWR.n1670 VPWR.n1164 6.04494
R11739 VPWR.n1279 VPWR.n1277 6.04494
R11740 VPWR.n1487 VPWR.n1271 6.04494
R11741 VPWR.n1490 VPWR.n1270 6.04494
R11742 VPWR.n1499 VPWR.n1266 6.04494
R11743 VPWR.n1502 VPWR.n1265 6.04494
R11744 VPWR.n1513 VPWR.n1261 6.04494
R11745 VPWR.n1516 VPWR.n1260 6.04494
R11746 VPWR.n1522 VPWR.n1254 6.04494
R11747 VPWR.n1533 VPWR.n1253 6.04494
R11748 VPWR.n1530 VPWR.n1527 6.04494
R11749 VPWR.n1525 VPWR.n1524 6.04494
R11750 VPWR.n1589 VPWR.n1238 6.04494
R11751 VPWR.n1587 VPWR.n1239 6.04494
R11752 VPWR.n2764 VPWR.n85 6.04494
R11753 VPWR.n2773 VPWR.n80 6.04494
R11754 VPWR.n2776 VPWR.n79 6.04494
R11755 VPWR.n2785 VPWR.n74 6.04494
R11756 VPWR.n2788 VPWR.n73 6.04494
R11757 VPWR.n2797 VPWR.n68 6.04494
R11758 VPWR.n2800 VPWR.n67 6.04494
R11759 VPWR.n2809 VPWR.n62 6.04494
R11760 VPWR.n2812 VPWR.n61 6.04494
R11761 VPWR.n2821 VPWR.n56 6.04494
R11762 VPWR.n2824 VPWR.n55 6.04494
R11763 VPWR.n2833 VPWR.n50 6.04494
R11764 VPWR.n2836 VPWR.n49 6.04494
R11765 VPWR.n2845 VPWR.n44 6.04494
R11766 VPWR.n2847 VPWR.n43 6.04494
R11767 VPWR.n2761 VPWR.n86 6.04494
R11768 VPWR.n3128 VPWR.n20 5.59663
R11769 VPWR.n3131 VPWR.n3130 5.59663
R11770 VPWR.n3129 VPWR.n22 5.59425
R11771 VPWR.n3115 VPWR.n3114 5.59425
R11772 VPWR.n3074 VPWR.n3073 5.39628
R11773 VPWR.n3054 VPWR.n3053 5.39628
R11774 VPWR.n3035 VPWR.n3034 5.39628
R11775 VPWR.n3114 VPWR.n23 4.9938
R11776 VPWR VPWR.n3103 4.94464
R11777 VPWR.n2881 VPWR 4.72593
R11778 VPWR.n2879 VPWR 4.72593
R11779 VPWR.n2877 VPWR 4.72593
R11780 VPWR.n2875 VPWR 4.72593
R11781 VPWR.n2873 VPWR 4.72593
R11782 VPWR.n2871 VPWR 4.72593
R11783 VPWR.n2869 VPWR 4.72593
R11784 VPWR.n2867 VPWR 4.72593
R11785 VPWR.n2865 VPWR 4.72593
R11786 VPWR.n2863 VPWR 4.72593
R11787 VPWR.n2861 VPWR 4.72593
R11788 VPWR.n2859 VPWR 4.72593
R11789 VPWR.n2857 VPWR 4.72593
R11790 VPWR.n2855 VPWR 4.72593
R11791 VPWR.n2853 VPWR 4.72593
R11792 VPWR.n36 VPWR.n26 4.6505
R11793 VPWR.n3117 VPWR.n3116 4.6505
R11794 VPWR.n34 VPWR.n23 4.6505
R11795 VPWR.n3127 VPWR.n3126 4.6505
R11796 VPWR.n3113 VPWR.n3112 4.6505
R11797 VPWR.n3107 VPWR.n21 4.6505
R11798 VPWR.n1154 VPWR.n1153 4.55954
R11799 VPWR.n3129 VPWR.n3128 4.5005
R11800 VPWR.n857 VPWR.n813 4.5005
R11801 VPWR.n1968 VPWR.n717 4.5005
R11802 VPWR.n2049 VPWR.n2048 4.5005
R11803 VPWR.n2103 VPWR.n608 4.5005
R11804 VPWR.n2177 VPWR.n2176 4.5005
R11805 VPWR.n640 VPWR.n550 4.5005
R11806 VPWR.n2335 VPWR.n551 4.5005
R11807 VPWR.n2336 VPWR.n520 4.5005
R11808 VPWR.n2468 VPWR.n461 4.5005
R11809 VPWR.n2525 VPWR.n2524 4.5005
R11810 VPWR.n2510 VPWR.n437 4.5005
R11811 VPWR.n2461 VPWR.n2460 4.5005
R11812 VPWR.n2389 VPWR.n474 4.5005
R11813 VPWR.n2308 VPWR.n2307 4.5005
R11814 VPWR.n658 VPWR.n557 4.5005
R11815 VPWR.n2173 VPWR.n2172 4.5005
R11816 VPWR.n2091 VPWR.n609 4.5005
R11817 VPWR.n2053 VPWR.n2052 4.5005
R11818 VPWR.n1967 VPWR.n716 4.5005
R11819 VPWR.n1893 VPWR.n1892 4.5005
R11820 VPWR.n1885 VPWR.n749 4.5005
R11821 VPWR.n1980 VPWR.n1975 4.5005
R11822 VPWR.n1979 VPWR.n719 4.5005
R11823 VPWR.n2094 VPWR.n604 4.5005
R11824 VPWR.n2200 VPWR.n2199 4.5005
R11825 VPWR.n651 VPWR.n552 4.5005
R11826 VPWR.n2332 VPWR.n2331 4.5005
R11827 VPWR.n2382 VPWR.n463 4.5005
R11828 VPWR.n2504 VPWR.n464 4.5005
R11829 VPWR.n2507 VPWR.n2506 4.5005
R11830 VPWR.n2621 VPWR.n397 4.5005
R11831 VPWR.n441 VPWR.n396 4.5005
R11832 VPWR.n2629 VPWR.n2628 4.5005
R11833 VPWR.n2586 VPWR.n388 4.5005
R11834 VPWR.n2530 VPWR.n2529 4.5005
R11835 VPWR.n2438 VPWR.n460 4.5005
R11836 VPWR.n2303 VPWR.n517 4.5005
R11837 VPWR.n2304 VPWR.n559 4.5005
R11838 VPWR.n637 VPWR.n558 4.5005
R11839 VPWR.n2165 VPWR.n2164 4.5005
R11840 VPWR.n2110 VPWR.n612 4.5005
R11841 VPWR.n756 VPWR.n713 4.5005
R11842 VPWR.n1960 VPWR.n1959 4.5005
R11843 VPWR.n816 VPWR.n754 4.5005
R11844 VPWR.n1818 VPWR.n1817 4.5005
R11845 VPWR.n1819 VPWR.n811 4.5005
R11846 VPWR.n1827 VPWR.n1826 4.5005
R11847 VPWR.n1831 VPWR.n1830 4.5005
R11848 VPWR.n1842 VPWR.n1841 4.5005
R11849 VPWR.n824 VPWR.n748 4.5005
R11850 VPWR.n1984 VPWR.n1983 4.5005
R11851 VPWR.n2041 VPWR.n601 4.5005
R11852 VPWR.n2205 VPWR.n602 4.5005
R11853 VPWR.n2204 VPWR.n603 4.5005
R11854 VPWR.n643 VPWR.n548 4.5005
R11855 VPWR.n2341 VPWR.n549 4.5005
R11856 VPWR.n2340 VPWR.n523 4.5005
R11857 VPWR.n2473 VPWR.n432 4.5005
R11858 VPWR.n2639 VPWR.n433 4.5005
R11859 VPWR.n2638 VPWR.n434 4.5005
R11860 VPWR.n2585 VPWR.n387 4.5005
R11861 VPWR.n2454 VPWR.n457 4.5005
R11862 VPWR.n2455 VPWR.n476 4.5005
R11863 VPWR.n2396 VPWR.n475 4.5005
R11864 VPWR.n2284 VPWR.n2283 4.5005
R11865 VPWR.n665 VPWR.n574 4.5005
R11866 VPWR.n2161 VPWR.n2160 4.5005
R11867 VPWR.n2066 VPWR.n613 4.5005
R11868 VPWR.n2061 VPWR.n2060 4.5005
R11869 VPWR.n774 VPWR.n711 4.5005
R11870 VPWR.n1898 VPWR.n1897 4.5005
R11871 VPWR.n1795 VPWR.n810 4.5005
R11872 VPWR.n1846 VPWR.n1845 4.5005
R11873 VPWR.n1878 VPWR.n743 4.5005
R11874 VPWR.n2007 VPWR.n2006 4.5005
R11875 VPWR.n725 VPWR.n600 4.5005
R11876 VPWR.n2211 VPWR.n2210 4.5005
R11877 VPWR.n2192 VPWR.n577 4.5005
R11878 VPWR.n2270 VPWR.n2269 4.5005
R11879 VPWR.n2324 VPWR.n526 4.5005
R11880 VPWR.n2375 VPWR.n2374 4.5005
R11881 VPWR.n2480 VPWR.n431 4.5005
R11882 VPWR.n2643 VPWR.n2642 4.5005
R11883 VPWR.n2614 VPWR.n405 4.5005
R11884 VPWR.n2692 VPWR.n2691 4.5005
R11885 VPWR.n436 VPWR.n399 4.5005
R11886 VPWR.n2700 VPWR.n2699 4.5005
R11887 VPWR.n2704 VPWR.n2703 4.5005
R11888 VPWR.n439 VPWR.n390 4.5005
R11889 VPWR.n2712 VPWR.n2711 4.5005
R11890 VPWR.n2716 VPWR.n2715 4.5005
R11891 VPWR.n448 VPWR.n381 4.5005
R11892 VPWR.n2578 VPWR.n2577 4.5005
R11893 VPWR.n2537 VPWR.n446 4.5005
R11894 VPWR.n2446 VPWR.n2445 4.5005
R11895 VPWR.n514 VPWR.n479 4.5005
R11896 VPWR.n2280 VPWR.n564 4.5005
R11897 VPWR.n2279 VPWR.n576 4.5005
R11898 VPWR.n2153 VPWR.n575 4.5005
R11899 VPWR.n2118 VPWR.n2117 4.5005
R11900 VPWR.n2064 VPWR.n710 4.5005
R11901 VPWR.n779 VPWR.n709 4.5005
R11902 VPWR.n1811 VPWR.n807 4.5005
R11903 VPWR.n1812 VPWR.n863 4.5005
R11904 VPWR.n885 VPWR.n862 4.5005
R11905 VPWR.n1756 VPWR.n1755 4.5005
R11906 VPWR.n897 VPWR.n861 4.5005
R11907 VPWR.n1751 VPWR.n1750 4.5005
R11908 VPWR.n894 VPWR.n852 4.5005
R11909 VPWR.n1743 VPWR.n851 4.5005
R11910 VPWR.n905 VPWR.n848 4.5005
R11911 VPWR.n1736 VPWR.n847 4.5005
R11912 VPWR.n908 VPWR.n839 4.5005
R11913 VPWR.n1866 VPWR.n840 4.5005
R11914 VPWR.n1867 VPWR.n827 4.5005
R11915 VPWR.n745 VPWR.n728 4.5005
R11916 VPWR.n2034 VPWR.n2033 4.5005
R11917 VPWR.n2218 VPWR.n583 4.5005
R11918 VPWR.n2246 VPWR.n584 4.5005
R11919 VPWR.n2247 VPWR.n579 4.5005
R11920 VPWR.n2316 VPWR.n527 4.5005
R11921 VPWR.n2371 VPWR.n2370 4.5005
R11922 VPWR.n2481 VPWR.n428 4.5005
R11923 VPWR.n2651 VPWR.n2650 4.5005
R11924 VPWR.n2596 VPWR.n406 4.5005
R11925 VPWR.n2688 VPWR.n2687 4.5005
R11926 VPWR.n2724 VPWR.n2723 4.5005
R11927 VPWR.n2560 VPWR.n379 4.5005
R11928 VPWR.n2450 VPWR.n454 4.5005
R11929 VPWR.n2449 VPWR.n478 4.5005
R11930 VPWR.n2403 VPWR.n477 4.5005
R11931 VPWR.n2292 VPWR.n2291 4.5005
R11932 VPWR.n634 VPWR.n562 4.5005
R11933 VPWR.n2152 VPWR.n2151 4.5005
R11934 VPWR.n2083 VPWR.n617 4.5005
R11935 VPWR.n1951 VPWR.n759 4.5005
R11936 VPWR.n1952 VPWR.n758 4.5005
R11937 VPWR.n1905 VPWR.n757 4.5005
R11938 VPWR.n1803 VPWR.n1802 4.5005
R11939 VPWR.n1763 VPWR.n866 4.5005
R11940 VPWR.n1663 VPWR.n1662 4.5005
R11941 VPWR.n1482 VPWR.n1172 4.5005
R11942 VPWR.n1655 VPWR.n888 4.5005
R11943 VPWR.n1268 VPWR.n1210 4.5005
R11944 VPWR.n1648 VPWR.n892 4.5005
R11945 VPWR.n1263 VPWR.n1219 4.5005
R11946 VPWR.n1641 VPWR.n1640 4.5005
R11947 VPWR.n1636 VPWR.n1635 4.5005
R11948 VPWR.n1615 VPWR.n1614 4.5005
R11949 VPWR.n1701 VPWR.n1700 4.5005
R11950 VPWR.n1702 VPWR.n911 4.5005
R11951 VPWR.n1729 VPWR.n1728 4.5005
R11952 VPWR.n1853 VPWR.n838 4.5005
R11953 VPWR.n1871 VPWR.n1870 4.5005
R11954 VPWR.n1999 VPWR.n729 4.5005
R11955 VPWR.n2030 VPWR.n2029 4.5005
R11956 VPWR.n2219 VPWR.n585 4.5005
R11957 VPWR.n2243 VPWR.n2242 4.5005
R11958 VPWR.n2262 VPWR.n545 4.5005
R11959 VPWR.n2348 VPWR.n2347 4.5005
R11960 VPWR.n547 VPWR.n529 4.5005
R11961 VPWR.n2488 VPWR.n424 4.5005
R11962 VPWR.n2655 VPWR.n2654 4.5005
R11963 VPWR.n2607 VPWR.n427 4.5005
R11964 VPWR.n426 VPWR.n408 4.5005
R11965 VPWR.n312 VPWR.n47 4.5005
R11966 VPWR.n326 VPWR.n52 4.5005
R11967 VPWR.n309 VPWR.n53 4.5005
R11968 VPWR.n333 VPWR.n58 4.5005
R11969 VPWR.n306 VPWR.n59 4.5005
R11970 VPWR.n340 VPWR.n64 4.5005
R11971 VPWR.n303 VPWR.n65 4.5005
R11972 VPWR.n347 VPWR.n70 4.5005
R11973 VPWR.n300 VPWR.n71 4.5005
R11974 VPWR.n354 VPWR.n76 4.5005
R11975 VPWR.n297 VPWR.n77 4.5005
R11976 VPWR.n361 VPWR.n82 4.5005
R11977 VPWR.n2728 VPWR.n2727 4.5005
R11978 VPWR.n2550 VPWR.n378 4.5005
R11979 VPWR.n2545 VPWR.n2544 4.5005
R11980 VPWR.n2430 VPWR.n452 4.5005
R11981 VPWR.n2296 VPWR.n504 4.5005
R11982 VPWR.n2295 VPWR.n561 4.5005
R11983 VPWR.n676 VPWR.n560 4.5005
R11984 VPWR.n2147 VPWR.n2146 4.5005
R11985 VPWR.n2082 VPWR.n618 4.5005
R11986 VPWR.n1948 VPWR.n1947 4.5005
R11987 VPWR.n786 VPWR.n760 4.5005
R11988 VPWR.n1807 VPWR.n797 4.5005
R11989 VPWR.n1806 VPWR.n865 4.5005
R11990 VPWR.n876 VPWR.n864 4.5005
R11991 VPWR.n1196 VPWR.n1166 4.5005
R11992 VPWR.n1195 VPWR.n874 4.5005
R11993 VPWR.n1771 VPWR.n1770 4.5005
R11994 VPWR.n1784 VPWR.n795 4.5005
R11995 VPWR.n1913 VPWR.n1912 4.5005
R11996 VPWR.n768 VPWR.n764 4.5005
R11997 VPWR.n1930 VPWR.n1929 4.5005
R11998 VPWR.n2075 VPWR.n621 4.5005
R11999 VPWR.n2136 VPWR.n2135 4.5005
R12000 VPWR.n630 VPWR.n622 4.5005
R12001 VPWR.n686 VPWR.n502 4.5005
R12002 VPWR.n2411 VPWR.n2410 4.5005
R12003 VPWR.n2423 VPWR.n450 4.5005
R12004 VPWR.n2548 VPWR.n451 4.5005
R12005 VPWR.n2570 VPWR.n2567 4.5005
R12006 VPWR.n2569 VPWR.n374 4.5005
R12007 VPWR.n293 VPWR.n83 4.5005
R12008 VPWR.n319 VPWR.n46 4.5005
R12009 VPWR.n2680 VPWR.n2679 4.5005
R12010 VPWR.n2599 VPWR.n414 4.5005
R12011 VPWR.n2665 VPWR.n2664 4.5005
R12012 VPWR.n2489 VPWR.n419 4.5005
R12013 VPWR.n2363 VPWR.n2362 4.5005
R12014 VPWR.n2349 VPWR.n539 4.5005
R12015 VPWR.n2253 VPWR.n2252 4.5005
R12016 VPWR.n587 VPWR.n582 4.5005
R12017 VPWR.n2229 VPWR.n2228 4.5005
R12018 VPWR.n731 VPWR.n593 4.5005
R12019 VPWR.n2012 VPWR.n742 4.5005
R12020 VPWR.n2013 VPWR.n741 4.5005
R12021 VPWR.n1854 VPWR.n740 4.5005
R12022 VPWR.n1725 VPWR.n1724 4.5005
R12023 VPWR.n1715 VPWR.n1714 4.5005
R12024 VPWR.n1237 VPWR.n917 4.5005
R12025 VPWR.n1593 VPWR.n1592 4.5005
R12026 VPWR.n1528 VPWR.n930 4.5005
R12027 VPWR.n1597 VPWR.n1233 4.5005
R12028 VPWR.n1520 VPWR.n1231 4.5005
R12029 VPWR.n1518 VPWR.n1228 4.5005
R12030 VPWR.n1511 VPWR.n1510 4.5005
R12031 VPWR.n1505 VPWR.n1504 4.5005
R12032 VPWR.n1497 VPWR.n1496 4.5005
R12033 VPWR.n1493 VPWR.n1492 4.5005
R12034 VPWR.n1485 VPWR.n1484 4.5005
R12035 VPWR.n1664 VPWR.n1169 4.5005
R12036 VPWR.n1668 VPWR.n1667 4.5005
R12037 VPWR.n1167 VPWR.n1159 4.5005
R12038 VPWR.n1677 VPWR.n1676 4.5005
R12039 VPWR.n1189 VPWR.n872 4.5005
R12040 VPWR.n1774 VPWR.n873 4.5005
R12041 VPWR.n1778 VPWR.n1777 4.5005
R12042 VPWR.n800 VPWR.n765 4.5005
R12043 VPWR.n1921 VPWR.n793 4.5005
R12044 VPWR.n1926 VPWR.n1925 4.5005
R12045 VPWR.n2074 VPWR.n623 4.5005
R12046 VPWR.n2132 VPWR.n627 4.5005
R12047 VPWR.n2131 VPWR.n683 4.5005
R12048 VPWR.n702 VPWR.n699 4.5005
R12049 VPWR.n507 VPWR.n488 4.5005
R12050 VPWR.n2422 VPWR.n2421 4.5005
R12051 VPWR.n500 VPWR.n499 4.5005
R12052 VPWR.n2553 VPWR.n371 4.5005
R12053 VPWR.n2736 VPWR.n2735 4.5005
R12054 VPWR.n369 VPWR.n368 4.5005
R12055 VPWR.n2759 VPWR.n2758 4.5005
R12056 VPWR.n2767 VPWR.n2766 4.5005
R12057 VPWR.n2771 VPWR.n2770 4.5005
R12058 VPWR.n2779 VPWR.n2778 4.5005
R12059 VPWR.n2783 VPWR.n2782 4.5005
R12060 VPWR.n2791 VPWR.n2790 4.5005
R12061 VPWR.n2795 VPWR.n2794 4.5005
R12062 VPWR.n2803 VPWR.n2802 4.5005
R12063 VPWR.n2807 VPWR.n2806 4.5005
R12064 VPWR.n2815 VPWR.n2814 4.5005
R12065 VPWR.n2819 VPWR.n2818 4.5005
R12066 VPWR.n2827 VPWR.n2826 4.5005
R12067 VPWR.n2831 VPWR.n2830 4.5005
R12068 VPWR.n2839 VPWR.n2838 4.5005
R12069 VPWR.n2843 VPWR.n2842 4.5005
R12070 VPWR.n2883 VPWR.n2849 4.5005
R12071 VPWR.n315 VPWR.n41 4.5005
R12072 VPWR.n2676 VPWR.n2675 4.5005
R12073 VPWR.n2671 VPWR.n417 4.5005
R12074 VPWR.n421 VPWR.n416 4.5005
R12075 VPWR.n2496 VPWR.n2495 4.5005
R12076 VPWR.n535 VPWR.n465 4.5005
R12077 VPWR.n2356 VPWR.n2355 4.5005
R12078 VPWR.n2256 VPWR.n541 4.5005
R12079 VPWR.n2236 VPWR.n2235 4.5005
R12080 VPWR.n595 VPWR.n590 4.5005
R12081 VPWR.n2023 VPWR.n2022 4.5005
R12082 VPWR.n2019 VPWR.n738 4.5005
R12083 VPWR.n832 VPWR.n737 4.5005
R12084 VPWR.n1861 VPWR.n1860 4.5005
R12085 VPWR.n1717 VPWR.n841 4.5005
R12086 VPWR.n1684 VPWR.n920 4.5005
R12087 VPWR.n1683 VPWR.n940 4.5005
R12088 VPWR.n2917 VPWR 4.49965
R12089 VPWR.n19 VPWR.n18 4.20017
R12090 VPWR.n963 VPWR.n962 4.20017
R12091 VPWR.n987 VPWR.n986 4.20017
R12092 VPWR.n1010 VPWR.n1009 4.20017
R12093 VPWR.n1045 VPWR.n1044 4.20017
R12094 VPWR.n1084 VPWR.n1083 4.20017
R12095 VPWR.n1122 VPWR.n1121 4.20017
R12096 VPWR.n3102 VPWR 4.14027
R12097 VPWR.n3086 VPWR 4.14027
R12098 VPWR.n3067 VPWR 4.14027
R12099 VPWR.n3047 VPWR 4.14027
R12100 VPWR.n3028 VPWR 4.14027
R12101 VPWR.n2992 VPWR 4.14027
R12102 VPWR.n2954 VPWR 4.14027
R12103 VPWR.n2882 VPWR.n2881 4.0005
R12104 VPWR.n3005 VPWR.n3002 3.76521
R12105 VPWR.n2969 VPWR.n2965 3.76521
R12106 VPWR.n2932 VPWR.n2928 3.76521
R12107 VPWR.n2900 VPWR.n2899 3.76521
R12108 VPWR.n37 VPWR 3.57245
R12109 VPWR.n857 VPWR.n856 3.4105
R12110 VPWR.n1956 VPWR.n717 3.4105
R12111 VPWR.n2050 VPWR.n2049 3.4105
R12112 VPWR.n705 VPWR.n608 3.4105
R12113 VPWR.n2176 VPWR.n2175 3.4105
R12114 VPWR.n2274 VPWR.n550 3.4105
R12115 VPWR.n2335 VPWR.n2334 3.4105
R12116 VPWR.n2337 VPWR.n2336 3.4105
R12117 VPWR.n2458 VPWR.n461 3.4105
R12118 VPWR.n2526 VPWR.n2525 3.4105
R12119 VPWR.n2631 VPWR.n396 3.4105
R12120 VPWR.n2630 VPWR.n2629 3.4105
R12121 VPWR.n2527 VPWR.n437 3.4105
R12122 VPWR.n2460 VPWR.n2459 3.4105
R12123 VPWR.n2301 VPWR.n474 3.4105
R12124 VPWR.n2307 VPWR.n2306 3.4105
R12125 VPWR.n2275 VPWR.n557 3.4105
R12126 VPWR.n2174 VPWR.n2173 3.4105
R12127 VPWR.n706 VPWR.n609 3.4105
R12128 VPWR.n2052 VPWR.n2051 3.4105
R12129 VPWR.n1957 VPWR.n716 3.4105
R12130 VPWR.n1894 VPWR.n1893 3.4105
R12131 VPWR.n1815 VPWR.n811 3.4105
R12132 VPWR.n1828 VPWR.n1827 3.4105
R12133 VPWR.n1830 VPWR.n1829 3.4105
R12134 VPWR.n855 VPWR.n749 3.4105
R12135 VPWR.n1981 VPWR.n1980 3.4105
R12136 VPWR.n1979 VPWR.n1978 3.4105
R12137 VPWR.n704 VPWR.n604 3.4105
R12138 VPWR.n2201 VPWR.n2200 3.4105
R12139 VPWR.n2273 VPWR.n552 3.4105
R12140 VPWR.n2333 VPWR.n2332 3.4105
R12141 VPWR.n2338 VPWR.n463 3.4105
R12142 VPWR.n2504 VPWR.n2503 3.4105
R12143 VPWR.n2506 VPWR.n2505 3.4105
R12144 VPWR.n2632 VPWR.n397 3.4105
R12145 VPWR.n2574 VPWR.n388 3.4105
R12146 VPWR.n2529 VPWR.n2528 3.4105
R12147 VPWR.n2457 VPWR.n460 3.4105
R12148 VPWR.n2303 VPWR.n2302 3.4105
R12149 VPWR.n2305 VPWR.n2304 3.4105
R12150 VPWR.n2276 VPWR.n558 3.4105
R12151 VPWR.n2164 VPWR.n2163 3.4105
R12152 VPWR.n707 VPWR.n612 3.4105
R12153 VPWR.n756 VPWR.n755 3.4105
R12154 VPWR.n1959 VPWR.n1958 3.4105
R12155 VPWR.n1895 VPWR.n754 3.4105
R12156 VPWR.n1817 VPWR.n1816 3.4105
R12157 VPWR.n1843 VPWR.n1842 3.4105
R12158 VPWR.n854 VPWR.n748 3.4105
R12159 VPWR.n1983 VPWR.n1982 3.4105
R12160 VPWR.n1977 VPWR.n601 3.4105
R12161 VPWR.n2206 VPWR.n2205 3.4105
R12162 VPWR.n2204 VPWR.n2203 3.4105
R12163 VPWR.n2272 VPWR.n548 3.4105
R12164 VPWR.n2342 VPWR.n2341 3.4105
R12165 VPWR.n2340 VPWR.n2339 3.4105
R12166 VPWR.n2502 VPWR.n432 3.4105
R12167 VPWR.n2640 VPWR.n2639 3.4105
R12168 VPWR.n2638 VPWR.n2637 3.4105
R12169 VPWR.n436 VPWR.n435 3.4105
R12170 VPWR.n2701 VPWR.n2700 3.4105
R12171 VPWR.n2703 VPWR.n2702 3.4105
R12172 VPWR.n439 VPWR.n438 3.4105
R12173 VPWR.n2713 VPWR.n2712 3.4105
R12174 VPWR.n2715 VPWR.n2714 3.4105
R12175 VPWR.n2575 VPWR.n387 3.4105
R12176 VPWR.n2454 VPWR.n2453 3.4105
R12177 VPWR.n2456 VPWR.n2455 3.4105
R12178 VPWR.n2300 VPWR.n475 3.4105
R12179 VPWR.n2283 VPWR.n2282 3.4105
R12180 VPWR.n2277 VPWR.n574 3.4105
R12181 VPWR.n2162 VPWR.n2161 3.4105
R12182 VPWR.n708 VPWR.n613 3.4105
R12183 VPWR.n2062 VPWR.n2061 3.4105
R12184 VPWR.n1955 VPWR.n711 3.4105
R12185 VPWR.n1897 VPWR.n1896 3.4105
R12186 VPWR.n1814 VPWR.n810 3.4105
R12187 VPWR.n1755 VPWR.n1754 3.4105
R12188 VPWR.n1753 VPWR.n861 3.4105
R12189 VPWR.n1752 VPWR.n1751 3.4105
R12190 VPWR.n912 VPWR.n852 3.4105
R12191 VPWR.n913 VPWR.n851 3.4105
R12192 VPWR.n914 VPWR.n848 3.4105
R12193 VPWR.n915 VPWR.n847 3.4105
R12194 VPWR.n1845 VPWR.n1844 3.4105
R12195 VPWR.n853 VPWR.n743 3.4105
R12196 VPWR.n2008 VPWR.n2007 3.4105
R12197 VPWR.n1976 VPWR.n600 3.4105
R12198 VPWR.n2210 VPWR.n2209 3.4105
R12199 VPWR.n2202 VPWR.n577 3.4105
R12200 VPWR.n2271 VPWR.n2270 3.4105
R12201 VPWR.n2343 VPWR.n526 3.4105
R12202 VPWR.n2374 VPWR.n2373 3.4105
R12203 VPWR.n2501 VPWR.n431 3.4105
R12204 VPWR.n2642 VPWR.n2641 3.4105
R12205 VPWR.n2636 VPWR.n405 3.4105
R12206 VPWR.n2691 VPWR.n2690 3.4105
R12207 VPWR.n448 VPWR.n447 3.4105
R12208 VPWR.n2577 VPWR.n2576 3.4105
R12209 VPWR.n2452 VPWR.n446 3.4105
R12210 VPWR.n2447 VPWR.n2446 3.4105
R12211 VPWR.n2299 VPWR.n479 3.4105
R12212 VPWR.n2281 VPWR.n2280 3.4105
R12213 VPWR.n2279 VPWR.n2278 3.4105
R12214 VPWR.n2149 VPWR.n575 3.4105
R12215 VPWR.n2119 VPWR.n2118 3.4105
R12216 VPWR.n2064 VPWR.n2063 3.4105
R12217 VPWR.n1954 VPWR.n709 3.4105
R12218 VPWR.n1811 VPWR.n1810 3.4105
R12219 VPWR.n1813 VPWR.n1812 3.4105
R12220 VPWR.n891 VPWR.n862 3.4105
R12221 VPWR.n916 VPWR.n839 3.4105
R12222 VPWR.n1866 VPWR.n1865 3.4105
R12223 VPWR.n1868 VPWR.n1867 3.4105
R12224 VPWR.n2009 VPWR.n728 3.4105
R12225 VPWR.n2033 VPWR.n2032 3.4105
R12226 VPWR.n2208 VPWR.n583 3.4105
R12227 VPWR.n2246 VPWR.n2245 3.4105
R12228 VPWR.n2248 VPWR.n2247 3.4105
R12229 VPWR.n2344 VPWR.n527 3.4105
R12230 VPWR.n2372 VPWR.n2371 3.4105
R12231 VPWR.n2500 VPWR.n428 3.4105
R12232 VPWR.n2652 VPWR.n2651 3.4105
R12233 VPWR.n2635 VPWR.n406 3.4105
R12234 VPWR.n2689 VPWR.n2688 3.4105
R12235 VPWR.n2742 VPWR.n52 3.4105
R12236 VPWR.n2743 VPWR.n53 3.4105
R12237 VPWR.n2744 VPWR.n58 3.4105
R12238 VPWR.n2745 VPWR.n59 3.4105
R12239 VPWR.n2746 VPWR.n64 3.4105
R12240 VPWR.n2747 VPWR.n65 3.4105
R12241 VPWR.n2748 VPWR.n70 3.4105
R12242 VPWR.n2749 VPWR.n71 3.4105
R12243 VPWR.n2750 VPWR.n76 3.4105
R12244 VPWR.n2751 VPWR.n77 3.4105
R12245 VPWR.n2725 VPWR.n2724 3.4105
R12246 VPWR.n2573 VPWR.n379 3.4105
R12247 VPWR.n2451 VPWR.n2450 3.4105
R12248 VPWR.n2449 VPWR.n2448 3.4105
R12249 VPWR.n2298 VPWR.n477 3.4105
R12250 VPWR.n2293 VPWR.n2292 3.4105
R12251 VPWR.n2127 VPWR.n562 3.4105
R12252 VPWR.n2151 VPWR.n2150 3.4105
R12253 VPWR.n2120 VPWR.n617 3.4105
R12254 VPWR.n1951 VPWR.n1950 3.4105
R12255 VPWR.n1953 VPWR.n1952 3.4105
R12256 VPWR.n1809 VPWR.n757 3.4105
R12257 VPWR.n1804 VPWR.n1803 3.4105
R12258 VPWR.n890 VPWR.n866 3.4105
R12259 VPWR.n1728 VPWR.n1727 3.4105
R12260 VPWR.n1864 VPWR.n838 3.4105
R12261 VPWR.n1870 VPWR.n1869 3.4105
R12262 VPWR.n2010 VPWR.n729 3.4105
R12263 VPWR.n2031 VPWR.n2030 3.4105
R12264 VPWR.n2207 VPWR.n585 3.4105
R12265 VPWR.n2244 VPWR.n2243 3.4105
R12266 VPWR.n2249 VPWR.n545 3.4105
R12267 VPWR.n2347 VPWR.n2346 3.4105
R12268 VPWR.n547 VPWR.n546 3.4105
R12269 VPWR.n2499 VPWR.n424 3.4105
R12270 VPWR.n2654 VPWR.n2653 3.4105
R12271 VPWR.n2634 VPWR.n427 3.4105
R12272 VPWR.n426 VPWR.n425 3.4105
R12273 VPWR.n2741 VPWR.n47 3.4105
R12274 VPWR.n2752 VPWR.n82 3.4105
R12275 VPWR.n2727 VPWR.n2726 3.4105
R12276 VPWR.n2572 VPWR.n378 3.4105
R12277 VPWR.n2546 VPWR.n2545 3.4105
R12278 VPWR.n2418 VPWR.n452 3.4105
R12279 VPWR.n2297 VPWR.n2296 3.4105
R12280 VPWR.n2295 VPWR.n2294 3.4105
R12281 VPWR.n2128 VPWR.n560 3.4105
R12282 VPWR.n2148 VPWR.n2147 3.4105
R12283 VPWR.n2121 VPWR.n618 3.4105
R12284 VPWR.n1949 VPWR.n1948 3.4105
R12285 VPWR.n1918 VPWR.n760 3.4105
R12286 VPWR.n1808 VPWR.n1807 3.4105
R12287 VPWR.n1806 VPWR.n1805 3.4105
R12288 VPWR.n889 VPWR.n864 3.4105
R12289 VPWR.n1422 VPWR.n1166 3.4105
R12290 VPWR.n1663 VPWR.n1170 3.4105
R12291 VPWR.n1482 VPWR.n1481 3.4105
R12292 VPWR.n1479 VPWR.n888 3.4105
R12293 VPWR.n1477 VPWR.n1268 3.4105
R12294 VPWR.n1475 VPWR.n892 3.4105
R12295 VPWR.n1473 VPWR.n1263 3.4105
R12296 VPWR.n1640 VPWR.n1639 3.4105
R12297 VPWR.n1637 VPWR.n1636 3.4105
R12298 VPWR.n1614 VPWR.n1613 3.4105
R12299 VPWR.n1700 VPWR.n1699 3.4105
R12300 VPWR.n1697 VPWR.n911 3.4105
R12301 VPWR.n1431 VPWR.n874 3.4105
R12302 VPWR.n1772 VPWR.n1771 3.4105
R12303 VPWR.n1775 VPWR.n795 3.4105
R12304 VPWR.n1914 VPWR.n1913 3.4105
R12305 VPWR.n1919 VPWR.n764 3.4105
R12306 VPWR.n1929 VPWR.n1928 3.4105
R12307 VPWR.n2122 VPWR.n621 3.4105
R12308 VPWR.n2135 VPWR.n2134 3.4105
R12309 VPWR.n2129 VPWR.n622 3.4105
R12310 VPWR.n700 VPWR.n502 3.4105
R12311 VPWR.n2412 VPWR.n2411 3.4105
R12312 VPWR.n2419 VPWR.n450 3.4105
R12313 VPWR.n2548 VPWR.n2547 3.4105
R12314 VPWR.n2571 VPWR.n2570 3.4105
R12315 VPWR.n2569 VPWR.n2568 3.4105
R12316 VPWR.n2753 VPWR.n83 3.4105
R12317 VPWR.n2768 VPWR.n2767 3.4105
R12318 VPWR.n2770 VPWR.n2769 3.4105
R12319 VPWR.n2780 VPWR.n2779 3.4105
R12320 VPWR.n2782 VPWR.n2781 3.4105
R12321 VPWR.n2792 VPWR.n2791 3.4105
R12322 VPWR.n2794 VPWR.n2793 3.4105
R12323 VPWR.n2804 VPWR.n2803 3.4105
R12324 VPWR.n2806 VPWR.n2805 3.4105
R12325 VPWR.n2816 VPWR.n2815 3.4105
R12326 VPWR.n2818 VPWR.n2817 3.4105
R12327 VPWR.n2828 VPWR.n2827 3.4105
R12328 VPWR.n2830 VPWR.n2829 3.4105
R12329 VPWR.n2840 VPWR.n2839 3.4105
R12330 VPWR.n2842 VPWR.n2841 3.4105
R12331 VPWR.n2740 VPWR.n46 3.4105
R12332 VPWR.n2679 VPWR.n2678 3.4105
R12333 VPWR.n2633 VPWR.n414 3.4105
R12334 VPWR.n2666 VPWR.n2665 3.4105
R12335 VPWR.n2498 VPWR.n419 3.4105
R12336 VPWR.n2362 VPWR.n2361 3.4105
R12337 VPWR.n2345 VPWR.n539 3.4105
R12338 VPWR.n2252 VPWR.n2251 3.4105
R12339 VPWR.n591 VPWR.n582 3.4105
R12340 VPWR.n2230 VPWR.n2229 3.4105
R12341 VPWR.n2020 VPWR.n593 3.4105
R12342 VPWR.n2012 VPWR.n2011 3.4105
R12343 VPWR.n2014 VPWR.n2013 3.4105
R12344 VPWR.n1863 VPWR.n740 3.4105
R12345 VPWR.n1726 VPWR.n1725 3.4105
R12346 VPWR.n1715 VPWR.n918 3.4105
R12347 VPWR.n1429 VPWR.n872 3.4105
R12348 VPWR.n1774 VPWR.n1773 3.4105
R12349 VPWR.n1777 VPWR.n1776 3.4105
R12350 VPWR.n1915 VPWR.n765 3.4105
R12351 VPWR.n1921 VPWR.n1920 3.4105
R12352 VPWR.n1927 VPWR.n1926 3.4105
R12353 VPWR.n2123 VPWR.n623 3.4105
R12354 VPWR.n2133 VPWR.n2132 3.4105
R12355 VPWR.n2131 VPWR.n2130 3.4105
R12356 VPWR.n702 VPWR.n701 3.4105
R12357 VPWR.n2413 VPWR.n488 3.4105
R12358 VPWR.n2421 VPWR.n2420 3.4105
R12359 VPWR.n2415 VPWR.n500 3.4105
R12360 VPWR.n449 VPWR.n371 3.4105
R12361 VPWR.n2737 VPWR.n2736 3.4105
R12362 VPWR.n2754 VPWR.n369 3.4105
R12363 VPWR.n2758 VPWR.n2757 3.4105
R12364 VPWR.n2884 VPWR.n2883 3.4105
R12365 VPWR.n2739 VPWR.n41 3.4105
R12366 VPWR.n2677 VPWR.n2676 3.4105
R12367 VPWR.n2671 VPWR.n2670 3.4105
R12368 VPWR.n2667 VPWR.n416 3.4105
R12369 VPWR.n2497 VPWR.n2496 3.4105
R12370 VPWR.n2360 VPWR.n465 3.4105
R12371 VPWR.n2357 VPWR.n2356 3.4105
R12372 VPWR.n2250 VPWR.n541 3.4105
R12373 VPWR.n2235 VPWR.n2234 3.4105
R12374 VPWR.n2231 VPWR.n590 3.4105
R12375 VPWR.n2022 VPWR.n2021 3.4105
R12376 VPWR.n2019 VPWR.n2018 3.4105
R12377 VPWR.n2015 VPWR.n737 3.4105
R12378 VPWR.n1862 VPWR.n1861 3.4105
R12379 VPWR.n937 VPWR.n841 3.4105
R12380 VPWR.n1685 VPWR.n1684 3.4105
R12381 VPWR.n1683 VPWR.n1682 3.4105
R12382 VPWR.n1234 VPWR.n917 3.4105
R12383 VPWR.n1594 VPWR.n1593 3.4105
R12384 VPWR.n1595 VPWR.n930 3.4105
R12385 VPWR.n1597 VPWR.n1596 3.4105
R12386 VPWR.n1507 VPWR.n1231 3.4105
R12387 VPWR.n1508 VPWR.n1228 3.4105
R12388 VPWR.n1510 VPWR.n1509 3.4105
R12389 VPWR.n1506 VPWR.n1505 3.4105
R12390 VPWR.n1496 VPWR.n1495 3.4105
R12391 VPWR.n1494 VPWR.n1493 3.4105
R12392 VPWR.n1484 VPWR.n1483 3.4105
R12393 VPWR.n1665 VPWR.n1664 3.4105
R12394 VPWR.n1667 VPWR.n1666 3.4105
R12395 VPWR.n1168 VPWR.n1167 3.4105
R12396 VPWR.n1678 VPWR.n1677 3.4105
R12397 VPWR.n1053 VPWR.n1049 3.38874
R12398 VPWR.n1092 VPWR.n1088 3.38874
R12399 VPWR.n1129 VPWR.n1125 3.38874
R12400 VPWR.n2855 VPWR.n2853 3.36211
R12401 VPWR.n2857 VPWR.n2855 3.36211
R12402 VPWR.n2859 VPWR.n2857 3.36211
R12403 VPWR.n2861 VPWR.n2859 3.36211
R12404 VPWR.n2863 VPWR.n2861 3.36211
R12405 VPWR.n2865 VPWR.n2863 3.36211
R12406 VPWR.n2867 VPWR.n2865 3.36211
R12407 VPWR.n2869 VPWR.n2867 3.36211
R12408 VPWR.n2871 VPWR.n2869 3.36211
R12409 VPWR.n2873 VPWR.n2871 3.36211
R12410 VPWR.n2875 VPWR.n2873 3.36211
R12411 VPWR.n2877 VPWR.n2875 3.36211
R12412 VPWR.n2879 VPWR.n2877 3.36211
R12413 VPWR.n2881 VPWR.n2879 3.36211
R12414 VPWR.t415 VPWR.t1799 3.35739
R12415 VPWR.t1873 VPWR.t706 3.35739
R12416 VPWR.n1510 VPWR.n1263 3.28012
R12417 VPWR.n1505 VPWR.n892 3.28012
R12418 VPWR.n1640 VPWR.n1228 3.28012
R12419 VPWR.n1496 VPWR.n1268 3.28012
R12420 VPWR.n1636 VPWR.n1231 3.28012
R12421 VPWR.n1493 VPWR.n888 3.28012
R12422 VPWR.n1614 VPWR.n1597 3.28012
R12423 VPWR.n1484 VPWR.n1482 3.28012
R12424 VPWR.n1700 VPWR.n930 3.28012
R12425 VPWR.n1664 VPWR.n1663 3.28012
R12426 VPWR.n1593 VPWR.n911 3.28012
R12427 VPWR.n1667 VPWR.n1166 3.28012
R12428 VPWR.n1167 VPWR.n874 3.28012
R12429 VPWR.n1715 VPWR.n917 3.28012
R12430 VPWR.n1677 VPWR.n872 3.28012
R12431 VPWR.n1684 VPWR.n1683 3.28012
R12432 VPWR.n2839 VPWR.n47 3.235
R12433 VPWR.n2830 VPWR.n52 3.235
R12434 VPWR.n2827 VPWR.n53 3.235
R12435 VPWR.n2818 VPWR.n58 3.235
R12436 VPWR.n2815 VPWR.n59 3.235
R12437 VPWR.n2806 VPWR.n64 3.235
R12438 VPWR.n2803 VPWR.n65 3.235
R12439 VPWR.n2794 VPWR.n70 3.235
R12440 VPWR.n2791 VPWR.n71 3.235
R12441 VPWR.n2782 VPWR.n76 3.235
R12442 VPWR.n2779 VPWR.n77 3.235
R12443 VPWR.n2770 VPWR.n82 3.235
R12444 VPWR.n2767 VPWR.n83 3.235
R12445 VPWR.n2842 VPWR.n46 3.235
R12446 VPWR.n2758 VPWR.n369 3.235
R12447 VPWR.n2883 VPWR.n41 3.21882
R12448 VPWR.n1032 VPWR.n1030 3.01226
R12449 VPWR.n1263 VPWR.n852 2.94005
R12450 VPWR.n1751 VPWR.n892 2.94005
R12451 VPWR.n1640 VPWR.n851 2.94005
R12452 VPWR.n1268 VPWR.n861 2.94005
R12453 VPWR.n1636 VPWR.n848 2.94005
R12454 VPWR.n1755 VPWR.n888 2.94005
R12455 VPWR.n1614 VPWR.n847 2.94005
R12456 VPWR.n1482 VPWR.n862 2.94005
R12457 VPWR.n1700 VPWR.n839 2.94005
R12458 VPWR.n1663 VPWR.n866 2.94005
R12459 VPWR.n1728 VPWR.n911 2.94005
R12460 VPWR.n1166 VPWR.n864 2.94005
R12461 VPWR.n1771 VPWR.n874 2.94005
R12462 VPWR.n1725 VPWR.n1715 2.94005
R12463 VPWR.n1774 VPWR.n872 2.94005
R12464 VPWR.n1684 VPWR.n841 2.94005
R12465 VPWR.n2691 VPWR.n53 2.89493
R12466 VPWR.n436 VPWR.n58 2.89493
R12467 VPWR.n2700 VPWR.n59 2.89493
R12468 VPWR.n2700 VPWR.n397 2.89493
R12469 VPWR.n2703 VPWR.n64 2.89493
R12470 VPWR.n2703 VPWR.n396 2.89493
R12471 VPWR.n1827 VPWR.n852 2.89493
R12472 VPWR.n1827 VPWR.n857 2.89493
R12473 VPWR.n857 VPWR.n717 2.89493
R12474 VPWR.n2049 VPWR.n717 2.89493
R12475 VPWR.n2049 VPWR.n608 2.89493
R12476 VPWR.n2176 VPWR.n608 2.89493
R12477 VPWR.n2176 VPWR.n550 2.89493
R12478 VPWR.n2335 VPWR.n550 2.89493
R12479 VPWR.n2336 VPWR.n2335 2.89493
R12480 VPWR.n2336 VPWR.n461 2.89493
R12481 VPWR.n2525 VPWR.n461 2.89493
R12482 VPWR.n2525 VPWR.n396 2.89493
R12483 VPWR.n439 VPWR.n65 2.89493
R12484 VPWR.n2629 VPWR.n439 2.89493
R12485 VPWR.n2629 VPWR.n437 2.89493
R12486 VPWR.n2460 VPWR.n437 2.89493
R12487 VPWR.n2460 VPWR.n474 2.89493
R12488 VPWR.n2307 VPWR.n474 2.89493
R12489 VPWR.n2307 VPWR.n557 2.89493
R12490 VPWR.n2173 VPWR.n557 2.89493
R12491 VPWR.n2173 VPWR.n609 2.89493
R12492 VPWR.n2052 VPWR.n609 2.89493
R12493 VPWR.n2052 VPWR.n716 2.89493
R12494 VPWR.n1893 VPWR.n716 2.89493
R12495 VPWR.n1893 VPWR.n811 2.89493
R12496 VPWR.n1751 VPWR.n811 2.89493
R12497 VPWR.n1830 VPWR.n851 2.89493
R12498 VPWR.n1830 VPWR.n749 2.89493
R12499 VPWR.n1980 VPWR.n749 2.89493
R12500 VPWR.n1980 VPWR.n1979 2.89493
R12501 VPWR.n1979 VPWR.n604 2.89493
R12502 VPWR.n2200 VPWR.n604 2.89493
R12503 VPWR.n2200 VPWR.n552 2.89493
R12504 VPWR.n2332 VPWR.n552 2.89493
R12505 VPWR.n2332 VPWR.n463 2.89493
R12506 VPWR.n2504 VPWR.n463 2.89493
R12507 VPWR.n2506 VPWR.n2504 2.89493
R12508 VPWR.n2506 VPWR.n397 2.89493
R12509 VPWR.n2712 VPWR.n70 2.89493
R12510 VPWR.n2712 VPWR.n388 2.89493
R12511 VPWR.n2529 VPWR.n388 2.89493
R12512 VPWR.n2529 VPWR.n460 2.89493
R12513 VPWR.n2303 VPWR.n460 2.89493
R12514 VPWR.n2304 VPWR.n2303 2.89493
R12515 VPWR.n2304 VPWR.n558 2.89493
R12516 VPWR.n2164 VPWR.n558 2.89493
R12517 VPWR.n2164 VPWR.n612 2.89493
R12518 VPWR.n756 VPWR.n612 2.89493
R12519 VPWR.n1959 VPWR.n756 2.89493
R12520 VPWR.n1959 VPWR.n754 2.89493
R12521 VPWR.n1817 VPWR.n754 2.89493
R12522 VPWR.n1817 VPWR.n861 2.89493
R12523 VPWR.n1842 VPWR.n848 2.89493
R12524 VPWR.n1842 VPWR.n748 2.89493
R12525 VPWR.n1983 VPWR.n748 2.89493
R12526 VPWR.n1983 VPWR.n601 2.89493
R12527 VPWR.n2205 VPWR.n601 2.89493
R12528 VPWR.n2205 VPWR.n2204 2.89493
R12529 VPWR.n2204 VPWR.n548 2.89493
R12530 VPWR.n2341 VPWR.n548 2.89493
R12531 VPWR.n2341 VPWR.n2340 2.89493
R12532 VPWR.n2340 VPWR.n432 2.89493
R12533 VPWR.n2639 VPWR.n432 2.89493
R12534 VPWR.n2639 VPWR.n2638 2.89493
R12535 VPWR.n2638 VPWR.n436 2.89493
R12536 VPWR.n2715 VPWR.n71 2.89493
R12537 VPWR.n2715 VPWR.n387 2.89493
R12538 VPWR.n2454 VPWR.n387 2.89493
R12539 VPWR.n2455 VPWR.n2454 2.89493
R12540 VPWR.n2455 VPWR.n475 2.89493
R12541 VPWR.n2283 VPWR.n475 2.89493
R12542 VPWR.n2283 VPWR.n574 2.89493
R12543 VPWR.n2161 VPWR.n574 2.89493
R12544 VPWR.n2161 VPWR.n613 2.89493
R12545 VPWR.n2061 VPWR.n613 2.89493
R12546 VPWR.n2061 VPWR.n711 2.89493
R12547 VPWR.n1897 VPWR.n711 2.89493
R12548 VPWR.n1897 VPWR.n810 2.89493
R12549 VPWR.n1755 VPWR.n810 2.89493
R12550 VPWR.n1845 VPWR.n847 2.89493
R12551 VPWR.n1845 VPWR.n743 2.89493
R12552 VPWR.n2007 VPWR.n743 2.89493
R12553 VPWR.n2007 VPWR.n600 2.89493
R12554 VPWR.n2210 VPWR.n600 2.89493
R12555 VPWR.n2210 VPWR.n577 2.89493
R12556 VPWR.n2270 VPWR.n577 2.89493
R12557 VPWR.n2270 VPWR.n526 2.89493
R12558 VPWR.n2374 VPWR.n526 2.89493
R12559 VPWR.n2374 VPWR.n431 2.89493
R12560 VPWR.n2642 VPWR.n431 2.89493
R12561 VPWR.n2642 VPWR.n405 2.89493
R12562 VPWR.n2691 VPWR.n405 2.89493
R12563 VPWR.n448 VPWR.n76 2.89493
R12564 VPWR.n2577 VPWR.n448 2.89493
R12565 VPWR.n2577 VPWR.n446 2.89493
R12566 VPWR.n2446 VPWR.n446 2.89493
R12567 VPWR.n2446 VPWR.n479 2.89493
R12568 VPWR.n2280 VPWR.n479 2.89493
R12569 VPWR.n2280 VPWR.n2279 2.89493
R12570 VPWR.n2279 VPWR.n575 2.89493
R12571 VPWR.n2118 VPWR.n575 2.89493
R12572 VPWR.n2118 VPWR.n2064 2.89493
R12573 VPWR.n2064 VPWR.n709 2.89493
R12574 VPWR.n1811 VPWR.n709 2.89493
R12575 VPWR.n1812 VPWR.n1811 2.89493
R12576 VPWR.n1812 VPWR.n862 2.89493
R12577 VPWR.n1866 VPWR.n839 2.89493
R12578 VPWR.n1867 VPWR.n1866 2.89493
R12579 VPWR.n1867 VPWR.n728 2.89493
R12580 VPWR.n2033 VPWR.n728 2.89493
R12581 VPWR.n2033 VPWR.n583 2.89493
R12582 VPWR.n2246 VPWR.n583 2.89493
R12583 VPWR.n2247 VPWR.n2246 2.89493
R12584 VPWR.n2247 VPWR.n527 2.89493
R12585 VPWR.n2371 VPWR.n527 2.89493
R12586 VPWR.n2371 VPWR.n428 2.89493
R12587 VPWR.n2651 VPWR.n428 2.89493
R12588 VPWR.n2651 VPWR.n406 2.89493
R12589 VPWR.n2688 VPWR.n406 2.89493
R12590 VPWR.n2688 VPWR.n52 2.89493
R12591 VPWR.n2724 VPWR.n77 2.89493
R12592 VPWR.n2724 VPWR.n379 2.89493
R12593 VPWR.n2450 VPWR.n379 2.89493
R12594 VPWR.n2450 VPWR.n2449 2.89493
R12595 VPWR.n2449 VPWR.n477 2.89493
R12596 VPWR.n2292 VPWR.n477 2.89493
R12597 VPWR.n2292 VPWR.n562 2.89493
R12598 VPWR.n2151 VPWR.n562 2.89493
R12599 VPWR.n2151 VPWR.n617 2.89493
R12600 VPWR.n1951 VPWR.n617 2.89493
R12601 VPWR.n1952 VPWR.n1951 2.89493
R12602 VPWR.n1952 VPWR.n757 2.89493
R12603 VPWR.n1803 VPWR.n757 2.89493
R12604 VPWR.n1803 VPWR.n866 2.89493
R12605 VPWR.n1728 VPWR.n838 2.89493
R12606 VPWR.n1870 VPWR.n838 2.89493
R12607 VPWR.n1870 VPWR.n729 2.89493
R12608 VPWR.n2030 VPWR.n729 2.89493
R12609 VPWR.n2030 VPWR.n585 2.89493
R12610 VPWR.n2243 VPWR.n585 2.89493
R12611 VPWR.n2243 VPWR.n545 2.89493
R12612 VPWR.n2347 VPWR.n545 2.89493
R12613 VPWR.n2347 VPWR.n547 2.89493
R12614 VPWR.n547 VPWR.n424 2.89493
R12615 VPWR.n2654 VPWR.n424 2.89493
R12616 VPWR.n2654 VPWR.n427 2.89493
R12617 VPWR.n427 VPWR.n426 2.89493
R12618 VPWR.n426 VPWR.n47 2.89493
R12619 VPWR.n2727 VPWR.n82 2.89493
R12620 VPWR.n2727 VPWR.n378 2.89493
R12621 VPWR.n2545 VPWR.n378 2.89493
R12622 VPWR.n2545 VPWR.n452 2.89493
R12623 VPWR.n2296 VPWR.n452 2.89493
R12624 VPWR.n2296 VPWR.n2295 2.89493
R12625 VPWR.n2295 VPWR.n560 2.89493
R12626 VPWR.n2147 VPWR.n560 2.89493
R12627 VPWR.n2147 VPWR.n618 2.89493
R12628 VPWR.n1948 VPWR.n618 2.89493
R12629 VPWR.n1948 VPWR.n760 2.89493
R12630 VPWR.n1807 VPWR.n760 2.89493
R12631 VPWR.n1807 VPWR.n1806 2.89493
R12632 VPWR.n1806 VPWR.n864 2.89493
R12633 VPWR.n1771 VPWR.n795 2.89493
R12634 VPWR.n1913 VPWR.n795 2.89493
R12635 VPWR.n1913 VPWR.n764 2.89493
R12636 VPWR.n1929 VPWR.n764 2.89493
R12637 VPWR.n1929 VPWR.n621 2.89493
R12638 VPWR.n2135 VPWR.n621 2.89493
R12639 VPWR.n2135 VPWR.n622 2.89493
R12640 VPWR.n622 VPWR.n502 2.89493
R12641 VPWR.n2411 VPWR.n502 2.89493
R12642 VPWR.n2411 VPWR.n450 2.89493
R12643 VPWR.n2548 VPWR.n450 2.89493
R12644 VPWR.n2570 VPWR.n2548 2.89493
R12645 VPWR.n2570 VPWR.n2569 2.89493
R12646 VPWR.n2569 VPWR.n83 2.89493
R12647 VPWR.n2679 VPWR.n46 2.89493
R12648 VPWR.n2679 VPWR.n414 2.89493
R12649 VPWR.n2665 VPWR.n414 2.89493
R12650 VPWR.n2665 VPWR.n419 2.89493
R12651 VPWR.n2362 VPWR.n419 2.89493
R12652 VPWR.n2362 VPWR.n539 2.89493
R12653 VPWR.n2252 VPWR.n539 2.89493
R12654 VPWR.n2252 VPWR.n582 2.89493
R12655 VPWR.n2229 VPWR.n582 2.89493
R12656 VPWR.n2229 VPWR.n593 2.89493
R12657 VPWR.n2012 VPWR.n593 2.89493
R12658 VPWR.n2013 VPWR.n2012 2.89493
R12659 VPWR.n2013 VPWR.n740 2.89493
R12660 VPWR.n1725 VPWR.n740 2.89493
R12661 VPWR.n1777 VPWR.n1774 2.89493
R12662 VPWR.n1777 VPWR.n765 2.89493
R12663 VPWR.n1921 VPWR.n765 2.89493
R12664 VPWR.n1926 VPWR.n1921 2.89493
R12665 VPWR.n1926 VPWR.n623 2.89493
R12666 VPWR.n2132 VPWR.n623 2.89493
R12667 VPWR.n2132 VPWR.n2131 2.89493
R12668 VPWR.n2131 VPWR.n702 2.89493
R12669 VPWR.n702 VPWR.n488 2.89493
R12670 VPWR.n2421 VPWR.n488 2.89493
R12671 VPWR.n2421 VPWR.n500 2.89493
R12672 VPWR.n500 VPWR.n371 2.89493
R12673 VPWR.n2736 VPWR.n371 2.89493
R12674 VPWR.n2736 VPWR.n369 2.89493
R12675 VPWR.n2676 VPWR.n41 2.89493
R12676 VPWR.n2676 VPWR.n2671 2.89493
R12677 VPWR.n2671 VPWR.n416 2.89493
R12678 VPWR.n2496 VPWR.n416 2.89493
R12679 VPWR.n2496 VPWR.n465 2.89493
R12680 VPWR.n2356 VPWR.n465 2.89493
R12681 VPWR.n2356 VPWR.n541 2.89493
R12682 VPWR.n2235 VPWR.n541 2.89493
R12683 VPWR.n2235 VPWR.n590 2.89493
R12684 VPWR.n2022 VPWR.n590 2.89493
R12685 VPWR.n2022 VPWR.n2019 2.89493
R12686 VPWR.n2019 VPWR.n737 2.89493
R12687 VPWR.n1861 VPWR.n737 2.89493
R12688 VPWR.n1861 VPWR.n841 2.89493
R12689 VPWR.n1036 VPWR.n1012 2.63579
R12690 VPWR.n3105 VPWR.t222 2.48308
R12691 VPWR.n3020 VPWR.n3019 2.25932
R12692 VPWR.n1680 VPWR.n1154 2.06026
R12693 VPWR.n1681 VPWR.n1680 1.78803
R12694 VPWR.n1685 VPWR.n939 1.32852
R12695 VPWR.n2668 VPWR.n2667 1.32852
R12696 VPWR.n2497 VPWR.n418 1.32852
R12697 VPWR.n2360 VPWR.n2359 1.32852
R12698 VPWR.n2358 VPWR.n2357 1.32852
R12699 VPWR.n2250 VPWR.n540 1.32852
R12700 VPWR.n2234 VPWR.n2233 1.32852
R12701 VPWR.n2232 VPWR.n2231 1.32852
R12702 VPWR.n2021 VPWR.n592 1.32852
R12703 VPWR.n2018 VPWR.n2017 1.32852
R12704 VPWR.n2016 VPWR.n2015 1.32852
R12705 VPWR.n2670 VPWR.n2669 1.32852
R12706 VPWR.n1862 VPWR.n739 1.32852
R12707 VPWR.n2677 VPWR.n415 1.32852
R12708 VPWR.n938 VPWR.n937 1.32852
R12709 VPWR.n2739 VPWR.n40 1.32852
R12710 VPWR.n2885 VPWR.n2884 1.32852
R12711 VPWR.n1682 VPWR.n1681 1.32852
R12712 VPWR.n3127 VPWR.n23 1.29068
R12713 VPWR.n3113 VPWR.n21 1.28175
R12714 VPWR VPWR.n1156 1.25994
R12715 VPWR.n2755 VPWR 1.25994
R12716 VPWR.n2738 VPWR 1.25994
R12717 VPWR VPWR.n370 1.25994
R12718 VPWR.n2416 VPWR 1.25994
R12719 VPWR VPWR.n2417 1.25994
R12720 VPWR.n2414 VPWR 1.25994
R12721 VPWR VPWR.n501 1.25994
R12722 VPWR VPWR.n2126 1.25994
R12723 VPWR.n2125 VPWR 1.25994
R12724 VPWR.n2124 VPWR 1.25994
R12725 VPWR VPWR.n703 1.25994
R12726 VPWR VPWR.n1917 1.25994
R12727 VPWR.n1916 VPWR 1.25994
R12728 VPWR VPWR.n794 1.25994
R12729 VPWR.n1155 VPWR 1.25994
R12730 VPWR VPWR.n2756 1.25994
R12731 VPWR.n1679 VPWR 1.25994
R12732 VPWR.n2886 VPWR.n2885 1.144
R12733 VPWR VPWR.n498 1.04685
R12734 VPWR.n453 VPWR 1.04685
R12735 VPWR VPWR.n2543 1.04685
R12736 VPWR.n2538 VPWR 1.04685
R12737 VPWR VPWR.n2536 1.04685
R12738 VPWR.n2531 VPWR 1.04685
R12739 VPWR.n2511 VPWR 1.04685
R12740 VPWR VPWR.n462 1.04685
R12741 VPWR VPWR.n2663 1.04685
R12742 VPWR VPWR.n420 1.04685
R12743 VPWR.n2656 VPWR 1.04685
R12744 VPWR.n2649 VPWR 1.04685
R12745 VPWR.n2644 VPWR 1.04685
R12746 VPWR.n2518 VPWR 1.04685
R12747 VPWR VPWR.n2523 1.04685
R12748 VPWR.n2424 VPWR 1.04685
R12749 VPWR.n2429 VPWR 1.04685
R12750 VPWR.n2431 VPWR 1.04685
R12751 VPWR.n480 VPWR 1.04685
R12752 VPWR VPWR.n2444 1.04685
R12753 VPWR.n2439 VPWR 1.04685
R12754 VPWR.n2462 VPWR 1.04685
R12755 VPWR.n2467 VPWR 1.04685
R12756 VPWR.n2494 VPWR 1.04685
R12757 VPWR.n2490 VPWR 1.04685
R12758 VPWR.n2487 VPWR 1.04685
R12759 VPWR.n2482 VPWR 1.04685
R12760 VPWR.n2479 VPWR 1.04685
R12761 VPWR.n2474 VPWR 1.04685
R12762 VPWR.n2469 VPWR 1.04685
R12763 VPWR VPWR.n503 1.04685
R12764 VPWR VPWR.n2409 1.04685
R12765 VPWR.n2404 VPWR 1.04685
R12766 VPWR VPWR.n2402 1.04685
R12767 VPWR.n2397 VPWR 1.04685
R12768 VPWR VPWR.n2395 1.04685
R12769 VPWR.n2390 VPWR 1.04685
R12770 VPWR VPWR.n2388 1.04685
R12771 VPWR VPWR.n538 1.04685
R12772 VPWR.n2364 VPWR 1.04685
R12773 VPWR VPWR.n2369 1.04685
R12774 VPWR.n528 VPWR 1.04685
R12775 VPWR.n2376 VPWR 1.04685
R12776 VPWR VPWR.n2381 1.04685
R12777 VPWR.n2383 VPWR 1.04685
R12778 VPWR VPWR.n698 1.04685
R12779 VPWR.n693 VPWR 1.04685
R12780 VPWR.n563 VPWR 1.04685
R12781 VPWR VPWR.n2290 1.04685
R12782 VPWR.n2285 VPWR 1.04685
R12783 VPWR VPWR.n573 1.04685
R12784 VPWR VPWR.n556 1.04685
R12785 VPWR.n2309 VPWR 1.04685
R12786 VPWR.n2354 VPWR 1.04685
R12787 VPWR.n2350 VPWR 1.04685
R12788 VPWR VPWR.n544 1.04685
R12789 VPWR VPWR.n2323 1.04685
R12790 VPWR.n2325 VPWR 1.04685
R12791 VPWR VPWR.n2330 1.04685
R12792 VPWR.n553 VPWR 1.04685
R12793 VPWR VPWR.n682 1.04685
R12794 VPWR.n677 VPWR 1.04685
R12795 VPWR VPWR.n675 1.04685
R12796 VPWR.n670 VPWR 1.04685
R12797 VPWR.n666 VPWR 1.04685
R12798 VPWR VPWR.n664 1.04685
R12799 VPWR.n659 VPWR 1.04685
R12800 VPWR VPWR.n657 1.04685
R12801 VPWR.n2257 VPWR 1.04685
R12802 VPWR VPWR.n2261 1.04685
R12803 VPWR.n2263 VPWR 1.04685
R12804 VPWR VPWR.n2268 1.04685
R12805 VPWR VPWR.n578 1.04685
R12806 VPWR VPWR.n650 1.04685
R12807 VPWR.n652 VPWR 1.04685
R12808 VPWR.n2137 VPWR 1.04685
R12809 VPWR.n2145 VPWR 1.04685
R12810 VPWR VPWR.n616 1.04685
R12811 VPWR.n2154 VPWR 1.04685
R12812 VPWR.n2159 VPWR 1.04685
R12813 VPWR.n2166 VPWR 1.04685
R12814 VPWR.n2171 VPWR 1.04685
R12815 VPWR.n2178 VPWR 1.04685
R12816 VPWR.n2237 VPWR 1.04685
R12817 VPWR VPWR.n2241 1.04685
R12818 VPWR.n586 VPWR 1.04685
R12819 VPWR VPWR.n2191 1.04685
R12820 VPWR.n2193 VPWR 1.04685
R12821 VPWR VPWR.n2198 1.04685
R12822 VPWR VPWR.n605 1.04685
R12823 VPWR.n2076 VPWR 1.04685
R12824 VPWR.n2081 VPWR 1.04685
R12825 VPWR.n2084 VPWR 1.04685
R12826 VPWR VPWR.n2065 1.04685
R12827 VPWR VPWR.n2116 1.04685
R12828 VPWR.n2111 VPWR 1.04685
R12829 VPWR VPWR.n2109 1.04685
R12830 VPWR.n2104 VPWR 1.04685
R12831 VPWR VPWR.n2227 1.04685
R12832 VPWR VPWR.n594 1.04685
R12833 VPWR.n2220 VPWR 1.04685
R12834 VPWR.n2217 VPWR 1.04685
R12835 VPWR.n2212 VPWR 1.04685
R12836 VPWR.n2097 VPWR 1.04685
R12837 VPWR VPWR.n2102 1.04685
R12838 VPWR.n1931 VPWR 1.04685
R12839 VPWR VPWR.n761 1.04685
R12840 VPWR VPWR.n1946 1.04685
R12841 VPWR.n1941 VPWR 1.04685
R12842 VPWR.n712 VPWR 1.04685
R12843 VPWR VPWR.n2059 1.04685
R12844 VPWR.n2054 VPWR 1.04685
R12845 VPWR.n718 VPWR 1.04685
R12846 VPWR.n2024 VPWR 1.04685
R12847 VPWR VPWR.n2028 1.04685
R12848 VPWR.n730 VPWR 1.04685
R12849 VPWR.n2035 VPWR 1.04685
R12850 VPWR VPWR.n2040 1.04685
R12851 VPWR.n2042 VPWR 1.04685
R12852 VPWR VPWR.n2047 1.04685
R12853 VPWR VPWR.n792 1.04685
R12854 VPWR.n787 VPWR 1.04685
R12855 VPWR VPWR.n785 1.04685
R12856 VPWR.n780 VPWR 1.04685
R12857 VPWR VPWR.n778 1.04685
R12858 VPWR.n1961 VPWR 1.04685
R12859 VPWR.n1966 VPWR 1.04685
R12860 VPWR.n1969 VPWR 1.04685
R12861 VPWR.n1994 VPWR 1.04685
R12862 VPWR VPWR.n1998 1.04685
R12863 VPWR.n2000 VPWR 1.04685
R12864 VPWR VPWR.n2005 1.04685
R12865 VPWR VPWR.n744 1.04685
R12866 VPWR.n1985 VPWR 1.04685
R12867 VPWR.n1974 VPWR 1.04685
R12868 VPWR VPWR.n796 1.04685
R12869 VPWR VPWR.n1911 1.04685
R12870 VPWR.n1906 VPWR 1.04685
R12871 VPWR VPWR.n1904 1.04685
R12872 VPWR.n1899 VPWR 1.04685
R12873 VPWR.n817 VPWR 1.04685
R12874 VPWR VPWR.n812 1.04685
R12875 VPWR VPWR.n1891 1.04685
R12876 VPWR.n833 VPWR 1.04685
R12877 VPWR VPWR.n837 1.04685
R12878 VPWR.n1872 VPWR 1.04685
R12879 VPWR VPWR.n1877 1.04685
R12880 VPWR.n1879 VPWR 1.04685
R12881 VPWR VPWR.n1884 1.04685
R12882 VPWR.n1886 VPWR 1.04685
R12883 VPWR VPWR.n2549 1.04685
R12884 VPWR VPWR.n2566 1.04685
R12885 VPWR.n2561 VPWR 1.04685
R12886 VPWR.n2579 VPWR 1.04685
R12887 VPWR.n2584 VPWR 1.04685
R12888 VPWR.n2587 VPWR 1.04685
R12889 VPWR.n2602 VPWR 1.04685
R12890 VPWR VPWR.n2606 1.04685
R12891 VPWR.n2608 VPWR 1.04685
R12892 VPWR VPWR.n2613 1.04685
R12893 VPWR.n2615 VPWR 1.04685
R12894 VPWR VPWR.n2620 1.04685
R12895 VPWR.n2622 VPWR 1.04685
R12896 VPWR VPWR.n2627 1.04685
R12897 VPWR VPWR.n440 1.04685
R12898 VPWR.n1783 VPWR 1.04685
R12899 VPWR.n1785 VPWR 1.04685
R12900 VPWR.n867 VPWR 1.04685
R12901 VPWR VPWR.n1801 1.04685
R12902 VPWR.n1796 VPWR 1.04685
R12903 VPWR VPWR.n860 1.04685
R12904 VPWR.n1820 VPWR 1.04685
R12905 VPWR.n1825 VPWR 1.04685
R12906 VPWR.n1832 VPWR 1.04685
R12907 VPWR.n1840 VPWR 1.04685
R12908 VPWR.n1859 VPWR 1.04685
R12909 VPWR.n1855 VPWR 1.04685
R12910 VPWR.n1852 VPWR 1.04685
R12911 VPWR.n1847 VPWR 1.04685
R12912 VPWR VPWR.n846 1.04685
R12913 VPWR VPWR.n2734 1.04685
R12914 VPWR.n2729 VPWR 1.04685
R12915 VPWR.n380 VPWR 1.04685
R12916 VPWR VPWR.n2722 1.04685
R12917 VPWR.n2674 VPWR 1.04685
R12918 VPWR.n2681 VPWR 1.04685
R12919 VPWR VPWR.n2686 1.04685
R12920 VPWR.n407 VPWR 1.04685
R12921 VPWR.n2693 VPWR 1.04685
R12922 VPWR VPWR.n2698 1.04685
R12923 VPWR.n398 VPWR 1.04685
R12924 VPWR.n2705 VPWR 1.04685
R12925 VPWR VPWR.n2710 1.04685
R12926 VPWR.n389 VPWR 1.04685
R12927 VPWR.n2717 VPWR 1.04685
R12928 VPWR.n875 VPWR 1.04685
R12929 VPWR VPWR.n1769 1.04685
R12930 VPWR.n1764 VPWR 1.04685
R12931 VPWR VPWR.n1762 1.04685
R12932 VPWR.n1757 VPWR 1.04685
R12933 VPWR.n898 VPWR 1.04685
R12934 VPWR VPWR.n893 1.04685
R12935 VPWR VPWR.n1749 1.04685
R12936 VPWR.n1744 VPWR 1.04685
R12937 VPWR VPWR.n1742 1.04685
R12938 VPWR.n1737 VPWR 1.04685
R12939 VPWR VPWR.n1735 1.04685
R12940 VPWR VPWR.n1723 1.04685
R12941 VPWR.n1716 VPWR 1.04685
R12942 VPWR.n1730 VPWR 1.04685
R12943 VPWR.n1194 VPWR 1.04685
R12944 VPWR.n1197 VPWR 1.04685
R12945 VPWR VPWR.n1171 1.04685
R12946 VPWR VPWR.n1661 1.04685
R12947 VPWR.n1656 VPWR 1.04685
R12948 VPWR VPWR.n1654 1.04685
R12949 VPWR.n1649 VPWR 1.04685
R12950 VPWR VPWR.n1647 1.04685
R12951 VPWR.n1642 VPWR 1.04685
R12952 VPWR.n1232 VPWR 1.04685
R12953 VPWR VPWR.n1634 1.04685
R12954 VPWR VPWR.n929 1.04685
R12955 VPWR.n1703 VPWR 1.04685
R12956 VPWR VPWR.n1713 1.04685
R12957 VPWR VPWR.n919 1.04685
R12958 VPWR VPWR.n367 1.04685
R12959 VPWR.n362 VPWR 1.04685
R12960 VPWR VPWR.n318 1.04685
R12961 VPWR.n320 VPWR 1.04685
R12962 VPWR VPWR.n325 1.04685
R12963 VPWR.n327 VPWR 1.04685
R12964 VPWR VPWR.n332 1.04685
R12965 VPWR.n334 VPWR 1.04685
R12966 VPWR VPWR.n339 1.04685
R12967 VPWR.n341 VPWR 1.04685
R12968 VPWR VPWR.n346 1.04685
R12969 VPWR.n348 VPWR 1.04685
R12970 VPWR VPWR.n353 1.04685
R12971 VPWR.n355 VPWR 1.04685
R12972 VPWR VPWR.n360 1.04685
R12973 VPWR VPWR.n84 1.04524
R12974 VPWR VPWR.n81 1.04524
R12975 VPWR VPWR.n78 1.04524
R12976 VPWR VPWR.n75 1.04524
R12977 VPWR VPWR.n72 1.04524
R12978 VPWR VPWR.n69 1.04524
R12979 VPWR VPWR.n66 1.04524
R12980 VPWR VPWR.n63 1.04524
R12981 VPWR VPWR.n60 1.04524
R12982 VPWR VPWR.n57 1.04524
R12983 VPWR VPWR.n54 1.04524
R12984 VPWR VPWR.n51 1.04524
R12985 VPWR VPWR.n48 1.04524
R12986 VPWR VPWR.n45 1.04524
R12987 VPWR VPWR.n42 1.04524
R12988 VPWR.n1585 VPWR 1.04524
R12989 VPWR VPWR.n1591 1.04524
R12990 VPWR VPWR.n1246 1.04524
R12991 VPWR.n1247 VPWR 1.04524
R12992 VPWR.n1535 VPWR 1.04524
R12993 VPWR.n1519 VPWR 1.04524
R12994 VPWR VPWR.n1259 1.04524
R12995 VPWR VPWR.n1262 1.04524
R12996 VPWR VPWR.n1264 1.04524
R12997 VPWR VPWR.n1267 1.04524
R12998 VPWR VPWR.n1269 1.04524
R12999 VPWR.n1415 VPWR 1.04524
R13000 VPWR.n1281 VPWR 1.04524
R13001 VPWR.n1165 VPWR 1.04524
R13002 VPWR VPWR.n1675 1.04524
R13003 VPWR VPWR.n42 0.900028
R13004 VPWR.n1585 VPWR 0.900028
R13005 VPWR.n1297 VPWR.n1157 0.880079
R13006 VPWR.n2760 VPWR.n290 0.880079
R13007 VPWR.n1591 VPWR.n1236 0.878476
R13008 VPWR.n1566 VPWR.n1246 0.878476
R13009 VPWR.n1554 VPWR.n1247 0.878476
R13010 VPWR.n1539 VPWR.n1535 0.878476
R13011 VPWR.n1519 VPWR.n1258 0.878476
R13012 VPWR.n1359 VPWR.n1259 0.878476
R13013 VPWR.n1370 VPWR.n1262 0.878476
R13014 VPWR.n1381 VPWR.n1264 0.878476
R13015 VPWR.n1392 VPWR.n1267 0.878476
R13016 VPWR.n1403 VPWR.n1269 0.878476
R13017 VPWR.n1415 VPWR.n1414 0.878476
R13018 VPWR.n1329 VPWR.n1281 0.878476
R13019 VPWR.n1317 VPWR.n1165 0.878476
R13020 VPWR.n1675 VPWR.n1158 0.878476
R13021 VPWR.n271 VPWR.n84 0.878476
R13022 VPWR.n268 VPWR.n81 0.878476
R13023 VPWR.n256 VPWR.n78 0.878476
R13024 VPWR.n237 VPWR.n75 0.878476
R13025 VPWR.n234 VPWR.n72 0.878476
R13026 VPWR.n222 VPWR.n69 0.878476
R13027 VPWR.n203 VPWR.n66 0.878476
R13028 VPWR.n200 VPWR.n63 0.878476
R13029 VPWR.n188 VPWR.n60 0.878476
R13030 VPWR.n169 VPWR.n57 0.878476
R13031 VPWR.n166 VPWR.n54 0.878476
R13032 VPWR.n154 VPWR.n51 0.878476
R13033 VPWR.n135 VPWR.n48 0.878476
R13034 VPWR.n132 VPWR.n45 0.878476
R13035 VPWR.n3126 VPWR.n3125 0.711611
R13036 VPWR.n34 VPWR.n33 0.711611
R13037 VPWR.n1299 VPWR.n1297 0.675548
R13038 VPWR.n1283 VPWR.n1158 0.675548
R13039 VPWR.n1319 VPWR.n1317 0.675548
R13040 VPWR.n1331 VPWR.n1329 0.675548
R13041 VPWR.n1414 VPWR.n1413 0.675548
R13042 VPWR.n1403 VPWR.n1402 0.675548
R13043 VPWR.n1392 VPWR.n1391 0.675548
R13044 VPWR.n1381 VPWR.n1380 0.675548
R13045 VPWR.n1370 VPWR.n1369 0.675548
R13046 VPWR.n1359 VPWR.n1358 0.675548
R13047 VPWR.n1258 VPWR.n1257 0.675548
R13048 VPWR.n1539 VPWR.n1538 0.675548
R13049 VPWR.n1556 VPWR.n1554 0.675548
R13050 VPWR.n1568 VPWR.n1566 0.675548
R13051 VPWR.n1241 VPWR.n1236 0.675548
R13052 VPWR.n132 VPWR.n131 0.675548
R13053 VPWR.n137 VPWR.n135 0.675548
R13054 VPWR.n154 VPWR.n153 0.675548
R13055 VPWR.n166 VPWR.n165 0.675548
R13056 VPWR.n171 VPWR.n169 0.675548
R13057 VPWR.n188 VPWR.n187 0.675548
R13058 VPWR.n200 VPWR.n199 0.675548
R13059 VPWR.n205 VPWR.n203 0.675548
R13060 VPWR.n222 VPWR.n221 0.675548
R13061 VPWR.n234 VPWR.n233 0.675548
R13062 VPWR.n239 VPWR.n237 0.675548
R13063 VPWR.n256 VPWR.n255 0.675548
R13064 VPWR.n268 VPWR.n267 0.675548
R13065 VPWR.n273 VPWR.n271 0.675548
R13066 VPWR.n290 VPWR.n289 0.675548
R13067 VPWR.n3095 VPWR.n3094 0.672385
R13068 VPWR.n3079 VPWR.n3074 0.672385
R13069 VPWR.n3059 VPWR.n3054 0.672385
R13070 VPWR.n3040 VPWR.n3035 0.672385
R13071 VPWR.n3116 VPWR.n36 0.654518
R13072 VPWR.n7 VPWR 0.63497
R13073 VPWR.n950 VPWR 0.63497
R13074 VPWR.n973 VPWR 0.63497
R13075 VPWR.n997 VPWR 0.63497
R13076 VPWR.n3122 VPWR.n26 0.573634
R13077 VPWR.n3118 VPWR.n3117 0.573634
R13078 VPWR VPWR.n3131 0.541783
R13079 VPWR.n2851 VPWR 0.499542
R13080 VPWR.n3130 VPWR.n21 0.498268
R13081 VPWR.n3128 VPWR.n3127 0.493804
R13082 VPWR.n1296 VPWR.n1294 0.404056
R13083 VPWR.n1305 VPWR.n1304 0.404056
R13084 VPWR.n1316 VPWR.n1314 0.404056
R13085 VPWR.n1328 VPWR.n1326 0.404056
R13086 VPWR.n1337 VPWR.n1336 0.404056
R13087 VPWR.n1408 VPWR.n1405 0.404056
R13088 VPWR.n1397 VPWR.n1394 0.404056
R13089 VPWR.n1386 VPWR.n1383 0.404056
R13090 VPWR.n1375 VPWR.n1372 0.404056
R13091 VPWR.n1364 VPWR.n1361 0.404056
R13092 VPWR.n1353 VPWR.n1350 0.404056
R13093 VPWR.n1542 VPWR.n1541 0.404056
R13094 VPWR.n1553 VPWR.n1551 0.404056
R13095 VPWR.n1565 VPWR.n1563 0.404056
R13096 VPWR.n1574 VPWR.n1573 0.404056
R13097 VPWR.n1584 VPWR.n1582 0.404056
R13098 VPWR.n97 VPWR.n92 0.404056
R13099 VPWR.n126 VPWR.n123 0.404056
R13100 VPWR.n141 VPWR.n134 0.404056
R13101 VPWR.n148 VPWR.n118 0.404056
R13102 VPWR.n160 VPWR.n156 0.404056
R13103 VPWR.n175 VPWR.n168 0.404056
R13104 VPWR.n182 VPWR.n113 0.404056
R13105 VPWR.n194 VPWR.n190 0.404056
R13106 VPWR.n209 VPWR.n202 0.404056
R13107 VPWR.n216 VPWR.n108 0.404056
R13108 VPWR.n228 VPWR.n224 0.404056
R13109 VPWR.n243 VPWR.n236 0.404056
R13110 VPWR.n250 VPWR.n103 0.404056
R13111 VPWR.n262 VPWR.n258 0.404056
R13112 VPWR.n277 VPWR.n270 0.404056
R13113 VPWR.n284 VPWR.n88 0.404056
R13114 VPWR.n1578 VPWR.n1245 0.349144
R13115 VPWR.n1547 VPWR.n1245 0.349144
R13116 VPWR.n1547 VPWR.n1546 0.349144
R13117 VPWR.n1546 VPWR.n1250 0.349144
R13118 VPWR.n1346 VPWR.n1250 0.349144
R13119 VPWR.n1346 VPWR.n1345 0.349144
R13120 VPWR.n1345 VPWR.n1344 0.349144
R13121 VPWR.n1344 VPWR.n1343 0.349144
R13122 VPWR.n1343 VPWR.n1342 0.349144
R13123 VPWR.n1342 VPWR.n1341 0.349144
R13124 VPWR.n1341 VPWR.n1276 0.349144
R13125 VPWR.n1310 VPWR.n1276 0.349144
R13126 VPWR.n1310 VPWR.n1309 0.349144
R13127 VPWR.n282 VPWR.n281 0.349144
R13128 VPWR.n281 VPWR.n101 0.349144
R13129 VPWR.n248 VPWR.n101 0.349144
R13130 VPWR.n248 VPWR.n247 0.349144
R13131 VPWR.n247 VPWR.n106 0.349144
R13132 VPWR.n214 VPWR.n106 0.349144
R13133 VPWR.n214 VPWR.n213 0.349144
R13134 VPWR.n213 VPWR.n111 0.349144
R13135 VPWR.n180 VPWR.n111 0.349144
R13136 VPWR.n180 VPWR.n179 0.349144
R13137 VPWR.n179 VPWR.n116 0.349144
R13138 VPWR.n146 VPWR.n116 0.349144
R13139 VPWR.n146 VPWR.n145 0.349144
R13140 VPWR.n1427 VPWR.n1423 0.346131
R13141 VPWR.n1433 VPWR.n1421 0.346131
R13142 VPWR.n1694 VPWR.n1690 0.346131
R13143 VPWR.n1695 VPWR.n936 0.346131
R13144 VPWR.n1605 VPWR.n932 0.346131
R13145 VPWR.n1610 VPWR.n1606 0.346131
R13146 VPWR.n1611 VPWR.n1601 0.346131
R13147 VPWR.n1466 VPWR.n1230 0.346131
R13148 VPWR.n1471 VPWR.n1467 0.346131
R13149 VPWR.n1472 VPWR.n1462 0.346131
R13150 VPWR.n1458 VPWR.n1457 0.346131
R13151 VPWR.n1453 VPWR.n1452 0.346131
R13152 VPWR.n1448 VPWR.n1447 0.346131
R13153 VPWR.n1443 VPWR.n1442 0.346131
R13154 VPWR.n1438 VPWR.n1437 0.346131
R13155 VPWR.n2883 VPWR.n2882 0.300179
R13156 VPWR.n3103 VPWR.n38 0.298167
R13157 VPWR.n1294 VPWR.n1293 0.286958
R13158 VPWR.n1306 VPWR.n1305 0.286958
R13159 VPWR.n1314 VPWR.n1313 0.286958
R13160 VPWR.n1326 VPWR.n1325 0.286958
R13161 VPWR.n1338 VPWR.n1337 0.286958
R13162 VPWR.n1408 VPWR.n1407 0.286958
R13163 VPWR.n1397 VPWR.n1396 0.286958
R13164 VPWR.n1386 VPWR.n1385 0.286958
R13165 VPWR.n1375 VPWR.n1374 0.286958
R13166 VPWR.n1364 VPWR.n1363 0.286958
R13167 VPWR.n1353 VPWR.n1352 0.286958
R13168 VPWR.n1543 VPWR.n1542 0.286958
R13169 VPWR.n1551 VPWR.n1550 0.286958
R13170 VPWR.n1563 VPWR.n1562 0.286958
R13171 VPWR.n1575 VPWR.n1574 0.286958
R13172 VPWR.n1582 VPWR.n1581 0.286958
R13173 VPWR.n98 VPWR.n97 0.286958
R13174 VPWR.n126 VPWR.n125 0.286958
R13175 VPWR.n142 VPWR.n141 0.286958
R13176 VPWR.n148 VPWR.n119 0.286958
R13177 VPWR.n160 VPWR.n157 0.286958
R13178 VPWR.n176 VPWR.n175 0.286958
R13179 VPWR.n182 VPWR.n114 0.286958
R13180 VPWR.n194 VPWR.n191 0.286958
R13181 VPWR.n210 VPWR.n209 0.286958
R13182 VPWR.n216 VPWR.n109 0.286958
R13183 VPWR.n228 VPWR.n225 0.286958
R13184 VPWR.n244 VPWR.n243 0.286958
R13185 VPWR.n250 VPWR.n104 0.286958
R13186 VPWR.n262 VPWR.n259 0.286958
R13187 VPWR.n278 VPWR.n277 0.286958
R13188 VPWR.n284 VPWR.n89 0.286958
R13189 VPWR.n2882 VPWR 0.2505
R13190 VPWR VPWR.n2754 0.249238
R13191 VPWR VPWR.n2753 0.249238
R13192 VPWR VPWR.n2752 0.249238
R13193 VPWR VPWR.n2751 0.249238
R13194 VPWR VPWR.n2737 0.249238
R13195 VPWR.n2568 VPWR 0.249238
R13196 VPWR.n2726 VPWR 0.249238
R13197 VPWR VPWR.n2725 0.249238
R13198 VPWR.n447 VPWR 0.249238
R13199 VPWR.n2714 VPWR 0.249238
R13200 VPWR.n449 VPWR 0.249238
R13201 VPWR.n2571 VPWR 0.249238
R13202 VPWR.n2572 VPWR 0.249238
R13203 VPWR.n2573 VPWR 0.249238
R13204 VPWR.n2576 VPWR 0.249238
R13205 VPWR VPWR.n2575 0.249238
R13206 VPWR VPWR.n2574 0.249238
R13207 VPWR.n2630 VPWR 0.249238
R13208 VPWR VPWR.n2415 0.249238
R13209 VPWR.n2547 VPWR 0.249238
R13210 VPWR VPWR.n2546 0.249238
R13211 VPWR.n2451 VPWR 0.249238
R13212 VPWR.n2452 VPWR 0.249238
R13213 VPWR.n2453 VPWR 0.249238
R13214 VPWR.n2528 VPWR 0.249238
R13215 VPWR VPWR.n2527 0.249238
R13216 VPWR VPWR.n2526 0.249238
R13217 VPWR.n2667 VPWR 0.249238
R13218 VPWR.n2666 VPWR 0.249238
R13219 VPWR.n2653 VPWR 0.249238
R13220 VPWR.n2652 VPWR 0.249238
R13221 VPWR.n2641 VPWR 0.249238
R13222 VPWR.n2640 VPWR 0.249238
R13223 VPWR.n2505 VPWR 0.249238
R13224 VPWR.n2420 VPWR 0.249238
R13225 VPWR VPWR.n2419 0.249238
R13226 VPWR VPWR.n2418 0.249238
R13227 VPWR.n2448 VPWR 0.249238
R13228 VPWR VPWR.n2447 0.249238
R13229 VPWR.n2456 VPWR 0.249238
R13230 VPWR.n2457 VPWR 0.249238
R13231 VPWR.n2459 VPWR 0.249238
R13232 VPWR VPWR.n2458 0.249238
R13233 VPWR VPWR.n2497 0.249238
R13234 VPWR VPWR.n2498 0.249238
R13235 VPWR VPWR.n2499 0.249238
R13236 VPWR VPWR.n2500 0.249238
R13237 VPWR VPWR.n2501 0.249238
R13238 VPWR VPWR.n2502 0.249238
R13239 VPWR.n2503 VPWR 0.249238
R13240 VPWR VPWR.n2413 0.249238
R13241 VPWR VPWR.n2412 0.249238
R13242 VPWR.n2297 VPWR 0.249238
R13243 VPWR.n2298 VPWR 0.249238
R13244 VPWR.n2299 VPWR 0.249238
R13245 VPWR.n2300 VPWR 0.249238
R13246 VPWR.n2302 VPWR 0.249238
R13247 VPWR VPWR.n2301 0.249238
R13248 VPWR.n2337 VPWR 0.249238
R13249 VPWR VPWR.n2360 0.249238
R13250 VPWR.n2361 VPWR 0.249238
R13251 VPWR.n546 VPWR 0.249238
R13252 VPWR VPWR.n2372 0.249238
R13253 VPWR.n2373 VPWR 0.249238
R13254 VPWR.n2339 VPWR 0.249238
R13255 VPWR.n2338 VPWR 0.249238
R13256 VPWR.n701 VPWR 0.249238
R13257 VPWR VPWR.n700 0.249238
R13258 VPWR.n2294 VPWR 0.249238
R13259 VPWR VPWR.n2293 0.249238
R13260 VPWR.n2281 VPWR 0.249238
R13261 VPWR.n2282 VPWR 0.249238
R13262 VPWR.n2305 VPWR 0.249238
R13263 VPWR.n2306 VPWR 0.249238
R13264 VPWR.n2334 VPWR 0.249238
R13265 VPWR.n2357 VPWR 0.249238
R13266 VPWR VPWR.n2345 0.249238
R13267 VPWR.n2346 VPWR 0.249238
R13268 VPWR.n2344 VPWR 0.249238
R13269 VPWR.n2343 VPWR 0.249238
R13270 VPWR.n2342 VPWR 0.249238
R13271 VPWR VPWR.n2333 0.249238
R13272 VPWR.n2130 VPWR 0.249238
R13273 VPWR VPWR.n2129 0.249238
R13274 VPWR VPWR.n2128 0.249238
R13275 VPWR VPWR.n2127 0.249238
R13276 VPWR.n2278 VPWR 0.249238
R13277 VPWR VPWR.n2277 0.249238
R13278 VPWR VPWR.n2276 0.249238
R13279 VPWR VPWR.n2275 0.249238
R13280 VPWR VPWR.n2274 0.249238
R13281 VPWR VPWR.n2250 0.249238
R13282 VPWR.n2251 VPWR 0.249238
R13283 VPWR.n2249 VPWR 0.249238
R13284 VPWR.n2248 VPWR 0.249238
R13285 VPWR VPWR.n2271 0.249238
R13286 VPWR VPWR.n2272 0.249238
R13287 VPWR VPWR.n2273 0.249238
R13288 VPWR.n2133 VPWR 0.249238
R13289 VPWR.n2134 VPWR 0.249238
R13290 VPWR.n2148 VPWR 0.249238
R13291 VPWR.n2150 VPWR 0.249238
R13292 VPWR VPWR.n2149 0.249238
R13293 VPWR.n2162 VPWR 0.249238
R13294 VPWR.n2163 VPWR 0.249238
R13295 VPWR.n2174 VPWR 0.249238
R13296 VPWR.n2175 VPWR 0.249238
R13297 VPWR.n2234 VPWR 0.249238
R13298 VPWR.n591 VPWR 0.249238
R13299 VPWR VPWR.n2244 0.249238
R13300 VPWR.n2245 VPWR 0.249238
R13301 VPWR VPWR.n2202 0.249238
R13302 VPWR.n2203 VPWR 0.249238
R13303 VPWR.n2201 VPWR 0.249238
R13304 VPWR VPWR.n2123 0.249238
R13305 VPWR VPWR.n2122 0.249238
R13306 VPWR VPWR.n2121 0.249238
R13307 VPWR VPWR.n2120 0.249238
R13308 VPWR VPWR.n2119 0.249238
R13309 VPWR VPWR.n708 0.249238
R13310 VPWR VPWR.n707 0.249238
R13311 VPWR VPWR.n706 0.249238
R13312 VPWR VPWR.n705 0.249238
R13313 VPWR.n2231 VPWR 0.249238
R13314 VPWR.n2230 VPWR 0.249238
R13315 VPWR VPWR.n2207 0.249238
R13316 VPWR VPWR.n2208 0.249238
R13317 VPWR.n2209 VPWR 0.249238
R13318 VPWR.n2206 VPWR 0.249238
R13319 VPWR VPWR.n704 0.249238
R13320 VPWR.n1927 VPWR 0.249238
R13321 VPWR.n1928 VPWR 0.249238
R13322 VPWR.n1949 VPWR 0.249238
R13323 VPWR.n1950 VPWR 0.249238
R13324 VPWR.n2063 VPWR 0.249238
R13325 VPWR VPWR.n2062 0.249238
R13326 VPWR.n755 VPWR 0.249238
R13327 VPWR.n2051 VPWR 0.249238
R13328 VPWR VPWR.n2050 0.249238
R13329 VPWR.n2021 VPWR 0.249238
R13330 VPWR.n2020 VPWR 0.249238
R13331 VPWR VPWR.n2031 0.249238
R13332 VPWR.n2032 VPWR 0.249238
R13333 VPWR VPWR.n1976 0.249238
R13334 VPWR VPWR.n1977 0.249238
R13335 VPWR.n1978 VPWR 0.249238
R13336 VPWR.n1920 VPWR 0.249238
R13337 VPWR VPWR.n1919 0.249238
R13338 VPWR VPWR.n1918 0.249238
R13339 VPWR.n1953 VPWR 0.249238
R13340 VPWR.n1954 VPWR 0.249238
R13341 VPWR.n1955 VPWR 0.249238
R13342 VPWR.n1958 VPWR 0.249238
R13343 VPWR VPWR.n1957 0.249238
R13344 VPWR VPWR.n1956 0.249238
R13345 VPWR.n2018 VPWR 0.249238
R13346 VPWR.n2011 VPWR 0.249238
R13347 VPWR.n2010 VPWR 0.249238
R13348 VPWR.n2009 VPWR 0.249238
R13349 VPWR.n2008 VPWR 0.249238
R13350 VPWR.n1982 VPWR 0.249238
R13351 VPWR.n1981 VPWR 0.249238
R13352 VPWR VPWR.n1915 0.249238
R13353 VPWR VPWR.n1914 0.249238
R13354 VPWR.n1808 VPWR 0.249238
R13355 VPWR.n1809 VPWR 0.249238
R13356 VPWR.n1810 VPWR 0.249238
R13357 VPWR.n1896 VPWR 0.249238
R13358 VPWR VPWR.n1895 0.249238
R13359 VPWR VPWR.n1894 0.249238
R13360 VPWR.n856 VPWR 0.249238
R13361 VPWR.n2015 VPWR 0.249238
R13362 VPWR.n2014 VPWR 0.249238
R13363 VPWR.n1869 VPWR 0.249238
R13364 VPWR.n1868 VPWR 0.249238
R13365 VPWR VPWR.n853 0.249238
R13366 VPWR VPWR.n854 0.249238
R13367 VPWR VPWR.n855 0.249238
R13368 VPWR.n2670 VPWR 0.249238
R13369 VPWR VPWR.n2633 0.249238
R13370 VPWR VPWR.n2634 0.249238
R13371 VPWR VPWR.n2635 0.249238
R13372 VPWR VPWR.n2636 0.249238
R13373 VPWR.n2637 VPWR 0.249238
R13374 VPWR.n2632 VPWR 0.249238
R13375 VPWR.n2631 VPWR 0.249238
R13376 VPWR.n1776 VPWR 0.249238
R13377 VPWR VPWR.n1775 0.249238
R13378 VPWR.n1805 VPWR 0.249238
R13379 VPWR VPWR.n1804 0.249238
R13380 VPWR.n1813 VPWR 0.249238
R13381 VPWR.n1814 VPWR 0.249238
R13382 VPWR.n1816 VPWR 0.249238
R13383 VPWR VPWR.n1815 0.249238
R13384 VPWR.n1828 VPWR 0.249238
R13385 VPWR.n1829 VPWR 0.249238
R13386 VPWR VPWR.n1862 0.249238
R13387 VPWR VPWR.n1863 0.249238
R13388 VPWR VPWR.n1864 0.249238
R13389 VPWR.n1865 VPWR 0.249238
R13390 VPWR.n1844 VPWR 0.249238
R13391 VPWR.n1843 VPWR 0.249238
R13392 VPWR VPWR.n2677 0.249238
R13393 VPWR.n2678 VPWR 0.249238
R13394 VPWR.n425 VPWR 0.249238
R13395 VPWR VPWR.n2689 0.249238
R13396 VPWR.n2690 VPWR 0.249238
R13397 VPWR.n435 VPWR 0.249238
R13398 VPWR VPWR.n2701 0.249238
R13399 VPWR.n2702 VPWR 0.249238
R13400 VPWR.n438 VPWR 0.249238
R13401 VPWR VPWR.n2713 0.249238
R13402 VPWR.n1773 VPWR 0.249238
R13403 VPWR VPWR.n1772 0.249238
R13404 VPWR.n889 VPWR 0.249238
R13405 VPWR.n890 VPWR 0.249238
R13406 VPWR.n891 VPWR 0.249238
R13407 VPWR.n1754 VPWR 0.249238
R13408 VPWR VPWR.n1753 0.249238
R13409 VPWR VPWR.n1752 0.249238
R13410 VPWR.n912 VPWR 0.249238
R13411 VPWR.n913 VPWR 0.249238
R13412 VPWR.n914 VPWR 0.249238
R13413 VPWR.n915 VPWR 0.249238
R13414 VPWR.n937 VPWR 0.249238
R13415 VPWR VPWR.n1726 0.249238
R13416 VPWR.n1727 VPWR 0.249238
R13417 VPWR.n916 VPWR 0.249238
R13418 VPWR VPWR.n2739 0.249238
R13419 VPWR VPWR.n2740 0.249238
R13420 VPWR VPWR.n2741 0.249238
R13421 VPWR VPWR.n2742 0.249238
R13422 VPWR VPWR.n2743 0.249238
R13423 VPWR VPWR.n2744 0.249238
R13424 VPWR VPWR.n2745 0.249238
R13425 VPWR VPWR.n2746 0.249238
R13426 VPWR VPWR.n2747 0.249238
R13427 VPWR VPWR.n2748 0.249238
R13428 VPWR VPWR.n2749 0.249238
R13429 VPWR VPWR.n2750 0.249238
R13430 VPWR.n2757 VPWR 0.249238
R13431 VPWR.n2768 VPWR 0.249238
R13432 VPWR.n2769 VPWR 0.249238
R13433 VPWR.n2780 VPWR 0.249238
R13434 VPWR.n2781 VPWR 0.249238
R13435 VPWR.n2792 VPWR 0.249238
R13436 VPWR.n2793 VPWR 0.249238
R13437 VPWR.n2804 VPWR 0.249238
R13438 VPWR.n2805 VPWR 0.249238
R13439 VPWR.n2816 VPWR 0.249238
R13440 VPWR.n2817 VPWR 0.249238
R13441 VPWR.n2828 VPWR 0.249238
R13442 VPWR.n2829 VPWR 0.249238
R13443 VPWR.n2840 VPWR 0.249238
R13444 VPWR.n2841 VPWR 0.249238
R13445 VPWR.n2884 VPWR 0.249238
R13446 VPWR.n1682 VPWR 0.249238
R13447 VPWR VPWR.n1234 0.249238
R13448 VPWR VPWR.n1594 0.249238
R13449 VPWR VPWR.n1595 0.249238
R13450 VPWR.n1596 VPWR 0.249238
R13451 VPWR VPWR.n1507 0.249238
R13452 VPWR VPWR.n1508 0.249238
R13453 VPWR.n1509 VPWR 0.249238
R13454 VPWR.n1506 VPWR 0.249238
R13455 VPWR.n1495 VPWR 0.249238
R13456 VPWR.n1494 VPWR 0.249238
R13457 VPWR.n1483 VPWR 0.249238
R13458 VPWR VPWR.n1665 0.249238
R13459 VPWR.n1666 VPWR 0.249238
R13460 VPWR.n1168 VPWR 0.249238
R13461 VPWR VPWR.n1678 0.249238
R13462 VPWR.n36 VPWR.n22 0.242688
R13463 VPWR.n3102 VPWR.n3086 0.213567
R13464 VPWR.n3086 VPWR.n3067 0.213567
R13465 VPWR.n3067 VPWR.n3047 0.213567
R13466 VPWR.n3047 VPWR.n3028 0.213567
R13467 VPWR.n3028 VPWR.n2992 0.213567
R13468 VPWR.n2992 VPWR.n2954 0.213567
R13469 VPWR.n2954 VPWR.n2917 0.213567
R13470 VPWR.n1154 VPWR.n1122 0.213567
R13471 VPWR.n1122 VPWR.n1084 0.213567
R13472 VPWR.n1084 VPWR.n1045 0.213567
R13473 VPWR.n1045 VPWR.n1010 0.213567
R13474 VPWR.n1010 VPWR.n987 0.213567
R13475 VPWR.n987 VPWR.n963 0.213567
R13476 VPWR.n963 VPWR.n19 0.213567
R13477 VPWR.n3116 VPWR.n3115 0.189116
R13478 VPWR.n3131 VPWR.n20 0.182233
R13479 VPWR.n1680 VPWR.n1679 0.179202
R13480 VPWR.n1679 VPWR.n1156 0.154425
R13481 VPWR.n1156 VPWR.n1155 0.154425
R13482 VPWR.n1155 VPWR.n794 0.154425
R13483 VPWR.n1916 VPWR.n794 0.154425
R13484 VPWR.n1917 VPWR.n1916 0.154425
R13485 VPWR.n1917 VPWR.n703 0.154425
R13486 VPWR.n2124 VPWR.n703 0.154425
R13487 VPWR.n2125 VPWR.n2124 0.154425
R13488 VPWR.n2126 VPWR.n2125 0.154425
R13489 VPWR.n2126 VPWR.n501 0.154425
R13490 VPWR.n2414 VPWR.n501 0.154425
R13491 VPWR.n2417 VPWR.n2414 0.154425
R13492 VPWR.n2417 VPWR.n2416 0.154425
R13493 VPWR.n2416 VPWR.n370 0.154425
R13494 VPWR.n2738 VPWR.n370 0.154425
R13495 VPWR.n2755 VPWR.n2738 0.154425
R13496 VPWR.n2756 VPWR.n2755 0.154425
R13497 VPWR.n1681 VPWR.n939 0.154425
R13498 VPWR.n939 VPWR.n938 0.154425
R13499 VPWR.n938 VPWR.n739 0.154425
R13500 VPWR.n2016 VPWR.n739 0.154425
R13501 VPWR.n2017 VPWR.n2016 0.154425
R13502 VPWR.n2017 VPWR.n592 0.154425
R13503 VPWR.n2232 VPWR.n592 0.154425
R13504 VPWR.n2233 VPWR.n2232 0.154425
R13505 VPWR.n2233 VPWR.n540 0.154425
R13506 VPWR.n2358 VPWR.n540 0.154425
R13507 VPWR.n2359 VPWR.n2358 0.154425
R13508 VPWR.n2359 VPWR.n418 0.154425
R13509 VPWR.n2668 VPWR.n418 0.154425
R13510 VPWR.n2669 VPWR.n2668 0.154425
R13511 VPWR.n2669 VPWR.n415 0.154425
R13512 VPWR.n415 VPWR.n40 0.154425
R13513 VPWR.n2885 VPWR.n40 0.154425
R13514 VPWR.n8 VPWR.n7 0.147771
R13515 VPWR.n951 VPWR.n950 0.147771
R13516 VPWR.n974 VPWR.n973 0.147771
R13517 VPWR.n998 VPWR.n997 0.147771
R13518 VPWR.n3103 VPWR.n3102 0.145025
R13519 VPWR.n1293 VPWR 0.135917
R13520 VPWR.n1306 VPWR 0.135917
R13521 VPWR.n1313 VPWR 0.135917
R13522 VPWR.n1325 VPWR 0.135917
R13523 VPWR.n1338 VPWR 0.135917
R13524 VPWR.n1407 VPWR 0.135917
R13525 VPWR.n1396 VPWR 0.135917
R13526 VPWR.n1385 VPWR 0.135917
R13527 VPWR.n1374 VPWR 0.135917
R13528 VPWR.n1363 VPWR 0.135917
R13529 VPWR.n1352 VPWR 0.135917
R13530 VPWR.n1543 VPWR 0.135917
R13531 VPWR.n1550 VPWR 0.135917
R13532 VPWR.n1562 VPWR 0.135917
R13533 VPWR.n1575 VPWR 0.135917
R13534 VPWR.n1581 VPWR 0.135917
R13535 VPWR.n98 VPWR 0.135917
R13536 VPWR.n125 VPWR 0.135917
R13537 VPWR.n142 VPWR 0.135917
R13538 VPWR.n119 VPWR 0.135917
R13539 VPWR.n157 VPWR 0.135917
R13540 VPWR.n176 VPWR 0.135917
R13541 VPWR.n114 VPWR 0.135917
R13542 VPWR.n191 VPWR 0.135917
R13543 VPWR.n210 VPWR 0.135917
R13544 VPWR.n109 VPWR 0.135917
R13545 VPWR.n225 VPWR 0.135917
R13546 VPWR.n244 VPWR 0.135917
R13547 VPWR.n104 VPWR 0.135917
R13548 VPWR.n259 VPWR 0.135917
R13549 VPWR.n278 VPWR 0.135917
R13550 VPWR.n89 VPWR 0.135917
R13551 VPWR.n38 VPWR.n37 0.123287
R13552 VPWR.n18 VPWR.n0 0.120292
R13553 VPWR.n14 VPWR.n0 0.120292
R13554 VPWR.n9 VPWR.n8 0.120292
R13555 VPWR.n962 VPWR.n941 0.120292
R13556 VPWR.n958 VPWR.n941 0.120292
R13557 VPWR.n952 VPWR.n951 0.120292
R13558 VPWR.n986 VPWR.n964 0.120292
R13559 VPWR.n981 VPWR.n964 0.120292
R13560 VPWR.n975 VPWR.n974 0.120292
R13561 VPWR.n1009 VPWR.n988 0.120292
R13562 VPWR.n1005 VPWR.n988 0.120292
R13563 VPWR.n999 VPWR.n998 0.120292
R13564 VPWR.n1041 VPWR.n1040 0.120292
R13565 VPWR.n1034 VPWR.n1013 0.120292
R13566 VPWR.n1027 VPWR.n1013 0.120292
R13567 VPWR.n1027 VPWR.n1026 0.120292
R13568 VPWR.n1025 VPWR.n1017 0.120292
R13569 VPWR.n1020 VPWR.n1017 0.120292
R13570 VPWR.n1020 VPWR.n1019 0.120292
R13571 VPWR.n1079 VPWR.n1078 0.120292
R13572 VPWR.n1072 VPWR.n1071 0.120292
R13573 VPWR.n1071 VPWR.n1048 0.120292
R13574 VPWR.n1064 VPWR.n1048 0.120292
R13575 VPWR.n1064 VPWR.n1063 0.120292
R13576 VPWR.n1063 VPWR.n1062 0.120292
R13577 VPWR.n1062 VPWR.n1050 0.120292
R13578 VPWR.n1056 VPWR.n1050 0.120292
R13579 VPWR.n1056 VPWR.n1055 0.120292
R13580 VPWR.n1118 VPWR.n1117 0.120292
R13581 VPWR.n1111 VPWR.n1110 0.120292
R13582 VPWR.n1110 VPWR.n1087 0.120292
R13583 VPWR.n1103 VPWR.n1087 0.120292
R13584 VPWR.n1103 VPWR.n1102 0.120292
R13585 VPWR.n1102 VPWR.n1101 0.120292
R13586 VPWR.n1101 VPWR.n1089 0.120292
R13587 VPWR.n1095 VPWR.n1089 0.120292
R13588 VPWR.n1095 VPWR.n1094 0.120292
R13589 VPWR.n1148 VPWR.n1147 0.120292
R13590 VPWR.n1147 VPWR.n1124 0.120292
R13591 VPWR.n1140 VPWR.n1124 0.120292
R13592 VPWR.n1140 VPWR.n1139 0.120292
R13593 VPWR.n1139 VPWR.n1138 0.120292
R13594 VPWR.n1138 VPWR.n1126 0.120292
R13595 VPWR.n1132 VPWR.n1126 0.120292
R13596 VPWR.n1132 VPWR.n1131 0.120292
R13597 VPWR.n3101 VPWR.n3087 0.120292
R13598 VPWR.n3085 VPWR.n3068 0.120292
R13599 VPWR.n3066 VPWR.n3048 0.120292
R13600 VPWR.n3046 VPWR.n3029 0.120292
R13601 VPWR.n3008 VPWR.n3007 0.120292
R13602 VPWR.n3009 VPWR.n3008 0.120292
R13603 VPWR.n3009 VPWR.n3000 0.120292
R13604 VPWR.n3014 VPWR.n3000 0.120292
R13605 VPWR.n3015 VPWR.n3014 0.120292
R13606 VPWR.n3015 VPWR.n2996 0.120292
R13607 VPWR.n3021 VPWR.n2996 0.120292
R13608 VPWR.n3023 VPWR.n2993 0.120292
R13609 VPWR.n3027 VPWR.n2993 0.120292
R13610 VPWR.n2972 VPWR.n2971 0.120292
R13611 VPWR.n2973 VPWR.n2972 0.120292
R13612 VPWR.n2973 VPWR.n2962 0.120292
R13613 VPWR.n2978 VPWR.n2962 0.120292
R13614 VPWR.n2979 VPWR.n2978 0.120292
R13615 VPWR.n2979 VPWR.n2958 0.120292
R13616 VPWR.n2984 VPWR.n2958 0.120292
R13617 VPWR.n2986 VPWR.n2955 0.120292
R13618 VPWR.n2991 VPWR.n2955 0.120292
R13619 VPWR.n2935 VPWR.n2934 0.120292
R13620 VPWR.n2936 VPWR.n2935 0.120292
R13621 VPWR.n2936 VPWR.n2925 0.120292
R13622 VPWR.n2941 VPWR.n2925 0.120292
R13623 VPWR.n2942 VPWR.n2941 0.120292
R13624 VPWR.n2942 VPWR.n2921 0.120292
R13625 VPWR.n2947 VPWR.n2921 0.120292
R13626 VPWR.n2949 VPWR.n2918 0.120292
R13627 VPWR.n2953 VPWR.n2918 0.120292
R13628 VPWR.n2897 VPWR.n2893 0.120292
R13629 VPWR.n2905 VPWR.n2893 0.120292
R13630 VPWR.n2906 VPWR.n2905 0.120292
R13631 VPWR.n2907 VPWR.n2906 0.120292
R13632 VPWR.n2907 VPWR.n2889 0.120292
R13633 VPWR.n2912 VPWR.n2889 0.120292
R13634 VPWR.n2913 VPWR.n2912 0.120292
R13635 VPWR VPWR.n1580 0.118556
R13636 VPWR.n1576 VPWR 0.118556
R13637 VPWR VPWR.n1561 0.118556
R13638 VPWR VPWR.n1549 0.118556
R13639 VPWR.n1544 VPWR 0.118556
R13640 VPWR VPWR.n1351 0.118556
R13641 VPWR VPWR.n1362 0.118556
R13642 VPWR VPWR.n1373 0.118556
R13643 VPWR VPWR.n1384 0.118556
R13644 VPWR VPWR.n1395 0.118556
R13645 VPWR VPWR.n1406 0.118556
R13646 VPWR.n1339 VPWR 0.118556
R13647 VPWR VPWR.n1324 0.118556
R13648 VPWR VPWR.n1312 0.118556
R13649 VPWR.n1307 VPWR 0.118556
R13650 VPWR VPWR.n1292 0.118556
R13651 VPWR.n90 VPWR 0.118556
R13652 VPWR.n279 VPWR 0.118556
R13653 VPWR.n260 VPWR 0.118556
R13654 VPWR.n105 VPWR 0.118556
R13655 VPWR.n245 VPWR 0.118556
R13656 VPWR.n226 VPWR 0.118556
R13657 VPWR.n110 VPWR 0.118556
R13658 VPWR.n211 VPWR 0.118556
R13659 VPWR.n192 VPWR 0.118556
R13660 VPWR.n115 VPWR 0.118556
R13661 VPWR.n177 VPWR 0.118556
R13662 VPWR.n158 VPWR 0.118556
R13663 VPWR.n120 VPWR 0.118556
R13664 VPWR.n143 VPWR 0.118556
R13665 VPWR.n99 VPWR 0.118556
R13666 VPWR VPWR.n124 0.118556
R13667 VPWR.n1431 VPWR.n1430 0.108238
R13668 VPWR.n1429 VPWR.n1428 0.108238
R13669 VPWR.n1686 VPWR.n1685 0.108238
R13670 VPWR.n1432 VPWR.n1422 0.108238
R13671 VPWR.n1417 VPWR.n1170 0.108238
R13672 VPWR.n1481 VPWR.n1416 0.108238
R13673 VPWR.n1480 VPWR.n1479 0.108238
R13674 VPWR.n1478 VPWR.n1477 0.108238
R13675 VPWR.n1476 VPWR.n1475 0.108238
R13676 VPWR.n1474 VPWR.n1473 0.108238
R13677 VPWR.n1639 VPWR.n1229 0.108238
R13678 VPWR.n1638 VPWR.n1637 0.108238
R13679 VPWR.n1613 VPWR.n1612 0.108238
R13680 VPWR.n1699 VPWR.n931 0.108238
R13681 VPWR.n1698 VPWR.n1697 0.108238
R13682 VPWR.n1696 VPWR.n918 0.108238
R13683 VPWR VPWR.n1429 0.100405
R13684 VPWR.n2754 VPWR 0.100405
R13685 VPWR.n2753 VPWR 0.100405
R13686 VPWR.n2752 VPWR 0.100405
R13687 VPWR.n2737 VPWR 0.100405
R13688 VPWR.n2568 VPWR 0.100405
R13689 VPWR.n2726 VPWR 0.100405
R13690 VPWR.n2725 VPWR 0.100405
R13691 VPWR.n447 VPWR 0.100405
R13692 VPWR VPWR.n449 0.100405
R13693 VPWR VPWR.n2571 0.100405
R13694 VPWR VPWR.n2572 0.100405
R13695 VPWR VPWR.n2573 0.100405
R13696 VPWR.n2576 VPWR 0.100405
R13697 VPWR.n2575 VPWR 0.100405
R13698 VPWR.n2574 VPWR 0.100405
R13699 VPWR.n2415 VPWR 0.100405
R13700 VPWR.n2547 VPWR 0.100405
R13701 VPWR.n2546 VPWR 0.100405
R13702 VPWR VPWR.n2451 0.100405
R13703 VPWR VPWR.n2452 0.100405
R13704 VPWR.n2453 VPWR 0.100405
R13705 VPWR.n2528 VPWR 0.100405
R13706 VPWR.n2527 VPWR 0.100405
R13707 VPWR VPWR.n2666 0.100405
R13708 VPWR.n2653 VPWR 0.100405
R13709 VPWR VPWR.n2652 0.100405
R13710 VPWR.n2641 VPWR 0.100405
R13711 VPWR VPWR.n2640 0.100405
R13712 VPWR.n2505 VPWR 0.100405
R13713 VPWR.n2526 VPWR 0.100405
R13714 VPWR.n2420 VPWR 0.100405
R13715 VPWR.n2419 VPWR 0.100405
R13716 VPWR.n2418 VPWR 0.100405
R13717 VPWR.n2448 VPWR 0.100405
R13718 VPWR.n2447 VPWR 0.100405
R13719 VPWR VPWR.n2456 0.100405
R13720 VPWR VPWR.n2457 0.100405
R13721 VPWR.n2459 VPWR 0.100405
R13722 VPWR.n2498 VPWR 0.100405
R13723 VPWR.n2499 VPWR 0.100405
R13724 VPWR.n2500 VPWR 0.100405
R13725 VPWR.n2501 VPWR 0.100405
R13726 VPWR.n2502 VPWR 0.100405
R13727 VPWR.n2503 VPWR 0.100405
R13728 VPWR.n2458 VPWR 0.100405
R13729 VPWR.n2413 VPWR 0.100405
R13730 VPWR.n2412 VPWR 0.100405
R13731 VPWR VPWR.n2297 0.100405
R13732 VPWR VPWR.n2298 0.100405
R13733 VPWR VPWR.n2299 0.100405
R13734 VPWR VPWR.n2300 0.100405
R13735 VPWR.n2302 VPWR 0.100405
R13736 VPWR.n2301 VPWR 0.100405
R13737 VPWR.n2361 VPWR 0.100405
R13738 VPWR.n546 VPWR 0.100405
R13739 VPWR.n2372 VPWR 0.100405
R13740 VPWR.n2373 VPWR 0.100405
R13741 VPWR.n2339 VPWR 0.100405
R13742 VPWR VPWR.n2338 0.100405
R13743 VPWR VPWR.n2337 0.100405
R13744 VPWR.n701 VPWR 0.100405
R13745 VPWR.n700 VPWR 0.100405
R13746 VPWR.n2294 VPWR 0.100405
R13747 VPWR.n2293 VPWR 0.100405
R13748 VPWR VPWR.n2281 0.100405
R13749 VPWR.n2282 VPWR 0.100405
R13750 VPWR VPWR.n2305 0.100405
R13751 VPWR.n2306 VPWR 0.100405
R13752 VPWR.n2345 VPWR 0.100405
R13753 VPWR.n2346 VPWR 0.100405
R13754 VPWR VPWR.n2344 0.100405
R13755 VPWR VPWR.n2343 0.100405
R13756 VPWR VPWR.n2342 0.100405
R13757 VPWR.n2333 VPWR 0.100405
R13758 VPWR.n2334 VPWR 0.100405
R13759 VPWR.n2130 VPWR 0.100405
R13760 VPWR.n2129 VPWR 0.100405
R13761 VPWR.n2128 VPWR 0.100405
R13762 VPWR.n2127 VPWR 0.100405
R13763 VPWR.n2278 VPWR 0.100405
R13764 VPWR.n2277 VPWR 0.100405
R13765 VPWR.n2276 VPWR 0.100405
R13766 VPWR.n2275 VPWR 0.100405
R13767 VPWR.n2251 VPWR 0.100405
R13768 VPWR VPWR.n2249 0.100405
R13769 VPWR VPWR.n2248 0.100405
R13770 VPWR.n2271 VPWR 0.100405
R13771 VPWR.n2272 VPWR 0.100405
R13772 VPWR.n2273 VPWR 0.100405
R13773 VPWR.n2274 VPWR 0.100405
R13774 VPWR VPWR.n2133 0.100405
R13775 VPWR.n2134 VPWR 0.100405
R13776 VPWR VPWR.n2148 0.100405
R13777 VPWR.n2150 VPWR 0.100405
R13778 VPWR.n2149 VPWR 0.100405
R13779 VPWR VPWR.n2162 0.100405
R13780 VPWR.n2163 VPWR 0.100405
R13781 VPWR VPWR.n2174 0.100405
R13782 VPWR VPWR.n591 0.100405
R13783 VPWR.n2244 VPWR 0.100405
R13784 VPWR.n2245 VPWR 0.100405
R13785 VPWR.n2202 VPWR 0.100405
R13786 VPWR.n2203 VPWR 0.100405
R13787 VPWR VPWR.n2201 0.100405
R13788 VPWR.n2175 VPWR 0.100405
R13789 VPWR.n2123 VPWR 0.100405
R13790 VPWR.n2122 VPWR 0.100405
R13791 VPWR.n2121 VPWR 0.100405
R13792 VPWR.n2120 VPWR 0.100405
R13793 VPWR.n2119 VPWR 0.100405
R13794 VPWR.n708 VPWR 0.100405
R13795 VPWR.n707 VPWR 0.100405
R13796 VPWR.n706 VPWR 0.100405
R13797 VPWR VPWR.n2230 0.100405
R13798 VPWR.n2207 VPWR 0.100405
R13799 VPWR.n2208 VPWR 0.100405
R13800 VPWR.n2209 VPWR 0.100405
R13801 VPWR VPWR.n2206 0.100405
R13802 VPWR.n704 VPWR 0.100405
R13803 VPWR.n705 VPWR 0.100405
R13804 VPWR VPWR.n1927 0.100405
R13805 VPWR.n1928 VPWR 0.100405
R13806 VPWR VPWR.n1949 0.100405
R13807 VPWR.n1950 VPWR 0.100405
R13808 VPWR.n2063 VPWR 0.100405
R13809 VPWR.n2062 VPWR 0.100405
R13810 VPWR.n755 VPWR 0.100405
R13811 VPWR.n2051 VPWR 0.100405
R13812 VPWR VPWR.n2020 0.100405
R13813 VPWR.n2031 VPWR 0.100405
R13814 VPWR.n2032 VPWR 0.100405
R13815 VPWR.n1976 VPWR 0.100405
R13816 VPWR.n1977 VPWR 0.100405
R13817 VPWR.n1978 VPWR 0.100405
R13818 VPWR.n2050 VPWR 0.100405
R13819 VPWR.n1920 VPWR 0.100405
R13820 VPWR.n1919 VPWR 0.100405
R13821 VPWR.n1918 VPWR 0.100405
R13822 VPWR VPWR.n1953 0.100405
R13823 VPWR VPWR.n1954 0.100405
R13824 VPWR VPWR.n1955 0.100405
R13825 VPWR.n1958 VPWR 0.100405
R13826 VPWR.n1957 VPWR 0.100405
R13827 VPWR.n2011 VPWR 0.100405
R13828 VPWR VPWR.n2010 0.100405
R13829 VPWR VPWR.n2009 0.100405
R13830 VPWR VPWR.n2008 0.100405
R13831 VPWR.n1982 VPWR 0.100405
R13832 VPWR VPWR.n1981 0.100405
R13833 VPWR.n1956 VPWR 0.100405
R13834 VPWR.n1915 VPWR 0.100405
R13835 VPWR.n1914 VPWR 0.100405
R13836 VPWR VPWR.n1808 0.100405
R13837 VPWR VPWR.n1809 0.100405
R13838 VPWR.n1810 VPWR 0.100405
R13839 VPWR.n1896 VPWR 0.100405
R13840 VPWR.n1895 VPWR 0.100405
R13841 VPWR.n1894 VPWR 0.100405
R13842 VPWR VPWR.n2014 0.100405
R13843 VPWR.n1869 VPWR 0.100405
R13844 VPWR VPWR.n1868 0.100405
R13845 VPWR.n853 VPWR 0.100405
R13846 VPWR.n854 VPWR 0.100405
R13847 VPWR.n855 VPWR 0.100405
R13848 VPWR.n856 VPWR 0.100405
R13849 VPWR.n2633 VPWR 0.100405
R13850 VPWR.n2634 VPWR 0.100405
R13851 VPWR.n2635 VPWR 0.100405
R13852 VPWR.n2636 VPWR 0.100405
R13853 VPWR.n2637 VPWR 0.100405
R13854 VPWR VPWR.n2632 0.100405
R13855 VPWR VPWR.n2631 0.100405
R13856 VPWR VPWR.n2630 0.100405
R13857 VPWR.n1776 VPWR 0.100405
R13858 VPWR.n1775 VPWR 0.100405
R13859 VPWR.n1805 VPWR 0.100405
R13860 VPWR.n1804 VPWR 0.100405
R13861 VPWR VPWR.n1813 0.100405
R13862 VPWR VPWR.n1814 0.100405
R13863 VPWR.n1816 VPWR 0.100405
R13864 VPWR.n1815 VPWR 0.100405
R13865 VPWR VPWR.n1828 0.100405
R13866 VPWR.n1863 VPWR 0.100405
R13867 VPWR.n1864 VPWR 0.100405
R13868 VPWR.n1865 VPWR 0.100405
R13869 VPWR.n1844 VPWR 0.100405
R13870 VPWR VPWR.n1843 0.100405
R13871 VPWR.n1829 VPWR 0.100405
R13872 VPWR.n2678 VPWR 0.100405
R13873 VPWR.n425 VPWR 0.100405
R13874 VPWR.n2689 VPWR 0.100405
R13875 VPWR.n2690 VPWR 0.100405
R13876 VPWR.n435 VPWR 0.100405
R13877 VPWR.n2701 VPWR 0.100405
R13878 VPWR.n2702 VPWR 0.100405
R13879 VPWR.n438 VPWR 0.100405
R13880 VPWR.n2713 VPWR 0.100405
R13881 VPWR.n2714 VPWR 0.100405
R13882 VPWR.n1773 VPWR 0.100405
R13883 VPWR.n1772 VPWR 0.100405
R13884 VPWR VPWR.n889 0.100405
R13885 VPWR VPWR.n890 0.100405
R13886 VPWR VPWR.n891 0.100405
R13887 VPWR.n1754 VPWR 0.100405
R13888 VPWR.n1753 VPWR 0.100405
R13889 VPWR.n1752 VPWR 0.100405
R13890 VPWR VPWR.n912 0.100405
R13891 VPWR VPWR.n913 0.100405
R13892 VPWR VPWR.n914 0.100405
R13893 VPWR.n1726 VPWR 0.100405
R13894 VPWR.n1727 VPWR 0.100405
R13895 VPWR VPWR.n916 0.100405
R13896 VPWR VPWR.n915 0.100405
R13897 VPWR.n2740 VPWR 0.100405
R13898 VPWR.n2741 VPWR 0.100405
R13899 VPWR.n2742 VPWR 0.100405
R13900 VPWR.n2743 VPWR 0.100405
R13901 VPWR.n2744 VPWR 0.100405
R13902 VPWR.n2745 VPWR 0.100405
R13903 VPWR.n2746 VPWR 0.100405
R13904 VPWR.n2747 VPWR 0.100405
R13905 VPWR.n2748 VPWR 0.100405
R13906 VPWR.n2749 VPWR 0.100405
R13907 VPWR.n2750 VPWR 0.100405
R13908 VPWR.n2751 VPWR 0.100405
R13909 VPWR.n1422 VPWR 0.100405
R13910 VPWR VPWR.n1170 0.100405
R13911 VPWR.n1481 VPWR 0.100405
R13912 VPWR.n1479 VPWR 0.100405
R13913 VPWR.n1477 VPWR 0.100405
R13914 VPWR.n1475 VPWR 0.100405
R13915 VPWR.n1473 VPWR 0.100405
R13916 VPWR.n1639 VPWR 0.100405
R13917 VPWR.n1637 VPWR 0.100405
R13918 VPWR.n1613 VPWR 0.100405
R13919 VPWR.n1699 VPWR 0.100405
R13920 VPWR.n1697 VPWR 0.100405
R13921 VPWR VPWR.n918 0.100405
R13922 VPWR VPWR.n1431 0.100405
R13923 VPWR.n2757 VPWR 0.100405
R13924 VPWR VPWR.n2768 0.100405
R13925 VPWR.n2769 VPWR 0.100405
R13926 VPWR VPWR.n2780 0.100405
R13927 VPWR.n2781 VPWR 0.100405
R13928 VPWR VPWR.n2792 0.100405
R13929 VPWR.n2793 VPWR 0.100405
R13930 VPWR VPWR.n2804 0.100405
R13931 VPWR.n2805 VPWR 0.100405
R13932 VPWR VPWR.n2816 0.100405
R13933 VPWR.n2817 VPWR 0.100405
R13934 VPWR VPWR.n2828 0.100405
R13935 VPWR.n2829 VPWR 0.100405
R13936 VPWR VPWR.n2840 0.100405
R13937 VPWR.n2841 VPWR 0.100405
R13938 VPWR.n1234 VPWR 0.100405
R13939 VPWR.n1594 VPWR 0.100405
R13940 VPWR.n1595 VPWR 0.100405
R13941 VPWR.n1596 VPWR 0.100405
R13942 VPWR.n1507 VPWR 0.100405
R13943 VPWR.n1508 VPWR 0.100405
R13944 VPWR.n1509 VPWR 0.100405
R13945 VPWR VPWR.n1506 0.100405
R13946 VPWR.n1495 VPWR 0.100405
R13947 VPWR VPWR.n1494 0.100405
R13948 VPWR.n1483 VPWR 0.100405
R13949 VPWR.n1665 VPWR 0.100405
R13950 VPWR.n1666 VPWR 0.100405
R13951 VPWR VPWR.n1168 0.100405
R13952 VPWR.n1678 VPWR 0.100405
R13953 VPWR VPWR.n3087 0.0994583
R13954 VPWR VPWR.n3068 0.0994583
R13955 VPWR VPWR.n1034 0.0981562
R13956 VPWR.n1079 VPWR 0.0981562
R13957 VPWR.n1118 VPWR 0.0981562
R13958 VPWR.n9 VPWR 0.0968542
R13959 VPWR.n952 VPWR 0.0968542
R13960 VPWR.n975 VPWR 0.0968542
R13961 VPWR.n999 VPWR 0.0968542
R13962 VPWR.n1041 VPWR 0.0968542
R13963 VPWR VPWR.n3048 0.0968542
R13964 VPWR VPWR.n3029 0.0968542
R13965 VPWR.n3007 VPWR 0.0968542
R13966 VPWR.n2971 VPWR 0.0968542
R13967 VPWR.n2934 VPWR 0.0968542
R13968 VPWR.n2897 VPWR 0.0968542
R13969 VPWR.n1430 VPWR 0.0945
R13970 VPWR.n1428 VPWR 0.0945
R13971 VPWR VPWR.n1417 0.0945
R13972 VPWR.n1416 VPWR 0.0945
R13973 VPWR VPWR.n1480 0.0945
R13974 VPWR VPWR.n1478 0.0945
R13975 VPWR VPWR.n1476 0.0945
R13976 VPWR VPWR.n1474 0.0945
R13977 VPWR VPWR.n1229 0.0945
R13978 VPWR VPWR.n1638 0.0945
R13979 VPWR.n1612 VPWR 0.0945
R13980 VPWR VPWR.n931 0.0945
R13981 VPWR VPWR.n1698 0.0945
R13982 VPWR VPWR.n1696 0.0945
R13983 VPWR.n1686 VPWR 0.0945
R13984 VPWR.n1432 VPWR 0.0945
R13985 VPWR.n37 VPWR.n20 0.0939125
R13986 VPWR.n1291 VPWR 0.093504
R13987 VPWR.n1302 VPWR 0.093504
R13988 VPWR.n1286 VPWR 0.093504
R13989 VPWR.n1322 VPWR 0.093504
R13990 VPWR.n1334 VPWR 0.093504
R13991 VPWR VPWR.n1410 0.093504
R13992 VPWR VPWR.n1399 0.093504
R13993 VPWR VPWR.n1388 0.093504
R13994 VPWR VPWR.n1377 0.093504
R13995 VPWR VPWR.n1366 0.093504
R13996 VPWR VPWR.n1355 0.093504
R13997 VPWR VPWR.n1252 0.093504
R13998 VPWR VPWR.n1249 0.093504
R13999 VPWR.n1559 VPWR 0.093504
R14000 VPWR.n1571 VPWR 0.093504
R14001 VPWR.n1244 VPWR 0.093504
R14002 VPWR.n96 VPWR 0.093504
R14003 VPWR VPWR.n128 0.093504
R14004 VPWR.n140 VPWR 0.093504
R14005 VPWR VPWR.n150 0.093504
R14006 VPWR VPWR.n162 0.093504
R14007 VPWR.n174 VPWR 0.093504
R14008 VPWR VPWR.n184 0.093504
R14009 VPWR VPWR.n196 0.093504
R14010 VPWR.n208 VPWR 0.093504
R14011 VPWR VPWR.n218 0.093504
R14012 VPWR VPWR.n230 0.093504
R14013 VPWR.n242 VPWR 0.093504
R14014 VPWR VPWR.n252 0.093504
R14015 VPWR VPWR.n264 0.093504
R14016 VPWR.n276 VPWR 0.093504
R14017 VPWR VPWR.n286 0.093504
R14018 VPWR.n2887 VPWR 0.0849042
R14019 VPWR.n1292 VPWR.n1287 0.0845517
R14020 VPWR.n1308 VPWR.n1307 0.0845517
R14021 VPWR.n1312 VPWR.n1311 0.0845517
R14022 VPWR.n1324 VPWR.n1323 0.0845517
R14023 VPWR.n1340 VPWR.n1339 0.0845517
R14024 VPWR.n1406 VPWR.n1272 0.0845517
R14025 VPWR.n1395 VPWR.n1273 0.0845517
R14026 VPWR.n1384 VPWR.n1274 0.0845517
R14027 VPWR.n1373 VPWR.n1275 0.0845517
R14028 VPWR.n1362 VPWR.n1347 0.0845517
R14029 VPWR.n1351 VPWR.n1348 0.0845517
R14030 VPWR.n1545 VPWR.n1544 0.0845517
R14031 VPWR.n1549 VPWR.n1548 0.0845517
R14032 VPWR.n1561 VPWR.n1560 0.0845517
R14033 VPWR.n1577 VPWR.n1576 0.0845517
R14034 VPWR.n1580 VPWR.n1579 0.0845517
R14035 VPWR.n100 VPWR.n99 0.0845517
R14036 VPWR.n124 VPWR.n121 0.0845517
R14037 VPWR.n144 VPWR.n143 0.0845517
R14038 VPWR.n147 VPWR.n120 0.0845517
R14039 VPWR.n159 VPWR.n158 0.0845517
R14040 VPWR.n178 VPWR.n177 0.0845517
R14041 VPWR.n181 VPWR.n115 0.0845517
R14042 VPWR.n193 VPWR.n192 0.0845517
R14043 VPWR.n212 VPWR.n211 0.0845517
R14044 VPWR.n215 VPWR.n110 0.0845517
R14045 VPWR.n227 VPWR.n226 0.0845517
R14046 VPWR.n246 VPWR.n245 0.0845517
R14047 VPWR.n249 VPWR.n105 0.0845517
R14048 VPWR.n261 VPWR.n260 0.0845517
R14049 VPWR.n280 VPWR.n279 0.0845517
R14050 VPWR.n283 VPWR.n90 0.0845517
R14051 VPWR.n1428 VPWR.n1427 0.0740128
R14052 VPWR.n1430 VPWR.n1423 0.071
R14053 VPWR.n1438 VPWR.n1417 0.071
R14054 VPWR.n1443 VPWR.n1416 0.071
R14055 VPWR.n1480 VPWR.n1448 0.071
R14056 VPWR.n1478 VPWR.n1453 0.071
R14057 VPWR.n1476 VPWR.n1458 0.071
R14058 VPWR.n1474 VPWR.n1472 0.071
R14059 VPWR.n1467 VPWR.n1229 0.071
R14060 VPWR.n1638 VPWR.n1230 0.071
R14061 VPWR.n1612 VPWR.n1611 0.071
R14062 VPWR.n1606 VPWR.n931 0.071
R14063 VPWR.n1698 VPWR.n932 0.071
R14064 VPWR.n1696 VPWR.n1695 0.071
R14065 VPWR.n1690 VPWR.n1686 0.071
R14066 VPWR.n1433 VPWR.n1432 0.071
R14067 VPWR VPWR.n1289 0.0678077
R14068 VPWR VPWR.n1300 0.0678077
R14069 VPWR VPWR.n1284 0.0678077
R14070 VPWR VPWR.n1320 0.0678077
R14071 VPWR VPWR.n1332 0.0678077
R14072 VPWR.n1411 VPWR 0.0678077
R14073 VPWR.n1400 VPWR 0.0678077
R14074 VPWR.n1389 VPWR 0.0678077
R14075 VPWR.n1378 VPWR 0.0678077
R14076 VPWR.n1367 VPWR 0.0678077
R14077 VPWR.n1356 VPWR 0.0678077
R14078 VPWR.n1255 VPWR 0.0678077
R14079 VPWR.n1536 VPWR 0.0678077
R14080 VPWR VPWR.n1557 0.0678077
R14081 VPWR VPWR.n1569 0.0678077
R14082 VPWR VPWR.n1242 0.0678077
R14083 VPWR VPWR.n94 0.0678077
R14084 VPWR.n129 VPWR 0.0678077
R14085 VPWR VPWR.n138 0.0678077
R14086 VPWR.n151 VPWR 0.0678077
R14087 VPWR.n163 VPWR 0.0678077
R14088 VPWR VPWR.n172 0.0678077
R14089 VPWR.n185 VPWR 0.0678077
R14090 VPWR.n197 VPWR 0.0678077
R14091 VPWR VPWR.n206 0.0678077
R14092 VPWR.n219 VPWR 0.0678077
R14093 VPWR.n231 VPWR 0.0678077
R14094 VPWR VPWR.n240 0.0678077
R14095 VPWR.n253 VPWR 0.0678077
R14096 VPWR.n265 VPWR 0.0678077
R14097 VPWR VPWR.n274 0.0678077
R14098 VPWR.n287 VPWR 0.0678077
R14099 VPWR.n3115 VPWR 0.063
R14100 VPWR VPWR.n1296 0.063
R14101 VPWR.n1304 VPWR 0.063
R14102 VPWR VPWR.n1316 0.063
R14103 VPWR VPWR.n1328 0.063
R14104 VPWR.n1336 VPWR 0.063
R14105 VPWR.n1405 VPWR 0.063
R14106 VPWR.n1394 VPWR 0.063
R14107 VPWR.n1383 VPWR 0.063
R14108 VPWR.n1372 VPWR 0.063
R14109 VPWR.n1361 VPWR 0.063
R14110 VPWR.n1350 VPWR 0.063
R14111 VPWR.n1541 VPWR 0.063
R14112 VPWR VPWR.n1553 0.063
R14113 VPWR VPWR.n1565 0.063
R14114 VPWR.n1573 VPWR 0.063
R14115 VPWR VPWR.n1584 0.063
R14116 VPWR.n123 VPWR 0.063
R14117 VPWR.n134 VPWR 0.063
R14118 VPWR VPWR.n118 0.063
R14119 VPWR.n156 VPWR 0.063
R14120 VPWR.n168 VPWR 0.063
R14121 VPWR VPWR.n113 0.063
R14122 VPWR.n190 VPWR 0.063
R14123 VPWR.n202 VPWR 0.063
R14124 VPWR VPWR.n108 0.063
R14125 VPWR.n224 VPWR 0.063
R14126 VPWR.n236 VPWR 0.063
R14127 VPWR VPWR.n103 0.063
R14128 VPWR.n258 VPWR 0.063
R14129 VPWR.n270 VPWR 0.063
R14130 VPWR VPWR.n88 0.063
R14131 VPWR.n92 VPWR 0.063
R14132 VPWR.n1289 VPWR 0.0608448
R14133 VPWR.n1300 VPWR 0.0608448
R14134 VPWR.n1284 VPWR 0.0608448
R14135 VPWR.n1320 VPWR 0.0608448
R14136 VPWR.n1332 VPWR 0.0608448
R14137 VPWR.n1411 VPWR 0.0608448
R14138 VPWR.n1400 VPWR 0.0608448
R14139 VPWR.n1389 VPWR 0.0608448
R14140 VPWR.n1378 VPWR 0.0608448
R14141 VPWR.n1367 VPWR 0.0608448
R14142 VPWR.n1356 VPWR 0.0608448
R14143 VPWR.n1255 VPWR 0.0608448
R14144 VPWR.n1536 VPWR 0.0608448
R14145 VPWR.n1557 VPWR 0.0608448
R14146 VPWR.n1569 VPWR 0.0608448
R14147 VPWR.n1242 VPWR 0.0608448
R14148 VPWR.n94 VPWR 0.0608448
R14149 VPWR.n129 VPWR 0.0608448
R14150 VPWR.n138 VPWR 0.0608448
R14151 VPWR.n151 VPWR 0.0608448
R14152 VPWR.n163 VPWR 0.0608448
R14153 VPWR.n172 VPWR 0.0608448
R14154 VPWR.n185 VPWR 0.0608448
R14155 VPWR.n197 VPWR 0.0608448
R14156 VPWR.n206 VPWR 0.0608448
R14157 VPWR.n219 VPWR 0.0608448
R14158 VPWR.n231 VPWR 0.0608448
R14159 VPWR.n240 VPWR 0.0608448
R14160 VPWR.n253 VPWR 0.0608448
R14161 VPWR.n265 VPWR 0.0608448
R14162 VPWR.n274 VPWR 0.0608448
R14163 VPWR.n287 VPWR 0.0608448
R14164 VPWR VPWR.n13 0.0603958
R14165 VPWR VPWR.n12 0.0603958
R14166 VPWR VPWR.n957 0.0603958
R14167 VPWR VPWR.n956 0.0603958
R14168 VPWR VPWR.n980 0.0603958
R14169 VPWR VPWR.n979 0.0603958
R14170 VPWR VPWR.n1004 0.0603958
R14171 VPWR VPWR.n1003 0.0603958
R14172 VPWR.n1040 VPWR 0.0603958
R14173 VPWR VPWR.n1039 0.0603958
R14174 VPWR.n1035 VPWR 0.0603958
R14175 VPWR.n1026 VPWR 0.0603958
R14176 VPWR VPWR.n1025 0.0603958
R14177 VPWR.n1078 VPWR 0.0603958
R14178 VPWR VPWR.n1077 0.0603958
R14179 VPWR.n1072 VPWR 0.0603958
R14180 VPWR.n1117 VPWR 0.0603958
R14181 VPWR VPWR.n1116 0.0603958
R14182 VPWR.n1111 VPWR 0.0603958
R14183 VPWR.n1148 VPWR 0.0603958
R14184 VPWR VPWR.n3089 0.0603958
R14185 VPWR VPWR.n3088 0.0603958
R14186 VPWR VPWR.n3101 0.0603958
R14187 VPWR.n3080 VPWR 0.0603958
R14188 VPWR.n3081 VPWR 0.0603958
R14189 VPWR VPWR.n3085 0.0603958
R14190 VPWR.n3060 VPWR 0.0603958
R14191 VPWR.n3061 VPWR 0.0603958
R14192 VPWR VPWR.n3066 0.0603958
R14193 VPWR.n3041 VPWR 0.0603958
R14194 VPWR.n3042 VPWR 0.0603958
R14195 VPWR VPWR.n3046 0.0603958
R14196 VPWR.n3022 VPWR 0.0603958
R14197 VPWR.n3023 VPWR 0.0603958
R14198 VPWR VPWR.n2984 0.0603958
R14199 VPWR.n2985 VPWR 0.0603958
R14200 VPWR.n2986 VPWR 0.0603958
R14201 VPWR VPWR.n2947 0.0603958
R14202 VPWR.n2948 VPWR 0.0603958
R14203 VPWR.n2949 VPWR 0.0603958
R14204 VPWR.n2913 VPWR 0.0603958
R14205 VPWR.n2916 VPWR 0.0603958
R14206 VPWR.n1436 VPWR.n1435 0.0599512
R14207 VPWR.n1420 VPWR.n1419 0.0599512
R14208 VPWR.n1426 VPWR.n1425 0.0599512
R14209 VPWR.n1441 VPWR.n1440 0.0599512
R14210 VPWR.n1446 VPWR.n1445 0.0599512
R14211 VPWR.n1451 VPWR.n1450 0.0599512
R14212 VPWR.n1456 VPWR.n1455 0.0599512
R14213 VPWR.n1461 VPWR.n1460 0.0599512
R14214 VPWR.n1470 VPWR.n1469 0.0599512
R14215 VPWR.n1465 VPWR.n1464 0.0599512
R14216 VPWR.n1600 VPWR.n1599 0.0599512
R14217 VPWR.n1609 VPWR.n1608 0.0599512
R14218 VPWR.n1604 VPWR.n1603 0.0599512
R14219 VPWR.n935 VPWR.n934 0.0599512
R14220 VPWR.n1693 VPWR.n1692 0.0599512
R14221 VPWR.n1689 VPWR.n1688 0.0599512
R14222 VPWR.n1294 VPWR.n1291 0.0565345
R14223 VPWR.n1292 VPWR 0.0565345
R14224 VPWR.n1305 VPWR.n1302 0.0565345
R14225 VPWR.n1307 VPWR 0.0565345
R14226 VPWR.n1314 VPWR.n1286 0.0565345
R14227 VPWR.n1312 VPWR 0.0565345
R14228 VPWR.n1326 VPWR.n1322 0.0565345
R14229 VPWR.n1324 VPWR 0.0565345
R14230 VPWR.n1337 VPWR.n1334 0.0565345
R14231 VPWR.n1339 VPWR 0.0565345
R14232 VPWR.n1410 VPWR.n1408 0.0565345
R14233 VPWR.n1406 VPWR 0.0565345
R14234 VPWR.n1399 VPWR.n1397 0.0565345
R14235 VPWR.n1395 VPWR 0.0565345
R14236 VPWR.n1388 VPWR.n1386 0.0565345
R14237 VPWR.n1384 VPWR 0.0565345
R14238 VPWR.n1377 VPWR.n1375 0.0565345
R14239 VPWR.n1373 VPWR 0.0565345
R14240 VPWR.n1366 VPWR.n1364 0.0565345
R14241 VPWR.n1362 VPWR 0.0565345
R14242 VPWR.n1355 VPWR.n1353 0.0565345
R14243 VPWR.n1351 VPWR 0.0565345
R14244 VPWR.n1542 VPWR.n1252 0.0565345
R14245 VPWR.n1544 VPWR 0.0565345
R14246 VPWR.n1551 VPWR.n1249 0.0565345
R14247 VPWR.n1549 VPWR 0.0565345
R14248 VPWR.n1563 VPWR.n1559 0.0565345
R14249 VPWR.n1561 VPWR 0.0565345
R14250 VPWR.n1574 VPWR.n1571 0.0565345
R14251 VPWR.n1576 VPWR 0.0565345
R14252 VPWR.n1582 VPWR.n1244 0.0565345
R14253 VPWR.n1580 VPWR 0.0565345
R14254 VPWR.n97 VPWR.n96 0.0565345
R14255 VPWR.n99 VPWR 0.0565345
R14256 VPWR.n128 VPWR.n126 0.0565345
R14257 VPWR.n124 VPWR 0.0565345
R14258 VPWR.n141 VPWR.n140 0.0565345
R14259 VPWR.n143 VPWR 0.0565345
R14260 VPWR.n150 VPWR.n148 0.0565345
R14261 VPWR.n120 VPWR 0.0565345
R14262 VPWR.n162 VPWR.n160 0.0565345
R14263 VPWR.n158 VPWR 0.0565345
R14264 VPWR.n175 VPWR.n174 0.0565345
R14265 VPWR.n177 VPWR 0.0565345
R14266 VPWR.n184 VPWR.n182 0.0565345
R14267 VPWR.n115 VPWR 0.0565345
R14268 VPWR.n196 VPWR.n194 0.0565345
R14269 VPWR.n192 VPWR 0.0565345
R14270 VPWR.n209 VPWR.n208 0.0565345
R14271 VPWR.n211 VPWR 0.0565345
R14272 VPWR.n218 VPWR.n216 0.0565345
R14273 VPWR.n110 VPWR 0.0565345
R14274 VPWR.n230 VPWR.n228 0.0565345
R14275 VPWR.n226 VPWR 0.0565345
R14276 VPWR.n243 VPWR.n242 0.0565345
R14277 VPWR.n245 VPWR 0.0565345
R14278 VPWR.n252 VPWR.n250 0.0565345
R14279 VPWR.n105 VPWR 0.0565345
R14280 VPWR.n264 VPWR.n262 0.0565345
R14281 VPWR.n260 VPWR 0.0565345
R14282 VPWR.n277 VPWR.n276 0.0565345
R14283 VPWR.n279 VPWR 0.0565345
R14284 VPWR.n286 VPWR.n284 0.0565345
R14285 VPWR.n90 VPWR 0.0565345
R14286 VPWR.n1435 VPWR 0.0469286
R14287 VPWR.n1419 VPWR 0.0469286
R14288 VPWR.n1425 VPWR 0.0469286
R14289 VPWR.n1440 VPWR 0.0469286
R14290 VPWR.n1445 VPWR 0.0469286
R14291 VPWR.n1450 VPWR 0.0469286
R14292 VPWR.n1455 VPWR 0.0469286
R14293 VPWR.n1460 VPWR 0.0469286
R14294 VPWR.n1469 VPWR 0.0469286
R14295 VPWR.n1464 VPWR 0.0469286
R14296 VPWR.n1599 VPWR 0.0469286
R14297 VPWR.n1608 VPWR 0.0469286
R14298 VPWR.n1603 VPWR 0.0469286
R14299 VPWR.n934 VPWR 0.0469286
R14300 VPWR.n1692 VPWR 0.0469286
R14301 VPWR.n1688 VPWR 0.0469286
R14302 VPWR.n1435 VPWR 0.0401341
R14303 VPWR.n1419 VPWR 0.0401341
R14304 VPWR.n1425 VPWR 0.0401341
R14305 VPWR.n1440 VPWR 0.0401341
R14306 VPWR.n1445 VPWR 0.0401341
R14307 VPWR.n1450 VPWR 0.0401341
R14308 VPWR.n1455 VPWR 0.0401341
R14309 VPWR.n1460 VPWR 0.0401341
R14310 VPWR.n1469 VPWR 0.0401341
R14311 VPWR.n1464 VPWR 0.0401341
R14312 VPWR.n1599 VPWR 0.0401341
R14313 VPWR.n1608 VPWR 0.0401341
R14314 VPWR.n1603 VPWR 0.0401341
R14315 VPWR.n934 VPWR 0.0401341
R14316 VPWR.n1692 VPWR 0.0401341
R14317 VPWR.n1688 VPWR 0.0401341
R14318 VPWR.n13 VPWR 0.0382604
R14319 VPWR.n957 VPWR 0.0382604
R14320 VPWR.n980 VPWR 0.0382604
R14321 VPWR.n1004 VPWR 0.0382604
R14322 VPWR.n1039 VPWR 0.0382604
R14323 VPWR.n1077 VPWR 0.0382604
R14324 VPWR.n1116 VPWR 0.0382604
R14325 VPWR.n1153 VPWR 0.0382604
R14326 VPWR.n39 VPWR 0.0375125
R14327 VPWR.n39 VPWR 0.0373589
R14328 VPWR.n1294 VPWR.n1287 0.0349828
R14329 VPWR.n1308 VPWR.n1305 0.0349828
R14330 VPWR.n1314 VPWR.n1311 0.0349828
R14331 VPWR.n1326 VPWR.n1323 0.0349828
R14332 VPWR.n1340 VPWR.n1337 0.0349828
R14333 VPWR.n1408 VPWR.n1272 0.0349828
R14334 VPWR.n1397 VPWR.n1273 0.0349828
R14335 VPWR.n1386 VPWR.n1274 0.0349828
R14336 VPWR.n1375 VPWR.n1275 0.0349828
R14337 VPWR.n1364 VPWR.n1347 0.0349828
R14338 VPWR.n1353 VPWR.n1348 0.0349828
R14339 VPWR.n1545 VPWR.n1542 0.0349828
R14340 VPWR.n1551 VPWR.n1548 0.0349828
R14341 VPWR.n1563 VPWR.n1560 0.0349828
R14342 VPWR.n1577 VPWR.n1574 0.0349828
R14343 VPWR.n1582 VPWR.n1579 0.0349828
R14344 VPWR.n100 VPWR.n97 0.0349828
R14345 VPWR.n126 VPWR.n121 0.0349828
R14346 VPWR.n144 VPWR.n141 0.0349828
R14347 VPWR.n148 VPWR.n147 0.0349828
R14348 VPWR.n160 VPWR.n159 0.0349828
R14349 VPWR.n178 VPWR.n175 0.0349828
R14350 VPWR.n182 VPWR.n181 0.0349828
R14351 VPWR.n194 VPWR.n193 0.0349828
R14352 VPWR.n212 VPWR.n209 0.0349828
R14353 VPWR.n216 VPWR.n215 0.0349828
R14354 VPWR.n228 VPWR.n227 0.0349828
R14355 VPWR.n246 VPWR.n243 0.0349828
R14356 VPWR.n250 VPWR.n249 0.0349828
R14357 VPWR.n262 VPWR.n261 0.0349828
R14358 VPWR.n280 VPWR.n277 0.0349828
R14359 VPWR.n284 VPWR.n283 0.0349828
R14360 VPWR.n499 VPWR 0.0341538
R14361 VPWR VPWR.n451 0.0341538
R14362 VPWR.n2544 VPWR 0.0341538
R14363 VPWR VPWR.n454 0.0341538
R14364 VPWR.n2537 VPWR 0.0341538
R14365 VPWR VPWR.n457 0.0341538
R14366 VPWR.n2530 VPWR 0.0341538
R14367 VPWR.n2510 VPWR 0.0341538
R14368 VPWR.n421 VPWR 0.0341538
R14369 VPWR.n2664 VPWR 0.0341538
R14370 VPWR.n2655 VPWR 0.0341538
R14371 VPWR.n2650 VPWR 0.0341538
R14372 VPWR.n2643 VPWR 0.0341538
R14373 VPWR.n433 VPWR 0.0341538
R14374 VPWR VPWR.n2507 0.0341538
R14375 VPWR.n2524 VPWR 0.0341538
R14376 VPWR VPWR.n2422 0.0341538
R14377 VPWR.n2423 VPWR 0.0341538
R14378 VPWR VPWR.n2430 0.0341538
R14379 VPWR VPWR.n478 0.0341538
R14380 VPWR.n2445 VPWR 0.0341538
R14381 VPWR VPWR.n476 0.0341538
R14382 VPWR.n2438 VPWR 0.0341538
R14383 VPWR.n2461 VPWR 0.0341538
R14384 VPWR.n2495 VPWR 0.0341538
R14385 VPWR.n2489 VPWR 0.0341538
R14386 VPWR VPWR.n2488 0.0341538
R14387 VPWR.n2481 VPWR 0.0341538
R14388 VPWR VPWR.n2480 0.0341538
R14389 VPWR.n2473 VPWR 0.0341538
R14390 VPWR VPWR.n464 0.0341538
R14391 VPWR VPWR.n2468 0.0341538
R14392 VPWR.n507 VPWR 0.0341538
R14393 VPWR.n2410 VPWR 0.0341538
R14394 VPWR VPWR.n504 0.0341538
R14395 VPWR.n2403 VPWR 0.0341538
R14396 VPWR VPWR.n514 0.0341538
R14397 VPWR.n2396 VPWR 0.0341538
R14398 VPWR VPWR.n517 0.0341538
R14399 VPWR.n2389 VPWR 0.0341538
R14400 VPWR.n535 VPWR 0.0341538
R14401 VPWR.n2363 VPWR 0.0341538
R14402 VPWR VPWR.n529 0.0341538
R14403 VPWR.n2370 VPWR 0.0341538
R14404 VPWR.n2375 VPWR 0.0341538
R14405 VPWR VPWR.n523 0.0341538
R14406 VPWR.n2382 VPWR 0.0341538
R14407 VPWR VPWR.n520 0.0341538
R14408 VPWR.n699 VPWR 0.0341538
R14409 VPWR VPWR.n686 0.0341538
R14410 VPWR VPWR.n561 0.0341538
R14411 VPWR.n2291 VPWR 0.0341538
R14412 VPWR VPWR.n564 0.0341538
R14413 VPWR.n2284 VPWR 0.0341538
R14414 VPWR.n559 VPWR 0.0341538
R14415 VPWR VPWR.n2308 0.0341538
R14416 VPWR.n2355 VPWR 0.0341538
R14417 VPWR.n2349 VPWR 0.0341538
R14418 VPWR VPWR.n2348 0.0341538
R14419 VPWR.n2316 VPWR 0.0341538
R14420 VPWR.n2324 VPWR 0.0341538
R14421 VPWR VPWR.n549 0.0341538
R14422 VPWR.n2331 VPWR 0.0341538
R14423 VPWR VPWR.n551 0.0341538
R14424 VPWR.n683 VPWR 0.0341538
R14425 VPWR VPWR.n630 0.0341538
R14426 VPWR.n676 VPWR 0.0341538
R14427 VPWR VPWR.n634 0.0341538
R14428 VPWR VPWR.n576 0.0341538
R14429 VPWR.n665 VPWR 0.0341538
R14430 VPWR VPWR.n637 0.0341538
R14431 VPWR.n658 VPWR 0.0341538
R14432 VPWR.n2256 VPWR 0.0341538
R14433 VPWR VPWR.n2253 0.0341538
R14434 VPWR.n2262 VPWR 0.0341538
R14435 VPWR VPWR.n579 0.0341538
R14436 VPWR.n2269 VPWR 0.0341538
R14437 VPWR.n643 VPWR 0.0341538
R14438 VPWR.n651 VPWR 0.0341538
R14439 VPWR VPWR.n640 0.0341538
R14440 VPWR.n627 VPWR 0.0341538
R14441 VPWR.n2136 VPWR 0.0341538
R14442 VPWR.n2146 VPWR 0.0341538
R14443 VPWR VPWR.n2152 0.0341538
R14444 VPWR.n2153 VPWR 0.0341538
R14445 VPWR.n2160 VPWR 0.0341538
R14446 VPWR.n2165 VPWR 0.0341538
R14447 VPWR.n2172 VPWR 0.0341538
R14448 VPWR.n2236 VPWR 0.0341538
R14449 VPWR VPWR.n587 0.0341538
R14450 VPWR.n2242 VPWR 0.0341538
R14451 VPWR VPWR.n584 0.0341538
R14452 VPWR.n2192 VPWR 0.0341538
R14453 VPWR VPWR.n603 0.0341538
R14454 VPWR.n2199 VPWR 0.0341538
R14455 VPWR.n2177 VPWR 0.0341538
R14456 VPWR VPWR.n2074 0.0341538
R14457 VPWR.n2075 VPWR 0.0341538
R14458 VPWR VPWR.n2082 0.0341538
R14459 VPWR.n2083 VPWR 0.0341538
R14460 VPWR.n2117 VPWR 0.0341538
R14461 VPWR VPWR.n2066 0.0341538
R14462 VPWR.n2110 VPWR 0.0341538
R14463 VPWR VPWR.n2091 0.0341538
R14464 VPWR.n595 VPWR 0.0341538
R14465 VPWR.n2228 VPWR 0.0341538
R14466 VPWR.n2219 VPWR 0.0341538
R14467 VPWR VPWR.n2218 0.0341538
R14468 VPWR.n2211 VPWR 0.0341538
R14469 VPWR.n602 VPWR 0.0341538
R14470 VPWR VPWR.n2094 0.0341538
R14471 VPWR.n2103 VPWR 0.0341538
R14472 VPWR.n1925 VPWR 0.0341538
R14473 VPWR.n1930 VPWR 0.0341538
R14474 VPWR.n1947 VPWR 0.0341538
R14475 VPWR VPWR.n759 0.0341538
R14476 VPWR VPWR.n710 0.0341538
R14477 VPWR.n2060 VPWR 0.0341538
R14478 VPWR VPWR.n713 0.0341538
R14479 VPWR.n2053 VPWR 0.0341538
R14480 VPWR.n2023 VPWR 0.0341538
R14481 VPWR VPWR.n731 0.0341538
R14482 VPWR.n2029 VPWR 0.0341538
R14483 VPWR.n2034 VPWR 0.0341538
R14484 VPWR VPWR.n725 0.0341538
R14485 VPWR.n2041 VPWR 0.0341538
R14486 VPWR VPWR.n719 0.0341538
R14487 VPWR.n2048 VPWR 0.0341538
R14488 VPWR.n793 VPWR 0.0341538
R14489 VPWR VPWR.n768 0.0341538
R14490 VPWR.n786 VPWR 0.0341538
R14491 VPWR VPWR.n758 0.0341538
R14492 VPWR.n779 VPWR 0.0341538
R14493 VPWR.n774 VPWR 0.0341538
R14494 VPWR.n1960 VPWR 0.0341538
R14495 VPWR VPWR.n1967 0.0341538
R14496 VPWR.n738 VPWR 0.0341538
R14497 VPWR VPWR.n742 0.0341538
R14498 VPWR.n1999 VPWR 0.0341538
R14499 VPWR VPWR.n745 0.0341538
R14500 VPWR.n2006 VPWR 0.0341538
R14501 VPWR.n1984 VPWR 0.0341538
R14502 VPWR.n1975 VPWR 0.0341538
R14503 VPWR.n1968 VPWR 0.0341538
R14504 VPWR.n800 VPWR 0.0341538
R14505 VPWR.n1912 VPWR 0.0341538
R14506 VPWR VPWR.n797 0.0341538
R14507 VPWR.n1905 VPWR 0.0341538
R14508 VPWR VPWR.n807 0.0341538
R14509 VPWR.n1898 VPWR 0.0341538
R14510 VPWR.n816 VPWR 0.0341538
R14511 VPWR.n1892 VPWR 0.0341538
R14512 VPWR.n832 VPWR 0.0341538
R14513 VPWR VPWR.n741 0.0341538
R14514 VPWR.n1871 VPWR 0.0341538
R14515 VPWR VPWR.n827 0.0341538
R14516 VPWR.n1878 VPWR 0.0341538
R14517 VPWR VPWR.n824 0.0341538
R14518 VPWR.n1885 VPWR 0.0341538
R14519 VPWR VPWR.n813 0.0341538
R14520 VPWR.n2553 VPWR 0.0341538
R14521 VPWR.n2567 VPWR 0.0341538
R14522 VPWR VPWR.n2550 0.0341538
R14523 VPWR.n2560 VPWR 0.0341538
R14524 VPWR.n2578 VPWR 0.0341538
R14525 VPWR VPWR.n2585 0.0341538
R14526 VPWR.n417 VPWR 0.0341538
R14527 VPWR VPWR.n2599 0.0341538
R14528 VPWR.n2607 VPWR 0.0341538
R14529 VPWR VPWR.n2596 0.0341538
R14530 VPWR.n2614 VPWR 0.0341538
R14531 VPWR VPWR.n434 0.0341538
R14532 VPWR.n2621 VPWR 0.0341538
R14533 VPWR VPWR.n441 0.0341538
R14534 VPWR.n2628 VPWR 0.0341538
R14535 VPWR.n2586 VPWR 0.0341538
R14536 VPWR.n1778 VPWR 0.0341538
R14537 VPWR VPWR.n1784 0.0341538
R14538 VPWR VPWR.n865 0.0341538
R14539 VPWR.n1802 VPWR 0.0341538
R14540 VPWR VPWR.n863 0.0341538
R14541 VPWR.n1795 VPWR 0.0341538
R14542 VPWR VPWR.n1818 0.0341538
R14543 VPWR.n1819 VPWR 0.0341538
R14544 VPWR.n1826 VPWR 0.0341538
R14545 VPWR.n1831 VPWR 0.0341538
R14546 VPWR.n1860 VPWR 0.0341538
R14547 VPWR.n1854 VPWR 0.0341538
R14548 VPWR VPWR.n1853 0.0341538
R14549 VPWR VPWR.n840 0.0341538
R14550 VPWR VPWR.n1846 0.0341538
R14551 VPWR.n1841 VPWR 0.0341538
R14552 VPWR.n2735 VPWR 0.0341538
R14553 VPWR VPWR.n374 0.0341538
R14554 VPWR.n2728 VPWR 0.0341538
R14555 VPWR.n2723 VPWR 0.0341538
R14556 VPWR.n2675 VPWR 0.0341538
R14557 VPWR.n2680 VPWR 0.0341538
R14558 VPWR VPWR.n408 0.0341538
R14559 VPWR.n2687 VPWR 0.0341538
R14560 VPWR.n2692 VPWR 0.0341538
R14561 VPWR VPWR.n399 0.0341538
R14562 VPWR.n2699 VPWR 0.0341538
R14563 VPWR.n2704 VPWR 0.0341538
R14564 VPWR VPWR.n390 0.0341538
R14565 VPWR.n2711 VPWR 0.0341538
R14566 VPWR.n2716 VPWR 0.0341538
R14567 VPWR VPWR.n381 0.0341538
R14568 VPWR VPWR.n873 0.0341538
R14569 VPWR.n1770 VPWR 0.0341538
R14570 VPWR VPWR.n876 0.0341538
R14571 VPWR.n1763 VPWR 0.0341538
R14572 VPWR VPWR.n885 0.0341538
R14573 VPWR.n1756 VPWR 0.0341538
R14574 VPWR.n897 VPWR 0.0341538
R14575 VPWR.n1750 VPWR 0.0341538
R14576 VPWR VPWR.n894 0.0341538
R14577 VPWR.n1743 VPWR 0.0341538
R14578 VPWR VPWR.n905 0.0341538
R14579 VPWR.n1736 VPWR 0.0341538
R14580 VPWR.n1717 VPWR 0.0341538
R14581 VPWR.n1724 VPWR 0.0341538
R14582 VPWR.n1729 VPWR 0.0341538
R14583 VPWR VPWR.n908 0.0341538
R14584 VPWR.n1189 VPWR 0.0341538
R14585 VPWR VPWR.n1195 0.0341538
R14586 VPWR.n1196 VPWR 0.0341538
R14587 VPWR.n1662 VPWR 0.0341538
R14588 VPWR VPWR.n1172 0.0341538
R14589 VPWR.n1655 VPWR 0.0341538
R14590 VPWR VPWR.n1210 0.0341538
R14591 VPWR.n1648 VPWR 0.0341538
R14592 VPWR VPWR.n1219 0.0341538
R14593 VPWR.n1641 VPWR 0.0341538
R14594 VPWR.n1635 VPWR 0.0341538
R14595 VPWR.n1615 VPWR 0.0341538
R14596 VPWR VPWR.n1701 0.0341538
R14597 VPWR.n920 VPWR 0.0341538
R14598 VPWR.n1714 VPWR 0.0341538
R14599 VPWR.n1702 VPWR 0.0341538
R14600 VPWR.n368 VPWR 0.0341538
R14601 VPWR VPWR.n293 0.0341538
R14602 VPWR.n315 VPWR 0.0341538
R14603 VPWR.n319 VPWR 0.0341538
R14604 VPWR VPWR.n312 0.0341538
R14605 VPWR.n326 VPWR 0.0341538
R14606 VPWR VPWR.n309 0.0341538
R14607 VPWR.n333 VPWR 0.0341538
R14608 VPWR VPWR.n306 0.0341538
R14609 VPWR.n340 VPWR 0.0341538
R14610 VPWR VPWR.n303 0.0341538
R14611 VPWR.n347 VPWR 0.0341538
R14612 VPWR VPWR.n300 0.0341538
R14613 VPWR.n354 VPWR 0.0341538
R14614 VPWR VPWR.n297 0.0341538
R14615 VPWR.n361 VPWR 0.0341538
R14616 VPWR.n940 VPWR 0.0341538
R14617 VPWR VPWR.n1237 0.0341538
R14618 VPWR.n1592 VPWR 0.0341538
R14619 VPWR.n1528 VPWR 0.0341538
R14620 VPWR VPWR.n1233 0.0341538
R14621 VPWR.n1520 VPWR 0.0341538
R14622 VPWR VPWR.n1518 0.0341538
R14623 VPWR.n1511 VPWR 0.0341538
R14624 VPWR.n1504 VPWR 0.0341538
R14625 VPWR.n1497 VPWR 0.0341538
R14626 VPWR.n1492 VPWR 0.0341538
R14627 VPWR.n1485 VPWR 0.0341538
R14628 VPWR VPWR.n1169 0.0341538
R14629 VPWR.n1668 VPWR 0.0341538
R14630 VPWR VPWR.n1159 0.0341538
R14631 VPWR.n1676 VPWR 0.0341538
R14632 VPWR.n2759 VPWR 0.0341538
R14633 VPWR.n2766 VPWR 0.0341538
R14634 VPWR.n2771 VPWR 0.0341538
R14635 VPWR.n2778 VPWR 0.0341538
R14636 VPWR.n2783 VPWR 0.0341538
R14637 VPWR.n2790 VPWR 0.0341538
R14638 VPWR.n2795 VPWR 0.0341538
R14639 VPWR.n2802 VPWR 0.0341538
R14640 VPWR.n2807 VPWR 0.0341538
R14641 VPWR.n2814 VPWR 0.0341538
R14642 VPWR.n2819 VPWR 0.0341538
R14643 VPWR.n2826 VPWR 0.0341538
R14644 VPWR.n2831 VPWR 0.0341538
R14645 VPWR.n2838 VPWR 0.0341538
R14646 VPWR.n2843 VPWR 0.0341538
R14647 VPWR.n2849 VPWR 0.0341538
R14648 VPWR.n2917 VPWR.n2887 0.0320292
R14649 VPWR VPWR.n22 0.03175
R14650 VPWR.n3089 VPWR 0.03175
R14651 VPWR VPWR.n3080 0.03175
R14652 VPWR VPWR.n3060 0.03175
R14653 VPWR VPWR.n3041 0.03175
R14654 VPWR VPWR.n3022 0.03175
R14655 VPWR VPWR.n2985 0.03175
R14656 VPWR VPWR.n2948 0.03175
R14657 VPWR VPWR.n2916 0.03175
R14658 VPWR.n2887 VPWR.n2886 0.0240975
R14659 VPWR.n2886 VPWR.n39 0.0240975
R14660 VPWR.n38 VPWR 0.024
R14661 VPWR.n14 VPWR 0.0239375
R14662 VPWR.n12 VPWR 0.0239375
R14663 VPWR.n958 VPWR 0.0239375
R14664 VPWR.n956 VPWR 0.0239375
R14665 VPWR.n979 VPWR 0.0239375
R14666 VPWR.n1003 VPWR 0.0239375
R14667 VPWR.n3042 VPWR 0.0239375
R14668 VPWR.n1044 VPWR 0.0226354
R14669 VPWR.n1035 VPWR 0.0226354
R14670 VPWR.n1121 VPWR 0.0226354
R14671 VPWR.n3061 VPWR 0.0226354
R14672 VPWR VPWR.n3021 0.0226354
R14673 VPWR VPWR.n2991 0.0226354
R14674 VPWR VPWR.n2953 0.0226354
R14675 VPWR.n1297 VPWR 0.0220517
R14676 VPWR VPWR.n1158 0.0220517
R14677 VPWR.n1317 VPWR 0.0220517
R14678 VPWR.n1329 VPWR 0.0220517
R14679 VPWR.n1414 VPWR 0.0220517
R14680 VPWR VPWR.n1403 0.0220517
R14681 VPWR VPWR.n1392 0.0220517
R14682 VPWR VPWR.n1381 0.0220517
R14683 VPWR VPWR.n1370 0.0220517
R14684 VPWR VPWR.n1359 0.0220517
R14685 VPWR VPWR.n1258 0.0220517
R14686 VPWR VPWR.n1539 0.0220517
R14687 VPWR.n1554 VPWR 0.0220517
R14688 VPWR.n1566 VPWR 0.0220517
R14689 VPWR VPWR.n1236 0.0220517
R14690 VPWR VPWR.n132 0.0220517
R14691 VPWR.n135 VPWR 0.0220517
R14692 VPWR VPWR.n154 0.0220517
R14693 VPWR VPWR.n166 0.0220517
R14694 VPWR.n169 VPWR 0.0220517
R14695 VPWR VPWR.n188 0.0220517
R14696 VPWR VPWR.n200 0.0220517
R14697 VPWR.n203 VPWR 0.0220517
R14698 VPWR VPWR.n222 0.0220517
R14699 VPWR VPWR.n234 0.0220517
R14700 VPWR.n237 VPWR 0.0220517
R14701 VPWR VPWR.n256 0.0220517
R14702 VPWR VPWR.n268 0.0220517
R14703 VPWR.n271 VPWR 0.0220517
R14704 VPWR.n290 VPWR 0.0220517
R14705 VPWR.n981 VPWR 0.0213333
R14706 VPWR.n1005 VPWR 0.0213333
R14707 VPWR.n1019 VPWR 0.0213333
R14708 VPWR.n1083 VPWR 0.0213333
R14709 VPWR.n1055 VPWR 0.0213333
R14710 VPWR.n1094 VPWR 0.0213333
R14711 VPWR.n1131 VPWR 0.0213333
R14712 VPWR.n3095 VPWR 0.0213333
R14713 VPWR.n3088 VPWR 0.0213333
R14714 VPWR VPWR.n3079 0.0213333
R14715 VPWR.n3081 VPWR 0.0213333
R14716 VPWR VPWR.n3059 0.0213333
R14717 VPWR VPWR.n3040 0.0213333
R14718 VPWR VPWR.n3027 0.0213333
R14719 VPWR.n2756 VPWR 0.0196917
R14720 VPWR.n2851 VPWR 0.0143889
R14721 VPWR VPWR.n19 0.0099
R14722 VPWR.n498 VPWR.n451 0.00691026
R14723 VPWR.n2544 VPWR.n453 0.00691026
R14724 VPWR.n2543 VPWR.n454 0.00691026
R14725 VPWR.n2538 VPWR.n2537 0.00691026
R14726 VPWR.n2536 VPWR.n457 0.00691026
R14727 VPWR.n2531 VPWR.n2530 0.00691026
R14728 VPWR.n2511 VPWR.n2510 0.00691026
R14729 VPWR.n2663 VPWR.n421 0.00691026
R14730 VPWR.n2664 VPWR.n420 0.00691026
R14731 VPWR.n2656 VPWR.n2655 0.00691026
R14732 VPWR.n2650 VPWR.n2649 0.00691026
R14733 VPWR.n2644 VPWR.n2643 0.00691026
R14734 VPWR.n2518 VPWR.n433 0.00691026
R14735 VPWR.n2523 VPWR.n2507 0.00691026
R14736 VPWR.n2524 VPWR.n462 0.00691026
R14737 VPWR.n2424 VPWR.n2423 0.00691026
R14738 VPWR.n2430 VPWR.n2429 0.00691026
R14739 VPWR.n2431 VPWR.n478 0.00691026
R14740 VPWR.n2445 VPWR.n480 0.00691026
R14741 VPWR.n2444 VPWR.n476 0.00691026
R14742 VPWR.n2439 VPWR.n2438 0.00691026
R14743 VPWR.n2462 VPWR.n2461 0.00691026
R14744 VPWR.n2495 VPWR.n2494 0.00691026
R14745 VPWR.n2490 VPWR.n2489 0.00691026
R14746 VPWR.n2488 VPWR.n2487 0.00691026
R14747 VPWR.n2482 VPWR.n2481 0.00691026
R14748 VPWR.n2480 VPWR.n2479 0.00691026
R14749 VPWR.n2474 VPWR.n2473 0.00691026
R14750 VPWR.n2469 VPWR.n464 0.00691026
R14751 VPWR.n2468 VPWR.n2467 0.00691026
R14752 VPWR.n2410 VPWR.n503 0.00691026
R14753 VPWR.n2409 VPWR.n504 0.00691026
R14754 VPWR.n2404 VPWR.n2403 0.00691026
R14755 VPWR.n2402 VPWR.n514 0.00691026
R14756 VPWR.n2397 VPWR.n2396 0.00691026
R14757 VPWR.n2395 VPWR.n517 0.00691026
R14758 VPWR.n2390 VPWR.n2389 0.00691026
R14759 VPWR.n538 VPWR.n535 0.00691026
R14760 VPWR.n2364 VPWR.n2363 0.00691026
R14761 VPWR.n2369 VPWR.n529 0.00691026
R14762 VPWR.n2370 VPWR.n528 0.00691026
R14763 VPWR.n2376 VPWR.n2375 0.00691026
R14764 VPWR.n2381 VPWR.n523 0.00691026
R14765 VPWR.n2383 VPWR.n2382 0.00691026
R14766 VPWR.n2388 VPWR.n520 0.00691026
R14767 VPWR.n698 VPWR.n686 0.00691026
R14768 VPWR.n693 VPWR.n561 0.00691026
R14769 VPWR.n2291 VPWR.n563 0.00691026
R14770 VPWR.n2290 VPWR.n564 0.00691026
R14771 VPWR.n2285 VPWR.n2284 0.00691026
R14772 VPWR.n573 VPWR.n559 0.00691026
R14773 VPWR.n2308 VPWR.n556 0.00691026
R14774 VPWR.n2355 VPWR.n2354 0.00691026
R14775 VPWR.n2350 VPWR.n2349 0.00691026
R14776 VPWR.n2348 VPWR.n544 0.00691026
R14777 VPWR.n2323 VPWR.n2316 0.00691026
R14778 VPWR.n2325 VPWR.n2324 0.00691026
R14779 VPWR.n2330 VPWR.n549 0.00691026
R14780 VPWR.n2331 VPWR.n553 0.00691026
R14781 VPWR.n2309 VPWR.n551 0.00691026
R14782 VPWR.n682 VPWR.n630 0.00691026
R14783 VPWR.n677 VPWR.n676 0.00691026
R14784 VPWR.n675 VPWR.n634 0.00691026
R14785 VPWR.n670 VPWR.n576 0.00691026
R14786 VPWR.n666 VPWR.n665 0.00691026
R14787 VPWR.n664 VPWR.n637 0.00691026
R14788 VPWR.n659 VPWR.n658 0.00691026
R14789 VPWR.n2257 VPWR.n2256 0.00691026
R14790 VPWR.n2261 VPWR.n2253 0.00691026
R14791 VPWR.n2263 VPWR.n2262 0.00691026
R14792 VPWR.n2268 VPWR.n579 0.00691026
R14793 VPWR.n2269 VPWR.n578 0.00691026
R14794 VPWR.n650 VPWR.n643 0.00691026
R14795 VPWR.n652 VPWR.n651 0.00691026
R14796 VPWR.n657 VPWR.n640 0.00691026
R14797 VPWR.n2137 VPWR.n2136 0.00691026
R14798 VPWR.n2146 VPWR.n2145 0.00691026
R14799 VPWR.n2152 VPWR.n616 0.00691026
R14800 VPWR.n2154 VPWR.n2153 0.00691026
R14801 VPWR.n2160 VPWR.n2159 0.00691026
R14802 VPWR.n2166 VPWR.n2165 0.00691026
R14803 VPWR.n2172 VPWR.n2171 0.00691026
R14804 VPWR.n2237 VPWR.n2236 0.00691026
R14805 VPWR.n2241 VPWR.n587 0.00691026
R14806 VPWR.n2242 VPWR.n586 0.00691026
R14807 VPWR.n2191 VPWR.n584 0.00691026
R14808 VPWR.n2193 VPWR.n2192 0.00691026
R14809 VPWR.n2198 VPWR.n603 0.00691026
R14810 VPWR.n2199 VPWR.n605 0.00691026
R14811 VPWR.n2178 VPWR.n2177 0.00691026
R14812 VPWR.n2076 VPWR.n2075 0.00691026
R14813 VPWR.n2082 VPWR.n2081 0.00691026
R14814 VPWR.n2084 VPWR.n2083 0.00691026
R14815 VPWR.n2117 VPWR.n2065 0.00691026
R14816 VPWR.n2116 VPWR.n2066 0.00691026
R14817 VPWR.n2111 VPWR.n2110 0.00691026
R14818 VPWR.n2109 VPWR.n2091 0.00691026
R14819 VPWR.n2227 VPWR.n595 0.00691026
R14820 VPWR.n2228 VPWR.n594 0.00691026
R14821 VPWR.n2220 VPWR.n2219 0.00691026
R14822 VPWR.n2218 VPWR.n2217 0.00691026
R14823 VPWR.n2212 VPWR.n2211 0.00691026
R14824 VPWR.n2097 VPWR.n602 0.00691026
R14825 VPWR.n2102 VPWR.n2094 0.00691026
R14826 VPWR.n2104 VPWR.n2103 0.00691026
R14827 VPWR.n1931 VPWR.n1930 0.00691026
R14828 VPWR.n1947 VPWR.n761 0.00691026
R14829 VPWR.n1946 VPWR.n759 0.00691026
R14830 VPWR.n1941 VPWR.n710 0.00691026
R14831 VPWR.n2060 VPWR.n712 0.00691026
R14832 VPWR.n2059 VPWR.n713 0.00691026
R14833 VPWR.n2054 VPWR.n2053 0.00691026
R14834 VPWR.n2024 VPWR.n2023 0.00691026
R14835 VPWR.n2028 VPWR.n731 0.00691026
R14836 VPWR.n2029 VPWR.n730 0.00691026
R14837 VPWR.n2035 VPWR.n2034 0.00691026
R14838 VPWR.n2040 VPWR.n725 0.00691026
R14839 VPWR.n2042 VPWR.n2041 0.00691026
R14840 VPWR.n2047 VPWR.n719 0.00691026
R14841 VPWR.n2048 VPWR.n718 0.00691026
R14842 VPWR.n792 VPWR.n768 0.00691026
R14843 VPWR.n787 VPWR.n786 0.00691026
R14844 VPWR.n785 VPWR.n758 0.00691026
R14845 VPWR.n780 VPWR.n779 0.00691026
R14846 VPWR.n778 VPWR.n774 0.00691026
R14847 VPWR.n1961 VPWR.n1960 0.00691026
R14848 VPWR.n1967 VPWR.n1966 0.00691026
R14849 VPWR.n1994 VPWR.n738 0.00691026
R14850 VPWR.n1998 VPWR.n742 0.00691026
R14851 VPWR.n2000 VPWR.n1999 0.00691026
R14852 VPWR.n2005 VPWR.n745 0.00691026
R14853 VPWR.n2006 VPWR.n744 0.00691026
R14854 VPWR.n1985 VPWR.n1984 0.00691026
R14855 VPWR.n1975 VPWR.n1974 0.00691026
R14856 VPWR.n1969 VPWR.n1968 0.00691026
R14857 VPWR.n1912 VPWR.n796 0.00691026
R14858 VPWR.n1911 VPWR.n797 0.00691026
R14859 VPWR.n1906 VPWR.n1905 0.00691026
R14860 VPWR.n1904 VPWR.n807 0.00691026
R14861 VPWR.n1899 VPWR.n1898 0.00691026
R14862 VPWR.n817 VPWR.n816 0.00691026
R14863 VPWR.n1892 VPWR.n812 0.00691026
R14864 VPWR.n833 VPWR.n832 0.00691026
R14865 VPWR.n837 VPWR.n741 0.00691026
R14866 VPWR.n1872 VPWR.n1871 0.00691026
R14867 VPWR.n1877 VPWR.n827 0.00691026
R14868 VPWR.n1879 VPWR.n1878 0.00691026
R14869 VPWR.n1884 VPWR.n824 0.00691026
R14870 VPWR.n1886 VPWR.n1885 0.00691026
R14871 VPWR.n1891 VPWR.n813 0.00691026
R14872 VPWR.n2567 VPWR.n2549 0.00691026
R14873 VPWR.n2566 VPWR.n2550 0.00691026
R14874 VPWR.n2561 VPWR.n2560 0.00691026
R14875 VPWR.n2579 VPWR.n2578 0.00691026
R14876 VPWR.n2585 VPWR.n2584 0.00691026
R14877 VPWR.n2602 VPWR.n417 0.00691026
R14878 VPWR.n2606 VPWR.n2599 0.00691026
R14879 VPWR.n2608 VPWR.n2607 0.00691026
R14880 VPWR.n2613 VPWR.n2596 0.00691026
R14881 VPWR.n2615 VPWR.n2614 0.00691026
R14882 VPWR.n2620 VPWR.n434 0.00691026
R14883 VPWR.n2622 VPWR.n2621 0.00691026
R14884 VPWR.n2627 VPWR.n441 0.00691026
R14885 VPWR.n2628 VPWR.n440 0.00691026
R14886 VPWR.n2587 VPWR.n2586 0.00691026
R14887 VPWR.n1784 VPWR.n1783 0.00691026
R14888 VPWR.n1785 VPWR.n865 0.00691026
R14889 VPWR.n1802 VPWR.n867 0.00691026
R14890 VPWR.n1801 VPWR.n863 0.00691026
R14891 VPWR.n1796 VPWR.n1795 0.00691026
R14892 VPWR.n1818 VPWR.n860 0.00691026
R14893 VPWR.n1820 VPWR.n1819 0.00691026
R14894 VPWR.n1826 VPWR.n1825 0.00691026
R14895 VPWR.n1832 VPWR.n1831 0.00691026
R14896 VPWR.n1860 VPWR.n1859 0.00691026
R14897 VPWR.n1855 VPWR.n1854 0.00691026
R14898 VPWR.n1853 VPWR.n1852 0.00691026
R14899 VPWR.n1847 VPWR.n840 0.00691026
R14900 VPWR.n1846 VPWR.n846 0.00691026
R14901 VPWR.n1841 VPWR.n1840 0.00691026
R14902 VPWR.n2734 VPWR.n374 0.00691026
R14903 VPWR.n2729 VPWR.n2728 0.00691026
R14904 VPWR.n2723 VPWR.n380 0.00691026
R14905 VPWR.n2675 VPWR.n2674 0.00691026
R14906 VPWR.n2681 VPWR.n2680 0.00691026
R14907 VPWR.n2686 VPWR.n408 0.00691026
R14908 VPWR.n2687 VPWR.n407 0.00691026
R14909 VPWR.n2693 VPWR.n2692 0.00691026
R14910 VPWR.n2698 VPWR.n399 0.00691026
R14911 VPWR.n2699 VPWR.n398 0.00691026
R14912 VPWR.n2705 VPWR.n2704 0.00691026
R14913 VPWR.n2710 VPWR.n390 0.00691026
R14914 VPWR.n2711 VPWR.n389 0.00691026
R14915 VPWR.n2717 VPWR.n2716 0.00691026
R14916 VPWR.n2722 VPWR.n381 0.00691026
R14917 VPWR.n1770 VPWR.n875 0.00691026
R14918 VPWR.n1769 VPWR.n876 0.00691026
R14919 VPWR.n1764 VPWR.n1763 0.00691026
R14920 VPWR.n1762 VPWR.n885 0.00691026
R14921 VPWR.n1757 VPWR.n1756 0.00691026
R14922 VPWR.n898 VPWR.n897 0.00691026
R14923 VPWR.n1750 VPWR.n893 0.00691026
R14924 VPWR.n1749 VPWR.n894 0.00691026
R14925 VPWR.n1744 VPWR.n1743 0.00691026
R14926 VPWR.n1742 VPWR.n905 0.00691026
R14927 VPWR.n1737 VPWR.n1736 0.00691026
R14928 VPWR.n1723 VPWR.n1717 0.00691026
R14929 VPWR.n1724 VPWR.n1716 0.00691026
R14930 VPWR.n1730 VPWR.n1729 0.00691026
R14931 VPWR.n1735 VPWR.n908 0.00691026
R14932 VPWR.n1195 VPWR.n1194 0.00691026
R14933 VPWR.n1197 VPWR.n1196 0.00691026
R14934 VPWR.n1662 VPWR.n1171 0.00691026
R14935 VPWR.n1661 VPWR.n1172 0.00691026
R14936 VPWR.n1656 VPWR.n1655 0.00691026
R14937 VPWR.n1654 VPWR.n1210 0.00691026
R14938 VPWR.n1649 VPWR.n1648 0.00691026
R14939 VPWR.n1647 VPWR.n1219 0.00691026
R14940 VPWR.n1642 VPWR.n1641 0.00691026
R14941 VPWR.n1635 VPWR.n1232 0.00691026
R14942 VPWR.n1634 VPWR.n1615 0.00691026
R14943 VPWR.n1701 VPWR.n929 0.00691026
R14944 VPWR.n1713 VPWR.n920 0.00691026
R14945 VPWR.n1714 VPWR.n919 0.00691026
R14946 VPWR.n1703 VPWR.n1702 0.00691026
R14947 VPWR.n367 VPWR.n293 0.00691026
R14948 VPWR.n318 VPWR.n315 0.00691026
R14949 VPWR.n320 VPWR.n319 0.00691026
R14950 VPWR.n325 VPWR.n312 0.00691026
R14951 VPWR.n327 VPWR.n326 0.00691026
R14952 VPWR.n332 VPWR.n309 0.00691026
R14953 VPWR.n334 VPWR.n333 0.00691026
R14954 VPWR.n339 VPWR.n306 0.00691026
R14955 VPWR.n341 VPWR.n340 0.00691026
R14956 VPWR.n346 VPWR.n303 0.00691026
R14957 VPWR.n348 VPWR.n347 0.00691026
R14958 VPWR.n353 VPWR.n300 0.00691026
R14959 VPWR.n355 VPWR.n354 0.00691026
R14960 VPWR.n360 VPWR.n297 0.00691026
R14961 VPWR.n362 VPWR.n361 0.00691026
R14962 VPWR.n1586 VPWR.n940 0.00691026
R14963 VPWR.n1590 VPWR.n1237 0.00691026
R14964 VPWR.n1592 VPWR.n1235 0.00691026
R14965 VPWR.n1529 VPWR.n1528 0.00691026
R14966 VPWR.n1534 VPWR.n1233 0.00691026
R14967 VPWR.n1521 VPWR.n1520 0.00691026
R14968 VPWR.n1518 VPWR.n1517 0.00691026
R14969 VPWR.n1512 VPWR.n1511 0.00691026
R14970 VPWR.n1504 VPWR.n1503 0.00691026
R14971 VPWR.n1498 VPWR.n1497 0.00691026
R14972 VPWR.n1492 VPWR.n1491 0.00691026
R14973 VPWR.n1486 VPWR.n1485 0.00691026
R14974 VPWR.n1280 VPWR.n1169 0.00691026
R14975 VPWR.n1669 VPWR.n1668 0.00691026
R14976 VPWR.n1674 VPWR.n1159 0.00691026
R14977 VPWR.n1676 VPWR.n1157 0.00691026
R14978 VPWR.n2760 VPWR.n2759 0.00691026
R14979 VPWR.n2766 VPWR.n2765 0.00691026
R14980 VPWR.n2772 VPWR.n2771 0.00691026
R14981 VPWR.n2778 VPWR.n2777 0.00691026
R14982 VPWR.n2784 VPWR.n2783 0.00691026
R14983 VPWR.n2790 VPWR.n2789 0.00691026
R14984 VPWR.n2796 VPWR.n2795 0.00691026
R14985 VPWR.n2802 VPWR.n2801 0.00691026
R14986 VPWR.n2808 VPWR.n2807 0.00691026
R14987 VPWR.n2814 VPWR.n2813 0.00691026
R14988 VPWR.n2820 VPWR.n2819 0.00691026
R14989 VPWR.n2826 VPWR.n2825 0.00691026
R14990 VPWR.n2832 VPWR.n2831 0.00691026
R14991 VPWR.n2838 VPWR.n2837 0.00691026
R14992 VPWR.n2844 VPWR.n2843 0.00691026
R14993 VPWR.n2849 VPWR.n2848 0.00691026
R14994 VPWR.n1581 VPWR 0.00397222
R14995 VPWR VPWR.n1575 0.00397222
R14996 VPWR.n1562 VPWR 0.00397222
R14997 VPWR.n1550 VPWR 0.00397222
R14998 VPWR VPWR.n1543 0.00397222
R14999 VPWR.n1352 VPWR 0.00397222
R15000 VPWR.n1363 VPWR 0.00397222
R15001 VPWR.n1374 VPWR 0.00397222
R15002 VPWR.n1385 VPWR 0.00397222
R15003 VPWR.n1396 VPWR 0.00397222
R15004 VPWR.n1407 VPWR 0.00397222
R15005 VPWR VPWR.n1338 0.00397222
R15006 VPWR.n1325 VPWR 0.00397222
R15007 VPWR.n1313 VPWR 0.00397222
R15008 VPWR VPWR.n1306 0.00397222
R15009 VPWR.n1293 VPWR 0.00397222
R15010 VPWR VPWR.n89 0.00397222
R15011 VPWR VPWR.n278 0.00397222
R15012 VPWR VPWR.n259 0.00397222
R15013 VPWR VPWR.n104 0.00397222
R15014 VPWR VPWR.n244 0.00397222
R15015 VPWR VPWR.n225 0.00397222
R15016 VPWR VPWR.n109 0.00397222
R15017 VPWR VPWR.n210 0.00397222
R15018 VPWR VPWR.n191 0.00397222
R15019 VPWR VPWR.n114 0.00397222
R15020 VPWR VPWR.n176 0.00397222
R15021 VPWR VPWR.n157 0.00397222
R15022 VPWR VPWR.n119 0.00397222
R15023 VPWR VPWR.n142 0.00397222
R15024 VPWR VPWR.n98 0.00397222
R15025 VPWR.n125 VPWR 0.00397222
R15026 VPWR.n1423 VPWR.n1421 0.00351282
R15027 VPWR.n1695 VPWR.n1694 0.00351282
R15028 VPWR.n936 VPWR.n932 0.00351282
R15029 VPWR.n1606 VPWR.n1605 0.00351282
R15030 VPWR.n1611 VPWR.n1610 0.00351282
R15031 VPWR.n1601 VPWR.n1230 0.00351282
R15032 VPWR.n1467 VPWR.n1466 0.00351282
R15033 VPWR.n1472 VPWR.n1471 0.00351282
R15034 VPWR.n1462 VPWR.n1458 0.00351282
R15035 VPWR.n1457 VPWR.n1453 0.00351282
R15036 VPWR.n1452 VPWR.n1448 0.00351282
R15037 VPWR.n1447 VPWR.n1443 0.00351282
R15038 VPWR.n1442 VPWR.n1438 0.00351282
R15039 VPWR.n1437 VPWR.n1433 0.00351282
R15040 VPWR.n1300 VPWR.n1299 0.00265517
R15041 VPWR.n1284 VPWR.n1283 0.00265517
R15042 VPWR.n1320 VPWR.n1319 0.00265517
R15043 VPWR.n1332 VPWR.n1331 0.00265517
R15044 VPWR.n1413 VPWR.n1411 0.00265517
R15045 VPWR.n1402 VPWR.n1400 0.00265517
R15046 VPWR.n1391 VPWR.n1389 0.00265517
R15047 VPWR.n1380 VPWR.n1378 0.00265517
R15048 VPWR.n1369 VPWR.n1367 0.00265517
R15049 VPWR.n1358 VPWR.n1356 0.00265517
R15050 VPWR.n1257 VPWR.n1255 0.00265517
R15051 VPWR.n1538 VPWR.n1536 0.00265517
R15052 VPWR.n1557 VPWR.n1556 0.00265517
R15053 VPWR.n1569 VPWR.n1568 0.00265517
R15054 VPWR.n1242 VPWR.n1241 0.00265517
R15055 VPWR.n131 VPWR.n129 0.00265517
R15056 VPWR.n138 VPWR.n137 0.00265517
R15057 VPWR.n153 VPWR.n151 0.00265517
R15058 VPWR.n165 VPWR.n163 0.00265517
R15059 VPWR.n172 VPWR.n171 0.00265517
R15060 VPWR.n187 VPWR.n185 0.00265517
R15061 VPWR.n199 VPWR.n197 0.00265517
R15062 VPWR.n206 VPWR.n205 0.00265517
R15063 VPWR.n221 VPWR.n219 0.00265517
R15064 VPWR.n233 VPWR.n231 0.00265517
R15065 VPWR.n240 VPWR.n239 0.00265517
R15066 VPWR.n255 VPWR.n253 0.00265517
R15067 VPWR.n267 VPWR.n265 0.00265517
R15068 VPWR.n274 VPWR.n273 0.00265517
R15069 VPWR.n289 VPWR.n287 0.00265517
R15070 VPWR.n1586 VPWR.n1585 0.00210256
R15071 VPWR.n1591 VPWR.n1590 0.00210256
R15072 VPWR.n1246 VPWR.n1235 0.00210256
R15073 VPWR.n1529 VPWR.n1247 0.00210256
R15074 VPWR.n1535 VPWR.n1534 0.00210256
R15075 VPWR.n1521 VPWR.n1519 0.00210256
R15076 VPWR.n1517 VPWR.n1259 0.00210256
R15077 VPWR.n1512 VPWR.n1262 0.00210256
R15078 VPWR.n1503 VPWR.n1264 0.00210256
R15079 VPWR.n1498 VPWR.n1267 0.00210256
R15080 VPWR.n1491 VPWR.n1269 0.00210256
R15081 VPWR.n1486 VPWR.n1415 0.00210256
R15082 VPWR.n1281 VPWR.n1280 0.00210256
R15083 VPWR.n1669 VPWR.n1165 0.00210256
R15084 VPWR.n1675 VPWR.n1674 0.00210256
R15085 VPWR.n2765 VPWR.n84 0.00210256
R15086 VPWR.n2772 VPWR.n81 0.00210256
R15087 VPWR.n2777 VPWR.n78 0.00210256
R15088 VPWR.n2784 VPWR.n75 0.00210256
R15089 VPWR.n2789 VPWR.n72 0.00210256
R15090 VPWR.n2796 VPWR.n69 0.00210256
R15091 VPWR.n2801 VPWR.n66 0.00210256
R15092 VPWR.n2808 VPWR.n63 0.00210256
R15093 VPWR.n2813 VPWR.n60 0.00210256
R15094 VPWR.n2820 VPWR.n57 0.00210256
R15095 VPWR.n2825 VPWR.n54 0.00210256
R15096 VPWR.n2832 VPWR.n51 0.00210256
R15097 VPWR.n2837 VPWR.n48 0.00210256
R15098 VPWR.n2844 VPWR.n45 0.00210256
R15099 VPWR.n2848 VPWR.n42 0.00210256
R15100 Iout.n1020 Iout.t72 239.927
R15101 Iout.n509 Iout.t210 239.927
R15102 Iout.n513 Iout.t175 239.927
R15103 Iout.n507 Iout.t108 239.927
R15104 Iout.n504 Iout.t114 239.927
R15105 Iout.n500 Iout.t80 239.927
R15106 Iout.n192 Iout.t43 239.927
R15107 Iout.n195 Iout.t232 239.927
R15108 Iout.n199 Iout.t169 239.927
R15109 Iout.n202 Iout.t225 239.927
R15110 Iout.n206 Iout.t56 239.927
R15111 Iout.n210 Iout.t69 239.927
R15112 Iout.n214 Iout.t128 239.927
R15113 Iout.n218 Iout.t46 239.927
R15114 Iout.n222 Iout.t233 239.927
R15115 Iout.n226 Iout.t252 239.927
R15116 Iout.n232 Iout.t136 239.927
R15117 Iout.n235 Iout.t157 239.927
R15118 Iout.n238 Iout.t15 239.927
R15119 Iout.n241 Iout.t1 239.927
R15120 Iout.n244 Iout.t221 239.927
R15121 Iout.n247 Iout.t18 239.927
R15122 Iout.n250 Iout.t238 239.927
R15123 Iout.n255 Iout.t237 239.927
R15124 Iout.n252 Iout.t212 239.927
R15125 Iout.n489 Iout.t228 239.927
R15126 Iout.n494 Iout.t197 239.927
R15127 Iout.n491 Iout.t28 239.927
R15128 Iout.n519 Iout.t250 239.927
R15129 Iout.n149 Iout.t21 239.927
R15130 Iout.n146 Iout.t33 239.927
R15131 Iout.n1010 Iout.t176 239.927
R15132 Iout.n1007 Iout.t66 239.927
R15133 Iout.n140 Iout.t68 239.927
R15134 Iout.n143 Iout.t39 239.927
R15135 Iout.n525 Iout.t27 239.927
R15136 Iout.n480 Iout.t147 239.927
R15137 Iout.n483 Iout.t192 239.927
R15138 Iout.n478 Iout.t200 239.927
R15139 Iout.n259 Iout.t198 239.927
R15140 Iout.n186 Iout.t204 239.927
R15141 Iout.n271 Iout.t65 239.927
R15142 Iout.n180 Iout.t60 239.927
R15143 Iout.n283 Iout.t140 239.927
R15144 Iout.n174 Iout.t135 239.927
R15145 Iout.n168 Iout.t22 239.927
R15146 Iout.n301 Iout.t7 239.927
R15147 Iout.n289 Iout.t215 239.927
R15148 Iout.n177 Iout.t84 239.927
R15149 Iout.n277 Iout.t154 239.927
R15150 Iout.n183 Iout.t0 239.927
R15151 Iout.n265 Iout.t144 239.927
R15152 Iout.n189 Iout.t64 239.927
R15153 Iout.n472 Iout.t53 239.927
R15154 Iout.n469 Iout.t249 239.927
R15155 Iout.n156 Iout.t178 239.927
R15156 Iout.n531 Iout.t236 239.927
R15157 Iout.n534 Iout.t105 239.927
R15158 Iout.n536 Iout.t44 239.927
R15159 Iout.n133 Iout.t26 239.927
R15160 Iout.n136 Iout.t78 239.927
R15161 Iout.n542 Iout.t161 239.927
R15162 Iout.n460 Iout.t158 239.927
R15163 Iout.n463 Iout.t63 239.927
R15164 Iout.n458 Iout.t25 239.927
R15165 Iout.n305 Iout.t118 239.927
R15166 Iout.n308 Iout.t91 239.927
R15167 Iout.n311 Iout.t222 239.927
R15168 Iout.n314 Iout.t67 239.927
R15169 Iout.n317 Iout.t8 239.927
R15170 Iout.n320 Iout.t182 239.927
R15171 Iout.n392 Iout.t104 239.927
R15172 Iout.n378 Iout.t29 239.927
R15173 Iout.n376 Iout.t223 239.927
R15174 Iout.n394 Iout.t244 239.927
R15175 Iout.n408 Iout.t16 239.927
R15176 Iout.n410 Iout.t240 239.927
R15177 Iout.n424 Iout.t152 239.927
R15178 Iout.n426 Iout.t206 239.927
R15179 Iout.n447 Iout.t226 239.927
R15180 Iout.n452 Iout.t173 239.927
R15181 Iout.n449 Iout.t184 239.927
R15182 Iout.n548 Iout.t75 239.927
R15183 Iout.n130 Iout.t234 239.927
R15184 Iout.n559 Iout.t131 239.927
R15185 Iout.n557 Iout.t231 239.927
R15186 Iout.n554 Iout.t151 239.927
R15187 Iout.n434 Iout.t194 239.927
R15188 Iout.n438 Iout.t156 239.927
R15189 Iout.n441 Iout.t76 239.927
R15190 Iout.n432 Iout.t142 239.927
R15191 Iout.n418 Iout.t132 239.927
R15192 Iout.n416 Iout.t70 239.927
R15193 Iout.n402 Iout.t55 239.927
R15194 Iout.n357 Iout.t86 239.927
R15195 Iout.n360 Iout.t37 239.927
R15196 Iout.n363 Iout.t146 239.927
R15197 Iout.n366 Iout.t30 239.927
R15198 Iout.n354 Iout.t93 239.927
R15199 Iout.n351 Iout.t224 239.927
R15200 Iout.n348 Iout.t32 239.927
R15201 Iout.n345 Iout.t229 239.927
R15202 Iout.n342 Iout.t190 239.927
R15203 Iout.n339 Iout.t141 239.927
R15204 Iout.n336 Iout.t230 239.927
R15205 Iout.n333 Iout.t41 239.927
R15206 Iout.n117 Iout.t191 239.927
R15207 Iout.n582 Iout.t235 239.927
R15208 Iout.n111 Iout.t193 239.927
R15209 Iout.n594 Iout.t34 239.927
R15210 Iout.n105 Iout.t180 239.927
R15211 Iout.n606 Iout.t203 239.927
R15212 Iout.n99 Iout.t148 239.927
R15213 Iout.n618 Iout.t255 239.927
R15214 Iout.n624 Iout.t155 239.927
R15215 Iout.n90 Iout.t52 239.927
R15216 Iout.n636 Iout.t107 239.927
R15217 Iout.n81 Iout.t186 239.927
R15218 Iout.n648 Iout.t209 239.927
R15219 Iout.n96 Iout.t126 239.927
R15220 Iout.n612 Iout.t31 239.927
R15221 Iout.n102 Iout.t35 239.927
R15222 Iout.n600 Iout.t143 239.927
R15223 Iout.n108 Iout.t153 239.927
R15224 Iout.n588 Iout.t48 239.927
R15225 Iout.n687 Iout.t89 239.927
R15226 Iout.n684 Iout.t13 239.927
R15227 Iout.n681 Iout.t167 239.927
R15228 Iout.n678 Iout.t71 239.927
R15229 Iout.n675 Iout.t199 239.927
R15230 Iout.n672 Iout.t168 239.927
R15231 Iout.n747 Iout.t51 239.927
R15232 Iout.n50 Iout.t202 239.927
R15233 Iout.n759 Iout.t139 239.927
R15234 Iout.n44 Iout.t120 239.927
R15235 Iout.n771 Iout.t165 239.927
R15236 Iout.n42 Iout.t196 239.927
R15237 Iout.n56 Iout.t100 239.927
R15238 Iout.n735 Iout.t213 239.927
R15239 Iout.n62 Iout.t119 239.927
R15240 Iout.n723 Iout.t12 239.927
R15241 Iout.n717 Iout.t134 239.927
R15242 Iout.n65 Iout.t109 239.927
R15243 Iout.n729 Iout.t217 239.927
R15244 Iout.n59 Iout.t57 239.927
R15245 Iout.n805 Iout.t205 239.927
R15246 Iout.n808 Iout.t54 239.927
R15247 Iout.n811 Iout.t211 239.927
R15248 Iout.n814 Iout.t171 239.927
R15249 Iout.n817 Iout.t40 239.927
R15250 Iout.n820 Iout.t160 239.927
R15251 Iout.n823 Iout.t42 239.927
R15252 Iout.n802 Iout.t189 239.927
R15253 Iout.n799 Iout.t50 239.927
R15254 Iout.n890 Iout.t59 239.927
R15255 Iout.n888 Iout.t137 239.927
R15256 Iout.n881 Iout.t129 239.927
R15257 Iout.n869 Iout.t117 239.927
R15258 Iout.n867 Iout.t103 239.927
R15259 Iout.n855 Iout.t185 239.927
R15260 Iout.n853 Iout.t79 239.927
R15261 Iout.n841 Iout.t251 239.927
R15262 Iout.n839 Iout.t83 239.927
R15263 Iout.n827 Iout.t208 239.927
R15264 Iout.n883 Iout.t3 239.927
R15265 Iout.n895 Iout.t162 239.927
R15266 Iout.n897 Iout.t248 239.927
R15267 Iout.n909 Iout.t216 239.927
R15268 Iout.n911 Iout.t159 239.927
R15269 Iout.n923 Iout.t125 239.927
R15270 Iout.n926 Iout.t214 239.927
R15271 Iout.n22 Iout.t116 239.927
R15272 Iout.n876 Iout.t121 239.927
R15273 Iout.n874 Iout.t106 239.927
R15274 Iout.n862 Iout.t101 239.927
R15275 Iout.n860 Iout.t17 239.927
R15276 Iout.n848 Iout.t181 239.927
R15277 Iout.n846 Iout.t45 239.927
R15278 Iout.n834 Iout.t195 239.927
R15279 Iout.n832 Iout.t246 239.927
R15280 Iout.n902 Iout.t241 239.927
R15281 Iout.n904 Iout.t87 239.927
R15282 Iout.n916 Iout.t219 239.927
R15283 Iout.n918 Iout.t11 239.927
R15284 Iout.n931 Iout.t201 239.927
R15285 Iout.n934 Iout.t207 239.927
R15286 Iout.n796 Iout.t95 239.927
R15287 Iout.n793 Iout.t94 239.927
R15288 Iout.n790 Iout.t73 239.927
R15289 Iout.n787 Iout.t20 239.927
R15290 Iout.n784 Iout.t174 239.927
R15291 Iout.n781 Iout.t218 239.927
R15292 Iout.n938 Iout.t97 239.927
R15293 Iout.n741 Iout.t4 239.927
R15294 Iout.n53 Iout.t227 239.927
R15295 Iout.n753 Iout.t110 239.927
R15296 Iout.n47 Iout.t36 239.927
R15297 Iout.n765 Iout.t150 239.927
R15298 Iout.n38 Iout.t112 239.927
R15299 Iout.n777 Iout.t58 239.927
R15300 Iout.n71 Iout.t38 239.927
R15301 Iout.n705 Iout.t123 239.927
R15302 Iout.n77 Iout.t187 239.927
R15303 Iout.n944 Iout.t5 239.927
R15304 Iout.n19 Iout.t6 239.927
R15305 Iout.n68 Iout.t61 239.927
R15306 Iout.n711 Iout.t49 239.927
R15307 Iout.n74 Iout.t138 239.927
R15308 Iout.n699 Iout.t166 239.927
R15309 Iout.n950 Iout.t243 239.927
R15310 Iout.n953 Iout.t74 239.927
R15311 Iout.n669 Iout.t98 239.927
R15312 Iout.n666 Iout.t122 239.927
R15313 Iout.n663 Iout.t62 239.927
R15314 Iout.n660 Iout.t179 239.927
R15315 Iout.n657 Iout.t113 239.927
R15316 Iout.n654 Iout.t164 239.927
R15317 Iout.n690 Iout.t188 239.927
R15318 Iout.n695 Iout.t47 239.927
R15319 Iout.n692 Iout.t163 239.927
R15320 Iout.n957 Iout.t102 239.927
R15321 Iout.n114 Iout.t10 239.927
R15322 Iout.n576 Iout.t172 239.927
R15323 Iout.n573 Iout.t19 239.927
R15324 Iout.n963 Iout.t111 239.927
R15325 Iout.n14 Iout.t14 239.927
R15326 Iout.n93 Iout.t115 239.927
R15327 Iout.n630 Iout.t82 239.927
R15328 Iout.n87 Iout.t247 239.927
R15329 Iout.n642 Iout.t23 239.927
R15330 Iout.n85 Iout.t90 239.927
R15331 Iout.n563 Iout.t85 239.927
R15332 Iout.n969 Iout.t96 239.927
R15333 Iout.n972 Iout.t24 239.927
R15334 Iout.n569 Iout.t242 239.927
R15335 Iout.n123 Iout.t239 239.927
R15336 Iout.n120 Iout.t81 239.927
R15337 Iout.n976 Iout.t177 239.927
R15338 Iout.n400 Iout.t254 239.927
R15339 Iout.n386 Iout.t99 239.927
R15340 Iout.n384 Iout.t183 239.927
R15341 Iout.n370 Iout.t77 239.927
R15342 Iout.n982 Iout.t245 239.927
R15343 Iout.n9 Iout.t92 239.927
R15344 Iout.n127 Iout.t88 239.927
R15345 Iout.n988 Iout.t253 239.927
R15346 Iout.n991 Iout.t133 239.927
R15347 Iout.n323 Iout.t130 239.927
R15348 Iout.n326 Iout.t145 239.927
R15349 Iout.n329 Iout.t2 239.927
R15350 Iout.n995 Iout.t127 239.927
R15351 Iout.n1001 Iout.t9 239.927
R15352 Iout.n4 Iout.t170 239.927
R15353 Iout.n295 Iout.t149 239.927
R15354 Iout.n172 Iout.t124 239.927
R15355 Iout.n1014 Iout.t220 239.927
R15356 Iout.n1021 Iout.n1020 7.9105
R15357 Iout.n510 Iout.n509 7.9105
R15358 Iout.n514 Iout.n513 7.9105
R15359 Iout.n508 Iout.n507 7.9105
R15360 Iout.n505 Iout.n504 7.9105
R15361 Iout.n501 Iout.n500 7.9105
R15362 Iout.n193 Iout.n192 7.9105
R15363 Iout.n196 Iout.n195 7.9105
R15364 Iout.n200 Iout.n199 7.9105
R15365 Iout.n203 Iout.n202 7.9105
R15366 Iout.n207 Iout.n206 7.9105
R15367 Iout.n211 Iout.n210 7.9105
R15368 Iout.n215 Iout.n214 7.9105
R15369 Iout.n219 Iout.n218 7.9105
R15370 Iout.n223 Iout.n222 7.9105
R15371 Iout.n227 Iout.n226 7.9105
R15372 Iout.n233 Iout.n232 7.9105
R15373 Iout.n236 Iout.n235 7.9105
R15374 Iout.n239 Iout.n238 7.9105
R15375 Iout.n242 Iout.n241 7.9105
R15376 Iout.n245 Iout.n244 7.9105
R15377 Iout.n248 Iout.n247 7.9105
R15378 Iout.n251 Iout.n250 7.9105
R15379 Iout.n256 Iout.n255 7.9105
R15380 Iout.n253 Iout.n252 7.9105
R15381 Iout.n490 Iout.n489 7.9105
R15382 Iout.n495 Iout.n494 7.9105
R15383 Iout.n492 Iout.n491 7.9105
R15384 Iout.n520 Iout.n519 7.9105
R15385 Iout.n150 Iout.n149 7.9105
R15386 Iout.n147 Iout.n146 7.9105
R15387 Iout.n1011 Iout.n1010 7.9105
R15388 Iout.n1008 Iout.n1007 7.9105
R15389 Iout.n141 Iout.n140 7.9105
R15390 Iout.n144 Iout.n143 7.9105
R15391 Iout.n526 Iout.n525 7.9105
R15392 Iout.n481 Iout.n480 7.9105
R15393 Iout.n484 Iout.n483 7.9105
R15394 Iout.n479 Iout.n478 7.9105
R15395 Iout.n260 Iout.n259 7.9105
R15396 Iout.n187 Iout.n186 7.9105
R15397 Iout.n272 Iout.n271 7.9105
R15398 Iout.n181 Iout.n180 7.9105
R15399 Iout.n284 Iout.n283 7.9105
R15400 Iout.n175 Iout.n174 7.9105
R15401 Iout.n169 Iout.n168 7.9105
R15402 Iout.n302 Iout.n301 7.9105
R15403 Iout.n290 Iout.n289 7.9105
R15404 Iout.n178 Iout.n177 7.9105
R15405 Iout.n278 Iout.n277 7.9105
R15406 Iout.n184 Iout.n183 7.9105
R15407 Iout.n266 Iout.n265 7.9105
R15408 Iout.n190 Iout.n189 7.9105
R15409 Iout.n473 Iout.n472 7.9105
R15410 Iout.n470 Iout.n469 7.9105
R15411 Iout.n157 Iout.n156 7.9105
R15412 Iout.n532 Iout.n531 7.9105
R15413 Iout.n535 Iout.n534 7.9105
R15414 Iout.n537 Iout.n536 7.9105
R15415 Iout.n134 Iout.n133 7.9105
R15416 Iout.n137 Iout.n136 7.9105
R15417 Iout.n543 Iout.n542 7.9105
R15418 Iout.n461 Iout.n460 7.9105
R15419 Iout.n464 Iout.n463 7.9105
R15420 Iout.n459 Iout.n458 7.9105
R15421 Iout.n306 Iout.n305 7.9105
R15422 Iout.n309 Iout.n308 7.9105
R15423 Iout.n312 Iout.n311 7.9105
R15424 Iout.n315 Iout.n314 7.9105
R15425 Iout.n318 Iout.n317 7.9105
R15426 Iout.n321 Iout.n320 7.9105
R15427 Iout.n393 Iout.n392 7.9105
R15428 Iout.n379 Iout.n378 7.9105
R15429 Iout.n377 Iout.n376 7.9105
R15430 Iout.n395 Iout.n394 7.9105
R15431 Iout.n409 Iout.n408 7.9105
R15432 Iout.n411 Iout.n410 7.9105
R15433 Iout.n425 Iout.n424 7.9105
R15434 Iout.n427 Iout.n426 7.9105
R15435 Iout.n448 Iout.n447 7.9105
R15436 Iout.n453 Iout.n452 7.9105
R15437 Iout.n450 Iout.n449 7.9105
R15438 Iout.n549 Iout.n548 7.9105
R15439 Iout.n131 Iout.n130 7.9105
R15440 Iout.n560 Iout.n559 7.9105
R15441 Iout.n558 Iout.n557 7.9105
R15442 Iout.n555 Iout.n554 7.9105
R15443 Iout.n435 Iout.n434 7.9105
R15444 Iout.n439 Iout.n438 7.9105
R15445 Iout.n442 Iout.n441 7.9105
R15446 Iout.n433 Iout.n432 7.9105
R15447 Iout.n419 Iout.n418 7.9105
R15448 Iout.n417 Iout.n416 7.9105
R15449 Iout.n403 Iout.n402 7.9105
R15450 Iout.n358 Iout.n357 7.9105
R15451 Iout.n361 Iout.n360 7.9105
R15452 Iout.n364 Iout.n363 7.9105
R15453 Iout.n367 Iout.n366 7.9105
R15454 Iout.n355 Iout.n354 7.9105
R15455 Iout.n352 Iout.n351 7.9105
R15456 Iout.n349 Iout.n348 7.9105
R15457 Iout.n346 Iout.n345 7.9105
R15458 Iout.n343 Iout.n342 7.9105
R15459 Iout.n340 Iout.n339 7.9105
R15460 Iout.n337 Iout.n336 7.9105
R15461 Iout.n334 Iout.n333 7.9105
R15462 Iout.n118 Iout.n117 7.9105
R15463 Iout.n583 Iout.n582 7.9105
R15464 Iout.n112 Iout.n111 7.9105
R15465 Iout.n595 Iout.n594 7.9105
R15466 Iout.n106 Iout.n105 7.9105
R15467 Iout.n607 Iout.n606 7.9105
R15468 Iout.n100 Iout.n99 7.9105
R15469 Iout.n619 Iout.n618 7.9105
R15470 Iout.n625 Iout.n624 7.9105
R15471 Iout.n91 Iout.n90 7.9105
R15472 Iout.n637 Iout.n636 7.9105
R15473 Iout.n82 Iout.n81 7.9105
R15474 Iout.n649 Iout.n648 7.9105
R15475 Iout.n97 Iout.n96 7.9105
R15476 Iout.n613 Iout.n612 7.9105
R15477 Iout.n103 Iout.n102 7.9105
R15478 Iout.n601 Iout.n600 7.9105
R15479 Iout.n109 Iout.n108 7.9105
R15480 Iout.n589 Iout.n588 7.9105
R15481 Iout.n688 Iout.n687 7.9105
R15482 Iout.n685 Iout.n684 7.9105
R15483 Iout.n682 Iout.n681 7.9105
R15484 Iout.n679 Iout.n678 7.9105
R15485 Iout.n676 Iout.n675 7.9105
R15486 Iout.n673 Iout.n672 7.9105
R15487 Iout.n748 Iout.n747 7.9105
R15488 Iout.n51 Iout.n50 7.9105
R15489 Iout.n760 Iout.n759 7.9105
R15490 Iout.n45 Iout.n44 7.9105
R15491 Iout.n772 Iout.n771 7.9105
R15492 Iout.n43 Iout.n42 7.9105
R15493 Iout.n57 Iout.n56 7.9105
R15494 Iout.n736 Iout.n735 7.9105
R15495 Iout.n63 Iout.n62 7.9105
R15496 Iout.n724 Iout.n723 7.9105
R15497 Iout.n718 Iout.n717 7.9105
R15498 Iout.n66 Iout.n65 7.9105
R15499 Iout.n730 Iout.n729 7.9105
R15500 Iout.n60 Iout.n59 7.9105
R15501 Iout.n806 Iout.n805 7.9105
R15502 Iout.n809 Iout.n808 7.9105
R15503 Iout.n812 Iout.n811 7.9105
R15504 Iout.n815 Iout.n814 7.9105
R15505 Iout.n818 Iout.n817 7.9105
R15506 Iout.n821 Iout.n820 7.9105
R15507 Iout.n824 Iout.n823 7.9105
R15508 Iout.n803 Iout.n802 7.9105
R15509 Iout.n800 Iout.n799 7.9105
R15510 Iout.n891 Iout.n890 7.9105
R15511 Iout.n889 Iout.n888 7.9105
R15512 Iout.n882 Iout.n881 7.9105
R15513 Iout.n870 Iout.n869 7.9105
R15514 Iout.n868 Iout.n867 7.9105
R15515 Iout.n856 Iout.n855 7.9105
R15516 Iout.n854 Iout.n853 7.9105
R15517 Iout.n842 Iout.n841 7.9105
R15518 Iout.n840 Iout.n839 7.9105
R15519 Iout.n828 Iout.n827 7.9105
R15520 Iout.n884 Iout.n883 7.9105
R15521 Iout.n896 Iout.n895 7.9105
R15522 Iout.n898 Iout.n897 7.9105
R15523 Iout.n910 Iout.n909 7.9105
R15524 Iout.n912 Iout.n911 7.9105
R15525 Iout.n924 Iout.n923 7.9105
R15526 Iout.n927 Iout.n926 7.9105
R15527 Iout.n23 Iout.n22 7.9105
R15528 Iout.n877 Iout.n876 7.9105
R15529 Iout.n875 Iout.n874 7.9105
R15530 Iout.n863 Iout.n862 7.9105
R15531 Iout.n861 Iout.n860 7.9105
R15532 Iout.n849 Iout.n848 7.9105
R15533 Iout.n847 Iout.n846 7.9105
R15534 Iout.n835 Iout.n834 7.9105
R15535 Iout.n833 Iout.n832 7.9105
R15536 Iout.n903 Iout.n902 7.9105
R15537 Iout.n905 Iout.n904 7.9105
R15538 Iout.n917 Iout.n916 7.9105
R15539 Iout.n919 Iout.n918 7.9105
R15540 Iout.n932 Iout.n931 7.9105
R15541 Iout.n935 Iout.n934 7.9105
R15542 Iout.n797 Iout.n796 7.9105
R15543 Iout.n794 Iout.n793 7.9105
R15544 Iout.n791 Iout.n790 7.9105
R15545 Iout.n788 Iout.n787 7.9105
R15546 Iout.n785 Iout.n784 7.9105
R15547 Iout.n782 Iout.n781 7.9105
R15548 Iout.n939 Iout.n938 7.9105
R15549 Iout.n742 Iout.n741 7.9105
R15550 Iout.n54 Iout.n53 7.9105
R15551 Iout.n754 Iout.n753 7.9105
R15552 Iout.n48 Iout.n47 7.9105
R15553 Iout.n766 Iout.n765 7.9105
R15554 Iout.n39 Iout.n38 7.9105
R15555 Iout.n778 Iout.n777 7.9105
R15556 Iout.n72 Iout.n71 7.9105
R15557 Iout.n706 Iout.n705 7.9105
R15558 Iout.n78 Iout.n77 7.9105
R15559 Iout.n945 Iout.n944 7.9105
R15560 Iout.n20 Iout.n19 7.9105
R15561 Iout.n69 Iout.n68 7.9105
R15562 Iout.n712 Iout.n711 7.9105
R15563 Iout.n75 Iout.n74 7.9105
R15564 Iout.n700 Iout.n699 7.9105
R15565 Iout.n951 Iout.n950 7.9105
R15566 Iout.n954 Iout.n953 7.9105
R15567 Iout.n670 Iout.n669 7.9105
R15568 Iout.n667 Iout.n666 7.9105
R15569 Iout.n664 Iout.n663 7.9105
R15570 Iout.n661 Iout.n660 7.9105
R15571 Iout.n658 Iout.n657 7.9105
R15572 Iout.n655 Iout.n654 7.9105
R15573 Iout.n691 Iout.n690 7.9105
R15574 Iout.n696 Iout.n695 7.9105
R15575 Iout.n693 Iout.n692 7.9105
R15576 Iout.n958 Iout.n957 7.9105
R15577 Iout.n115 Iout.n114 7.9105
R15578 Iout.n577 Iout.n576 7.9105
R15579 Iout.n574 Iout.n573 7.9105
R15580 Iout.n964 Iout.n963 7.9105
R15581 Iout.n15 Iout.n14 7.9105
R15582 Iout.n94 Iout.n93 7.9105
R15583 Iout.n631 Iout.n630 7.9105
R15584 Iout.n88 Iout.n87 7.9105
R15585 Iout.n643 Iout.n642 7.9105
R15586 Iout.n86 Iout.n85 7.9105
R15587 Iout.n564 Iout.n563 7.9105
R15588 Iout.n970 Iout.n969 7.9105
R15589 Iout.n973 Iout.n972 7.9105
R15590 Iout.n570 Iout.n569 7.9105
R15591 Iout.n124 Iout.n123 7.9105
R15592 Iout.n121 Iout.n120 7.9105
R15593 Iout.n977 Iout.n976 7.9105
R15594 Iout.n401 Iout.n400 7.9105
R15595 Iout.n387 Iout.n386 7.9105
R15596 Iout.n385 Iout.n384 7.9105
R15597 Iout.n371 Iout.n370 7.9105
R15598 Iout.n983 Iout.n982 7.9105
R15599 Iout.n10 Iout.n9 7.9105
R15600 Iout.n128 Iout.n127 7.9105
R15601 Iout.n989 Iout.n988 7.9105
R15602 Iout.n992 Iout.n991 7.9105
R15603 Iout.n324 Iout.n323 7.9105
R15604 Iout.n327 Iout.n326 7.9105
R15605 Iout.n330 Iout.n329 7.9105
R15606 Iout.n996 Iout.n995 7.9105
R15607 Iout.n1002 Iout.n1001 7.9105
R15608 Iout.n5 Iout.n4 7.9105
R15609 Iout.n296 Iout.n295 7.9105
R15610 Iout.n173 Iout.n172 7.9105
R15611 Iout.n1015 Iout.n1014 7.9105
R15612 Iout.n886 Iout.n885 3.86101
R15613 Iout.n880 Iout.n879 3.86101
R15614 Iout.n894 Iout.n893 3.86101
R15615 Iout.n872 Iout.n871 3.86101
R15616 Iout.n900 Iout.n899 3.86101
R15617 Iout.n866 Iout.n865 3.86101
R15618 Iout.n908 Iout.n907 3.86101
R15619 Iout.n858 Iout.n857 3.86101
R15620 Iout.n914 Iout.n913 3.86101
R15621 Iout.n852 Iout.n851 3.86101
R15622 Iout.n922 Iout.n921 3.86101
R15623 Iout.n844 Iout.n843 3.86101
R15624 Iout.n929 Iout.n928 3.86101
R15625 Iout.n838 Iout.n837 3.86101
R15626 Iout.n925 Iout.n21 3.86101
R15627 Iout.n830 Iout.n829 3.86101
R15628 Iout.n879 Iout.n878 3.4105
R15629 Iout.n887 Iout.n886 3.4105
R15630 Iout.n893 Iout.n892 3.4105
R15631 Iout.n798 Iout.n28 3.4105
R15632 Iout.n801 Iout.n29 3.4105
R15633 Iout.n804 Iout.n30 3.4105
R15634 Iout.n807 Iout.n31 3.4105
R15635 Iout.n873 Iout.n872 3.4105
R15636 Iout.n744 Iout.n743 3.4105
R15637 Iout.n740 Iout.n739 3.4105
R15638 Iout.n732 Iout.n731 3.4105
R15639 Iout.n728 Iout.n727 3.4105
R15640 Iout.n720 Iout.n719 3.4105
R15641 Iout.n795 Iout.n27 3.4105
R15642 Iout.n901 Iout.n900 3.4105
R15643 Iout.n722 Iout.n721 3.4105
R15644 Iout.n726 Iout.n725 3.4105
R15645 Iout.n734 Iout.n733 3.4105
R15646 Iout.n738 Iout.n737 3.4105
R15647 Iout.n746 Iout.n745 3.4105
R15648 Iout.n750 Iout.n749 3.4105
R15649 Iout.n752 Iout.n751 3.4105
R15650 Iout.n810 Iout.n32 3.4105
R15651 Iout.n865 Iout.n864 3.4105
R15652 Iout.n668 Iout.n55 3.4105
R15653 Iout.n671 Iout.n58 3.4105
R15654 Iout.n674 Iout.n61 3.4105
R15655 Iout.n677 Iout.n64 3.4105
R15656 Iout.n680 Iout.n67 3.4105
R15657 Iout.n683 Iout.n70 3.4105
R15658 Iout.n686 Iout.n73 3.4105
R15659 Iout.n714 Iout.n713 3.4105
R15660 Iout.n716 Iout.n715 3.4105
R15661 Iout.n792 Iout.n26 3.4105
R15662 Iout.n907 Iout.n906 3.4105
R15663 Iout.n587 Iout.n586 3.4105
R15664 Iout.n591 Iout.n590 3.4105
R15665 Iout.n599 Iout.n598 3.4105
R15666 Iout.n603 Iout.n602 3.4105
R15667 Iout.n611 Iout.n610 3.4105
R15668 Iout.n615 Iout.n614 3.4105
R15669 Iout.n623 Iout.n622 3.4105
R15670 Iout.n627 Iout.n626 3.4105
R15671 Iout.n665 Iout.n52 3.4105
R15672 Iout.n758 Iout.n757 3.4105
R15673 Iout.n756 Iout.n755 3.4105
R15674 Iout.n813 Iout.n33 3.4105
R15675 Iout.n859 Iout.n858 3.4105
R15676 Iout.n629 Iout.n628 3.4105
R15677 Iout.n621 Iout.n620 3.4105
R15678 Iout.n617 Iout.n616 3.4105
R15679 Iout.n609 Iout.n608 3.4105
R15680 Iout.n605 Iout.n604 3.4105
R15681 Iout.n597 Iout.n596 3.4105
R15682 Iout.n593 Iout.n592 3.4105
R15683 Iout.n585 Iout.n584 3.4105
R15684 Iout.n581 Iout.n580 3.4105
R15685 Iout.n579 Iout.n578 3.4105
R15686 Iout.n689 Iout.n76 3.4105
R15687 Iout.n710 Iout.n709 3.4105
R15688 Iout.n708 Iout.n707 3.4105
R15689 Iout.n789 Iout.n25 3.4105
R15690 Iout.n915 Iout.n914 3.4105
R15691 Iout.n572 Iout.n571 3.4105
R15692 Iout.n335 Iout.n116 3.4105
R15693 Iout.n338 Iout.n113 3.4105
R15694 Iout.n341 Iout.n110 3.4105
R15695 Iout.n344 Iout.n107 3.4105
R15696 Iout.n347 Iout.n104 3.4105
R15697 Iout.n350 Iout.n101 3.4105
R15698 Iout.n353 Iout.n98 3.4105
R15699 Iout.n356 Iout.n95 3.4105
R15700 Iout.n359 Iout.n92 3.4105
R15701 Iout.n633 Iout.n632 3.4105
R15702 Iout.n635 Iout.n634 3.4105
R15703 Iout.n662 Iout.n49 3.4105
R15704 Iout.n762 Iout.n761 3.4105
R15705 Iout.n764 Iout.n763 3.4105
R15706 Iout.n816 Iout.n34 3.4105
R15707 Iout.n851 Iout.n850 3.4105
R15708 Iout.n399 Iout.n398 3.4105
R15709 Iout.n405 Iout.n404 3.4105
R15710 Iout.n415 Iout.n414 3.4105
R15711 Iout.n421 Iout.n420 3.4105
R15712 Iout.n431 Iout.n430 3.4105
R15713 Iout.n444 Iout.n443 3.4105
R15714 Iout.n440 Iout.n159 3.4105
R15715 Iout.n437 Iout.n436 3.4105
R15716 Iout.n553 Iout.n552 3.4105
R15717 Iout.n556 Iout.n119 3.4105
R15718 Iout.n562 Iout.n561 3.4105
R15719 Iout.n568 Iout.n567 3.4105
R15720 Iout.n566 Iout.n565 3.4105
R15721 Iout.n575 Iout.n79 3.4105
R15722 Iout.n698 Iout.n697 3.4105
R15723 Iout.n702 Iout.n701 3.4105
R15724 Iout.n704 Iout.n703 3.4105
R15725 Iout.n786 Iout.n24 3.4105
R15726 Iout.n921 Iout.n920 3.4105
R15727 Iout.n129 Iout.n125 3.4105
R15728 Iout.n547 Iout.n546 3.4105
R15729 Iout.n551 Iout.n550 3.4105
R15730 Iout.n451 Iout.n158 3.4105
R15731 Iout.n455 Iout.n454 3.4105
R15732 Iout.n446 Iout.n445 3.4105
R15733 Iout.n429 Iout.n428 3.4105
R15734 Iout.n423 Iout.n422 3.4105
R15735 Iout.n413 Iout.n412 3.4105
R15736 Iout.n407 Iout.n406 3.4105
R15737 Iout.n397 Iout.n396 3.4105
R15738 Iout.n391 Iout.n390 3.4105
R15739 Iout.n389 Iout.n388 3.4105
R15740 Iout.n362 Iout.n89 3.4105
R15741 Iout.n641 Iout.n640 3.4105
R15742 Iout.n639 Iout.n638 3.4105
R15743 Iout.n659 Iout.n46 3.4105
R15744 Iout.n770 Iout.n769 3.4105
R15745 Iout.n768 Iout.n767 3.4105
R15746 Iout.n819 Iout.n35 3.4105
R15747 Iout.n845 Iout.n844 3.4105
R15748 Iout.n325 Iout.n165 3.4105
R15749 Iout.n322 Iout.n164 3.4105
R15750 Iout.n319 Iout.n163 3.4105
R15751 Iout.n316 Iout.n162 3.4105
R15752 Iout.n313 Iout.n161 3.4105
R15753 Iout.n310 Iout.n160 3.4105
R15754 Iout.n307 Iout.n155 3.4105
R15755 Iout.n457 Iout.n456 3.4105
R15756 Iout.n466 Iout.n465 3.4105
R15757 Iout.n462 Iout.n126 3.4105
R15758 Iout.n545 Iout.n544 3.4105
R15759 Iout.n541 Iout.n540 3.4105
R15760 Iout.n135 Iout.n3 3.4105
R15761 Iout.n987 Iout.n986 3.4105
R15762 Iout.n985 Iout.n984 3.4105
R15763 Iout.n122 Iout.n8 3.4105
R15764 Iout.n968 Iout.n967 3.4105
R15765 Iout.n966 Iout.n965 3.4105
R15766 Iout.n694 Iout.n13 3.4105
R15767 Iout.n949 Iout.n948 3.4105
R15768 Iout.n947 Iout.n946 3.4105
R15769 Iout.n783 Iout.n18 3.4105
R15770 Iout.n930 Iout.n929 3.4105
R15771 Iout.n1004 Iout.n1003 3.4105
R15772 Iout.n539 Iout.n538 3.4105
R15773 Iout.n533 Iout.n132 3.4105
R15774 Iout.n530 Iout.n529 3.4105
R15775 Iout.n468 Iout.n467 3.4105
R15776 Iout.n471 Iout.n153 3.4105
R15777 Iout.n475 Iout.n474 3.4105
R15778 Iout.n264 Iout.n263 3.4105
R15779 Iout.n268 Iout.n267 3.4105
R15780 Iout.n276 Iout.n275 3.4105
R15781 Iout.n280 Iout.n279 3.4105
R15782 Iout.n288 Iout.n287 3.4105
R15783 Iout.n292 Iout.n291 3.4105
R15784 Iout.n300 Iout.n299 3.4105
R15785 Iout.n328 Iout.n166 3.4105
R15786 Iout.n381 Iout.n380 3.4105
R15787 Iout.n383 Iout.n382 3.4105
R15788 Iout.n365 Iout.n83 3.4105
R15789 Iout.n645 Iout.n644 3.4105
R15790 Iout.n647 Iout.n646 3.4105
R15791 Iout.n656 Iout.n40 3.4105
R15792 Iout.n774 Iout.n773 3.4105
R15793 Iout.n776 Iout.n775 3.4105
R15794 Iout.n822 Iout.n36 3.4105
R15795 Iout.n837 Iout.n836 3.4105
R15796 Iout.n298 Iout.n297 3.4105
R15797 Iout.n294 Iout.n293 3.4105
R15798 Iout.n286 Iout.n285 3.4105
R15799 Iout.n282 Iout.n281 3.4105
R15800 Iout.n274 Iout.n273 3.4105
R15801 Iout.n270 Iout.n269 3.4105
R15802 Iout.n262 Iout.n261 3.4105
R15803 Iout.n477 Iout.n476 3.4105
R15804 Iout.n486 Iout.n485 3.4105
R15805 Iout.n482 Iout.n151 3.4105
R15806 Iout.n528 Iout.n527 3.4105
R15807 Iout.n524 Iout.n523 3.4105
R15808 Iout.n142 Iout.n138 3.4105
R15809 Iout.n1006 Iout.n1005 3.4105
R15810 Iout.n1009 Iout.n0 3.4105
R15811 Iout.n1000 Iout.n999 3.4105
R15812 Iout.n998 Iout.n997 3.4105
R15813 Iout.n990 Iout.n6 3.4105
R15814 Iout.n981 Iout.n980 3.4105
R15815 Iout.n979 Iout.n978 3.4105
R15816 Iout.n971 Iout.n11 3.4105
R15817 Iout.n962 Iout.n961 3.4105
R15818 Iout.n960 Iout.n959 3.4105
R15819 Iout.n952 Iout.n16 3.4105
R15820 Iout.n943 Iout.n942 3.4105
R15821 Iout.n941 Iout.n940 3.4105
R15822 Iout.n933 Iout.n21 3.4105
R15823 Iout.n1017 Iout.n1016 3.4105
R15824 Iout.n148 Iout.n2 3.4105
R15825 Iout.n518 Iout.n517 3.4105
R15826 Iout.n522 Iout.n521 3.4105
R15827 Iout.n493 Iout.n139 3.4105
R15828 Iout.n497 Iout.n496 3.4105
R15829 Iout.n488 Iout.n487 3.4105
R15830 Iout.n254 Iout.n154 3.4105
R15831 Iout.n258 Iout.n257 3.4105
R15832 Iout.n249 Iout.n188 3.4105
R15833 Iout.n246 Iout.n185 3.4105
R15834 Iout.n243 Iout.n182 3.4105
R15835 Iout.n240 Iout.n179 3.4105
R15836 Iout.n237 Iout.n176 3.4105
R15837 Iout.n234 Iout.n170 3.4105
R15838 Iout.n231 Iout.n230 3.4105
R15839 Iout.n171 Iout.n167 3.4105
R15840 Iout.n304 Iout.n303 3.4105
R15841 Iout.n332 Iout.n331 3.4105
R15842 Iout.n375 Iout.n374 3.4105
R15843 Iout.n373 Iout.n372 3.4105
R15844 Iout.n369 Iout.n368 3.4105
R15845 Iout.n84 Iout.n80 3.4105
R15846 Iout.n651 Iout.n650 3.4105
R15847 Iout.n653 Iout.n652 3.4105
R15848 Iout.n41 Iout.n37 3.4105
R15849 Iout.n780 Iout.n779 3.4105
R15850 Iout.n826 Iout.n825 3.4105
R15851 Iout.n831 Iout.n830 3.4105
R15852 Iout.n229 Iout.n228 3.4105
R15853 Iout.n225 Iout.n224 3.4105
R15854 Iout.n221 Iout.n220 3.4105
R15855 Iout.n217 Iout.n216 3.4105
R15856 Iout.n213 Iout.n212 3.4105
R15857 Iout.n209 Iout.n208 3.4105
R15858 Iout.n205 Iout.n204 3.4105
R15859 Iout.n201 Iout.n191 3.4105
R15860 Iout.n198 Iout.n197 3.4105
R15861 Iout.n194 Iout.n152 3.4105
R15862 Iout.n499 Iout.n498 3.4105
R15863 Iout.n503 Iout.n502 3.4105
R15864 Iout.n506 Iout.n145 3.4105
R15865 Iout.n516 Iout.n515 3.4105
R15866 Iout.n512 Iout.n511 3.4105
R15867 Iout.n1019 Iout.n1018 3.4105
R15868 Iout.n936 Iout.n23 1.43848
R15869 Iout.n936 Iout.n935 1.34612
R15870 Iout.n939 Iout.n937 1.34612
R15871 Iout.n20 Iout.n17 1.34612
R15872 Iout.n955 Iout.n954 1.34612
R15873 Iout.n958 Iout.n956 1.34612
R15874 Iout.n15 Iout.n12 1.34612
R15875 Iout.n974 Iout.n973 1.34612
R15876 Iout.n977 Iout.n975 1.34612
R15877 Iout.n10 Iout.n7 1.34612
R15878 Iout.n993 Iout.n992 1.34612
R15879 Iout.n996 Iout.n994 1.34612
R15880 Iout.n5 Iout.n1 1.34612
R15881 Iout.n1012 Iout.n1011 1.34612
R15882 Iout.n1015 Iout.n1013 1.34612
R15883 Iout.n1022 Iout.n1021 1.34612
R15884 Iout.n197 Iout.n154 0.451012
R15885 Iout.n476 Iout.n154 0.451012
R15886 Iout.n476 Iout.n475 0.451012
R15887 Iout.n475 Iout.n155 0.451012
R15888 Iout.n445 Iout.n155 0.451012
R15889 Iout.n445 Iout.n444 0.451012
R15890 Iout.n444 Iout.n107 0.451012
R15891 Iout.n604 Iout.n107 0.451012
R15892 Iout.n604 Iout.n603 0.451012
R15893 Iout.n603 Iout.n64 0.451012
R15894 Iout.n733 Iout.n64 0.451012
R15895 Iout.n733 Iout.n732 0.451012
R15896 Iout.n732 Iout.n29 0.451012
R15897 Iout.n886 Iout.n29 0.451012
R15898 Iout.n258 Iout.n191 0.451012
R15899 Iout.n262 Iout.n258 0.451012
R15900 Iout.n263 Iout.n262 0.451012
R15901 Iout.n263 Iout.n160 0.451012
R15902 Iout.n429 Iout.n160 0.451012
R15903 Iout.n430 Iout.n429 0.451012
R15904 Iout.n430 Iout.n104 0.451012
R15905 Iout.n609 Iout.n104 0.451012
R15906 Iout.n610 Iout.n609 0.451012
R15907 Iout.n610 Iout.n61 0.451012
R15908 Iout.n738 Iout.n61 0.451012
R15909 Iout.n739 Iout.n738 0.451012
R15910 Iout.n739 Iout.n30 0.451012
R15911 Iout.n879 Iout.n30 0.451012
R15912 Iout.n487 Iout.n152 0.451012
R15913 Iout.n487 Iout.n486 0.451012
R15914 Iout.n486 Iout.n153 0.451012
R15915 Iout.n456 Iout.n153 0.451012
R15916 Iout.n456 Iout.n455 0.451012
R15917 Iout.n455 Iout.n159 0.451012
R15918 Iout.n159 Iout.n110 0.451012
R15919 Iout.n597 Iout.n110 0.451012
R15920 Iout.n598 Iout.n597 0.451012
R15921 Iout.n598 Iout.n67 0.451012
R15922 Iout.n726 Iout.n67 0.451012
R15923 Iout.n727 Iout.n726 0.451012
R15924 Iout.n727 Iout.n28 0.451012
R15925 Iout.n893 Iout.n28 0.451012
R15926 Iout.n204 Iout.n188 0.451012
R15927 Iout.n269 Iout.n188 0.451012
R15928 Iout.n269 Iout.n268 0.451012
R15929 Iout.n268 Iout.n161 0.451012
R15930 Iout.n422 Iout.n161 0.451012
R15931 Iout.n422 Iout.n421 0.451012
R15932 Iout.n421 Iout.n101 0.451012
R15933 Iout.n616 Iout.n101 0.451012
R15934 Iout.n616 Iout.n615 0.451012
R15935 Iout.n615 Iout.n58 0.451012
R15936 Iout.n745 Iout.n58 0.451012
R15937 Iout.n745 Iout.n744 0.451012
R15938 Iout.n744 Iout.n31 0.451012
R15939 Iout.n872 Iout.n31 0.451012
R15940 Iout.n498 Iout.n497 0.451012
R15941 Iout.n497 Iout.n151 0.451012
R15942 Iout.n467 Iout.n151 0.451012
R15943 Iout.n467 Iout.n466 0.451012
R15944 Iout.n466 Iout.n158 0.451012
R15945 Iout.n436 Iout.n158 0.451012
R15946 Iout.n436 Iout.n113 0.451012
R15947 Iout.n592 Iout.n113 0.451012
R15948 Iout.n592 Iout.n591 0.451012
R15949 Iout.n591 Iout.n70 0.451012
R15950 Iout.n721 Iout.n70 0.451012
R15951 Iout.n721 Iout.n720 0.451012
R15952 Iout.n720 Iout.n27 0.451012
R15953 Iout.n900 Iout.n27 0.451012
R15954 Iout.n208 Iout.n185 0.451012
R15955 Iout.n274 Iout.n185 0.451012
R15956 Iout.n275 Iout.n274 0.451012
R15957 Iout.n275 Iout.n162 0.451012
R15958 Iout.n413 Iout.n162 0.451012
R15959 Iout.n414 Iout.n413 0.451012
R15960 Iout.n414 Iout.n98 0.451012
R15961 Iout.n621 Iout.n98 0.451012
R15962 Iout.n622 Iout.n621 0.451012
R15963 Iout.n622 Iout.n55 0.451012
R15964 Iout.n750 Iout.n55 0.451012
R15965 Iout.n751 Iout.n750 0.451012
R15966 Iout.n751 Iout.n32 0.451012
R15967 Iout.n865 Iout.n32 0.451012
R15968 Iout.n502 Iout.n139 0.451012
R15969 Iout.n528 Iout.n139 0.451012
R15970 Iout.n529 Iout.n528 0.451012
R15971 Iout.n529 Iout.n126 0.451012
R15972 Iout.n551 Iout.n126 0.451012
R15973 Iout.n552 Iout.n551 0.451012
R15974 Iout.n552 Iout.n116 0.451012
R15975 Iout.n585 Iout.n116 0.451012
R15976 Iout.n586 Iout.n585 0.451012
R15977 Iout.n586 Iout.n73 0.451012
R15978 Iout.n714 Iout.n73 0.451012
R15979 Iout.n715 Iout.n714 0.451012
R15980 Iout.n715 Iout.n26 0.451012
R15981 Iout.n907 Iout.n26 0.451012
R15982 Iout.n212 Iout.n182 0.451012
R15983 Iout.n281 Iout.n182 0.451012
R15984 Iout.n281 Iout.n280 0.451012
R15985 Iout.n280 Iout.n163 0.451012
R15986 Iout.n406 Iout.n163 0.451012
R15987 Iout.n406 Iout.n405 0.451012
R15988 Iout.n405 Iout.n95 0.451012
R15989 Iout.n628 Iout.n95 0.451012
R15990 Iout.n628 Iout.n627 0.451012
R15991 Iout.n627 Iout.n52 0.451012
R15992 Iout.n757 Iout.n52 0.451012
R15993 Iout.n757 Iout.n756 0.451012
R15994 Iout.n756 Iout.n33 0.451012
R15995 Iout.n858 Iout.n33 0.451012
R15996 Iout.n522 Iout.n145 0.451012
R15997 Iout.n523 Iout.n522 0.451012
R15998 Iout.n523 Iout.n132 0.451012
R15999 Iout.n545 Iout.n132 0.451012
R16000 Iout.n546 Iout.n545 0.451012
R16001 Iout.n546 Iout.n119 0.451012
R16002 Iout.n572 Iout.n119 0.451012
R16003 Iout.n580 Iout.n572 0.451012
R16004 Iout.n580 Iout.n579 0.451012
R16005 Iout.n579 Iout.n76 0.451012
R16006 Iout.n709 Iout.n76 0.451012
R16007 Iout.n709 Iout.n708 0.451012
R16008 Iout.n708 Iout.n25 0.451012
R16009 Iout.n914 Iout.n25 0.451012
R16010 Iout.n216 Iout.n179 0.451012
R16011 Iout.n286 Iout.n179 0.451012
R16012 Iout.n287 Iout.n286 0.451012
R16013 Iout.n287 Iout.n164 0.451012
R16014 Iout.n397 Iout.n164 0.451012
R16015 Iout.n398 Iout.n397 0.451012
R16016 Iout.n398 Iout.n92 0.451012
R16017 Iout.n633 Iout.n92 0.451012
R16018 Iout.n634 Iout.n633 0.451012
R16019 Iout.n634 Iout.n49 0.451012
R16020 Iout.n762 Iout.n49 0.451012
R16021 Iout.n763 Iout.n762 0.451012
R16022 Iout.n763 Iout.n34 0.451012
R16023 Iout.n851 Iout.n34 0.451012
R16024 Iout.n517 Iout.n516 0.451012
R16025 Iout.n517 Iout.n138 0.451012
R16026 Iout.n539 Iout.n138 0.451012
R16027 Iout.n540 Iout.n539 0.451012
R16028 Iout.n540 Iout.n125 0.451012
R16029 Iout.n562 Iout.n125 0.451012
R16030 Iout.n567 Iout.n562 0.451012
R16031 Iout.n567 Iout.n566 0.451012
R16032 Iout.n566 Iout.n79 0.451012
R16033 Iout.n698 Iout.n79 0.451012
R16034 Iout.n702 Iout.n698 0.451012
R16035 Iout.n703 Iout.n702 0.451012
R16036 Iout.n703 Iout.n24 0.451012
R16037 Iout.n921 Iout.n24 0.451012
R16038 Iout.n220 Iout.n176 0.451012
R16039 Iout.n293 Iout.n176 0.451012
R16040 Iout.n293 Iout.n292 0.451012
R16041 Iout.n292 Iout.n165 0.451012
R16042 Iout.n390 Iout.n165 0.451012
R16043 Iout.n390 Iout.n389 0.451012
R16044 Iout.n389 Iout.n89 0.451012
R16045 Iout.n640 Iout.n89 0.451012
R16046 Iout.n640 Iout.n639 0.451012
R16047 Iout.n639 Iout.n46 0.451012
R16048 Iout.n769 Iout.n46 0.451012
R16049 Iout.n769 Iout.n768 0.451012
R16050 Iout.n768 Iout.n35 0.451012
R16051 Iout.n844 Iout.n35 0.451012
R16052 Iout.n511 Iout.n2 0.451012
R16053 Iout.n1005 Iout.n2 0.451012
R16054 Iout.n1005 Iout.n1004 0.451012
R16055 Iout.n1004 Iout.n3 0.451012
R16056 Iout.n986 Iout.n3 0.451012
R16057 Iout.n986 Iout.n985 0.451012
R16058 Iout.n985 Iout.n8 0.451012
R16059 Iout.n967 Iout.n8 0.451012
R16060 Iout.n967 Iout.n966 0.451012
R16061 Iout.n966 Iout.n13 0.451012
R16062 Iout.n948 Iout.n13 0.451012
R16063 Iout.n948 Iout.n947 0.451012
R16064 Iout.n947 Iout.n18 0.451012
R16065 Iout.n929 Iout.n18 0.451012
R16066 Iout.n224 Iout.n170 0.451012
R16067 Iout.n298 Iout.n170 0.451012
R16068 Iout.n299 Iout.n298 0.451012
R16069 Iout.n299 Iout.n166 0.451012
R16070 Iout.n381 Iout.n166 0.451012
R16071 Iout.n382 Iout.n381 0.451012
R16072 Iout.n382 Iout.n83 0.451012
R16073 Iout.n645 Iout.n83 0.451012
R16074 Iout.n646 Iout.n645 0.451012
R16075 Iout.n646 Iout.n40 0.451012
R16076 Iout.n774 Iout.n40 0.451012
R16077 Iout.n775 Iout.n774 0.451012
R16078 Iout.n775 Iout.n36 0.451012
R16079 Iout.n837 Iout.n36 0.451012
R16080 Iout.n1018 Iout.n1017 0.451012
R16081 Iout.n1017 Iout.n0 0.451012
R16082 Iout.n999 Iout.n0 0.451012
R16083 Iout.n999 Iout.n998 0.451012
R16084 Iout.n998 Iout.n6 0.451012
R16085 Iout.n980 Iout.n6 0.451012
R16086 Iout.n980 Iout.n979 0.451012
R16087 Iout.n979 Iout.n11 0.451012
R16088 Iout.n961 Iout.n11 0.451012
R16089 Iout.n961 Iout.n960 0.451012
R16090 Iout.n960 Iout.n16 0.451012
R16091 Iout.n942 Iout.n16 0.451012
R16092 Iout.n942 Iout.n941 0.451012
R16093 Iout.n941 Iout.n21 0.451012
R16094 Iout.n230 Iout.n229 0.451012
R16095 Iout.n230 Iout.n167 0.451012
R16096 Iout.n304 Iout.n167 0.451012
R16097 Iout.n332 Iout.n304 0.451012
R16098 Iout.n374 Iout.n332 0.451012
R16099 Iout.n374 Iout.n373 0.451012
R16100 Iout.n373 Iout.n369 0.451012
R16101 Iout.n369 Iout.n80 0.451012
R16102 Iout.n651 Iout.n80 0.451012
R16103 Iout.n652 Iout.n651 0.451012
R16104 Iout.n652 Iout.n37 0.451012
R16105 Iout.n780 Iout.n37 0.451012
R16106 Iout.n826 Iout.n780 0.451012
R16107 Iout.n830 Iout.n826 0.451012
R16108 Iout.n231 Iout 0.2919
R16109 Iout.n303 Iout 0.2919
R16110 Iout Iout.n300 0.2919
R16111 Iout.n375 Iout 0.2919
R16112 Iout.n380 Iout 0.2919
R16113 Iout.n391 Iout 0.2919
R16114 Iout.n368 Iout 0.2919
R16115 Iout Iout.n365 0.2919
R16116 Iout Iout.n362 0.2919
R16117 Iout Iout.n359 0.2919
R16118 Iout.n650 Iout 0.2919
R16119 Iout Iout.n647 0.2919
R16120 Iout.n638 Iout 0.2919
R16121 Iout Iout.n635 0.2919
R16122 Iout.n626 Iout 0.2919
R16123 Iout.n41 Iout 0.2919
R16124 Iout.n773 Iout 0.2919
R16125 Iout Iout.n770 0.2919
R16126 Iout.n761 Iout 0.2919
R16127 Iout Iout.n758 0.2919
R16128 Iout.n749 Iout 0.2919
R16129 Iout.n825 Iout 0.2919
R16130 Iout Iout.n822 0.2919
R16131 Iout Iout.n819 0.2919
R16132 Iout Iout.n816 0.2919
R16133 Iout Iout.n813 0.2919
R16134 Iout Iout.n810 0.2919
R16135 Iout Iout.n807 0.2919
R16136 Iout.n829 Iout 0.2919
R16137 Iout.n838 Iout 0.2919
R16138 Iout.n843 Iout 0.2919
R16139 Iout.n852 Iout 0.2919
R16140 Iout.n857 Iout 0.2919
R16141 Iout.n866 Iout 0.2919
R16142 Iout.n871 Iout 0.2919
R16143 Iout.n880 Iout 0.2919
R16144 Iout Iout.n925 0.2919
R16145 Iout.n928 Iout 0.2919
R16146 Iout.n922 Iout 0.2919
R16147 Iout.n913 Iout 0.2919
R16148 Iout.n908 Iout 0.2919
R16149 Iout.n899 Iout 0.2919
R16150 Iout.n894 Iout 0.2919
R16151 Iout.n885 Iout 0.2919
R16152 Iout.n831 Iout 0.2919
R16153 Iout.n836 Iout 0.2919
R16154 Iout.n845 Iout 0.2919
R16155 Iout.n850 Iout 0.2919
R16156 Iout.n859 Iout 0.2919
R16157 Iout.n864 Iout 0.2919
R16158 Iout.n873 Iout 0.2919
R16159 Iout.n878 Iout 0.2919
R16160 Iout.n887 Iout 0.2919
R16161 Iout.n892 Iout 0.2919
R16162 Iout.n933 Iout 0.2919
R16163 Iout.n930 Iout 0.2919
R16164 Iout.n920 Iout 0.2919
R16165 Iout.n915 Iout 0.2919
R16166 Iout.n906 Iout 0.2919
R16167 Iout.n901 Iout 0.2919
R16168 Iout.n940 Iout 0.2919
R16169 Iout Iout.n783 0.2919
R16170 Iout Iout.n786 0.2919
R16171 Iout Iout.n789 0.2919
R16172 Iout Iout.n792 0.2919
R16173 Iout Iout.n795 0.2919
R16174 Iout Iout.n798 0.2919
R16175 Iout Iout.n801 0.2919
R16176 Iout Iout.n804 0.2919
R16177 Iout.n779 Iout 0.2919
R16178 Iout Iout.n776 0.2919
R16179 Iout.n767 Iout 0.2919
R16180 Iout Iout.n764 0.2919
R16181 Iout.n755 Iout 0.2919
R16182 Iout Iout.n752 0.2919
R16183 Iout.n743 Iout 0.2919
R16184 Iout Iout.n740 0.2919
R16185 Iout.n731 Iout 0.2919
R16186 Iout Iout.n728 0.2919
R16187 Iout.n719 Iout 0.2919
R16188 Iout Iout.n943 0.2919
R16189 Iout.n946 Iout 0.2919
R16190 Iout Iout.n704 0.2919
R16191 Iout.n707 Iout 0.2919
R16192 Iout Iout.n716 0.2919
R16193 Iout.n952 Iout 0.2919
R16194 Iout.n949 Iout 0.2919
R16195 Iout.n701 Iout 0.2919
R16196 Iout Iout.n710 0.2919
R16197 Iout.n713 Iout 0.2919
R16198 Iout Iout.n722 0.2919
R16199 Iout.n725 Iout 0.2919
R16200 Iout Iout.n734 0.2919
R16201 Iout.n737 Iout 0.2919
R16202 Iout Iout.n746 0.2919
R16203 Iout.n653 Iout 0.2919
R16204 Iout.n656 Iout 0.2919
R16205 Iout.n659 Iout 0.2919
R16206 Iout.n662 Iout 0.2919
R16207 Iout.n665 Iout 0.2919
R16208 Iout.n668 Iout 0.2919
R16209 Iout.n671 Iout 0.2919
R16210 Iout.n674 Iout 0.2919
R16211 Iout.n677 Iout 0.2919
R16212 Iout.n680 Iout 0.2919
R16213 Iout.n683 Iout 0.2919
R16214 Iout.n686 Iout 0.2919
R16215 Iout.n959 Iout 0.2919
R16216 Iout Iout.n694 0.2919
R16217 Iout.n697 Iout 0.2919
R16218 Iout.n689 Iout 0.2919
R16219 Iout Iout.n962 0.2919
R16220 Iout.n965 Iout 0.2919
R16221 Iout Iout.n575 0.2919
R16222 Iout.n578 Iout 0.2919
R16223 Iout Iout.n587 0.2919
R16224 Iout.n590 Iout 0.2919
R16225 Iout Iout.n599 0.2919
R16226 Iout.n602 Iout 0.2919
R16227 Iout Iout.n611 0.2919
R16228 Iout.n614 Iout 0.2919
R16229 Iout Iout.n623 0.2919
R16230 Iout.n84 Iout 0.2919
R16231 Iout.n644 Iout 0.2919
R16232 Iout Iout.n641 0.2919
R16233 Iout.n632 Iout 0.2919
R16234 Iout Iout.n629 0.2919
R16235 Iout.n620 Iout 0.2919
R16236 Iout Iout.n617 0.2919
R16237 Iout.n608 Iout 0.2919
R16238 Iout Iout.n605 0.2919
R16239 Iout.n596 Iout 0.2919
R16240 Iout Iout.n593 0.2919
R16241 Iout.n584 Iout 0.2919
R16242 Iout Iout.n581 0.2919
R16243 Iout.n971 Iout 0.2919
R16244 Iout.n968 Iout 0.2919
R16245 Iout.n565 Iout 0.2919
R16246 Iout.n978 Iout 0.2919
R16247 Iout Iout.n122 0.2919
R16248 Iout Iout.n568 0.2919
R16249 Iout.n571 Iout 0.2919
R16250 Iout Iout.n335 0.2919
R16251 Iout Iout.n338 0.2919
R16252 Iout Iout.n341 0.2919
R16253 Iout Iout.n344 0.2919
R16254 Iout Iout.n347 0.2919
R16255 Iout Iout.n350 0.2919
R16256 Iout Iout.n353 0.2919
R16257 Iout Iout.n356 0.2919
R16258 Iout.n372 Iout 0.2919
R16259 Iout.n383 Iout 0.2919
R16260 Iout.n388 Iout 0.2919
R16261 Iout.n399 Iout 0.2919
R16262 Iout.n404 Iout 0.2919
R16263 Iout.n415 Iout 0.2919
R16264 Iout.n420 Iout 0.2919
R16265 Iout.n431 Iout 0.2919
R16266 Iout.n443 Iout 0.2919
R16267 Iout Iout.n440 0.2919
R16268 Iout Iout.n437 0.2919
R16269 Iout.n553 Iout 0.2919
R16270 Iout.n556 Iout 0.2919
R16271 Iout.n561 Iout 0.2919
R16272 Iout Iout.n981 0.2919
R16273 Iout.n984 Iout 0.2919
R16274 Iout.n990 Iout 0.2919
R16275 Iout.n987 Iout 0.2919
R16276 Iout Iout.n129 0.2919
R16277 Iout Iout.n547 0.2919
R16278 Iout.n550 Iout 0.2919
R16279 Iout Iout.n451 0.2919
R16280 Iout.n454 Iout 0.2919
R16281 Iout.n446 Iout 0.2919
R16282 Iout.n428 Iout 0.2919
R16283 Iout.n423 Iout 0.2919
R16284 Iout.n412 Iout 0.2919
R16285 Iout.n407 Iout 0.2919
R16286 Iout.n396 Iout 0.2919
R16287 Iout.n331 Iout 0.2919
R16288 Iout Iout.n328 0.2919
R16289 Iout Iout.n325 0.2919
R16290 Iout Iout.n322 0.2919
R16291 Iout Iout.n319 0.2919
R16292 Iout Iout.n316 0.2919
R16293 Iout Iout.n313 0.2919
R16294 Iout Iout.n310 0.2919
R16295 Iout Iout.n307 0.2919
R16296 Iout.n457 Iout 0.2919
R16297 Iout.n465 Iout 0.2919
R16298 Iout Iout.n462 0.2919
R16299 Iout.n544 Iout 0.2919
R16300 Iout Iout.n541 0.2919
R16301 Iout Iout.n135 0.2919
R16302 Iout.n997 Iout 0.2919
R16303 Iout Iout.n1000 0.2919
R16304 Iout.n1003 Iout 0.2919
R16305 Iout.n538 Iout 0.2919
R16306 Iout.n533 Iout 0.2919
R16307 Iout.n530 Iout 0.2919
R16308 Iout Iout.n468 0.2919
R16309 Iout Iout.n471 0.2919
R16310 Iout.n474 Iout 0.2919
R16311 Iout Iout.n264 0.2919
R16312 Iout.n267 Iout 0.2919
R16313 Iout Iout.n276 0.2919
R16314 Iout.n279 Iout 0.2919
R16315 Iout Iout.n288 0.2919
R16316 Iout.n291 Iout 0.2919
R16317 Iout.n171 Iout 0.2919
R16318 Iout.n297 Iout 0.2919
R16319 Iout Iout.n294 0.2919
R16320 Iout.n285 Iout 0.2919
R16321 Iout Iout.n282 0.2919
R16322 Iout.n273 Iout 0.2919
R16323 Iout Iout.n270 0.2919
R16324 Iout.n261 Iout 0.2919
R16325 Iout.n477 Iout 0.2919
R16326 Iout.n485 Iout 0.2919
R16327 Iout Iout.n482 0.2919
R16328 Iout.n527 Iout 0.2919
R16329 Iout Iout.n524 0.2919
R16330 Iout Iout.n142 0.2919
R16331 Iout.n1006 Iout 0.2919
R16332 Iout.n1009 Iout 0.2919
R16333 Iout.n1016 Iout 0.2919
R16334 Iout Iout.n148 0.2919
R16335 Iout Iout.n518 0.2919
R16336 Iout.n521 Iout 0.2919
R16337 Iout Iout.n493 0.2919
R16338 Iout.n496 Iout 0.2919
R16339 Iout.n488 Iout 0.2919
R16340 Iout Iout.n254 0.2919
R16341 Iout.n257 Iout 0.2919
R16342 Iout.n249 Iout 0.2919
R16343 Iout.n246 Iout 0.2919
R16344 Iout.n243 Iout 0.2919
R16345 Iout.n240 Iout 0.2919
R16346 Iout.n237 Iout 0.2919
R16347 Iout.n234 Iout 0.2919
R16348 Iout.n228 Iout 0.2919
R16349 Iout Iout.n225 0.2919
R16350 Iout Iout.n221 0.2919
R16351 Iout Iout.n217 0.2919
R16352 Iout Iout.n213 0.2919
R16353 Iout Iout.n209 0.2919
R16354 Iout Iout.n205 0.2919
R16355 Iout Iout.n201 0.2919
R16356 Iout Iout.n198 0.2919
R16357 Iout Iout.n194 0.2919
R16358 Iout.n499 Iout 0.2919
R16359 Iout.n503 Iout 0.2919
R16360 Iout.n506 Iout 0.2919
R16361 Iout.n515 Iout 0.2919
R16362 Iout Iout.n512 0.2919
R16363 Iout.n1019 Iout 0.2919
R16364 Iout.n1013 Iout.n1012 0.092855
R16365 Iout.n1012 Iout.n1 0.092855
R16366 Iout.n994 Iout.n1 0.092855
R16367 Iout.n994 Iout.n993 0.092855
R16368 Iout.n993 Iout.n7 0.092855
R16369 Iout.n975 Iout.n7 0.092855
R16370 Iout.n975 Iout.n974 0.092855
R16371 Iout.n974 Iout.n12 0.092855
R16372 Iout.n956 Iout.n12 0.092855
R16373 Iout.n956 Iout.n955 0.092855
R16374 Iout.n955 Iout.n17 0.092855
R16375 Iout.n937 Iout.n17 0.092855
R16376 Iout.n937 Iout.n936 0.092855
R16377 Iout.n197 Iout 0.0818902
R16378 Iout.n191 Iout 0.0818902
R16379 Iout.n152 Iout 0.0818902
R16380 Iout.n204 Iout 0.0818902
R16381 Iout.n498 Iout 0.0818902
R16382 Iout.n208 Iout 0.0818902
R16383 Iout.n502 Iout 0.0818902
R16384 Iout.n212 Iout 0.0818902
R16385 Iout.n145 Iout 0.0818902
R16386 Iout.n216 Iout 0.0818902
R16387 Iout.n516 Iout 0.0818902
R16388 Iout.n220 Iout 0.0818902
R16389 Iout.n511 Iout 0.0818902
R16390 Iout.n224 Iout 0.0818902
R16391 Iout.n1018 Iout 0.0818902
R16392 Iout.n229 Iout 0.0818902
R16393 Iout.n1013 Iout 0.072645
R16394 Iout.n302 Iout 0.0532071
R16395 Iout Iout.n377 0.0532071
R16396 Iout.n379 Iout 0.0532071
R16397 Iout.n367 Iout 0.0532071
R16398 Iout.n364 Iout 0.0532071
R16399 Iout.n361 Iout 0.0532071
R16400 Iout.n649 Iout 0.0532071
R16401 Iout Iout.n82 0.0532071
R16402 Iout.n637 Iout 0.0532071
R16403 Iout Iout.n91 0.0532071
R16404 Iout Iout.n43 0.0532071
R16405 Iout.n772 Iout 0.0532071
R16406 Iout Iout.n45 0.0532071
R16407 Iout.n760 Iout 0.0532071
R16408 Iout Iout.n51 0.0532071
R16409 Iout.n824 Iout 0.0532071
R16410 Iout.n821 Iout 0.0532071
R16411 Iout.n818 Iout 0.0532071
R16412 Iout.n815 Iout 0.0532071
R16413 Iout.n812 Iout 0.0532071
R16414 Iout.n809 Iout 0.0532071
R16415 Iout.n828 Iout 0.0532071
R16416 Iout Iout.n840 0.0532071
R16417 Iout.n842 Iout 0.0532071
R16418 Iout Iout.n854 0.0532071
R16419 Iout.n856 Iout 0.0532071
R16420 Iout Iout.n868 0.0532071
R16421 Iout.n870 Iout 0.0532071
R16422 Iout.n927 Iout 0.0532071
R16423 Iout Iout.n924 0.0532071
R16424 Iout.n912 Iout 0.0532071
R16425 Iout Iout.n910 0.0532071
R16426 Iout.n898 Iout 0.0532071
R16427 Iout Iout.n896 0.0532071
R16428 Iout.n884 Iout 0.0532071
R16429 Iout Iout.n882 0.0532071
R16430 Iout Iout.n833 0.0532071
R16431 Iout.n835 Iout 0.0532071
R16432 Iout Iout.n847 0.0532071
R16433 Iout.n849 Iout 0.0532071
R16434 Iout Iout.n861 0.0532071
R16435 Iout.n863 Iout 0.0532071
R16436 Iout Iout.n875 0.0532071
R16437 Iout.n877 Iout 0.0532071
R16438 Iout Iout.n889 0.0532071
R16439 Iout Iout.n932 0.0532071
R16440 Iout.n919 Iout 0.0532071
R16441 Iout Iout.n917 0.0532071
R16442 Iout.n905 Iout 0.0532071
R16443 Iout Iout.n903 0.0532071
R16444 Iout.n891 Iout 0.0532071
R16445 Iout.n782 Iout 0.0532071
R16446 Iout.n785 Iout 0.0532071
R16447 Iout.n788 Iout 0.0532071
R16448 Iout.n791 Iout 0.0532071
R16449 Iout.n794 Iout 0.0532071
R16450 Iout.n797 Iout 0.0532071
R16451 Iout.n800 Iout 0.0532071
R16452 Iout.n803 Iout 0.0532071
R16453 Iout.n806 Iout 0.0532071
R16454 Iout.n778 Iout 0.0532071
R16455 Iout Iout.n39 0.0532071
R16456 Iout.n766 Iout 0.0532071
R16457 Iout Iout.n48 0.0532071
R16458 Iout.n754 Iout 0.0532071
R16459 Iout Iout.n54 0.0532071
R16460 Iout.n742 Iout 0.0532071
R16461 Iout Iout.n60 0.0532071
R16462 Iout.n730 Iout 0.0532071
R16463 Iout Iout.n66 0.0532071
R16464 Iout.n945 Iout 0.0532071
R16465 Iout.n78 Iout 0.0532071
R16466 Iout.n706 Iout 0.0532071
R16467 Iout Iout.n72 0.0532071
R16468 Iout.n718 Iout 0.0532071
R16469 Iout Iout.n951 0.0532071
R16470 Iout.n700 Iout 0.0532071
R16471 Iout Iout.n75 0.0532071
R16472 Iout.n712 Iout 0.0532071
R16473 Iout Iout.n69 0.0532071
R16474 Iout.n724 Iout 0.0532071
R16475 Iout Iout.n63 0.0532071
R16476 Iout.n736 Iout 0.0532071
R16477 Iout Iout.n57 0.0532071
R16478 Iout.n748 Iout 0.0532071
R16479 Iout Iout.n655 0.0532071
R16480 Iout Iout.n658 0.0532071
R16481 Iout Iout.n661 0.0532071
R16482 Iout Iout.n664 0.0532071
R16483 Iout Iout.n667 0.0532071
R16484 Iout Iout.n670 0.0532071
R16485 Iout Iout.n673 0.0532071
R16486 Iout Iout.n676 0.0532071
R16487 Iout Iout.n679 0.0532071
R16488 Iout Iout.n682 0.0532071
R16489 Iout Iout.n685 0.0532071
R16490 Iout.n693 Iout 0.0532071
R16491 Iout.n696 Iout 0.0532071
R16492 Iout Iout.n691 0.0532071
R16493 Iout Iout.n688 0.0532071
R16494 Iout.n964 Iout 0.0532071
R16495 Iout.n574 Iout 0.0532071
R16496 Iout.n577 Iout 0.0532071
R16497 Iout Iout.n115 0.0532071
R16498 Iout.n589 Iout 0.0532071
R16499 Iout Iout.n109 0.0532071
R16500 Iout.n601 Iout 0.0532071
R16501 Iout Iout.n103 0.0532071
R16502 Iout.n613 Iout 0.0532071
R16503 Iout Iout.n97 0.0532071
R16504 Iout.n625 Iout 0.0532071
R16505 Iout Iout.n86 0.0532071
R16506 Iout.n643 Iout 0.0532071
R16507 Iout Iout.n88 0.0532071
R16508 Iout.n631 Iout 0.0532071
R16509 Iout Iout.n94 0.0532071
R16510 Iout.n619 Iout 0.0532071
R16511 Iout Iout.n100 0.0532071
R16512 Iout.n607 Iout 0.0532071
R16513 Iout Iout.n106 0.0532071
R16514 Iout.n595 Iout 0.0532071
R16515 Iout Iout.n112 0.0532071
R16516 Iout.n583 Iout 0.0532071
R16517 Iout Iout.n970 0.0532071
R16518 Iout.n564 Iout 0.0532071
R16519 Iout Iout.n118 0.0532071
R16520 Iout.n121 Iout 0.0532071
R16521 Iout.n124 Iout 0.0532071
R16522 Iout.n570 Iout 0.0532071
R16523 Iout.n334 Iout 0.0532071
R16524 Iout.n337 Iout 0.0532071
R16525 Iout.n340 Iout 0.0532071
R16526 Iout.n343 Iout 0.0532071
R16527 Iout.n346 Iout 0.0532071
R16528 Iout.n349 Iout 0.0532071
R16529 Iout.n352 Iout 0.0532071
R16530 Iout.n355 Iout 0.0532071
R16531 Iout.n358 Iout 0.0532071
R16532 Iout.n371 Iout 0.0532071
R16533 Iout Iout.n385 0.0532071
R16534 Iout.n387 Iout 0.0532071
R16535 Iout Iout.n401 0.0532071
R16536 Iout.n403 Iout 0.0532071
R16537 Iout Iout.n417 0.0532071
R16538 Iout.n419 Iout 0.0532071
R16539 Iout Iout.n433 0.0532071
R16540 Iout.n442 Iout 0.0532071
R16541 Iout.n439 Iout 0.0532071
R16542 Iout.n435 Iout 0.0532071
R16543 Iout Iout.n555 0.0532071
R16544 Iout Iout.n558 0.0532071
R16545 Iout.n983 Iout 0.0532071
R16546 Iout.n560 Iout 0.0532071
R16547 Iout Iout.n989 0.0532071
R16548 Iout.n128 Iout 0.0532071
R16549 Iout.n131 Iout 0.0532071
R16550 Iout.n549 Iout 0.0532071
R16551 Iout.n450 Iout 0.0532071
R16552 Iout.n453 Iout 0.0532071
R16553 Iout Iout.n448 0.0532071
R16554 Iout.n427 Iout 0.0532071
R16555 Iout Iout.n425 0.0532071
R16556 Iout.n411 Iout 0.0532071
R16557 Iout Iout.n409 0.0532071
R16558 Iout.n395 Iout 0.0532071
R16559 Iout Iout.n393 0.0532071
R16560 Iout.n330 Iout 0.0532071
R16561 Iout.n327 Iout 0.0532071
R16562 Iout.n324 Iout 0.0532071
R16563 Iout.n321 Iout 0.0532071
R16564 Iout.n318 Iout 0.0532071
R16565 Iout.n315 Iout 0.0532071
R16566 Iout.n312 Iout 0.0532071
R16567 Iout.n309 Iout 0.0532071
R16568 Iout.n306 Iout 0.0532071
R16569 Iout Iout.n459 0.0532071
R16570 Iout.n464 Iout 0.0532071
R16571 Iout.n461 Iout 0.0532071
R16572 Iout.n543 Iout 0.0532071
R16573 Iout.n137 Iout 0.0532071
R16574 Iout.n134 Iout 0.0532071
R16575 Iout.n1002 Iout 0.0532071
R16576 Iout.n537 Iout 0.0532071
R16577 Iout Iout.n535 0.0532071
R16578 Iout Iout.n532 0.0532071
R16579 Iout.n157 Iout 0.0532071
R16580 Iout.n470 Iout 0.0532071
R16581 Iout.n473 Iout 0.0532071
R16582 Iout.n190 Iout 0.0532071
R16583 Iout.n266 Iout 0.0532071
R16584 Iout Iout.n184 0.0532071
R16585 Iout.n278 Iout 0.0532071
R16586 Iout Iout.n178 0.0532071
R16587 Iout.n290 Iout 0.0532071
R16588 Iout Iout.n169 0.0532071
R16589 Iout Iout.n173 0.0532071
R16590 Iout.n296 Iout 0.0532071
R16591 Iout Iout.n175 0.0532071
R16592 Iout.n284 Iout 0.0532071
R16593 Iout Iout.n181 0.0532071
R16594 Iout.n272 Iout 0.0532071
R16595 Iout Iout.n187 0.0532071
R16596 Iout.n260 Iout 0.0532071
R16597 Iout Iout.n479 0.0532071
R16598 Iout.n484 Iout 0.0532071
R16599 Iout.n481 Iout 0.0532071
R16600 Iout.n526 Iout 0.0532071
R16601 Iout.n144 Iout 0.0532071
R16602 Iout.n141 Iout 0.0532071
R16603 Iout Iout.n1008 0.0532071
R16604 Iout.n147 Iout 0.0532071
R16605 Iout.n150 Iout 0.0532071
R16606 Iout.n520 Iout 0.0532071
R16607 Iout.n492 Iout 0.0532071
R16608 Iout.n495 Iout 0.0532071
R16609 Iout Iout.n490 0.0532071
R16610 Iout.n253 Iout 0.0532071
R16611 Iout.n256 Iout 0.0532071
R16612 Iout Iout.n251 0.0532071
R16613 Iout Iout.n248 0.0532071
R16614 Iout Iout.n245 0.0532071
R16615 Iout Iout.n242 0.0532071
R16616 Iout Iout.n239 0.0532071
R16617 Iout Iout.n236 0.0532071
R16618 Iout Iout.n233 0.0532071
R16619 Iout.n227 Iout 0.0532071
R16620 Iout.n223 Iout 0.0532071
R16621 Iout.n219 Iout 0.0532071
R16622 Iout.n215 Iout 0.0532071
R16623 Iout.n211 Iout 0.0532071
R16624 Iout.n207 Iout 0.0532071
R16625 Iout.n203 Iout 0.0532071
R16626 Iout.n200 Iout 0.0532071
R16627 Iout.n196 Iout 0.0532071
R16628 Iout.n193 Iout 0.0532071
R16629 Iout Iout.n501 0.0532071
R16630 Iout Iout.n505 0.0532071
R16631 Iout Iout.n508 0.0532071
R16632 Iout.n514 Iout 0.0532071
R16633 Iout.n510 Iout 0.0532071
R16634 Iout.n1020 Iout 0.03925
R16635 Iout.n509 Iout 0.03925
R16636 Iout.n513 Iout 0.03925
R16637 Iout.n507 Iout 0.03925
R16638 Iout.n504 Iout 0.03925
R16639 Iout.n500 Iout 0.03925
R16640 Iout.n192 Iout 0.03925
R16641 Iout.n195 Iout 0.03925
R16642 Iout.n199 Iout 0.03925
R16643 Iout.n202 Iout 0.03925
R16644 Iout.n206 Iout 0.03925
R16645 Iout.n210 Iout 0.03925
R16646 Iout.n214 Iout 0.03925
R16647 Iout.n218 Iout 0.03925
R16648 Iout.n222 Iout 0.03925
R16649 Iout.n226 Iout 0.03925
R16650 Iout.n232 Iout 0.03925
R16651 Iout.n235 Iout 0.03925
R16652 Iout.n238 Iout 0.03925
R16653 Iout.n241 Iout 0.03925
R16654 Iout.n244 Iout 0.03925
R16655 Iout.n247 Iout 0.03925
R16656 Iout.n250 Iout 0.03925
R16657 Iout.n255 Iout 0.03925
R16658 Iout.n252 Iout 0.03925
R16659 Iout.n489 Iout 0.03925
R16660 Iout.n494 Iout 0.03925
R16661 Iout.n491 Iout 0.03925
R16662 Iout.n519 Iout 0.03925
R16663 Iout.n149 Iout 0.03925
R16664 Iout.n146 Iout 0.03925
R16665 Iout.n1010 Iout 0.03925
R16666 Iout.n1007 Iout 0.03925
R16667 Iout.n140 Iout 0.03925
R16668 Iout.n143 Iout 0.03925
R16669 Iout.n525 Iout 0.03925
R16670 Iout.n480 Iout 0.03925
R16671 Iout.n483 Iout 0.03925
R16672 Iout.n478 Iout 0.03925
R16673 Iout.n259 Iout 0.03925
R16674 Iout.n186 Iout 0.03925
R16675 Iout.n271 Iout 0.03925
R16676 Iout.n180 Iout 0.03925
R16677 Iout.n283 Iout 0.03925
R16678 Iout.n174 Iout 0.03925
R16679 Iout.n168 Iout 0.03925
R16680 Iout.n301 Iout 0.03925
R16681 Iout.n289 Iout 0.03925
R16682 Iout.n177 Iout 0.03925
R16683 Iout.n277 Iout 0.03925
R16684 Iout.n183 Iout 0.03925
R16685 Iout.n265 Iout 0.03925
R16686 Iout.n189 Iout 0.03925
R16687 Iout.n472 Iout 0.03925
R16688 Iout.n469 Iout 0.03925
R16689 Iout.n156 Iout 0.03925
R16690 Iout.n531 Iout 0.03925
R16691 Iout.n534 Iout 0.03925
R16692 Iout.n536 Iout 0.03925
R16693 Iout.n133 Iout 0.03925
R16694 Iout.n136 Iout 0.03925
R16695 Iout.n542 Iout 0.03925
R16696 Iout.n460 Iout 0.03925
R16697 Iout.n463 Iout 0.03925
R16698 Iout.n458 Iout 0.03925
R16699 Iout.n305 Iout 0.03925
R16700 Iout.n308 Iout 0.03925
R16701 Iout.n311 Iout 0.03925
R16702 Iout.n314 Iout 0.03925
R16703 Iout.n317 Iout 0.03925
R16704 Iout.n320 Iout 0.03925
R16705 Iout.n392 Iout 0.03925
R16706 Iout.n378 Iout 0.03925
R16707 Iout.n376 Iout 0.03925
R16708 Iout.n394 Iout 0.03925
R16709 Iout.n408 Iout 0.03925
R16710 Iout.n410 Iout 0.03925
R16711 Iout.n424 Iout 0.03925
R16712 Iout.n426 Iout 0.03925
R16713 Iout.n447 Iout 0.03925
R16714 Iout.n452 Iout 0.03925
R16715 Iout.n449 Iout 0.03925
R16716 Iout.n548 Iout 0.03925
R16717 Iout.n130 Iout 0.03925
R16718 Iout.n559 Iout 0.03925
R16719 Iout.n557 Iout 0.03925
R16720 Iout.n554 Iout 0.03925
R16721 Iout.n434 Iout 0.03925
R16722 Iout.n438 Iout 0.03925
R16723 Iout.n441 Iout 0.03925
R16724 Iout.n432 Iout 0.03925
R16725 Iout.n418 Iout 0.03925
R16726 Iout.n416 Iout 0.03925
R16727 Iout.n402 Iout 0.03925
R16728 Iout.n357 Iout 0.03925
R16729 Iout.n360 Iout 0.03925
R16730 Iout.n363 Iout 0.03925
R16731 Iout.n366 Iout 0.03925
R16732 Iout.n354 Iout 0.03925
R16733 Iout.n351 Iout 0.03925
R16734 Iout.n348 Iout 0.03925
R16735 Iout.n345 Iout 0.03925
R16736 Iout.n342 Iout 0.03925
R16737 Iout.n339 Iout 0.03925
R16738 Iout.n336 Iout 0.03925
R16739 Iout.n333 Iout 0.03925
R16740 Iout.n117 Iout 0.03925
R16741 Iout.n582 Iout 0.03925
R16742 Iout.n111 Iout 0.03925
R16743 Iout.n594 Iout 0.03925
R16744 Iout.n105 Iout 0.03925
R16745 Iout.n606 Iout 0.03925
R16746 Iout.n99 Iout 0.03925
R16747 Iout.n618 Iout 0.03925
R16748 Iout.n624 Iout 0.03925
R16749 Iout.n90 Iout 0.03925
R16750 Iout.n636 Iout 0.03925
R16751 Iout.n81 Iout 0.03925
R16752 Iout.n648 Iout 0.03925
R16753 Iout.n96 Iout 0.03925
R16754 Iout.n612 Iout 0.03925
R16755 Iout.n102 Iout 0.03925
R16756 Iout.n600 Iout 0.03925
R16757 Iout.n108 Iout 0.03925
R16758 Iout.n588 Iout 0.03925
R16759 Iout.n687 Iout 0.03925
R16760 Iout.n684 Iout 0.03925
R16761 Iout.n681 Iout 0.03925
R16762 Iout.n678 Iout 0.03925
R16763 Iout.n675 Iout 0.03925
R16764 Iout.n672 Iout 0.03925
R16765 Iout.n747 Iout 0.03925
R16766 Iout.n50 Iout 0.03925
R16767 Iout.n759 Iout 0.03925
R16768 Iout.n44 Iout 0.03925
R16769 Iout.n771 Iout 0.03925
R16770 Iout.n42 Iout 0.03925
R16771 Iout.n56 Iout 0.03925
R16772 Iout.n735 Iout 0.03925
R16773 Iout.n62 Iout 0.03925
R16774 Iout.n723 Iout 0.03925
R16775 Iout.n717 Iout 0.03925
R16776 Iout.n65 Iout 0.03925
R16777 Iout.n729 Iout 0.03925
R16778 Iout.n59 Iout 0.03925
R16779 Iout.n805 Iout 0.03925
R16780 Iout.n808 Iout 0.03925
R16781 Iout.n811 Iout 0.03925
R16782 Iout.n814 Iout 0.03925
R16783 Iout.n817 Iout 0.03925
R16784 Iout.n820 Iout 0.03925
R16785 Iout.n823 Iout 0.03925
R16786 Iout.n802 Iout 0.03925
R16787 Iout.n799 Iout 0.03925
R16788 Iout.n890 Iout 0.03925
R16789 Iout.n888 Iout 0.03925
R16790 Iout.n881 Iout 0.03925
R16791 Iout.n869 Iout 0.03925
R16792 Iout.n867 Iout 0.03925
R16793 Iout.n855 Iout 0.03925
R16794 Iout.n853 Iout 0.03925
R16795 Iout.n841 Iout 0.03925
R16796 Iout.n839 Iout 0.03925
R16797 Iout.n827 Iout 0.03925
R16798 Iout.n883 Iout 0.03925
R16799 Iout.n895 Iout 0.03925
R16800 Iout.n897 Iout 0.03925
R16801 Iout.n909 Iout 0.03925
R16802 Iout.n911 Iout 0.03925
R16803 Iout.n923 Iout 0.03925
R16804 Iout.n926 Iout 0.03925
R16805 Iout.n22 Iout 0.03925
R16806 Iout.n876 Iout 0.03925
R16807 Iout.n874 Iout 0.03925
R16808 Iout.n862 Iout 0.03925
R16809 Iout.n860 Iout 0.03925
R16810 Iout.n848 Iout 0.03925
R16811 Iout.n846 Iout 0.03925
R16812 Iout.n834 Iout 0.03925
R16813 Iout.n832 Iout 0.03925
R16814 Iout.n902 Iout 0.03925
R16815 Iout.n904 Iout 0.03925
R16816 Iout.n916 Iout 0.03925
R16817 Iout.n918 Iout 0.03925
R16818 Iout.n931 Iout 0.03925
R16819 Iout.n934 Iout 0.03925
R16820 Iout.n796 Iout 0.03925
R16821 Iout.n793 Iout 0.03925
R16822 Iout.n790 Iout 0.03925
R16823 Iout.n787 Iout 0.03925
R16824 Iout.n784 Iout 0.03925
R16825 Iout.n781 Iout 0.03925
R16826 Iout.n938 Iout 0.03925
R16827 Iout.n741 Iout 0.03925
R16828 Iout.n53 Iout 0.03925
R16829 Iout.n753 Iout 0.03925
R16830 Iout.n47 Iout 0.03925
R16831 Iout.n765 Iout 0.03925
R16832 Iout.n38 Iout 0.03925
R16833 Iout.n777 Iout 0.03925
R16834 Iout.n71 Iout 0.03925
R16835 Iout.n705 Iout 0.03925
R16836 Iout.n77 Iout 0.03925
R16837 Iout.n944 Iout 0.03925
R16838 Iout.n19 Iout 0.03925
R16839 Iout.n68 Iout 0.03925
R16840 Iout.n711 Iout 0.03925
R16841 Iout.n74 Iout 0.03925
R16842 Iout.n699 Iout 0.03925
R16843 Iout.n950 Iout 0.03925
R16844 Iout.n953 Iout 0.03925
R16845 Iout.n669 Iout 0.03925
R16846 Iout.n666 Iout 0.03925
R16847 Iout.n663 Iout 0.03925
R16848 Iout.n660 Iout 0.03925
R16849 Iout.n657 Iout 0.03925
R16850 Iout.n654 Iout 0.03925
R16851 Iout.n690 Iout 0.03925
R16852 Iout.n695 Iout 0.03925
R16853 Iout.n692 Iout 0.03925
R16854 Iout.n957 Iout 0.03925
R16855 Iout.n114 Iout 0.03925
R16856 Iout.n576 Iout 0.03925
R16857 Iout.n573 Iout 0.03925
R16858 Iout.n963 Iout 0.03925
R16859 Iout.n14 Iout 0.03925
R16860 Iout.n93 Iout 0.03925
R16861 Iout.n630 Iout 0.03925
R16862 Iout.n87 Iout 0.03925
R16863 Iout.n642 Iout 0.03925
R16864 Iout.n85 Iout 0.03925
R16865 Iout.n563 Iout 0.03925
R16866 Iout.n969 Iout 0.03925
R16867 Iout.n972 Iout 0.03925
R16868 Iout.n569 Iout 0.03925
R16869 Iout.n123 Iout 0.03925
R16870 Iout.n120 Iout 0.03925
R16871 Iout.n976 Iout 0.03925
R16872 Iout.n400 Iout 0.03925
R16873 Iout.n386 Iout 0.03925
R16874 Iout.n384 Iout 0.03925
R16875 Iout.n370 Iout 0.03925
R16876 Iout.n982 Iout 0.03925
R16877 Iout.n9 Iout 0.03925
R16878 Iout.n127 Iout 0.03925
R16879 Iout.n988 Iout 0.03925
R16880 Iout.n991 Iout 0.03925
R16881 Iout.n323 Iout 0.03925
R16882 Iout.n326 Iout 0.03925
R16883 Iout.n329 Iout 0.03925
R16884 Iout.n995 Iout 0.03925
R16885 Iout.n1001 Iout 0.03925
R16886 Iout.n4 Iout 0.03925
R16887 Iout.n295 Iout 0.03925
R16888 Iout.n172 Iout 0.03925
R16889 Iout.n1014 Iout 0.03925
R16890 Iout.n1022 Iout 0.02071
R16891 Iout Iout.n1022 0.00379
R16892 Iout.n303 Iout.n302 0.00105952
R16893 Iout.n377 Iout.n375 0.00105952
R16894 Iout.n380 Iout.n379 0.00105952
R16895 Iout.n368 Iout.n367 0.00105952
R16896 Iout.n365 Iout.n364 0.00105952
R16897 Iout.n362 Iout.n361 0.00105952
R16898 Iout.n650 Iout.n649 0.00105952
R16899 Iout.n647 Iout.n82 0.00105952
R16900 Iout.n638 Iout.n637 0.00105952
R16901 Iout.n635 Iout.n91 0.00105952
R16902 Iout.n43 Iout.n41 0.00105952
R16903 Iout.n773 Iout.n772 0.00105952
R16904 Iout.n770 Iout.n45 0.00105952
R16905 Iout.n761 Iout.n760 0.00105952
R16906 Iout.n758 Iout.n51 0.00105952
R16907 Iout.n825 Iout.n824 0.00105952
R16908 Iout.n822 Iout.n821 0.00105952
R16909 Iout.n819 Iout.n818 0.00105952
R16910 Iout.n816 Iout.n815 0.00105952
R16911 Iout.n813 Iout.n812 0.00105952
R16912 Iout.n810 Iout.n809 0.00105952
R16913 Iout.n829 Iout.n828 0.00105952
R16914 Iout.n840 Iout.n838 0.00105952
R16915 Iout.n843 Iout.n842 0.00105952
R16916 Iout.n854 Iout.n852 0.00105952
R16917 Iout.n857 Iout.n856 0.00105952
R16918 Iout.n868 Iout.n866 0.00105952
R16919 Iout.n871 Iout.n870 0.00105952
R16920 Iout.n925 Iout.n23 0.00105952
R16921 Iout.n928 Iout.n927 0.00105952
R16922 Iout.n924 Iout.n922 0.00105952
R16923 Iout.n913 Iout.n912 0.00105952
R16924 Iout.n910 Iout.n908 0.00105952
R16925 Iout.n899 Iout.n898 0.00105952
R16926 Iout.n896 Iout.n894 0.00105952
R16927 Iout.n885 Iout.n884 0.00105952
R16928 Iout.n882 Iout.n880 0.00105952
R16929 Iout.n833 Iout.n831 0.00105952
R16930 Iout.n836 Iout.n835 0.00105952
R16931 Iout.n847 Iout.n845 0.00105952
R16932 Iout.n850 Iout.n849 0.00105952
R16933 Iout.n861 Iout.n859 0.00105952
R16934 Iout.n864 Iout.n863 0.00105952
R16935 Iout.n875 Iout.n873 0.00105952
R16936 Iout.n878 Iout.n877 0.00105952
R16937 Iout.n889 Iout.n887 0.00105952
R16938 Iout.n935 Iout.n933 0.00105952
R16939 Iout.n932 Iout.n930 0.00105952
R16940 Iout.n920 Iout.n919 0.00105952
R16941 Iout.n917 Iout.n915 0.00105952
R16942 Iout.n906 Iout.n905 0.00105952
R16943 Iout.n903 Iout.n901 0.00105952
R16944 Iout.n892 Iout.n891 0.00105952
R16945 Iout.n940 Iout.n939 0.00105952
R16946 Iout.n783 Iout.n782 0.00105952
R16947 Iout.n786 Iout.n785 0.00105952
R16948 Iout.n789 Iout.n788 0.00105952
R16949 Iout.n792 Iout.n791 0.00105952
R16950 Iout.n795 Iout.n794 0.00105952
R16951 Iout.n798 Iout.n797 0.00105952
R16952 Iout.n801 Iout.n800 0.00105952
R16953 Iout.n804 Iout.n803 0.00105952
R16954 Iout.n807 Iout.n806 0.00105952
R16955 Iout.n779 Iout.n778 0.00105952
R16956 Iout.n776 Iout.n39 0.00105952
R16957 Iout.n767 Iout.n766 0.00105952
R16958 Iout.n764 Iout.n48 0.00105952
R16959 Iout.n755 Iout.n754 0.00105952
R16960 Iout.n752 Iout.n54 0.00105952
R16961 Iout.n743 Iout.n742 0.00105952
R16962 Iout.n740 Iout.n60 0.00105952
R16963 Iout.n731 Iout.n730 0.00105952
R16964 Iout.n728 Iout.n66 0.00105952
R16965 Iout.n943 Iout.n20 0.00105952
R16966 Iout.n946 Iout.n945 0.00105952
R16967 Iout.n704 Iout.n78 0.00105952
R16968 Iout.n707 Iout.n706 0.00105952
R16969 Iout.n716 Iout.n72 0.00105952
R16970 Iout.n719 Iout.n718 0.00105952
R16971 Iout.n954 Iout.n952 0.00105952
R16972 Iout.n951 Iout.n949 0.00105952
R16973 Iout.n701 Iout.n700 0.00105952
R16974 Iout.n710 Iout.n75 0.00105952
R16975 Iout.n713 Iout.n712 0.00105952
R16976 Iout.n722 Iout.n69 0.00105952
R16977 Iout.n725 Iout.n724 0.00105952
R16978 Iout.n734 Iout.n63 0.00105952
R16979 Iout.n737 Iout.n736 0.00105952
R16980 Iout.n746 Iout.n57 0.00105952
R16981 Iout.n749 Iout.n748 0.00105952
R16982 Iout.n655 Iout.n653 0.00105952
R16983 Iout.n658 Iout.n656 0.00105952
R16984 Iout.n661 Iout.n659 0.00105952
R16985 Iout.n664 Iout.n662 0.00105952
R16986 Iout.n667 Iout.n665 0.00105952
R16987 Iout.n670 Iout.n668 0.00105952
R16988 Iout.n673 Iout.n671 0.00105952
R16989 Iout.n676 Iout.n674 0.00105952
R16990 Iout.n679 Iout.n677 0.00105952
R16991 Iout.n682 Iout.n680 0.00105952
R16992 Iout.n685 Iout.n683 0.00105952
R16993 Iout.n959 Iout.n958 0.00105952
R16994 Iout.n694 Iout.n693 0.00105952
R16995 Iout.n697 Iout.n696 0.00105952
R16996 Iout.n691 Iout.n689 0.00105952
R16997 Iout.n688 Iout.n686 0.00105952
R16998 Iout.n962 Iout.n15 0.00105952
R16999 Iout.n965 Iout.n964 0.00105952
R17000 Iout.n575 Iout.n574 0.00105952
R17001 Iout.n578 Iout.n577 0.00105952
R17002 Iout.n587 Iout.n115 0.00105952
R17003 Iout.n590 Iout.n589 0.00105952
R17004 Iout.n599 Iout.n109 0.00105952
R17005 Iout.n602 Iout.n601 0.00105952
R17006 Iout.n611 Iout.n103 0.00105952
R17007 Iout.n614 Iout.n613 0.00105952
R17008 Iout.n623 Iout.n97 0.00105952
R17009 Iout.n626 Iout.n625 0.00105952
R17010 Iout.n86 Iout.n84 0.00105952
R17011 Iout.n644 Iout.n643 0.00105952
R17012 Iout.n641 Iout.n88 0.00105952
R17013 Iout.n632 Iout.n631 0.00105952
R17014 Iout.n629 Iout.n94 0.00105952
R17015 Iout.n620 Iout.n619 0.00105952
R17016 Iout.n617 Iout.n100 0.00105952
R17017 Iout.n608 Iout.n607 0.00105952
R17018 Iout.n605 Iout.n106 0.00105952
R17019 Iout.n596 Iout.n595 0.00105952
R17020 Iout.n593 Iout.n112 0.00105952
R17021 Iout.n584 Iout.n583 0.00105952
R17022 Iout.n973 Iout.n971 0.00105952
R17023 Iout.n970 Iout.n968 0.00105952
R17024 Iout.n565 Iout.n564 0.00105952
R17025 Iout.n581 Iout.n118 0.00105952
R17026 Iout.n978 Iout.n977 0.00105952
R17027 Iout.n122 Iout.n121 0.00105952
R17028 Iout.n568 Iout.n124 0.00105952
R17029 Iout.n571 Iout.n570 0.00105952
R17030 Iout.n335 Iout.n334 0.00105952
R17031 Iout.n338 Iout.n337 0.00105952
R17032 Iout.n341 Iout.n340 0.00105952
R17033 Iout.n344 Iout.n343 0.00105952
R17034 Iout.n347 Iout.n346 0.00105952
R17035 Iout.n350 Iout.n349 0.00105952
R17036 Iout.n353 Iout.n352 0.00105952
R17037 Iout.n356 Iout.n355 0.00105952
R17038 Iout.n359 Iout.n358 0.00105952
R17039 Iout.n372 Iout.n371 0.00105952
R17040 Iout.n385 Iout.n383 0.00105952
R17041 Iout.n388 Iout.n387 0.00105952
R17042 Iout.n401 Iout.n399 0.00105952
R17043 Iout.n404 Iout.n403 0.00105952
R17044 Iout.n417 Iout.n415 0.00105952
R17045 Iout.n420 Iout.n419 0.00105952
R17046 Iout.n433 Iout.n431 0.00105952
R17047 Iout.n443 Iout.n442 0.00105952
R17048 Iout.n440 Iout.n439 0.00105952
R17049 Iout.n437 Iout.n435 0.00105952
R17050 Iout.n555 Iout.n553 0.00105952
R17051 Iout.n558 Iout.n556 0.00105952
R17052 Iout.n981 Iout.n10 0.00105952
R17053 Iout.n984 Iout.n983 0.00105952
R17054 Iout.n561 Iout.n560 0.00105952
R17055 Iout.n992 Iout.n990 0.00105952
R17056 Iout.n989 Iout.n987 0.00105952
R17057 Iout.n129 Iout.n128 0.00105952
R17058 Iout.n547 Iout.n131 0.00105952
R17059 Iout.n550 Iout.n549 0.00105952
R17060 Iout.n451 Iout.n450 0.00105952
R17061 Iout.n454 Iout.n453 0.00105952
R17062 Iout.n448 Iout.n446 0.00105952
R17063 Iout.n428 Iout.n427 0.00105952
R17064 Iout.n425 Iout.n423 0.00105952
R17065 Iout.n412 Iout.n411 0.00105952
R17066 Iout.n409 Iout.n407 0.00105952
R17067 Iout.n396 Iout.n395 0.00105952
R17068 Iout.n393 Iout.n391 0.00105952
R17069 Iout.n331 Iout.n330 0.00105952
R17070 Iout.n328 Iout.n327 0.00105952
R17071 Iout.n325 Iout.n324 0.00105952
R17072 Iout.n322 Iout.n321 0.00105952
R17073 Iout.n319 Iout.n318 0.00105952
R17074 Iout.n316 Iout.n315 0.00105952
R17075 Iout.n313 Iout.n312 0.00105952
R17076 Iout.n310 Iout.n309 0.00105952
R17077 Iout.n307 Iout.n306 0.00105952
R17078 Iout.n459 Iout.n457 0.00105952
R17079 Iout.n465 Iout.n464 0.00105952
R17080 Iout.n462 Iout.n461 0.00105952
R17081 Iout.n544 Iout.n543 0.00105952
R17082 Iout.n541 Iout.n137 0.00105952
R17083 Iout.n997 Iout.n996 0.00105952
R17084 Iout.n135 Iout.n134 0.00105952
R17085 Iout.n1000 Iout.n5 0.00105952
R17086 Iout.n1003 Iout.n1002 0.00105952
R17087 Iout.n538 Iout.n537 0.00105952
R17088 Iout.n535 Iout.n533 0.00105952
R17089 Iout.n532 Iout.n530 0.00105952
R17090 Iout.n468 Iout.n157 0.00105952
R17091 Iout.n471 Iout.n470 0.00105952
R17092 Iout.n474 Iout.n473 0.00105952
R17093 Iout.n264 Iout.n190 0.00105952
R17094 Iout.n267 Iout.n266 0.00105952
R17095 Iout.n276 Iout.n184 0.00105952
R17096 Iout.n279 Iout.n278 0.00105952
R17097 Iout.n288 Iout.n178 0.00105952
R17098 Iout.n291 Iout.n290 0.00105952
R17099 Iout.n300 Iout.n169 0.00105952
R17100 Iout.n173 Iout.n171 0.00105952
R17101 Iout.n297 Iout.n296 0.00105952
R17102 Iout.n294 Iout.n175 0.00105952
R17103 Iout.n285 Iout.n284 0.00105952
R17104 Iout.n282 Iout.n181 0.00105952
R17105 Iout.n273 Iout.n272 0.00105952
R17106 Iout.n270 Iout.n187 0.00105952
R17107 Iout.n261 Iout.n260 0.00105952
R17108 Iout.n479 Iout.n477 0.00105952
R17109 Iout.n485 Iout.n484 0.00105952
R17110 Iout.n482 Iout.n481 0.00105952
R17111 Iout.n527 Iout.n526 0.00105952
R17112 Iout.n524 Iout.n144 0.00105952
R17113 Iout.n142 Iout.n141 0.00105952
R17114 Iout.n1008 Iout.n1006 0.00105952
R17115 Iout.n1011 Iout.n1009 0.00105952
R17116 Iout.n1016 Iout.n1015 0.00105952
R17117 Iout.n148 Iout.n147 0.00105952
R17118 Iout.n518 Iout.n150 0.00105952
R17119 Iout.n521 Iout.n520 0.00105952
R17120 Iout.n493 Iout.n492 0.00105952
R17121 Iout.n496 Iout.n495 0.00105952
R17122 Iout.n490 Iout.n488 0.00105952
R17123 Iout.n254 Iout.n253 0.00105952
R17124 Iout.n257 Iout.n256 0.00105952
R17125 Iout.n251 Iout.n249 0.00105952
R17126 Iout.n248 Iout.n246 0.00105952
R17127 Iout.n245 Iout.n243 0.00105952
R17128 Iout.n242 Iout.n240 0.00105952
R17129 Iout.n239 Iout.n237 0.00105952
R17130 Iout.n236 Iout.n234 0.00105952
R17131 Iout.n233 Iout.n231 0.00105952
R17132 Iout.n228 Iout.n227 0.00105952
R17133 Iout.n225 Iout.n223 0.00105952
R17134 Iout.n221 Iout.n219 0.00105952
R17135 Iout.n217 Iout.n215 0.00105952
R17136 Iout.n213 Iout.n211 0.00105952
R17137 Iout.n209 Iout.n207 0.00105952
R17138 Iout.n205 Iout.n203 0.00105952
R17139 Iout.n201 Iout.n200 0.00105952
R17140 Iout.n198 Iout.n196 0.00105952
R17141 Iout.n194 Iout.n193 0.00105952
R17142 Iout.n501 Iout.n499 0.00105952
R17143 Iout.n505 Iout.n503 0.00105952
R17144 Iout.n508 Iout.n506 0.00105952
R17145 Iout.n515 Iout.n514 0.00105952
R17146 Iout.n512 Iout.n510 0.00105952
R17147 Iout.n1021 Iout.n1019 0.00105952
R17148 XThC.Tn[10].n55 XThC.Tn[10].n54 256.103
R17149 XThC.Tn[10].n59 XThC.Tn[10].n57 243.68
R17150 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R17151 XThC.Tn[10].n59 XThC.Tn[10].n58 205.28
R17152 XThC.Tn[10].n55 XThC.Tn[10].n53 202.095
R17153 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R17154 XThC.Tn[10].n5 XThC.Tn[10].n3 161.406
R17155 XThC.Tn[10].n8 XThC.Tn[10].n6 161.406
R17156 XThC.Tn[10].n11 XThC.Tn[10].n9 161.406
R17157 XThC.Tn[10].n14 XThC.Tn[10].n12 161.406
R17158 XThC.Tn[10].n17 XThC.Tn[10].n15 161.406
R17159 XThC.Tn[10].n20 XThC.Tn[10].n18 161.406
R17160 XThC.Tn[10].n23 XThC.Tn[10].n21 161.406
R17161 XThC.Tn[10].n26 XThC.Tn[10].n24 161.406
R17162 XThC.Tn[10].n29 XThC.Tn[10].n27 161.406
R17163 XThC.Tn[10].n32 XThC.Tn[10].n30 161.406
R17164 XThC.Tn[10].n35 XThC.Tn[10].n33 161.406
R17165 XThC.Tn[10].n38 XThC.Tn[10].n36 161.406
R17166 XThC.Tn[10].n41 XThC.Tn[10].n39 161.406
R17167 XThC.Tn[10].n44 XThC.Tn[10].n42 161.406
R17168 XThC.Tn[10].n47 XThC.Tn[10].n45 161.406
R17169 XThC.Tn[10].n50 XThC.Tn[10].n48 161.406
R17170 XThC.Tn[10].n3 XThC.Tn[10].t36 161.202
R17171 XThC.Tn[10].n6 XThC.Tn[10].t21 161.202
R17172 XThC.Tn[10].n9 XThC.Tn[10].t23 161.202
R17173 XThC.Tn[10].n12 XThC.Tn[10].t25 161.202
R17174 XThC.Tn[10].n15 XThC.Tn[10].t14 161.202
R17175 XThC.Tn[10].n18 XThC.Tn[10].t15 161.202
R17176 XThC.Tn[10].n21 XThC.Tn[10].t28 161.202
R17177 XThC.Tn[10].n24 XThC.Tn[10].t37 161.202
R17178 XThC.Tn[10].n27 XThC.Tn[10].t39 161.202
R17179 XThC.Tn[10].n30 XThC.Tn[10].t26 161.202
R17180 XThC.Tn[10].n33 XThC.Tn[10].t27 161.202
R17181 XThC.Tn[10].n36 XThC.Tn[10].t40 161.202
R17182 XThC.Tn[10].n39 XThC.Tn[10].t16 161.202
R17183 XThC.Tn[10].n42 XThC.Tn[10].t19 161.202
R17184 XThC.Tn[10].n45 XThC.Tn[10].t32 161.202
R17185 XThC.Tn[10].n48 XThC.Tn[10].t42 161.202
R17186 XThC.Tn[10].n3 XThC.Tn[10].t38 145.137
R17187 XThC.Tn[10].n6 XThC.Tn[10].t24 145.137
R17188 XThC.Tn[10].n9 XThC.Tn[10].t29 145.137
R17189 XThC.Tn[10].n12 XThC.Tn[10].t30 145.137
R17190 XThC.Tn[10].n15 XThC.Tn[10].t17 145.137
R17191 XThC.Tn[10].n18 XThC.Tn[10].t18 145.137
R17192 XThC.Tn[10].n21 XThC.Tn[10].t34 145.137
R17193 XThC.Tn[10].n24 XThC.Tn[10].t41 145.137
R17194 XThC.Tn[10].n27 XThC.Tn[10].t43 145.137
R17195 XThC.Tn[10].n30 XThC.Tn[10].t31 145.137
R17196 XThC.Tn[10].n33 XThC.Tn[10].t33 145.137
R17197 XThC.Tn[10].n36 XThC.Tn[10].t12 145.137
R17198 XThC.Tn[10].n39 XThC.Tn[10].t20 145.137
R17199 XThC.Tn[10].n42 XThC.Tn[10].t22 145.137
R17200 XThC.Tn[10].n45 XThC.Tn[10].t35 145.137
R17201 XThC.Tn[10].n48 XThC.Tn[10].t13 145.137
R17202 XThC.Tn[10].n53 XThC.Tn[10].t5 26.5955
R17203 XThC.Tn[10].n53 XThC.Tn[10].t4 26.5955
R17204 XThC.Tn[10].n57 XThC.Tn[10].t1 26.5955
R17205 XThC.Tn[10].n57 XThC.Tn[10].t8 26.5955
R17206 XThC.Tn[10].n58 XThC.Tn[10].t11 26.5955
R17207 XThC.Tn[10].n58 XThC.Tn[10].t9 26.5955
R17208 XThC.Tn[10].n54 XThC.Tn[10].t7 26.5955
R17209 XThC.Tn[10].n54 XThC.Tn[10].t0 26.5955
R17210 XThC.Tn[10].n1 XThC.Tn[10].t10 24.9236
R17211 XThC.Tn[10].n1 XThC.Tn[10].t3 24.9236
R17212 XThC.Tn[10].n0 XThC.Tn[10].t2 24.9236
R17213 XThC.Tn[10].n0 XThC.Tn[10].t6 24.9236
R17214 XThC.Tn[10] XThC.Tn[10].n59 22.9652
R17215 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R17216 XThC.Tn[10].n56 XThC.Tn[10].n55 13.9299
R17217 XThC.Tn[10] XThC.Tn[10].n56 13.9299
R17218 XThC.Tn[10].n52 XThC.Tn[10].n51 5.13256
R17219 XThC.Tn[10].n56 XThC.Tn[10].n52 2.99115
R17220 XThC.Tn[10].n56 XThC.Tn[10] 2.87153
R17221 XThC.Tn[10].n52 XThC.Tn[10] 2.2734
R17222 XThC.Tn[10].n51 XThC.Tn[10] 2.26343
R17223 XThC.Tn[10].n8 XThC.Tn[10] 0.931056
R17224 XThC.Tn[10].n11 XThC.Tn[10] 0.931056
R17225 XThC.Tn[10].n14 XThC.Tn[10] 0.931056
R17226 XThC.Tn[10].n17 XThC.Tn[10] 0.931056
R17227 XThC.Tn[10].n20 XThC.Tn[10] 0.931056
R17228 XThC.Tn[10].n23 XThC.Tn[10] 0.931056
R17229 XThC.Tn[10].n26 XThC.Tn[10] 0.931056
R17230 XThC.Tn[10].n29 XThC.Tn[10] 0.931056
R17231 XThC.Tn[10].n32 XThC.Tn[10] 0.931056
R17232 XThC.Tn[10].n35 XThC.Tn[10] 0.931056
R17233 XThC.Tn[10].n38 XThC.Tn[10] 0.931056
R17234 XThC.Tn[10].n41 XThC.Tn[10] 0.931056
R17235 XThC.Tn[10].n44 XThC.Tn[10] 0.931056
R17236 XThC.Tn[10].n47 XThC.Tn[10] 0.931056
R17237 XThC.Tn[10].n50 XThC.Tn[10] 0.931056
R17238 XThC.Tn[10] XThC.Tn[10].n5 0.396333
R17239 XThC.Tn[10] XThC.Tn[10].n8 0.396333
R17240 XThC.Tn[10] XThC.Tn[10].n11 0.396333
R17241 XThC.Tn[10] XThC.Tn[10].n14 0.396333
R17242 XThC.Tn[10] XThC.Tn[10].n17 0.396333
R17243 XThC.Tn[10] XThC.Tn[10].n20 0.396333
R17244 XThC.Tn[10] XThC.Tn[10].n23 0.396333
R17245 XThC.Tn[10] XThC.Tn[10].n26 0.396333
R17246 XThC.Tn[10] XThC.Tn[10].n29 0.396333
R17247 XThC.Tn[10] XThC.Tn[10].n32 0.396333
R17248 XThC.Tn[10] XThC.Tn[10].n35 0.396333
R17249 XThC.Tn[10] XThC.Tn[10].n38 0.396333
R17250 XThC.Tn[10] XThC.Tn[10].n41 0.396333
R17251 XThC.Tn[10] XThC.Tn[10].n44 0.396333
R17252 XThC.Tn[10] XThC.Tn[10].n47 0.396333
R17253 XThC.Tn[10] XThC.Tn[10].n50 0.396333
R17254 XThC.Tn[10].n4 XThC.Tn[10] 0.104667
R17255 XThC.Tn[10].n7 XThC.Tn[10] 0.104667
R17256 XThC.Tn[10].n10 XThC.Tn[10] 0.104667
R17257 XThC.Tn[10].n13 XThC.Tn[10] 0.104667
R17258 XThC.Tn[10].n16 XThC.Tn[10] 0.104667
R17259 XThC.Tn[10].n19 XThC.Tn[10] 0.104667
R17260 XThC.Tn[10].n22 XThC.Tn[10] 0.104667
R17261 XThC.Tn[10].n25 XThC.Tn[10] 0.104667
R17262 XThC.Tn[10].n28 XThC.Tn[10] 0.104667
R17263 XThC.Tn[10].n31 XThC.Tn[10] 0.104667
R17264 XThC.Tn[10].n34 XThC.Tn[10] 0.104667
R17265 XThC.Tn[10].n37 XThC.Tn[10] 0.104667
R17266 XThC.Tn[10].n40 XThC.Tn[10] 0.104667
R17267 XThC.Tn[10].n43 XThC.Tn[10] 0.104667
R17268 XThC.Tn[10].n46 XThC.Tn[10] 0.104667
R17269 XThC.Tn[10].n49 XThC.Tn[10] 0.104667
R17270 XThC.Tn[10].n4 XThC.Tn[10] 0.0309878
R17271 XThC.Tn[10].n7 XThC.Tn[10] 0.0309878
R17272 XThC.Tn[10].n10 XThC.Tn[10] 0.0309878
R17273 XThC.Tn[10].n13 XThC.Tn[10] 0.0309878
R17274 XThC.Tn[10].n16 XThC.Tn[10] 0.0309878
R17275 XThC.Tn[10].n19 XThC.Tn[10] 0.0309878
R17276 XThC.Tn[10].n22 XThC.Tn[10] 0.0309878
R17277 XThC.Tn[10].n25 XThC.Tn[10] 0.0309878
R17278 XThC.Tn[10].n28 XThC.Tn[10] 0.0309878
R17279 XThC.Tn[10].n31 XThC.Tn[10] 0.0309878
R17280 XThC.Tn[10].n34 XThC.Tn[10] 0.0309878
R17281 XThC.Tn[10].n37 XThC.Tn[10] 0.0309878
R17282 XThC.Tn[10].n40 XThC.Tn[10] 0.0309878
R17283 XThC.Tn[10].n43 XThC.Tn[10] 0.0309878
R17284 XThC.Tn[10].n46 XThC.Tn[10] 0.0309878
R17285 XThC.Tn[10].n49 XThC.Tn[10] 0.0309878
R17286 XThC.Tn[10].n5 XThC.Tn[10].n4 0.027939
R17287 XThC.Tn[10].n8 XThC.Tn[10].n7 0.027939
R17288 XThC.Tn[10].n11 XThC.Tn[10].n10 0.027939
R17289 XThC.Tn[10].n14 XThC.Tn[10].n13 0.027939
R17290 XThC.Tn[10].n17 XThC.Tn[10].n16 0.027939
R17291 XThC.Tn[10].n20 XThC.Tn[10].n19 0.027939
R17292 XThC.Tn[10].n23 XThC.Tn[10].n22 0.027939
R17293 XThC.Tn[10].n26 XThC.Tn[10].n25 0.027939
R17294 XThC.Tn[10].n29 XThC.Tn[10].n28 0.027939
R17295 XThC.Tn[10].n32 XThC.Tn[10].n31 0.027939
R17296 XThC.Tn[10].n35 XThC.Tn[10].n34 0.027939
R17297 XThC.Tn[10].n38 XThC.Tn[10].n37 0.027939
R17298 XThC.Tn[10].n41 XThC.Tn[10].n40 0.027939
R17299 XThC.Tn[10].n44 XThC.Tn[10].n43 0.027939
R17300 XThC.Tn[10].n47 XThC.Tn[10].n46 0.027939
R17301 XThC.Tn[10].n50 XThC.Tn[10].n49 0.027939
R17302 XThC.Tn[10].n51 XThC.Tn[10] 0.00285068
R17303 XThR.XTBN.Y.n1 XThR.XTBN.Y.t60 212.081
R17304 XThR.XTBN.Y.n8 XThR.XTBN.Y.t12 212.081
R17305 XThR.XTBN.Y.n2 XThR.XTBN.Y.t81 212.081
R17306 XThR.XTBN.Y.n3 XThR.XTBN.Y.t121 212.081
R17307 XThR.XTBN.Y.n12 XThR.XTBN.Y.t115 212.081
R17308 XThR.XTBN.Y.n19 XThR.XTBN.Y.t65 212.081
R17309 XThR.XTBN.Y.n13 XThR.XTBN.Y.t21 212.081
R17310 XThR.XTBN.Y.n14 XThR.XTBN.Y.t57 212.081
R17311 XThR.XTBN.Y.n24 XThR.XTBN.Y.t27 212.081
R17312 XThR.XTBN.Y.n31 XThR.XTBN.Y.t96 212.081
R17313 XThR.XTBN.Y.n25 XThR.XTBN.Y.t46 212.081
R17314 XThR.XTBN.Y.n26 XThR.XTBN.Y.t89 212.081
R17315 XThR.XTBN.Y.n36 XThR.XTBN.Y.t80 212.081
R17316 XThR.XTBN.Y.n43 XThR.XTBN.Y.t31 212.081
R17317 XThR.XTBN.Y.n37 XThR.XTBN.Y.t102 212.081
R17318 XThR.XTBN.Y.n38 XThR.XTBN.Y.t25 212.081
R17319 XThR.XTBN.Y.n48 XThR.XTBN.Y.t85 212.081
R17320 XThR.XTBN.Y.n55 XThR.XTBN.Y.t33 212.081
R17321 XThR.XTBN.Y.n49 XThR.XTBN.Y.t105 212.081
R17322 XThR.XTBN.Y.n50 XThR.XTBN.Y.t26 212.081
R17323 XThR.XTBN.Y.n60 XThR.XTBN.Y.t54 212.081
R17324 XThR.XTBN.Y.n67 XThR.XTBN.Y.t5 212.081
R17325 XThR.XTBN.Y.n61 XThR.XTBN.Y.t73 212.081
R17326 XThR.XTBN.Y.n62 XThR.XTBN.Y.t114 212.081
R17327 XThR.XTBN.Y.n72 XThR.XTBN.Y.t49 212.081
R17328 XThR.XTBN.Y.n79 XThR.XTBN.Y.t119 212.081
R17329 XThR.XTBN.Y.n73 XThR.XTBN.Y.t69 212.081
R17330 XThR.XTBN.Y.n74 XThR.XTBN.Y.t108 212.081
R17331 XThR.XTBN.Y.n163 XThR.XTBN.Y.t41 212.081
R17332 XThR.XTBN.Y.n154 XThR.XTBN.Y.t113 212.081
R17333 XThR.XTBN.Y.n158 XThR.XTBN.Y.t34 212.081
R17334 XThR.XTBN.Y.n155 XThR.XTBN.Y.t72 212.081
R17335 XThR.XTBN.Y.n151 XThR.XTBN.Y.t19 212.081
R17336 XThR.XTBN.Y.n142 XThR.XTBN.Y.t86 212.081
R17337 XThR.XTBN.Y.n146 XThR.XTBN.Y.t6 212.081
R17338 XThR.XTBN.Y.n143 XThR.XTBN.Y.t43 212.081
R17339 XThR.XTBN.Y.n139 XThR.XTBN.Y.t45 212.081
R17340 XThR.XTBN.Y.n130 XThR.XTBN.Y.t117 212.081
R17341 XThR.XTBN.Y.n134 XThR.XTBN.Y.t36 212.081
R17342 XThR.XTBN.Y.n131 XThR.XTBN.Y.t75 212.081
R17343 XThR.XTBN.Y.n127 XThR.XTBN.Y.t100 212.081
R17344 XThR.XTBN.Y.n118 XThR.XTBN.Y.t50 212.081
R17345 XThR.XTBN.Y.n122 XThR.XTBN.Y.t92 212.081
R17346 XThR.XTBN.Y.n119 XThR.XTBN.Y.t13 212.081
R17347 XThR.XTBN.Y.n115 XThR.XTBN.Y.t15 212.081
R17348 XThR.XTBN.Y.n106 XThR.XTBN.Y.t83 212.081
R17349 XThR.XTBN.Y.n110 XThR.XTBN.Y.t123 212.081
R17350 XThR.XTBN.Y.n107 XThR.XTBN.Y.t39 212.081
R17351 XThR.XTBN.Y.n103 XThR.XTBN.Y.t66 212.081
R17352 XThR.XTBN.Y.n94 XThR.XTBN.Y.t23 212.081
R17353 XThR.XTBN.Y.n98 XThR.XTBN.Y.t59 212.081
R17354 XThR.XTBN.Y.n95 XThR.XTBN.Y.t97 212.081
R17355 XThR.XTBN.Y.n92 XThR.XTBN.Y.t99 212.081
R17356 XThR.XTBN.Y.n83 XThR.XTBN.Y.t87 212.081
R17357 XThR.XTBN.Y.n87 XThR.XTBN.Y.t77 212.081
R17358 XThR.XTBN.Y.n84 XThR.XTBN.Y.t68 212.081
R17359 XThR.XTBN.Y.n167 XThR.XTBN.Y.t63 212.081
R17360 XThR.XTBN.Y.n169 XThR.XTBN.Y.t106 212.081
R17361 XThR.XTBN.Y.n174 XThR.XTBN.Y.t56 212.081
R17362 XThR.XTBN.Y.n170 XThR.XTBN.Y.t7 212.081
R17363 XThR.XTBN.Y XThR.XTBN.Y.n180 203.923
R17364 XThR.XTBN.Y.n171 XThR.XTBN.Y.n170 188.516
R17365 XThR.XTBN.Y.n164 XThR.XTBN.Y.n163 180.482
R17366 XThR.XTBN.Y.n152 XThR.XTBN.Y.n151 180.482
R17367 XThR.XTBN.Y.n140 XThR.XTBN.Y.n139 180.482
R17368 XThR.XTBN.Y.n128 XThR.XTBN.Y.n127 180.482
R17369 XThR.XTBN.Y.n116 XThR.XTBN.Y.n115 180.482
R17370 XThR.XTBN.Y.n104 XThR.XTBN.Y.n103 180.482
R17371 XThR.XTBN.Y.n93 XThR.XTBN.Y.n92 180.482
R17372 XThR.XTBN.Y.n5 XThR.XTBN.Y.n4 173.761
R17373 XThR.XTBN.Y.n16 XThR.XTBN.Y.n15 173.761
R17374 XThR.XTBN.Y.n28 XThR.XTBN.Y.n27 173.761
R17375 XThR.XTBN.Y.n40 XThR.XTBN.Y.n39 173.761
R17376 XThR.XTBN.Y.n52 XThR.XTBN.Y.n51 173.761
R17377 XThR.XTBN.Y.n64 XThR.XTBN.Y.n63 173.761
R17378 XThR.XTBN.Y.n76 XThR.XTBN.Y.n75 173.761
R17379 XThR.XTBN.Y.n168 XThR.XTBN.Y 154.304
R17380 XThR.XTBN.Y.n10 XThR.XTBN.Y.n9 152
R17381 XThR.XTBN.Y.n7 XThR.XTBN.Y.n0 152
R17382 XThR.XTBN.Y.n6 XThR.XTBN.Y.n5 152
R17383 XThR.XTBN.Y.n17 XThR.XTBN.Y.n16 152
R17384 XThR.XTBN.Y.n18 XThR.XTBN.Y.n11 152
R17385 XThR.XTBN.Y.n21 XThR.XTBN.Y.n20 152
R17386 XThR.XTBN.Y.n29 XThR.XTBN.Y.n28 152
R17387 XThR.XTBN.Y.n30 XThR.XTBN.Y.n23 152
R17388 XThR.XTBN.Y.n33 XThR.XTBN.Y.n32 152
R17389 XThR.XTBN.Y.n41 XThR.XTBN.Y.n40 152
R17390 XThR.XTBN.Y.n42 XThR.XTBN.Y.n35 152
R17391 XThR.XTBN.Y.n45 XThR.XTBN.Y.n44 152
R17392 XThR.XTBN.Y.n53 XThR.XTBN.Y.n52 152
R17393 XThR.XTBN.Y.n54 XThR.XTBN.Y.n47 152
R17394 XThR.XTBN.Y.n57 XThR.XTBN.Y.n56 152
R17395 XThR.XTBN.Y.n65 XThR.XTBN.Y.n64 152
R17396 XThR.XTBN.Y.n66 XThR.XTBN.Y.n59 152
R17397 XThR.XTBN.Y.n69 XThR.XTBN.Y.n68 152
R17398 XThR.XTBN.Y.n77 XThR.XTBN.Y.n76 152
R17399 XThR.XTBN.Y.n78 XThR.XTBN.Y.n71 152
R17400 XThR.XTBN.Y.n81 XThR.XTBN.Y.n80 152
R17401 XThR.XTBN.Y.n157 XThR.XTBN.Y.n156 152
R17402 XThR.XTBN.Y.n160 XThR.XTBN.Y.n159 152
R17403 XThR.XTBN.Y.n162 XThR.XTBN.Y.n161 152
R17404 XThR.XTBN.Y.n145 XThR.XTBN.Y.n144 152
R17405 XThR.XTBN.Y.n148 XThR.XTBN.Y.n147 152
R17406 XThR.XTBN.Y.n150 XThR.XTBN.Y.n149 152
R17407 XThR.XTBN.Y.n133 XThR.XTBN.Y.n132 152
R17408 XThR.XTBN.Y.n136 XThR.XTBN.Y.n135 152
R17409 XThR.XTBN.Y.n138 XThR.XTBN.Y.n137 152
R17410 XThR.XTBN.Y.n121 XThR.XTBN.Y.n120 152
R17411 XThR.XTBN.Y.n124 XThR.XTBN.Y.n123 152
R17412 XThR.XTBN.Y.n126 XThR.XTBN.Y.n125 152
R17413 XThR.XTBN.Y.n109 XThR.XTBN.Y.n108 152
R17414 XThR.XTBN.Y.n112 XThR.XTBN.Y.n111 152
R17415 XThR.XTBN.Y.n114 XThR.XTBN.Y.n113 152
R17416 XThR.XTBN.Y.n97 XThR.XTBN.Y.n96 152
R17417 XThR.XTBN.Y.n100 XThR.XTBN.Y.n99 152
R17418 XThR.XTBN.Y.n102 XThR.XTBN.Y.n101 152
R17419 XThR.XTBN.Y.n86 XThR.XTBN.Y.n85 152
R17420 XThR.XTBN.Y.n89 XThR.XTBN.Y.n88 152
R17421 XThR.XTBN.Y.n91 XThR.XTBN.Y.n90 152
R17422 XThR.XTBN.Y.n173 XThR.XTBN.Y.n172 152
R17423 XThR.XTBN.Y.n176 XThR.XTBN.Y.n175 152
R17424 XThR.XTBN.Y.n1 XThR.XTBN.Y.t95 139.78
R17425 XThR.XTBN.Y.n8 XThR.XTBN.Y.t44 139.78
R17426 XThR.XTBN.Y.n2 XThR.XTBN.Y.t116 139.78
R17427 XThR.XTBN.Y.n3 XThR.XTBN.Y.t35 139.78
R17428 XThR.XTBN.Y.n12 XThR.XTBN.Y.t42 139.78
R17429 XThR.XTBN.Y.n19 XThR.XTBN.Y.t112 139.78
R17430 XThR.XTBN.Y.n13 XThR.XTBN.Y.t64 139.78
R17431 XThR.XTBN.Y.n14 XThR.XTBN.Y.t107 139.78
R17432 XThR.XTBN.Y.n24 XThR.XTBN.Y.t61 139.78
R17433 XThR.XTBN.Y.n31 XThR.XTBN.Y.t14 139.78
R17434 XThR.XTBN.Y.n25 XThR.XTBN.Y.t82 139.78
R17435 XThR.XTBN.Y.n26 XThR.XTBN.Y.t122 139.78
R17436 XThR.XTBN.Y.n36 XThR.XTBN.Y.t11 139.78
R17437 XThR.XTBN.Y.n43 XThR.XTBN.Y.t79 139.78
R17438 XThR.XTBN.Y.n37 XThR.XTBN.Y.t32 139.78
R17439 XThR.XTBN.Y.n38 XThR.XTBN.Y.t71 139.78
R17440 XThR.XTBN.Y.n48 XThR.XTBN.Y.t29 139.78
R17441 XThR.XTBN.Y.n55 XThR.XTBN.Y.t98 139.78
R17442 XThR.XTBN.Y.n49 XThR.XTBN.Y.t47 139.78
R17443 XThR.XTBN.Y.n50 XThR.XTBN.Y.t90 139.78
R17444 XThR.XTBN.Y.n60 XThR.XTBN.Y.t8 139.78
R17445 XThR.XTBN.Y.n67 XThR.XTBN.Y.t74 139.78
R17446 XThR.XTBN.Y.n61 XThR.XTBN.Y.t28 139.78
R17447 XThR.XTBN.Y.n62 XThR.XTBN.Y.t67 139.78
R17448 XThR.XTBN.Y.n72 XThR.XTBN.Y.t111 139.78
R17449 XThR.XTBN.Y.n79 XThR.XTBN.Y.t62 139.78
R17450 XThR.XTBN.Y.n73 XThR.XTBN.Y.t18 139.78
R17451 XThR.XTBN.Y.n74 XThR.XTBN.Y.t53 139.78
R17452 XThR.XTBN.Y.n163 XThR.XTBN.Y.t101 139.78
R17453 XThR.XTBN.Y.n154 XThR.XTBN.Y.t52 139.78
R17454 XThR.XTBN.Y.n158 XThR.XTBN.Y.t93 139.78
R17455 XThR.XTBN.Y.n155 XThR.XTBN.Y.t16 139.78
R17456 XThR.XTBN.Y.n151 XThR.XTBN.Y.t88 139.78
R17457 XThR.XTBN.Y.n142 XThR.XTBN.Y.t37 139.78
R17458 XThR.XTBN.Y.n146 XThR.XTBN.Y.t76 139.78
R17459 XThR.XTBN.Y.n143 XThR.XTBN.Y.t118 139.78
R17460 XThR.XTBN.Y.n139 XThR.XTBN.Y.t104 139.78
R17461 XThR.XTBN.Y.n130 XThR.XTBN.Y.t55 139.78
R17462 XThR.XTBN.Y.n134 XThR.XTBN.Y.t94 139.78
R17463 XThR.XTBN.Y.n131 XThR.XTBN.Y.t17 139.78
R17464 XThR.XTBN.Y.n127 XThR.XTBN.Y.t51 139.78
R17465 XThR.XTBN.Y.n118 XThR.XTBN.Y.t4 139.78
R17466 XThR.XTBN.Y.n122 XThR.XTBN.Y.t40 139.78
R17467 XThR.XTBN.Y.n119 XThR.XTBN.Y.t84 139.78
R17468 XThR.XTBN.Y.n115 XThR.XTBN.Y.t38 139.78
R17469 XThR.XTBN.Y.n106 XThR.XTBN.Y.t109 139.78
R17470 XThR.XTBN.Y.n110 XThR.XTBN.Y.t30 139.78
R17471 XThR.XTBN.Y.n107 XThR.XTBN.Y.t70 139.78
R17472 XThR.XTBN.Y.n103 XThR.XTBN.Y.t24 139.78
R17473 XThR.XTBN.Y.n94 XThR.XTBN.Y.t91 139.78
R17474 XThR.XTBN.Y.n98 XThR.XTBN.Y.t10 139.78
R17475 XThR.XTBN.Y.n95 XThR.XTBN.Y.t48 139.78
R17476 XThR.XTBN.Y.n92 XThR.XTBN.Y.t20 139.78
R17477 XThR.XTBN.Y.n83 XThR.XTBN.Y.t120 139.78
R17478 XThR.XTBN.Y.n87 XThR.XTBN.Y.t110 139.78
R17479 XThR.XTBN.Y.n84 XThR.XTBN.Y.t103 139.78
R17480 XThR.XTBN.Y.n167 XThR.XTBN.Y.t22 139.78
R17481 XThR.XTBN.Y.n169 XThR.XTBN.Y.t58 139.78
R17482 XThR.XTBN.Y.n174 XThR.XTBN.Y.t9 139.78
R17483 XThR.XTBN.Y.n170 XThR.XTBN.Y.t78 139.78
R17484 XThR.XTBN.Y.n184 XThR.XTBN.Y.n183 101.489
R17485 XThR.XTBN.Y.n179 XThR.XTBN.Y 58.2909
R17486 XThR.XTBN.Y.n7 XThR.XTBN.Y.n6 49.6611
R17487 XThR.XTBN.Y.n18 XThR.XTBN.Y.n17 49.6611
R17488 XThR.XTBN.Y.n30 XThR.XTBN.Y.n29 49.6611
R17489 XThR.XTBN.Y.n42 XThR.XTBN.Y.n41 49.6611
R17490 XThR.XTBN.Y.n54 XThR.XTBN.Y.n53 49.6611
R17491 XThR.XTBN.Y.n66 XThR.XTBN.Y.n65 49.6611
R17492 XThR.XTBN.Y.n78 XThR.XTBN.Y.n77 49.6611
R17493 XThR.XTBN.Y.n9 XThR.XTBN.Y.n8 44.549
R17494 XThR.XTBN.Y.n20 XThR.XTBN.Y.n19 44.549
R17495 XThR.XTBN.Y.n32 XThR.XTBN.Y.n31 44.549
R17496 XThR.XTBN.Y.n44 XThR.XTBN.Y.n43 44.549
R17497 XThR.XTBN.Y.n56 XThR.XTBN.Y.n55 44.549
R17498 XThR.XTBN.Y.n68 XThR.XTBN.Y.n67 44.549
R17499 XThR.XTBN.Y.n80 XThR.XTBN.Y.n79 44.549
R17500 XThR.XTBN.Y.n4 XThR.XTBN.Y.n2 43.0884
R17501 XThR.XTBN.Y.n15 XThR.XTBN.Y.n13 43.0884
R17502 XThR.XTBN.Y.n27 XThR.XTBN.Y.n25 43.0884
R17503 XThR.XTBN.Y.n39 XThR.XTBN.Y.n37 43.0884
R17504 XThR.XTBN.Y.n51 XThR.XTBN.Y.n49 43.0884
R17505 XThR.XTBN.Y.n63 XThR.XTBN.Y.n61 43.0884
R17506 XThR.XTBN.Y.n75 XThR.XTBN.Y.n73 43.0884
R17507 XThR.XTBN.Y.n163 XThR.XTBN.Y.n162 30.6732
R17508 XThR.XTBN.Y.n162 XThR.XTBN.Y.n154 30.6732
R17509 XThR.XTBN.Y.n159 XThR.XTBN.Y.n154 30.6732
R17510 XThR.XTBN.Y.n159 XThR.XTBN.Y.n158 30.6732
R17511 XThR.XTBN.Y.n158 XThR.XTBN.Y.n157 30.6732
R17512 XThR.XTBN.Y.n157 XThR.XTBN.Y.n155 30.6732
R17513 XThR.XTBN.Y.n151 XThR.XTBN.Y.n150 30.6732
R17514 XThR.XTBN.Y.n150 XThR.XTBN.Y.n142 30.6732
R17515 XThR.XTBN.Y.n147 XThR.XTBN.Y.n142 30.6732
R17516 XThR.XTBN.Y.n147 XThR.XTBN.Y.n146 30.6732
R17517 XThR.XTBN.Y.n146 XThR.XTBN.Y.n145 30.6732
R17518 XThR.XTBN.Y.n145 XThR.XTBN.Y.n143 30.6732
R17519 XThR.XTBN.Y.n139 XThR.XTBN.Y.n138 30.6732
R17520 XThR.XTBN.Y.n138 XThR.XTBN.Y.n130 30.6732
R17521 XThR.XTBN.Y.n135 XThR.XTBN.Y.n130 30.6732
R17522 XThR.XTBN.Y.n135 XThR.XTBN.Y.n134 30.6732
R17523 XThR.XTBN.Y.n134 XThR.XTBN.Y.n133 30.6732
R17524 XThR.XTBN.Y.n133 XThR.XTBN.Y.n131 30.6732
R17525 XThR.XTBN.Y.n127 XThR.XTBN.Y.n126 30.6732
R17526 XThR.XTBN.Y.n126 XThR.XTBN.Y.n118 30.6732
R17527 XThR.XTBN.Y.n123 XThR.XTBN.Y.n118 30.6732
R17528 XThR.XTBN.Y.n123 XThR.XTBN.Y.n122 30.6732
R17529 XThR.XTBN.Y.n122 XThR.XTBN.Y.n121 30.6732
R17530 XThR.XTBN.Y.n121 XThR.XTBN.Y.n119 30.6732
R17531 XThR.XTBN.Y.n115 XThR.XTBN.Y.n114 30.6732
R17532 XThR.XTBN.Y.n114 XThR.XTBN.Y.n106 30.6732
R17533 XThR.XTBN.Y.n111 XThR.XTBN.Y.n106 30.6732
R17534 XThR.XTBN.Y.n111 XThR.XTBN.Y.n110 30.6732
R17535 XThR.XTBN.Y.n110 XThR.XTBN.Y.n109 30.6732
R17536 XThR.XTBN.Y.n109 XThR.XTBN.Y.n107 30.6732
R17537 XThR.XTBN.Y.n103 XThR.XTBN.Y.n102 30.6732
R17538 XThR.XTBN.Y.n102 XThR.XTBN.Y.n94 30.6732
R17539 XThR.XTBN.Y.n99 XThR.XTBN.Y.n94 30.6732
R17540 XThR.XTBN.Y.n99 XThR.XTBN.Y.n98 30.6732
R17541 XThR.XTBN.Y.n98 XThR.XTBN.Y.n97 30.6732
R17542 XThR.XTBN.Y.n97 XThR.XTBN.Y.n95 30.6732
R17543 XThR.XTBN.Y.n92 XThR.XTBN.Y.n91 30.6732
R17544 XThR.XTBN.Y.n91 XThR.XTBN.Y.n83 30.6732
R17545 XThR.XTBN.Y.n88 XThR.XTBN.Y.n83 30.6732
R17546 XThR.XTBN.Y.n88 XThR.XTBN.Y.n87 30.6732
R17547 XThR.XTBN.Y.n87 XThR.XTBN.Y.n86 30.6732
R17548 XThR.XTBN.Y.n86 XThR.XTBN.Y.n84 30.6732
R17549 XThR.XTBN.Y.n168 XThR.XTBN.Y.n167 30.6732
R17550 XThR.XTBN.Y.n169 XThR.XTBN.Y.n168 30.6732
R17551 XThR.XTBN.Y.n175 XThR.XTBN.Y.n169 30.6732
R17552 XThR.XTBN.Y.n175 XThR.XTBN.Y.n174 30.6732
R17553 XThR.XTBN.Y.n174 XThR.XTBN.Y.n173 30.6732
R17554 XThR.XTBN.Y.n173 XThR.XTBN.Y.n170 30.6732
R17555 XThR.XTBN.Y.n180 XThR.XTBN.Y.t3 26.5955
R17556 XThR.XTBN.Y.n180 XThR.XTBN.Y.t2 26.5955
R17557 XThR.XTBN.Y.n183 XThR.XTBN.Y.t0 24.9236
R17558 XThR.XTBN.Y.n183 XThR.XTBN.Y.t1 24.9236
R17559 XThR.XTBN.Y.n10 XThR.XTBN.Y.n0 21.7605
R17560 XThR.XTBN.Y.n21 XThR.XTBN.Y.n11 21.7605
R17561 XThR.XTBN.Y.n33 XThR.XTBN.Y.n23 21.7605
R17562 XThR.XTBN.Y.n45 XThR.XTBN.Y.n35 21.7605
R17563 XThR.XTBN.Y.n57 XThR.XTBN.Y.n47 21.7605
R17564 XThR.XTBN.Y.n69 XThR.XTBN.Y.n59 21.7605
R17565 XThR.XTBN.Y.n81 XThR.XTBN.Y.n71 21.7605
R17566 XThR.XTBN.Y.n161 XThR.XTBN.Y 18.4325
R17567 XThR.XTBN.Y.n149 XThR.XTBN.Y 18.4325
R17568 XThR.XTBN.Y.n137 XThR.XTBN.Y 18.4325
R17569 XThR.XTBN.Y.n125 XThR.XTBN.Y 18.4325
R17570 XThR.XTBN.Y.n113 XThR.XTBN.Y 18.4325
R17571 XThR.XTBN.Y.n101 XThR.XTBN.Y 18.4325
R17572 XThR.XTBN.Y.n90 XThR.XTBN.Y 18.4325
R17573 XThR.XTBN.Y.n4 XThR.XTBN.Y.n3 18.2581
R17574 XThR.XTBN.Y.n15 XThR.XTBN.Y.n14 18.2581
R17575 XThR.XTBN.Y.n27 XThR.XTBN.Y.n26 18.2581
R17576 XThR.XTBN.Y.n39 XThR.XTBN.Y.n38 18.2581
R17577 XThR.XTBN.Y.n51 XThR.XTBN.Y.n50 18.2581
R17578 XThR.XTBN.Y.n63 XThR.XTBN.Y.n62 18.2581
R17579 XThR.XTBN.Y.n75 XThR.XTBN.Y.n74 18.2581
R17580 XThR.XTBN.Y.n5 XThR.XTBN.Y 17.6005
R17581 XThR.XTBN.Y.n16 XThR.XTBN.Y 17.6005
R17582 XThR.XTBN.Y.n28 XThR.XTBN.Y 17.6005
R17583 XThR.XTBN.Y.n40 XThR.XTBN.Y 17.6005
R17584 XThR.XTBN.Y.n52 XThR.XTBN.Y 17.6005
R17585 XThR.XTBN.Y.n64 XThR.XTBN.Y 17.6005
R17586 XThR.XTBN.Y.n76 XThR.XTBN.Y 17.6005
R17587 XThR.XTBN.Y.n22 XThR.XTBN.Y.n10 17.1655
R17588 XThR.XTBN.Y.n172 XThR.XTBN.Y 17.1525
R17589 XThR.XTBN.Y XThR.XTBN.Y.n171 17.1525
R17590 XThR.XTBN.Y.n105 XThR.XTBN.Y.n93 17.054
R17591 XThR.XTBN.Y.n9 XThR.XTBN.Y.n1 16.7975
R17592 XThR.XTBN.Y.n20 XThR.XTBN.Y.n12 16.7975
R17593 XThR.XTBN.Y.n32 XThR.XTBN.Y.n24 16.7975
R17594 XThR.XTBN.Y.n44 XThR.XTBN.Y.n36 16.7975
R17595 XThR.XTBN.Y.n56 XThR.XTBN.Y.n48 16.7975
R17596 XThR.XTBN.Y.n68 XThR.XTBN.Y.n60 16.7975
R17597 XThR.XTBN.Y.n80 XThR.XTBN.Y.n72 16.7975
R17598 XThR.XTBN.Y XThR.XTBN.Y.n160 16.3845
R17599 XThR.XTBN.Y XThR.XTBN.Y.n148 16.3845
R17600 XThR.XTBN.Y XThR.XTBN.Y.n136 16.3845
R17601 XThR.XTBN.Y XThR.XTBN.Y.n124 16.3845
R17602 XThR.XTBN.Y XThR.XTBN.Y.n112 16.3845
R17603 XThR.XTBN.Y XThR.XTBN.Y.n100 16.3845
R17604 XThR.XTBN.Y XThR.XTBN.Y.n89 16.3845
R17605 XThR.XTBN.Y.n22 XThR.XTBN.Y.n21 16.0405
R17606 XThR.XTBN.Y.n34 XThR.XTBN.Y.n33 16.0405
R17607 XThR.XTBN.Y.n46 XThR.XTBN.Y.n45 16.0405
R17608 XThR.XTBN.Y.n58 XThR.XTBN.Y.n57 16.0405
R17609 XThR.XTBN.Y.n70 XThR.XTBN.Y.n69 16.0405
R17610 XThR.XTBN.Y.n82 XThR.XTBN.Y.n81 16.0405
R17611 XThR.XTBN.Y.n165 XThR.XTBN.Y.n164 15.5925
R17612 XThR.XTBN.Y.n153 XThR.XTBN.Y.n152 15.5925
R17613 XThR.XTBN.Y.n141 XThR.XTBN.Y.n140 15.5925
R17614 XThR.XTBN.Y.n129 XThR.XTBN.Y.n128 15.5925
R17615 XThR.XTBN.Y.n117 XThR.XTBN.Y.n116 15.5925
R17616 XThR.XTBN.Y.n105 XThR.XTBN.Y.n104 15.5925
R17617 XThR.XTBN.Y.n156 XThR.XTBN.Y 14.3365
R17618 XThR.XTBN.Y.n144 XThR.XTBN.Y 14.3365
R17619 XThR.XTBN.Y.n132 XThR.XTBN.Y 14.3365
R17620 XThR.XTBN.Y.n120 XThR.XTBN.Y 14.3365
R17621 XThR.XTBN.Y.n108 XThR.XTBN.Y 14.3365
R17622 XThR.XTBN.Y.n96 XThR.XTBN.Y 14.3365
R17623 XThR.XTBN.Y.n85 XThR.XTBN.Y 14.3365
R17624 XThR.XTBN.Y XThR.XTBN.Y.n182 13.5685
R17625 XThR.XTBN.Y.n177 XThR.XTBN.Y.n176 12.2885
R17626 XThR.XTBN.Y XThR.XTBN.Y.n181 10.7525
R17627 XThR.XTBN.Y.n156 XThR.XTBN.Y 9.2165
R17628 XThR.XTBN.Y.n144 XThR.XTBN.Y 9.2165
R17629 XThR.XTBN.Y.n132 XThR.XTBN.Y 9.2165
R17630 XThR.XTBN.Y.n120 XThR.XTBN.Y 9.2165
R17631 XThR.XTBN.Y.n108 XThR.XTBN.Y 9.2165
R17632 XThR.XTBN.Y.n96 XThR.XTBN.Y 9.2165
R17633 XThR.XTBN.Y.n85 XThR.XTBN.Y 9.2165
R17634 XThR.XTBN.Y.n160 XThR.XTBN.Y 7.1685
R17635 XThR.XTBN.Y.n148 XThR.XTBN.Y 7.1685
R17636 XThR.XTBN.Y.n136 XThR.XTBN.Y 7.1685
R17637 XThR.XTBN.Y.n124 XThR.XTBN.Y 7.1685
R17638 XThR.XTBN.Y.n112 XThR.XTBN.Y 7.1685
R17639 XThR.XTBN.Y.n100 XThR.XTBN.Y 7.1685
R17640 XThR.XTBN.Y.n89 XThR.XTBN.Y 7.1685
R17641 XThR.XTBN.Y.n177 XThR.XTBN.Y 6.9125
R17642 XThR.XTBN.Y.n181 XThR.XTBN.Y 6.6565
R17643 XThR.XTBN.Y.n6 XThR.XTBN.Y.n2 6.57323
R17644 XThR.XTBN.Y.n17 XThR.XTBN.Y.n13 6.57323
R17645 XThR.XTBN.Y.n29 XThR.XTBN.Y.n25 6.57323
R17646 XThR.XTBN.Y.n41 XThR.XTBN.Y.n37 6.57323
R17647 XThR.XTBN.Y.n53 XThR.XTBN.Y.n49 6.57323
R17648 XThR.XTBN.Y.n65 XThR.XTBN.Y.n61 6.57323
R17649 XThR.XTBN.Y.n77 XThR.XTBN.Y.n73 6.57323
R17650 XThR.XTBN.Y.n172 XThR.XTBN.Y 6.4005
R17651 XThR.XTBN.Y.n171 XThR.XTBN.Y 6.4005
R17652 XThR.XTBN.Y.n179 XThR.XTBN.Y.n178 5.74665
R17653 XThR.XTBN.Y.n178 XThR.XTBN.Y.n166 5.74569
R17654 XThR.XTBN.Y.n161 XThR.XTBN.Y 5.1205
R17655 XThR.XTBN.Y.n149 XThR.XTBN.Y 5.1205
R17656 XThR.XTBN.Y.n137 XThR.XTBN.Y 5.1205
R17657 XThR.XTBN.Y.n125 XThR.XTBN.Y 5.1205
R17658 XThR.XTBN.Y.n113 XThR.XTBN.Y 5.1205
R17659 XThR.XTBN.Y.n101 XThR.XTBN.Y 5.1205
R17660 XThR.XTBN.Y.n90 XThR.XTBN.Y 5.1205
R17661 XThR.XTBN.Y.n8 XThR.XTBN.Y.n7 5.11262
R17662 XThR.XTBN.Y.n19 XThR.XTBN.Y.n18 5.11262
R17663 XThR.XTBN.Y.n31 XThR.XTBN.Y.n30 5.11262
R17664 XThR.XTBN.Y.n43 XThR.XTBN.Y.n42 5.11262
R17665 XThR.XTBN.Y.n55 XThR.XTBN.Y.n54 5.11262
R17666 XThR.XTBN.Y.n67 XThR.XTBN.Y.n66 5.11262
R17667 XThR.XTBN.Y.n79 XThR.XTBN.Y.n78 5.11262
R17668 XThR.XTBN.Y.n182 XThR.XTBN.Y.n179 5.06717
R17669 XThR.XTBN.Y.n181 XThR.XTBN.Y 5.04292
R17670 XThR.XTBN.Y.n178 XThR.XTBN.Y.n177 4.6505
R17671 XThR.XTBN.Y.n176 XThR.XTBN.Y 4.3525
R17672 XThR.XTBN.Y XThR.XTBN.Y.n0 4.1605
R17673 XThR.XTBN.Y XThR.XTBN.Y.n11 4.1605
R17674 XThR.XTBN.Y XThR.XTBN.Y.n23 4.1605
R17675 XThR.XTBN.Y XThR.XTBN.Y.n35 4.1605
R17676 XThR.XTBN.Y XThR.XTBN.Y.n47 4.1605
R17677 XThR.XTBN.Y XThR.XTBN.Y.n59 4.1605
R17678 XThR.XTBN.Y XThR.XTBN.Y.n71 4.1605
R17679 XThR.XTBN.Y.n182 XThR.XTBN.Y 3.8405
R17680 XThR.XTBN.Y.n184 XThR.XTBN.Y 2.5605
R17681 XThR.XTBN.Y.n164 XThR.XTBN.Y 2.3045
R17682 XThR.XTBN.Y.n152 XThR.XTBN.Y 2.3045
R17683 XThR.XTBN.Y.n140 XThR.XTBN.Y 2.3045
R17684 XThR.XTBN.Y.n128 XThR.XTBN.Y 2.3045
R17685 XThR.XTBN.Y.n116 XThR.XTBN.Y 2.3045
R17686 XThR.XTBN.Y.n104 XThR.XTBN.Y 2.3045
R17687 XThR.XTBN.Y.n93 XThR.XTBN.Y 2.3045
R17688 XThR.XTBN.Y XThR.XTBN.Y.n184 1.93989
R17689 XThR.XTBN.Y.n166 XThR.XTBN.Y.n82 1.53415
R17690 XThR.XTBN.Y.n34 XThR.XTBN.Y.n22 1.49088
R17691 XThR.XTBN.Y.n58 XThR.XTBN.Y.n46 1.49088
R17692 XThR.XTBN.Y.n82 XThR.XTBN.Y.n70 1.48608
R17693 XThR.XTBN.Y.n153 XThR.XTBN.Y.n141 1.46204
R17694 XThR.XTBN.Y.n129 XThR.XTBN.Y.n117 1.46204
R17695 XThR.XTBN.Y.n166 XThR.XTBN.Y.n165 1.20723
R17696 XThR.XTBN.Y.n165 XThR.XTBN.Y.n153 1.15435
R17697 XThR.XTBN.Y.n141 XThR.XTBN.Y.n129 1.15435
R17698 XThR.XTBN.Y.n117 XThR.XTBN.Y.n105 1.15435
R17699 XThR.XTBN.Y.n70 XThR.XTBN.Y.n58 1.13031
R17700 XThR.XTBN.Y.n46 XThR.XTBN.Y.n34 1.1255
R17701 XThR.Tn[6].n2 XThR.Tn[6].n1 332.332
R17702 XThR.Tn[6].n2 XThR.Tn[6].n0 296.493
R17703 XThR.Tn[6] XThR.Tn[6].n82 161.363
R17704 XThR.Tn[6] XThR.Tn[6].n77 161.363
R17705 XThR.Tn[6] XThR.Tn[6].n72 161.363
R17706 XThR.Tn[6] XThR.Tn[6].n67 161.363
R17707 XThR.Tn[6] XThR.Tn[6].n62 161.363
R17708 XThR.Tn[6] XThR.Tn[6].n57 161.363
R17709 XThR.Tn[6] XThR.Tn[6].n52 161.363
R17710 XThR.Tn[6] XThR.Tn[6].n47 161.363
R17711 XThR.Tn[6] XThR.Tn[6].n42 161.363
R17712 XThR.Tn[6] XThR.Tn[6].n37 161.363
R17713 XThR.Tn[6] XThR.Tn[6].n32 161.363
R17714 XThR.Tn[6] XThR.Tn[6].n27 161.363
R17715 XThR.Tn[6] XThR.Tn[6].n22 161.363
R17716 XThR.Tn[6] XThR.Tn[6].n17 161.363
R17717 XThR.Tn[6] XThR.Tn[6].n12 161.363
R17718 XThR.Tn[6] XThR.Tn[6].n10 161.363
R17719 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R17720 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R17721 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R17722 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R17723 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R17724 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R17725 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R17726 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R17727 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R17728 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R17729 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R17730 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R17731 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R17732 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R17733 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R17734 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R17735 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R17736 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R17737 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R17738 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R17739 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R17740 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R17741 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R17742 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R17743 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R17744 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R17745 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R17746 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R17747 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R17748 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R17749 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R17750 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R17751 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R17752 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R17753 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R17754 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R17755 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R17756 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R17757 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R17758 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R17759 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R17760 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R17761 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R17762 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R17763 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R17764 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R17765 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R17766 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R17767 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R17768 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R17769 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R17770 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R17771 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R17772 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R17773 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R17774 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R17775 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R17776 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R17777 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R17778 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R17779 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R17780 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R17781 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R17782 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R17783 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R17784 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R17785 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R17786 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R17787 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R17788 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R17789 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R17790 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R17791 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R17792 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R17793 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R17794 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R17795 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R17796 XThR.Tn[6].n7 XThR.Tn[6].n5 135.249
R17797 XThR.Tn[6].n9 XThR.Tn[6].n3 98.982
R17798 XThR.Tn[6].n8 XThR.Tn[6].n4 98.982
R17799 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R17800 XThR.Tn[6].n9 XThR.Tn[6].n8 36.2672
R17801 XThR.Tn[6].n8 XThR.Tn[6].n7 36.2672
R17802 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R17803 XThR.Tn[6].n1 XThR.Tn[6].t6 26.5955
R17804 XThR.Tn[6].n1 XThR.Tn[6].t5 26.5955
R17805 XThR.Tn[6].n0 XThR.Tn[6].t7 26.5955
R17806 XThR.Tn[6].n0 XThR.Tn[6].t4 26.5955
R17807 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R17808 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R17809 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R17810 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R17811 XThR.Tn[6].n5 XThR.Tn[6].t0 24.9236
R17812 XThR.Tn[6].n5 XThR.Tn[6].t1 24.9236
R17813 XThR.Tn[6].n6 XThR.Tn[6].t3 24.9236
R17814 XThR.Tn[6].n6 XThR.Tn[6].t2 24.9236
R17815 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R17816 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R17817 XThR.Tn[6] XThR.Tn[6].n11 5.4407
R17818 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R17819 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R17820 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R17821 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R17822 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R17823 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R17824 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R17825 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R17826 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R17827 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R17828 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R17829 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R17830 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R17831 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R17832 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R17833 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R17834 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R17835 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R17836 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R17837 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R17838 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R17839 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R17840 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R17841 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R17842 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R17843 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R17844 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R17845 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R17846 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R17847 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R17848 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R17849 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R17850 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R17851 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R17852 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R17853 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R17854 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R17855 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R17856 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R17857 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R17858 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R17859 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R17860 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R17861 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R17862 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R17863 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R17864 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R17865 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R17866 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R17867 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R17868 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R17869 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R17870 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R17871 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R17872 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R17873 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R17874 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R17875 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R17876 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R17877 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R17878 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R17879 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R17880 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R17881 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R17882 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R17883 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R17884 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R17885 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R17886 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R17887 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R17888 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R17889 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R17890 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R17891 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R17892 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R17893 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R17894 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R17895 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R17896 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R17897 XThR.Tn[6] XThR.Tn[6].n87 0.038
R17898 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R17899 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R17900 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R17901 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R17902 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R17903 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R17904 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R17905 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R17906 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R17907 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R17908 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R17909 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R17910 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R17911 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R17912 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R17913 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R17914 XThR.Tn[14].n5 XThR.Tn[14].n4 256.103
R17915 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R17916 XThR.Tn[14].n88 XThR.Tn[14].n87 241.847
R17917 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R17918 XThR.Tn[14].n5 XThR.Tn[14].n3 202.095
R17919 XThR.Tn[14].n88 XThR.Tn[14].n86 185
R17920 XThR.Tn[14] XThR.Tn[14].n79 161.363
R17921 XThR.Tn[14] XThR.Tn[14].n74 161.363
R17922 XThR.Tn[14] XThR.Tn[14].n69 161.363
R17923 XThR.Tn[14] XThR.Tn[14].n64 161.363
R17924 XThR.Tn[14] XThR.Tn[14].n59 161.363
R17925 XThR.Tn[14] XThR.Tn[14].n54 161.363
R17926 XThR.Tn[14] XThR.Tn[14].n49 161.363
R17927 XThR.Tn[14] XThR.Tn[14].n44 161.363
R17928 XThR.Tn[14] XThR.Tn[14].n39 161.363
R17929 XThR.Tn[14] XThR.Tn[14].n34 161.363
R17930 XThR.Tn[14] XThR.Tn[14].n29 161.363
R17931 XThR.Tn[14] XThR.Tn[14].n24 161.363
R17932 XThR.Tn[14] XThR.Tn[14].n19 161.363
R17933 XThR.Tn[14] XThR.Tn[14].n14 161.363
R17934 XThR.Tn[14] XThR.Tn[14].n9 161.363
R17935 XThR.Tn[14] XThR.Tn[14].n7 161.363
R17936 XThR.Tn[14].n81 XThR.Tn[14].n80 161.3
R17937 XThR.Tn[14].n76 XThR.Tn[14].n75 161.3
R17938 XThR.Tn[14].n71 XThR.Tn[14].n70 161.3
R17939 XThR.Tn[14].n66 XThR.Tn[14].n65 161.3
R17940 XThR.Tn[14].n61 XThR.Tn[14].n60 161.3
R17941 XThR.Tn[14].n56 XThR.Tn[14].n55 161.3
R17942 XThR.Tn[14].n51 XThR.Tn[14].n50 161.3
R17943 XThR.Tn[14].n46 XThR.Tn[14].n45 161.3
R17944 XThR.Tn[14].n41 XThR.Tn[14].n40 161.3
R17945 XThR.Tn[14].n36 XThR.Tn[14].n35 161.3
R17946 XThR.Tn[14].n31 XThR.Tn[14].n30 161.3
R17947 XThR.Tn[14].n26 XThR.Tn[14].n25 161.3
R17948 XThR.Tn[14].n21 XThR.Tn[14].n20 161.3
R17949 XThR.Tn[14].n16 XThR.Tn[14].n15 161.3
R17950 XThR.Tn[14].n11 XThR.Tn[14].n10 161.3
R17951 XThR.Tn[14].n79 XThR.Tn[14].t51 161.106
R17952 XThR.Tn[14].n74 XThR.Tn[14].t58 161.106
R17953 XThR.Tn[14].n69 XThR.Tn[14].t39 161.106
R17954 XThR.Tn[14].n64 XThR.Tn[14].t22 161.106
R17955 XThR.Tn[14].n59 XThR.Tn[14].t49 161.106
R17956 XThR.Tn[14].n54 XThR.Tn[14].t12 161.106
R17957 XThR.Tn[14].n49 XThR.Tn[14].t56 161.106
R17958 XThR.Tn[14].n44 XThR.Tn[14].t36 161.106
R17959 XThR.Tn[14].n39 XThR.Tn[14].t19 161.106
R17960 XThR.Tn[14].n34 XThR.Tn[14].t25 161.106
R17961 XThR.Tn[14].n29 XThR.Tn[14].t73 161.106
R17962 XThR.Tn[14].n24 XThR.Tn[14].t38 161.106
R17963 XThR.Tn[14].n19 XThR.Tn[14].t72 161.106
R17964 XThR.Tn[14].n14 XThR.Tn[14].t54 161.106
R17965 XThR.Tn[14].n9 XThR.Tn[14].t13 161.106
R17966 XThR.Tn[14].n7 XThR.Tn[14].t62 161.106
R17967 XThR.Tn[14].n80 XThR.Tn[14].t32 159.978
R17968 XThR.Tn[14].n75 XThR.Tn[14].t37 159.978
R17969 XThR.Tn[14].n70 XThR.Tn[14].t20 159.978
R17970 XThR.Tn[14].n65 XThR.Tn[14].t68 159.978
R17971 XThR.Tn[14].n60 XThR.Tn[14].t30 159.978
R17972 XThR.Tn[14].n55 XThR.Tn[14].t55 159.978
R17973 XThR.Tn[14].n50 XThR.Tn[14].t35 159.978
R17974 XThR.Tn[14].n45 XThR.Tn[14].t16 159.978
R17975 XThR.Tn[14].n40 XThR.Tn[14].t66 159.978
R17976 XThR.Tn[14].n35 XThR.Tn[14].t71 159.978
R17977 XThR.Tn[14].n30 XThR.Tn[14].t53 159.978
R17978 XThR.Tn[14].n25 XThR.Tn[14].t18 159.978
R17979 XThR.Tn[14].n20 XThR.Tn[14].t52 159.978
R17980 XThR.Tn[14].n15 XThR.Tn[14].t34 159.978
R17981 XThR.Tn[14].n10 XThR.Tn[14].t60 159.978
R17982 XThR.Tn[14].n79 XThR.Tn[14].t41 145.038
R17983 XThR.Tn[14].n74 XThR.Tn[14].t65 145.038
R17984 XThR.Tn[14].n69 XThR.Tn[14].t45 145.038
R17985 XThR.Tn[14].n64 XThR.Tn[14].t26 145.038
R17986 XThR.Tn[14].n59 XThR.Tn[14].t59 145.038
R17987 XThR.Tn[14].n54 XThR.Tn[14].t40 145.038
R17988 XThR.Tn[14].n49 XThR.Tn[14].t46 145.038
R17989 XThR.Tn[14].n44 XThR.Tn[14].t27 145.038
R17990 XThR.Tn[14].n39 XThR.Tn[14].t23 145.038
R17991 XThR.Tn[14].n34 XThR.Tn[14].t57 145.038
R17992 XThR.Tn[14].n29 XThR.Tn[14].t15 145.038
R17993 XThR.Tn[14].n24 XThR.Tn[14].t44 145.038
R17994 XThR.Tn[14].n19 XThR.Tn[14].t14 145.038
R17995 XThR.Tn[14].n14 XThR.Tn[14].t64 145.038
R17996 XThR.Tn[14].n9 XThR.Tn[14].t24 145.038
R17997 XThR.Tn[14].n7 XThR.Tn[14].t69 145.038
R17998 XThR.Tn[14].n80 XThR.Tn[14].t43 143.911
R17999 XThR.Tn[14].n75 XThR.Tn[14].t70 143.911
R18000 XThR.Tn[14].n70 XThR.Tn[14].t48 143.911
R18001 XThR.Tn[14].n65 XThR.Tn[14].t31 143.911
R18002 XThR.Tn[14].n60 XThR.Tn[14].t63 143.911
R18003 XThR.Tn[14].n55 XThR.Tn[14].t42 143.911
R18004 XThR.Tn[14].n50 XThR.Tn[14].t50 143.911
R18005 XThR.Tn[14].n45 XThR.Tn[14].t33 143.911
R18006 XThR.Tn[14].n40 XThR.Tn[14].t29 143.911
R18007 XThR.Tn[14].n35 XThR.Tn[14].t61 143.911
R18008 XThR.Tn[14].n30 XThR.Tn[14].t21 143.911
R18009 XThR.Tn[14].n25 XThR.Tn[14].t47 143.911
R18010 XThR.Tn[14].n20 XThR.Tn[14].t17 143.911
R18011 XThR.Tn[14].n15 XThR.Tn[14].t67 143.911
R18012 XThR.Tn[14].n10 XThR.Tn[14].t28 143.911
R18013 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R18014 XThR.Tn[14].n3 XThR.Tn[14].t6 26.5955
R18015 XThR.Tn[14].n3 XThR.Tn[14].t7 26.5955
R18016 XThR.Tn[14].n4 XThR.Tn[14].t4 26.5955
R18017 XThR.Tn[14].n4 XThR.Tn[14].t5 26.5955
R18018 XThR.Tn[14].n0 XThR.Tn[14].t8 26.5955
R18019 XThR.Tn[14].n0 XThR.Tn[14].t9 26.5955
R18020 XThR.Tn[14].n1 XThR.Tn[14].t10 26.5955
R18021 XThR.Tn[14].n1 XThR.Tn[14].t11 26.5955
R18022 XThR.Tn[14].n86 XThR.Tn[14].t0 24.9236
R18023 XThR.Tn[14].n86 XThR.Tn[14].t1 24.9236
R18024 XThR.Tn[14].n87 XThR.Tn[14].t2 24.9236
R18025 XThR.Tn[14].n87 XThR.Tn[14].t3 24.9236
R18026 XThR.Tn[14] XThR.Tn[14].n88 18.8943
R18027 XThR.Tn[14].n6 XThR.Tn[14].n5 13.5534
R18028 XThR.Tn[14].n85 XThR.Tn[14] 8.47191
R18029 XThR.Tn[14] XThR.Tn[14].n85 6.34069
R18030 XThR.Tn[14] XThR.Tn[14].n8 5.4407
R18031 XThR.Tn[14].n13 XThR.Tn[14].n12 4.5005
R18032 XThR.Tn[14].n18 XThR.Tn[14].n17 4.5005
R18033 XThR.Tn[14].n23 XThR.Tn[14].n22 4.5005
R18034 XThR.Tn[14].n28 XThR.Tn[14].n27 4.5005
R18035 XThR.Tn[14].n33 XThR.Tn[14].n32 4.5005
R18036 XThR.Tn[14].n38 XThR.Tn[14].n37 4.5005
R18037 XThR.Tn[14].n43 XThR.Tn[14].n42 4.5005
R18038 XThR.Tn[14].n48 XThR.Tn[14].n47 4.5005
R18039 XThR.Tn[14].n53 XThR.Tn[14].n52 4.5005
R18040 XThR.Tn[14].n58 XThR.Tn[14].n57 4.5005
R18041 XThR.Tn[14].n63 XThR.Tn[14].n62 4.5005
R18042 XThR.Tn[14].n68 XThR.Tn[14].n67 4.5005
R18043 XThR.Tn[14].n73 XThR.Tn[14].n72 4.5005
R18044 XThR.Tn[14].n78 XThR.Tn[14].n77 4.5005
R18045 XThR.Tn[14].n83 XThR.Tn[14].n82 4.5005
R18046 XThR.Tn[14].n84 XThR.Tn[14] 3.70586
R18047 XThR.Tn[14].n13 XThR.Tn[14] 2.52282
R18048 XThR.Tn[14].n18 XThR.Tn[14] 2.52282
R18049 XThR.Tn[14].n23 XThR.Tn[14] 2.52282
R18050 XThR.Tn[14].n28 XThR.Tn[14] 2.52282
R18051 XThR.Tn[14].n33 XThR.Tn[14] 2.52282
R18052 XThR.Tn[14].n38 XThR.Tn[14] 2.52282
R18053 XThR.Tn[14].n43 XThR.Tn[14] 2.52282
R18054 XThR.Tn[14].n48 XThR.Tn[14] 2.52282
R18055 XThR.Tn[14].n53 XThR.Tn[14] 2.52282
R18056 XThR.Tn[14].n58 XThR.Tn[14] 2.52282
R18057 XThR.Tn[14].n63 XThR.Tn[14] 2.52282
R18058 XThR.Tn[14].n68 XThR.Tn[14] 2.52282
R18059 XThR.Tn[14].n73 XThR.Tn[14] 2.52282
R18060 XThR.Tn[14].n78 XThR.Tn[14] 2.52282
R18061 XThR.Tn[14].n83 XThR.Tn[14] 2.52282
R18062 XThR.Tn[14].n85 XThR.Tn[14] 1.79489
R18063 XThR.Tn[14].n6 XThR.Tn[14] 1.50638
R18064 XThR.Tn[14] XThR.Tn[14].n6 1.19676
R18065 XThR.Tn[14].n81 XThR.Tn[14] 1.08677
R18066 XThR.Tn[14].n76 XThR.Tn[14] 1.08677
R18067 XThR.Tn[14].n71 XThR.Tn[14] 1.08677
R18068 XThR.Tn[14].n66 XThR.Tn[14] 1.08677
R18069 XThR.Tn[14].n61 XThR.Tn[14] 1.08677
R18070 XThR.Tn[14].n56 XThR.Tn[14] 1.08677
R18071 XThR.Tn[14].n51 XThR.Tn[14] 1.08677
R18072 XThR.Tn[14].n46 XThR.Tn[14] 1.08677
R18073 XThR.Tn[14].n41 XThR.Tn[14] 1.08677
R18074 XThR.Tn[14].n36 XThR.Tn[14] 1.08677
R18075 XThR.Tn[14].n31 XThR.Tn[14] 1.08677
R18076 XThR.Tn[14].n26 XThR.Tn[14] 1.08677
R18077 XThR.Tn[14].n21 XThR.Tn[14] 1.08677
R18078 XThR.Tn[14].n16 XThR.Tn[14] 1.08677
R18079 XThR.Tn[14].n11 XThR.Tn[14] 1.08677
R18080 XThR.Tn[14] XThR.Tn[14].n13 0.839786
R18081 XThR.Tn[14] XThR.Tn[14].n18 0.839786
R18082 XThR.Tn[14] XThR.Tn[14].n23 0.839786
R18083 XThR.Tn[14] XThR.Tn[14].n28 0.839786
R18084 XThR.Tn[14] XThR.Tn[14].n33 0.839786
R18085 XThR.Tn[14] XThR.Tn[14].n38 0.839786
R18086 XThR.Tn[14] XThR.Tn[14].n43 0.839786
R18087 XThR.Tn[14] XThR.Tn[14].n48 0.839786
R18088 XThR.Tn[14] XThR.Tn[14].n53 0.839786
R18089 XThR.Tn[14] XThR.Tn[14].n58 0.839786
R18090 XThR.Tn[14] XThR.Tn[14].n63 0.839786
R18091 XThR.Tn[14] XThR.Tn[14].n68 0.839786
R18092 XThR.Tn[14] XThR.Tn[14].n73 0.839786
R18093 XThR.Tn[14] XThR.Tn[14].n78 0.839786
R18094 XThR.Tn[14] XThR.Tn[14].n83 0.839786
R18095 XThR.Tn[14].n8 XThR.Tn[14] 0.499542
R18096 XThR.Tn[14].n82 XThR.Tn[14] 0.063
R18097 XThR.Tn[14].n77 XThR.Tn[14] 0.063
R18098 XThR.Tn[14].n72 XThR.Tn[14] 0.063
R18099 XThR.Tn[14].n67 XThR.Tn[14] 0.063
R18100 XThR.Tn[14].n62 XThR.Tn[14] 0.063
R18101 XThR.Tn[14].n57 XThR.Tn[14] 0.063
R18102 XThR.Tn[14].n52 XThR.Tn[14] 0.063
R18103 XThR.Tn[14].n47 XThR.Tn[14] 0.063
R18104 XThR.Tn[14].n42 XThR.Tn[14] 0.063
R18105 XThR.Tn[14].n37 XThR.Tn[14] 0.063
R18106 XThR.Tn[14].n32 XThR.Tn[14] 0.063
R18107 XThR.Tn[14].n27 XThR.Tn[14] 0.063
R18108 XThR.Tn[14].n22 XThR.Tn[14] 0.063
R18109 XThR.Tn[14].n17 XThR.Tn[14] 0.063
R18110 XThR.Tn[14].n12 XThR.Tn[14] 0.063
R18111 XThR.Tn[14].n84 XThR.Tn[14] 0.0540714
R18112 XThR.Tn[14] XThR.Tn[14].n84 0.038
R18113 XThR.Tn[14].n8 XThR.Tn[14] 0.0143889
R18114 XThR.Tn[14].n82 XThR.Tn[14].n81 0.00771154
R18115 XThR.Tn[14].n77 XThR.Tn[14].n76 0.00771154
R18116 XThR.Tn[14].n72 XThR.Tn[14].n71 0.00771154
R18117 XThR.Tn[14].n67 XThR.Tn[14].n66 0.00771154
R18118 XThR.Tn[14].n62 XThR.Tn[14].n61 0.00771154
R18119 XThR.Tn[14].n57 XThR.Tn[14].n56 0.00771154
R18120 XThR.Tn[14].n52 XThR.Tn[14].n51 0.00771154
R18121 XThR.Tn[14].n47 XThR.Tn[14].n46 0.00771154
R18122 XThR.Tn[14].n42 XThR.Tn[14].n41 0.00771154
R18123 XThR.Tn[14].n37 XThR.Tn[14].n36 0.00771154
R18124 XThR.Tn[14].n32 XThR.Tn[14].n31 0.00771154
R18125 XThR.Tn[14].n27 XThR.Tn[14].n26 0.00771154
R18126 XThR.Tn[14].n22 XThR.Tn[14].n21 0.00771154
R18127 XThR.Tn[14].n17 XThR.Tn[14].n16 0.00771154
R18128 XThR.Tn[14].n12 XThR.Tn[14].n11 0.00771154
R18129 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R18130 XThR.Tn[12].n2 XThR.Tn[12].n1 243.679
R18131 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R18132 XThR.Tn[12].n2 XThR.Tn[12].n0 205.28
R18133 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R18134 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R18135 XThR.Tn[12] XThR.Tn[12].n78 161.363
R18136 XThR.Tn[12] XThR.Tn[12].n73 161.363
R18137 XThR.Tn[12] XThR.Tn[12].n68 161.363
R18138 XThR.Tn[12] XThR.Tn[12].n63 161.363
R18139 XThR.Tn[12] XThR.Tn[12].n58 161.363
R18140 XThR.Tn[12] XThR.Tn[12].n53 161.363
R18141 XThR.Tn[12] XThR.Tn[12].n48 161.363
R18142 XThR.Tn[12] XThR.Tn[12].n43 161.363
R18143 XThR.Tn[12] XThR.Tn[12].n38 161.363
R18144 XThR.Tn[12] XThR.Tn[12].n33 161.363
R18145 XThR.Tn[12] XThR.Tn[12].n28 161.363
R18146 XThR.Tn[12] XThR.Tn[12].n23 161.363
R18147 XThR.Tn[12] XThR.Tn[12].n18 161.363
R18148 XThR.Tn[12] XThR.Tn[12].n13 161.363
R18149 XThR.Tn[12] XThR.Tn[12].n8 161.363
R18150 XThR.Tn[12] XThR.Tn[12].n6 161.363
R18151 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R18152 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R18153 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R18154 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R18155 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R18156 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R18157 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R18158 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R18159 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R18160 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R18161 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R18162 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R18163 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R18164 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R18165 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R18166 XThR.Tn[12].n78 XThR.Tn[12].t18 161.106
R18167 XThR.Tn[12].n73 XThR.Tn[12].t24 161.106
R18168 XThR.Tn[12].n68 XThR.Tn[12].t67 161.106
R18169 XThR.Tn[12].n63 XThR.Tn[12].t52 161.106
R18170 XThR.Tn[12].n58 XThR.Tn[12].t16 161.106
R18171 XThR.Tn[12].n53 XThR.Tn[12].t40 161.106
R18172 XThR.Tn[12].n48 XThR.Tn[12].t22 161.106
R18173 XThR.Tn[12].n43 XThR.Tn[12].t65 161.106
R18174 XThR.Tn[12].n38 XThR.Tn[12].t51 161.106
R18175 XThR.Tn[12].n33 XThR.Tn[12].t56 161.106
R18176 XThR.Tn[12].n28 XThR.Tn[12].t39 161.106
R18177 XThR.Tn[12].n23 XThR.Tn[12].t66 161.106
R18178 XThR.Tn[12].n18 XThR.Tn[12].t38 161.106
R18179 XThR.Tn[12].n13 XThR.Tn[12].t20 161.106
R18180 XThR.Tn[12].n8 XThR.Tn[12].t43 161.106
R18181 XThR.Tn[12].n6 XThR.Tn[12].t28 161.106
R18182 XThR.Tn[12].n79 XThR.Tn[12].t58 159.978
R18183 XThR.Tn[12].n74 XThR.Tn[12].t62 159.978
R18184 XThR.Tn[12].n69 XThR.Tn[12].t47 159.978
R18185 XThR.Tn[12].n64 XThR.Tn[12].t31 159.978
R18186 XThR.Tn[12].n59 XThR.Tn[12].t55 159.978
R18187 XThR.Tn[12].n54 XThR.Tn[12].t19 159.978
R18188 XThR.Tn[12].n49 XThR.Tn[12].t61 159.978
R18189 XThR.Tn[12].n44 XThR.Tn[12].t44 159.978
R18190 XThR.Tn[12].n39 XThR.Tn[12].t29 159.978
R18191 XThR.Tn[12].n34 XThR.Tn[12].t37 159.978
R18192 XThR.Tn[12].n29 XThR.Tn[12].t17 159.978
R18193 XThR.Tn[12].n24 XThR.Tn[12].t46 159.978
R18194 XThR.Tn[12].n19 XThR.Tn[12].t15 159.978
R18195 XThR.Tn[12].n14 XThR.Tn[12].t60 159.978
R18196 XThR.Tn[12].n9 XThR.Tn[12].t21 159.978
R18197 XThR.Tn[12].n78 XThR.Tn[12].t69 145.038
R18198 XThR.Tn[12].n73 XThR.Tn[12].t32 145.038
R18199 XThR.Tn[12].n68 XThR.Tn[12].t73 145.038
R18200 XThR.Tn[12].n63 XThR.Tn[12].t57 145.038
R18201 XThR.Tn[12].n58 XThR.Tn[12].t25 145.038
R18202 XThR.Tn[12].n53 XThR.Tn[12].t68 145.038
R18203 XThR.Tn[12].n48 XThR.Tn[12].t12 145.038
R18204 XThR.Tn[12].n43 XThR.Tn[12].t59 145.038
R18205 XThR.Tn[12].n38 XThR.Tn[12].t54 145.038
R18206 XThR.Tn[12].n33 XThR.Tn[12].t23 145.038
R18207 XThR.Tn[12].n28 XThR.Tn[12].t48 145.038
R18208 XThR.Tn[12].n23 XThR.Tn[12].t70 145.038
R18209 XThR.Tn[12].n18 XThR.Tn[12].t45 145.038
R18210 XThR.Tn[12].n13 XThR.Tn[12].t30 145.038
R18211 XThR.Tn[12].n8 XThR.Tn[12].t53 145.038
R18212 XThR.Tn[12].n6 XThR.Tn[12].t36 145.038
R18213 XThR.Tn[12].n79 XThR.Tn[12].t27 143.911
R18214 XThR.Tn[12].n74 XThR.Tn[12].t50 143.911
R18215 XThR.Tn[12].n69 XThR.Tn[12].t34 143.911
R18216 XThR.Tn[12].n64 XThR.Tn[12].t13 143.911
R18217 XThR.Tn[12].n59 XThR.Tn[12].t42 143.911
R18218 XThR.Tn[12].n54 XThR.Tn[12].t26 143.911
R18219 XThR.Tn[12].n49 XThR.Tn[12].t35 143.911
R18220 XThR.Tn[12].n44 XThR.Tn[12].t14 143.911
R18221 XThR.Tn[12].n39 XThR.Tn[12].t72 143.911
R18222 XThR.Tn[12].n34 XThR.Tn[12].t41 143.911
R18223 XThR.Tn[12].n29 XThR.Tn[12].t64 143.911
R18224 XThR.Tn[12].n24 XThR.Tn[12].t33 143.911
R18225 XThR.Tn[12].n19 XThR.Tn[12].t63 143.911
R18226 XThR.Tn[12].n14 XThR.Tn[12].t49 143.911
R18227 XThR.Tn[12].n9 XThR.Tn[12].t71 143.911
R18228 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R18229 XThR.Tn[12].n85 XThR.Tn[12].t10 26.5955
R18230 XThR.Tn[12].n85 XThR.Tn[12].t8 26.5955
R18231 XThR.Tn[12].n86 XThR.Tn[12].t11 26.5955
R18232 XThR.Tn[12].n86 XThR.Tn[12].t9 26.5955
R18233 XThR.Tn[12].n0 XThR.Tn[12].t0 26.5955
R18234 XThR.Tn[12].n0 XThR.Tn[12].t2 26.5955
R18235 XThR.Tn[12].n1 XThR.Tn[12].t3 26.5955
R18236 XThR.Tn[12].n1 XThR.Tn[12].t1 26.5955
R18237 XThR.Tn[12].n4 XThR.Tn[12].t6 24.9236
R18238 XThR.Tn[12].n4 XThR.Tn[12].t4 24.9236
R18239 XThR.Tn[12].n3 XThR.Tn[12].t7 24.9236
R18240 XThR.Tn[12].n3 XThR.Tn[12].t5 24.9236
R18241 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R18242 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R18243 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R18244 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R18245 XThR.Tn[12] XThR.Tn[12].n7 5.4407
R18246 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R18247 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R18248 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R18249 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R18250 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R18251 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R18252 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R18253 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R18254 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R18255 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R18256 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R18257 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R18258 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R18259 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R18260 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R18261 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R18262 XThR.Tn[12].n12 XThR.Tn[12] 2.52282
R18263 XThR.Tn[12].n17 XThR.Tn[12] 2.52282
R18264 XThR.Tn[12].n22 XThR.Tn[12] 2.52282
R18265 XThR.Tn[12].n27 XThR.Tn[12] 2.52282
R18266 XThR.Tn[12].n32 XThR.Tn[12] 2.52282
R18267 XThR.Tn[12].n37 XThR.Tn[12] 2.52282
R18268 XThR.Tn[12].n42 XThR.Tn[12] 2.52282
R18269 XThR.Tn[12].n47 XThR.Tn[12] 2.52282
R18270 XThR.Tn[12].n52 XThR.Tn[12] 2.52282
R18271 XThR.Tn[12].n57 XThR.Tn[12] 2.52282
R18272 XThR.Tn[12].n62 XThR.Tn[12] 2.52282
R18273 XThR.Tn[12].n67 XThR.Tn[12] 2.52282
R18274 XThR.Tn[12].n72 XThR.Tn[12] 2.52282
R18275 XThR.Tn[12].n77 XThR.Tn[12] 2.52282
R18276 XThR.Tn[12].n82 XThR.Tn[12] 2.52282
R18277 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R18278 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R18279 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R18280 XThR.Tn[12].n80 XThR.Tn[12] 1.08677
R18281 XThR.Tn[12].n75 XThR.Tn[12] 1.08677
R18282 XThR.Tn[12].n70 XThR.Tn[12] 1.08677
R18283 XThR.Tn[12].n65 XThR.Tn[12] 1.08677
R18284 XThR.Tn[12].n60 XThR.Tn[12] 1.08677
R18285 XThR.Tn[12].n55 XThR.Tn[12] 1.08677
R18286 XThR.Tn[12].n50 XThR.Tn[12] 1.08677
R18287 XThR.Tn[12].n45 XThR.Tn[12] 1.08677
R18288 XThR.Tn[12].n40 XThR.Tn[12] 1.08677
R18289 XThR.Tn[12].n35 XThR.Tn[12] 1.08677
R18290 XThR.Tn[12].n30 XThR.Tn[12] 1.08677
R18291 XThR.Tn[12].n25 XThR.Tn[12] 1.08677
R18292 XThR.Tn[12].n20 XThR.Tn[12] 1.08677
R18293 XThR.Tn[12].n15 XThR.Tn[12] 1.08677
R18294 XThR.Tn[12].n10 XThR.Tn[12] 1.08677
R18295 XThR.Tn[12] XThR.Tn[12].n12 0.839786
R18296 XThR.Tn[12] XThR.Tn[12].n17 0.839786
R18297 XThR.Tn[12] XThR.Tn[12].n22 0.839786
R18298 XThR.Tn[12] XThR.Tn[12].n27 0.839786
R18299 XThR.Tn[12] XThR.Tn[12].n32 0.839786
R18300 XThR.Tn[12] XThR.Tn[12].n37 0.839786
R18301 XThR.Tn[12] XThR.Tn[12].n42 0.839786
R18302 XThR.Tn[12] XThR.Tn[12].n47 0.839786
R18303 XThR.Tn[12] XThR.Tn[12].n52 0.839786
R18304 XThR.Tn[12] XThR.Tn[12].n57 0.839786
R18305 XThR.Tn[12] XThR.Tn[12].n62 0.839786
R18306 XThR.Tn[12] XThR.Tn[12].n67 0.839786
R18307 XThR.Tn[12] XThR.Tn[12].n72 0.839786
R18308 XThR.Tn[12] XThR.Tn[12].n77 0.839786
R18309 XThR.Tn[12] XThR.Tn[12].n82 0.839786
R18310 XThR.Tn[12].n7 XThR.Tn[12] 0.499542
R18311 XThR.Tn[12].n81 XThR.Tn[12] 0.063
R18312 XThR.Tn[12].n76 XThR.Tn[12] 0.063
R18313 XThR.Tn[12].n71 XThR.Tn[12] 0.063
R18314 XThR.Tn[12].n66 XThR.Tn[12] 0.063
R18315 XThR.Tn[12].n61 XThR.Tn[12] 0.063
R18316 XThR.Tn[12].n56 XThR.Tn[12] 0.063
R18317 XThR.Tn[12].n51 XThR.Tn[12] 0.063
R18318 XThR.Tn[12].n46 XThR.Tn[12] 0.063
R18319 XThR.Tn[12].n41 XThR.Tn[12] 0.063
R18320 XThR.Tn[12].n36 XThR.Tn[12] 0.063
R18321 XThR.Tn[12].n31 XThR.Tn[12] 0.063
R18322 XThR.Tn[12].n26 XThR.Tn[12] 0.063
R18323 XThR.Tn[12].n21 XThR.Tn[12] 0.063
R18324 XThR.Tn[12].n16 XThR.Tn[12] 0.063
R18325 XThR.Tn[12].n11 XThR.Tn[12] 0.063
R18326 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R18327 XThR.Tn[12] XThR.Tn[12].n83 0.038
R18328 XThR.Tn[12].n7 XThR.Tn[12] 0.0143889
R18329 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00771154
R18330 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00771154
R18331 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00771154
R18332 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00771154
R18333 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00771154
R18334 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00771154
R18335 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00771154
R18336 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00771154
R18337 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00771154
R18338 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00771154
R18339 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00771154
R18340 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00771154
R18341 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00771154
R18342 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00771154
R18343 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00771154
R18344 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R18345 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R18346 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R18347 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R18348 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R18349 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R18350 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R18351 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R18352 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R18353 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R18354 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R18355 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R18356 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R18357 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R18358 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R18359 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R18360 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R18361 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R18362 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R18363 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R18364 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R18365 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R18366 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R18367 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R18368 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R18369 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R18370 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R18371 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R18372 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R18373 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R18374 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R18375 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R18376 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R18377 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R18378 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R18379 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R18380 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R18381 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R18382 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R18383 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R18384 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R18385 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R18386 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R18387 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R18388 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R18389 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R18390 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R18391 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R18392 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R18393 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R18394 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R18395 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R18396 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R18397 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R18398 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R18399 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R18400 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R18401 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R18402 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R18403 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R18404 XThC.XTBN.Y.n189 XThC.XTBN.Y.n188 208.965
R18405 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R18406 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R18407 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R18408 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R18409 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R18410 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R18411 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R18412 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R18413 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R18414 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R18415 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R18416 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R18417 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R18418 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R18419 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R18420 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R18421 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R18422 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R18423 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R18424 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R18425 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R18426 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R18427 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R18428 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R18429 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R18430 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R18431 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R18432 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R18433 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R18434 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R18435 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R18436 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R18437 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R18438 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R18439 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R18440 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R18441 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R18442 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R18443 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R18444 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R18445 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R18446 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R18447 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R18448 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R18449 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R18450 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R18451 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R18452 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R18453 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R18454 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R18455 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R18456 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R18457 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R18458 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R18459 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R18460 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R18461 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R18462 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R18463 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R18464 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R18465 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R18466 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R18467 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R18468 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R18469 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R18470 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R18471 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R18472 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R18473 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R18474 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R18475 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R18476 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R18477 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R18478 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R18479 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R18480 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R18481 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R18482 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R18483 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R18484 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R18485 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R18486 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R18487 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R18488 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R18489 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R18490 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R18491 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R18492 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R18493 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R18494 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R18495 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R18496 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R18497 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R18498 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R18499 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R18500 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R18501 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R18502 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R18503 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R18504 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R18505 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R18506 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R18507 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R18508 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R18509 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R18510 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R18511 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R18512 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R18513 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R18514 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R18515 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R18516 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R18517 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R18518 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R18519 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R18520 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R18521 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R18522 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R18523 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R18524 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R18525 XThC.XTBN.Y XThC.XTBN.Y.n192 96.8352
R18526 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R18527 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R18528 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R18529 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R18530 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R18531 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R18532 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R18533 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R18534 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R18535 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R18536 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R18537 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R18538 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R18539 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R18540 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R18541 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R18542 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R18543 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R18544 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R18545 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R18546 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R18547 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R18548 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R18549 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R18550 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R18551 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R18552 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R18553 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R18554 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R18555 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R18556 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R18557 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R18558 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R18559 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R18560 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R18561 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R18562 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R18563 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R18564 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R18565 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R18566 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R18567 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R18568 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R18569 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R18570 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R18571 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R18572 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R18573 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R18574 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R18575 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R18576 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R18577 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R18578 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R18579 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R18580 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R18581 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R18582 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R18583 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R18584 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R18585 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R18586 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R18587 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R18588 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R18589 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R18590 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R18591 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R18592 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R18593 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R18594 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R18595 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R18596 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 26.5955
R18597 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 26.5955
R18598 XThC.XTBN.Y.n192 XThC.XTBN.Y.t1 24.9236
R18599 XThC.XTBN.Y.n192 XThC.XTBN.Y.t0 24.9236
R18600 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R18601 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R18602 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R18603 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R18604 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R18605 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R18606 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R18607 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R18608 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R18609 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R18610 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R18611 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R18612 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R18613 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R18614 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R18615 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R18616 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R18617 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R18618 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R18619 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R18620 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R18621 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R18622 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R18623 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R18624 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R18625 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R18626 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R18627 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R18628 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R18629 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R18630 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R18631 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R18632 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R18633 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R18634 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R18635 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R18636 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R18637 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R18638 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R18639 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R18640 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R18641 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R18642 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R18643 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R18644 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R18645 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R18646 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R18647 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R18648 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R18649 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R18650 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R18651 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R18652 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R18653 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R18654 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R18655 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R18656 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R18657 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R18658 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R18659 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R18660 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R18661 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R18662 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R18663 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R18664 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R18665 XThC.XTBN.Y.n190 XThC.XTBN.Y 12.5445
R18666 XThC.XTBN.Y.n191 XThC.XTBN.Y 11.2645
R18667 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R18668 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R18669 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R18670 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R18671 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R18672 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R18673 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R18674 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R18675 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R18676 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R18677 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R18678 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R18679 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R18680 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R18681 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R18682 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R18683 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R18684 XThC.XTBN.Y.n191 XThC.XTBN.Y 6.1445
R18685 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R18686 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R18687 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R18688 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R18689 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R18690 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R18691 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R18692 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R18693 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R18694 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R18695 XThC.XTBN.Y XThC.XTBN.Y.n190 4.8645
R18696 XThC.XTBN.Y XThC.XTBN.Y.n191 4.65505
R18697 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R18698 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R18699 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R18700 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R18701 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R18702 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R18703 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R18704 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R18705 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R18706 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R18707 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R18708 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R18709 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R18710 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R18711 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R18712 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R18713 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R18714 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R18715 XThC.XTBN.Y XThC.XTBN.Y.n189 2.0485
R18716 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R18717 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R18718 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R18719 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R18720 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R18721 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R18722 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R18723 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R18724 XThC.XTBN.Y.n189 XThC.XTBN.Y 1.55202
R18725 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R18726 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R18727 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R18728 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R18729 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R18730 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R18731 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R18732 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R18733 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R18734 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R18735 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R18736 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R18737 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R18738 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R18739 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R18740 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R18741 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R18742 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R18743 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R18744 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R18745 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R18746 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R18747 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R18748 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R18749 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R18750 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R18751 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R18752 XThC.Tn[6].n12 XThC.Tn[6].n10 161.406
R18753 XThC.Tn[6].n15 XThC.Tn[6].n13 161.406
R18754 XThC.Tn[6].n18 XThC.Tn[6].n16 161.406
R18755 XThC.Tn[6].n21 XThC.Tn[6].n19 161.406
R18756 XThC.Tn[6].n24 XThC.Tn[6].n22 161.406
R18757 XThC.Tn[6].n27 XThC.Tn[6].n25 161.406
R18758 XThC.Tn[6].n30 XThC.Tn[6].n28 161.406
R18759 XThC.Tn[6].n33 XThC.Tn[6].n31 161.406
R18760 XThC.Tn[6].n36 XThC.Tn[6].n34 161.406
R18761 XThC.Tn[6].n39 XThC.Tn[6].n37 161.406
R18762 XThC.Tn[6].n42 XThC.Tn[6].n40 161.406
R18763 XThC.Tn[6].n45 XThC.Tn[6].n43 161.406
R18764 XThC.Tn[6].n48 XThC.Tn[6].n46 161.406
R18765 XThC.Tn[6].n51 XThC.Tn[6].n49 161.406
R18766 XThC.Tn[6].n54 XThC.Tn[6].n52 161.406
R18767 XThC.Tn[6].n57 XThC.Tn[6].n55 161.406
R18768 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R18769 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R18770 XThC.Tn[6].n16 XThC.Tn[6].t17 161.202
R18771 XThC.Tn[6].n19 XThC.Tn[6].t18 161.202
R18772 XThC.Tn[6].n22 XThC.Tn[6].t37 161.202
R18773 XThC.Tn[6].n25 XThC.Tn[6].t38 161.202
R18774 XThC.Tn[6].n28 XThC.Tn[6].t22 161.202
R18775 XThC.Tn[6].n31 XThC.Tn[6].t29 161.202
R18776 XThC.Tn[6].n34 XThC.Tn[6].t31 161.202
R18777 XThC.Tn[6].n37 XThC.Tn[6].t19 161.202
R18778 XThC.Tn[6].n40 XThC.Tn[6].t21 161.202
R18779 XThC.Tn[6].n43 XThC.Tn[6].t32 161.202
R18780 XThC.Tn[6].n46 XThC.Tn[6].t41 161.202
R18781 XThC.Tn[6].n49 XThC.Tn[6].t43 161.202
R18782 XThC.Tn[6].n52 XThC.Tn[6].t24 161.202
R18783 XThC.Tn[6].n55 XThC.Tn[6].t34 161.202
R18784 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R18785 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R18786 XThC.Tn[6].n16 XThC.Tn[6].t42 145.137
R18787 XThC.Tn[6].n19 XThC.Tn[6].t12 145.137
R18788 XThC.Tn[6].n22 XThC.Tn[6].t33 145.137
R18789 XThC.Tn[6].n25 XThC.Tn[6].t35 145.137
R18790 XThC.Tn[6].n28 XThC.Tn[6].t16 145.137
R18791 XThC.Tn[6].n31 XThC.Tn[6].t25 145.137
R18792 XThC.Tn[6].n34 XThC.Tn[6].t27 145.137
R18793 XThC.Tn[6].n37 XThC.Tn[6].t14 145.137
R18794 XThC.Tn[6].n40 XThC.Tn[6].t15 145.137
R18795 XThC.Tn[6].n43 XThC.Tn[6].t28 145.137
R18796 XThC.Tn[6].n46 XThC.Tn[6].t36 145.137
R18797 XThC.Tn[6].n49 XThC.Tn[6].t39 145.137
R18798 XThC.Tn[6].n52 XThC.Tn[6].t20 145.137
R18799 XThC.Tn[6].n55 XThC.Tn[6].t30 145.137
R18800 XThC.Tn[6].n5 XThC.Tn[6].n3 135.248
R18801 XThC.Tn[6].n5 XThC.Tn[6].n4 98.982
R18802 XThC.Tn[6].n7 XThC.Tn[6].n6 98.982
R18803 XThC.Tn[6].n9 XThC.Tn[6].n8 98.982
R18804 XThC.Tn[6].n7 XThC.Tn[6].n5 36.2672
R18805 XThC.Tn[6].n9 XThC.Tn[6].n7 36.2672
R18806 XThC.Tn[6].n59 XThC.Tn[6].n9 32.6405
R18807 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R18808 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R18809 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R18810 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R18811 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R18812 XThC.Tn[6].n3 XThC.Tn[6].t10 24.9236
R18813 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R18814 XThC.Tn[6].n4 XThC.Tn[6].t8 24.9236
R18815 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R18816 XThC.Tn[6].n6 XThC.Tn[6].t1 24.9236
R18817 XThC.Tn[6].n8 XThC.Tn[6].t0 24.9236
R18818 XThC.Tn[6].n8 XThC.Tn[6].t3 24.9236
R18819 XThC.Tn[6].n60 XThC.Tn[6].n2 18.5605
R18820 XThC.Tn[6].n60 XThC.Tn[6].n59 11.5205
R18821 XThC.Tn[6].n59 XThC.Tn[6].n58 3.18344
R18822 XThC.Tn[6].n58 XThC.Tn[6] 3.09179
R18823 XThC.Tn[6].n15 XThC.Tn[6] 0.931056
R18824 XThC.Tn[6].n18 XThC.Tn[6] 0.931056
R18825 XThC.Tn[6].n21 XThC.Tn[6] 0.931056
R18826 XThC.Tn[6].n24 XThC.Tn[6] 0.931056
R18827 XThC.Tn[6].n27 XThC.Tn[6] 0.931056
R18828 XThC.Tn[6].n30 XThC.Tn[6] 0.931056
R18829 XThC.Tn[6].n33 XThC.Tn[6] 0.931056
R18830 XThC.Tn[6].n36 XThC.Tn[6] 0.931056
R18831 XThC.Tn[6].n39 XThC.Tn[6] 0.931056
R18832 XThC.Tn[6].n42 XThC.Tn[6] 0.931056
R18833 XThC.Tn[6].n45 XThC.Tn[6] 0.931056
R18834 XThC.Tn[6].n48 XThC.Tn[6] 0.931056
R18835 XThC.Tn[6].n51 XThC.Tn[6] 0.931056
R18836 XThC.Tn[6].n54 XThC.Tn[6] 0.931056
R18837 XThC.Tn[6].n57 XThC.Tn[6] 0.931056
R18838 XThC.Tn[6] XThC.Tn[6].n60 0.6405
R18839 XThC.Tn[6] XThC.Tn[6].n12 0.396333
R18840 XThC.Tn[6] XThC.Tn[6].n15 0.396333
R18841 XThC.Tn[6] XThC.Tn[6].n18 0.396333
R18842 XThC.Tn[6] XThC.Tn[6].n21 0.396333
R18843 XThC.Tn[6] XThC.Tn[6].n24 0.396333
R18844 XThC.Tn[6] XThC.Tn[6].n27 0.396333
R18845 XThC.Tn[6] XThC.Tn[6].n30 0.396333
R18846 XThC.Tn[6] XThC.Tn[6].n33 0.396333
R18847 XThC.Tn[6] XThC.Tn[6].n36 0.396333
R18848 XThC.Tn[6] XThC.Tn[6].n39 0.396333
R18849 XThC.Tn[6] XThC.Tn[6].n42 0.396333
R18850 XThC.Tn[6] XThC.Tn[6].n45 0.396333
R18851 XThC.Tn[6] XThC.Tn[6].n48 0.396333
R18852 XThC.Tn[6] XThC.Tn[6].n51 0.396333
R18853 XThC.Tn[6] XThC.Tn[6].n54 0.396333
R18854 XThC.Tn[6] XThC.Tn[6].n57 0.396333
R18855 XThC.Tn[6].n11 XThC.Tn[6] 0.104667
R18856 XThC.Tn[6].n14 XThC.Tn[6] 0.104667
R18857 XThC.Tn[6].n17 XThC.Tn[6] 0.104667
R18858 XThC.Tn[6].n20 XThC.Tn[6] 0.104667
R18859 XThC.Tn[6].n23 XThC.Tn[6] 0.104667
R18860 XThC.Tn[6].n26 XThC.Tn[6] 0.104667
R18861 XThC.Tn[6].n29 XThC.Tn[6] 0.104667
R18862 XThC.Tn[6].n32 XThC.Tn[6] 0.104667
R18863 XThC.Tn[6].n35 XThC.Tn[6] 0.104667
R18864 XThC.Tn[6].n38 XThC.Tn[6] 0.104667
R18865 XThC.Tn[6].n41 XThC.Tn[6] 0.104667
R18866 XThC.Tn[6].n44 XThC.Tn[6] 0.104667
R18867 XThC.Tn[6].n47 XThC.Tn[6] 0.104667
R18868 XThC.Tn[6].n50 XThC.Tn[6] 0.104667
R18869 XThC.Tn[6].n53 XThC.Tn[6] 0.104667
R18870 XThC.Tn[6].n56 XThC.Tn[6] 0.104667
R18871 XThC.Tn[6].n11 XThC.Tn[6] 0.0309878
R18872 XThC.Tn[6].n14 XThC.Tn[6] 0.0309878
R18873 XThC.Tn[6].n17 XThC.Tn[6] 0.0309878
R18874 XThC.Tn[6].n20 XThC.Tn[6] 0.0309878
R18875 XThC.Tn[6].n23 XThC.Tn[6] 0.0309878
R18876 XThC.Tn[6].n26 XThC.Tn[6] 0.0309878
R18877 XThC.Tn[6].n29 XThC.Tn[6] 0.0309878
R18878 XThC.Tn[6].n32 XThC.Tn[6] 0.0309878
R18879 XThC.Tn[6].n35 XThC.Tn[6] 0.0309878
R18880 XThC.Tn[6].n38 XThC.Tn[6] 0.0309878
R18881 XThC.Tn[6].n41 XThC.Tn[6] 0.0309878
R18882 XThC.Tn[6].n44 XThC.Tn[6] 0.0309878
R18883 XThC.Tn[6].n47 XThC.Tn[6] 0.0309878
R18884 XThC.Tn[6].n50 XThC.Tn[6] 0.0309878
R18885 XThC.Tn[6].n53 XThC.Tn[6] 0.0309878
R18886 XThC.Tn[6].n56 XThC.Tn[6] 0.0309878
R18887 XThC.Tn[6].n12 XThC.Tn[6].n11 0.027939
R18888 XThC.Tn[6].n15 XThC.Tn[6].n14 0.027939
R18889 XThC.Tn[6].n18 XThC.Tn[6].n17 0.027939
R18890 XThC.Tn[6].n21 XThC.Tn[6].n20 0.027939
R18891 XThC.Tn[6].n24 XThC.Tn[6].n23 0.027939
R18892 XThC.Tn[6].n27 XThC.Tn[6].n26 0.027939
R18893 XThC.Tn[6].n30 XThC.Tn[6].n29 0.027939
R18894 XThC.Tn[6].n33 XThC.Tn[6].n32 0.027939
R18895 XThC.Tn[6].n36 XThC.Tn[6].n35 0.027939
R18896 XThC.Tn[6].n39 XThC.Tn[6].n38 0.027939
R18897 XThC.Tn[6].n42 XThC.Tn[6].n41 0.027939
R18898 XThC.Tn[6].n45 XThC.Tn[6].n44 0.027939
R18899 XThC.Tn[6].n48 XThC.Tn[6].n47 0.027939
R18900 XThC.Tn[6].n51 XThC.Tn[6].n50 0.027939
R18901 XThC.Tn[6].n54 XThC.Tn[6].n53 0.027939
R18902 XThC.Tn[6].n57 XThC.Tn[6].n56 0.027939
R18903 XThC.Tn[6].n58 XThC.Tn[6] 0.0140108
R18904 XThR.Tn[9].n8 XThR.Tn[9].n7 256.104
R18905 XThR.Tn[9].n5 XThR.Tn[9].n3 243.68
R18906 XThR.Tn[9].n2 XThR.Tn[9].n1 241.847
R18907 XThR.Tn[9].n5 XThR.Tn[9].n4 205.28
R18908 XThR.Tn[9].n8 XThR.Tn[9].n6 202.094
R18909 XThR.Tn[9].n2 XThR.Tn[9].n0 185
R18910 XThR.Tn[9] XThR.Tn[9].n82 161.363
R18911 XThR.Tn[9] XThR.Tn[9].n77 161.363
R18912 XThR.Tn[9] XThR.Tn[9].n72 161.363
R18913 XThR.Tn[9] XThR.Tn[9].n67 161.363
R18914 XThR.Tn[9] XThR.Tn[9].n62 161.363
R18915 XThR.Tn[9] XThR.Tn[9].n57 161.363
R18916 XThR.Tn[9] XThR.Tn[9].n52 161.363
R18917 XThR.Tn[9] XThR.Tn[9].n47 161.363
R18918 XThR.Tn[9] XThR.Tn[9].n42 161.363
R18919 XThR.Tn[9] XThR.Tn[9].n37 161.363
R18920 XThR.Tn[9] XThR.Tn[9].n32 161.363
R18921 XThR.Tn[9] XThR.Tn[9].n27 161.363
R18922 XThR.Tn[9] XThR.Tn[9].n22 161.363
R18923 XThR.Tn[9] XThR.Tn[9].n17 161.363
R18924 XThR.Tn[9] XThR.Tn[9].n12 161.363
R18925 XThR.Tn[9] XThR.Tn[9].n10 161.363
R18926 XThR.Tn[9].n84 XThR.Tn[9].n83 161.3
R18927 XThR.Tn[9].n79 XThR.Tn[9].n78 161.3
R18928 XThR.Tn[9].n74 XThR.Tn[9].n73 161.3
R18929 XThR.Tn[9].n69 XThR.Tn[9].n68 161.3
R18930 XThR.Tn[9].n64 XThR.Tn[9].n63 161.3
R18931 XThR.Tn[9].n59 XThR.Tn[9].n58 161.3
R18932 XThR.Tn[9].n54 XThR.Tn[9].n53 161.3
R18933 XThR.Tn[9].n49 XThR.Tn[9].n48 161.3
R18934 XThR.Tn[9].n44 XThR.Tn[9].n43 161.3
R18935 XThR.Tn[9].n39 XThR.Tn[9].n38 161.3
R18936 XThR.Tn[9].n34 XThR.Tn[9].n33 161.3
R18937 XThR.Tn[9].n29 XThR.Tn[9].n28 161.3
R18938 XThR.Tn[9].n24 XThR.Tn[9].n23 161.3
R18939 XThR.Tn[9].n19 XThR.Tn[9].n18 161.3
R18940 XThR.Tn[9].n14 XThR.Tn[9].n13 161.3
R18941 XThR.Tn[9].n82 XThR.Tn[9].t63 161.106
R18942 XThR.Tn[9].n77 XThR.Tn[9].t69 161.106
R18943 XThR.Tn[9].n72 XThR.Tn[9].t47 161.106
R18944 XThR.Tn[9].n67 XThR.Tn[9].t34 161.106
R18945 XThR.Tn[9].n62 XThR.Tn[9].t62 161.106
R18946 XThR.Tn[9].n57 XThR.Tn[9].t24 161.106
R18947 XThR.Tn[9].n52 XThR.Tn[9].t66 161.106
R18948 XThR.Tn[9].n47 XThR.Tn[9].t45 161.106
R18949 XThR.Tn[9].n42 XThR.Tn[9].t32 161.106
R18950 XThR.Tn[9].n37 XThR.Tn[9].t37 161.106
R18951 XThR.Tn[9].n32 XThR.Tn[9].t23 161.106
R18952 XThR.Tn[9].n27 XThR.Tn[9].t46 161.106
R18953 XThR.Tn[9].n22 XThR.Tn[9].t21 161.106
R18954 XThR.Tn[9].n17 XThR.Tn[9].t64 161.106
R18955 XThR.Tn[9].n12 XThR.Tn[9].t28 161.106
R18956 XThR.Tn[9].n10 XThR.Tn[9].t71 161.106
R18957 XThR.Tn[9].n83 XThR.Tn[9].t54 159.978
R18958 XThR.Tn[9].n78 XThR.Tn[9].t61 159.978
R18959 XThR.Tn[9].n73 XThR.Tn[9].t43 159.978
R18960 XThR.Tn[9].n68 XThR.Tn[9].t27 159.978
R18961 XThR.Tn[9].n63 XThR.Tn[9].t52 159.978
R18962 XThR.Tn[9].n58 XThR.Tn[9].t18 159.978
R18963 XThR.Tn[9].n53 XThR.Tn[9].t60 159.978
R18964 XThR.Tn[9].n48 XThR.Tn[9].t40 159.978
R18965 XThR.Tn[9].n43 XThR.Tn[9].t25 159.978
R18966 XThR.Tn[9].n38 XThR.Tn[9].t33 159.978
R18967 XThR.Tn[9].n33 XThR.Tn[9].t16 159.978
R18968 XThR.Tn[9].n28 XThR.Tn[9].t42 159.978
R18969 XThR.Tn[9].n23 XThR.Tn[9].t15 159.978
R18970 XThR.Tn[9].n18 XThR.Tn[9].t59 159.978
R18971 XThR.Tn[9].n13 XThR.Tn[9].t19 159.978
R18972 XThR.Tn[9].n82 XThR.Tn[9].t49 145.038
R18973 XThR.Tn[9].n77 XThR.Tn[9].t14 145.038
R18974 XThR.Tn[9].n72 XThR.Tn[9].t57 145.038
R18975 XThR.Tn[9].n67 XThR.Tn[9].t38 145.038
R18976 XThR.Tn[9].n62 XThR.Tn[9].t70 145.038
R18977 XThR.Tn[9].n57 XThR.Tn[9].t48 145.038
R18978 XThR.Tn[9].n52 XThR.Tn[9].t58 145.038
R18979 XThR.Tn[9].n47 XThR.Tn[9].t39 145.038
R18980 XThR.Tn[9].n42 XThR.Tn[9].t36 145.038
R18981 XThR.Tn[9].n37 XThR.Tn[9].t67 145.038
R18982 XThR.Tn[9].n32 XThR.Tn[9].t31 145.038
R18983 XThR.Tn[9].n27 XThR.Tn[9].t56 145.038
R18984 XThR.Tn[9].n22 XThR.Tn[9].t29 145.038
R18985 XThR.Tn[9].n17 XThR.Tn[9].t72 145.038
R18986 XThR.Tn[9].n12 XThR.Tn[9].t35 145.038
R18987 XThR.Tn[9].n10 XThR.Tn[9].t17 145.038
R18988 XThR.Tn[9].n83 XThR.Tn[9].t68 143.911
R18989 XThR.Tn[9].n78 XThR.Tn[9].t30 143.911
R18990 XThR.Tn[9].n73 XThR.Tn[9].t12 143.911
R18991 XThR.Tn[9].n68 XThR.Tn[9].t53 143.911
R18992 XThR.Tn[9].n63 XThR.Tn[9].t22 143.911
R18993 XThR.Tn[9].n58 XThR.Tn[9].t65 143.911
R18994 XThR.Tn[9].n53 XThR.Tn[9].t13 143.911
R18995 XThR.Tn[9].n48 XThR.Tn[9].t55 143.911
R18996 XThR.Tn[9].n43 XThR.Tn[9].t51 143.911
R18997 XThR.Tn[9].n38 XThR.Tn[9].t20 143.911
R18998 XThR.Tn[9].n33 XThR.Tn[9].t44 143.911
R18999 XThR.Tn[9].n28 XThR.Tn[9].t73 143.911
R19000 XThR.Tn[9].n23 XThR.Tn[9].t41 143.911
R19001 XThR.Tn[9].n18 XThR.Tn[9].t26 143.911
R19002 XThR.Tn[9].n13 XThR.Tn[9].t50 143.911
R19003 XThR.Tn[9] XThR.Tn[9].n5 35.7652
R19004 XThR.Tn[9].n6 XThR.Tn[9].t6 26.5955
R19005 XThR.Tn[9].n6 XThR.Tn[9].t4 26.5955
R19006 XThR.Tn[9].n7 XThR.Tn[9].t7 26.5955
R19007 XThR.Tn[9].n7 XThR.Tn[9].t5 26.5955
R19008 XThR.Tn[9].n3 XThR.Tn[9].t10 26.5955
R19009 XThR.Tn[9].n3 XThR.Tn[9].t8 26.5955
R19010 XThR.Tn[9].n4 XThR.Tn[9].t11 26.5955
R19011 XThR.Tn[9].n4 XThR.Tn[9].t9 26.5955
R19012 XThR.Tn[9].n0 XThR.Tn[9].t0 24.9236
R19013 XThR.Tn[9].n0 XThR.Tn[9].t2 24.9236
R19014 XThR.Tn[9].n1 XThR.Tn[9].t1 24.9236
R19015 XThR.Tn[9].n1 XThR.Tn[9].t3 24.9236
R19016 XThR.Tn[9] XThR.Tn[9].n2 22.9615
R19017 XThR.Tn[9].n9 XThR.Tn[9].n8 13.5534
R19018 XThR.Tn[9].n88 XThR.Tn[9] 7.97984
R19019 XThR.Tn[9] XThR.Tn[9].n11 5.4407
R19020 XThR.Tn[9].n16 XThR.Tn[9].n15 4.5005
R19021 XThR.Tn[9].n21 XThR.Tn[9].n20 4.5005
R19022 XThR.Tn[9].n26 XThR.Tn[9].n25 4.5005
R19023 XThR.Tn[9].n31 XThR.Tn[9].n30 4.5005
R19024 XThR.Tn[9].n36 XThR.Tn[9].n35 4.5005
R19025 XThR.Tn[9].n41 XThR.Tn[9].n40 4.5005
R19026 XThR.Tn[9].n46 XThR.Tn[9].n45 4.5005
R19027 XThR.Tn[9].n51 XThR.Tn[9].n50 4.5005
R19028 XThR.Tn[9].n56 XThR.Tn[9].n55 4.5005
R19029 XThR.Tn[9].n61 XThR.Tn[9].n60 4.5005
R19030 XThR.Tn[9].n66 XThR.Tn[9].n65 4.5005
R19031 XThR.Tn[9].n71 XThR.Tn[9].n70 4.5005
R19032 XThR.Tn[9].n76 XThR.Tn[9].n75 4.5005
R19033 XThR.Tn[9].n81 XThR.Tn[9].n80 4.5005
R19034 XThR.Tn[9].n86 XThR.Tn[9].n85 4.5005
R19035 XThR.Tn[9].n87 XThR.Tn[9] 3.70586
R19036 XThR.Tn[9].n88 XThR.Tn[9].n9 2.99115
R19037 XThR.Tn[9].n9 XThR.Tn[9] 2.87153
R19038 XThR.Tn[9].n16 XThR.Tn[9] 2.52282
R19039 XThR.Tn[9].n21 XThR.Tn[9] 2.52282
R19040 XThR.Tn[9].n26 XThR.Tn[9] 2.52282
R19041 XThR.Tn[9].n31 XThR.Tn[9] 2.52282
R19042 XThR.Tn[9].n36 XThR.Tn[9] 2.52282
R19043 XThR.Tn[9].n41 XThR.Tn[9] 2.52282
R19044 XThR.Tn[9].n46 XThR.Tn[9] 2.52282
R19045 XThR.Tn[9].n51 XThR.Tn[9] 2.52282
R19046 XThR.Tn[9].n56 XThR.Tn[9] 2.52282
R19047 XThR.Tn[9].n61 XThR.Tn[9] 2.52282
R19048 XThR.Tn[9].n66 XThR.Tn[9] 2.52282
R19049 XThR.Tn[9].n71 XThR.Tn[9] 2.52282
R19050 XThR.Tn[9].n76 XThR.Tn[9] 2.52282
R19051 XThR.Tn[9].n81 XThR.Tn[9] 2.52282
R19052 XThR.Tn[9].n86 XThR.Tn[9] 2.52282
R19053 XThR.Tn[9] XThR.Tn[9].n88 2.2734
R19054 XThR.Tn[9].n9 XThR.Tn[9] 1.50638
R19055 XThR.Tn[9].n84 XThR.Tn[9] 1.08677
R19056 XThR.Tn[9].n79 XThR.Tn[9] 1.08677
R19057 XThR.Tn[9].n74 XThR.Tn[9] 1.08677
R19058 XThR.Tn[9].n69 XThR.Tn[9] 1.08677
R19059 XThR.Tn[9].n64 XThR.Tn[9] 1.08677
R19060 XThR.Tn[9].n59 XThR.Tn[9] 1.08677
R19061 XThR.Tn[9].n54 XThR.Tn[9] 1.08677
R19062 XThR.Tn[9].n49 XThR.Tn[9] 1.08677
R19063 XThR.Tn[9].n44 XThR.Tn[9] 1.08677
R19064 XThR.Tn[9].n39 XThR.Tn[9] 1.08677
R19065 XThR.Tn[9].n34 XThR.Tn[9] 1.08677
R19066 XThR.Tn[9].n29 XThR.Tn[9] 1.08677
R19067 XThR.Tn[9].n24 XThR.Tn[9] 1.08677
R19068 XThR.Tn[9].n19 XThR.Tn[9] 1.08677
R19069 XThR.Tn[9].n14 XThR.Tn[9] 1.08677
R19070 XThR.Tn[9] XThR.Tn[9].n16 0.839786
R19071 XThR.Tn[9] XThR.Tn[9].n21 0.839786
R19072 XThR.Tn[9] XThR.Tn[9].n26 0.839786
R19073 XThR.Tn[9] XThR.Tn[9].n31 0.839786
R19074 XThR.Tn[9] XThR.Tn[9].n36 0.839786
R19075 XThR.Tn[9] XThR.Tn[9].n41 0.839786
R19076 XThR.Tn[9] XThR.Tn[9].n46 0.839786
R19077 XThR.Tn[9] XThR.Tn[9].n51 0.839786
R19078 XThR.Tn[9] XThR.Tn[9].n56 0.839786
R19079 XThR.Tn[9] XThR.Tn[9].n61 0.839786
R19080 XThR.Tn[9] XThR.Tn[9].n66 0.839786
R19081 XThR.Tn[9] XThR.Tn[9].n71 0.839786
R19082 XThR.Tn[9] XThR.Tn[9].n76 0.839786
R19083 XThR.Tn[9] XThR.Tn[9].n81 0.839786
R19084 XThR.Tn[9] XThR.Tn[9].n86 0.839786
R19085 XThR.Tn[9].n11 XThR.Tn[9] 0.499542
R19086 XThR.Tn[9].n85 XThR.Tn[9] 0.063
R19087 XThR.Tn[9].n80 XThR.Tn[9] 0.063
R19088 XThR.Tn[9].n75 XThR.Tn[9] 0.063
R19089 XThR.Tn[9].n70 XThR.Tn[9] 0.063
R19090 XThR.Tn[9].n65 XThR.Tn[9] 0.063
R19091 XThR.Tn[9].n60 XThR.Tn[9] 0.063
R19092 XThR.Tn[9].n55 XThR.Tn[9] 0.063
R19093 XThR.Tn[9].n50 XThR.Tn[9] 0.063
R19094 XThR.Tn[9].n45 XThR.Tn[9] 0.063
R19095 XThR.Tn[9].n40 XThR.Tn[9] 0.063
R19096 XThR.Tn[9].n35 XThR.Tn[9] 0.063
R19097 XThR.Tn[9].n30 XThR.Tn[9] 0.063
R19098 XThR.Tn[9].n25 XThR.Tn[9] 0.063
R19099 XThR.Tn[9].n20 XThR.Tn[9] 0.063
R19100 XThR.Tn[9].n15 XThR.Tn[9] 0.063
R19101 XThR.Tn[9].n87 XThR.Tn[9] 0.0540714
R19102 XThR.Tn[9] XThR.Tn[9].n87 0.038
R19103 XThR.Tn[9].n11 XThR.Tn[9] 0.0143889
R19104 XThR.Tn[9].n85 XThR.Tn[9].n84 0.00771154
R19105 XThR.Tn[9].n80 XThR.Tn[9].n79 0.00771154
R19106 XThR.Tn[9].n75 XThR.Tn[9].n74 0.00771154
R19107 XThR.Tn[9].n70 XThR.Tn[9].n69 0.00771154
R19108 XThR.Tn[9].n65 XThR.Tn[9].n64 0.00771154
R19109 XThR.Tn[9].n60 XThR.Tn[9].n59 0.00771154
R19110 XThR.Tn[9].n55 XThR.Tn[9].n54 0.00771154
R19111 XThR.Tn[9].n50 XThR.Tn[9].n49 0.00771154
R19112 XThR.Tn[9].n45 XThR.Tn[9].n44 0.00771154
R19113 XThR.Tn[9].n40 XThR.Tn[9].n39 0.00771154
R19114 XThR.Tn[9].n35 XThR.Tn[9].n34 0.00771154
R19115 XThR.Tn[9].n30 XThR.Tn[9].n29 0.00771154
R19116 XThR.Tn[9].n25 XThR.Tn[9].n24 0.00771154
R19117 XThR.Tn[9].n20 XThR.Tn[9].n19 0.00771154
R19118 XThR.Tn[9].n15 XThR.Tn[9].n14 0.00771154
R19119 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R19120 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R19121 XThC.Tn[5].n12 XThC.Tn[5].n10 161.406
R19122 XThC.Tn[5].n15 XThC.Tn[5].n13 161.406
R19123 XThC.Tn[5].n18 XThC.Tn[5].n16 161.406
R19124 XThC.Tn[5].n21 XThC.Tn[5].n19 161.406
R19125 XThC.Tn[5].n24 XThC.Tn[5].n22 161.406
R19126 XThC.Tn[5].n27 XThC.Tn[5].n25 161.406
R19127 XThC.Tn[5].n30 XThC.Tn[5].n28 161.406
R19128 XThC.Tn[5].n33 XThC.Tn[5].n31 161.406
R19129 XThC.Tn[5].n36 XThC.Tn[5].n34 161.406
R19130 XThC.Tn[5].n39 XThC.Tn[5].n37 161.406
R19131 XThC.Tn[5].n42 XThC.Tn[5].n40 161.406
R19132 XThC.Tn[5].n45 XThC.Tn[5].n43 161.406
R19133 XThC.Tn[5].n48 XThC.Tn[5].n46 161.406
R19134 XThC.Tn[5].n51 XThC.Tn[5].n49 161.406
R19135 XThC.Tn[5].n54 XThC.Tn[5].n52 161.406
R19136 XThC.Tn[5].n57 XThC.Tn[5].n55 161.406
R19137 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R19138 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R19139 XThC.Tn[5].n16 XThC.Tn[5].t23 161.202
R19140 XThC.Tn[5].n19 XThC.Tn[5].t24 161.202
R19141 XThC.Tn[5].n22 XThC.Tn[5].t13 161.202
R19142 XThC.Tn[5].n25 XThC.Tn[5].t14 161.202
R19143 XThC.Tn[5].n28 XThC.Tn[5].t27 161.202
R19144 XThC.Tn[5].n31 XThC.Tn[5].t35 161.202
R19145 XThC.Tn[5].n34 XThC.Tn[5].t37 161.202
R19146 XThC.Tn[5].n37 XThC.Tn[5].t25 161.202
R19147 XThC.Tn[5].n40 XThC.Tn[5].t26 161.202
R19148 XThC.Tn[5].n43 XThC.Tn[5].t39 161.202
R19149 XThC.Tn[5].n46 XThC.Tn[5].t16 161.202
R19150 XThC.Tn[5].n49 XThC.Tn[5].t18 161.202
R19151 XThC.Tn[5].n52 XThC.Tn[5].t30 161.202
R19152 XThC.Tn[5].n55 XThC.Tn[5].t41 161.202
R19153 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R19154 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R19155 XThC.Tn[5].n16 XThC.Tn[5].t36 145.137
R19156 XThC.Tn[5].n19 XThC.Tn[5].t38 145.137
R19157 XThC.Tn[5].n22 XThC.Tn[5].t28 145.137
R19158 XThC.Tn[5].n25 XThC.Tn[5].t29 145.137
R19159 XThC.Tn[5].n28 XThC.Tn[5].t43 145.137
R19160 XThC.Tn[5].n31 XThC.Tn[5].t17 145.137
R19161 XThC.Tn[5].n34 XThC.Tn[5].t20 145.137
R19162 XThC.Tn[5].n37 XThC.Tn[5].t40 145.137
R19163 XThC.Tn[5].n40 XThC.Tn[5].t42 145.137
R19164 XThC.Tn[5].n43 XThC.Tn[5].t21 145.137
R19165 XThC.Tn[5].n46 XThC.Tn[5].t31 145.137
R19166 XThC.Tn[5].n49 XThC.Tn[5].t32 145.137
R19167 XThC.Tn[5].n52 XThC.Tn[5].t12 145.137
R19168 XThC.Tn[5].n55 XThC.Tn[5].t22 145.137
R19169 XThC.Tn[5].n6 XThC.Tn[5].n4 135.249
R19170 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R19171 XThC.Tn[5].n6 XThC.Tn[5].n5 98.981
R19172 XThC.Tn[5].n8 XThC.Tn[5].n7 98.981
R19173 XThC.Tn[5].n8 XThC.Tn[5].n6 36.2672
R19174 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R19175 XThC.Tn[5].n59 XThC.Tn[5].n9 32.6405
R19176 XThC.Tn[5].n1 XThC.Tn[5].t5 26.5955
R19177 XThC.Tn[5].n1 XThC.Tn[5].t4 26.5955
R19178 XThC.Tn[5].n0 XThC.Tn[5].t7 26.5955
R19179 XThC.Tn[5].n0 XThC.Tn[5].t6 26.5955
R19180 XThC.Tn[5].n3 XThC.Tn[5].t1 24.9236
R19181 XThC.Tn[5].n3 XThC.Tn[5].t0 24.9236
R19182 XThC.Tn[5].n4 XThC.Tn[5].t8 24.9236
R19183 XThC.Tn[5].n4 XThC.Tn[5].t11 24.9236
R19184 XThC.Tn[5].n5 XThC.Tn[5].t10 24.9236
R19185 XThC.Tn[5].n5 XThC.Tn[5].t9 24.9236
R19186 XThC.Tn[5].n7 XThC.Tn[5].t3 24.9236
R19187 XThC.Tn[5].n7 XThC.Tn[5].t2 24.9236
R19188 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R19189 XThC.Tn[5] XThC.Tn[5].n59 6.7205
R19190 XThC.Tn[5].n58 XThC.Tn[5] 3.62266
R19191 XThC.Tn[5].n59 XThC.Tn[5].n58 3.18437
R19192 XThC.Tn[5].n15 XThC.Tn[5] 0.931056
R19193 XThC.Tn[5].n18 XThC.Tn[5] 0.931056
R19194 XThC.Tn[5].n21 XThC.Tn[5] 0.931056
R19195 XThC.Tn[5].n24 XThC.Tn[5] 0.931056
R19196 XThC.Tn[5].n27 XThC.Tn[5] 0.931056
R19197 XThC.Tn[5].n30 XThC.Tn[5] 0.931056
R19198 XThC.Tn[5].n33 XThC.Tn[5] 0.931056
R19199 XThC.Tn[5].n36 XThC.Tn[5] 0.931056
R19200 XThC.Tn[5].n39 XThC.Tn[5] 0.931056
R19201 XThC.Tn[5].n42 XThC.Tn[5] 0.931056
R19202 XThC.Tn[5].n45 XThC.Tn[5] 0.931056
R19203 XThC.Tn[5].n48 XThC.Tn[5] 0.931056
R19204 XThC.Tn[5].n51 XThC.Tn[5] 0.931056
R19205 XThC.Tn[5].n54 XThC.Tn[5] 0.931056
R19206 XThC.Tn[5].n57 XThC.Tn[5] 0.931056
R19207 XThC.Tn[5] XThC.Tn[5].n12 0.396333
R19208 XThC.Tn[5] XThC.Tn[5].n15 0.396333
R19209 XThC.Tn[5] XThC.Tn[5].n18 0.396333
R19210 XThC.Tn[5] XThC.Tn[5].n21 0.396333
R19211 XThC.Tn[5] XThC.Tn[5].n24 0.396333
R19212 XThC.Tn[5] XThC.Tn[5].n27 0.396333
R19213 XThC.Tn[5] XThC.Tn[5].n30 0.396333
R19214 XThC.Tn[5] XThC.Tn[5].n33 0.396333
R19215 XThC.Tn[5] XThC.Tn[5].n36 0.396333
R19216 XThC.Tn[5] XThC.Tn[5].n39 0.396333
R19217 XThC.Tn[5] XThC.Tn[5].n42 0.396333
R19218 XThC.Tn[5] XThC.Tn[5].n45 0.396333
R19219 XThC.Tn[5] XThC.Tn[5].n48 0.396333
R19220 XThC.Tn[5] XThC.Tn[5].n51 0.396333
R19221 XThC.Tn[5] XThC.Tn[5].n54 0.396333
R19222 XThC.Tn[5] XThC.Tn[5].n57 0.396333
R19223 XThC.Tn[5].n11 XThC.Tn[5] 0.104667
R19224 XThC.Tn[5].n14 XThC.Tn[5] 0.104667
R19225 XThC.Tn[5].n17 XThC.Tn[5] 0.104667
R19226 XThC.Tn[5].n20 XThC.Tn[5] 0.104667
R19227 XThC.Tn[5].n23 XThC.Tn[5] 0.104667
R19228 XThC.Tn[5].n26 XThC.Tn[5] 0.104667
R19229 XThC.Tn[5].n29 XThC.Tn[5] 0.104667
R19230 XThC.Tn[5].n32 XThC.Tn[5] 0.104667
R19231 XThC.Tn[5].n35 XThC.Tn[5] 0.104667
R19232 XThC.Tn[5].n38 XThC.Tn[5] 0.104667
R19233 XThC.Tn[5].n41 XThC.Tn[5] 0.104667
R19234 XThC.Tn[5].n44 XThC.Tn[5] 0.104667
R19235 XThC.Tn[5].n47 XThC.Tn[5] 0.104667
R19236 XThC.Tn[5].n50 XThC.Tn[5] 0.104667
R19237 XThC.Tn[5].n53 XThC.Tn[5] 0.104667
R19238 XThC.Tn[5].n56 XThC.Tn[5] 0.104667
R19239 XThC.Tn[5].n11 XThC.Tn[5] 0.0309878
R19240 XThC.Tn[5].n14 XThC.Tn[5] 0.0309878
R19241 XThC.Tn[5].n17 XThC.Tn[5] 0.0309878
R19242 XThC.Tn[5].n20 XThC.Tn[5] 0.0309878
R19243 XThC.Tn[5].n23 XThC.Tn[5] 0.0309878
R19244 XThC.Tn[5].n26 XThC.Tn[5] 0.0309878
R19245 XThC.Tn[5].n29 XThC.Tn[5] 0.0309878
R19246 XThC.Tn[5].n32 XThC.Tn[5] 0.0309878
R19247 XThC.Tn[5].n35 XThC.Tn[5] 0.0309878
R19248 XThC.Tn[5].n38 XThC.Tn[5] 0.0309878
R19249 XThC.Tn[5].n41 XThC.Tn[5] 0.0309878
R19250 XThC.Tn[5].n44 XThC.Tn[5] 0.0309878
R19251 XThC.Tn[5].n47 XThC.Tn[5] 0.0309878
R19252 XThC.Tn[5].n50 XThC.Tn[5] 0.0309878
R19253 XThC.Tn[5].n53 XThC.Tn[5] 0.0309878
R19254 XThC.Tn[5].n56 XThC.Tn[5] 0.0309878
R19255 XThC.Tn[5].n12 XThC.Tn[5].n11 0.027939
R19256 XThC.Tn[5].n15 XThC.Tn[5].n14 0.027939
R19257 XThC.Tn[5].n18 XThC.Tn[5].n17 0.027939
R19258 XThC.Tn[5].n21 XThC.Tn[5].n20 0.027939
R19259 XThC.Tn[5].n24 XThC.Tn[5].n23 0.027939
R19260 XThC.Tn[5].n27 XThC.Tn[5].n26 0.027939
R19261 XThC.Tn[5].n30 XThC.Tn[5].n29 0.027939
R19262 XThC.Tn[5].n33 XThC.Tn[5].n32 0.027939
R19263 XThC.Tn[5].n36 XThC.Tn[5].n35 0.027939
R19264 XThC.Tn[5].n39 XThC.Tn[5].n38 0.027939
R19265 XThC.Tn[5].n42 XThC.Tn[5].n41 0.027939
R19266 XThC.Tn[5].n45 XThC.Tn[5].n44 0.027939
R19267 XThC.Tn[5].n48 XThC.Tn[5].n47 0.027939
R19268 XThC.Tn[5].n51 XThC.Tn[5].n50 0.027939
R19269 XThC.Tn[5].n54 XThC.Tn[5].n53 0.027939
R19270 XThC.Tn[5].n57 XThC.Tn[5].n56 0.027939
R19271 XThC.Tn[5].n58 XThC.Tn[5] 0.0129681
R19272 XThC.Tn[9].n2 XThC.Tn[9].n1 265.341
R19273 XThC.Tn[9].n5 XThC.Tn[9].n3 243.68
R19274 XThC.Tn[9].n58 XThC.Tn[9].n56 241.847
R19275 XThC.Tn[9].n5 XThC.Tn[9].n4 205.28
R19276 XThC.Tn[9].n2 XThC.Tn[9].n0 202.094
R19277 XThC.Tn[9].n58 XThC.Tn[9].n57 185
R19278 XThC.Tn[9].n9 XThC.Tn[9].n7 161.406
R19279 XThC.Tn[9].n12 XThC.Tn[9].n10 161.406
R19280 XThC.Tn[9].n15 XThC.Tn[9].n13 161.406
R19281 XThC.Tn[9].n18 XThC.Tn[9].n16 161.406
R19282 XThC.Tn[9].n21 XThC.Tn[9].n19 161.406
R19283 XThC.Tn[9].n24 XThC.Tn[9].n22 161.406
R19284 XThC.Tn[9].n27 XThC.Tn[9].n25 161.406
R19285 XThC.Tn[9].n30 XThC.Tn[9].n28 161.406
R19286 XThC.Tn[9].n33 XThC.Tn[9].n31 161.406
R19287 XThC.Tn[9].n36 XThC.Tn[9].n34 161.406
R19288 XThC.Tn[9].n39 XThC.Tn[9].n37 161.406
R19289 XThC.Tn[9].n42 XThC.Tn[9].n40 161.406
R19290 XThC.Tn[9].n45 XThC.Tn[9].n43 161.406
R19291 XThC.Tn[9].n48 XThC.Tn[9].n46 161.406
R19292 XThC.Tn[9].n51 XThC.Tn[9].n49 161.406
R19293 XThC.Tn[9].n54 XThC.Tn[9].n52 161.406
R19294 XThC.Tn[9].n7 XThC.Tn[9].t12 161.202
R19295 XThC.Tn[9].n10 XThC.Tn[9].t30 161.202
R19296 XThC.Tn[9].n13 XThC.Tn[9].t34 161.202
R19297 XThC.Tn[9].n16 XThC.Tn[9].t35 161.202
R19298 XThC.Tn[9].n19 XThC.Tn[9].t24 161.202
R19299 XThC.Tn[9].n22 XThC.Tn[9].t25 161.202
R19300 XThC.Tn[9].n25 XThC.Tn[9].t38 161.202
R19301 XThC.Tn[9].n28 XThC.Tn[9].t14 161.202
R19302 XThC.Tn[9].n31 XThC.Tn[9].t16 161.202
R19303 XThC.Tn[9].n34 XThC.Tn[9].t36 161.202
R19304 XThC.Tn[9].n37 XThC.Tn[9].t37 161.202
R19305 XThC.Tn[9].n40 XThC.Tn[9].t18 161.202
R19306 XThC.Tn[9].n43 XThC.Tn[9].t27 161.202
R19307 XThC.Tn[9].n46 XThC.Tn[9].t29 161.202
R19308 XThC.Tn[9].n49 XThC.Tn[9].t41 161.202
R19309 XThC.Tn[9].n52 XThC.Tn[9].t20 161.202
R19310 XThC.Tn[9].n7 XThC.Tn[9].t26 145.137
R19311 XThC.Tn[9].n10 XThC.Tn[9].t13 145.137
R19312 XThC.Tn[9].n13 XThC.Tn[9].t15 145.137
R19313 XThC.Tn[9].n16 XThC.Tn[9].t17 145.137
R19314 XThC.Tn[9].n19 XThC.Tn[9].t39 145.137
R19315 XThC.Tn[9].n22 XThC.Tn[9].t40 145.137
R19316 XThC.Tn[9].n25 XThC.Tn[9].t22 145.137
R19317 XThC.Tn[9].n28 XThC.Tn[9].t28 145.137
R19318 XThC.Tn[9].n31 XThC.Tn[9].t31 145.137
R19319 XThC.Tn[9].n34 XThC.Tn[9].t19 145.137
R19320 XThC.Tn[9].n37 XThC.Tn[9].t21 145.137
R19321 XThC.Tn[9].n40 XThC.Tn[9].t32 145.137
R19322 XThC.Tn[9].n43 XThC.Tn[9].t42 145.137
R19323 XThC.Tn[9].n46 XThC.Tn[9].t43 145.137
R19324 XThC.Tn[9].n49 XThC.Tn[9].t23 145.137
R19325 XThC.Tn[9].n52 XThC.Tn[9].t33 145.137
R19326 XThC.Tn[9].n1 XThC.Tn[9].t6 26.5955
R19327 XThC.Tn[9].n1 XThC.Tn[9].t5 26.5955
R19328 XThC.Tn[9].n0 XThC.Tn[9].t4 26.5955
R19329 XThC.Tn[9].n0 XThC.Tn[9].t7 26.5955
R19330 XThC.Tn[9].n3 XThC.Tn[9].t9 26.5955
R19331 XThC.Tn[9].n3 XThC.Tn[9].t8 26.5955
R19332 XThC.Tn[9].n4 XThC.Tn[9].t11 26.5955
R19333 XThC.Tn[9].n4 XThC.Tn[9].t10 26.5955
R19334 XThC.Tn[9].n56 XThC.Tn[9].t1 24.9236
R19335 XThC.Tn[9].n56 XThC.Tn[9].t0 24.9236
R19336 XThC.Tn[9].n57 XThC.Tn[9].t2 24.9236
R19337 XThC.Tn[9].n57 XThC.Tn[9].t3 24.9236
R19338 XThC.Tn[9] XThC.Tn[9].n5 22.9652
R19339 XThC.Tn[9] XThC.Tn[9].n58 18.8943
R19340 XThC.Tn[9].n6 XThC.Tn[9].n2 13.9299
R19341 XThC.Tn[9].n6 XThC.Tn[9] 13.9299
R19342 XThC.Tn[9] XThC.Tn[9].n55 6.34069
R19343 XThC.Tn[9].n55 XThC.Tn[9] 5.13485
R19344 XThC.Tn[9].n55 XThC.Tn[9] 1.79489
R19345 XThC.Tn[9] XThC.Tn[9].n6 1.19676
R19346 XThC.Tn[9].n12 XThC.Tn[9] 0.931056
R19347 XThC.Tn[9].n15 XThC.Tn[9] 0.931056
R19348 XThC.Tn[9].n18 XThC.Tn[9] 0.931056
R19349 XThC.Tn[9].n21 XThC.Tn[9] 0.931056
R19350 XThC.Tn[9].n24 XThC.Tn[9] 0.931056
R19351 XThC.Tn[9].n27 XThC.Tn[9] 0.931056
R19352 XThC.Tn[9].n30 XThC.Tn[9] 0.931056
R19353 XThC.Tn[9].n33 XThC.Tn[9] 0.931056
R19354 XThC.Tn[9].n36 XThC.Tn[9] 0.931056
R19355 XThC.Tn[9].n39 XThC.Tn[9] 0.931056
R19356 XThC.Tn[9].n42 XThC.Tn[9] 0.931056
R19357 XThC.Tn[9].n45 XThC.Tn[9] 0.931056
R19358 XThC.Tn[9].n48 XThC.Tn[9] 0.931056
R19359 XThC.Tn[9].n51 XThC.Tn[9] 0.931056
R19360 XThC.Tn[9].n54 XThC.Tn[9] 0.931056
R19361 XThC.Tn[9] XThC.Tn[9].n9 0.396333
R19362 XThC.Tn[9] XThC.Tn[9].n12 0.396333
R19363 XThC.Tn[9] XThC.Tn[9].n15 0.396333
R19364 XThC.Tn[9] XThC.Tn[9].n18 0.396333
R19365 XThC.Tn[9] XThC.Tn[9].n21 0.396333
R19366 XThC.Tn[9] XThC.Tn[9].n24 0.396333
R19367 XThC.Tn[9] XThC.Tn[9].n27 0.396333
R19368 XThC.Tn[9] XThC.Tn[9].n30 0.396333
R19369 XThC.Tn[9] XThC.Tn[9].n33 0.396333
R19370 XThC.Tn[9] XThC.Tn[9].n36 0.396333
R19371 XThC.Tn[9] XThC.Tn[9].n39 0.396333
R19372 XThC.Tn[9] XThC.Tn[9].n42 0.396333
R19373 XThC.Tn[9] XThC.Tn[9].n45 0.396333
R19374 XThC.Tn[9] XThC.Tn[9].n48 0.396333
R19375 XThC.Tn[9] XThC.Tn[9].n51 0.396333
R19376 XThC.Tn[9] XThC.Tn[9].n54 0.396333
R19377 XThC.Tn[9].n8 XThC.Tn[9] 0.104667
R19378 XThC.Tn[9].n11 XThC.Tn[9] 0.104667
R19379 XThC.Tn[9].n14 XThC.Tn[9] 0.104667
R19380 XThC.Tn[9].n17 XThC.Tn[9] 0.104667
R19381 XThC.Tn[9].n20 XThC.Tn[9] 0.104667
R19382 XThC.Tn[9].n23 XThC.Tn[9] 0.104667
R19383 XThC.Tn[9].n26 XThC.Tn[9] 0.104667
R19384 XThC.Tn[9].n29 XThC.Tn[9] 0.104667
R19385 XThC.Tn[9].n32 XThC.Tn[9] 0.104667
R19386 XThC.Tn[9].n35 XThC.Tn[9] 0.104667
R19387 XThC.Tn[9].n38 XThC.Tn[9] 0.104667
R19388 XThC.Tn[9].n41 XThC.Tn[9] 0.104667
R19389 XThC.Tn[9].n44 XThC.Tn[9] 0.104667
R19390 XThC.Tn[9].n47 XThC.Tn[9] 0.104667
R19391 XThC.Tn[9].n50 XThC.Tn[9] 0.104667
R19392 XThC.Tn[9].n53 XThC.Tn[9] 0.104667
R19393 XThC.Tn[9].n8 XThC.Tn[9] 0.0309878
R19394 XThC.Tn[9].n11 XThC.Tn[9] 0.0309878
R19395 XThC.Tn[9].n14 XThC.Tn[9] 0.0309878
R19396 XThC.Tn[9].n17 XThC.Tn[9] 0.0309878
R19397 XThC.Tn[9].n20 XThC.Tn[9] 0.0309878
R19398 XThC.Tn[9].n23 XThC.Tn[9] 0.0309878
R19399 XThC.Tn[9].n26 XThC.Tn[9] 0.0309878
R19400 XThC.Tn[9].n29 XThC.Tn[9] 0.0309878
R19401 XThC.Tn[9].n32 XThC.Tn[9] 0.0309878
R19402 XThC.Tn[9].n35 XThC.Tn[9] 0.0309878
R19403 XThC.Tn[9].n38 XThC.Tn[9] 0.0309878
R19404 XThC.Tn[9].n41 XThC.Tn[9] 0.0309878
R19405 XThC.Tn[9].n44 XThC.Tn[9] 0.0309878
R19406 XThC.Tn[9].n47 XThC.Tn[9] 0.0309878
R19407 XThC.Tn[9].n50 XThC.Tn[9] 0.0309878
R19408 XThC.Tn[9].n53 XThC.Tn[9] 0.0309878
R19409 XThC.Tn[9].n9 XThC.Tn[9].n8 0.027939
R19410 XThC.Tn[9].n12 XThC.Tn[9].n11 0.027939
R19411 XThC.Tn[9].n15 XThC.Tn[9].n14 0.027939
R19412 XThC.Tn[9].n18 XThC.Tn[9].n17 0.027939
R19413 XThC.Tn[9].n21 XThC.Tn[9].n20 0.027939
R19414 XThC.Tn[9].n24 XThC.Tn[9].n23 0.027939
R19415 XThC.Tn[9].n27 XThC.Tn[9].n26 0.027939
R19416 XThC.Tn[9].n30 XThC.Tn[9].n29 0.027939
R19417 XThC.Tn[9].n33 XThC.Tn[9].n32 0.027939
R19418 XThC.Tn[9].n36 XThC.Tn[9].n35 0.027939
R19419 XThC.Tn[9].n39 XThC.Tn[9].n38 0.027939
R19420 XThC.Tn[9].n42 XThC.Tn[9].n41 0.027939
R19421 XThC.Tn[9].n45 XThC.Tn[9].n44 0.027939
R19422 XThC.Tn[9].n48 XThC.Tn[9].n47 0.027939
R19423 XThC.Tn[9].n51 XThC.Tn[9].n50 0.027939
R19424 XThC.Tn[9].n54 XThC.Tn[9].n53 0.027939
R19425 XThC.Tn[11].n54 XThC.Tn[11].n53 265.341
R19426 XThC.Tn[11].n58 XThC.Tn[11].n57 243.68
R19427 XThC.Tn[11].n2 XThC.Tn[11].n0 241.847
R19428 XThC.Tn[11].n58 XThC.Tn[11].n56 205.28
R19429 XThC.Tn[11].n54 XThC.Tn[11].n52 202.094
R19430 XThC.Tn[11].n2 XThC.Tn[11].n1 185
R19431 XThC.Tn[11].n5 XThC.Tn[11].n3 161.406
R19432 XThC.Tn[11].n8 XThC.Tn[11].n6 161.406
R19433 XThC.Tn[11].n11 XThC.Tn[11].n9 161.406
R19434 XThC.Tn[11].n14 XThC.Tn[11].n12 161.406
R19435 XThC.Tn[11].n17 XThC.Tn[11].n15 161.406
R19436 XThC.Tn[11].n20 XThC.Tn[11].n18 161.406
R19437 XThC.Tn[11].n23 XThC.Tn[11].n21 161.406
R19438 XThC.Tn[11].n26 XThC.Tn[11].n24 161.406
R19439 XThC.Tn[11].n29 XThC.Tn[11].n27 161.406
R19440 XThC.Tn[11].n32 XThC.Tn[11].n30 161.406
R19441 XThC.Tn[11].n35 XThC.Tn[11].n33 161.406
R19442 XThC.Tn[11].n38 XThC.Tn[11].n36 161.406
R19443 XThC.Tn[11].n41 XThC.Tn[11].n39 161.406
R19444 XThC.Tn[11].n44 XThC.Tn[11].n42 161.406
R19445 XThC.Tn[11].n47 XThC.Tn[11].n45 161.406
R19446 XThC.Tn[11].n50 XThC.Tn[11].n48 161.406
R19447 XThC.Tn[11].n3 XThC.Tn[11].t18 161.202
R19448 XThC.Tn[11].n6 XThC.Tn[11].t35 161.202
R19449 XThC.Tn[11].n9 XThC.Tn[11].t37 161.202
R19450 XThC.Tn[11].n12 XThC.Tn[11].t39 161.202
R19451 XThC.Tn[11].n15 XThC.Tn[11].t28 161.202
R19452 XThC.Tn[11].n18 XThC.Tn[11].t29 161.202
R19453 XThC.Tn[11].n21 XThC.Tn[11].t42 161.202
R19454 XThC.Tn[11].n24 XThC.Tn[11].t19 161.202
R19455 XThC.Tn[11].n27 XThC.Tn[11].t21 161.202
R19456 XThC.Tn[11].n30 XThC.Tn[11].t40 161.202
R19457 XThC.Tn[11].n33 XThC.Tn[11].t41 161.202
R19458 XThC.Tn[11].n36 XThC.Tn[11].t22 161.202
R19459 XThC.Tn[11].n39 XThC.Tn[11].t30 161.202
R19460 XThC.Tn[11].n42 XThC.Tn[11].t33 161.202
R19461 XThC.Tn[11].n45 XThC.Tn[11].t14 161.202
R19462 XThC.Tn[11].n48 XThC.Tn[11].t24 161.202
R19463 XThC.Tn[11].n3 XThC.Tn[11].t20 145.137
R19464 XThC.Tn[11].n6 XThC.Tn[11].t38 145.137
R19465 XThC.Tn[11].n9 XThC.Tn[11].t43 145.137
R19466 XThC.Tn[11].n12 XThC.Tn[11].t12 145.137
R19467 XThC.Tn[11].n15 XThC.Tn[11].t31 145.137
R19468 XThC.Tn[11].n18 XThC.Tn[11].t32 145.137
R19469 XThC.Tn[11].n21 XThC.Tn[11].t16 145.137
R19470 XThC.Tn[11].n24 XThC.Tn[11].t23 145.137
R19471 XThC.Tn[11].n27 XThC.Tn[11].t25 145.137
R19472 XThC.Tn[11].n30 XThC.Tn[11].t13 145.137
R19473 XThC.Tn[11].n33 XThC.Tn[11].t15 145.137
R19474 XThC.Tn[11].n36 XThC.Tn[11].t26 145.137
R19475 XThC.Tn[11].n39 XThC.Tn[11].t34 145.137
R19476 XThC.Tn[11].n42 XThC.Tn[11].t36 145.137
R19477 XThC.Tn[11].n45 XThC.Tn[11].t17 145.137
R19478 XThC.Tn[11].n48 XThC.Tn[11].t27 145.137
R19479 XThC.Tn[11].n53 XThC.Tn[11].t5 26.5955
R19480 XThC.Tn[11].n53 XThC.Tn[11].t7 26.5955
R19481 XThC.Tn[11].n52 XThC.Tn[11].t11 26.5955
R19482 XThC.Tn[11].n52 XThC.Tn[11].t8 26.5955
R19483 XThC.Tn[11].n56 XThC.Tn[11].t2 26.5955
R19484 XThC.Tn[11].n56 XThC.Tn[11].t1 26.5955
R19485 XThC.Tn[11].n57 XThC.Tn[11].t0 26.5955
R19486 XThC.Tn[11].n57 XThC.Tn[11].t3 26.5955
R19487 XThC.Tn[11].n1 XThC.Tn[11].t4 24.9236
R19488 XThC.Tn[11].n1 XThC.Tn[11].t10 24.9236
R19489 XThC.Tn[11].n0 XThC.Tn[11].t6 24.9236
R19490 XThC.Tn[11].n0 XThC.Tn[11].t9 24.9236
R19491 XThC.Tn[11] XThC.Tn[11].n58 22.9652
R19492 XThC.Tn[11] XThC.Tn[11].n2 18.8943
R19493 XThC.Tn[11].n55 XThC.Tn[11].n54 13.9299
R19494 XThC.Tn[11] XThC.Tn[11].n55 13.9299
R19495 XThC.Tn[11].n51 XThC.Tn[11] 6.34069
R19496 XThC.Tn[11].n51 XThC.Tn[11] 5.13485
R19497 XThC.Tn[11] XThC.Tn[11].n51 1.79489
R19498 XThC.Tn[11].n55 XThC.Tn[11] 1.19676
R19499 XThC.Tn[11].n8 XThC.Tn[11] 0.931056
R19500 XThC.Tn[11].n11 XThC.Tn[11] 0.931056
R19501 XThC.Tn[11].n14 XThC.Tn[11] 0.931056
R19502 XThC.Tn[11].n17 XThC.Tn[11] 0.931056
R19503 XThC.Tn[11].n20 XThC.Tn[11] 0.931056
R19504 XThC.Tn[11].n23 XThC.Tn[11] 0.931056
R19505 XThC.Tn[11].n26 XThC.Tn[11] 0.931056
R19506 XThC.Tn[11].n29 XThC.Tn[11] 0.931056
R19507 XThC.Tn[11].n32 XThC.Tn[11] 0.931056
R19508 XThC.Tn[11].n35 XThC.Tn[11] 0.931056
R19509 XThC.Tn[11].n38 XThC.Tn[11] 0.931056
R19510 XThC.Tn[11].n41 XThC.Tn[11] 0.931056
R19511 XThC.Tn[11].n44 XThC.Tn[11] 0.931056
R19512 XThC.Tn[11].n47 XThC.Tn[11] 0.931056
R19513 XThC.Tn[11].n50 XThC.Tn[11] 0.931056
R19514 XThC.Tn[11] XThC.Tn[11].n5 0.396333
R19515 XThC.Tn[11] XThC.Tn[11].n8 0.396333
R19516 XThC.Tn[11] XThC.Tn[11].n11 0.396333
R19517 XThC.Tn[11] XThC.Tn[11].n14 0.396333
R19518 XThC.Tn[11] XThC.Tn[11].n17 0.396333
R19519 XThC.Tn[11] XThC.Tn[11].n20 0.396333
R19520 XThC.Tn[11] XThC.Tn[11].n23 0.396333
R19521 XThC.Tn[11] XThC.Tn[11].n26 0.396333
R19522 XThC.Tn[11] XThC.Tn[11].n29 0.396333
R19523 XThC.Tn[11] XThC.Tn[11].n32 0.396333
R19524 XThC.Tn[11] XThC.Tn[11].n35 0.396333
R19525 XThC.Tn[11] XThC.Tn[11].n38 0.396333
R19526 XThC.Tn[11] XThC.Tn[11].n41 0.396333
R19527 XThC.Tn[11] XThC.Tn[11].n44 0.396333
R19528 XThC.Tn[11] XThC.Tn[11].n47 0.396333
R19529 XThC.Tn[11] XThC.Tn[11].n50 0.396333
R19530 XThC.Tn[11].n4 XThC.Tn[11] 0.104667
R19531 XThC.Tn[11].n7 XThC.Tn[11] 0.104667
R19532 XThC.Tn[11].n10 XThC.Tn[11] 0.104667
R19533 XThC.Tn[11].n13 XThC.Tn[11] 0.104667
R19534 XThC.Tn[11].n16 XThC.Tn[11] 0.104667
R19535 XThC.Tn[11].n19 XThC.Tn[11] 0.104667
R19536 XThC.Tn[11].n22 XThC.Tn[11] 0.104667
R19537 XThC.Tn[11].n25 XThC.Tn[11] 0.104667
R19538 XThC.Tn[11].n28 XThC.Tn[11] 0.104667
R19539 XThC.Tn[11].n31 XThC.Tn[11] 0.104667
R19540 XThC.Tn[11].n34 XThC.Tn[11] 0.104667
R19541 XThC.Tn[11].n37 XThC.Tn[11] 0.104667
R19542 XThC.Tn[11].n40 XThC.Tn[11] 0.104667
R19543 XThC.Tn[11].n43 XThC.Tn[11] 0.104667
R19544 XThC.Tn[11].n46 XThC.Tn[11] 0.104667
R19545 XThC.Tn[11].n49 XThC.Tn[11] 0.104667
R19546 XThC.Tn[11].n4 XThC.Tn[11] 0.0309878
R19547 XThC.Tn[11].n7 XThC.Tn[11] 0.0309878
R19548 XThC.Tn[11].n10 XThC.Tn[11] 0.0309878
R19549 XThC.Tn[11].n13 XThC.Tn[11] 0.0309878
R19550 XThC.Tn[11].n16 XThC.Tn[11] 0.0309878
R19551 XThC.Tn[11].n19 XThC.Tn[11] 0.0309878
R19552 XThC.Tn[11].n22 XThC.Tn[11] 0.0309878
R19553 XThC.Tn[11].n25 XThC.Tn[11] 0.0309878
R19554 XThC.Tn[11].n28 XThC.Tn[11] 0.0309878
R19555 XThC.Tn[11].n31 XThC.Tn[11] 0.0309878
R19556 XThC.Tn[11].n34 XThC.Tn[11] 0.0309878
R19557 XThC.Tn[11].n37 XThC.Tn[11] 0.0309878
R19558 XThC.Tn[11].n40 XThC.Tn[11] 0.0309878
R19559 XThC.Tn[11].n43 XThC.Tn[11] 0.0309878
R19560 XThC.Tn[11].n46 XThC.Tn[11] 0.0309878
R19561 XThC.Tn[11].n49 XThC.Tn[11] 0.0309878
R19562 XThC.Tn[11].n5 XThC.Tn[11].n4 0.027939
R19563 XThC.Tn[11].n8 XThC.Tn[11].n7 0.027939
R19564 XThC.Tn[11].n11 XThC.Tn[11].n10 0.027939
R19565 XThC.Tn[11].n14 XThC.Tn[11].n13 0.027939
R19566 XThC.Tn[11].n17 XThC.Tn[11].n16 0.027939
R19567 XThC.Tn[11].n20 XThC.Tn[11].n19 0.027939
R19568 XThC.Tn[11].n23 XThC.Tn[11].n22 0.027939
R19569 XThC.Tn[11].n26 XThC.Tn[11].n25 0.027939
R19570 XThC.Tn[11].n29 XThC.Tn[11].n28 0.027939
R19571 XThC.Tn[11].n32 XThC.Tn[11].n31 0.027939
R19572 XThC.Tn[11].n35 XThC.Tn[11].n34 0.027939
R19573 XThC.Tn[11].n38 XThC.Tn[11].n37 0.027939
R19574 XThC.Tn[11].n41 XThC.Tn[11].n40 0.027939
R19575 XThC.Tn[11].n44 XThC.Tn[11].n43 0.027939
R19576 XThC.Tn[11].n47 XThC.Tn[11].n46 0.027939
R19577 XThC.Tn[11].n50 XThC.Tn[11].n49 0.027939
R19578 XThC.Tn[12].n5 XThC.Tn[12].n4 256.104
R19579 XThC.Tn[12].n8 XThC.Tn[12].n6 243.68
R19580 XThC.Tn[12].n2 XThC.Tn[12].n1 241.847
R19581 XThC.Tn[12].n8 XThC.Tn[12].n7 205.28
R19582 XThC.Tn[12].n5 XThC.Tn[12].n3 202.095
R19583 XThC.Tn[12].n2 XThC.Tn[12].n0 185
R19584 XThC.Tn[12].n12 XThC.Tn[12].n10 161.406
R19585 XThC.Tn[12].n15 XThC.Tn[12].n13 161.406
R19586 XThC.Tn[12].n18 XThC.Tn[12].n16 161.406
R19587 XThC.Tn[12].n21 XThC.Tn[12].n19 161.406
R19588 XThC.Tn[12].n24 XThC.Tn[12].n22 161.406
R19589 XThC.Tn[12].n27 XThC.Tn[12].n25 161.406
R19590 XThC.Tn[12].n30 XThC.Tn[12].n28 161.406
R19591 XThC.Tn[12].n33 XThC.Tn[12].n31 161.406
R19592 XThC.Tn[12].n36 XThC.Tn[12].n34 161.406
R19593 XThC.Tn[12].n39 XThC.Tn[12].n37 161.406
R19594 XThC.Tn[12].n42 XThC.Tn[12].n40 161.406
R19595 XThC.Tn[12].n45 XThC.Tn[12].n43 161.406
R19596 XThC.Tn[12].n48 XThC.Tn[12].n46 161.406
R19597 XThC.Tn[12].n51 XThC.Tn[12].n49 161.406
R19598 XThC.Tn[12].n54 XThC.Tn[12].n52 161.406
R19599 XThC.Tn[12].n57 XThC.Tn[12].n55 161.406
R19600 XThC.Tn[12].n10 XThC.Tn[12].t35 161.202
R19601 XThC.Tn[12].n13 XThC.Tn[12].t20 161.202
R19602 XThC.Tn[12].n16 XThC.Tn[12].t22 161.202
R19603 XThC.Tn[12].n19 XThC.Tn[12].t24 161.202
R19604 XThC.Tn[12].n22 XThC.Tn[12].t13 161.202
R19605 XThC.Tn[12].n25 XThC.Tn[12].t14 161.202
R19606 XThC.Tn[12].n28 XThC.Tn[12].t27 161.202
R19607 XThC.Tn[12].n31 XThC.Tn[12].t36 161.202
R19608 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R19609 XThC.Tn[12].n37 XThC.Tn[12].t25 161.202
R19610 XThC.Tn[12].n40 XThC.Tn[12].t26 161.202
R19611 XThC.Tn[12].n43 XThC.Tn[12].t39 161.202
R19612 XThC.Tn[12].n46 XThC.Tn[12].t15 161.202
R19613 XThC.Tn[12].n49 XThC.Tn[12].t18 161.202
R19614 XThC.Tn[12].n52 XThC.Tn[12].t31 161.202
R19615 XThC.Tn[12].n55 XThC.Tn[12].t41 161.202
R19616 XThC.Tn[12].n10 XThC.Tn[12].t37 145.137
R19617 XThC.Tn[12].n13 XThC.Tn[12].t23 145.137
R19618 XThC.Tn[12].n16 XThC.Tn[12].t28 145.137
R19619 XThC.Tn[12].n19 XThC.Tn[12].t29 145.137
R19620 XThC.Tn[12].n22 XThC.Tn[12].t16 145.137
R19621 XThC.Tn[12].n25 XThC.Tn[12].t17 145.137
R19622 XThC.Tn[12].n28 XThC.Tn[12].t33 145.137
R19623 XThC.Tn[12].n31 XThC.Tn[12].t40 145.137
R19624 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R19625 XThC.Tn[12].n37 XThC.Tn[12].t30 145.137
R19626 XThC.Tn[12].n40 XThC.Tn[12].t32 145.137
R19627 XThC.Tn[12].n43 XThC.Tn[12].t43 145.137
R19628 XThC.Tn[12].n46 XThC.Tn[12].t19 145.137
R19629 XThC.Tn[12].n49 XThC.Tn[12].t21 145.137
R19630 XThC.Tn[12].n52 XThC.Tn[12].t34 145.137
R19631 XThC.Tn[12].n55 XThC.Tn[12].t12 145.137
R19632 XThC.Tn[12].n3 XThC.Tn[12].t5 26.5955
R19633 XThC.Tn[12].n3 XThC.Tn[12].t6 26.5955
R19634 XThC.Tn[12].n4 XThC.Tn[12].t4 26.5955
R19635 XThC.Tn[12].n4 XThC.Tn[12].t7 26.5955
R19636 XThC.Tn[12].n6 XThC.Tn[12].t9 26.5955
R19637 XThC.Tn[12].n6 XThC.Tn[12].t8 26.5955
R19638 XThC.Tn[12].n7 XThC.Tn[12].t11 26.5955
R19639 XThC.Tn[12].n7 XThC.Tn[12].t10 26.5955
R19640 XThC.Tn[12].n0 XThC.Tn[12].t1 24.9236
R19641 XThC.Tn[12].n0 XThC.Tn[12].t0 24.9236
R19642 XThC.Tn[12].n1 XThC.Tn[12].t3 24.9236
R19643 XThC.Tn[12].n1 XThC.Tn[12].t2 24.9236
R19644 XThC.Tn[12] XThC.Tn[12].n8 22.9652
R19645 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R19646 XThC.Tn[12].n9 XThC.Tn[12].n5 13.9299
R19647 XThC.Tn[12].n9 XThC.Tn[12] 13.9299
R19648 XThC.Tn[12].n59 XThC.Tn[12].n58 5.13244
R19649 XThC.Tn[12].n58 XThC.Tn[12] 3.8444
R19650 XThC.Tn[12].n59 XThC.Tn[12].n9 2.99115
R19651 XThC.Tn[12].n9 XThC.Tn[12] 2.87153
R19652 XThC.Tn[12] XThC.Tn[12].n59 2.2734
R19653 XThC.Tn[12].n15 XThC.Tn[12] 0.931056
R19654 XThC.Tn[12].n18 XThC.Tn[12] 0.931056
R19655 XThC.Tn[12].n21 XThC.Tn[12] 0.931056
R19656 XThC.Tn[12].n24 XThC.Tn[12] 0.931056
R19657 XThC.Tn[12].n27 XThC.Tn[12] 0.931056
R19658 XThC.Tn[12].n30 XThC.Tn[12] 0.931056
R19659 XThC.Tn[12].n33 XThC.Tn[12] 0.931056
R19660 XThC.Tn[12].n36 XThC.Tn[12] 0.931056
R19661 XThC.Tn[12].n39 XThC.Tn[12] 0.931056
R19662 XThC.Tn[12].n42 XThC.Tn[12] 0.931056
R19663 XThC.Tn[12].n45 XThC.Tn[12] 0.931056
R19664 XThC.Tn[12].n48 XThC.Tn[12] 0.931056
R19665 XThC.Tn[12].n51 XThC.Tn[12] 0.931056
R19666 XThC.Tn[12].n54 XThC.Tn[12] 0.931056
R19667 XThC.Tn[12].n57 XThC.Tn[12] 0.931056
R19668 XThC.Tn[12] XThC.Tn[12].n12 0.396333
R19669 XThC.Tn[12] XThC.Tn[12].n15 0.396333
R19670 XThC.Tn[12] XThC.Tn[12].n18 0.396333
R19671 XThC.Tn[12] XThC.Tn[12].n21 0.396333
R19672 XThC.Tn[12] XThC.Tn[12].n24 0.396333
R19673 XThC.Tn[12] XThC.Tn[12].n27 0.396333
R19674 XThC.Tn[12] XThC.Tn[12].n30 0.396333
R19675 XThC.Tn[12] XThC.Tn[12].n33 0.396333
R19676 XThC.Tn[12] XThC.Tn[12].n36 0.396333
R19677 XThC.Tn[12] XThC.Tn[12].n39 0.396333
R19678 XThC.Tn[12] XThC.Tn[12].n42 0.396333
R19679 XThC.Tn[12] XThC.Tn[12].n45 0.396333
R19680 XThC.Tn[12] XThC.Tn[12].n48 0.396333
R19681 XThC.Tn[12] XThC.Tn[12].n51 0.396333
R19682 XThC.Tn[12] XThC.Tn[12].n54 0.396333
R19683 XThC.Tn[12] XThC.Tn[12].n57 0.396333
R19684 XThC.Tn[12].n11 XThC.Tn[12] 0.104667
R19685 XThC.Tn[12].n14 XThC.Tn[12] 0.104667
R19686 XThC.Tn[12].n17 XThC.Tn[12] 0.104667
R19687 XThC.Tn[12].n20 XThC.Tn[12] 0.104667
R19688 XThC.Tn[12].n23 XThC.Tn[12] 0.104667
R19689 XThC.Tn[12].n26 XThC.Tn[12] 0.104667
R19690 XThC.Tn[12].n29 XThC.Tn[12] 0.104667
R19691 XThC.Tn[12].n32 XThC.Tn[12] 0.104667
R19692 XThC.Tn[12].n35 XThC.Tn[12] 0.104667
R19693 XThC.Tn[12].n38 XThC.Tn[12] 0.104667
R19694 XThC.Tn[12].n41 XThC.Tn[12] 0.104667
R19695 XThC.Tn[12].n44 XThC.Tn[12] 0.104667
R19696 XThC.Tn[12].n47 XThC.Tn[12] 0.104667
R19697 XThC.Tn[12].n50 XThC.Tn[12] 0.104667
R19698 XThC.Tn[12].n53 XThC.Tn[12] 0.104667
R19699 XThC.Tn[12].n56 XThC.Tn[12] 0.104667
R19700 XThC.Tn[12].n11 XThC.Tn[12] 0.0309878
R19701 XThC.Tn[12].n14 XThC.Tn[12] 0.0309878
R19702 XThC.Tn[12].n17 XThC.Tn[12] 0.0309878
R19703 XThC.Tn[12].n20 XThC.Tn[12] 0.0309878
R19704 XThC.Tn[12].n23 XThC.Tn[12] 0.0309878
R19705 XThC.Tn[12].n26 XThC.Tn[12] 0.0309878
R19706 XThC.Tn[12].n29 XThC.Tn[12] 0.0309878
R19707 XThC.Tn[12].n32 XThC.Tn[12] 0.0309878
R19708 XThC.Tn[12].n35 XThC.Tn[12] 0.0309878
R19709 XThC.Tn[12].n38 XThC.Tn[12] 0.0309878
R19710 XThC.Tn[12].n41 XThC.Tn[12] 0.0309878
R19711 XThC.Tn[12].n44 XThC.Tn[12] 0.0309878
R19712 XThC.Tn[12].n47 XThC.Tn[12] 0.0309878
R19713 XThC.Tn[12].n50 XThC.Tn[12] 0.0309878
R19714 XThC.Tn[12].n53 XThC.Tn[12] 0.0309878
R19715 XThC.Tn[12].n56 XThC.Tn[12] 0.0309878
R19716 XThC.Tn[12].n12 XThC.Tn[12].n11 0.027939
R19717 XThC.Tn[12].n15 XThC.Tn[12].n14 0.027939
R19718 XThC.Tn[12].n18 XThC.Tn[12].n17 0.027939
R19719 XThC.Tn[12].n21 XThC.Tn[12].n20 0.027939
R19720 XThC.Tn[12].n24 XThC.Tn[12].n23 0.027939
R19721 XThC.Tn[12].n27 XThC.Tn[12].n26 0.027939
R19722 XThC.Tn[12].n30 XThC.Tn[12].n29 0.027939
R19723 XThC.Tn[12].n33 XThC.Tn[12].n32 0.027939
R19724 XThC.Tn[12].n36 XThC.Tn[12].n35 0.027939
R19725 XThC.Tn[12].n39 XThC.Tn[12].n38 0.027939
R19726 XThC.Tn[12].n42 XThC.Tn[12].n41 0.027939
R19727 XThC.Tn[12].n45 XThC.Tn[12].n44 0.027939
R19728 XThC.Tn[12].n48 XThC.Tn[12].n47 0.027939
R19729 XThC.Tn[12].n51 XThC.Tn[12].n50 0.027939
R19730 XThC.Tn[12].n54 XThC.Tn[12].n53 0.027939
R19731 XThC.Tn[12].n57 XThC.Tn[12].n56 0.027939
R19732 XThC.Tn[12].n58 XThC.Tn[12] 0.00316553
R19733 XThC.Tn[13].n55 XThC.Tn[13].n54 265.341
R19734 XThC.Tn[13].n59 XThC.Tn[13].n57 243.68
R19735 XThC.Tn[13].n2 XThC.Tn[13].n0 241.847
R19736 XThC.Tn[13].n59 XThC.Tn[13].n58 205.28
R19737 XThC.Tn[13].n55 XThC.Tn[13].n53 202.094
R19738 XThC.Tn[13].n2 XThC.Tn[13].n1 185
R19739 XThC.Tn[13].n5 XThC.Tn[13].n3 161.406
R19740 XThC.Tn[13].n8 XThC.Tn[13].n6 161.406
R19741 XThC.Tn[13].n11 XThC.Tn[13].n9 161.406
R19742 XThC.Tn[13].n14 XThC.Tn[13].n12 161.406
R19743 XThC.Tn[13].n17 XThC.Tn[13].n15 161.406
R19744 XThC.Tn[13].n20 XThC.Tn[13].n18 161.406
R19745 XThC.Tn[13].n23 XThC.Tn[13].n21 161.406
R19746 XThC.Tn[13].n26 XThC.Tn[13].n24 161.406
R19747 XThC.Tn[13].n29 XThC.Tn[13].n27 161.406
R19748 XThC.Tn[13].n32 XThC.Tn[13].n30 161.406
R19749 XThC.Tn[13].n35 XThC.Tn[13].n33 161.406
R19750 XThC.Tn[13].n38 XThC.Tn[13].n36 161.406
R19751 XThC.Tn[13].n41 XThC.Tn[13].n39 161.406
R19752 XThC.Tn[13].n44 XThC.Tn[13].n42 161.406
R19753 XThC.Tn[13].n47 XThC.Tn[13].n45 161.406
R19754 XThC.Tn[13].n50 XThC.Tn[13].n48 161.406
R19755 XThC.Tn[13].n3 XThC.Tn[13].t27 161.202
R19756 XThC.Tn[13].n6 XThC.Tn[13].t12 161.202
R19757 XThC.Tn[13].n9 XThC.Tn[13].t14 161.202
R19758 XThC.Tn[13].n12 XThC.Tn[13].t16 161.202
R19759 XThC.Tn[13].n15 XThC.Tn[13].t37 161.202
R19760 XThC.Tn[13].n18 XThC.Tn[13].t38 161.202
R19761 XThC.Tn[13].n21 XThC.Tn[13].t19 161.202
R19762 XThC.Tn[13].n24 XThC.Tn[13].t28 161.202
R19763 XThC.Tn[13].n27 XThC.Tn[13].t30 161.202
R19764 XThC.Tn[13].n30 XThC.Tn[13].t17 161.202
R19765 XThC.Tn[13].n33 XThC.Tn[13].t18 161.202
R19766 XThC.Tn[13].n36 XThC.Tn[13].t31 161.202
R19767 XThC.Tn[13].n39 XThC.Tn[13].t39 161.202
R19768 XThC.Tn[13].n42 XThC.Tn[13].t42 161.202
R19769 XThC.Tn[13].n45 XThC.Tn[13].t23 161.202
R19770 XThC.Tn[13].n48 XThC.Tn[13].t33 161.202
R19771 XThC.Tn[13].n3 XThC.Tn[13].t29 145.137
R19772 XThC.Tn[13].n6 XThC.Tn[13].t15 145.137
R19773 XThC.Tn[13].n9 XThC.Tn[13].t20 145.137
R19774 XThC.Tn[13].n12 XThC.Tn[13].t21 145.137
R19775 XThC.Tn[13].n15 XThC.Tn[13].t40 145.137
R19776 XThC.Tn[13].n18 XThC.Tn[13].t41 145.137
R19777 XThC.Tn[13].n21 XThC.Tn[13].t25 145.137
R19778 XThC.Tn[13].n24 XThC.Tn[13].t32 145.137
R19779 XThC.Tn[13].n27 XThC.Tn[13].t34 145.137
R19780 XThC.Tn[13].n30 XThC.Tn[13].t22 145.137
R19781 XThC.Tn[13].n33 XThC.Tn[13].t24 145.137
R19782 XThC.Tn[13].n36 XThC.Tn[13].t35 145.137
R19783 XThC.Tn[13].n39 XThC.Tn[13].t43 145.137
R19784 XThC.Tn[13].n42 XThC.Tn[13].t13 145.137
R19785 XThC.Tn[13].n45 XThC.Tn[13].t26 145.137
R19786 XThC.Tn[13].n48 XThC.Tn[13].t36 145.137
R19787 XThC.Tn[13].n57 XThC.Tn[13].t1 26.5955
R19788 XThC.Tn[13].n57 XThC.Tn[13].t0 26.5955
R19789 XThC.Tn[13].n54 XThC.Tn[13].t8 26.5955
R19790 XThC.Tn[13].n54 XThC.Tn[13].t11 26.5955
R19791 XThC.Tn[13].n53 XThC.Tn[13].t10 26.5955
R19792 XThC.Tn[13].n53 XThC.Tn[13].t9 26.5955
R19793 XThC.Tn[13].n58 XThC.Tn[13].t3 26.5955
R19794 XThC.Tn[13].n58 XThC.Tn[13].t2 26.5955
R19795 XThC.Tn[13].n1 XThC.Tn[13].t4 24.9236
R19796 XThC.Tn[13].n1 XThC.Tn[13].t6 24.9236
R19797 XThC.Tn[13].n0 XThC.Tn[13].t7 24.9236
R19798 XThC.Tn[13].n0 XThC.Tn[13].t5 24.9236
R19799 XThC.Tn[13] XThC.Tn[13].n59 22.9652
R19800 XThC.Tn[13] XThC.Tn[13].n2 18.8943
R19801 XThC.Tn[13].n56 XThC.Tn[13].n55 13.9299
R19802 XThC.Tn[13] XThC.Tn[13].n56 13.9299
R19803 XThC.Tn[13].n52 XThC.Tn[13] 6.34069
R19804 XThC.Tn[13].n52 XThC.Tn[13].n51 5.13021
R19805 XThC.Tn[13].n51 XThC.Tn[13] 4.03795
R19806 XThC.Tn[13] XThC.Tn[13].n52 1.79489
R19807 XThC.Tn[13].n56 XThC.Tn[13] 1.19676
R19808 XThC.Tn[13].n8 XThC.Tn[13] 0.931056
R19809 XThC.Tn[13].n11 XThC.Tn[13] 0.931056
R19810 XThC.Tn[13].n14 XThC.Tn[13] 0.931056
R19811 XThC.Tn[13].n17 XThC.Tn[13] 0.931056
R19812 XThC.Tn[13].n20 XThC.Tn[13] 0.931056
R19813 XThC.Tn[13].n23 XThC.Tn[13] 0.931056
R19814 XThC.Tn[13].n26 XThC.Tn[13] 0.931056
R19815 XThC.Tn[13].n29 XThC.Tn[13] 0.931056
R19816 XThC.Tn[13].n32 XThC.Tn[13] 0.931056
R19817 XThC.Tn[13].n35 XThC.Tn[13] 0.931056
R19818 XThC.Tn[13].n38 XThC.Tn[13] 0.931056
R19819 XThC.Tn[13].n41 XThC.Tn[13] 0.931056
R19820 XThC.Tn[13].n44 XThC.Tn[13] 0.931056
R19821 XThC.Tn[13].n47 XThC.Tn[13] 0.931056
R19822 XThC.Tn[13].n50 XThC.Tn[13] 0.931056
R19823 XThC.Tn[13] XThC.Tn[13].n5 0.396333
R19824 XThC.Tn[13] XThC.Tn[13].n8 0.396333
R19825 XThC.Tn[13] XThC.Tn[13].n11 0.396333
R19826 XThC.Tn[13] XThC.Tn[13].n14 0.396333
R19827 XThC.Tn[13] XThC.Tn[13].n17 0.396333
R19828 XThC.Tn[13] XThC.Tn[13].n20 0.396333
R19829 XThC.Tn[13] XThC.Tn[13].n23 0.396333
R19830 XThC.Tn[13] XThC.Tn[13].n26 0.396333
R19831 XThC.Tn[13] XThC.Tn[13].n29 0.396333
R19832 XThC.Tn[13] XThC.Tn[13].n32 0.396333
R19833 XThC.Tn[13] XThC.Tn[13].n35 0.396333
R19834 XThC.Tn[13] XThC.Tn[13].n38 0.396333
R19835 XThC.Tn[13] XThC.Tn[13].n41 0.396333
R19836 XThC.Tn[13] XThC.Tn[13].n44 0.396333
R19837 XThC.Tn[13] XThC.Tn[13].n47 0.396333
R19838 XThC.Tn[13] XThC.Tn[13].n50 0.396333
R19839 XThC.Tn[13].n4 XThC.Tn[13] 0.104667
R19840 XThC.Tn[13].n7 XThC.Tn[13] 0.104667
R19841 XThC.Tn[13].n10 XThC.Tn[13] 0.104667
R19842 XThC.Tn[13].n13 XThC.Tn[13] 0.104667
R19843 XThC.Tn[13].n16 XThC.Tn[13] 0.104667
R19844 XThC.Tn[13].n19 XThC.Tn[13] 0.104667
R19845 XThC.Tn[13].n22 XThC.Tn[13] 0.104667
R19846 XThC.Tn[13].n25 XThC.Tn[13] 0.104667
R19847 XThC.Tn[13].n28 XThC.Tn[13] 0.104667
R19848 XThC.Tn[13].n31 XThC.Tn[13] 0.104667
R19849 XThC.Tn[13].n34 XThC.Tn[13] 0.104667
R19850 XThC.Tn[13].n37 XThC.Tn[13] 0.104667
R19851 XThC.Tn[13].n40 XThC.Tn[13] 0.104667
R19852 XThC.Tn[13].n43 XThC.Tn[13] 0.104667
R19853 XThC.Tn[13].n46 XThC.Tn[13] 0.104667
R19854 XThC.Tn[13].n49 XThC.Tn[13] 0.104667
R19855 XThC.Tn[13].n4 XThC.Tn[13] 0.0309878
R19856 XThC.Tn[13].n7 XThC.Tn[13] 0.0309878
R19857 XThC.Tn[13].n10 XThC.Tn[13] 0.0309878
R19858 XThC.Tn[13].n13 XThC.Tn[13] 0.0309878
R19859 XThC.Tn[13].n16 XThC.Tn[13] 0.0309878
R19860 XThC.Tn[13].n19 XThC.Tn[13] 0.0309878
R19861 XThC.Tn[13].n22 XThC.Tn[13] 0.0309878
R19862 XThC.Tn[13].n25 XThC.Tn[13] 0.0309878
R19863 XThC.Tn[13].n28 XThC.Tn[13] 0.0309878
R19864 XThC.Tn[13].n31 XThC.Tn[13] 0.0309878
R19865 XThC.Tn[13].n34 XThC.Tn[13] 0.0309878
R19866 XThC.Tn[13].n37 XThC.Tn[13] 0.0309878
R19867 XThC.Tn[13].n40 XThC.Tn[13] 0.0309878
R19868 XThC.Tn[13].n43 XThC.Tn[13] 0.0309878
R19869 XThC.Tn[13].n46 XThC.Tn[13] 0.0309878
R19870 XThC.Tn[13].n49 XThC.Tn[13] 0.0309878
R19871 XThC.Tn[13].n5 XThC.Tn[13].n4 0.027939
R19872 XThC.Tn[13].n8 XThC.Tn[13].n7 0.027939
R19873 XThC.Tn[13].n11 XThC.Tn[13].n10 0.027939
R19874 XThC.Tn[13].n14 XThC.Tn[13].n13 0.027939
R19875 XThC.Tn[13].n17 XThC.Tn[13].n16 0.027939
R19876 XThC.Tn[13].n20 XThC.Tn[13].n19 0.027939
R19877 XThC.Tn[13].n23 XThC.Tn[13].n22 0.027939
R19878 XThC.Tn[13].n26 XThC.Tn[13].n25 0.027939
R19879 XThC.Tn[13].n29 XThC.Tn[13].n28 0.027939
R19880 XThC.Tn[13].n32 XThC.Tn[13].n31 0.027939
R19881 XThC.Tn[13].n35 XThC.Tn[13].n34 0.027939
R19882 XThC.Tn[13].n38 XThC.Tn[13].n37 0.027939
R19883 XThC.Tn[13].n41 XThC.Tn[13].n40 0.027939
R19884 XThC.Tn[13].n44 XThC.Tn[13].n43 0.027939
R19885 XThC.Tn[13].n47 XThC.Tn[13].n46 0.027939
R19886 XThC.Tn[13].n50 XThC.Tn[13].n49 0.027939
R19887 XThC.Tn[13].n51 XThC.Tn[13] 0.00548355
R19888 XThC.Tn[0].n59 XThC.Tn[0].n58 332.332
R19889 XThC.Tn[0].n59 XThC.Tn[0].n57 296.493
R19890 XThC.Tn[0].n9 XThC.Tn[0].n7 161.406
R19891 XThC.Tn[0].n12 XThC.Tn[0].n10 161.406
R19892 XThC.Tn[0].n15 XThC.Tn[0].n13 161.406
R19893 XThC.Tn[0].n18 XThC.Tn[0].n16 161.406
R19894 XThC.Tn[0].n21 XThC.Tn[0].n19 161.406
R19895 XThC.Tn[0].n24 XThC.Tn[0].n22 161.406
R19896 XThC.Tn[0].n27 XThC.Tn[0].n25 161.406
R19897 XThC.Tn[0].n30 XThC.Tn[0].n28 161.406
R19898 XThC.Tn[0].n33 XThC.Tn[0].n31 161.406
R19899 XThC.Tn[0].n36 XThC.Tn[0].n34 161.406
R19900 XThC.Tn[0].n39 XThC.Tn[0].n37 161.406
R19901 XThC.Tn[0].n42 XThC.Tn[0].n40 161.406
R19902 XThC.Tn[0].n45 XThC.Tn[0].n43 161.406
R19903 XThC.Tn[0].n48 XThC.Tn[0].n46 161.406
R19904 XThC.Tn[0].n51 XThC.Tn[0].n49 161.406
R19905 XThC.Tn[0].n54 XThC.Tn[0].n52 161.406
R19906 XThC.Tn[0].n7 XThC.Tn[0].t22 161.202
R19907 XThC.Tn[0].n10 XThC.Tn[0].t41 161.202
R19908 XThC.Tn[0].n13 XThC.Tn[0].t12 161.202
R19909 XThC.Tn[0].n16 XThC.Tn[0].t13 161.202
R19910 XThC.Tn[0].n19 XThC.Tn[0].t32 161.202
R19911 XThC.Tn[0].n22 XThC.Tn[0].t34 161.202
R19912 XThC.Tn[0].n25 XThC.Tn[0].t17 161.202
R19913 XThC.Tn[0].n28 XThC.Tn[0].t25 161.202
R19914 XThC.Tn[0].n31 XThC.Tn[0].t26 161.202
R19915 XThC.Tn[0].n34 XThC.Tn[0].t15 161.202
R19916 XThC.Tn[0].n37 XThC.Tn[0].t16 161.202
R19917 XThC.Tn[0].n40 XThC.Tn[0].t27 161.202
R19918 XThC.Tn[0].n43 XThC.Tn[0].t36 161.202
R19919 XThC.Tn[0].n46 XThC.Tn[0].t38 161.202
R19920 XThC.Tn[0].n49 XThC.Tn[0].t19 161.202
R19921 XThC.Tn[0].n52 XThC.Tn[0].t29 161.202
R19922 XThC.Tn[0].n7 XThC.Tn[0].t18 145.137
R19923 XThC.Tn[0].n10 XThC.Tn[0].t35 145.137
R19924 XThC.Tn[0].n13 XThC.Tn[0].t37 145.137
R19925 XThC.Tn[0].n16 XThC.Tn[0].t39 145.137
R19926 XThC.Tn[0].n19 XThC.Tn[0].t28 145.137
R19927 XThC.Tn[0].n22 XThC.Tn[0].t30 145.137
R19928 XThC.Tn[0].n25 XThC.Tn[0].t43 145.137
R19929 XThC.Tn[0].n28 XThC.Tn[0].t20 145.137
R19930 XThC.Tn[0].n31 XThC.Tn[0].t21 145.137
R19931 XThC.Tn[0].n34 XThC.Tn[0].t40 145.137
R19932 XThC.Tn[0].n37 XThC.Tn[0].t42 145.137
R19933 XThC.Tn[0].n40 XThC.Tn[0].t23 145.137
R19934 XThC.Tn[0].n43 XThC.Tn[0].t31 145.137
R19935 XThC.Tn[0].n46 XThC.Tn[0].t33 145.137
R19936 XThC.Tn[0].n49 XThC.Tn[0].t14 145.137
R19937 XThC.Tn[0].n52 XThC.Tn[0].t24 145.137
R19938 XThC.Tn[0].n2 XThC.Tn[0].n0 135.248
R19939 XThC.Tn[0].n2 XThC.Tn[0].n1 98.982
R19940 XThC.Tn[0].n4 XThC.Tn[0].n3 98.982
R19941 XThC.Tn[0].n6 XThC.Tn[0].n5 98.982
R19942 XThC.Tn[0].n4 XThC.Tn[0].n2 36.2672
R19943 XThC.Tn[0].n6 XThC.Tn[0].n4 36.2672
R19944 XThC.Tn[0].n56 XThC.Tn[0].n6 32.6405
R19945 XThC.Tn[0].n57 XThC.Tn[0].t1 26.5955
R19946 XThC.Tn[0].n57 XThC.Tn[0].t0 26.5955
R19947 XThC.Tn[0].n58 XThC.Tn[0].t3 26.5955
R19948 XThC.Tn[0].n58 XThC.Tn[0].t2 26.5955
R19949 XThC.Tn[0].n0 XThC.Tn[0].t11 24.9236
R19950 XThC.Tn[0].n0 XThC.Tn[0].t8 24.9236
R19951 XThC.Tn[0].n1 XThC.Tn[0].t9 24.9236
R19952 XThC.Tn[0].n1 XThC.Tn[0].t10 24.9236
R19953 XThC.Tn[0].n3 XThC.Tn[0].t7 24.9236
R19954 XThC.Tn[0].n3 XThC.Tn[0].t6 24.9236
R19955 XThC.Tn[0].n5 XThC.Tn[0].t5 24.9236
R19956 XThC.Tn[0].n5 XThC.Tn[0].t4 24.9236
R19957 XThC.Tn[0].n60 XThC.Tn[0].n59 18.5605
R19958 XThC.Tn[0].n60 XThC.Tn[0].n56 11.5205
R19959 XThC.Tn[0].n56 XThC.Tn[0].n55 3.16389
R19960 XThC.Tn[0].n12 XThC.Tn[0] 0.931056
R19961 XThC.Tn[0].n15 XThC.Tn[0] 0.931056
R19962 XThC.Tn[0].n18 XThC.Tn[0] 0.931056
R19963 XThC.Tn[0].n21 XThC.Tn[0] 0.931056
R19964 XThC.Tn[0].n24 XThC.Tn[0] 0.931056
R19965 XThC.Tn[0].n27 XThC.Tn[0] 0.931056
R19966 XThC.Tn[0].n30 XThC.Tn[0] 0.931056
R19967 XThC.Tn[0].n33 XThC.Tn[0] 0.931056
R19968 XThC.Tn[0].n36 XThC.Tn[0] 0.931056
R19969 XThC.Tn[0].n39 XThC.Tn[0] 0.931056
R19970 XThC.Tn[0].n42 XThC.Tn[0] 0.931056
R19971 XThC.Tn[0].n45 XThC.Tn[0] 0.931056
R19972 XThC.Tn[0].n48 XThC.Tn[0] 0.931056
R19973 XThC.Tn[0].n51 XThC.Tn[0] 0.931056
R19974 XThC.Tn[0].n54 XThC.Tn[0] 0.931056
R19975 XThC.Tn[0] XThC.Tn[0].n60 0.6405
R19976 XThC.Tn[0] XThC.Tn[0].n9 0.396333
R19977 XThC.Tn[0] XThC.Tn[0].n12 0.396333
R19978 XThC.Tn[0] XThC.Tn[0].n15 0.396333
R19979 XThC.Tn[0] XThC.Tn[0].n18 0.396333
R19980 XThC.Tn[0] XThC.Tn[0].n21 0.396333
R19981 XThC.Tn[0] XThC.Tn[0].n24 0.396333
R19982 XThC.Tn[0] XThC.Tn[0].n27 0.396333
R19983 XThC.Tn[0] XThC.Tn[0].n30 0.396333
R19984 XThC.Tn[0] XThC.Tn[0].n33 0.396333
R19985 XThC.Tn[0] XThC.Tn[0].n36 0.396333
R19986 XThC.Tn[0] XThC.Tn[0].n39 0.396333
R19987 XThC.Tn[0] XThC.Tn[0].n42 0.396333
R19988 XThC.Tn[0] XThC.Tn[0].n45 0.396333
R19989 XThC.Tn[0] XThC.Tn[0].n48 0.396333
R19990 XThC.Tn[0] XThC.Tn[0].n51 0.396333
R19991 XThC.Tn[0] XThC.Tn[0].n54 0.396333
R19992 XThC.Tn[0].n55 XThC.Tn[0] 0.243556
R19993 XThC.Tn[0].n8 XThC.Tn[0] 0.104667
R19994 XThC.Tn[0].n11 XThC.Tn[0] 0.104667
R19995 XThC.Tn[0].n14 XThC.Tn[0] 0.104667
R19996 XThC.Tn[0].n17 XThC.Tn[0] 0.104667
R19997 XThC.Tn[0].n20 XThC.Tn[0] 0.104667
R19998 XThC.Tn[0].n23 XThC.Tn[0] 0.104667
R19999 XThC.Tn[0].n26 XThC.Tn[0] 0.104667
R20000 XThC.Tn[0].n29 XThC.Tn[0] 0.104667
R20001 XThC.Tn[0].n32 XThC.Tn[0] 0.104667
R20002 XThC.Tn[0].n35 XThC.Tn[0] 0.104667
R20003 XThC.Tn[0].n38 XThC.Tn[0] 0.104667
R20004 XThC.Tn[0].n41 XThC.Tn[0] 0.104667
R20005 XThC.Tn[0].n44 XThC.Tn[0] 0.104667
R20006 XThC.Tn[0].n47 XThC.Tn[0] 0.104667
R20007 XThC.Tn[0].n50 XThC.Tn[0] 0.104667
R20008 XThC.Tn[0].n53 XThC.Tn[0] 0.104667
R20009 XThC.Tn[0].n55 XThC.Tn[0] 0.0326429
R20010 XThC.Tn[0].n8 XThC.Tn[0] 0.0309878
R20011 XThC.Tn[0].n11 XThC.Tn[0] 0.0309878
R20012 XThC.Tn[0].n14 XThC.Tn[0] 0.0309878
R20013 XThC.Tn[0].n17 XThC.Tn[0] 0.0309878
R20014 XThC.Tn[0].n20 XThC.Tn[0] 0.0309878
R20015 XThC.Tn[0].n23 XThC.Tn[0] 0.0309878
R20016 XThC.Tn[0].n26 XThC.Tn[0] 0.0309878
R20017 XThC.Tn[0].n29 XThC.Tn[0] 0.0309878
R20018 XThC.Tn[0].n32 XThC.Tn[0] 0.0309878
R20019 XThC.Tn[0].n35 XThC.Tn[0] 0.0309878
R20020 XThC.Tn[0].n38 XThC.Tn[0] 0.0309878
R20021 XThC.Tn[0].n41 XThC.Tn[0] 0.0309878
R20022 XThC.Tn[0].n44 XThC.Tn[0] 0.0309878
R20023 XThC.Tn[0].n47 XThC.Tn[0] 0.0309878
R20024 XThC.Tn[0].n50 XThC.Tn[0] 0.0309878
R20025 XThC.Tn[0].n53 XThC.Tn[0] 0.0309878
R20026 XThC.Tn[0].n9 XThC.Tn[0].n8 0.027939
R20027 XThC.Tn[0].n12 XThC.Tn[0].n11 0.027939
R20028 XThC.Tn[0].n15 XThC.Tn[0].n14 0.027939
R20029 XThC.Tn[0].n18 XThC.Tn[0].n17 0.027939
R20030 XThC.Tn[0].n21 XThC.Tn[0].n20 0.027939
R20031 XThC.Tn[0].n24 XThC.Tn[0].n23 0.027939
R20032 XThC.Tn[0].n27 XThC.Tn[0].n26 0.027939
R20033 XThC.Tn[0].n30 XThC.Tn[0].n29 0.027939
R20034 XThC.Tn[0].n33 XThC.Tn[0].n32 0.027939
R20035 XThC.Tn[0].n36 XThC.Tn[0].n35 0.027939
R20036 XThC.Tn[0].n39 XThC.Tn[0].n38 0.027939
R20037 XThC.Tn[0].n42 XThC.Tn[0].n41 0.027939
R20038 XThC.Tn[0].n45 XThC.Tn[0].n44 0.027939
R20039 XThC.Tn[0].n48 XThC.Tn[0].n47 0.027939
R20040 XThC.Tn[0].n51 XThC.Tn[0].n50 0.027939
R20041 XThC.Tn[0].n54 XThC.Tn[0].n53 0.027939
R20042 XThC.XTB4.Y.t0 XThC.XTB4.Y.n21 268.738
R20043 XThC.XTB4.Y.n22 XThC.XTB4.Y.t0 268.077
R20044 XThC.XTB4.Y.n0 XThC.XTB4.Y.t1 235.56
R20045 XThC.XTB4.Y.n4 XThC.XTB4.Y.t3 212.081
R20046 XThC.XTB4.Y.n3 XThC.XTB4.Y.t2 212.081
R20047 XThC.XTB4.Y.n9 XThC.XTB4.Y.t17 212.081
R20048 XThC.XTB4.Y.n1 XThC.XTB4.Y.t13 212.081
R20049 XThC.XTB4.Y.n13 XThC.XTB4.Y.t8 212.081
R20050 XThC.XTB4.Y.n14 XThC.XTB4.Y.t12 212.081
R20051 XThC.XTB4.Y.n16 XThC.XTB4.Y.t6 212.081
R20052 XThC.XTB4.Y.n12 XThC.XTB4.Y.t16 212.081
R20053 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 173.761
R20054 XThC.XTB4.Y.n15 XThC.XTB4.Y 158.656
R20055 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 152
R20056 XThC.XTB4.Y.n6 XThC.XTB4.Y.n2 152
R20057 XThC.XTB4.Y.n11 XThC.XTB4.Y.n10 152
R20058 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 152
R20059 XThC.XTB4.Y.n4 XThC.XTB4.Y.t14 139.78
R20060 XThC.XTB4.Y.n3 XThC.XTB4.Y.t10 139.78
R20061 XThC.XTB4.Y.n9 XThC.XTB4.Y.t7 139.78
R20062 XThC.XTB4.Y.n1 XThC.XTB4.Y.t4 139.78
R20063 XThC.XTB4.Y.n13 XThC.XTB4.Y.t11 139.78
R20064 XThC.XTB4.Y.n14 XThC.XTB4.Y.t15 139.78
R20065 XThC.XTB4.Y.n16 XThC.XTB4.Y.t9 139.78
R20066 XThC.XTB4.Y.n12 XThC.XTB4.Y.t5 139.78
R20067 XThC.XTB4.Y.n20 XThC.XTB4.Y.n11 72.9296
R20068 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 61.346
R20069 XThC.XTB4.Y.n8 XThC.XTB4.Y.n2 49.6611
R20070 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 45.2793
R20071 XThC.XTB4.Y.n5 XThC.XTB4.Y.n3 42.3581
R20072 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 38.1854
R20073 XThC.XTB4.Y.n17 XThC.XTB4.Y.n12 30.6732
R20074 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 30.6732
R20075 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R20076 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R20077 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 21.7605
R20078 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 18.9884
R20079 XThC.XTB4.Y XThC.XTB4.Y.n22 17.8682
R20080 XThC.XTB4.Y.n10 XThC.XTB4.Y.n1 16.0672
R20081 XThC.XTB4.Y.n18 XThC.XTB4.Y 14.7905
R20082 XThC.XTB4.Y.n11 XThC.XTB4.Y 11.5205
R20083 XThC.XTB4.Y.n21 XThC.XTB4.Y.n20 10.353
R20084 XThC.XTB4.Y.n7 XThC.XTB4.Y 10.2405
R20085 XThC.XTB4.Y.n3 XThC.XTB4.Y.n2 7.30353
R20086 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 7.24578
R20087 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 4.38232
R20088 XThC.XTB4.Y.n22 XThC.XTB4.Y.n21 3.29747
R20089 XThC.XTB4.Y XThC.XTB4.Y.n0 2.22659
R20090 XThC.XTB4.Y.n0 XThC.XTB4.Y 1.55202
R20091 XThC.XTB4.Y.n19 XThC.XTB4.Y 0.966538
R20092 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R20093 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R20094 XThR.Tn[3] XThR.Tn[3].n82 161.363
R20095 XThR.Tn[3] XThR.Tn[3].n77 161.363
R20096 XThR.Tn[3] XThR.Tn[3].n72 161.363
R20097 XThR.Tn[3] XThR.Tn[3].n67 161.363
R20098 XThR.Tn[3] XThR.Tn[3].n62 161.363
R20099 XThR.Tn[3] XThR.Tn[3].n57 161.363
R20100 XThR.Tn[3] XThR.Tn[3].n52 161.363
R20101 XThR.Tn[3] XThR.Tn[3].n47 161.363
R20102 XThR.Tn[3] XThR.Tn[3].n42 161.363
R20103 XThR.Tn[3] XThR.Tn[3].n37 161.363
R20104 XThR.Tn[3] XThR.Tn[3].n32 161.363
R20105 XThR.Tn[3] XThR.Tn[3].n27 161.363
R20106 XThR.Tn[3] XThR.Tn[3].n22 161.363
R20107 XThR.Tn[3] XThR.Tn[3].n17 161.363
R20108 XThR.Tn[3] XThR.Tn[3].n12 161.363
R20109 XThR.Tn[3] XThR.Tn[3].n10 161.363
R20110 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R20111 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R20112 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R20113 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R20114 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R20115 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R20116 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R20117 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R20118 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R20119 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R20120 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R20121 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R20122 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R20123 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R20124 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R20125 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R20126 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R20127 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R20128 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R20129 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R20130 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R20131 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R20132 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R20133 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R20134 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R20135 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R20136 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R20137 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R20138 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R20139 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R20140 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R20141 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R20142 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R20143 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R20144 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R20145 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R20146 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R20147 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R20148 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R20149 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R20150 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R20151 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R20152 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R20153 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R20154 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R20155 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R20156 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R20157 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R20158 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R20159 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R20160 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R20161 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R20162 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R20163 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R20164 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R20165 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R20166 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R20167 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R20168 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R20169 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R20170 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R20171 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R20172 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R20173 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R20174 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R20175 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R20176 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R20177 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R20178 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R20179 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R20180 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R20181 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R20182 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R20183 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R20184 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R20185 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R20186 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R20187 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R20188 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R20189 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R20190 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R20191 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R20192 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R20193 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R20194 XThR.Tn[3].n1 XThR.Tn[3].t8 26.5955
R20195 XThR.Tn[3].n1 XThR.Tn[3].t11 26.5955
R20196 XThR.Tn[3].n0 XThR.Tn[3].t9 26.5955
R20197 XThR.Tn[3].n0 XThR.Tn[3].t10 26.5955
R20198 XThR.Tn[3].n3 XThR.Tn[3].t7 24.9236
R20199 XThR.Tn[3].n3 XThR.Tn[3].t4 24.9236
R20200 XThR.Tn[3].n4 XThR.Tn[3].t6 24.9236
R20201 XThR.Tn[3].n4 XThR.Tn[3].t5 24.9236
R20202 XThR.Tn[3].n5 XThR.Tn[3].t0 24.9236
R20203 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R20204 XThR.Tn[3].n6 XThR.Tn[3].t3 24.9236
R20205 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R20206 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R20207 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R20208 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R20209 XThR.Tn[3] XThR.Tn[3].n11 5.4407
R20210 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R20211 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R20212 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R20213 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R20214 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R20215 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R20216 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R20217 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R20218 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R20219 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R20220 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R20221 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R20222 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R20223 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R20224 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R20225 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R20226 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R20227 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R20228 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R20229 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R20230 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R20231 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R20232 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R20233 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R20234 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R20235 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R20236 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R20237 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R20238 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R20239 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R20240 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R20241 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R20242 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R20243 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R20244 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R20245 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R20246 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R20247 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R20248 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R20249 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R20250 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R20251 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R20252 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R20253 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R20254 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R20255 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R20256 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R20257 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R20258 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R20259 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R20260 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R20261 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R20262 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R20263 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R20264 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R20265 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R20266 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R20267 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R20268 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R20269 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R20270 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R20271 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R20272 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R20273 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R20274 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R20275 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R20276 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R20277 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R20278 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R20279 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R20280 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R20281 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R20282 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R20283 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R20284 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R20285 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R20286 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R20287 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R20288 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R20289 XThR.Tn[3] XThR.Tn[3].n87 0.038
R20290 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R20291 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R20292 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R20293 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R20294 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R20295 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R20296 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R20297 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R20298 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R20299 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R20300 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R20301 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R20302 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R20303 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R20304 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R20305 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R20306 XThR.Tn[5].n88 XThR.Tn[5].n87 332.332
R20307 XThR.Tn[5].n88 XThR.Tn[5].n86 296.493
R20308 XThR.Tn[5] XThR.Tn[5].n79 161.363
R20309 XThR.Tn[5] XThR.Tn[5].n74 161.363
R20310 XThR.Tn[5] XThR.Tn[5].n69 161.363
R20311 XThR.Tn[5] XThR.Tn[5].n64 161.363
R20312 XThR.Tn[5] XThR.Tn[5].n59 161.363
R20313 XThR.Tn[5] XThR.Tn[5].n54 161.363
R20314 XThR.Tn[5] XThR.Tn[5].n49 161.363
R20315 XThR.Tn[5] XThR.Tn[5].n44 161.363
R20316 XThR.Tn[5] XThR.Tn[5].n39 161.363
R20317 XThR.Tn[5] XThR.Tn[5].n34 161.363
R20318 XThR.Tn[5] XThR.Tn[5].n29 161.363
R20319 XThR.Tn[5] XThR.Tn[5].n24 161.363
R20320 XThR.Tn[5] XThR.Tn[5].n19 161.363
R20321 XThR.Tn[5] XThR.Tn[5].n14 161.363
R20322 XThR.Tn[5] XThR.Tn[5].n9 161.363
R20323 XThR.Tn[5] XThR.Tn[5].n7 161.363
R20324 XThR.Tn[5].n81 XThR.Tn[5].n80 161.3
R20325 XThR.Tn[5].n76 XThR.Tn[5].n75 161.3
R20326 XThR.Tn[5].n71 XThR.Tn[5].n70 161.3
R20327 XThR.Tn[5].n66 XThR.Tn[5].n65 161.3
R20328 XThR.Tn[5].n61 XThR.Tn[5].n60 161.3
R20329 XThR.Tn[5].n56 XThR.Tn[5].n55 161.3
R20330 XThR.Tn[5].n51 XThR.Tn[5].n50 161.3
R20331 XThR.Tn[5].n46 XThR.Tn[5].n45 161.3
R20332 XThR.Tn[5].n41 XThR.Tn[5].n40 161.3
R20333 XThR.Tn[5].n36 XThR.Tn[5].n35 161.3
R20334 XThR.Tn[5].n31 XThR.Tn[5].n30 161.3
R20335 XThR.Tn[5].n26 XThR.Tn[5].n25 161.3
R20336 XThR.Tn[5].n21 XThR.Tn[5].n20 161.3
R20337 XThR.Tn[5].n16 XThR.Tn[5].n15 161.3
R20338 XThR.Tn[5].n11 XThR.Tn[5].n10 161.3
R20339 XThR.Tn[5].n79 XThR.Tn[5].t62 161.106
R20340 XThR.Tn[5].n74 XThR.Tn[5].t70 161.106
R20341 XThR.Tn[5].n69 XThR.Tn[5].t52 161.106
R20342 XThR.Tn[5].n64 XThR.Tn[5].t35 161.106
R20343 XThR.Tn[5].n59 XThR.Tn[5].t60 161.106
R20344 XThR.Tn[5].n54 XThR.Tn[5].t24 161.106
R20345 XThR.Tn[5].n49 XThR.Tn[5].t68 161.106
R20346 XThR.Tn[5].n44 XThR.Tn[5].t49 161.106
R20347 XThR.Tn[5].n39 XThR.Tn[5].t32 161.106
R20348 XThR.Tn[5].n34 XThR.Tn[5].t40 161.106
R20349 XThR.Tn[5].n29 XThR.Tn[5].t22 161.106
R20350 XThR.Tn[5].n24 XThR.Tn[5].t51 161.106
R20351 XThR.Tn[5].n19 XThR.Tn[5].t21 161.106
R20352 XThR.Tn[5].n14 XThR.Tn[5].t66 161.106
R20353 XThR.Tn[5].n9 XThR.Tn[5].t26 161.106
R20354 XThR.Tn[5].n7 XThR.Tn[5].t72 161.106
R20355 XThR.Tn[5].n80 XThR.Tn[5].t59 159.978
R20356 XThR.Tn[5].n75 XThR.Tn[5].t64 159.978
R20357 XThR.Tn[5].n70 XThR.Tn[5].t47 159.978
R20358 XThR.Tn[5].n65 XThR.Tn[5].t31 159.978
R20359 XThR.Tn[5].n60 XThR.Tn[5].t57 159.978
R20360 XThR.Tn[5].n55 XThR.Tn[5].t20 159.978
R20361 XThR.Tn[5].n50 XThR.Tn[5].t63 159.978
R20362 XThR.Tn[5].n45 XThR.Tn[5].t45 159.978
R20363 XThR.Tn[5].n40 XThR.Tn[5].t29 159.978
R20364 XThR.Tn[5].n35 XThR.Tn[5].t37 159.978
R20365 XThR.Tn[5].n30 XThR.Tn[5].t19 159.978
R20366 XThR.Tn[5].n25 XThR.Tn[5].t46 159.978
R20367 XThR.Tn[5].n20 XThR.Tn[5].t18 159.978
R20368 XThR.Tn[5].n15 XThR.Tn[5].t61 159.978
R20369 XThR.Tn[5].n10 XThR.Tn[5].t23 159.978
R20370 XThR.Tn[5].n79 XThR.Tn[5].t54 145.038
R20371 XThR.Tn[5].n74 XThR.Tn[5].t12 145.038
R20372 XThR.Tn[5].n69 XThR.Tn[5].t56 145.038
R20373 XThR.Tn[5].n64 XThR.Tn[5].t41 145.038
R20374 XThR.Tn[5].n59 XThR.Tn[5].t71 145.038
R20375 XThR.Tn[5].n54 XThR.Tn[5].t53 145.038
R20376 XThR.Tn[5].n49 XThR.Tn[5].t58 145.038
R20377 XThR.Tn[5].n44 XThR.Tn[5].t42 145.038
R20378 XThR.Tn[5].n39 XThR.Tn[5].t38 145.038
R20379 XThR.Tn[5].n34 XThR.Tn[5].t69 145.038
R20380 XThR.Tn[5].n29 XThR.Tn[5].t30 145.038
R20381 XThR.Tn[5].n24 XThR.Tn[5].t55 145.038
R20382 XThR.Tn[5].n19 XThR.Tn[5].t28 145.038
R20383 XThR.Tn[5].n14 XThR.Tn[5].t73 145.038
R20384 XThR.Tn[5].n9 XThR.Tn[5].t39 145.038
R20385 XThR.Tn[5].n7 XThR.Tn[5].t17 145.038
R20386 XThR.Tn[5].n80 XThR.Tn[5].t27 143.911
R20387 XThR.Tn[5].n75 XThR.Tn[5].t50 143.911
R20388 XThR.Tn[5].n70 XThR.Tn[5].t34 143.911
R20389 XThR.Tn[5].n65 XThR.Tn[5].t15 143.911
R20390 XThR.Tn[5].n60 XThR.Tn[5].t44 143.911
R20391 XThR.Tn[5].n55 XThR.Tn[5].t25 143.911
R20392 XThR.Tn[5].n50 XThR.Tn[5].t36 143.911
R20393 XThR.Tn[5].n45 XThR.Tn[5].t16 143.911
R20394 XThR.Tn[5].n40 XThR.Tn[5].t14 143.911
R20395 XThR.Tn[5].n35 XThR.Tn[5].t43 143.911
R20396 XThR.Tn[5].n30 XThR.Tn[5].t67 143.911
R20397 XThR.Tn[5].n25 XThR.Tn[5].t33 143.911
R20398 XThR.Tn[5].n20 XThR.Tn[5].t65 143.911
R20399 XThR.Tn[5].n15 XThR.Tn[5].t48 143.911
R20400 XThR.Tn[5].n10 XThR.Tn[5].t13 143.911
R20401 XThR.Tn[5].n2 XThR.Tn[5].n0 135.249
R20402 XThR.Tn[5].n2 XThR.Tn[5].n1 98.981
R20403 XThR.Tn[5].n4 XThR.Tn[5].n3 98.981
R20404 XThR.Tn[5].n6 XThR.Tn[5].n5 98.981
R20405 XThR.Tn[5].n4 XThR.Tn[5].n2 36.2672
R20406 XThR.Tn[5].n6 XThR.Tn[5].n4 36.2672
R20407 XThR.Tn[5].n85 XThR.Tn[5].n6 32.6405
R20408 XThR.Tn[5].n87 XThR.Tn[5].t1 26.5955
R20409 XThR.Tn[5].n87 XThR.Tn[5].t0 26.5955
R20410 XThR.Tn[5].n86 XThR.Tn[5].t2 26.5955
R20411 XThR.Tn[5].n86 XThR.Tn[5].t3 26.5955
R20412 XThR.Tn[5].n0 XThR.Tn[5].t8 24.9236
R20413 XThR.Tn[5].n0 XThR.Tn[5].t9 24.9236
R20414 XThR.Tn[5].n1 XThR.Tn[5].t11 24.9236
R20415 XThR.Tn[5].n1 XThR.Tn[5].t10 24.9236
R20416 XThR.Tn[5].n3 XThR.Tn[5].t6 24.9236
R20417 XThR.Tn[5].n3 XThR.Tn[5].t5 24.9236
R20418 XThR.Tn[5].n5 XThR.Tn[5].t7 24.9236
R20419 XThR.Tn[5].n5 XThR.Tn[5].t4 24.9236
R20420 XThR.Tn[5].n89 XThR.Tn[5].n88 18.5605
R20421 XThR.Tn[5].n89 XThR.Tn[5].n85 11.5205
R20422 XThR.Tn[5].n85 XThR.Tn[5] 5.71508
R20423 XThR.Tn[5] XThR.Tn[5].n8 5.4407
R20424 XThR.Tn[5].n13 XThR.Tn[5].n12 4.5005
R20425 XThR.Tn[5].n18 XThR.Tn[5].n17 4.5005
R20426 XThR.Tn[5].n23 XThR.Tn[5].n22 4.5005
R20427 XThR.Tn[5].n28 XThR.Tn[5].n27 4.5005
R20428 XThR.Tn[5].n33 XThR.Tn[5].n32 4.5005
R20429 XThR.Tn[5].n38 XThR.Tn[5].n37 4.5005
R20430 XThR.Tn[5].n43 XThR.Tn[5].n42 4.5005
R20431 XThR.Tn[5].n48 XThR.Tn[5].n47 4.5005
R20432 XThR.Tn[5].n53 XThR.Tn[5].n52 4.5005
R20433 XThR.Tn[5].n58 XThR.Tn[5].n57 4.5005
R20434 XThR.Tn[5].n63 XThR.Tn[5].n62 4.5005
R20435 XThR.Tn[5].n68 XThR.Tn[5].n67 4.5005
R20436 XThR.Tn[5].n73 XThR.Tn[5].n72 4.5005
R20437 XThR.Tn[5].n78 XThR.Tn[5].n77 4.5005
R20438 XThR.Tn[5].n83 XThR.Tn[5].n82 4.5005
R20439 XThR.Tn[5].n84 XThR.Tn[5] 3.70586
R20440 XThR.Tn[5].n13 XThR.Tn[5] 2.52282
R20441 XThR.Tn[5].n18 XThR.Tn[5] 2.52282
R20442 XThR.Tn[5].n23 XThR.Tn[5] 2.52282
R20443 XThR.Tn[5].n28 XThR.Tn[5] 2.52282
R20444 XThR.Tn[5].n33 XThR.Tn[5] 2.52282
R20445 XThR.Tn[5].n38 XThR.Tn[5] 2.52282
R20446 XThR.Tn[5].n43 XThR.Tn[5] 2.52282
R20447 XThR.Tn[5].n48 XThR.Tn[5] 2.52282
R20448 XThR.Tn[5].n53 XThR.Tn[5] 2.52282
R20449 XThR.Tn[5].n58 XThR.Tn[5] 2.52282
R20450 XThR.Tn[5].n63 XThR.Tn[5] 2.52282
R20451 XThR.Tn[5].n68 XThR.Tn[5] 2.52282
R20452 XThR.Tn[5].n73 XThR.Tn[5] 2.52282
R20453 XThR.Tn[5].n78 XThR.Tn[5] 2.52282
R20454 XThR.Tn[5].n83 XThR.Tn[5] 2.52282
R20455 XThR.Tn[5].n81 XThR.Tn[5] 1.08677
R20456 XThR.Tn[5].n76 XThR.Tn[5] 1.08677
R20457 XThR.Tn[5].n71 XThR.Tn[5] 1.08677
R20458 XThR.Tn[5].n66 XThR.Tn[5] 1.08677
R20459 XThR.Tn[5].n61 XThR.Tn[5] 1.08677
R20460 XThR.Tn[5].n56 XThR.Tn[5] 1.08677
R20461 XThR.Tn[5].n51 XThR.Tn[5] 1.08677
R20462 XThR.Tn[5].n46 XThR.Tn[5] 1.08677
R20463 XThR.Tn[5].n41 XThR.Tn[5] 1.08677
R20464 XThR.Tn[5].n36 XThR.Tn[5] 1.08677
R20465 XThR.Tn[5].n31 XThR.Tn[5] 1.08677
R20466 XThR.Tn[5].n26 XThR.Tn[5] 1.08677
R20467 XThR.Tn[5].n21 XThR.Tn[5] 1.08677
R20468 XThR.Tn[5].n16 XThR.Tn[5] 1.08677
R20469 XThR.Tn[5].n11 XThR.Tn[5] 1.08677
R20470 XThR.Tn[5] XThR.Tn[5].n13 0.839786
R20471 XThR.Tn[5] XThR.Tn[5].n18 0.839786
R20472 XThR.Tn[5] XThR.Tn[5].n23 0.839786
R20473 XThR.Tn[5] XThR.Tn[5].n28 0.839786
R20474 XThR.Tn[5] XThR.Tn[5].n33 0.839786
R20475 XThR.Tn[5] XThR.Tn[5].n38 0.839786
R20476 XThR.Tn[5] XThR.Tn[5].n43 0.839786
R20477 XThR.Tn[5] XThR.Tn[5].n48 0.839786
R20478 XThR.Tn[5] XThR.Tn[5].n53 0.839786
R20479 XThR.Tn[5] XThR.Tn[5].n58 0.839786
R20480 XThR.Tn[5] XThR.Tn[5].n63 0.839786
R20481 XThR.Tn[5] XThR.Tn[5].n68 0.839786
R20482 XThR.Tn[5] XThR.Tn[5].n73 0.839786
R20483 XThR.Tn[5] XThR.Tn[5].n78 0.839786
R20484 XThR.Tn[5] XThR.Tn[5].n83 0.839786
R20485 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R20486 XThR.Tn[5].n8 XThR.Tn[5] 0.499542
R20487 XThR.Tn[5].n82 XThR.Tn[5] 0.063
R20488 XThR.Tn[5].n77 XThR.Tn[5] 0.063
R20489 XThR.Tn[5].n72 XThR.Tn[5] 0.063
R20490 XThR.Tn[5].n67 XThR.Tn[5] 0.063
R20491 XThR.Tn[5].n62 XThR.Tn[5] 0.063
R20492 XThR.Tn[5].n57 XThR.Tn[5] 0.063
R20493 XThR.Tn[5].n52 XThR.Tn[5] 0.063
R20494 XThR.Tn[5].n47 XThR.Tn[5] 0.063
R20495 XThR.Tn[5].n42 XThR.Tn[5] 0.063
R20496 XThR.Tn[5].n37 XThR.Tn[5] 0.063
R20497 XThR.Tn[5].n32 XThR.Tn[5] 0.063
R20498 XThR.Tn[5].n27 XThR.Tn[5] 0.063
R20499 XThR.Tn[5].n22 XThR.Tn[5] 0.063
R20500 XThR.Tn[5].n17 XThR.Tn[5] 0.063
R20501 XThR.Tn[5].n12 XThR.Tn[5] 0.063
R20502 XThR.Tn[5].n84 XThR.Tn[5] 0.0540714
R20503 XThR.Tn[5] XThR.Tn[5].n84 0.038
R20504 XThR.Tn[5].n8 XThR.Tn[5] 0.0143889
R20505 XThR.Tn[5].n82 XThR.Tn[5].n81 0.00771154
R20506 XThR.Tn[5].n77 XThR.Tn[5].n76 0.00771154
R20507 XThR.Tn[5].n72 XThR.Tn[5].n71 0.00771154
R20508 XThR.Tn[5].n67 XThR.Tn[5].n66 0.00771154
R20509 XThR.Tn[5].n62 XThR.Tn[5].n61 0.00771154
R20510 XThR.Tn[5].n57 XThR.Tn[5].n56 0.00771154
R20511 XThR.Tn[5].n52 XThR.Tn[5].n51 0.00771154
R20512 XThR.Tn[5].n47 XThR.Tn[5].n46 0.00771154
R20513 XThR.Tn[5].n42 XThR.Tn[5].n41 0.00771154
R20514 XThR.Tn[5].n37 XThR.Tn[5].n36 0.00771154
R20515 XThR.Tn[5].n32 XThR.Tn[5].n31 0.00771154
R20516 XThR.Tn[5].n27 XThR.Tn[5].n26 0.00771154
R20517 XThR.Tn[5].n22 XThR.Tn[5].n21 0.00771154
R20518 XThR.Tn[5].n17 XThR.Tn[5].n16 0.00771154
R20519 XThR.Tn[5].n12 XThR.Tn[5].n11 0.00771154
R20520 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R20521 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R20522 XThC.Tn[4].n12 XThC.Tn[4].n10 161.406
R20523 XThC.Tn[4].n15 XThC.Tn[4].n13 161.406
R20524 XThC.Tn[4].n18 XThC.Tn[4].n16 161.406
R20525 XThC.Tn[4].n21 XThC.Tn[4].n19 161.406
R20526 XThC.Tn[4].n24 XThC.Tn[4].n22 161.406
R20527 XThC.Tn[4].n27 XThC.Tn[4].n25 161.406
R20528 XThC.Tn[4].n30 XThC.Tn[4].n28 161.406
R20529 XThC.Tn[4].n33 XThC.Tn[4].n31 161.406
R20530 XThC.Tn[4].n36 XThC.Tn[4].n34 161.406
R20531 XThC.Tn[4].n39 XThC.Tn[4].n37 161.406
R20532 XThC.Tn[4].n42 XThC.Tn[4].n40 161.406
R20533 XThC.Tn[4].n45 XThC.Tn[4].n43 161.406
R20534 XThC.Tn[4].n48 XThC.Tn[4].n46 161.406
R20535 XThC.Tn[4].n51 XThC.Tn[4].n49 161.406
R20536 XThC.Tn[4].n54 XThC.Tn[4].n52 161.406
R20537 XThC.Tn[4].n57 XThC.Tn[4].n55 161.406
R20538 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R20539 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R20540 XThC.Tn[4].n16 XThC.Tn[4].t13 161.202
R20541 XThC.Tn[4].n19 XThC.Tn[4].t15 161.202
R20542 XThC.Tn[4].n22 XThC.Tn[4].t36 161.202
R20543 XThC.Tn[4].n25 XThC.Tn[4].t37 161.202
R20544 XThC.Tn[4].n28 XThC.Tn[4].t18 161.202
R20545 XThC.Tn[4].n31 XThC.Tn[4].t27 161.202
R20546 XThC.Tn[4].n34 XThC.Tn[4].t29 161.202
R20547 XThC.Tn[4].n37 XThC.Tn[4].t16 161.202
R20548 XThC.Tn[4].n40 XThC.Tn[4].t17 161.202
R20549 XThC.Tn[4].n43 XThC.Tn[4].t30 161.202
R20550 XThC.Tn[4].n46 XThC.Tn[4].t38 161.202
R20551 XThC.Tn[4].n49 XThC.Tn[4].t41 161.202
R20552 XThC.Tn[4].n52 XThC.Tn[4].t22 161.202
R20553 XThC.Tn[4].n55 XThC.Tn[4].t32 161.202
R20554 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R20555 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R20556 XThC.Tn[4].n16 XThC.Tn[4].t19 145.137
R20557 XThC.Tn[4].n19 XThC.Tn[4].t20 145.137
R20558 XThC.Tn[4].n22 XThC.Tn[4].t39 145.137
R20559 XThC.Tn[4].n25 XThC.Tn[4].t40 145.137
R20560 XThC.Tn[4].n28 XThC.Tn[4].t24 145.137
R20561 XThC.Tn[4].n31 XThC.Tn[4].t31 145.137
R20562 XThC.Tn[4].n34 XThC.Tn[4].t33 145.137
R20563 XThC.Tn[4].n37 XThC.Tn[4].t21 145.137
R20564 XThC.Tn[4].n40 XThC.Tn[4].t23 145.137
R20565 XThC.Tn[4].n43 XThC.Tn[4].t34 145.137
R20566 XThC.Tn[4].n46 XThC.Tn[4].t42 145.137
R20567 XThC.Tn[4].n49 XThC.Tn[4].t12 145.137
R20568 XThC.Tn[4].n52 XThC.Tn[4].t25 145.137
R20569 XThC.Tn[4].n55 XThC.Tn[4].t35 145.137
R20570 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R20571 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R20572 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R20573 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R20574 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R20575 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R20576 XThC.Tn[4].n59 XThC.Tn[4].n9 32.6405
R20577 XThC.Tn[4].n1 XThC.Tn[4].t11 26.5955
R20578 XThC.Tn[4].n1 XThC.Tn[4].t10 26.5955
R20579 XThC.Tn[4].n0 XThC.Tn[4].t9 26.5955
R20580 XThC.Tn[4].n0 XThC.Tn[4].t8 26.5955
R20581 XThC.Tn[4].n3 XThC.Tn[4].t5 24.9236
R20582 XThC.Tn[4].n3 XThC.Tn[4].t4 24.9236
R20583 XThC.Tn[4].n4 XThC.Tn[4].t7 24.9236
R20584 XThC.Tn[4].n4 XThC.Tn[4].t6 24.9236
R20585 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R20586 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R20587 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R20588 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R20589 XThC.Tn[4].n60 XThC.Tn[4].n2 18.5605
R20590 XThC.Tn[4].n60 XThC.Tn[4].n59 11.5205
R20591 XThC.Tn[4].n58 XThC.Tn[4] 4.63701
R20592 XThC.Tn[4].n59 XThC.Tn[4].n58 3.1844
R20593 XThC.Tn[4].n15 XThC.Tn[4] 0.931056
R20594 XThC.Tn[4].n18 XThC.Tn[4] 0.931056
R20595 XThC.Tn[4].n21 XThC.Tn[4] 0.931056
R20596 XThC.Tn[4].n24 XThC.Tn[4] 0.931056
R20597 XThC.Tn[4].n27 XThC.Tn[4] 0.931056
R20598 XThC.Tn[4].n30 XThC.Tn[4] 0.931056
R20599 XThC.Tn[4].n33 XThC.Tn[4] 0.931056
R20600 XThC.Tn[4].n36 XThC.Tn[4] 0.931056
R20601 XThC.Tn[4].n39 XThC.Tn[4] 0.931056
R20602 XThC.Tn[4].n42 XThC.Tn[4] 0.931056
R20603 XThC.Tn[4].n45 XThC.Tn[4] 0.931056
R20604 XThC.Tn[4].n48 XThC.Tn[4] 0.931056
R20605 XThC.Tn[4].n51 XThC.Tn[4] 0.931056
R20606 XThC.Tn[4].n54 XThC.Tn[4] 0.931056
R20607 XThC.Tn[4].n57 XThC.Tn[4] 0.931056
R20608 XThC.Tn[4] XThC.Tn[4].n60 0.6405
R20609 XThC.Tn[4] XThC.Tn[4].n12 0.396333
R20610 XThC.Tn[4] XThC.Tn[4].n15 0.396333
R20611 XThC.Tn[4] XThC.Tn[4].n18 0.396333
R20612 XThC.Tn[4] XThC.Tn[4].n21 0.396333
R20613 XThC.Tn[4] XThC.Tn[4].n24 0.396333
R20614 XThC.Tn[4] XThC.Tn[4].n27 0.396333
R20615 XThC.Tn[4] XThC.Tn[4].n30 0.396333
R20616 XThC.Tn[4] XThC.Tn[4].n33 0.396333
R20617 XThC.Tn[4] XThC.Tn[4].n36 0.396333
R20618 XThC.Tn[4] XThC.Tn[4].n39 0.396333
R20619 XThC.Tn[4] XThC.Tn[4].n42 0.396333
R20620 XThC.Tn[4] XThC.Tn[4].n45 0.396333
R20621 XThC.Tn[4] XThC.Tn[4].n48 0.396333
R20622 XThC.Tn[4] XThC.Tn[4].n51 0.396333
R20623 XThC.Tn[4] XThC.Tn[4].n54 0.396333
R20624 XThC.Tn[4] XThC.Tn[4].n57 0.396333
R20625 XThC.Tn[4].n11 XThC.Tn[4] 0.104667
R20626 XThC.Tn[4].n14 XThC.Tn[4] 0.104667
R20627 XThC.Tn[4].n17 XThC.Tn[4] 0.104667
R20628 XThC.Tn[4].n20 XThC.Tn[4] 0.104667
R20629 XThC.Tn[4].n23 XThC.Tn[4] 0.104667
R20630 XThC.Tn[4].n26 XThC.Tn[4] 0.104667
R20631 XThC.Tn[4].n29 XThC.Tn[4] 0.104667
R20632 XThC.Tn[4].n32 XThC.Tn[4] 0.104667
R20633 XThC.Tn[4].n35 XThC.Tn[4] 0.104667
R20634 XThC.Tn[4].n38 XThC.Tn[4] 0.104667
R20635 XThC.Tn[4].n41 XThC.Tn[4] 0.104667
R20636 XThC.Tn[4].n44 XThC.Tn[4] 0.104667
R20637 XThC.Tn[4].n47 XThC.Tn[4] 0.104667
R20638 XThC.Tn[4].n50 XThC.Tn[4] 0.104667
R20639 XThC.Tn[4].n53 XThC.Tn[4] 0.104667
R20640 XThC.Tn[4].n56 XThC.Tn[4] 0.104667
R20641 XThC.Tn[4].n11 XThC.Tn[4] 0.0309878
R20642 XThC.Tn[4].n14 XThC.Tn[4] 0.0309878
R20643 XThC.Tn[4].n17 XThC.Tn[4] 0.0309878
R20644 XThC.Tn[4].n20 XThC.Tn[4] 0.0309878
R20645 XThC.Tn[4].n23 XThC.Tn[4] 0.0309878
R20646 XThC.Tn[4].n26 XThC.Tn[4] 0.0309878
R20647 XThC.Tn[4].n29 XThC.Tn[4] 0.0309878
R20648 XThC.Tn[4].n32 XThC.Tn[4] 0.0309878
R20649 XThC.Tn[4].n35 XThC.Tn[4] 0.0309878
R20650 XThC.Tn[4].n38 XThC.Tn[4] 0.0309878
R20651 XThC.Tn[4].n41 XThC.Tn[4] 0.0309878
R20652 XThC.Tn[4].n44 XThC.Tn[4] 0.0309878
R20653 XThC.Tn[4].n47 XThC.Tn[4] 0.0309878
R20654 XThC.Tn[4].n50 XThC.Tn[4] 0.0309878
R20655 XThC.Tn[4].n53 XThC.Tn[4] 0.0309878
R20656 XThC.Tn[4].n56 XThC.Tn[4] 0.0309878
R20657 XThC.Tn[4].n12 XThC.Tn[4].n11 0.027939
R20658 XThC.Tn[4].n15 XThC.Tn[4].n14 0.027939
R20659 XThC.Tn[4].n18 XThC.Tn[4].n17 0.027939
R20660 XThC.Tn[4].n21 XThC.Tn[4].n20 0.027939
R20661 XThC.Tn[4].n24 XThC.Tn[4].n23 0.027939
R20662 XThC.Tn[4].n27 XThC.Tn[4].n26 0.027939
R20663 XThC.Tn[4].n30 XThC.Tn[4].n29 0.027939
R20664 XThC.Tn[4].n33 XThC.Tn[4].n32 0.027939
R20665 XThC.Tn[4].n36 XThC.Tn[4].n35 0.027939
R20666 XThC.Tn[4].n39 XThC.Tn[4].n38 0.027939
R20667 XThC.Tn[4].n42 XThC.Tn[4].n41 0.027939
R20668 XThC.Tn[4].n45 XThC.Tn[4].n44 0.027939
R20669 XThC.Tn[4].n48 XThC.Tn[4].n47 0.027939
R20670 XThC.Tn[4].n51 XThC.Tn[4].n50 0.027939
R20671 XThC.Tn[4].n54 XThC.Tn[4].n53 0.027939
R20672 XThC.Tn[4].n57 XThC.Tn[4].n56 0.027939
R20673 XThC.Tn[4].n58 XThC.Tn[4] 0.0129465
R20674 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R20675 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R20676 XThC.Tn[2].n12 XThC.Tn[2].n10 161.406
R20677 XThC.Tn[2].n15 XThC.Tn[2].n13 161.406
R20678 XThC.Tn[2].n18 XThC.Tn[2].n16 161.406
R20679 XThC.Tn[2].n21 XThC.Tn[2].n19 161.406
R20680 XThC.Tn[2].n24 XThC.Tn[2].n22 161.406
R20681 XThC.Tn[2].n27 XThC.Tn[2].n25 161.406
R20682 XThC.Tn[2].n30 XThC.Tn[2].n28 161.406
R20683 XThC.Tn[2].n33 XThC.Tn[2].n31 161.406
R20684 XThC.Tn[2].n36 XThC.Tn[2].n34 161.406
R20685 XThC.Tn[2].n39 XThC.Tn[2].n37 161.406
R20686 XThC.Tn[2].n42 XThC.Tn[2].n40 161.406
R20687 XThC.Tn[2].n45 XThC.Tn[2].n43 161.406
R20688 XThC.Tn[2].n48 XThC.Tn[2].n46 161.406
R20689 XThC.Tn[2].n51 XThC.Tn[2].n49 161.406
R20690 XThC.Tn[2].n54 XThC.Tn[2].n52 161.406
R20691 XThC.Tn[2].n57 XThC.Tn[2].n55 161.406
R20692 XThC.Tn[2].n10 XThC.Tn[2].t18 161.202
R20693 XThC.Tn[2].n13 XThC.Tn[2].t35 161.202
R20694 XThC.Tn[2].n16 XThC.Tn[2].t37 161.202
R20695 XThC.Tn[2].n19 XThC.Tn[2].t39 161.202
R20696 XThC.Tn[2].n22 XThC.Tn[2].t28 161.202
R20697 XThC.Tn[2].n25 XThC.Tn[2].t29 161.202
R20698 XThC.Tn[2].n28 XThC.Tn[2].t42 161.202
R20699 XThC.Tn[2].n31 XThC.Tn[2].t19 161.202
R20700 XThC.Tn[2].n34 XThC.Tn[2].t21 161.202
R20701 XThC.Tn[2].n37 XThC.Tn[2].t40 161.202
R20702 XThC.Tn[2].n40 XThC.Tn[2].t41 161.202
R20703 XThC.Tn[2].n43 XThC.Tn[2].t22 161.202
R20704 XThC.Tn[2].n46 XThC.Tn[2].t30 161.202
R20705 XThC.Tn[2].n49 XThC.Tn[2].t33 161.202
R20706 XThC.Tn[2].n52 XThC.Tn[2].t14 161.202
R20707 XThC.Tn[2].n55 XThC.Tn[2].t24 161.202
R20708 XThC.Tn[2].n10 XThC.Tn[2].t20 145.137
R20709 XThC.Tn[2].n13 XThC.Tn[2].t38 145.137
R20710 XThC.Tn[2].n16 XThC.Tn[2].t43 145.137
R20711 XThC.Tn[2].n19 XThC.Tn[2].t12 145.137
R20712 XThC.Tn[2].n22 XThC.Tn[2].t31 145.137
R20713 XThC.Tn[2].n25 XThC.Tn[2].t32 145.137
R20714 XThC.Tn[2].n28 XThC.Tn[2].t16 145.137
R20715 XThC.Tn[2].n31 XThC.Tn[2].t23 145.137
R20716 XThC.Tn[2].n34 XThC.Tn[2].t25 145.137
R20717 XThC.Tn[2].n37 XThC.Tn[2].t13 145.137
R20718 XThC.Tn[2].n40 XThC.Tn[2].t15 145.137
R20719 XThC.Tn[2].n43 XThC.Tn[2].t26 145.137
R20720 XThC.Tn[2].n46 XThC.Tn[2].t34 145.137
R20721 XThC.Tn[2].n49 XThC.Tn[2].t36 145.137
R20722 XThC.Tn[2].n52 XThC.Tn[2].t17 145.137
R20723 XThC.Tn[2].n55 XThC.Tn[2].t27 145.137
R20724 XThC.Tn[2].n7 XThC.Tn[2].n6 135.248
R20725 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R20726 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R20727 XThC.Tn[2].n7 XThC.Tn[2].n5 98.982
R20728 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R20729 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R20730 XThC.Tn[2].n59 XThC.Tn[2].n9 32.6405
R20731 XThC.Tn[2].n1 XThC.Tn[2].t8 26.5955
R20732 XThC.Tn[2].n1 XThC.Tn[2].t7 26.5955
R20733 XThC.Tn[2].n0 XThC.Tn[2].t10 26.5955
R20734 XThC.Tn[2].n0 XThC.Tn[2].t9 26.5955
R20735 XThC.Tn[2].n3 XThC.Tn[2].t6 24.9236
R20736 XThC.Tn[2].n3 XThC.Tn[2].t5 24.9236
R20737 XThC.Tn[2].n4 XThC.Tn[2].t4 24.9236
R20738 XThC.Tn[2].n4 XThC.Tn[2].t3 24.9236
R20739 XThC.Tn[2].n5 XThC.Tn[2].t1 24.9236
R20740 XThC.Tn[2].n5 XThC.Tn[2].t2 24.9236
R20741 XThC.Tn[2].n6 XThC.Tn[2].t11 24.9236
R20742 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R20743 XThC.Tn[2].n60 XThC.Tn[2].n2 18.5605
R20744 XThC.Tn[2].n60 XThC.Tn[2].n59 11.5205
R20745 XThC.Tn[2].n58 XThC.Tn[2] 6.32799
R20746 XThC.Tn[2].n59 XThC.Tn[2].n58 3.18175
R20747 XThC.Tn[2].n15 XThC.Tn[2] 0.931056
R20748 XThC.Tn[2].n18 XThC.Tn[2] 0.931056
R20749 XThC.Tn[2].n21 XThC.Tn[2] 0.931056
R20750 XThC.Tn[2].n24 XThC.Tn[2] 0.931056
R20751 XThC.Tn[2].n27 XThC.Tn[2] 0.931056
R20752 XThC.Tn[2].n30 XThC.Tn[2] 0.931056
R20753 XThC.Tn[2].n33 XThC.Tn[2] 0.931056
R20754 XThC.Tn[2].n36 XThC.Tn[2] 0.931056
R20755 XThC.Tn[2].n39 XThC.Tn[2] 0.931056
R20756 XThC.Tn[2].n42 XThC.Tn[2] 0.931056
R20757 XThC.Tn[2].n45 XThC.Tn[2] 0.931056
R20758 XThC.Tn[2].n48 XThC.Tn[2] 0.931056
R20759 XThC.Tn[2].n51 XThC.Tn[2] 0.931056
R20760 XThC.Tn[2].n54 XThC.Tn[2] 0.931056
R20761 XThC.Tn[2].n57 XThC.Tn[2] 0.931056
R20762 XThC.Tn[2] XThC.Tn[2].n60 0.6405
R20763 XThC.Tn[2] XThC.Tn[2].n12 0.396333
R20764 XThC.Tn[2] XThC.Tn[2].n15 0.396333
R20765 XThC.Tn[2] XThC.Tn[2].n18 0.396333
R20766 XThC.Tn[2] XThC.Tn[2].n21 0.396333
R20767 XThC.Tn[2] XThC.Tn[2].n24 0.396333
R20768 XThC.Tn[2] XThC.Tn[2].n27 0.396333
R20769 XThC.Tn[2] XThC.Tn[2].n30 0.396333
R20770 XThC.Tn[2] XThC.Tn[2].n33 0.396333
R20771 XThC.Tn[2] XThC.Tn[2].n36 0.396333
R20772 XThC.Tn[2] XThC.Tn[2].n39 0.396333
R20773 XThC.Tn[2] XThC.Tn[2].n42 0.396333
R20774 XThC.Tn[2] XThC.Tn[2].n45 0.396333
R20775 XThC.Tn[2] XThC.Tn[2].n48 0.396333
R20776 XThC.Tn[2] XThC.Tn[2].n51 0.396333
R20777 XThC.Tn[2] XThC.Tn[2].n54 0.396333
R20778 XThC.Tn[2] XThC.Tn[2].n57 0.396333
R20779 XThC.Tn[2].n11 XThC.Tn[2] 0.104667
R20780 XThC.Tn[2].n14 XThC.Tn[2] 0.104667
R20781 XThC.Tn[2].n17 XThC.Tn[2] 0.104667
R20782 XThC.Tn[2].n20 XThC.Tn[2] 0.104667
R20783 XThC.Tn[2].n23 XThC.Tn[2] 0.104667
R20784 XThC.Tn[2].n26 XThC.Tn[2] 0.104667
R20785 XThC.Tn[2].n29 XThC.Tn[2] 0.104667
R20786 XThC.Tn[2].n32 XThC.Tn[2] 0.104667
R20787 XThC.Tn[2].n35 XThC.Tn[2] 0.104667
R20788 XThC.Tn[2].n38 XThC.Tn[2] 0.104667
R20789 XThC.Tn[2].n41 XThC.Tn[2] 0.104667
R20790 XThC.Tn[2].n44 XThC.Tn[2] 0.104667
R20791 XThC.Tn[2].n47 XThC.Tn[2] 0.104667
R20792 XThC.Tn[2].n50 XThC.Tn[2] 0.104667
R20793 XThC.Tn[2].n53 XThC.Tn[2] 0.104667
R20794 XThC.Tn[2].n56 XThC.Tn[2] 0.104667
R20795 XThC.Tn[2].n11 XThC.Tn[2] 0.0309878
R20796 XThC.Tn[2].n14 XThC.Tn[2] 0.0309878
R20797 XThC.Tn[2].n17 XThC.Tn[2] 0.0309878
R20798 XThC.Tn[2].n20 XThC.Tn[2] 0.0309878
R20799 XThC.Tn[2].n23 XThC.Tn[2] 0.0309878
R20800 XThC.Tn[2].n26 XThC.Tn[2] 0.0309878
R20801 XThC.Tn[2].n29 XThC.Tn[2] 0.0309878
R20802 XThC.Tn[2].n32 XThC.Tn[2] 0.0309878
R20803 XThC.Tn[2].n35 XThC.Tn[2] 0.0309878
R20804 XThC.Tn[2].n38 XThC.Tn[2] 0.0309878
R20805 XThC.Tn[2].n41 XThC.Tn[2] 0.0309878
R20806 XThC.Tn[2].n44 XThC.Tn[2] 0.0309878
R20807 XThC.Tn[2].n47 XThC.Tn[2] 0.0309878
R20808 XThC.Tn[2].n50 XThC.Tn[2] 0.0309878
R20809 XThC.Tn[2].n53 XThC.Tn[2] 0.0309878
R20810 XThC.Tn[2].n56 XThC.Tn[2] 0.0309878
R20811 XThC.Tn[2].n12 XThC.Tn[2].n11 0.027939
R20812 XThC.Tn[2].n15 XThC.Tn[2].n14 0.027939
R20813 XThC.Tn[2].n18 XThC.Tn[2].n17 0.027939
R20814 XThC.Tn[2].n21 XThC.Tn[2].n20 0.027939
R20815 XThC.Tn[2].n24 XThC.Tn[2].n23 0.027939
R20816 XThC.Tn[2].n27 XThC.Tn[2].n26 0.027939
R20817 XThC.Tn[2].n30 XThC.Tn[2].n29 0.027939
R20818 XThC.Tn[2].n33 XThC.Tn[2].n32 0.027939
R20819 XThC.Tn[2].n36 XThC.Tn[2].n35 0.027939
R20820 XThC.Tn[2].n39 XThC.Tn[2].n38 0.027939
R20821 XThC.Tn[2].n42 XThC.Tn[2].n41 0.027939
R20822 XThC.Tn[2].n45 XThC.Tn[2].n44 0.027939
R20823 XThC.Tn[2].n48 XThC.Tn[2].n47 0.027939
R20824 XThC.Tn[2].n51 XThC.Tn[2].n50 0.027939
R20825 XThC.Tn[2].n54 XThC.Tn[2].n53 0.027939
R20826 XThC.Tn[2].n57 XThC.Tn[2].n56 0.027939
R20827 XThC.Tn[2].n58 XThC.Tn[2] 0.0156819
R20828 Vbias.t4 Vbias.n512 313.474
R20829 Vbias.t6 Vbias.n518 313.464
R20830 Vbias.n516 Vbias.t4 313.13
R20831 Vbias.n522 Vbias.t6 313.13
R20832 Vbias.n515 Vbias.n514 299.471
R20833 Vbias.n521 Vbias.n520 299.471
R20834 Vbias.n515 Vbias.n513 299.144
R20835 Vbias.n521 Vbias.n519 299.144
R20836 Vbias.n509 Vbias.t187 119.309
R20837 Vbias.n507 Vbias.t30 119.309
R20838 Vbias.n505 Vbias.t18 119.309
R20839 Vbias.n503 Vbias.t254 119.309
R20840 Vbias.n501 Vbias.t101 119.309
R20841 Vbias.n499 Vbias.t81 119.309
R20842 Vbias.n497 Vbias.t252 119.309
R20843 Vbias.n495 Vbias.t175 119.309
R20844 Vbias.n493 Vbias.t153 119.309
R20845 Vbias.n491 Vbias.t66 119.309
R20846 Vbias.n489 Vbias.t233 119.309
R20847 Vbias.n487 Vbias.t147 119.309
R20848 Vbias.n485 Vbias.t62 119.309
R20849 Vbias.n483 Vbias.t47 119.309
R20850 Vbias.n481 Vbias.t207 119.309
R20851 Vbias.n480 Vbias.t135 119.309
R20852 Vbias.n477 Vbias.t116 119.309
R20853 Vbias.n475 Vbias.t216 119.309
R20854 Vbias.n473 Vbias.t199 119.309
R20855 Vbias.n471 Vbias.t179 119.309
R20856 Vbias.n469 Vbias.t31 119.309
R20857 Vbias.n467 Vbias.t264 119.309
R20858 Vbias.n465 Vbias.t177 119.309
R20859 Vbias.n463 Vbias.t102 119.309
R20860 Vbias.n461 Vbias.t82 119.309
R20861 Vbias.n459 Vbias.t253 119.309
R20862 Vbias.n457 Vbias.t162 119.309
R20863 Vbias.n455 Vbias.t75 119.309
R20864 Vbias.n453 Vbias.t248 119.309
R20865 Vbias.n451 Vbias.t235 119.309
R20866 Vbias.n449 Vbias.t136 119.309
R20867 Vbias.n448 Vbias.t63 119.309
R20868 Vbias.n445 Vbias.t152 119.309
R20869 Vbias.n443 Vbias.t244 119.309
R20870 Vbias.n441 Vbias.t231 119.309
R20871 Vbias.n439 Vbias.t211 119.309
R20872 Vbias.n437 Vbias.t58 119.309
R20873 Vbias.n435 Vbias.t38 119.309
R20874 Vbias.n433 Vbias.t205 119.309
R20875 Vbias.n431 Vbias.t131 119.309
R20876 Vbias.n429 Vbias.t108 119.309
R20877 Vbias.n427 Vbias.t24 119.309
R20878 Vbias.n425 Vbias.t189 119.309
R20879 Vbias.n423 Vbias.t105 119.309
R20880 Vbias.n421 Vbias.t20 119.309
R20881 Vbias.n419 Vbias.t267 119.309
R20882 Vbias.n417 Vbias.t166 119.309
R20883 Vbias.n416 Vbias.t93 119.309
R20884 Vbias.n413 Vbias.t79 119.309
R20885 Vbias.n411 Vbias.t171 119.309
R20886 Vbias.n409 Vbias.t159 119.309
R20887 Vbias.n407 Vbias.t139 119.309
R20888 Vbias.n405 Vbias.t245 119.309
R20889 Vbias.n403 Vbias.t223 119.309
R20890 Vbias.n401 Vbias.t132 119.309
R20891 Vbias.n399 Vbias.t59 119.309
R20892 Vbias.n397 Vbias.t39 119.309
R20893 Vbias.n395 Vbias.t206 119.309
R20894 Vbias.n393 Vbias.t118 119.309
R20895 Vbias.n391 Vbias.t35 119.309
R20896 Vbias.n389 Vbias.t202 119.309
R20897 Vbias.n387 Vbias.t191 119.309
R20898 Vbias.n385 Vbias.t94 119.309
R20899 Vbias.n384 Vbias.t22 119.309
R20900 Vbias.n381 Vbias.t261 119.309
R20901 Vbias.n379 Vbias.t98 119.309
R20902 Vbias.n377 Vbias.t87 119.309
R20903 Vbias.n375 Vbias.t68 119.309
R20904 Vbias.n373 Vbias.t172 119.309
R20905 Vbias.n371 Vbias.t150 119.309
R20906 Vbias.n369 Vbias.t60 119.309
R20907 Vbias.n367 Vbias.t246 119.309
R20908 Vbias.n365 Vbias.t225 119.309
R20909 Vbias.n363 Vbias.t133 119.309
R20910 Vbias.n361 Vbias.t46 119.309
R20911 Vbias.n359 Vbias.t219 119.309
R20912 Vbias.n357 Vbias.t130 119.309
R20913 Vbias.n355 Vbias.t119 119.309
R20914 Vbias.n353 Vbias.t23 119.309
R20915 Vbias.n352 Vbias.t204 119.309
R20916 Vbias.n349 Vbias.t182 119.309
R20917 Vbias.n347 Vbias.t26 119.309
R20918 Vbias.n345 Vbias.t13 119.309
R20919 Vbias.n343 Vbias.t249 119.309
R20920 Vbias.n341 Vbias.t96 119.309
R20921 Vbias.n339 Vbias.t71 119.309
R20922 Vbias.n337 Vbias.t242 119.309
R20923 Vbias.n335 Vbias.t169 119.309
R20924 Vbias.n333 Vbias.t144 119.309
R20925 Vbias.n331 Vbias.t56 119.309
R20926 Vbias.n329 Vbias.t227 119.309
R20927 Vbias.n327 Vbias.t141 119.309
R20928 Vbias.n325 Vbias.t54 119.309
R20929 Vbias.n323 Vbias.t43 119.309
R20930 Vbias.n321 Vbias.t201 119.309
R20931 Vbias.n320 Vbias.t127 119.309
R20932 Vbias.n317 Vbias.t111 119.309
R20933 Vbias.n315 Vbias.t210 119.309
R20934 Vbias.n313 Vbias.t193 119.309
R20935 Vbias.n311 Vbias.t174 119.309
R20936 Vbias.n309 Vbias.t27 119.309
R20937 Vbias.n307 Vbias.t257 119.309
R20938 Vbias.n305 Vbias.t170 119.309
R20939 Vbias.n303 Vbias.t97 119.309
R20940 Vbias.n301 Vbias.t74 119.309
R20941 Vbias.n299 Vbias.t243 119.309
R20942 Vbias.n297 Vbias.t156 119.309
R20943 Vbias.n295 Vbias.t69 119.309
R20944 Vbias.n293 Vbias.t241 119.309
R20945 Vbias.n291 Vbias.t228 119.309
R20946 Vbias.n289 Vbias.t128 119.309
R20947 Vbias.n288 Vbias.t55 119.309
R20948 Vbias.n285 Vbias.t143 119.309
R20949 Vbias.n283 Vbias.t238 119.309
R20950 Vbias.n281 Vbias.t226 119.309
R20951 Vbias.n279 Vbias.t203 119.309
R20952 Vbias.n277 Vbias.t50 119.309
R20953 Vbias.n275 Vbias.t33 119.309
R20954 Vbias.n273 Vbias.t196 119.309
R20955 Vbias.n271 Vbias.t124 119.309
R20956 Vbias.n269 Vbias.t104 119.309
R20957 Vbias.n267 Vbias.t17 119.309
R20958 Vbias.n265 Vbias.t185 119.309
R20959 Vbias.n263 Vbias.t99 119.309
R20960 Vbias.n261 Vbias.t14 119.309
R20961 Vbias.n259 Vbias.t263 119.309
R20962 Vbias.n257 Vbias.t160 119.309
R20963 Vbias.n256 Vbias.t88 119.309
R20964 Vbias.n253 Vbias.t70 119.309
R20965 Vbias.n251 Vbias.t167 119.309
R20966 Vbias.n249 Vbias.t155 119.309
R20967 Vbias.n247 Vbias.t129 119.309
R20968 Vbias.n245 Vbias.t239 119.309
R20969 Vbias.n243 Vbias.t217 119.309
R20970 Vbias.n241 Vbias.t125 119.309
R20971 Vbias.n239 Vbias.t51 119.309
R20972 Vbias.n237 Vbias.t34 119.309
R20973 Vbias.n235 Vbias.t198 119.309
R20974 Vbias.n233 Vbias.t113 119.309
R20975 Vbias.n231 Vbias.t29 119.309
R20976 Vbias.n229 Vbias.t194 119.309
R20977 Vbias.n227 Vbias.t186 119.309
R20978 Vbias.n225 Vbias.t89 119.309
R20979 Vbias.n224 Vbias.t15 119.309
R20980 Vbias.n221 Vbias.t256 119.309
R20981 Vbias.n219 Vbias.t95 119.309
R20982 Vbias.n217 Vbias.t86 119.309
R20983 Vbias.n215 Vbias.t57 119.309
R20984 Vbias.n213 Vbias.t168 119.309
R20985 Vbias.n211 Vbias.t142 119.309
R20986 Vbias.n209 Vbias.t52 119.309
R20987 Vbias.n207 Vbias.t240 119.309
R20988 Vbias.n205 Vbias.t218 119.309
R20989 Vbias.n203 Vbias.t126 119.309
R20990 Vbias.n201 Vbias.t42 119.309
R20991 Vbias.n199 Vbias.t214 119.309
R20992 Vbias.n197 Vbias.t123 119.309
R20993 Vbias.n195 Vbias.t114 119.309
R20994 Vbias.n193 Vbias.t16 119.309
R20995 Vbias.n192 Vbias.t195 119.309
R20996 Vbias.n189 Vbias.t115 119.309
R20997 Vbias.n187 Vbias.t213 119.309
R20998 Vbias.n185 Vbias.t197 119.309
R20999 Vbias.n183 Vbias.t178 119.309
R21000 Vbias.n181 Vbias.t28 119.309
R21001 Vbias.n179 Vbias.t262 119.309
R21002 Vbias.n177 Vbias.t173 119.309
R21003 Vbias.n175 Vbias.t100 119.309
R21004 Vbias.n173 Vbias.t80 119.309
R21005 Vbias.n171 Vbias.t250 119.309
R21006 Vbias.n169 Vbias.t161 119.309
R21007 Vbias.n167 Vbias.t72 119.309
R21008 Vbias.n165 Vbias.t247 119.309
R21009 Vbias.n163 Vbias.t232 119.309
R21010 Vbias.n161 Vbias.t134 119.309
R21011 Vbias.n160 Vbias.t61 119.309
R21012 Vbias.n157 Vbias.t255 119.309
R21013 Vbias.n155 Vbias.t91 119.309
R21014 Vbias.n153 Vbias.t84 119.309
R21015 Vbias.n151 Vbias.t53 119.309
R21016 Vbias.n149 Vbias.t165 119.309
R21017 Vbias.n147 Vbias.t140 119.309
R21018 Vbias.n145 Vbias.t49 119.309
R21019 Vbias.n143 Vbias.t237 119.309
R21020 Vbias.n141 Vbias.t215 119.309
R21021 Vbias.n139 Vbias.t122 119.309
R21022 Vbias.n137 Vbias.t40 119.309
R21023 Vbias.n135 Vbias.t212 119.309
R21024 Vbias.n133 Vbias.t121 119.309
R21025 Vbias.n131 Vbias.t109 119.309
R21026 Vbias.n129 Vbias.t12 119.309
R21027 Vbias.n128 Vbias.t192 119.309
R21028 Vbias.n125 Vbias.t92 119.309
R21029 Vbias.n123 Vbias.t181 119.309
R21030 Vbias.n121 Vbias.t176 119.309
R21031 Vbias.n119 Vbias.t154 119.309
R21032 Vbias.n117 Vbias.t258 119.309
R21033 Vbias.n115 Vbias.t234 119.309
R21034 Vbias.n113 Vbias.t149 119.309
R21035 Vbias.n111 Vbias.t76 119.309
R21036 Vbias.n109 Vbias.t48 119.309
R21037 Vbias.n107 Vbias.t224 119.309
R21038 Vbias.n105 Vbias.t137 119.309
R21039 Vbias.n103 Vbias.t44 119.309
R21040 Vbias.n101 Vbias.t220 119.309
R21041 Vbias.n99 Vbias.t209 119.309
R21042 Vbias.n97 Vbias.t106 119.309
R21043 Vbias.n96 Vbias.t36 119.309
R21044 Vbias.n93 Vbias.t19 119.309
R21045 Vbias.n91 Vbias.t110 119.309
R21046 Vbias.n89 Vbias.t103 119.309
R21047 Vbias.n87 Vbias.t83 119.309
R21048 Vbias.n85 Vbias.t183 119.309
R21049 Vbias.n83 Vbias.t163 119.309
R21050 Vbias.n81 Vbias.t77 119.309
R21051 Vbias.n79 Vbias.t259 119.309
R21052 Vbias.n77 Vbias.t236 119.309
R21053 Vbias.n75 Vbias.t151 119.309
R21054 Vbias.n73 Vbias.t64 119.309
R21055 Vbias.n71 Vbias.t230 119.309
R21056 Vbias.n69 Vbias.t145 119.309
R21057 Vbias.n67 Vbias.t138 119.309
R21058 Vbias.n65 Vbias.t37 119.309
R21059 Vbias.n64 Vbias.t221 119.309
R21060 Vbias.n61 Vbias.t200 119.309
R21061 Vbias.n59 Vbias.t41 119.309
R21062 Vbias.n57 Vbias.t32 119.309
R21063 Vbias.n55 Vbias.t265 119.309
R21064 Vbias.n53 Vbias.t112 119.309
R21065 Vbias.n51 Vbias.t90 119.309
R21066 Vbias.n49 Vbias.t260 119.309
R21067 Vbias.n47 Vbias.t184 119.309
R21068 Vbias.n45 Vbias.t164 119.309
R21069 Vbias.n43 Vbias.t78 119.309
R21070 Vbias.n41 Vbias.t251 119.309
R21071 Vbias.n39 Vbias.t158 119.309
R21072 Vbias.n37 Vbias.t73 119.309
R21073 Vbias.n35 Vbias.t65 119.309
R21074 Vbias.n33 Vbias.t222 119.309
R21075 Vbias.n32 Vbias.t146 119.309
R21076 Vbias.n29 Vbias.t67 119.309
R21077 Vbias.n27 Vbias.t157 119.309
R21078 Vbias.n25 Vbias.t148 119.309
R21079 Vbias.n23 Vbias.t120 119.309
R21080 Vbias.n21 Vbias.t229 119.309
R21081 Vbias.n19 Vbias.t208 119.309
R21082 Vbias.n17 Vbias.t117 119.309
R21083 Vbias.n15 Vbias.t45 119.309
R21084 Vbias.n13 Vbias.t25 119.309
R21085 Vbias.n11 Vbias.t190 119.309
R21086 Vbias.n9 Vbias.t107 119.309
R21087 Vbias.n7 Vbias.t21 119.309
R21088 Vbias.n5 Vbias.t188 119.309
R21089 Vbias.n3 Vbias.t180 119.309
R21090 Vbias.n1 Vbias.t85 119.309
R21091 Vbias.n0 Vbias.t266 119.309
R21092 Vbias.n513 Vbias.t8 53.3064
R21093 Vbias.n513 Vbias.t3 53.3064
R21094 Vbias.n519 Vbias.t10 53.3064
R21095 Vbias.n519 Vbias.t11 53.3064
R21096 Vbias.n512 Vbias.t5 34.1153
R21097 Vbias.n518 Vbias.t7 34.1153
R21098 Vbias.n514 Vbias.t2 33.6064
R21099 Vbias.n514 Vbias.t9 33.6064
R21100 Vbias.n520 Vbias.t1 33.6064
R21101 Vbias.n520 Vbias.t0 33.6064
R21102 Vbias Vbias.n480 8.00727
R21103 Vbias Vbias.n448 8.00727
R21104 Vbias Vbias.n416 8.00727
R21105 Vbias Vbias.n384 8.00727
R21106 Vbias Vbias.n352 8.00727
R21107 Vbias Vbias.n320 8.00727
R21108 Vbias Vbias.n288 8.00727
R21109 Vbias Vbias.n256 8.00727
R21110 Vbias Vbias.n224 8.00727
R21111 Vbias Vbias.n192 8.00727
R21112 Vbias Vbias.n160 8.00727
R21113 Vbias Vbias.n128 8.00727
R21114 Vbias Vbias.n96 8.00727
R21115 Vbias Vbias.n64 8.00727
R21116 Vbias Vbias.n32 8.00727
R21117 Vbias Vbias.n0 8.00727
R21118 Vbias.n510 Vbias.n509 7.9105
R21119 Vbias.n508 Vbias.n507 7.9105
R21120 Vbias.n506 Vbias.n505 7.9105
R21121 Vbias.n504 Vbias.n503 7.9105
R21122 Vbias.n502 Vbias.n501 7.9105
R21123 Vbias.n500 Vbias.n499 7.9105
R21124 Vbias.n498 Vbias.n497 7.9105
R21125 Vbias.n496 Vbias.n495 7.9105
R21126 Vbias.n494 Vbias.n493 7.9105
R21127 Vbias.n492 Vbias.n491 7.9105
R21128 Vbias.n490 Vbias.n489 7.9105
R21129 Vbias.n488 Vbias.n487 7.9105
R21130 Vbias.n486 Vbias.n485 7.9105
R21131 Vbias.n484 Vbias.n483 7.9105
R21132 Vbias.n482 Vbias.n481 7.9105
R21133 Vbias.n478 Vbias.n477 7.9105
R21134 Vbias.n476 Vbias.n475 7.9105
R21135 Vbias.n474 Vbias.n473 7.9105
R21136 Vbias.n472 Vbias.n471 7.9105
R21137 Vbias.n470 Vbias.n469 7.9105
R21138 Vbias.n468 Vbias.n467 7.9105
R21139 Vbias.n466 Vbias.n465 7.9105
R21140 Vbias.n464 Vbias.n463 7.9105
R21141 Vbias.n462 Vbias.n461 7.9105
R21142 Vbias.n460 Vbias.n459 7.9105
R21143 Vbias.n458 Vbias.n457 7.9105
R21144 Vbias.n456 Vbias.n455 7.9105
R21145 Vbias.n454 Vbias.n453 7.9105
R21146 Vbias.n452 Vbias.n451 7.9105
R21147 Vbias.n450 Vbias.n449 7.9105
R21148 Vbias.n446 Vbias.n445 7.9105
R21149 Vbias.n444 Vbias.n443 7.9105
R21150 Vbias.n442 Vbias.n441 7.9105
R21151 Vbias.n440 Vbias.n439 7.9105
R21152 Vbias.n438 Vbias.n437 7.9105
R21153 Vbias.n436 Vbias.n435 7.9105
R21154 Vbias.n434 Vbias.n433 7.9105
R21155 Vbias.n432 Vbias.n431 7.9105
R21156 Vbias.n430 Vbias.n429 7.9105
R21157 Vbias.n428 Vbias.n427 7.9105
R21158 Vbias.n426 Vbias.n425 7.9105
R21159 Vbias.n424 Vbias.n423 7.9105
R21160 Vbias.n422 Vbias.n421 7.9105
R21161 Vbias.n420 Vbias.n419 7.9105
R21162 Vbias.n418 Vbias.n417 7.9105
R21163 Vbias.n414 Vbias.n413 7.9105
R21164 Vbias.n412 Vbias.n411 7.9105
R21165 Vbias.n410 Vbias.n409 7.9105
R21166 Vbias.n408 Vbias.n407 7.9105
R21167 Vbias.n406 Vbias.n405 7.9105
R21168 Vbias.n404 Vbias.n403 7.9105
R21169 Vbias.n402 Vbias.n401 7.9105
R21170 Vbias.n400 Vbias.n399 7.9105
R21171 Vbias.n398 Vbias.n397 7.9105
R21172 Vbias.n396 Vbias.n395 7.9105
R21173 Vbias.n394 Vbias.n393 7.9105
R21174 Vbias.n392 Vbias.n391 7.9105
R21175 Vbias.n390 Vbias.n389 7.9105
R21176 Vbias.n388 Vbias.n387 7.9105
R21177 Vbias.n386 Vbias.n385 7.9105
R21178 Vbias.n382 Vbias.n381 7.9105
R21179 Vbias.n380 Vbias.n379 7.9105
R21180 Vbias.n378 Vbias.n377 7.9105
R21181 Vbias.n376 Vbias.n375 7.9105
R21182 Vbias.n374 Vbias.n373 7.9105
R21183 Vbias.n372 Vbias.n371 7.9105
R21184 Vbias.n370 Vbias.n369 7.9105
R21185 Vbias.n368 Vbias.n367 7.9105
R21186 Vbias.n366 Vbias.n365 7.9105
R21187 Vbias.n364 Vbias.n363 7.9105
R21188 Vbias.n362 Vbias.n361 7.9105
R21189 Vbias.n360 Vbias.n359 7.9105
R21190 Vbias.n358 Vbias.n357 7.9105
R21191 Vbias.n356 Vbias.n355 7.9105
R21192 Vbias.n354 Vbias.n353 7.9105
R21193 Vbias.n350 Vbias.n349 7.9105
R21194 Vbias.n348 Vbias.n347 7.9105
R21195 Vbias.n346 Vbias.n345 7.9105
R21196 Vbias.n344 Vbias.n343 7.9105
R21197 Vbias.n342 Vbias.n341 7.9105
R21198 Vbias.n340 Vbias.n339 7.9105
R21199 Vbias.n338 Vbias.n337 7.9105
R21200 Vbias.n336 Vbias.n335 7.9105
R21201 Vbias.n334 Vbias.n333 7.9105
R21202 Vbias.n332 Vbias.n331 7.9105
R21203 Vbias.n330 Vbias.n329 7.9105
R21204 Vbias.n328 Vbias.n327 7.9105
R21205 Vbias.n326 Vbias.n325 7.9105
R21206 Vbias.n324 Vbias.n323 7.9105
R21207 Vbias.n322 Vbias.n321 7.9105
R21208 Vbias.n318 Vbias.n317 7.9105
R21209 Vbias.n316 Vbias.n315 7.9105
R21210 Vbias.n314 Vbias.n313 7.9105
R21211 Vbias.n312 Vbias.n311 7.9105
R21212 Vbias.n310 Vbias.n309 7.9105
R21213 Vbias.n308 Vbias.n307 7.9105
R21214 Vbias.n306 Vbias.n305 7.9105
R21215 Vbias.n304 Vbias.n303 7.9105
R21216 Vbias.n302 Vbias.n301 7.9105
R21217 Vbias.n300 Vbias.n299 7.9105
R21218 Vbias.n298 Vbias.n297 7.9105
R21219 Vbias.n296 Vbias.n295 7.9105
R21220 Vbias.n294 Vbias.n293 7.9105
R21221 Vbias.n292 Vbias.n291 7.9105
R21222 Vbias.n290 Vbias.n289 7.9105
R21223 Vbias.n286 Vbias.n285 7.9105
R21224 Vbias.n284 Vbias.n283 7.9105
R21225 Vbias.n282 Vbias.n281 7.9105
R21226 Vbias.n280 Vbias.n279 7.9105
R21227 Vbias.n278 Vbias.n277 7.9105
R21228 Vbias.n276 Vbias.n275 7.9105
R21229 Vbias.n274 Vbias.n273 7.9105
R21230 Vbias.n272 Vbias.n271 7.9105
R21231 Vbias.n270 Vbias.n269 7.9105
R21232 Vbias.n268 Vbias.n267 7.9105
R21233 Vbias.n266 Vbias.n265 7.9105
R21234 Vbias.n264 Vbias.n263 7.9105
R21235 Vbias.n262 Vbias.n261 7.9105
R21236 Vbias.n260 Vbias.n259 7.9105
R21237 Vbias.n258 Vbias.n257 7.9105
R21238 Vbias.n254 Vbias.n253 7.9105
R21239 Vbias.n252 Vbias.n251 7.9105
R21240 Vbias.n250 Vbias.n249 7.9105
R21241 Vbias.n248 Vbias.n247 7.9105
R21242 Vbias.n246 Vbias.n245 7.9105
R21243 Vbias.n244 Vbias.n243 7.9105
R21244 Vbias.n242 Vbias.n241 7.9105
R21245 Vbias.n240 Vbias.n239 7.9105
R21246 Vbias.n238 Vbias.n237 7.9105
R21247 Vbias.n236 Vbias.n235 7.9105
R21248 Vbias.n234 Vbias.n233 7.9105
R21249 Vbias.n232 Vbias.n231 7.9105
R21250 Vbias.n230 Vbias.n229 7.9105
R21251 Vbias.n228 Vbias.n227 7.9105
R21252 Vbias.n226 Vbias.n225 7.9105
R21253 Vbias.n222 Vbias.n221 7.9105
R21254 Vbias.n220 Vbias.n219 7.9105
R21255 Vbias.n218 Vbias.n217 7.9105
R21256 Vbias.n216 Vbias.n215 7.9105
R21257 Vbias.n214 Vbias.n213 7.9105
R21258 Vbias.n212 Vbias.n211 7.9105
R21259 Vbias.n210 Vbias.n209 7.9105
R21260 Vbias.n208 Vbias.n207 7.9105
R21261 Vbias.n206 Vbias.n205 7.9105
R21262 Vbias.n204 Vbias.n203 7.9105
R21263 Vbias.n202 Vbias.n201 7.9105
R21264 Vbias.n200 Vbias.n199 7.9105
R21265 Vbias.n198 Vbias.n197 7.9105
R21266 Vbias.n196 Vbias.n195 7.9105
R21267 Vbias.n194 Vbias.n193 7.9105
R21268 Vbias.n190 Vbias.n189 7.9105
R21269 Vbias.n188 Vbias.n187 7.9105
R21270 Vbias.n186 Vbias.n185 7.9105
R21271 Vbias.n184 Vbias.n183 7.9105
R21272 Vbias.n182 Vbias.n181 7.9105
R21273 Vbias.n180 Vbias.n179 7.9105
R21274 Vbias.n178 Vbias.n177 7.9105
R21275 Vbias.n176 Vbias.n175 7.9105
R21276 Vbias.n174 Vbias.n173 7.9105
R21277 Vbias.n172 Vbias.n171 7.9105
R21278 Vbias.n170 Vbias.n169 7.9105
R21279 Vbias.n168 Vbias.n167 7.9105
R21280 Vbias.n166 Vbias.n165 7.9105
R21281 Vbias.n164 Vbias.n163 7.9105
R21282 Vbias.n162 Vbias.n161 7.9105
R21283 Vbias.n158 Vbias.n157 7.9105
R21284 Vbias.n156 Vbias.n155 7.9105
R21285 Vbias.n154 Vbias.n153 7.9105
R21286 Vbias.n152 Vbias.n151 7.9105
R21287 Vbias.n150 Vbias.n149 7.9105
R21288 Vbias.n148 Vbias.n147 7.9105
R21289 Vbias.n146 Vbias.n145 7.9105
R21290 Vbias.n144 Vbias.n143 7.9105
R21291 Vbias.n142 Vbias.n141 7.9105
R21292 Vbias.n140 Vbias.n139 7.9105
R21293 Vbias.n138 Vbias.n137 7.9105
R21294 Vbias.n136 Vbias.n135 7.9105
R21295 Vbias.n134 Vbias.n133 7.9105
R21296 Vbias.n132 Vbias.n131 7.9105
R21297 Vbias.n130 Vbias.n129 7.9105
R21298 Vbias.n126 Vbias.n125 7.9105
R21299 Vbias.n124 Vbias.n123 7.9105
R21300 Vbias.n122 Vbias.n121 7.9105
R21301 Vbias.n120 Vbias.n119 7.9105
R21302 Vbias.n118 Vbias.n117 7.9105
R21303 Vbias.n116 Vbias.n115 7.9105
R21304 Vbias.n114 Vbias.n113 7.9105
R21305 Vbias.n112 Vbias.n111 7.9105
R21306 Vbias.n110 Vbias.n109 7.9105
R21307 Vbias.n108 Vbias.n107 7.9105
R21308 Vbias.n106 Vbias.n105 7.9105
R21309 Vbias.n104 Vbias.n103 7.9105
R21310 Vbias.n102 Vbias.n101 7.9105
R21311 Vbias.n100 Vbias.n99 7.9105
R21312 Vbias.n98 Vbias.n97 7.9105
R21313 Vbias.n94 Vbias.n93 7.9105
R21314 Vbias.n92 Vbias.n91 7.9105
R21315 Vbias.n90 Vbias.n89 7.9105
R21316 Vbias.n88 Vbias.n87 7.9105
R21317 Vbias.n86 Vbias.n85 7.9105
R21318 Vbias.n84 Vbias.n83 7.9105
R21319 Vbias.n82 Vbias.n81 7.9105
R21320 Vbias.n80 Vbias.n79 7.9105
R21321 Vbias.n78 Vbias.n77 7.9105
R21322 Vbias.n76 Vbias.n75 7.9105
R21323 Vbias.n74 Vbias.n73 7.9105
R21324 Vbias.n72 Vbias.n71 7.9105
R21325 Vbias.n70 Vbias.n69 7.9105
R21326 Vbias.n68 Vbias.n67 7.9105
R21327 Vbias.n66 Vbias.n65 7.9105
R21328 Vbias.n62 Vbias.n61 7.9105
R21329 Vbias.n60 Vbias.n59 7.9105
R21330 Vbias.n58 Vbias.n57 7.9105
R21331 Vbias.n56 Vbias.n55 7.9105
R21332 Vbias.n54 Vbias.n53 7.9105
R21333 Vbias.n52 Vbias.n51 7.9105
R21334 Vbias.n50 Vbias.n49 7.9105
R21335 Vbias.n48 Vbias.n47 7.9105
R21336 Vbias.n46 Vbias.n45 7.9105
R21337 Vbias.n44 Vbias.n43 7.9105
R21338 Vbias.n42 Vbias.n41 7.9105
R21339 Vbias.n40 Vbias.n39 7.9105
R21340 Vbias.n38 Vbias.n37 7.9105
R21341 Vbias.n36 Vbias.n35 7.9105
R21342 Vbias.n34 Vbias.n33 7.9105
R21343 Vbias.n30 Vbias.n29 7.9105
R21344 Vbias.n28 Vbias.n27 7.9105
R21345 Vbias.n26 Vbias.n25 7.9105
R21346 Vbias.n24 Vbias.n23 7.9105
R21347 Vbias.n22 Vbias.n21 7.9105
R21348 Vbias.n20 Vbias.n19 7.9105
R21349 Vbias.n18 Vbias.n17 7.9105
R21350 Vbias.n16 Vbias.n15 7.9105
R21351 Vbias.n14 Vbias.n13 7.9105
R21352 Vbias.n12 Vbias.n11 7.9105
R21353 Vbias.n10 Vbias.n9 7.9105
R21354 Vbias.n8 Vbias.n7 7.9105
R21355 Vbias.n6 Vbias.n5 7.9105
R21356 Vbias.n4 Vbias.n3 7.9105
R21357 Vbias.n2 Vbias.n1 7.9105
R21358 Vbias.n524 Vbias 6.41494
R21359 Vbias.n516 Vbias.n515 2.87046
R21360 Vbias.n522 Vbias.n521 2.87046
R21361 Vbias.n511 Vbias 1.6647
R21362 Vbias.n479 Vbias 1.6647
R21363 Vbias.n447 Vbias 1.6647
R21364 Vbias.n415 Vbias 1.6647
R21365 Vbias.n383 Vbias 1.6647
R21366 Vbias.n351 Vbias 1.6647
R21367 Vbias.n319 Vbias 1.6647
R21368 Vbias.n287 Vbias 1.6647
R21369 Vbias.n255 Vbias 1.6647
R21370 Vbias.n223 Vbias 1.6647
R21371 Vbias.n191 Vbias 1.6647
R21372 Vbias.n159 Vbias 1.6647
R21373 Vbias.n127 Vbias 1.6647
R21374 Vbias.n95 Vbias 1.6647
R21375 Vbias.n63 Vbias 1.6647
R21376 Vbias.n31 Vbias 1.6647
R21377 Vbias.n524 Vbias.n511 0.5692
R21378 Vbias.n63 Vbias.n31 0.410967
R21379 Vbias.n95 Vbias.n63 0.410967
R21380 Vbias.n127 Vbias.n95 0.410967
R21381 Vbias.n159 Vbias.n127 0.410967
R21382 Vbias.n191 Vbias.n159 0.410967
R21383 Vbias.n223 Vbias.n191 0.410967
R21384 Vbias.n255 Vbias.n223 0.410967
R21385 Vbias.n287 Vbias.n255 0.410967
R21386 Vbias.n319 Vbias.n287 0.410967
R21387 Vbias.n351 Vbias.n319 0.410967
R21388 Vbias.n383 Vbias.n351 0.410967
R21389 Vbias.n415 Vbias.n383 0.410967
R21390 Vbias.n447 Vbias.n415 0.410967
R21391 Vbias.n479 Vbias.n447 0.410967
R21392 Vbias.n511 Vbias.n479 0.410967
R21393 Vbias.n31 Vbias 0.383811
R21394 Vbias.n482 Vbias 0.252372
R21395 Vbias.n484 Vbias 0.252372
R21396 Vbias.n486 Vbias 0.252372
R21397 Vbias.n488 Vbias 0.252372
R21398 Vbias.n490 Vbias 0.252372
R21399 Vbias.n492 Vbias 0.252372
R21400 Vbias.n494 Vbias 0.252372
R21401 Vbias.n496 Vbias 0.252372
R21402 Vbias.n498 Vbias 0.252372
R21403 Vbias.n500 Vbias 0.252372
R21404 Vbias.n502 Vbias 0.252372
R21405 Vbias.n504 Vbias 0.252372
R21406 Vbias.n506 Vbias 0.252372
R21407 Vbias.n508 Vbias 0.252372
R21408 Vbias.n510 Vbias 0.252372
R21409 Vbias.n450 Vbias 0.252372
R21410 Vbias.n452 Vbias 0.252372
R21411 Vbias.n454 Vbias 0.252372
R21412 Vbias.n456 Vbias 0.252372
R21413 Vbias.n458 Vbias 0.252372
R21414 Vbias.n460 Vbias 0.252372
R21415 Vbias.n462 Vbias 0.252372
R21416 Vbias.n464 Vbias 0.252372
R21417 Vbias.n466 Vbias 0.252372
R21418 Vbias.n468 Vbias 0.252372
R21419 Vbias.n470 Vbias 0.252372
R21420 Vbias.n472 Vbias 0.252372
R21421 Vbias.n474 Vbias 0.252372
R21422 Vbias.n476 Vbias 0.252372
R21423 Vbias.n478 Vbias 0.252372
R21424 Vbias.n418 Vbias 0.252372
R21425 Vbias.n420 Vbias 0.252372
R21426 Vbias.n422 Vbias 0.252372
R21427 Vbias.n424 Vbias 0.252372
R21428 Vbias.n426 Vbias 0.252372
R21429 Vbias.n428 Vbias 0.252372
R21430 Vbias.n430 Vbias 0.252372
R21431 Vbias.n432 Vbias 0.252372
R21432 Vbias.n434 Vbias 0.252372
R21433 Vbias.n436 Vbias 0.252372
R21434 Vbias.n438 Vbias 0.252372
R21435 Vbias.n440 Vbias 0.252372
R21436 Vbias.n442 Vbias 0.252372
R21437 Vbias.n444 Vbias 0.252372
R21438 Vbias.n446 Vbias 0.252372
R21439 Vbias.n386 Vbias 0.252372
R21440 Vbias.n388 Vbias 0.252372
R21441 Vbias.n390 Vbias 0.252372
R21442 Vbias.n392 Vbias 0.252372
R21443 Vbias.n394 Vbias 0.252372
R21444 Vbias.n396 Vbias 0.252372
R21445 Vbias.n398 Vbias 0.252372
R21446 Vbias.n400 Vbias 0.252372
R21447 Vbias.n402 Vbias 0.252372
R21448 Vbias.n404 Vbias 0.252372
R21449 Vbias.n406 Vbias 0.252372
R21450 Vbias.n408 Vbias 0.252372
R21451 Vbias.n410 Vbias 0.252372
R21452 Vbias.n412 Vbias 0.252372
R21453 Vbias.n414 Vbias 0.252372
R21454 Vbias.n354 Vbias 0.252372
R21455 Vbias.n356 Vbias 0.252372
R21456 Vbias.n358 Vbias 0.252372
R21457 Vbias.n360 Vbias 0.252372
R21458 Vbias.n362 Vbias 0.252372
R21459 Vbias.n364 Vbias 0.252372
R21460 Vbias.n366 Vbias 0.252372
R21461 Vbias.n368 Vbias 0.252372
R21462 Vbias.n370 Vbias 0.252372
R21463 Vbias.n372 Vbias 0.252372
R21464 Vbias.n374 Vbias 0.252372
R21465 Vbias.n376 Vbias 0.252372
R21466 Vbias.n378 Vbias 0.252372
R21467 Vbias.n380 Vbias 0.252372
R21468 Vbias.n382 Vbias 0.252372
R21469 Vbias.n322 Vbias 0.252372
R21470 Vbias.n324 Vbias 0.252372
R21471 Vbias.n326 Vbias 0.252372
R21472 Vbias.n328 Vbias 0.252372
R21473 Vbias.n330 Vbias 0.252372
R21474 Vbias.n332 Vbias 0.252372
R21475 Vbias.n334 Vbias 0.252372
R21476 Vbias.n336 Vbias 0.252372
R21477 Vbias.n338 Vbias 0.252372
R21478 Vbias.n340 Vbias 0.252372
R21479 Vbias.n342 Vbias 0.252372
R21480 Vbias.n344 Vbias 0.252372
R21481 Vbias.n346 Vbias 0.252372
R21482 Vbias.n348 Vbias 0.252372
R21483 Vbias.n350 Vbias 0.252372
R21484 Vbias.n290 Vbias 0.252372
R21485 Vbias.n292 Vbias 0.252372
R21486 Vbias.n294 Vbias 0.252372
R21487 Vbias.n296 Vbias 0.252372
R21488 Vbias.n298 Vbias 0.252372
R21489 Vbias.n300 Vbias 0.252372
R21490 Vbias.n302 Vbias 0.252372
R21491 Vbias.n304 Vbias 0.252372
R21492 Vbias.n306 Vbias 0.252372
R21493 Vbias.n308 Vbias 0.252372
R21494 Vbias.n310 Vbias 0.252372
R21495 Vbias.n312 Vbias 0.252372
R21496 Vbias.n314 Vbias 0.252372
R21497 Vbias.n316 Vbias 0.252372
R21498 Vbias.n318 Vbias 0.252372
R21499 Vbias.n258 Vbias 0.252372
R21500 Vbias.n260 Vbias 0.252372
R21501 Vbias.n262 Vbias 0.252372
R21502 Vbias.n264 Vbias 0.252372
R21503 Vbias.n266 Vbias 0.252372
R21504 Vbias.n268 Vbias 0.252372
R21505 Vbias.n270 Vbias 0.252372
R21506 Vbias.n272 Vbias 0.252372
R21507 Vbias.n274 Vbias 0.252372
R21508 Vbias.n276 Vbias 0.252372
R21509 Vbias.n278 Vbias 0.252372
R21510 Vbias.n280 Vbias 0.252372
R21511 Vbias.n282 Vbias 0.252372
R21512 Vbias.n284 Vbias 0.252372
R21513 Vbias.n286 Vbias 0.252372
R21514 Vbias.n226 Vbias 0.252372
R21515 Vbias.n228 Vbias 0.252372
R21516 Vbias.n230 Vbias 0.252372
R21517 Vbias.n232 Vbias 0.252372
R21518 Vbias.n234 Vbias 0.252372
R21519 Vbias.n236 Vbias 0.252372
R21520 Vbias.n238 Vbias 0.252372
R21521 Vbias.n240 Vbias 0.252372
R21522 Vbias.n242 Vbias 0.252372
R21523 Vbias.n244 Vbias 0.252372
R21524 Vbias.n246 Vbias 0.252372
R21525 Vbias.n248 Vbias 0.252372
R21526 Vbias.n250 Vbias 0.252372
R21527 Vbias.n252 Vbias 0.252372
R21528 Vbias.n254 Vbias 0.252372
R21529 Vbias.n194 Vbias 0.252372
R21530 Vbias.n196 Vbias 0.252372
R21531 Vbias.n198 Vbias 0.252372
R21532 Vbias.n200 Vbias 0.252372
R21533 Vbias.n202 Vbias 0.252372
R21534 Vbias.n204 Vbias 0.252372
R21535 Vbias.n206 Vbias 0.252372
R21536 Vbias.n208 Vbias 0.252372
R21537 Vbias.n210 Vbias 0.252372
R21538 Vbias.n212 Vbias 0.252372
R21539 Vbias.n214 Vbias 0.252372
R21540 Vbias.n216 Vbias 0.252372
R21541 Vbias.n218 Vbias 0.252372
R21542 Vbias.n220 Vbias 0.252372
R21543 Vbias.n222 Vbias 0.252372
R21544 Vbias.n162 Vbias 0.252372
R21545 Vbias.n164 Vbias 0.252372
R21546 Vbias.n166 Vbias 0.252372
R21547 Vbias.n168 Vbias 0.252372
R21548 Vbias.n170 Vbias 0.252372
R21549 Vbias.n172 Vbias 0.252372
R21550 Vbias.n174 Vbias 0.252372
R21551 Vbias.n176 Vbias 0.252372
R21552 Vbias.n178 Vbias 0.252372
R21553 Vbias.n180 Vbias 0.252372
R21554 Vbias.n182 Vbias 0.252372
R21555 Vbias.n184 Vbias 0.252372
R21556 Vbias.n186 Vbias 0.252372
R21557 Vbias.n188 Vbias 0.252372
R21558 Vbias.n190 Vbias 0.252372
R21559 Vbias.n130 Vbias 0.252372
R21560 Vbias.n132 Vbias 0.252372
R21561 Vbias.n134 Vbias 0.252372
R21562 Vbias.n136 Vbias 0.252372
R21563 Vbias.n138 Vbias 0.252372
R21564 Vbias.n140 Vbias 0.252372
R21565 Vbias.n142 Vbias 0.252372
R21566 Vbias.n144 Vbias 0.252372
R21567 Vbias.n146 Vbias 0.252372
R21568 Vbias.n148 Vbias 0.252372
R21569 Vbias.n150 Vbias 0.252372
R21570 Vbias.n152 Vbias 0.252372
R21571 Vbias.n154 Vbias 0.252372
R21572 Vbias.n156 Vbias 0.252372
R21573 Vbias.n158 Vbias 0.252372
R21574 Vbias.n98 Vbias 0.252372
R21575 Vbias.n100 Vbias 0.252372
R21576 Vbias.n102 Vbias 0.252372
R21577 Vbias.n104 Vbias 0.252372
R21578 Vbias.n106 Vbias 0.252372
R21579 Vbias.n108 Vbias 0.252372
R21580 Vbias.n110 Vbias 0.252372
R21581 Vbias.n112 Vbias 0.252372
R21582 Vbias.n114 Vbias 0.252372
R21583 Vbias.n116 Vbias 0.252372
R21584 Vbias.n118 Vbias 0.252372
R21585 Vbias.n120 Vbias 0.252372
R21586 Vbias.n122 Vbias 0.252372
R21587 Vbias.n124 Vbias 0.252372
R21588 Vbias.n126 Vbias 0.252372
R21589 Vbias.n66 Vbias 0.252372
R21590 Vbias.n68 Vbias 0.252372
R21591 Vbias.n70 Vbias 0.252372
R21592 Vbias.n72 Vbias 0.252372
R21593 Vbias.n74 Vbias 0.252372
R21594 Vbias.n76 Vbias 0.252372
R21595 Vbias.n78 Vbias 0.252372
R21596 Vbias.n80 Vbias 0.252372
R21597 Vbias.n82 Vbias 0.252372
R21598 Vbias.n84 Vbias 0.252372
R21599 Vbias.n86 Vbias 0.252372
R21600 Vbias.n88 Vbias 0.252372
R21601 Vbias.n90 Vbias 0.252372
R21602 Vbias.n92 Vbias 0.252372
R21603 Vbias.n94 Vbias 0.252372
R21604 Vbias.n34 Vbias 0.252372
R21605 Vbias.n36 Vbias 0.252372
R21606 Vbias.n38 Vbias 0.252372
R21607 Vbias.n40 Vbias 0.252372
R21608 Vbias.n42 Vbias 0.252372
R21609 Vbias.n44 Vbias 0.252372
R21610 Vbias.n46 Vbias 0.252372
R21611 Vbias.n48 Vbias 0.252372
R21612 Vbias.n50 Vbias 0.252372
R21613 Vbias.n52 Vbias 0.252372
R21614 Vbias.n54 Vbias 0.252372
R21615 Vbias.n56 Vbias 0.252372
R21616 Vbias.n58 Vbias 0.252372
R21617 Vbias.n60 Vbias 0.252372
R21618 Vbias.n62 Vbias 0.252372
R21619 Vbias.n2 Vbias 0.252372
R21620 Vbias.n4 Vbias 0.252372
R21621 Vbias.n6 Vbias 0.252372
R21622 Vbias.n8 Vbias 0.252372
R21623 Vbias.n10 Vbias 0.252372
R21624 Vbias.n12 Vbias 0.252372
R21625 Vbias.n14 Vbias 0.252372
R21626 Vbias.n16 Vbias 0.252372
R21627 Vbias.n18 Vbias 0.252372
R21628 Vbias.n20 Vbias 0.252372
R21629 Vbias.n22 Vbias 0.252372
R21630 Vbias.n24 Vbias 0.252372
R21631 Vbias.n26 Vbias 0.252372
R21632 Vbias.n28 Vbias 0.252372
R21633 Vbias.n30 Vbias 0.252372
R21634 Vbias Vbias.n524 0.237067
R21635 Vbias.n517 Vbias.n512 0.215542
R21636 Vbias.n523 Vbias.n518 0.215542
R21637 Vbias Vbias.n517 0.175939
R21638 Vbias.n517 Vbias.n516 0.150018
R21639 Vbias.n523 Vbias.n522 0.150018
R21640 Vbias Vbias.n523 0.127693
R21641 Vbias Vbias.n482 0.0972718
R21642 Vbias Vbias.n484 0.0972718
R21643 Vbias Vbias.n486 0.0972718
R21644 Vbias Vbias.n488 0.0972718
R21645 Vbias Vbias.n490 0.0972718
R21646 Vbias Vbias.n492 0.0972718
R21647 Vbias Vbias.n494 0.0972718
R21648 Vbias Vbias.n496 0.0972718
R21649 Vbias Vbias.n498 0.0972718
R21650 Vbias Vbias.n500 0.0972718
R21651 Vbias Vbias.n502 0.0972718
R21652 Vbias Vbias.n504 0.0972718
R21653 Vbias Vbias.n506 0.0972718
R21654 Vbias Vbias.n508 0.0972718
R21655 Vbias Vbias.n510 0.0972718
R21656 Vbias Vbias.n450 0.0972718
R21657 Vbias Vbias.n452 0.0972718
R21658 Vbias Vbias.n454 0.0972718
R21659 Vbias Vbias.n456 0.0972718
R21660 Vbias Vbias.n458 0.0972718
R21661 Vbias Vbias.n460 0.0972718
R21662 Vbias Vbias.n462 0.0972718
R21663 Vbias Vbias.n464 0.0972718
R21664 Vbias Vbias.n466 0.0972718
R21665 Vbias Vbias.n468 0.0972718
R21666 Vbias Vbias.n470 0.0972718
R21667 Vbias Vbias.n472 0.0972718
R21668 Vbias Vbias.n474 0.0972718
R21669 Vbias Vbias.n476 0.0972718
R21670 Vbias Vbias.n478 0.0972718
R21671 Vbias Vbias.n418 0.0972718
R21672 Vbias Vbias.n420 0.0972718
R21673 Vbias Vbias.n422 0.0972718
R21674 Vbias Vbias.n424 0.0972718
R21675 Vbias Vbias.n426 0.0972718
R21676 Vbias Vbias.n428 0.0972718
R21677 Vbias Vbias.n430 0.0972718
R21678 Vbias Vbias.n432 0.0972718
R21679 Vbias Vbias.n434 0.0972718
R21680 Vbias Vbias.n436 0.0972718
R21681 Vbias Vbias.n438 0.0972718
R21682 Vbias Vbias.n440 0.0972718
R21683 Vbias Vbias.n442 0.0972718
R21684 Vbias Vbias.n444 0.0972718
R21685 Vbias Vbias.n446 0.0972718
R21686 Vbias Vbias.n386 0.0972718
R21687 Vbias Vbias.n388 0.0972718
R21688 Vbias Vbias.n390 0.0972718
R21689 Vbias Vbias.n392 0.0972718
R21690 Vbias Vbias.n394 0.0972718
R21691 Vbias Vbias.n396 0.0972718
R21692 Vbias Vbias.n398 0.0972718
R21693 Vbias Vbias.n400 0.0972718
R21694 Vbias Vbias.n402 0.0972718
R21695 Vbias Vbias.n404 0.0972718
R21696 Vbias Vbias.n406 0.0972718
R21697 Vbias Vbias.n408 0.0972718
R21698 Vbias Vbias.n410 0.0972718
R21699 Vbias Vbias.n412 0.0972718
R21700 Vbias Vbias.n414 0.0972718
R21701 Vbias Vbias.n354 0.0972718
R21702 Vbias Vbias.n356 0.0972718
R21703 Vbias Vbias.n358 0.0972718
R21704 Vbias Vbias.n360 0.0972718
R21705 Vbias Vbias.n362 0.0972718
R21706 Vbias Vbias.n364 0.0972718
R21707 Vbias Vbias.n366 0.0972718
R21708 Vbias Vbias.n368 0.0972718
R21709 Vbias Vbias.n370 0.0972718
R21710 Vbias Vbias.n372 0.0972718
R21711 Vbias Vbias.n374 0.0972718
R21712 Vbias Vbias.n376 0.0972718
R21713 Vbias Vbias.n378 0.0972718
R21714 Vbias Vbias.n380 0.0972718
R21715 Vbias Vbias.n382 0.0972718
R21716 Vbias Vbias.n322 0.0972718
R21717 Vbias Vbias.n324 0.0972718
R21718 Vbias Vbias.n326 0.0972718
R21719 Vbias Vbias.n328 0.0972718
R21720 Vbias Vbias.n330 0.0972718
R21721 Vbias Vbias.n332 0.0972718
R21722 Vbias Vbias.n334 0.0972718
R21723 Vbias Vbias.n336 0.0972718
R21724 Vbias Vbias.n338 0.0972718
R21725 Vbias Vbias.n340 0.0972718
R21726 Vbias Vbias.n342 0.0972718
R21727 Vbias Vbias.n344 0.0972718
R21728 Vbias Vbias.n346 0.0972718
R21729 Vbias Vbias.n348 0.0972718
R21730 Vbias Vbias.n350 0.0972718
R21731 Vbias Vbias.n290 0.0972718
R21732 Vbias Vbias.n292 0.0972718
R21733 Vbias Vbias.n294 0.0972718
R21734 Vbias Vbias.n296 0.0972718
R21735 Vbias Vbias.n298 0.0972718
R21736 Vbias Vbias.n300 0.0972718
R21737 Vbias Vbias.n302 0.0972718
R21738 Vbias Vbias.n304 0.0972718
R21739 Vbias Vbias.n306 0.0972718
R21740 Vbias Vbias.n308 0.0972718
R21741 Vbias Vbias.n310 0.0972718
R21742 Vbias Vbias.n312 0.0972718
R21743 Vbias Vbias.n314 0.0972718
R21744 Vbias Vbias.n316 0.0972718
R21745 Vbias Vbias.n318 0.0972718
R21746 Vbias Vbias.n258 0.0972718
R21747 Vbias Vbias.n260 0.0972718
R21748 Vbias Vbias.n262 0.0972718
R21749 Vbias Vbias.n264 0.0972718
R21750 Vbias Vbias.n266 0.0972718
R21751 Vbias Vbias.n268 0.0972718
R21752 Vbias Vbias.n270 0.0972718
R21753 Vbias Vbias.n272 0.0972718
R21754 Vbias Vbias.n274 0.0972718
R21755 Vbias Vbias.n276 0.0972718
R21756 Vbias Vbias.n278 0.0972718
R21757 Vbias Vbias.n280 0.0972718
R21758 Vbias Vbias.n282 0.0972718
R21759 Vbias Vbias.n284 0.0972718
R21760 Vbias Vbias.n286 0.0972718
R21761 Vbias Vbias.n226 0.0972718
R21762 Vbias Vbias.n228 0.0972718
R21763 Vbias Vbias.n230 0.0972718
R21764 Vbias Vbias.n232 0.0972718
R21765 Vbias Vbias.n234 0.0972718
R21766 Vbias Vbias.n236 0.0972718
R21767 Vbias Vbias.n238 0.0972718
R21768 Vbias Vbias.n240 0.0972718
R21769 Vbias Vbias.n242 0.0972718
R21770 Vbias Vbias.n244 0.0972718
R21771 Vbias Vbias.n246 0.0972718
R21772 Vbias Vbias.n248 0.0972718
R21773 Vbias Vbias.n250 0.0972718
R21774 Vbias Vbias.n252 0.0972718
R21775 Vbias Vbias.n254 0.0972718
R21776 Vbias Vbias.n194 0.0972718
R21777 Vbias Vbias.n196 0.0972718
R21778 Vbias Vbias.n198 0.0972718
R21779 Vbias Vbias.n200 0.0972718
R21780 Vbias Vbias.n202 0.0972718
R21781 Vbias Vbias.n204 0.0972718
R21782 Vbias Vbias.n206 0.0972718
R21783 Vbias Vbias.n208 0.0972718
R21784 Vbias Vbias.n210 0.0972718
R21785 Vbias Vbias.n212 0.0972718
R21786 Vbias Vbias.n214 0.0972718
R21787 Vbias Vbias.n216 0.0972718
R21788 Vbias Vbias.n218 0.0972718
R21789 Vbias Vbias.n220 0.0972718
R21790 Vbias Vbias.n222 0.0972718
R21791 Vbias Vbias.n162 0.0972718
R21792 Vbias Vbias.n164 0.0972718
R21793 Vbias Vbias.n166 0.0972718
R21794 Vbias Vbias.n168 0.0972718
R21795 Vbias Vbias.n170 0.0972718
R21796 Vbias Vbias.n172 0.0972718
R21797 Vbias Vbias.n174 0.0972718
R21798 Vbias Vbias.n176 0.0972718
R21799 Vbias Vbias.n178 0.0972718
R21800 Vbias Vbias.n180 0.0972718
R21801 Vbias Vbias.n182 0.0972718
R21802 Vbias Vbias.n184 0.0972718
R21803 Vbias Vbias.n186 0.0972718
R21804 Vbias Vbias.n188 0.0972718
R21805 Vbias Vbias.n190 0.0972718
R21806 Vbias Vbias.n130 0.0972718
R21807 Vbias Vbias.n132 0.0972718
R21808 Vbias Vbias.n134 0.0972718
R21809 Vbias Vbias.n136 0.0972718
R21810 Vbias Vbias.n138 0.0972718
R21811 Vbias Vbias.n140 0.0972718
R21812 Vbias Vbias.n142 0.0972718
R21813 Vbias Vbias.n144 0.0972718
R21814 Vbias Vbias.n146 0.0972718
R21815 Vbias Vbias.n148 0.0972718
R21816 Vbias Vbias.n150 0.0972718
R21817 Vbias Vbias.n152 0.0972718
R21818 Vbias Vbias.n154 0.0972718
R21819 Vbias Vbias.n156 0.0972718
R21820 Vbias Vbias.n158 0.0972718
R21821 Vbias Vbias.n98 0.0972718
R21822 Vbias Vbias.n100 0.0972718
R21823 Vbias Vbias.n102 0.0972718
R21824 Vbias Vbias.n104 0.0972718
R21825 Vbias Vbias.n106 0.0972718
R21826 Vbias Vbias.n108 0.0972718
R21827 Vbias Vbias.n110 0.0972718
R21828 Vbias Vbias.n112 0.0972718
R21829 Vbias Vbias.n114 0.0972718
R21830 Vbias Vbias.n116 0.0972718
R21831 Vbias Vbias.n118 0.0972718
R21832 Vbias Vbias.n120 0.0972718
R21833 Vbias Vbias.n122 0.0972718
R21834 Vbias Vbias.n124 0.0972718
R21835 Vbias Vbias.n126 0.0972718
R21836 Vbias Vbias.n66 0.0972718
R21837 Vbias Vbias.n68 0.0972718
R21838 Vbias Vbias.n70 0.0972718
R21839 Vbias Vbias.n72 0.0972718
R21840 Vbias Vbias.n74 0.0972718
R21841 Vbias Vbias.n76 0.0972718
R21842 Vbias Vbias.n78 0.0972718
R21843 Vbias Vbias.n80 0.0972718
R21844 Vbias Vbias.n82 0.0972718
R21845 Vbias Vbias.n84 0.0972718
R21846 Vbias Vbias.n86 0.0972718
R21847 Vbias Vbias.n88 0.0972718
R21848 Vbias Vbias.n90 0.0972718
R21849 Vbias Vbias.n92 0.0972718
R21850 Vbias Vbias.n94 0.0972718
R21851 Vbias Vbias.n34 0.0972718
R21852 Vbias Vbias.n36 0.0972718
R21853 Vbias Vbias.n38 0.0972718
R21854 Vbias Vbias.n40 0.0972718
R21855 Vbias Vbias.n42 0.0972718
R21856 Vbias Vbias.n44 0.0972718
R21857 Vbias Vbias.n46 0.0972718
R21858 Vbias Vbias.n48 0.0972718
R21859 Vbias Vbias.n50 0.0972718
R21860 Vbias Vbias.n52 0.0972718
R21861 Vbias Vbias.n54 0.0972718
R21862 Vbias Vbias.n56 0.0972718
R21863 Vbias Vbias.n58 0.0972718
R21864 Vbias Vbias.n60 0.0972718
R21865 Vbias Vbias.n62 0.0972718
R21866 Vbias Vbias.n2 0.0972718
R21867 Vbias Vbias.n4 0.0972718
R21868 Vbias Vbias.n6 0.0972718
R21869 Vbias Vbias.n8 0.0972718
R21870 Vbias Vbias.n10 0.0972718
R21871 Vbias Vbias.n12 0.0972718
R21872 Vbias Vbias.n14 0.0972718
R21873 Vbias Vbias.n16 0.0972718
R21874 Vbias Vbias.n18 0.0972718
R21875 Vbias Vbias.n20 0.0972718
R21876 Vbias Vbias.n22 0.0972718
R21877 Vbias Vbias.n24 0.0972718
R21878 Vbias Vbias.n26 0.0972718
R21879 Vbias Vbias.n28 0.0972718
R21880 Vbias Vbias.n30 0.0972718
R21881 Vbias.n509 Vbias 0.0489375
R21882 Vbias.n507 Vbias 0.0489375
R21883 Vbias.n505 Vbias 0.0489375
R21884 Vbias.n503 Vbias 0.0489375
R21885 Vbias.n501 Vbias 0.0489375
R21886 Vbias.n499 Vbias 0.0489375
R21887 Vbias.n497 Vbias 0.0489375
R21888 Vbias.n495 Vbias 0.0489375
R21889 Vbias.n493 Vbias 0.0489375
R21890 Vbias.n491 Vbias 0.0489375
R21891 Vbias.n489 Vbias 0.0489375
R21892 Vbias.n487 Vbias 0.0489375
R21893 Vbias.n485 Vbias 0.0489375
R21894 Vbias.n483 Vbias 0.0489375
R21895 Vbias.n481 Vbias 0.0489375
R21896 Vbias.n480 Vbias 0.0489375
R21897 Vbias.n477 Vbias 0.0489375
R21898 Vbias.n475 Vbias 0.0489375
R21899 Vbias.n473 Vbias 0.0489375
R21900 Vbias.n471 Vbias 0.0489375
R21901 Vbias.n469 Vbias 0.0489375
R21902 Vbias.n467 Vbias 0.0489375
R21903 Vbias.n465 Vbias 0.0489375
R21904 Vbias.n463 Vbias 0.0489375
R21905 Vbias.n461 Vbias 0.0489375
R21906 Vbias.n459 Vbias 0.0489375
R21907 Vbias.n457 Vbias 0.0489375
R21908 Vbias.n455 Vbias 0.0489375
R21909 Vbias.n453 Vbias 0.0489375
R21910 Vbias.n451 Vbias 0.0489375
R21911 Vbias.n449 Vbias 0.0489375
R21912 Vbias.n448 Vbias 0.0489375
R21913 Vbias.n445 Vbias 0.0489375
R21914 Vbias.n443 Vbias 0.0489375
R21915 Vbias.n441 Vbias 0.0489375
R21916 Vbias.n439 Vbias 0.0489375
R21917 Vbias.n437 Vbias 0.0489375
R21918 Vbias.n435 Vbias 0.0489375
R21919 Vbias.n433 Vbias 0.0489375
R21920 Vbias.n431 Vbias 0.0489375
R21921 Vbias.n429 Vbias 0.0489375
R21922 Vbias.n427 Vbias 0.0489375
R21923 Vbias.n425 Vbias 0.0489375
R21924 Vbias.n423 Vbias 0.0489375
R21925 Vbias.n421 Vbias 0.0489375
R21926 Vbias.n419 Vbias 0.0489375
R21927 Vbias.n417 Vbias 0.0489375
R21928 Vbias.n416 Vbias 0.0489375
R21929 Vbias.n413 Vbias 0.0489375
R21930 Vbias.n411 Vbias 0.0489375
R21931 Vbias.n409 Vbias 0.0489375
R21932 Vbias.n407 Vbias 0.0489375
R21933 Vbias.n405 Vbias 0.0489375
R21934 Vbias.n403 Vbias 0.0489375
R21935 Vbias.n401 Vbias 0.0489375
R21936 Vbias.n399 Vbias 0.0489375
R21937 Vbias.n397 Vbias 0.0489375
R21938 Vbias.n395 Vbias 0.0489375
R21939 Vbias.n393 Vbias 0.0489375
R21940 Vbias.n391 Vbias 0.0489375
R21941 Vbias.n389 Vbias 0.0489375
R21942 Vbias.n387 Vbias 0.0489375
R21943 Vbias.n385 Vbias 0.0489375
R21944 Vbias.n384 Vbias 0.0489375
R21945 Vbias.n381 Vbias 0.0489375
R21946 Vbias.n379 Vbias 0.0489375
R21947 Vbias.n377 Vbias 0.0489375
R21948 Vbias.n375 Vbias 0.0489375
R21949 Vbias.n373 Vbias 0.0489375
R21950 Vbias.n371 Vbias 0.0489375
R21951 Vbias.n369 Vbias 0.0489375
R21952 Vbias.n367 Vbias 0.0489375
R21953 Vbias.n365 Vbias 0.0489375
R21954 Vbias.n363 Vbias 0.0489375
R21955 Vbias.n361 Vbias 0.0489375
R21956 Vbias.n359 Vbias 0.0489375
R21957 Vbias.n357 Vbias 0.0489375
R21958 Vbias.n355 Vbias 0.0489375
R21959 Vbias.n353 Vbias 0.0489375
R21960 Vbias.n352 Vbias 0.0489375
R21961 Vbias.n349 Vbias 0.0489375
R21962 Vbias.n347 Vbias 0.0489375
R21963 Vbias.n345 Vbias 0.0489375
R21964 Vbias.n343 Vbias 0.0489375
R21965 Vbias.n341 Vbias 0.0489375
R21966 Vbias.n339 Vbias 0.0489375
R21967 Vbias.n337 Vbias 0.0489375
R21968 Vbias.n335 Vbias 0.0489375
R21969 Vbias.n333 Vbias 0.0489375
R21970 Vbias.n331 Vbias 0.0489375
R21971 Vbias.n329 Vbias 0.0489375
R21972 Vbias.n327 Vbias 0.0489375
R21973 Vbias.n325 Vbias 0.0489375
R21974 Vbias.n323 Vbias 0.0489375
R21975 Vbias.n321 Vbias 0.0489375
R21976 Vbias.n320 Vbias 0.0489375
R21977 Vbias.n317 Vbias 0.0489375
R21978 Vbias.n315 Vbias 0.0489375
R21979 Vbias.n313 Vbias 0.0489375
R21980 Vbias.n311 Vbias 0.0489375
R21981 Vbias.n309 Vbias 0.0489375
R21982 Vbias.n307 Vbias 0.0489375
R21983 Vbias.n305 Vbias 0.0489375
R21984 Vbias.n303 Vbias 0.0489375
R21985 Vbias.n301 Vbias 0.0489375
R21986 Vbias.n299 Vbias 0.0489375
R21987 Vbias.n297 Vbias 0.0489375
R21988 Vbias.n295 Vbias 0.0489375
R21989 Vbias.n293 Vbias 0.0489375
R21990 Vbias.n291 Vbias 0.0489375
R21991 Vbias.n289 Vbias 0.0489375
R21992 Vbias.n288 Vbias 0.0489375
R21993 Vbias.n285 Vbias 0.0489375
R21994 Vbias.n283 Vbias 0.0489375
R21995 Vbias.n281 Vbias 0.0489375
R21996 Vbias.n279 Vbias 0.0489375
R21997 Vbias.n277 Vbias 0.0489375
R21998 Vbias.n275 Vbias 0.0489375
R21999 Vbias.n273 Vbias 0.0489375
R22000 Vbias.n271 Vbias 0.0489375
R22001 Vbias.n269 Vbias 0.0489375
R22002 Vbias.n267 Vbias 0.0489375
R22003 Vbias.n265 Vbias 0.0489375
R22004 Vbias.n263 Vbias 0.0489375
R22005 Vbias.n261 Vbias 0.0489375
R22006 Vbias.n259 Vbias 0.0489375
R22007 Vbias.n257 Vbias 0.0489375
R22008 Vbias.n256 Vbias 0.0489375
R22009 Vbias.n253 Vbias 0.0489375
R22010 Vbias.n251 Vbias 0.0489375
R22011 Vbias.n249 Vbias 0.0489375
R22012 Vbias.n247 Vbias 0.0489375
R22013 Vbias.n245 Vbias 0.0489375
R22014 Vbias.n243 Vbias 0.0489375
R22015 Vbias.n241 Vbias 0.0489375
R22016 Vbias.n239 Vbias 0.0489375
R22017 Vbias.n237 Vbias 0.0489375
R22018 Vbias.n235 Vbias 0.0489375
R22019 Vbias.n233 Vbias 0.0489375
R22020 Vbias.n231 Vbias 0.0489375
R22021 Vbias.n229 Vbias 0.0489375
R22022 Vbias.n227 Vbias 0.0489375
R22023 Vbias.n225 Vbias 0.0489375
R22024 Vbias.n224 Vbias 0.0489375
R22025 Vbias.n221 Vbias 0.0489375
R22026 Vbias.n219 Vbias 0.0489375
R22027 Vbias.n217 Vbias 0.0489375
R22028 Vbias.n215 Vbias 0.0489375
R22029 Vbias.n213 Vbias 0.0489375
R22030 Vbias.n211 Vbias 0.0489375
R22031 Vbias.n209 Vbias 0.0489375
R22032 Vbias.n207 Vbias 0.0489375
R22033 Vbias.n205 Vbias 0.0489375
R22034 Vbias.n203 Vbias 0.0489375
R22035 Vbias.n201 Vbias 0.0489375
R22036 Vbias.n199 Vbias 0.0489375
R22037 Vbias.n197 Vbias 0.0489375
R22038 Vbias.n195 Vbias 0.0489375
R22039 Vbias.n193 Vbias 0.0489375
R22040 Vbias.n192 Vbias 0.0489375
R22041 Vbias.n189 Vbias 0.0489375
R22042 Vbias.n187 Vbias 0.0489375
R22043 Vbias.n185 Vbias 0.0489375
R22044 Vbias.n183 Vbias 0.0489375
R22045 Vbias.n181 Vbias 0.0489375
R22046 Vbias.n179 Vbias 0.0489375
R22047 Vbias.n177 Vbias 0.0489375
R22048 Vbias.n175 Vbias 0.0489375
R22049 Vbias.n173 Vbias 0.0489375
R22050 Vbias.n171 Vbias 0.0489375
R22051 Vbias.n169 Vbias 0.0489375
R22052 Vbias.n167 Vbias 0.0489375
R22053 Vbias.n165 Vbias 0.0489375
R22054 Vbias.n163 Vbias 0.0489375
R22055 Vbias.n161 Vbias 0.0489375
R22056 Vbias.n160 Vbias 0.0489375
R22057 Vbias.n157 Vbias 0.0489375
R22058 Vbias.n155 Vbias 0.0489375
R22059 Vbias.n153 Vbias 0.0489375
R22060 Vbias.n151 Vbias 0.0489375
R22061 Vbias.n149 Vbias 0.0489375
R22062 Vbias.n147 Vbias 0.0489375
R22063 Vbias.n145 Vbias 0.0489375
R22064 Vbias.n143 Vbias 0.0489375
R22065 Vbias.n141 Vbias 0.0489375
R22066 Vbias.n139 Vbias 0.0489375
R22067 Vbias.n137 Vbias 0.0489375
R22068 Vbias.n135 Vbias 0.0489375
R22069 Vbias.n133 Vbias 0.0489375
R22070 Vbias.n131 Vbias 0.0489375
R22071 Vbias.n129 Vbias 0.0489375
R22072 Vbias.n128 Vbias 0.0489375
R22073 Vbias.n125 Vbias 0.0489375
R22074 Vbias.n123 Vbias 0.0489375
R22075 Vbias.n121 Vbias 0.0489375
R22076 Vbias.n119 Vbias 0.0489375
R22077 Vbias.n117 Vbias 0.0489375
R22078 Vbias.n115 Vbias 0.0489375
R22079 Vbias.n113 Vbias 0.0489375
R22080 Vbias.n111 Vbias 0.0489375
R22081 Vbias.n109 Vbias 0.0489375
R22082 Vbias.n107 Vbias 0.0489375
R22083 Vbias.n105 Vbias 0.0489375
R22084 Vbias.n103 Vbias 0.0489375
R22085 Vbias.n101 Vbias 0.0489375
R22086 Vbias.n99 Vbias 0.0489375
R22087 Vbias.n97 Vbias 0.0489375
R22088 Vbias.n96 Vbias 0.0489375
R22089 Vbias.n93 Vbias 0.0489375
R22090 Vbias.n91 Vbias 0.0489375
R22091 Vbias.n89 Vbias 0.0489375
R22092 Vbias.n87 Vbias 0.0489375
R22093 Vbias.n85 Vbias 0.0489375
R22094 Vbias.n83 Vbias 0.0489375
R22095 Vbias.n81 Vbias 0.0489375
R22096 Vbias.n79 Vbias 0.0489375
R22097 Vbias.n77 Vbias 0.0489375
R22098 Vbias.n75 Vbias 0.0489375
R22099 Vbias.n73 Vbias 0.0489375
R22100 Vbias.n71 Vbias 0.0489375
R22101 Vbias.n69 Vbias 0.0489375
R22102 Vbias.n67 Vbias 0.0489375
R22103 Vbias.n65 Vbias 0.0489375
R22104 Vbias.n64 Vbias 0.0489375
R22105 Vbias.n61 Vbias 0.0489375
R22106 Vbias.n59 Vbias 0.0489375
R22107 Vbias.n57 Vbias 0.0489375
R22108 Vbias.n55 Vbias 0.0489375
R22109 Vbias.n53 Vbias 0.0489375
R22110 Vbias.n51 Vbias 0.0489375
R22111 Vbias.n49 Vbias 0.0489375
R22112 Vbias.n47 Vbias 0.0489375
R22113 Vbias.n45 Vbias 0.0489375
R22114 Vbias.n43 Vbias 0.0489375
R22115 Vbias.n41 Vbias 0.0489375
R22116 Vbias.n39 Vbias 0.0489375
R22117 Vbias.n37 Vbias 0.0489375
R22118 Vbias.n35 Vbias 0.0489375
R22119 Vbias.n33 Vbias 0.0489375
R22120 Vbias.n32 Vbias 0.0489375
R22121 Vbias.n29 Vbias 0.0489375
R22122 Vbias.n27 Vbias 0.0489375
R22123 Vbias.n25 Vbias 0.0489375
R22124 Vbias.n23 Vbias 0.0489375
R22125 Vbias.n21 Vbias 0.0489375
R22126 Vbias.n19 Vbias 0.0489375
R22127 Vbias.n17 Vbias 0.0489375
R22128 Vbias.n15 Vbias 0.0489375
R22129 Vbias.n13 Vbias 0.0489375
R22130 Vbias.n11 Vbias 0.0489375
R22131 Vbias.n9 Vbias 0.0489375
R22132 Vbias.n7 Vbias 0.0489375
R22133 Vbias.n5 Vbias 0.0489375
R22134 Vbias.n3 Vbias 0.0489375
R22135 Vbias.n1 Vbias 0.0489375
R22136 Vbias.n0 Vbias 0.0489375
R22137 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R22138 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R22139 XThC.Tn[1].n12 XThC.Tn[1].n10 161.406
R22140 XThC.Tn[1].n15 XThC.Tn[1].n13 161.406
R22141 XThC.Tn[1].n18 XThC.Tn[1].n16 161.406
R22142 XThC.Tn[1].n21 XThC.Tn[1].n19 161.406
R22143 XThC.Tn[1].n24 XThC.Tn[1].n22 161.406
R22144 XThC.Tn[1].n27 XThC.Tn[1].n25 161.406
R22145 XThC.Tn[1].n30 XThC.Tn[1].n28 161.406
R22146 XThC.Tn[1].n33 XThC.Tn[1].n31 161.406
R22147 XThC.Tn[1].n36 XThC.Tn[1].n34 161.406
R22148 XThC.Tn[1].n39 XThC.Tn[1].n37 161.406
R22149 XThC.Tn[1].n42 XThC.Tn[1].n40 161.406
R22150 XThC.Tn[1].n45 XThC.Tn[1].n43 161.406
R22151 XThC.Tn[1].n48 XThC.Tn[1].n46 161.406
R22152 XThC.Tn[1].n51 XThC.Tn[1].n49 161.406
R22153 XThC.Tn[1].n54 XThC.Tn[1].n52 161.406
R22154 XThC.Tn[1].n57 XThC.Tn[1].n55 161.406
R22155 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R22156 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R22157 XThC.Tn[1].n16 XThC.Tn[1].t16 161.202
R22158 XThC.Tn[1].n19 XThC.Tn[1].t18 161.202
R22159 XThC.Tn[1].n22 XThC.Tn[1].t39 161.202
R22160 XThC.Tn[1].n25 XThC.Tn[1].t40 161.202
R22161 XThC.Tn[1].n28 XThC.Tn[1].t21 161.202
R22162 XThC.Tn[1].n31 XThC.Tn[1].t30 161.202
R22163 XThC.Tn[1].n34 XThC.Tn[1].t32 161.202
R22164 XThC.Tn[1].n37 XThC.Tn[1].t19 161.202
R22165 XThC.Tn[1].n40 XThC.Tn[1].t20 161.202
R22166 XThC.Tn[1].n43 XThC.Tn[1].t33 161.202
R22167 XThC.Tn[1].n46 XThC.Tn[1].t41 161.202
R22168 XThC.Tn[1].n49 XThC.Tn[1].t12 161.202
R22169 XThC.Tn[1].n52 XThC.Tn[1].t25 161.202
R22170 XThC.Tn[1].n55 XThC.Tn[1].t35 161.202
R22171 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R22172 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R22173 XThC.Tn[1].n16 XThC.Tn[1].t22 145.137
R22174 XThC.Tn[1].n19 XThC.Tn[1].t23 145.137
R22175 XThC.Tn[1].n22 XThC.Tn[1].t42 145.137
R22176 XThC.Tn[1].n25 XThC.Tn[1].t43 145.137
R22177 XThC.Tn[1].n28 XThC.Tn[1].t27 145.137
R22178 XThC.Tn[1].n31 XThC.Tn[1].t34 145.137
R22179 XThC.Tn[1].n34 XThC.Tn[1].t36 145.137
R22180 XThC.Tn[1].n37 XThC.Tn[1].t24 145.137
R22181 XThC.Tn[1].n40 XThC.Tn[1].t26 145.137
R22182 XThC.Tn[1].n43 XThC.Tn[1].t37 145.137
R22183 XThC.Tn[1].n46 XThC.Tn[1].t13 145.137
R22184 XThC.Tn[1].n49 XThC.Tn[1].t15 145.137
R22185 XThC.Tn[1].n52 XThC.Tn[1].t28 145.137
R22186 XThC.Tn[1].n55 XThC.Tn[1].t38 145.137
R22187 XThC.Tn[1].n7 XThC.Tn[1].n6 135.249
R22188 XThC.Tn[1].n9 XThC.Tn[1].n3 98.981
R22189 XThC.Tn[1].n8 XThC.Tn[1].n4 98.981
R22190 XThC.Tn[1].n7 XThC.Tn[1].n5 98.981
R22191 XThC.Tn[1].n9 XThC.Tn[1].n8 36.2672
R22192 XThC.Tn[1].n8 XThC.Tn[1].n7 36.2672
R22193 XThC.Tn[1].n59 XThC.Tn[1].n9 32.6405
R22194 XThC.Tn[1].n1 XThC.Tn[1].t9 26.5955
R22195 XThC.Tn[1].n1 XThC.Tn[1].t8 26.5955
R22196 XThC.Tn[1].n0 XThC.Tn[1].t11 26.5955
R22197 XThC.Tn[1].n0 XThC.Tn[1].t10 26.5955
R22198 XThC.Tn[1].n3 XThC.Tn[1].t5 24.9236
R22199 XThC.Tn[1].n3 XThC.Tn[1].t4 24.9236
R22200 XThC.Tn[1].n4 XThC.Tn[1].t7 24.9236
R22201 XThC.Tn[1].n4 XThC.Tn[1].t6 24.9236
R22202 XThC.Tn[1].n5 XThC.Tn[1].t1 24.9236
R22203 XThC.Tn[1].n5 XThC.Tn[1].t0 24.9236
R22204 XThC.Tn[1].n6 XThC.Tn[1].t3 24.9236
R22205 XThC.Tn[1].n6 XThC.Tn[1].t2 24.9236
R22206 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R22207 XThC.Tn[1].n58 XThC.Tn[1] 7.29217
R22208 XThC.Tn[1] XThC.Tn[1].n59 6.7205
R22209 XThC.Tn[1].n59 XThC.Tn[1].n58 3.13711
R22210 XThC.Tn[1].n15 XThC.Tn[1] 0.931056
R22211 XThC.Tn[1].n18 XThC.Tn[1] 0.931056
R22212 XThC.Tn[1].n21 XThC.Tn[1] 0.931056
R22213 XThC.Tn[1].n24 XThC.Tn[1] 0.931056
R22214 XThC.Tn[1].n27 XThC.Tn[1] 0.931056
R22215 XThC.Tn[1].n30 XThC.Tn[1] 0.931056
R22216 XThC.Tn[1].n33 XThC.Tn[1] 0.931056
R22217 XThC.Tn[1].n36 XThC.Tn[1] 0.931056
R22218 XThC.Tn[1].n39 XThC.Tn[1] 0.931056
R22219 XThC.Tn[1].n42 XThC.Tn[1] 0.931056
R22220 XThC.Tn[1].n45 XThC.Tn[1] 0.931056
R22221 XThC.Tn[1].n48 XThC.Tn[1] 0.931056
R22222 XThC.Tn[1].n51 XThC.Tn[1] 0.931056
R22223 XThC.Tn[1].n54 XThC.Tn[1] 0.931056
R22224 XThC.Tn[1].n57 XThC.Tn[1] 0.931056
R22225 XThC.Tn[1] XThC.Tn[1].n12 0.396333
R22226 XThC.Tn[1] XThC.Tn[1].n15 0.396333
R22227 XThC.Tn[1] XThC.Tn[1].n18 0.396333
R22228 XThC.Tn[1] XThC.Tn[1].n21 0.396333
R22229 XThC.Tn[1] XThC.Tn[1].n24 0.396333
R22230 XThC.Tn[1] XThC.Tn[1].n27 0.396333
R22231 XThC.Tn[1] XThC.Tn[1].n30 0.396333
R22232 XThC.Tn[1] XThC.Tn[1].n33 0.396333
R22233 XThC.Tn[1] XThC.Tn[1].n36 0.396333
R22234 XThC.Tn[1] XThC.Tn[1].n39 0.396333
R22235 XThC.Tn[1] XThC.Tn[1].n42 0.396333
R22236 XThC.Tn[1] XThC.Tn[1].n45 0.396333
R22237 XThC.Tn[1] XThC.Tn[1].n48 0.396333
R22238 XThC.Tn[1] XThC.Tn[1].n51 0.396333
R22239 XThC.Tn[1] XThC.Tn[1].n54 0.396333
R22240 XThC.Tn[1] XThC.Tn[1].n57 0.396333
R22241 XThC.Tn[1].n11 XThC.Tn[1] 0.104667
R22242 XThC.Tn[1].n14 XThC.Tn[1] 0.104667
R22243 XThC.Tn[1].n17 XThC.Tn[1] 0.104667
R22244 XThC.Tn[1].n20 XThC.Tn[1] 0.104667
R22245 XThC.Tn[1].n23 XThC.Tn[1] 0.104667
R22246 XThC.Tn[1].n26 XThC.Tn[1] 0.104667
R22247 XThC.Tn[1].n29 XThC.Tn[1] 0.104667
R22248 XThC.Tn[1].n32 XThC.Tn[1] 0.104667
R22249 XThC.Tn[1].n35 XThC.Tn[1] 0.104667
R22250 XThC.Tn[1].n38 XThC.Tn[1] 0.104667
R22251 XThC.Tn[1].n41 XThC.Tn[1] 0.104667
R22252 XThC.Tn[1].n44 XThC.Tn[1] 0.104667
R22253 XThC.Tn[1].n47 XThC.Tn[1] 0.104667
R22254 XThC.Tn[1].n50 XThC.Tn[1] 0.104667
R22255 XThC.Tn[1].n53 XThC.Tn[1] 0.104667
R22256 XThC.Tn[1].n56 XThC.Tn[1] 0.104667
R22257 XThC.Tn[1].n58 XThC.Tn[1] 0.0594286
R22258 XThC.Tn[1].n11 XThC.Tn[1] 0.0309878
R22259 XThC.Tn[1].n14 XThC.Tn[1] 0.0309878
R22260 XThC.Tn[1].n17 XThC.Tn[1] 0.0309878
R22261 XThC.Tn[1].n20 XThC.Tn[1] 0.0309878
R22262 XThC.Tn[1].n23 XThC.Tn[1] 0.0309878
R22263 XThC.Tn[1].n26 XThC.Tn[1] 0.0309878
R22264 XThC.Tn[1].n29 XThC.Tn[1] 0.0309878
R22265 XThC.Tn[1].n32 XThC.Tn[1] 0.0309878
R22266 XThC.Tn[1].n35 XThC.Tn[1] 0.0309878
R22267 XThC.Tn[1].n38 XThC.Tn[1] 0.0309878
R22268 XThC.Tn[1].n41 XThC.Tn[1] 0.0309878
R22269 XThC.Tn[1].n44 XThC.Tn[1] 0.0309878
R22270 XThC.Tn[1].n47 XThC.Tn[1] 0.0309878
R22271 XThC.Tn[1].n50 XThC.Tn[1] 0.0309878
R22272 XThC.Tn[1].n53 XThC.Tn[1] 0.0309878
R22273 XThC.Tn[1].n56 XThC.Tn[1] 0.0309878
R22274 XThC.Tn[1].n12 XThC.Tn[1].n11 0.027939
R22275 XThC.Tn[1].n15 XThC.Tn[1].n14 0.027939
R22276 XThC.Tn[1].n18 XThC.Tn[1].n17 0.027939
R22277 XThC.Tn[1].n21 XThC.Tn[1].n20 0.027939
R22278 XThC.Tn[1].n24 XThC.Tn[1].n23 0.027939
R22279 XThC.Tn[1].n27 XThC.Tn[1].n26 0.027939
R22280 XThC.Tn[1].n30 XThC.Tn[1].n29 0.027939
R22281 XThC.Tn[1].n33 XThC.Tn[1].n32 0.027939
R22282 XThC.Tn[1].n36 XThC.Tn[1].n35 0.027939
R22283 XThC.Tn[1].n39 XThC.Tn[1].n38 0.027939
R22284 XThC.Tn[1].n42 XThC.Tn[1].n41 0.027939
R22285 XThC.Tn[1].n45 XThC.Tn[1].n44 0.027939
R22286 XThC.Tn[1].n48 XThC.Tn[1].n47 0.027939
R22287 XThC.Tn[1].n51 XThC.Tn[1].n50 0.027939
R22288 XThC.Tn[1].n54 XThC.Tn[1].n53 0.027939
R22289 XThC.Tn[1].n57 XThC.Tn[1].n56 0.027939
R22290 XThC.Tn[3].n2 XThC.Tn[3].n1 332.332
R22291 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R22292 XThC.Tn[3].n12 XThC.Tn[3].n10 161.406
R22293 XThC.Tn[3].n15 XThC.Tn[3].n13 161.406
R22294 XThC.Tn[3].n18 XThC.Tn[3].n16 161.406
R22295 XThC.Tn[3].n21 XThC.Tn[3].n19 161.406
R22296 XThC.Tn[3].n24 XThC.Tn[3].n22 161.406
R22297 XThC.Tn[3].n27 XThC.Tn[3].n25 161.406
R22298 XThC.Tn[3].n30 XThC.Tn[3].n28 161.406
R22299 XThC.Tn[3].n33 XThC.Tn[3].n31 161.406
R22300 XThC.Tn[3].n36 XThC.Tn[3].n34 161.406
R22301 XThC.Tn[3].n39 XThC.Tn[3].n37 161.406
R22302 XThC.Tn[3].n42 XThC.Tn[3].n40 161.406
R22303 XThC.Tn[3].n45 XThC.Tn[3].n43 161.406
R22304 XThC.Tn[3].n48 XThC.Tn[3].n46 161.406
R22305 XThC.Tn[3].n51 XThC.Tn[3].n49 161.406
R22306 XThC.Tn[3].n54 XThC.Tn[3].n52 161.406
R22307 XThC.Tn[3].n57 XThC.Tn[3].n55 161.406
R22308 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R22309 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R22310 XThC.Tn[3].n16 XThC.Tn[3].t29 161.202
R22311 XThC.Tn[3].n19 XThC.Tn[3].t31 161.202
R22312 XThC.Tn[3].n22 XThC.Tn[3].t20 161.202
R22313 XThC.Tn[3].n25 XThC.Tn[3].t21 161.202
R22314 XThC.Tn[3].n28 XThC.Tn[3].t34 161.202
R22315 XThC.Tn[3].n31 XThC.Tn[3].t43 161.202
R22316 XThC.Tn[3].n34 XThC.Tn[3].t13 161.202
R22317 XThC.Tn[3].n37 XThC.Tn[3].t32 161.202
R22318 XThC.Tn[3].n40 XThC.Tn[3].t33 161.202
R22319 XThC.Tn[3].n43 XThC.Tn[3].t14 161.202
R22320 XThC.Tn[3].n46 XThC.Tn[3].t22 161.202
R22321 XThC.Tn[3].n49 XThC.Tn[3].t25 161.202
R22322 XThC.Tn[3].n52 XThC.Tn[3].t38 161.202
R22323 XThC.Tn[3].n55 XThC.Tn[3].t16 161.202
R22324 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R22325 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R22326 XThC.Tn[3].n16 XThC.Tn[3].t35 145.137
R22327 XThC.Tn[3].n19 XThC.Tn[3].t36 145.137
R22328 XThC.Tn[3].n22 XThC.Tn[3].t23 145.137
R22329 XThC.Tn[3].n25 XThC.Tn[3].t24 145.137
R22330 XThC.Tn[3].n28 XThC.Tn[3].t40 145.137
R22331 XThC.Tn[3].n31 XThC.Tn[3].t15 145.137
R22332 XThC.Tn[3].n34 XThC.Tn[3].t17 145.137
R22333 XThC.Tn[3].n37 XThC.Tn[3].t37 145.137
R22334 XThC.Tn[3].n40 XThC.Tn[3].t39 145.137
R22335 XThC.Tn[3].n43 XThC.Tn[3].t18 145.137
R22336 XThC.Tn[3].n46 XThC.Tn[3].t26 145.137
R22337 XThC.Tn[3].n49 XThC.Tn[3].t28 145.137
R22338 XThC.Tn[3].n52 XThC.Tn[3].t41 145.137
R22339 XThC.Tn[3].n55 XThC.Tn[3].t19 145.137
R22340 XThC.Tn[3].n6 XThC.Tn[3].n4 135.249
R22341 XThC.Tn[3].n9 XThC.Tn[3].n3 98.981
R22342 XThC.Tn[3].n6 XThC.Tn[3].n5 98.981
R22343 XThC.Tn[3].n8 XThC.Tn[3].n7 98.981
R22344 XThC.Tn[3].n8 XThC.Tn[3].n6 36.2672
R22345 XThC.Tn[3].n9 XThC.Tn[3].n8 36.2672
R22346 XThC.Tn[3].n58 XThC.Tn[3].n9 32.6405
R22347 XThC.Tn[3].n1 XThC.Tn[3].t7 26.5955
R22348 XThC.Tn[3].n1 XThC.Tn[3].t6 26.5955
R22349 XThC.Tn[3].n0 XThC.Tn[3].t5 26.5955
R22350 XThC.Tn[3].n0 XThC.Tn[3].t4 26.5955
R22351 XThC.Tn[3].n3 XThC.Tn[3].t1 24.9236
R22352 XThC.Tn[3].n3 XThC.Tn[3].t0 24.9236
R22353 XThC.Tn[3].n4 XThC.Tn[3].t11 24.9236
R22354 XThC.Tn[3].n4 XThC.Tn[3].t10 24.9236
R22355 XThC.Tn[3].n5 XThC.Tn[3].t9 24.9236
R22356 XThC.Tn[3].n5 XThC.Tn[3].t8 24.9236
R22357 XThC.Tn[3].n7 XThC.Tn[3].t3 24.9236
R22358 XThC.Tn[3].n7 XThC.Tn[3].t2 24.9236
R22359 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R22360 XThC.Tn[3] XThC.Tn[3].n58 6.7205
R22361 XThC.Tn[3].n58 XThC.Tn[3] 3.19574
R22362 XThC.Tn[3].n15 XThC.Tn[3] 0.931056
R22363 XThC.Tn[3].n18 XThC.Tn[3] 0.931056
R22364 XThC.Tn[3].n21 XThC.Tn[3] 0.931056
R22365 XThC.Tn[3].n24 XThC.Tn[3] 0.931056
R22366 XThC.Tn[3].n27 XThC.Tn[3] 0.931056
R22367 XThC.Tn[3].n30 XThC.Tn[3] 0.931056
R22368 XThC.Tn[3].n33 XThC.Tn[3] 0.931056
R22369 XThC.Tn[3].n36 XThC.Tn[3] 0.931056
R22370 XThC.Tn[3].n39 XThC.Tn[3] 0.931056
R22371 XThC.Tn[3].n42 XThC.Tn[3] 0.931056
R22372 XThC.Tn[3].n45 XThC.Tn[3] 0.931056
R22373 XThC.Tn[3].n48 XThC.Tn[3] 0.931056
R22374 XThC.Tn[3].n51 XThC.Tn[3] 0.931056
R22375 XThC.Tn[3].n54 XThC.Tn[3] 0.931056
R22376 XThC.Tn[3].n57 XThC.Tn[3] 0.931056
R22377 XThC.Tn[3] XThC.Tn[3].n12 0.396333
R22378 XThC.Tn[3] XThC.Tn[3].n15 0.396333
R22379 XThC.Tn[3] XThC.Tn[3].n18 0.396333
R22380 XThC.Tn[3] XThC.Tn[3].n21 0.396333
R22381 XThC.Tn[3] XThC.Tn[3].n24 0.396333
R22382 XThC.Tn[3] XThC.Tn[3].n27 0.396333
R22383 XThC.Tn[3] XThC.Tn[3].n30 0.396333
R22384 XThC.Tn[3] XThC.Tn[3].n33 0.396333
R22385 XThC.Tn[3] XThC.Tn[3].n36 0.396333
R22386 XThC.Tn[3] XThC.Tn[3].n39 0.396333
R22387 XThC.Tn[3] XThC.Tn[3].n42 0.396333
R22388 XThC.Tn[3] XThC.Tn[3].n45 0.396333
R22389 XThC.Tn[3] XThC.Tn[3].n48 0.396333
R22390 XThC.Tn[3] XThC.Tn[3].n51 0.396333
R22391 XThC.Tn[3] XThC.Tn[3].n54 0.396333
R22392 XThC.Tn[3] XThC.Tn[3].n57 0.396333
R22393 XThC.Tn[3].n11 XThC.Tn[3] 0.104667
R22394 XThC.Tn[3].n14 XThC.Tn[3] 0.104667
R22395 XThC.Tn[3].n17 XThC.Tn[3] 0.104667
R22396 XThC.Tn[3].n20 XThC.Tn[3] 0.104667
R22397 XThC.Tn[3].n23 XThC.Tn[3] 0.104667
R22398 XThC.Tn[3].n26 XThC.Tn[3] 0.104667
R22399 XThC.Tn[3].n29 XThC.Tn[3] 0.104667
R22400 XThC.Tn[3].n32 XThC.Tn[3] 0.104667
R22401 XThC.Tn[3].n35 XThC.Tn[3] 0.104667
R22402 XThC.Tn[3].n38 XThC.Tn[3] 0.104667
R22403 XThC.Tn[3].n41 XThC.Tn[3] 0.104667
R22404 XThC.Tn[3].n44 XThC.Tn[3] 0.104667
R22405 XThC.Tn[3].n47 XThC.Tn[3] 0.104667
R22406 XThC.Tn[3].n50 XThC.Tn[3] 0.104667
R22407 XThC.Tn[3].n53 XThC.Tn[3] 0.104667
R22408 XThC.Tn[3].n56 XThC.Tn[3] 0.104667
R22409 XThC.Tn[3].n11 XThC.Tn[3] 0.0309878
R22410 XThC.Tn[3].n14 XThC.Tn[3] 0.0309878
R22411 XThC.Tn[3].n17 XThC.Tn[3] 0.0309878
R22412 XThC.Tn[3].n20 XThC.Tn[3] 0.0309878
R22413 XThC.Tn[3].n23 XThC.Tn[3] 0.0309878
R22414 XThC.Tn[3].n26 XThC.Tn[3] 0.0309878
R22415 XThC.Tn[3].n29 XThC.Tn[3] 0.0309878
R22416 XThC.Tn[3].n32 XThC.Tn[3] 0.0309878
R22417 XThC.Tn[3].n35 XThC.Tn[3] 0.0309878
R22418 XThC.Tn[3].n38 XThC.Tn[3] 0.0309878
R22419 XThC.Tn[3].n41 XThC.Tn[3] 0.0309878
R22420 XThC.Tn[3].n44 XThC.Tn[3] 0.0309878
R22421 XThC.Tn[3].n47 XThC.Tn[3] 0.0309878
R22422 XThC.Tn[3].n50 XThC.Tn[3] 0.0309878
R22423 XThC.Tn[3].n53 XThC.Tn[3] 0.0309878
R22424 XThC.Tn[3].n56 XThC.Tn[3] 0.0309878
R22425 XThC.Tn[3].n12 XThC.Tn[3].n11 0.027939
R22426 XThC.Tn[3].n15 XThC.Tn[3].n14 0.027939
R22427 XThC.Tn[3].n18 XThC.Tn[3].n17 0.027939
R22428 XThC.Tn[3].n21 XThC.Tn[3].n20 0.027939
R22429 XThC.Tn[3].n24 XThC.Tn[3].n23 0.027939
R22430 XThC.Tn[3].n27 XThC.Tn[3].n26 0.027939
R22431 XThC.Tn[3].n30 XThC.Tn[3].n29 0.027939
R22432 XThC.Tn[3].n33 XThC.Tn[3].n32 0.027939
R22433 XThC.Tn[3].n36 XThC.Tn[3].n35 0.027939
R22434 XThC.Tn[3].n39 XThC.Tn[3].n38 0.027939
R22435 XThC.Tn[3].n42 XThC.Tn[3].n41 0.027939
R22436 XThC.Tn[3].n45 XThC.Tn[3].n44 0.027939
R22437 XThC.Tn[3].n48 XThC.Tn[3].n47 0.027939
R22438 XThC.Tn[3].n51 XThC.Tn[3].n50 0.027939
R22439 XThC.Tn[3].n54 XThC.Tn[3].n53 0.027939
R22440 XThC.Tn[3].n57 XThC.Tn[3].n56 0.027939
R22441 XThR.Tn[10].n5 XThR.Tn[10].n4 256.103
R22442 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R22443 XThR.Tn[10].n88 XThR.Tn[10].n87 241.847
R22444 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R22445 XThR.Tn[10].n5 XThR.Tn[10].n3 202.095
R22446 XThR.Tn[10].n88 XThR.Tn[10].n86 185
R22447 XThR.Tn[10] XThR.Tn[10].n79 161.363
R22448 XThR.Tn[10] XThR.Tn[10].n74 161.363
R22449 XThR.Tn[10] XThR.Tn[10].n69 161.363
R22450 XThR.Tn[10] XThR.Tn[10].n64 161.363
R22451 XThR.Tn[10] XThR.Tn[10].n59 161.363
R22452 XThR.Tn[10] XThR.Tn[10].n54 161.363
R22453 XThR.Tn[10] XThR.Tn[10].n49 161.363
R22454 XThR.Tn[10] XThR.Tn[10].n44 161.363
R22455 XThR.Tn[10] XThR.Tn[10].n39 161.363
R22456 XThR.Tn[10] XThR.Tn[10].n34 161.363
R22457 XThR.Tn[10] XThR.Tn[10].n29 161.363
R22458 XThR.Tn[10] XThR.Tn[10].n24 161.363
R22459 XThR.Tn[10] XThR.Tn[10].n19 161.363
R22460 XThR.Tn[10] XThR.Tn[10].n14 161.363
R22461 XThR.Tn[10] XThR.Tn[10].n9 161.363
R22462 XThR.Tn[10] XThR.Tn[10].n7 161.363
R22463 XThR.Tn[10].n81 XThR.Tn[10].n80 161.3
R22464 XThR.Tn[10].n76 XThR.Tn[10].n75 161.3
R22465 XThR.Tn[10].n71 XThR.Tn[10].n70 161.3
R22466 XThR.Tn[10].n66 XThR.Tn[10].n65 161.3
R22467 XThR.Tn[10].n61 XThR.Tn[10].n60 161.3
R22468 XThR.Tn[10].n56 XThR.Tn[10].n55 161.3
R22469 XThR.Tn[10].n51 XThR.Tn[10].n50 161.3
R22470 XThR.Tn[10].n46 XThR.Tn[10].n45 161.3
R22471 XThR.Tn[10].n41 XThR.Tn[10].n40 161.3
R22472 XThR.Tn[10].n36 XThR.Tn[10].n35 161.3
R22473 XThR.Tn[10].n31 XThR.Tn[10].n30 161.3
R22474 XThR.Tn[10].n26 XThR.Tn[10].n25 161.3
R22475 XThR.Tn[10].n21 XThR.Tn[10].n20 161.3
R22476 XThR.Tn[10].n16 XThR.Tn[10].n15 161.3
R22477 XThR.Tn[10].n11 XThR.Tn[10].n10 161.3
R22478 XThR.Tn[10].n79 XThR.Tn[10].t37 161.106
R22479 XThR.Tn[10].n74 XThR.Tn[10].t45 161.106
R22480 XThR.Tn[10].n69 XThR.Tn[10].t27 161.106
R22481 XThR.Tn[10].n64 XThR.Tn[10].t72 161.106
R22482 XThR.Tn[10].n59 XThR.Tn[10].t35 161.106
R22483 XThR.Tn[10].n54 XThR.Tn[10].t61 161.106
R22484 XThR.Tn[10].n49 XThR.Tn[10].t43 161.106
R22485 XThR.Tn[10].n44 XThR.Tn[10].t24 161.106
R22486 XThR.Tn[10].n39 XThR.Tn[10].t69 161.106
R22487 XThR.Tn[10].n34 XThR.Tn[10].t15 161.106
R22488 XThR.Tn[10].n29 XThR.Tn[10].t59 161.106
R22489 XThR.Tn[10].n24 XThR.Tn[10].t26 161.106
R22490 XThR.Tn[10].n19 XThR.Tn[10].t58 161.106
R22491 XThR.Tn[10].n14 XThR.Tn[10].t41 161.106
R22492 XThR.Tn[10].n9 XThR.Tn[10].t63 161.106
R22493 XThR.Tn[10].n7 XThR.Tn[10].t47 161.106
R22494 XThR.Tn[10].n80 XThR.Tn[10].t34 159.978
R22495 XThR.Tn[10].n75 XThR.Tn[10].t39 159.978
R22496 XThR.Tn[10].n70 XThR.Tn[10].t22 159.978
R22497 XThR.Tn[10].n65 XThR.Tn[10].t68 159.978
R22498 XThR.Tn[10].n60 XThR.Tn[10].t32 159.978
R22499 XThR.Tn[10].n55 XThR.Tn[10].t57 159.978
R22500 XThR.Tn[10].n50 XThR.Tn[10].t38 159.978
R22501 XThR.Tn[10].n45 XThR.Tn[10].t20 159.978
R22502 XThR.Tn[10].n40 XThR.Tn[10].t66 159.978
R22503 XThR.Tn[10].n35 XThR.Tn[10].t12 159.978
R22504 XThR.Tn[10].n30 XThR.Tn[10].t56 159.978
R22505 XThR.Tn[10].n25 XThR.Tn[10].t21 159.978
R22506 XThR.Tn[10].n20 XThR.Tn[10].t55 159.978
R22507 XThR.Tn[10].n15 XThR.Tn[10].t36 159.978
R22508 XThR.Tn[10].n10 XThR.Tn[10].t60 159.978
R22509 XThR.Tn[10].n79 XThR.Tn[10].t29 145.038
R22510 XThR.Tn[10].n74 XThR.Tn[10].t49 145.038
R22511 XThR.Tn[10].n69 XThR.Tn[10].t31 145.038
R22512 XThR.Tn[10].n64 XThR.Tn[10].t16 145.038
R22513 XThR.Tn[10].n59 XThR.Tn[10].t46 145.038
R22514 XThR.Tn[10].n54 XThR.Tn[10].t28 145.038
R22515 XThR.Tn[10].n49 XThR.Tn[10].t33 145.038
R22516 XThR.Tn[10].n44 XThR.Tn[10].t17 145.038
R22517 XThR.Tn[10].n39 XThR.Tn[10].t14 145.038
R22518 XThR.Tn[10].n34 XThR.Tn[10].t44 145.038
R22519 XThR.Tn[10].n29 XThR.Tn[10].t67 145.038
R22520 XThR.Tn[10].n24 XThR.Tn[10].t30 145.038
R22521 XThR.Tn[10].n19 XThR.Tn[10].t65 145.038
R22522 XThR.Tn[10].n14 XThR.Tn[10].t48 145.038
R22523 XThR.Tn[10].n9 XThR.Tn[10].t13 145.038
R22524 XThR.Tn[10].n7 XThR.Tn[10].t54 145.038
R22525 XThR.Tn[10].n80 XThR.Tn[10].t64 143.911
R22526 XThR.Tn[10].n75 XThR.Tn[10].t25 143.911
R22527 XThR.Tn[10].n70 XThR.Tn[10].t71 143.911
R22528 XThR.Tn[10].n65 XThR.Tn[10].t52 143.911
R22529 XThR.Tn[10].n60 XThR.Tn[10].t19 143.911
R22530 XThR.Tn[10].n55 XThR.Tn[10].t62 143.911
R22531 XThR.Tn[10].n50 XThR.Tn[10].t73 143.911
R22532 XThR.Tn[10].n45 XThR.Tn[10].t53 143.911
R22533 XThR.Tn[10].n40 XThR.Tn[10].t51 143.911
R22534 XThR.Tn[10].n35 XThR.Tn[10].t18 143.911
R22535 XThR.Tn[10].n30 XThR.Tn[10].t42 143.911
R22536 XThR.Tn[10].n25 XThR.Tn[10].t70 143.911
R22537 XThR.Tn[10].n20 XThR.Tn[10].t40 143.911
R22538 XThR.Tn[10].n15 XThR.Tn[10].t23 143.911
R22539 XThR.Tn[10].n10 XThR.Tn[10].t50 143.911
R22540 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R22541 XThR.Tn[10].n3 XThR.Tn[10].t6 26.5955
R22542 XThR.Tn[10].n3 XThR.Tn[10].t4 26.5955
R22543 XThR.Tn[10].n4 XThR.Tn[10].t7 26.5955
R22544 XThR.Tn[10].n4 XThR.Tn[10].t5 26.5955
R22545 XThR.Tn[10].n0 XThR.Tn[10].t10 26.5955
R22546 XThR.Tn[10].n0 XThR.Tn[10].t8 26.5955
R22547 XThR.Tn[10].n1 XThR.Tn[10].t11 26.5955
R22548 XThR.Tn[10].n1 XThR.Tn[10].t9 26.5955
R22549 XThR.Tn[10].n86 XThR.Tn[10].t0 24.9236
R22550 XThR.Tn[10].n86 XThR.Tn[10].t2 24.9236
R22551 XThR.Tn[10].n87 XThR.Tn[10].t1 24.9236
R22552 XThR.Tn[10].n87 XThR.Tn[10].t3 24.9236
R22553 XThR.Tn[10] XThR.Tn[10].n88 18.8943
R22554 XThR.Tn[10].n6 XThR.Tn[10].n5 13.5534
R22555 XThR.Tn[10].n85 XThR.Tn[10] 7.84567
R22556 XThR.Tn[10] XThR.Tn[10].n85 6.34069
R22557 XThR.Tn[10] XThR.Tn[10].n8 5.4407
R22558 XThR.Tn[10].n13 XThR.Tn[10].n12 4.5005
R22559 XThR.Tn[10].n18 XThR.Tn[10].n17 4.5005
R22560 XThR.Tn[10].n23 XThR.Tn[10].n22 4.5005
R22561 XThR.Tn[10].n28 XThR.Tn[10].n27 4.5005
R22562 XThR.Tn[10].n33 XThR.Tn[10].n32 4.5005
R22563 XThR.Tn[10].n38 XThR.Tn[10].n37 4.5005
R22564 XThR.Tn[10].n43 XThR.Tn[10].n42 4.5005
R22565 XThR.Tn[10].n48 XThR.Tn[10].n47 4.5005
R22566 XThR.Tn[10].n53 XThR.Tn[10].n52 4.5005
R22567 XThR.Tn[10].n58 XThR.Tn[10].n57 4.5005
R22568 XThR.Tn[10].n63 XThR.Tn[10].n62 4.5005
R22569 XThR.Tn[10].n68 XThR.Tn[10].n67 4.5005
R22570 XThR.Tn[10].n73 XThR.Tn[10].n72 4.5005
R22571 XThR.Tn[10].n78 XThR.Tn[10].n77 4.5005
R22572 XThR.Tn[10].n83 XThR.Tn[10].n82 4.5005
R22573 XThR.Tn[10].n84 XThR.Tn[10] 3.70586
R22574 XThR.Tn[10].n13 XThR.Tn[10] 2.52282
R22575 XThR.Tn[10].n18 XThR.Tn[10] 2.52282
R22576 XThR.Tn[10].n23 XThR.Tn[10] 2.52282
R22577 XThR.Tn[10].n28 XThR.Tn[10] 2.52282
R22578 XThR.Tn[10].n33 XThR.Tn[10] 2.52282
R22579 XThR.Tn[10].n38 XThR.Tn[10] 2.52282
R22580 XThR.Tn[10].n43 XThR.Tn[10] 2.52282
R22581 XThR.Tn[10].n48 XThR.Tn[10] 2.52282
R22582 XThR.Tn[10].n53 XThR.Tn[10] 2.52282
R22583 XThR.Tn[10].n58 XThR.Tn[10] 2.52282
R22584 XThR.Tn[10].n63 XThR.Tn[10] 2.52282
R22585 XThR.Tn[10].n68 XThR.Tn[10] 2.52282
R22586 XThR.Tn[10].n73 XThR.Tn[10] 2.52282
R22587 XThR.Tn[10].n78 XThR.Tn[10] 2.52282
R22588 XThR.Tn[10].n83 XThR.Tn[10] 2.52282
R22589 XThR.Tn[10].n85 XThR.Tn[10] 1.79489
R22590 XThR.Tn[10].n6 XThR.Tn[10] 1.50638
R22591 XThR.Tn[10] XThR.Tn[10].n6 1.19676
R22592 XThR.Tn[10].n81 XThR.Tn[10] 1.08677
R22593 XThR.Tn[10].n76 XThR.Tn[10] 1.08677
R22594 XThR.Tn[10].n71 XThR.Tn[10] 1.08677
R22595 XThR.Tn[10].n66 XThR.Tn[10] 1.08677
R22596 XThR.Tn[10].n61 XThR.Tn[10] 1.08677
R22597 XThR.Tn[10].n56 XThR.Tn[10] 1.08677
R22598 XThR.Tn[10].n51 XThR.Tn[10] 1.08677
R22599 XThR.Tn[10].n46 XThR.Tn[10] 1.08677
R22600 XThR.Tn[10].n41 XThR.Tn[10] 1.08677
R22601 XThR.Tn[10].n36 XThR.Tn[10] 1.08677
R22602 XThR.Tn[10].n31 XThR.Tn[10] 1.08677
R22603 XThR.Tn[10].n26 XThR.Tn[10] 1.08677
R22604 XThR.Tn[10].n21 XThR.Tn[10] 1.08677
R22605 XThR.Tn[10].n16 XThR.Tn[10] 1.08677
R22606 XThR.Tn[10].n11 XThR.Tn[10] 1.08677
R22607 XThR.Tn[10] XThR.Tn[10].n13 0.839786
R22608 XThR.Tn[10] XThR.Tn[10].n18 0.839786
R22609 XThR.Tn[10] XThR.Tn[10].n23 0.839786
R22610 XThR.Tn[10] XThR.Tn[10].n28 0.839786
R22611 XThR.Tn[10] XThR.Tn[10].n33 0.839786
R22612 XThR.Tn[10] XThR.Tn[10].n38 0.839786
R22613 XThR.Tn[10] XThR.Tn[10].n43 0.839786
R22614 XThR.Tn[10] XThR.Tn[10].n48 0.839786
R22615 XThR.Tn[10] XThR.Tn[10].n53 0.839786
R22616 XThR.Tn[10] XThR.Tn[10].n58 0.839786
R22617 XThR.Tn[10] XThR.Tn[10].n63 0.839786
R22618 XThR.Tn[10] XThR.Tn[10].n68 0.839786
R22619 XThR.Tn[10] XThR.Tn[10].n73 0.839786
R22620 XThR.Tn[10] XThR.Tn[10].n78 0.839786
R22621 XThR.Tn[10] XThR.Tn[10].n83 0.839786
R22622 XThR.Tn[10].n8 XThR.Tn[10] 0.499542
R22623 XThR.Tn[10].n82 XThR.Tn[10] 0.063
R22624 XThR.Tn[10].n77 XThR.Tn[10] 0.063
R22625 XThR.Tn[10].n72 XThR.Tn[10] 0.063
R22626 XThR.Tn[10].n67 XThR.Tn[10] 0.063
R22627 XThR.Tn[10].n62 XThR.Tn[10] 0.063
R22628 XThR.Tn[10].n57 XThR.Tn[10] 0.063
R22629 XThR.Tn[10].n52 XThR.Tn[10] 0.063
R22630 XThR.Tn[10].n47 XThR.Tn[10] 0.063
R22631 XThR.Tn[10].n42 XThR.Tn[10] 0.063
R22632 XThR.Tn[10].n37 XThR.Tn[10] 0.063
R22633 XThR.Tn[10].n32 XThR.Tn[10] 0.063
R22634 XThR.Tn[10].n27 XThR.Tn[10] 0.063
R22635 XThR.Tn[10].n22 XThR.Tn[10] 0.063
R22636 XThR.Tn[10].n17 XThR.Tn[10] 0.063
R22637 XThR.Tn[10].n12 XThR.Tn[10] 0.063
R22638 XThR.Tn[10].n84 XThR.Tn[10] 0.0540714
R22639 XThR.Tn[10] XThR.Tn[10].n84 0.038
R22640 XThR.Tn[10].n8 XThR.Tn[10] 0.0143889
R22641 XThR.Tn[10].n82 XThR.Tn[10].n81 0.00771154
R22642 XThR.Tn[10].n77 XThR.Tn[10].n76 0.00771154
R22643 XThR.Tn[10].n72 XThR.Tn[10].n71 0.00771154
R22644 XThR.Tn[10].n67 XThR.Tn[10].n66 0.00771154
R22645 XThR.Tn[10].n62 XThR.Tn[10].n61 0.00771154
R22646 XThR.Tn[10].n57 XThR.Tn[10].n56 0.00771154
R22647 XThR.Tn[10].n52 XThR.Tn[10].n51 0.00771154
R22648 XThR.Tn[10].n47 XThR.Tn[10].n46 0.00771154
R22649 XThR.Tn[10].n42 XThR.Tn[10].n41 0.00771154
R22650 XThR.Tn[10].n37 XThR.Tn[10].n36 0.00771154
R22651 XThR.Tn[10].n32 XThR.Tn[10].n31 0.00771154
R22652 XThR.Tn[10].n27 XThR.Tn[10].n26 0.00771154
R22653 XThR.Tn[10].n22 XThR.Tn[10].n21 0.00771154
R22654 XThR.Tn[10].n17 XThR.Tn[10].n16 0.00771154
R22655 XThR.Tn[10].n12 XThR.Tn[10].n11 0.00771154
R22656 XThC.Tn[14].n55 XThC.Tn[14].n54 256.104
R22657 XThC.Tn[14].n59 XThC.Tn[14].n58 243.679
R22658 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22659 XThC.Tn[14].n59 XThC.Tn[14].n57 205.28
R22660 XThC.Tn[14].n55 XThC.Tn[14].n53 202.095
R22661 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22662 XThC.Tn[14].n5 XThC.Tn[14].n3 161.406
R22663 XThC.Tn[14].n8 XThC.Tn[14].n6 161.406
R22664 XThC.Tn[14].n11 XThC.Tn[14].n9 161.406
R22665 XThC.Tn[14].n14 XThC.Tn[14].n12 161.406
R22666 XThC.Tn[14].n17 XThC.Tn[14].n15 161.406
R22667 XThC.Tn[14].n20 XThC.Tn[14].n18 161.406
R22668 XThC.Tn[14].n23 XThC.Tn[14].n21 161.406
R22669 XThC.Tn[14].n26 XThC.Tn[14].n24 161.406
R22670 XThC.Tn[14].n29 XThC.Tn[14].n27 161.406
R22671 XThC.Tn[14].n32 XThC.Tn[14].n30 161.406
R22672 XThC.Tn[14].n35 XThC.Tn[14].n33 161.406
R22673 XThC.Tn[14].n38 XThC.Tn[14].n36 161.406
R22674 XThC.Tn[14].n41 XThC.Tn[14].n39 161.406
R22675 XThC.Tn[14].n44 XThC.Tn[14].n42 161.406
R22676 XThC.Tn[14].n47 XThC.Tn[14].n45 161.406
R22677 XThC.Tn[14].n50 XThC.Tn[14].n48 161.406
R22678 XThC.Tn[14].n3 XThC.Tn[14].t38 161.202
R22679 XThC.Tn[14].n6 XThC.Tn[14].t22 161.202
R22680 XThC.Tn[14].n9 XThC.Tn[14].t25 161.202
R22681 XThC.Tn[14].n12 XThC.Tn[14].t26 161.202
R22682 XThC.Tn[14].n15 XThC.Tn[14].t14 161.202
R22683 XThC.Tn[14].n18 XThC.Tn[14].t17 161.202
R22684 XThC.Tn[14].n21 XThC.Tn[14].t31 161.202
R22685 XThC.Tn[14].n24 XThC.Tn[14].t39 161.202
R22686 XThC.Tn[14].n27 XThC.Tn[14].t41 161.202
R22687 XThC.Tn[14].n30 XThC.Tn[14].t27 161.202
R22688 XThC.Tn[14].n33 XThC.Tn[14].t30 161.202
R22689 XThC.Tn[14].n36 XThC.Tn[14].t42 161.202
R22690 XThC.Tn[14].n39 XThC.Tn[14].t19 161.202
R22691 XThC.Tn[14].n42 XThC.Tn[14].t21 161.202
R22692 XThC.Tn[14].n45 XThC.Tn[14].t33 161.202
R22693 XThC.Tn[14].n48 XThC.Tn[14].t12 161.202
R22694 XThC.Tn[14].n3 XThC.Tn[14].t43 145.137
R22695 XThC.Tn[14].n6 XThC.Tn[14].t29 145.137
R22696 XThC.Tn[14].n9 XThC.Tn[14].t32 145.137
R22697 XThC.Tn[14].n12 XThC.Tn[14].t34 145.137
R22698 XThC.Tn[14].n15 XThC.Tn[14].t20 145.137
R22699 XThC.Tn[14].n18 XThC.Tn[14].t23 145.137
R22700 XThC.Tn[14].n21 XThC.Tn[14].t37 145.137
R22701 XThC.Tn[14].n24 XThC.Tn[14].t13 145.137
R22702 XThC.Tn[14].n27 XThC.Tn[14].t15 145.137
R22703 XThC.Tn[14].n30 XThC.Tn[14].t35 145.137
R22704 XThC.Tn[14].n33 XThC.Tn[14].t36 145.137
R22705 XThC.Tn[14].n36 XThC.Tn[14].t16 145.137
R22706 XThC.Tn[14].n39 XThC.Tn[14].t24 145.137
R22707 XThC.Tn[14].n42 XThC.Tn[14].t28 145.137
R22708 XThC.Tn[14].n45 XThC.Tn[14].t40 145.137
R22709 XThC.Tn[14].n48 XThC.Tn[14].t18 145.137
R22710 XThC.Tn[14].n53 XThC.Tn[14].t8 26.5955
R22711 XThC.Tn[14].n53 XThC.Tn[14].t9 26.5955
R22712 XThC.Tn[14].n54 XThC.Tn[14].t11 26.5955
R22713 XThC.Tn[14].n54 XThC.Tn[14].t10 26.5955
R22714 XThC.Tn[14].n57 XThC.Tn[14].t1 26.5955
R22715 XThC.Tn[14].n57 XThC.Tn[14].t0 26.5955
R22716 XThC.Tn[14].n58 XThC.Tn[14].t3 26.5955
R22717 XThC.Tn[14].n58 XThC.Tn[14].t2 26.5955
R22718 XThC.Tn[14].n1 XThC.Tn[14].t5 24.9236
R22719 XThC.Tn[14].n1 XThC.Tn[14].t7 24.9236
R22720 XThC.Tn[14].n0 XThC.Tn[14].t4 24.9236
R22721 XThC.Tn[14].n0 XThC.Tn[14].t6 24.9236
R22722 XThC.Tn[14] XThC.Tn[14].n59 22.9652
R22723 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22724 XThC.Tn[14].n56 XThC.Tn[14].n55 13.9299
R22725 XThC.Tn[14] XThC.Tn[14].n56 13.9299
R22726 XThC.Tn[14].n51 XThC.Tn[14] 5.65386
R22727 XThC.Tn[14].n52 XThC.Tn[14].n51 5.13312
R22728 XThC.Tn[14].n56 XThC.Tn[14].n52 2.99115
R22729 XThC.Tn[14].n56 XThC.Tn[14] 2.87153
R22730 XThC.Tn[14].n52 XThC.Tn[14] 2.2734
R22731 XThC.Tn[14].n8 XThC.Tn[14] 0.931056
R22732 XThC.Tn[14].n11 XThC.Tn[14] 0.931056
R22733 XThC.Tn[14].n14 XThC.Tn[14] 0.931056
R22734 XThC.Tn[14].n17 XThC.Tn[14] 0.931056
R22735 XThC.Tn[14].n20 XThC.Tn[14] 0.931056
R22736 XThC.Tn[14].n23 XThC.Tn[14] 0.931056
R22737 XThC.Tn[14].n26 XThC.Tn[14] 0.931056
R22738 XThC.Tn[14].n29 XThC.Tn[14] 0.931056
R22739 XThC.Tn[14].n32 XThC.Tn[14] 0.931056
R22740 XThC.Tn[14].n35 XThC.Tn[14] 0.931056
R22741 XThC.Tn[14].n38 XThC.Tn[14] 0.931056
R22742 XThC.Tn[14].n41 XThC.Tn[14] 0.931056
R22743 XThC.Tn[14].n44 XThC.Tn[14] 0.931056
R22744 XThC.Tn[14].n47 XThC.Tn[14] 0.931056
R22745 XThC.Tn[14].n50 XThC.Tn[14] 0.931056
R22746 XThC.Tn[14] XThC.Tn[14].n5 0.396333
R22747 XThC.Tn[14] XThC.Tn[14].n8 0.396333
R22748 XThC.Tn[14] XThC.Tn[14].n11 0.396333
R22749 XThC.Tn[14] XThC.Tn[14].n14 0.396333
R22750 XThC.Tn[14] XThC.Tn[14].n17 0.396333
R22751 XThC.Tn[14] XThC.Tn[14].n20 0.396333
R22752 XThC.Tn[14] XThC.Tn[14].n23 0.396333
R22753 XThC.Tn[14] XThC.Tn[14].n26 0.396333
R22754 XThC.Tn[14] XThC.Tn[14].n29 0.396333
R22755 XThC.Tn[14] XThC.Tn[14].n32 0.396333
R22756 XThC.Tn[14] XThC.Tn[14].n35 0.396333
R22757 XThC.Tn[14] XThC.Tn[14].n38 0.396333
R22758 XThC.Tn[14] XThC.Tn[14].n41 0.396333
R22759 XThC.Tn[14] XThC.Tn[14].n44 0.396333
R22760 XThC.Tn[14] XThC.Tn[14].n47 0.396333
R22761 XThC.Tn[14] XThC.Tn[14].n50 0.396333
R22762 XThC.Tn[14].n4 XThC.Tn[14] 0.104667
R22763 XThC.Tn[14].n7 XThC.Tn[14] 0.104667
R22764 XThC.Tn[14].n10 XThC.Tn[14] 0.104667
R22765 XThC.Tn[14].n13 XThC.Tn[14] 0.104667
R22766 XThC.Tn[14].n16 XThC.Tn[14] 0.104667
R22767 XThC.Tn[14].n19 XThC.Tn[14] 0.104667
R22768 XThC.Tn[14].n22 XThC.Tn[14] 0.104667
R22769 XThC.Tn[14].n25 XThC.Tn[14] 0.104667
R22770 XThC.Tn[14].n28 XThC.Tn[14] 0.104667
R22771 XThC.Tn[14].n31 XThC.Tn[14] 0.104667
R22772 XThC.Tn[14].n34 XThC.Tn[14] 0.104667
R22773 XThC.Tn[14].n37 XThC.Tn[14] 0.104667
R22774 XThC.Tn[14].n40 XThC.Tn[14] 0.104667
R22775 XThC.Tn[14].n43 XThC.Tn[14] 0.104667
R22776 XThC.Tn[14].n46 XThC.Tn[14] 0.104667
R22777 XThC.Tn[14].n49 XThC.Tn[14] 0.104667
R22778 XThC.Tn[14].n4 XThC.Tn[14] 0.0309878
R22779 XThC.Tn[14].n7 XThC.Tn[14] 0.0309878
R22780 XThC.Tn[14].n10 XThC.Tn[14] 0.0309878
R22781 XThC.Tn[14].n13 XThC.Tn[14] 0.0309878
R22782 XThC.Tn[14].n16 XThC.Tn[14] 0.0309878
R22783 XThC.Tn[14].n19 XThC.Tn[14] 0.0309878
R22784 XThC.Tn[14].n22 XThC.Tn[14] 0.0309878
R22785 XThC.Tn[14].n25 XThC.Tn[14] 0.0309878
R22786 XThC.Tn[14].n28 XThC.Tn[14] 0.0309878
R22787 XThC.Tn[14].n31 XThC.Tn[14] 0.0309878
R22788 XThC.Tn[14].n34 XThC.Tn[14] 0.0309878
R22789 XThC.Tn[14].n37 XThC.Tn[14] 0.0309878
R22790 XThC.Tn[14].n40 XThC.Tn[14] 0.0309878
R22791 XThC.Tn[14].n43 XThC.Tn[14] 0.0309878
R22792 XThC.Tn[14].n46 XThC.Tn[14] 0.0309878
R22793 XThC.Tn[14].n49 XThC.Tn[14] 0.0309878
R22794 XThC.Tn[14].n5 XThC.Tn[14].n4 0.027939
R22795 XThC.Tn[14].n8 XThC.Tn[14].n7 0.027939
R22796 XThC.Tn[14].n11 XThC.Tn[14].n10 0.027939
R22797 XThC.Tn[14].n14 XThC.Tn[14].n13 0.027939
R22798 XThC.Tn[14].n17 XThC.Tn[14].n16 0.027939
R22799 XThC.Tn[14].n20 XThC.Tn[14].n19 0.027939
R22800 XThC.Tn[14].n23 XThC.Tn[14].n22 0.027939
R22801 XThC.Tn[14].n26 XThC.Tn[14].n25 0.027939
R22802 XThC.Tn[14].n29 XThC.Tn[14].n28 0.027939
R22803 XThC.Tn[14].n32 XThC.Tn[14].n31 0.027939
R22804 XThC.Tn[14].n35 XThC.Tn[14].n34 0.027939
R22805 XThC.Tn[14].n38 XThC.Tn[14].n37 0.027939
R22806 XThC.Tn[14].n41 XThC.Tn[14].n40 0.027939
R22807 XThC.Tn[14].n44 XThC.Tn[14].n43 0.027939
R22808 XThC.Tn[14].n47 XThC.Tn[14].n46 0.027939
R22809 XThC.Tn[14].n50 XThC.Tn[14].n49 0.027939
R22810 XThC.Tn[14].n51 XThC.Tn[14] 0.00250754
R22811 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R22812 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R22813 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R22814 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R22815 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R22816 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R22817 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R22818 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R22819 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R22820 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22821 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22822 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22823 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22824 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22825 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22826 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22827 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22828 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22829 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22830 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22831 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22832 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22833 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22834 XThC.XTB1.Y.n0 XThC.XTB1.Y.t1 132.067
R22835 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22836 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22837 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22838 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22839 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22840 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22841 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22842 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22843 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22844 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22845 XThC.XTB1.Y.n2 XThC.XTB1.Y.t2 26.5955
R22846 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22847 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22848 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22849 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22850 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22851 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22852 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22853 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22854 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22855 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22856 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22857 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22858 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22859 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22860 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22861 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22862 XThC.Tn[8].n56 XThC.Tn[8].n55 256.104
R22863 XThC.Tn[8].n60 XThC.Tn[8].n59 243.679
R22864 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22865 XThC.Tn[8].n60 XThC.Tn[8].n58 205.28
R22866 XThC.Tn[8].n56 XThC.Tn[8].n54 202.095
R22867 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22868 XThC.Tn[8].n5 XThC.Tn[8].n3 161.406
R22869 XThC.Tn[8].n8 XThC.Tn[8].n6 161.406
R22870 XThC.Tn[8].n11 XThC.Tn[8].n9 161.406
R22871 XThC.Tn[8].n14 XThC.Tn[8].n12 161.406
R22872 XThC.Tn[8].n17 XThC.Tn[8].n15 161.406
R22873 XThC.Tn[8].n20 XThC.Tn[8].n18 161.406
R22874 XThC.Tn[8].n23 XThC.Tn[8].n21 161.406
R22875 XThC.Tn[8].n26 XThC.Tn[8].n24 161.406
R22876 XThC.Tn[8].n29 XThC.Tn[8].n27 161.406
R22877 XThC.Tn[8].n32 XThC.Tn[8].n30 161.406
R22878 XThC.Tn[8].n35 XThC.Tn[8].n33 161.406
R22879 XThC.Tn[8].n38 XThC.Tn[8].n36 161.406
R22880 XThC.Tn[8].n41 XThC.Tn[8].n39 161.406
R22881 XThC.Tn[8].n44 XThC.Tn[8].n42 161.406
R22882 XThC.Tn[8].n47 XThC.Tn[8].n45 161.406
R22883 XThC.Tn[8].n50 XThC.Tn[8].n48 161.406
R22884 XThC.Tn[8].n3 XThC.Tn[8].t41 161.202
R22885 XThC.Tn[8].n6 XThC.Tn[8].t26 161.202
R22886 XThC.Tn[8].n9 XThC.Tn[8].t28 161.202
R22887 XThC.Tn[8].n12 XThC.Tn[8].t30 161.202
R22888 XThC.Tn[8].n15 XThC.Tn[8].t19 161.202
R22889 XThC.Tn[8].n18 XThC.Tn[8].t20 161.202
R22890 XThC.Tn[8].n21 XThC.Tn[8].t33 161.202
R22891 XThC.Tn[8].n24 XThC.Tn[8].t42 161.202
R22892 XThC.Tn[8].n27 XThC.Tn[8].t12 161.202
R22893 XThC.Tn[8].n30 XThC.Tn[8].t31 161.202
R22894 XThC.Tn[8].n33 XThC.Tn[8].t32 161.202
R22895 XThC.Tn[8].n36 XThC.Tn[8].t13 161.202
R22896 XThC.Tn[8].n39 XThC.Tn[8].t21 161.202
R22897 XThC.Tn[8].n42 XThC.Tn[8].t24 161.202
R22898 XThC.Tn[8].n45 XThC.Tn[8].t37 161.202
R22899 XThC.Tn[8].n48 XThC.Tn[8].t15 161.202
R22900 XThC.Tn[8].n3 XThC.Tn[8].t43 145.137
R22901 XThC.Tn[8].n6 XThC.Tn[8].t29 145.137
R22902 XThC.Tn[8].n9 XThC.Tn[8].t34 145.137
R22903 XThC.Tn[8].n12 XThC.Tn[8].t35 145.137
R22904 XThC.Tn[8].n15 XThC.Tn[8].t22 145.137
R22905 XThC.Tn[8].n18 XThC.Tn[8].t23 145.137
R22906 XThC.Tn[8].n21 XThC.Tn[8].t39 145.137
R22907 XThC.Tn[8].n24 XThC.Tn[8].t14 145.137
R22908 XThC.Tn[8].n27 XThC.Tn[8].t16 145.137
R22909 XThC.Tn[8].n30 XThC.Tn[8].t36 145.137
R22910 XThC.Tn[8].n33 XThC.Tn[8].t38 145.137
R22911 XThC.Tn[8].n36 XThC.Tn[8].t17 145.137
R22912 XThC.Tn[8].n39 XThC.Tn[8].t25 145.137
R22913 XThC.Tn[8].n42 XThC.Tn[8].t27 145.137
R22914 XThC.Tn[8].n45 XThC.Tn[8].t40 145.137
R22915 XThC.Tn[8].n48 XThC.Tn[8].t18 145.137
R22916 XThC.Tn[8].n54 XThC.Tn[8].t9 26.5955
R22917 XThC.Tn[8].n54 XThC.Tn[8].t10 26.5955
R22918 XThC.Tn[8].n55 XThC.Tn[8].t8 26.5955
R22919 XThC.Tn[8].n55 XThC.Tn[8].t11 26.5955
R22920 XThC.Tn[8].n58 XThC.Tn[8].t2 26.5955
R22921 XThC.Tn[8].n58 XThC.Tn[8].t1 26.5955
R22922 XThC.Tn[8].n59 XThC.Tn[8].t0 26.5955
R22923 XThC.Tn[8].n59 XThC.Tn[8].t3 26.5955
R22924 XThC.Tn[8].n1 XThC.Tn[8].t7 24.9236
R22925 XThC.Tn[8].n1 XThC.Tn[8].t6 24.9236
R22926 XThC.Tn[8].n0 XThC.Tn[8].t5 24.9236
R22927 XThC.Tn[8].n0 XThC.Tn[8].t4 24.9236
R22928 XThC.Tn[8] XThC.Tn[8].n60 22.9652
R22929 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22930 XThC.Tn[8].n57 XThC.Tn[8].n56 13.9299
R22931 XThC.Tn[8] XThC.Tn[8].n57 13.9299
R22932 XThC.Tn[8].n53 XThC.Tn[8].n52 5.09639
R22933 XThC.Tn[8].n57 XThC.Tn[8].n53 2.99115
R22934 XThC.Tn[8].n57 XThC.Tn[8] 2.87153
R22935 XThC.Tn[8].n53 XThC.Tn[8] 2.2734
R22936 XThC.Tn[8].n51 XThC.Tn[8] 1.14336
R22937 XThC.Tn[8].n8 XThC.Tn[8] 0.931056
R22938 XThC.Tn[8].n11 XThC.Tn[8] 0.931056
R22939 XThC.Tn[8].n14 XThC.Tn[8] 0.931056
R22940 XThC.Tn[8].n17 XThC.Tn[8] 0.931056
R22941 XThC.Tn[8].n20 XThC.Tn[8] 0.931056
R22942 XThC.Tn[8].n23 XThC.Tn[8] 0.931056
R22943 XThC.Tn[8].n26 XThC.Tn[8] 0.931056
R22944 XThC.Tn[8].n29 XThC.Tn[8] 0.931056
R22945 XThC.Tn[8].n32 XThC.Tn[8] 0.931056
R22946 XThC.Tn[8].n35 XThC.Tn[8] 0.931056
R22947 XThC.Tn[8].n38 XThC.Tn[8] 0.931056
R22948 XThC.Tn[8].n41 XThC.Tn[8] 0.931056
R22949 XThC.Tn[8].n44 XThC.Tn[8] 0.931056
R22950 XThC.Tn[8].n47 XThC.Tn[8] 0.931056
R22951 XThC.Tn[8].n50 XThC.Tn[8] 0.931056
R22952 XThC.Tn[8] XThC.Tn[8].n5 0.396333
R22953 XThC.Tn[8] XThC.Tn[8].n8 0.396333
R22954 XThC.Tn[8] XThC.Tn[8].n11 0.396333
R22955 XThC.Tn[8] XThC.Tn[8].n14 0.396333
R22956 XThC.Tn[8] XThC.Tn[8].n17 0.396333
R22957 XThC.Tn[8] XThC.Tn[8].n20 0.396333
R22958 XThC.Tn[8] XThC.Tn[8].n23 0.396333
R22959 XThC.Tn[8] XThC.Tn[8].n26 0.396333
R22960 XThC.Tn[8] XThC.Tn[8].n29 0.396333
R22961 XThC.Tn[8] XThC.Tn[8].n32 0.396333
R22962 XThC.Tn[8] XThC.Tn[8].n35 0.396333
R22963 XThC.Tn[8] XThC.Tn[8].n38 0.396333
R22964 XThC.Tn[8] XThC.Tn[8].n41 0.396333
R22965 XThC.Tn[8] XThC.Tn[8].n44 0.396333
R22966 XThC.Tn[8] XThC.Tn[8].n47 0.396333
R22967 XThC.Tn[8] XThC.Tn[8].n50 0.396333
R22968 XThC.Tn[8].n52 XThC.Tn[8].n51 0.166125
R22969 XThC.Tn[8].n4 XThC.Tn[8] 0.104667
R22970 XThC.Tn[8].n7 XThC.Tn[8] 0.104667
R22971 XThC.Tn[8].n10 XThC.Tn[8] 0.104667
R22972 XThC.Tn[8].n13 XThC.Tn[8] 0.104667
R22973 XThC.Tn[8].n16 XThC.Tn[8] 0.104667
R22974 XThC.Tn[8].n19 XThC.Tn[8] 0.104667
R22975 XThC.Tn[8].n22 XThC.Tn[8] 0.104667
R22976 XThC.Tn[8].n25 XThC.Tn[8] 0.104667
R22977 XThC.Tn[8].n28 XThC.Tn[8] 0.104667
R22978 XThC.Tn[8].n31 XThC.Tn[8] 0.104667
R22979 XThC.Tn[8].n34 XThC.Tn[8] 0.104667
R22980 XThC.Tn[8].n37 XThC.Tn[8] 0.104667
R22981 XThC.Tn[8].n40 XThC.Tn[8] 0.104667
R22982 XThC.Tn[8].n43 XThC.Tn[8] 0.104667
R22983 XThC.Tn[8].n46 XThC.Tn[8] 0.104667
R22984 XThC.Tn[8].n49 XThC.Tn[8] 0.104667
R22985 XThC.Tn[8].n52 XThC.Tn[8] 0.0389615
R22986 XThC.Tn[8].n51 XThC.Tn[8] 0.038
R22987 XThC.Tn[8].n4 XThC.Tn[8] 0.0309878
R22988 XThC.Tn[8].n7 XThC.Tn[8] 0.0309878
R22989 XThC.Tn[8].n10 XThC.Tn[8] 0.0309878
R22990 XThC.Tn[8].n13 XThC.Tn[8] 0.0309878
R22991 XThC.Tn[8].n16 XThC.Tn[8] 0.0309878
R22992 XThC.Tn[8].n19 XThC.Tn[8] 0.0309878
R22993 XThC.Tn[8].n22 XThC.Tn[8] 0.0309878
R22994 XThC.Tn[8].n25 XThC.Tn[8] 0.0309878
R22995 XThC.Tn[8].n28 XThC.Tn[8] 0.0309878
R22996 XThC.Tn[8].n31 XThC.Tn[8] 0.0309878
R22997 XThC.Tn[8].n34 XThC.Tn[8] 0.0309878
R22998 XThC.Tn[8].n37 XThC.Tn[8] 0.0309878
R22999 XThC.Tn[8].n40 XThC.Tn[8] 0.0309878
R23000 XThC.Tn[8].n43 XThC.Tn[8] 0.0309878
R23001 XThC.Tn[8].n46 XThC.Tn[8] 0.0309878
R23002 XThC.Tn[8].n49 XThC.Tn[8] 0.0309878
R23003 XThC.Tn[8].n5 XThC.Tn[8].n4 0.027939
R23004 XThC.Tn[8].n8 XThC.Tn[8].n7 0.027939
R23005 XThC.Tn[8].n11 XThC.Tn[8].n10 0.027939
R23006 XThC.Tn[8].n14 XThC.Tn[8].n13 0.027939
R23007 XThC.Tn[8].n17 XThC.Tn[8].n16 0.027939
R23008 XThC.Tn[8].n20 XThC.Tn[8].n19 0.027939
R23009 XThC.Tn[8].n23 XThC.Tn[8].n22 0.027939
R23010 XThC.Tn[8].n26 XThC.Tn[8].n25 0.027939
R23011 XThC.Tn[8].n29 XThC.Tn[8].n28 0.027939
R23012 XThC.Tn[8].n32 XThC.Tn[8].n31 0.027939
R23013 XThC.Tn[8].n35 XThC.Tn[8].n34 0.027939
R23014 XThC.Tn[8].n38 XThC.Tn[8].n37 0.027939
R23015 XThC.Tn[8].n41 XThC.Tn[8].n40 0.027939
R23016 XThC.Tn[8].n44 XThC.Tn[8].n43 0.027939
R23017 XThC.Tn[8].n47 XThC.Tn[8].n46 0.027939
R23018 XThC.Tn[8].n50 XThC.Tn[8].n49 0.027939
R23019 XThR.Tn[1].n2 XThR.Tn[1].n1 332.332
R23020 XThR.Tn[1].n2 XThR.Tn[1].n0 296.493
R23021 XThR.Tn[1] XThR.Tn[1].n82 161.363
R23022 XThR.Tn[1] XThR.Tn[1].n77 161.363
R23023 XThR.Tn[1] XThR.Tn[1].n72 161.363
R23024 XThR.Tn[1] XThR.Tn[1].n67 161.363
R23025 XThR.Tn[1] XThR.Tn[1].n62 161.363
R23026 XThR.Tn[1] XThR.Tn[1].n57 161.363
R23027 XThR.Tn[1] XThR.Tn[1].n52 161.363
R23028 XThR.Tn[1] XThR.Tn[1].n47 161.363
R23029 XThR.Tn[1] XThR.Tn[1].n42 161.363
R23030 XThR.Tn[1] XThR.Tn[1].n37 161.363
R23031 XThR.Tn[1] XThR.Tn[1].n32 161.363
R23032 XThR.Tn[1] XThR.Tn[1].n27 161.363
R23033 XThR.Tn[1] XThR.Tn[1].n22 161.363
R23034 XThR.Tn[1] XThR.Tn[1].n17 161.363
R23035 XThR.Tn[1] XThR.Tn[1].n12 161.363
R23036 XThR.Tn[1] XThR.Tn[1].n10 161.363
R23037 XThR.Tn[1].n84 XThR.Tn[1].n83 161.3
R23038 XThR.Tn[1].n79 XThR.Tn[1].n78 161.3
R23039 XThR.Tn[1].n74 XThR.Tn[1].n73 161.3
R23040 XThR.Tn[1].n69 XThR.Tn[1].n68 161.3
R23041 XThR.Tn[1].n64 XThR.Tn[1].n63 161.3
R23042 XThR.Tn[1].n59 XThR.Tn[1].n58 161.3
R23043 XThR.Tn[1].n54 XThR.Tn[1].n53 161.3
R23044 XThR.Tn[1].n49 XThR.Tn[1].n48 161.3
R23045 XThR.Tn[1].n44 XThR.Tn[1].n43 161.3
R23046 XThR.Tn[1].n39 XThR.Tn[1].n38 161.3
R23047 XThR.Tn[1].n34 XThR.Tn[1].n33 161.3
R23048 XThR.Tn[1].n29 XThR.Tn[1].n28 161.3
R23049 XThR.Tn[1].n24 XThR.Tn[1].n23 161.3
R23050 XThR.Tn[1].n19 XThR.Tn[1].n18 161.3
R23051 XThR.Tn[1].n14 XThR.Tn[1].n13 161.3
R23052 XThR.Tn[1].n82 XThR.Tn[1].t70 161.106
R23053 XThR.Tn[1].n77 XThR.Tn[1].t14 161.106
R23054 XThR.Tn[1].n72 XThR.Tn[1].t56 161.106
R23055 XThR.Tn[1].n67 XThR.Tn[1].t42 161.106
R23056 XThR.Tn[1].n62 XThR.Tn[1].t68 161.106
R23057 XThR.Tn[1].n57 XThR.Tn[1].t31 161.106
R23058 XThR.Tn[1].n52 XThR.Tn[1].t12 161.106
R23059 XThR.Tn[1].n47 XThR.Tn[1].t54 161.106
R23060 XThR.Tn[1].n42 XThR.Tn[1].t41 161.106
R23061 XThR.Tn[1].n37 XThR.Tn[1].t46 161.106
R23062 XThR.Tn[1].n32 XThR.Tn[1].t29 161.106
R23063 XThR.Tn[1].n27 XThR.Tn[1].t55 161.106
R23064 XThR.Tn[1].n22 XThR.Tn[1].t28 161.106
R23065 XThR.Tn[1].n17 XThR.Tn[1].t73 161.106
R23066 XThR.Tn[1].n12 XThR.Tn[1].t34 161.106
R23067 XThR.Tn[1].n10 XThR.Tn[1].t18 161.106
R23068 XThR.Tn[1].n83 XThR.Tn[1].t66 159.978
R23069 XThR.Tn[1].n78 XThR.Tn[1].t72 159.978
R23070 XThR.Tn[1].n73 XThR.Tn[1].t52 159.978
R23071 XThR.Tn[1].n68 XThR.Tn[1].t39 159.978
R23072 XThR.Tn[1].n63 XThR.Tn[1].t63 159.978
R23073 XThR.Tn[1].n58 XThR.Tn[1].t27 159.978
R23074 XThR.Tn[1].n53 XThR.Tn[1].t71 159.978
R23075 XThR.Tn[1].n48 XThR.Tn[1].t49 159.978
R23076 XThR.Tn[1].n43 XThR.Tn[1].t36 159.978
R23077 XThR.Tn[1].n38 XThR.Tn[1].t43 159.978
R23078 XThR.Tn[1].n33 XThR.Tn[1].t26 159.978
R23079 XThR.Tn[1].n28 XThR.Tn[1].t51 159.978
R23080 XThR.Tn[1].n23 XThR.Tn[1].t25 159.978
R23081 XThR.Tn[1].n18 XThR.Tn[1].t69 159.978
R23082 XThR.Tn[1].n13 XThR.Tn[1].t30 159.978
R23083 XThR.Tn[1].n82 XThR.Tn[1].t58 145.038
R23084 XThR.Tn[1].n77 XThR.Tn[1].t20 145.038
R23085 XThR.Tn[1].n72 XThR.Tn[1].t62 145.038
R23086 XThR.Tn[1].n67 XThR.Tn[1].t47 145.038
R23087 XThR.Tn[1].n62 XThR.Tn[1].t15 145.038
R23088 XThR.Tn[1].n57 XThR.Tn[1].t57 145.038
R23089 XThR.Tn[1].n52 XThR.Tn[1].t64 145.038
R23090 XThR.Tn[1].n47 XThR.Tn[1].t48 145.038
R23091 XThR.Tn[1].n42 XThR.Tn[1].t45 145.038
R23092 XThR.Tn[1].n37 XThR.Tn[1].t13 145.038
R23093 XThR.Tn[1].n32 XThR.Tn[1].t37 145.038
R23094 XThR.Tn[1].n27 XThR.Tn[1].t59 145.038
R23095 XThR.Tn[1].n22 XThR.Tn[1].t35 145.038
R23096 XThR.Tn[1].n17 XThR.Tn[1].t19 145.038
R23097 XThR.Tn[1].n12 XThR.Tn[1].t44 145.038
R23098 XThR.Tn[1].n10 XThR.Tn[1].t24 145.038
R23099 XThR.Tn[1].n83 XThR.Tn[1].t17 143.911
R23100 XThR.Tn[1].n78 XThR.Tn[1].t40 143.911
R23101 XThR.Tn[1].n73 XThR.Tn[1].t22 143.911
R23102 XThR.Tn[1].n68 XThR.Tn[1].t65 143.911
R23103 XThR.Tn[1].n63 XThR.Tn[1].t33 143.911
R23104 XThR.Tn[1].n58 XThR.Tn[1].t16 143.911
R23105 XThR.Tn[1].n53 XThR.Tn[1].t23 143.911
R23106 XThR.Tn[1].n48 XThR.Tn[1].t67 143.911
R23107 XThR.Tn[1].n43 XThR.Tn[1].t60 143.911
R23108 XThR.Tn[1].n38 XThR.Tn[1].t32 143.911
R23109 XThR.Tn[1].n33 XThR.Tn[1].t53 143.911
R23110 XThR.Tn[1].n28 XThR.Tn[1].t21 143.911
R23111 XThR.Tn[1].n23 XThR.Tn[1].t50 143.911
R23112 XThR.Tn[1].n18 XThR.Tn[1].t38 143.911
R23113 XThR.Tn[1].n13 XThR.Tn[1].t61 143.911
R23114 XThR.Tn[1].n7 XThR.Tn[1].n6 135.249
R23115 XThR.Tn[1].n9 XThR.Tn[1].n3 98.981
R23116 XThR.Tn[1].n8 XThR.Tn[1].n4 98.981
R23117 XThR.Tn[1].n7 XThR.Tn[1].n5 98.981
R23118 XThR.Tn[1].n9 XThR.Tn[1].n8 36.2672
R23119 XThR.Tn[1].n8 XThR.Tn[1].n7 36.2672
R23120 XThR.Tn[1].n88 XThR.Tn[1].n9 32.6405
R23121 XThR.Tn[1].n1 XThR.Tn[1].t11 26.5955
R23122 XThR.Tn[1].n1 XThR.Tn[1].t10 26.5955
R23123 XThR.Tn[1].n0 XThR.Tn[1].t8 26.5955
R23124 XThR.Tn[1].n0 XThR.Tn[1].t9 26.5955
R23125 XThR.Tn[1].n3 XThR.Tn[1].t7 24.9236
R23126 XThR.Tn[1].n3 XThR.Tn[1].t4 24.9236
R23127 XThR.Tn[1].n4 XThR.Tn[1].t6 24.9236
R23128 XThR.Tn[1].n4 XThR.Tn[1].t5 24.9236
R23129 XThR.Tn[1].n5 XThR.Tn[1].t2 24.9236
R23130 XThR.Tn[1].n5 XThR.Tn[1].t1 24.9236
R23131 XThR.Tn[1].n6 XThR.Tn[1].t3 24.9236
R23132 XThR.Tn[1].n6 XThR.Tn[1].t0 24.9236
R23133 XThR.Tn[1].n89 XThR.Tn[1].n2 18.5605
R23134 XThR.Tn[1].n89 XThR.Tn[1].n88 11.5205
R23135 XThR.Tn[1].n88 XThR.Tn[1] 6.42118
R23136 XThR.Tn[1] XThR.Tn[1].n11 5.4407
R23137 XThR.Tn[1].n16 XThR.Tn[1].n15 4.5005
R23138 XThR.Tn[1].n21 XThR.Tn[1].n20 4.5005
R23139 XThR.Tn[1].n26 XThR.Tn[1].n25 4.5005
R23140 XThR.Tn[1].n31 XThR.Tn[1].n30 4.5005
R23141 XThR.Tn[1].n36 XThR.Tn[1].n35 4.5005
R23142 XThR.Tn[1].n41 XThR.Tn[1].n40 4.5005
R23143 XThR.Tn[1].n46 XThR.Tn[1].n45 4.5005
R23144 XThR.Tn[1].n51 XThR.Tn[1].n50 4.5005
R23145 XThR.Tn[1].n56 XThR.Tn[1].n55 4.5005
R23146 XThR.Tn[1].n61 XThR.Tn[1].n60 4.5005
R23147 XThR.Tn[1].n66 XThR.Tn[1].n65 4.5005
R23148 XThR.Tn[1].n71 XThR.Tn[1].n70 4.5005
R23149 XThR.Tn[1].n76 XThR.Tn[1].n75 4.5005
R23150 XThR.Tn[1].n81 XThR.Tn[1].n80 4.5005
R23151 XThR.Tn[1].n86 XThR.Tn[1].n85 4.5005
R23152 XThR.Tn[1].n87 XThR.Tn[1] 3.70586
R23153 XThR.Tn[1].n16 XThR.Tn[1] 2.52282
R23154 XThR.Tn[1].n21 XThR.Tn[1] 2.52282
R23155 XThR.Tn[1].n26 XThR.Tn[1] 2.52282
R23156 XThR.Tn[1].n31 XThR.Tn[1] 2.52282
R23157 XThR.Tn[1].n36 XThR.Tn[1] 2.52282
R23158 XThR.Tn[1].n41 XThR.Tn[1] 2.52282
R23159 XThR.Tn[1].n46 XThR.Tn[1] 2.52282
R23160 XThR.Tn[1].n51 XThR.Tn[1] 2.52282
R23161 XThR.Tn[1].n56 XThR.Tn[1] 2.52282
R23162 XThR.Tn[1].n61 XThR.Tn[1] 2.52282
R23163 XThR.Tn[1].n66 XThR.Tn[1] 2.52282
R23164 XThR.Tn[1].n71 XThR.Tn[1] 2.52282
R23165 XThR.Tn[1].n76 XThR.Tn[1] 2.52282
R23166 XThR.Tn[1].n81 XThR.Tn[1] 2.52282
R23167 XThR.Tn[1].n86 XThR.Tn[1] 2.52282
R23168 XThR.Tn[1].n84 XThR.Tn[1] 1.08677
R23169 XThR.Tn[1].n79 XThR.Tn[1] 1.08677
R23170 XThR.Tn[1].n74 XThR.Tn[1] 1.08677
R23171 XThR.Tn[1].n69 XThR.Tn[1] 1.08677
R23172 XThR.Tn[1].n64 XThR.Tn[1] 1.08677
R23173 XThR.Tn[1].n59 XThR.Tn[1] 1.08677
R23174 XThR.Tn[1].n54 XThR.Tn[1] 1.08677
R23175 XThR.Tn[1].n49 XThR.Tn[1] 1.08677
R23176 XThR.Tn[1].n44 XThR.Tn[1] 1.08677
R23177 XThR.Tn[1].n39 XThR.Tn[1] 1.08677
R23178 XThR.Tn[1].n34 XThR.Tn[1] 1.08677
R23179 XThR.Tn[1].n29 XThR.Tn[1] 1.08677
R23180 XThR.Tn[1].n24 XThR.Tn[1] 1.08677
R23181 XThR.Tn[1].n19 XThR.Tn[1] 1.08677
R23182 XThR.Tn[1].n14 XThR.Tn[1] 1.08677
R23183 XThR.Tn[1] XThR.Tn[1].n16 0.839786
R23184 XThR.Tn[1] XThR.Tn[1].n21 0.839786
R23185 XThR.Tn[1] XThR.Tn[1].n26 0.839786
R23186 XThR.Tn[1] XThR.Tn[1].n31 0.839786
R23187 XThR.Tn[1] XThR.Tn[1].n36 0.839786
R23188 XThR.Tn[1] XThR.Tn[1].n41 0.839786
R23189 XThR.Tn[1] XThR.Tn[1].n46 0.839786
R23190 XThR.Tn[1] XThR.Tn[1].n51 0.839786
R23191 XThR.Tn[1] XThR.Tn[1].n56 0.839786
R23192 XThR.Tn[1] XThR.Tn[1].n61 0.839786
R23193 XThR.Tn[1] XThR.Tn[1].n66 0.839786
R23194 XThR.Tn[1] XThR.Tn[1].n71 0.839786
R23195 XThR.Tn[1] XThR.Tn[1].n76 0.839786
R23196 XThR.Tn[1] XThR.Tn[1].n81 0.839786
R23197 XThR.Tn[1] XThR.Tn[1].n86 0.839786
R23198 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R23199 XThR.Tn[1].n11 XThR.Tn[1] 0.499542
R23200 XThR.Tn[1].n85 XThR.Tn[1] 0.063
R23201 XThR.Tn[1].n80 XThR.Tn[1] 0.063
R23202 XThR.Tn[1].n75 XThR.Tn[1] 0.063
R23203 XThR.Tn[1].n70 XThR.Tn[1] 0.063
R23204 XThR.Tn[1].n65 XThR.Tn[1] 0.063
R23205 XThR.Tn[1].n60 XThR.Tn[1] 0.063
R23206 XThR.Tn[1].n55 XThR.Tn[1] 0.063
R23207 XThR.Tn[1].n50 XThR.Tn[1] 0.063
R23208 XThR.Tn[1].n45 XThR.Tn[1] 0.063
R23209 XThR.Tn[1].n40 XThR.Tn[1] 0.063
R23210 XThR.Tn[1].n35 XThR.Tn[1] 0.063
R23211 XThR.Tn[1].n30 XThR.Tn[1] 0.063
R23212 XThR.Tn[1].n25 XThR.Tn[1] 0.063
R23213 XThR.Tn[1].n20 XThR.Tn[1] 0.063
R23214 XThR.Tn[1].n15 XThR.Tn[1] 0.063
R23215 XThR.Tn[1].n87 XThR.Tn[1] 0.0540714
R23216 XThR.Tn[1] XThR.Tn[1].n87 0.038
R23217 XThR.Tn[1].n11 XThR.Tn[1] 0.0143889
R23218 XThR.Tn[1].n85 XThR.Tn[1].n84 0.00771154
R23219 XThR.Tn[1].n80 XThR.Tn[1].n79 0.00771154
R23220 XThR.Tn[1].n75 XThR.Tn[1].n74 0.00771154
R23221 XThR.Tn[1].n70 XThR.Tn[1].n69 0.00771154
R23222 XThR.Tn[1].n65 XThR.Tn[1].n64 0.00771154
R23223 XThR.Tn[1].n60 XThR.Tn[1].n59 0.00771154
R23224 XThR.Tn[1].n55 XThR.Tn[1].n54 0.00771154
R23225 XThR.Tn[1].n50 XThR.Tn[1].n49 0.00771154
R23226 XThR.Tn[1].n45 XThR.Tn[1].n44 0.00771154
R23227 XThR.Tn[1].n40 XThR.Tn[1].n39 0.00771154
R23228 XThR.Tn[1].n35 XThR.Tn[1].n34 0.00771154
R23229 XThR.Tn[1].n30 XThR.Tn[1].n29 0.00771154
R23230 XThR.Tn[1].n25 XThR.Tn[1].n24 0.00771154
R23231 XThR.Tn[1].n20 XThR.Tn[1].n19 0.00771154
R23232 XThR.Tn[1].n15 XThR.Tn[1].n14 0.00771154
R23233 XThC.Tn[7].n2 XThC.Tn[7].n1 255.096
R23234 XThC.Tn[7].n55 XThC.Tn[7].n53 236.589
R23235 XThC.Tn[7].n2 XThC.Tn[7].n0 201.845
R23236 XThC.Tn[7].n55 XThC.Tn[7].n54 200.321
R23237 XThC.Tn[7].n5 XThC.Tn[7].n3 161.406
R23238 XThC.Tn[7].n8 XThC.Tn[7].n6 161.406
R23239 XThC.Tn[7].n11 XThC.Tn[7].n9 161.406
R23240 XThC.Tn[7].n14 XThC.Tn[7].n12 161.406
R23241 XThC.Tn[7].n17 XThC.Tn[7].n15 161.406
R23242 XThC.Tn[7].n20 XThC.Tn[7].n18 161.406
R23243 XThC.Tn[7].n23 XThC.Tn[7].n21 161.406
R23244 XThC.Tn[7].n26 XThC.Tn[7].n24 161.406
R23245 XThC.Tn[7].n29 XThC.Tn[7].n27 161.406
R23246 XThC.Tn[7].n32 XThC.Tn[7].n30 161.406
R23247 XThC.Tn[7].n35 XThC.Tn[7].n33 161.406
R23248 XThC.Tn[7].n38 XThC.Tn[7].n36 161.406
R23249 XThC.Tn[7].n41 XThC.Tn[7].n39 161.406
R23250 XThC.Tn[7].n44 XThC.Tn[7].n42 161.406
R23251 XThC.Tn[7].n47 XThC.Tn[7].n45 161.406
R23252 XThC.Tn[7].n50 XThC.Tn[7].n48 161.406
R23253 XThC.Tn[7].n3 XThC.Tn[7].t11 161.202
R23254 XThC.Tn[7].n6 XThC.Tn[7].t30 161.202
R23255 XThC.Tn[7].n9 XThC.Tn[7].t34 161.202
R23256 XThC.Tn[7].n12 XThC.Tn[7].t35 161.202
R23257 XThC.Tn[7].n15 XThC.Tn[7].t22 161.202
R23258 XThC.Tn[7].n18 XThC.Tn[7].t23 161.202
R23259 XThC.Tn[7].n21 XThC.Tn[7].t39 161.202
R23260 XThC.Tn[7].n24 XThC.Tn[7].t14 161.202
R23261 XThC.Tn[7].n27 XThC.Tn[7].t16 161.202
R23262 XThC.Tn[7].n30 XThC.Tn[7].t36 161.202
R23263 XThC.Tn[7].n33 XThC.Tn[7].t38 161.202
R23264 XThC.Tn[7].n36 XThC.Tn[7].t17 161.202
R23265 XThC.Tn[7].n39 XThC.Tn[7].t26 161.202
R23266 XThC.Tn[7].n42 XThC.Tn[7].t28 161.202
R23267 XThC.Tn[7].n45 XThC.Tn[7].t9 161.202
R23268 XThC.Tn[7].n48 XThC.Tn[7].t19 161.202
R23269 XThC.Tn[7].n3 XThC.Tn[7].t8 145.137
R23270 XThC.Tn[7].n6 XThC.Tn[7].t25 145.137
R23271 XThC.Tn[7].n9 XThC.Tn[7].t27 145.137
R23272 XThC.Tn[7].n12 XThC.Tn[7].t29 145.137
R23273 XThC.Tn[7].n15 XThC.Tn[7].t18 145.137
R23274 XThC.Tn[7].n18 XThC.Tn[7].t20 145.137
R23275 XThC.Tn[7].n21 XThC.Tn[7].t33 145.137
R23276 XThC.Tn[7].n24 XThC.Tn[7].t10 145.137
R23277 XThC.Tn[7].n27 XThC.Tn[7].t12 145.137
R23278 XThC.Tn[7].n30 XThC.Tn[7].t31 145.137
R23279 XThC.Tn[7].n33 XThC.Tn[7].t32 145.137
R23280 XThC.Tn[7].n36 XThC.Tn[7].t13 145.137
R23281 XThC.Tn[7].n39 XThC.Tn[7].t21 145.137
R23282 XThC.Tn[7].n42 XThC.Tn[7].t24 145.137
R23283 XThC.Tn[7].n45 XThC.Tn[7].t37 145.137
R23284 XThC.Tn[7].n48 XThC.Tn[7].t15 145.137
R23285 XThC.Tn[7].n0 XThC.Tn[7].t4 26.5955
R23286 XThC.Tn[7].n0 XThC.Tn[7].t7 26.5955
R23287 XThC.Tn[7].n1 XThC.Tn[7].t6 26.5955
R23288 XThC.Tn[7].n1 XThC.Tn[7].t5 26.5955
R23289 XThC.Tn[7] XThC.Tn[7].n2 26.5002
R23290 XThC.Tn[7].n53 XThC.Tn[7].t2 24.9236
R23291 XThC.Tn[7].n53 XThC.Tn[7].t1 24.9236
R23292 XThC.Tn[7].n54 XThC.Tn[7].t0 24.9236
R23293 XThC.Tn[7].n54 XThC.Tn[7].t3 24.9236
R23294 XThC.Tn[7].n56 XThC.Tn[7].n55 12.0894
R23295 XThC.Tn[7].n56 XThC.Tn[7] 9.64206
R23296 XThC.Tn[7].n52 XThC.Tn[7] 8.14595
R23297 XThC.Tn[7].n52 XThC.Tn[7].n51 3.36239
R23298 XThC.Tn[7] XThC.Tn[7].n52 3.15894
R23299 XThC.Tn[7].n51 XThC.Tn[7] 2.07622
R23300 XThC.Tn[7] XThC.Tn[7].n56 1.66284
R23301 XThC.Tn[7].n8 XThC.Tn[7] 0.931056
R23302 XThC.Tn[7].n11 XThC.Tn[7] 0.931056
R23303 XThC.Tn[7].n14 XThC.Tn[7] 0.931056
R23304 XThC.Tn[7].n17 XThC.Tn[7] 0.931056
R23305 XThC.Tn[7].n20 XThC.Tn[7] 0.931056
R23306 XThC.Tn[7].n23 XThC.Tn[7] 0.931056
R23307 XThC.Tn[7].n26 XThC.Tn[7] 0.931056
R23308 XThC.Tn[7].n29 XThC.Tn[7] 0.931056
R23309 XThC.Tn[7].n32 XThC.Tn[7] 0.931056
R23310 XThC.Tn[7].n35 XThC.Tn[7] 0.931056
R23311 XThC.Tn[7].n38 XThC.Tn[7] 0.931056
R23312 XThC.Tn[7].n41 XThC.Tn[7] 0.931056
R23313 XThC.Tn[7].n44 XThC.Tn[7] 0.931056
R23314 XThC.Tn[7].n47 XThC.Tn[7] 0.931056
R23315 XThC.Tn[7].n50 XThC.Tn[7] 0.931056
R23316 XThC.Tn[7] XThC.Tn[7].n5 0.396333
R23317 XThC.Tn[7] XThC.Tn[7].n8 0.396333
R23318 XThC.Tn[7] XThC.Tn[7].n11 0.396333
R23319 XThC.Tn[7] XThC.Tn[7].n14 0.396333
R23320 XThC.Tn[7] XThC.Tn[7].n17 0.396333
R23321 XThC.Tn[7] XThC.Tn[7].n20 0.396333
R23322 XThC.Tn[7] XThC.Tn[7].n23 0.396333
R23323 XThC.Tn[7] XThC.Tn[7].n26 0.396333
R23324 XThC.Tn[7] XThC.Tn[7].n29 0.396333
R23325 XThC.Tn[7] XThC.Tn[7].n32 0.396333
R23326 XThC.Tn[7] XThC.Tn[7].n35 0.396333
R23327 XThC.Tn[7] XThC.Tn[7].n38 0.396333
R23328 XThC.Tn[7] XThC.Tn[7].n41 0.396333
R23329 XThC.Tn[7] XThC.Tn[7].n44 0.396333
R23330 XThC.Tn[7] XThC.Tn[7].n47 0.396333
R23331 XThC.Tn[7] XThC.Tn[7].n50 0.396333
R23332 XThC.Tn[7].n4 XThC.Tn[7] 0.104667
R23333 XThC.Tn[7].n7 XThC.Tn[7] 0.104667
R23334 XThC.Tn[7].n10 XThC.Tn[7] 0.104667
R23335 XThC.Tn[7].n13 XThC.Tn[7] 0.104667
R23336 XThC.Tn[7].n16 XThC.Tn[7] 0.104667
R23337 XThC.Tn[7].n19 XThC.Tn[7] 0.104667
R23338 XThC.Tn[7].n22 XThC.Tn[7] 0.104667
R23339 XThC.Tn[7].n25 XThC.Tn[7] 0.104667
R23340 XThC.Tn[7].n28 XThC.Tn[7] 0.104667
R23341 XThC.Tn[7].n31 XThC.Tn[7] 0.104667
R23342 XThC.Tn[7].n34 XThC.Tn[7] 0.104667
R23343 XThC.Tn[7].n37 XThC.Tn[7] 0.104667
R23344 XThC.Tn[7].n40 XThC.Tn[7] 0.104667
R23345 XThC.Tn[7].n43 XThC.Tn[7] 0.104667
R23346 XThC.Tn[7].n46 XThC.Tn[7] 0.104667
R23347 XThC.Tn[7].n49 XThC.Tn[7] 0.104667
R23348 XThC.Tn[7].n4 XThC.Tn[7] 0.0309878
R23349 XThC.Tn[7].n7 XThC.Tn[7] 0.0309878
R23350 XThC.Tn[7].n10 XThC.Tn[7] 0.0309878
R23351 XThC.Tn[7].n13 XThC.Tn[7] 0.0309878
R23352 XThC.Tn[7].n16 XThC.Tn[7] 0.0309878
R23353 XThC.Tn[7].n19 XThC.Tn[7] 0.0309878
R23354 XThC.Tn[7].n22 XThC.Tn[7] 0.0309878
R23355 XThC.Tn[7].n25 XThC.Tn[7] 0.0309878
R23356 XThC.Tn[7].n28 XThC.Tn[7] 0.0309878
R23357 XThC.Tn[7].n31 XThC.Tn[7] 0.0309878
R23358 XThC.Tn[7].n34 XThC.Tn[7] 0.0309878
R23359 XThC.Tn[7].n37 XThC.Tn[7] 0.0309878
R23360 XThC.Tn[7].n40 XThC.Tn[7] 0.0309878
R23361 XThC.Tn[7].n43 XThC.Tn[7] 0.0309878
R23362 XThC.Tn[7].n46 XThC.Tn[7] 0.0309878
R23363 XThC.Tn[7].n49 XThC.Tn[7] 0.0309878
R23364 XThC.Tn[7].n5 XThC.Tn[7].n4 0.027939
R23365 XThC.Tn[7].n8 XThC.Tn[7].n7 0.027939
R23366 XThC.Tn[7].n11 XThC.Tn[7].n10 0.027939
R23367 XThC.Tn[7].n14 XThC.Tn[7].n13 0.027939
R23368 XThC.Tn[7].n17 XThC.Tn[7].n16 0.027939
R23369 XThC.Tn[7].n20 XThC.Tn[7].n19 0.027939
R23370 XThC.Tn[7].n23 XThC.Tn[7].n22 0.027939
R23371 XThC.Tn[7].n26 XThC.Tn[7].n25 0.027939
R23372 XThC.Tn[7].n29 XThC.Tn[7].n28 0.027939
R23373 XThC.Tn[7].n32 XThC.Tn[7].n31 0.027939
R23374 XThC.Tn[7].n35 XThC.Tn[7].n34 0.027939
R23375 XThC.Tn[7].n38 XThC.Tn[7].n37 0.027939
R23376 XThC.Tn[7].n41 XThC.Tn[7].n40 0.027939
R23377 XThC.Tn[7].n44 XThC.Tn[7].n43 0.027939
R23378 XThC.Tn[7].n47 XThC.Tn[7].n46 0.027939
R23379 XThC.Tn[7].n50 XThC.Tn[7].n49 0.027939
R23380 XThC.Tn[7].n51 XThC.Tn[7] 0.00240908
R23381 XThR.Tn[4].n2 XThR.Tn[4].n1 332.334
R23382 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R23383 XThR.Tn[4] XThR.Tn[4].n82 161.363
R23384 XThR.Tn[4] XThR.Tn[4].n77 161.363
R23385 XThR.Tn[4] XThR.Tn[4].n72 161.363
R23386 XThR.Tn[4] XThR.Tn[4].n67 161.363
R23387 XThR.Tn[4] XThR.Tn[4].n62 161.363
R23388 XThR.Tn[4] XThR.Tn[4].n57 161.363
R23389 XThR.Tn[4] XThR.Tn[4].n52 161.363
R23390 XThR.Tn[4] XThR.Tn[4].n47 161.363
R23391 XThR.Tn[4] XThR.Tn[4].n42 161.363
R23392 XThR.Tn[4] XThR.Tn[4].n37 161.363
R23393 XThR.Tn[4] XThR.Tn[4].n32 161.363
R23394 XThR.Tn[4] XThR.Tn[4].n27 161.363
R23395 XThR.Tn[4] XThR.Tn[4].n22 161.363
R23396 XThR.Tn[4] XThR.Tn[4].n17 161.363
R23397 XThR.Tn[4] XThR.Tn[4].n12 161.363
R23398 XThR.Tn[4] XThR.Tn[4].n10 161.363
R23399 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R23400 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R23401 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R23402 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R23403 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R23404 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R23405 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R23406 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R23407 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R23408 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R23409 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R23410 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R23411 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R23412 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R23413 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R23414 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R23415 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R23416 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R23417 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R23418 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R23419 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R23420 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R23421 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R23422 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R23423 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R23424 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R23425 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R23426 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R23427 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R23428 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R23429 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R23430 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R23431 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R23432 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R23433 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R23434 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R23435 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R23436 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R23437 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R23438 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R23439 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R23440 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R23441 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R23442 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R23443 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R23444 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R23445 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R23446 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R23447 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R23448 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R23449 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R23450 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R23451 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R23452 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R23453 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R23454 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R23455 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R23456 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R23457 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R23458 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R23459 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R23460 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R23461 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R23462 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R23463 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R23464 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R23465 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R23466 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R23467 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R23468 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R23469 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R23470 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R23471 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R23472 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R23473 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R23474 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R23475 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R23476 XThR.Tn[4].n5 XThR.Tn[4].n3 135.249
R23477 XThR.Tn[4].n5 XThR.Tn[4].n4 98.982
R23478 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R23479 XThR.Tn[4].n9 XThR.Tn[4].n8 98.982
R23480 XThR.Tn[4].n7 XThR.Tn[4].n5 36.2672
R23481 XThR.Tn[4].n9 XThR.Tn[4].n7 36.2672
R23482 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R23483 XThR.Tn[4].n0 XThR.Tn[4].t1 26.5955
R23484 XThR.Tn[4].n0 XThR.Tn[4].t2 26.5955
R23485 XThR.Tn[4].n1 XThR.Tn[4].t0 26.5955
R23486 XThR.Tn[4].n1 XThR.Tn[4].t3 26.5955
R23487 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R23488 XThR.Tn[4].n3 XThR.Tn[4].t9 24.9236
R23489 XThR.Tn[4].n4 XThR.Tn[4].t11 24.9236
R23490 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R23491 XThR.Tn[4].n6 XThR.Tn[4].t6 24.9236
R23492 XThR.Tn[4].n6 XThR.Tn[4].t5 24.9236
R23493 XThR.Tn[4].n8 XThR.Tn[4].t7 24.9236
R23494 XThR.Tn[4].n8 XThR.Tn[4].t4 24.9236
R23495 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R23496 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R23497 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R23498 XThR.Tn[4] XThR.Tn[4].n11 5.4407
R23499 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R23500 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R23501 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R23502 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R23503 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R23504 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R23505 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R23506 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R23507 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R23508 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R23509 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R23510 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R23511 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R23512 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R23513 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R23514 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R23515 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R23516 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R23517 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R23518 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R23519 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R23520 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R23521 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R23522 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R23523 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R23524 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R23525 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R23526 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R23527 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R23528 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R23529 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R23530 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R23531 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R23532 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R23533 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R23534 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R23535 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R23536 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R23537 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R23538 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R23539 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R23540 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R23541 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R23542 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R23543 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R23544 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R23545 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R23546 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R23547 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R23548 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R23549 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R23550 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R23551 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R23552 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R23553 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R23554 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R23555 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R23556 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R23557 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R23558 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R23559 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R23560 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R23561 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R23562 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R23563 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R23564 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R23565 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R23566 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R23567 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R23568 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R23569 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R23570 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R23571 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R23572 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R23573 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R23574 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R23575 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R23576 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R23577 XThR.Tn[4] XThR.Tn[4].n87 0.038
R23578 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R23579 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R23580 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R23581 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R23582 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R23583 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R23584 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R23585 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R23586 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R23587 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R23588 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R23589 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R23590 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R23591 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R23592 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R23593 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R23594 XThR.Tn[11].n87 XThR.Tn[11].n86 256.103
R23595 XThR.Tn[11].n2 XThR.Tn[11].n0 243.68
R23596 XThR.Tn[11].n5 XThR.Tn[11].n3 241.847
R23597 XThR.Tn[11].n2 XThR.Tn[11].n1 205.28
R23598 XThR.Tn[11].n87 XThR.Tn[11].n85 202.094
R23599 XThR.Tn[11].n5 XThR.Tn[11].n4 185
R23600 XThR.Tn[11] XThR.Tn[11].n78 161.363
R23601 XThR.Tn[11] XThR.Tn[11].n73 161.363
R23602 XThR.Tn[11] XThR.Tn[11].n68 161.363
R23603 XThR.Tn[11] XThR.Tn[11].n63 161.363
R23604 XThR.Tn[11] XThR.Tn[11].n58 161.363
R23605 XThR.Tn[11] XThR.Tn[11].n53 161.363
R23606 XThR.Tn[11] XThR.Tn[11].n48 161.363
R23607 XThR.Tn[11] XThR.Tn[11].n43 161.363
R23608 XThR.Tn[11] XThR.Tn[11].n38 161.363
R23609 XThR.Tn[11] XThR.Tn[11].n33 161.363
R23610 XThR.Tn[11] XThR.Tn[11].n28 161.363
R23611 XThR.Tn[11] XThR.Tn[11].n23 161.363
R23612 XThR.Tn[11] XThR.Tn[11].n18 161.363
R23613 XThR.Tn[11] XThR.Tn[11].n13 161.363
R23614 XThR.Tn[11] XThR.Tn[11].n8 161.363
R23615 XThR.Tn[11] XThR.Tn[11].n6 161.363
R23616 XThR.Tn[11].n80 XThR.Tn[11].n79 161.3
R23617 XThR.Tn[11].n75 XThR.Tn[11].n74 161.3
R23618 XThR.Tn[11].n70 XThR.Tn[11].n69 161.3
R23619 XThR.Tn[11].n65 XThR.Tn[11].n64 161.3
R23620 XThR.Tn[11].n60 XThR.Tn[11].n59 161.3
R23621 XThR.Tn[11].n55 XThR.Tn[11].n54 161.3
R23622 XThR.Tn[11].n50 XThR.Tn[11].n49 161.3
R23623 XThR.Tn[11].n45 XThR.Tn[11].n44 161.3
R23624 XThR.Tn[11].n40 XThR.Tn[11].n39 161.3
R23625 XThR.Tn[11].n35 XThR.Tn[11].n34 161.3
R23626 XThR.Tn[11].n30 XThR.Tn[11].n29 161.3
R23627 XThR.Tn[11].n25 XThR.Tn[11].n24 161.3
R23628 XThR.Tn[11].n20 XThR.Tn[11].n19 161.3
R23629 XThR.Tn[11].n15 XThR.Tn[11].n14 161.3
R23630 XThR.Tn[11].n10 XThR.Tn[11].n9 161.3
R23631 XThR.Tn[11].n78 XThR.Tn[11].t40 161.106
R23632 XThR.Tn[11].n73 XThR.Tn[11].t46 161.106
R23633 XThR.Tn[11].n68 XThR.Tn[11].t24 161.106
R23634 XThR.Tn[11].n63 XThR.Tn[11].t73 161.106
R23635 XThR.Tn[11].n58 XThR.Tn[11].t39 161.106
R23636 XThR.Tn[11].n53 XThR.Tn[11].t63 161.106
R23637 XThR.Tn[11].n48 XThR.Tn[11].t43 161.106
R23638 XThR.Tn[11].n43 XThR.Tn[11].t22 161.106
R23639 XThR.Tn[11].n38 XThR.Tn[11].t71 161.106
R23640 XThR.Tn[11].n33 XThR.Tn[11].t14 161.106
R23641 XThR.Tn[11].n28 XThR.Tn[11].t62 161.106
R23642 XThR.Tn[11].n23 XThR.Tn[11].t23 161.106
R23643 XThR.Tn[11].n18 XThR.Tn[11].t60 161.106
R23644 XThR.Tn[11].n13 XThR.Tn[11].t41 161.106
R23645 XThR.Tn[11].n8 XThR.Tn[11].t67 161.106
R23646 XThR.Tn[11].n6 XThR.Tn[11].t48 161.106
R23647 XThR.Tn[11].n79 XThR.Tn[11].t31 159.978
R23648 XThR.Tn[11].n74 XThR.Tn[11].t38 159.978
R23649 XThR.Tn[11].n69 XThR.Tn[11].t20 159.978
R23650 XThR.Tn[11].n64 XThR.Tn[11].t66 159.978
R23651 XThR.Tn[11].n59 XThR.Tn[11].t29 159.978
R23652 XThR.Tn[11].n54 XThR.Tn[11].t57 159.978
R23653 XThR.Tn[11].n49 XThR.Tn[11].t37 159.978
R23654 XThR.Tn[11].n44 XThR.Tn[11].t17 159.978
R23655 XThR.Tn[11].n39 XThR.Tn[11].t64 159.978
R23656 XThR.Tn[11].n34 XThR.Tn[11].t72 159.978
R23657 XThR.Tn[11].n29 XThR.Tn[11].t55 159.978
R23658 XThR.Tn[11].n24 XThR.Tn[11].t19 159.978
R23659 XThR.Tn[11].n19 XThR.Tn[11].t54 159.978
R23660 XThR.Tn[11].n14 XThR.Tn[11].t36 159.978
R23661 XThR.Tn[11].n9 XThR.Tn[11].t58 159.978
R23662 XThR.Tn[11].n78 XThR.Tn[11].t26 145.038
R23663 XThR.Tn[11].n73 XThR.Tn[11].t53 145.038
R23664 XThR.Tn[11].n68 XThR.Tn[11].t34 145.038
R23665 XThR.Tn[11].n63 XThR.Tn[11].t15 145.038
R23666 XThR.Tn[11].n58 XThR.Tn[11].t47 145.038
R23667 XThR.Tn[11].n53 XThR.Tn[11].t25 145.038
R23668 XThR.Tn[11].n48 XThR.Tn[11].t35 145.038
R23669 XThR.Tn[11].n43 XThR.Tn[11].t16 145.038
R23670 XThR.Tn[11].n38 XThR.Tn[11].t13 145.038
R23671 XThR.Tn[11].n33 XThR.Tn[11].t44 145.038
R23672 XThR.Tn[11].n28 XThR.Tn[11].t70 145.038
R23673 XThR.Tn[11].n23 XThR.Tn[11].t33 145.038
R23674 XThR.Tn[11].n18 XThR.Tn[11].t68 145.038
R23675 XThR.Tn[11].n13 XThR.Tn[11].t49 145.038
R23676 XThR.Tn[11].n8 XThR.Tn[11].t12 145.038
R23677 XThR.Tn[11].n6 XThR.Tn[11].t56 145.038
R23678 XThR.Tn[11].n79 XThR.Tn[11].t45 143.911
R23679 XThR.Tn[11].n74 XThR.Tn[11].t69 143.911
R23680 XThR.Tn[11].n69 XThR.Tn[11].t51 143.911
R23681 XThR.Tn[11].n64 XThR.Tn[11].t30 143.911
R23682 XThR.Tn[11].n59 XThR.Tn[11].t61 143.911
R23683 XThR.Tn[11].n54 XThR.Tn[11].t42 143.911
R23684 XThR.Tn[11].n49 XThR.Tn[11].t52 143.911
R23685 XThR.Tn[11].n44 XThR.Tn[11].t32 143.911
R23686 XThR.Tn[11].n39 XThR.Tn[11].t28 143.911
R23687 XThR.Tn[11].n34 XThR.Tn[11].t59 143.911
R23688 XThR.Tn[11].n29 XThR.Tn[11].t21 143.911
R23689 XThR.Tn[11].n24 XThR.Tn[11].t50 143.911
R23690 XThR.Tn[11].n19 XThR.Tn[11].t18 143.911
R23691 XThR.Tn[11].n14 XThR.Tn[11].t65 143.911
R23692 XThR.Tn[11].n9 XThR.Tn[11].t27 143.911
R23693 XThR.Tn[11] XThR.Tn[11].n2 35.7652
R23694 XThR.Tn[11].n85 XThR.Tn[11].t0 26.5955
R23695 XThR.Tn[11].n85 XThR.Tn[11].t2 26.5955
R23696 XThR.Tn[11].n0 XThR.Tn[11].t8 26.5955
R23697 XThR.Tn[11].n0 XThR.Tn[11].t10 26.5955
R23698 XThR.Tn[11].n1 XThR.Tn[11].t9 26.5955
R23699 XThR.Tn[11].n1 XThR.Tn[11].t11 26.5955
R23700 XThR.Tn[11].n86 XThR.Tn[11].t1 26.5955
R23701 XThR.Tn[11].n86 XThR.Tn[11].t3 26.5955
R23702 XThR.Tn[11].n4 XThR.Tn[11].t6 24.9236
R23703 XThR.Tn[11].n4 XThR.Tn[11].t4 24.9236
R23704 XThR.Tn[11].n3 XThR.Tn[11].t7 24.9236
R23705 XThR.Tn[11].n3 XThR.Tn[11].t5 24.9236
R23706 XThR.Tn[11] XThR.Tn[11].n5 22.9615
R23707 XThR.Tn[11].n88 XThR.Tn[11].n87 13.5534
R23708 XThR.Tn[11].n84 XThR.Tn[11] 8.41462
R23709 XThR.Tn[11] XThR.Tn[11].n7 5.4407
R23710 XThR.Tn[11].n12 XThR.Tn[11].n11 4.5005
R23711 XThR.Tn[11].n17 XThR.Tn[11].n16 4.5005
R23712 XThR.Tn[11].n22 XThR.Tn[11].n21 4.5005
R23713 XThR.Tn[11].n27 XThR.Tn[11].n26 4.5005
R23714 XThR.Tn[11].n32 XThR.Tn[11].n31 4.5005
R23715 XThR.Tn[11].n37 XThR.Tn[11].n36 4.5005
R23716 XThR.Tn[11].n42 XThR.Tn[11].n41 4.5005
R23717 XThR.Tn[11].n47 XThR.Tn[11].n46 4.5005
R23718 XThR.Tn[11].n52 XThR.Tn[11].n51 4.5005
R23719 XThR.Tn[11].n57 XThR.Tn[11].n56 4.5005
R23720 XThR.Tn[11].n62 XThR.Tn[11].n61 4.5005
R23721 XThR.Tn[11].n67 XThR.Tn[11].n66 4.5005
R23722 XThR.Tn[11].n72 XThR.Tn[11].n71 4.5005
R23723 XThR.Tn[11].n77 XThR.Tn[11].n76 4.5005
R23724 XThR.Tn[11].n82 XThR.Tn[11].n81 4.5005
R23725 XThR.Tn[11].n83 XThR.Tn[11] 3.70586
R23726 XThR.Tn[11].n88 XThR.Tn[11].n84 2.99115
R23727 XThR.Tn[11].n88 XThR.Tn[11] 2.87153
R23728 XThR.Tn[11].n12 XThR.Tn[11] 2.52282
R23729 XThR.Tn[11].n17 XThR.Tn[11] 2.52282
R23730 XThR.Tn[11].n22 XThR.Tn[11] 2.52282
R23731 XThR.Tn[11].n27 XThR.Tn[11] 2.52282
R23732 XThR.Tn[11].n32 XThR.Tn[11] 2.52282
R23733 XThR.Tn[11].n37 XThR.Tn[11] 2.52282
R23734 XThR.Tn[11].n42 XThR.Tn[11] 2.52282
R23735 XThR.Tn[11].n47 XThR.Tn[11] 2.52282
R23736 XThR.Tn[11].n52 XThR.Tn[11] 2.52282
R23737 XThR.Tn[11].n57 XThR.Tn[11] 2.52282
R23738 XThR.Tn[11].n62 XThR.Tn[11] 2.52282
R23739 XThR.Tn[11].n67 XThR.Tn[11] 2.52282
R23740 XThR.Tn[11].n72 XThR.Tn[11] 2.52282
R23741 XThR.Tn[11].n77 XThR.Tn[11] 2.52282
R23742 XThR.Tn[11].n82 XThR.Tn[11] 2.52282
R23743 XThR.Tn[11].n84 XThR.Tn[11] 2.2734
R23744 XThR.Tn[11] XThR.Tn[11].n88 1.50638
R23745 XThR.Tn[11].n80 XThR.Tn[11] 1.08677
R23746 XThR.Tn[11].n75 XThR.Tn[11] 1.08677
R23747 XThR.Tn[11].n70 XThR.Tn[11] 1.08677
R23748 XThR.Tn[11].n65 XThR.Tn[11] 1.08677
R23749 XThR.Tn[11].n60 XThR.Tn[11] 1.08677
R23750 XThR.Tn[11].n55 XThR.Tn[11] 1.08677
R23751 XThR.Tn[11].n50 XThR.Tn[11] 1.08677
R23752 XThR.Tn[11].n45 XThR.Tn[11] 1.08677
R23753 XThR.Tn[11].n40 XThR.Tn[11] 1.08677
R23754 XThR.Tn[11].n35 XThR.Tn[11] 1.08677
R23755 XThR.Tn[11].n30 XThR.Tn[11] 1.08677
R23756 XThR.Tn[11].n25 XThR.Tn[11] 1.08677
R23757 XThR.Tn[11].n20 XThR.Tn[11] 1.08677
R23758 XThR.Tn[11].n15 XThR.Tn[11] 1.08677
R23759 XThR.Tn[11].n10 XThR.Tn[11] 1.08677
R23760 XThR.Tn[11] XThR.Tn[11].n12 0.839786
R23761 XThR.Tn[11] XThR.Tn[11].n17 0.839786
R23762 XThR.Tn[11] XThR.Tn[11].n22 0.839786
R23763 XThR.Tn[11] XThR.Tn[11].n27 0.839786
R23764 XThR.Tn[11] XThR.Tn[11].n32 0.839786
R23765 XThR.Tn[11] XThR.Tn[11].n37 0.839786
R23766 XThR.Tn[11] XThR.Tn[11].n42 0.839786
R23767 XThR.Tn[11] XThR.Tn[11].n47 0.839786
R23768 XThR.Tn[11] XThR.Tn[11].n52 0.839786
R23769 XThR.Tn[11] XThR.Tn[11].n57 0.839786
R23770 XThR.Tn[11] XThR.Tn[11].n62 0.839786
R23771 XThR.Tn[11] XThR.Tn[11].n67 0.839786
R23772 XThR.Tn[11] XThR.Tn[11].n72 0.839786
R23773 XThR.Tn[11] XThR.Tn[11].n77 0.839786
R23774 XThR.Tn[11] XThR.Tn[11].n82 0.839786
R23775 XThR.Tn[11].n7 XThR.Tn[11] 0.499542
R23776 XThR.Tn[11].n81 XThR.Tn[11] 0.063
R23777 XThR.Tn[11].n76 XThR.Tn[11] 0.063
R23778 XThR.Tn[11].n71 XThR.Tn[11] 0.063
R23779 XThR.Tn[11].n66 XThR.Tn[11] 0.063
R23780 XThR.Tn[11].n61 XThR.Tn[11] 0.063
R23781 XThR.Tn[11].n56 XThR.Tn[11] 0.063
R23782 XThR.Tn[11].n51 XThR.Tn[11] 0.063
R23783 XThR.Tn[11].n46 XThR.Tn[11] 0.063
R23784 XThR.Tn[11].n41 XThR.Tn[11] 0.063
R23785 XThR.Tn[11].n36 XThR.Tn[11] 0.063
R23786 XThR.Tn[11].n31 XThR.Tn[11] 0.063
R23787 XThR.Tn[11].n26 XThR.Tn[11] 0.063
R23788 XThR.Tn[11].n21 XThR.Tn[11] 0.063
R23789 XThR.Tn[11].n16 XThR.Tn[11] 0.063
R23790 XThR.Tn[11].n11 XThR.Tn[11] 0.063
R23791 XThR.Tn[11].n83 XThR.Tn[11] 0.0540714
R23792 XThR.Tn[11] XThR.Tn[11].n83 0.038
R23793 XThR.Tn[11].n7 XThR.Tn[11] 0.0143889
R23794 XThR.Tn[11].n81 XThR.Tn[11].n80 0.00771154
R23795 XThR.Tn[11].n76 XThR.Tn[11].n75 0.00771154
R23796 XThR.Tn[11].n71 XThR.Tn[11].n70 0.00771154
R23797 XThR.Tn[11].n66 XThR.Tn[11].n65 0.00771154
R23798 XThR.Tn[11].n61 XThR.Tn[11].n60 0.00771154
R23799 XThR.Tn[11].n56 XThR.Tn[11].n55 0.00771154
R23800 XThR.Tn[11].n51 XThR.Tn[11].n50 0.00771154
R23801 XThR.Tn[11].n46 XThR.Tn[11].n45 0.00771154
R23802 XThR.Tn[11].n41 XThR.Tn[11].n40 0.00771154
R23803 XThR.Tn[11].n36 XThR.Tn[11].n35 0.00771154
R23804 XThR.Tn[11].n31 XThR.Tn[11].n30 0.00771154
R23805 XThR.Tn[11].n26 XThR.Tn[11].n25 0.00771154
R23806 XThR.Tn[11].n21 XThR.Tn[11].n20 0.00771154
R23807 XThR.Tn[11].n16 XThR.Tn[11].n15 0.00771154
R23808 XThR.Tn[11].n11 XThR.Tn[11].n10 0.00771154
R23809 XThR.Tn[7].n5 XThR.Tn[7].n3 244.069
R23810 XThR.Tn[7].n2 XThR.Tn[7].n1 236.589
R23811 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23812 XThR.Tn[7].n2 XThR.Tn[7].n0 200.321
R23813 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23814 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23815 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23816 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23817 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23818 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23819 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23820 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23821 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23822 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23823 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23824 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23825 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23826 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23827 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23828 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23829 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23830 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23831 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23832 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23833 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23834 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23835 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23836 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23837 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23838 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23839 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23840 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23841 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23842 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23843 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23844 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23845 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23846 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23847 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23848 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23849 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23850 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23851 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23852 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23853 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23854 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23855 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23856 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23857 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23858 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23859 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23860 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23861 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23862 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23863 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23864 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23865 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23866 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23867 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23868 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23869 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23870 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23871 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23872 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23873 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23874 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23875 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23876 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23877 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23878 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23879 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23880 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23881 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23882 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23883 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23884 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23885 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23886 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23887 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23888 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23889 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23890 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23891 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23892 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23893 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23894 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23895 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23896 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23897 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23898 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23899 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23900 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23901 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23902 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23903 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23904 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23905 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23906 XThR.Tn[7].n4 XThR.Tn[7].t5 26.5955
R23907 XThR.Tn[7].n4 XThR.Tn[7].t4 26.5955
R23908 XThR.Tn[7].n3 XThR.Tn[7].t6 26.5955
R23909 XThR.Tn[7].n3 XThR.Tn[7].t7 26.5955
R23910 XThR.Tn[7].n0 XThR.Tn[7].t2 24.9236
R23911 XThR.Tn[7].n0 XThR.Tn[7].t1 24.9236
R23912 XThR.Tn[7].n1 XThR.Tn[7].t3 24.9236
R23913 XThR.Tn[7].n1 XThR.Tn[7].t0 24.9236
R23914 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23915 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23916 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23917 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23918 XThR.Tn[7] XThR.Tn[7].n8 5.4407
R23919 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23920 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23921 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23922 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23923 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23924 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23925 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23926 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23927 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23928 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23929 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23930 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23931 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23932 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23933 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23934 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23935 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23936 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23937 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23938 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23939 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23940 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23941 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23942 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23943 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23944 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23945 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23946 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23947 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23948 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23949 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23950 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23951 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23952 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23953 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23954 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23955 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23956 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23957 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23958 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23959 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23960 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23961 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23962 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23963 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23964 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23965 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23966 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23967 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23968 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23969 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23970 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23971 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23972 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23973 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23974 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23975 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23976 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23977 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23978 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23979 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23980 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23981 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23982 XThR.Tn[7].n6 XThR.Tn[7] 0.829611
R23983 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23984 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23985 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23986 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23987 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23988 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23989 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23990 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23991 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23992 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23993 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23994 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23995 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23996 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23997 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23998 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23999 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R24000 XThR.Tn[7] XThR.Tn[7].n84 0.038
R24001 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R24002 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R24003 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R24004 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R24005 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R24006 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R24007 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R24008 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R24009 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R24010 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R24011 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R24012 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R24013 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R24014 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R24015 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R24016 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R24017 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R24018 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R24019 XThR.Tn[0] XThR.Tn[0].n82 161.363
R24020 XThR.Tn[0] XThR.Tn[0].n77 161.363
R24021 XThR.Tn[0] XThR.Tn[0].n72 161.363
R24022 XThR.Tn[0] XThR.Tn[0].n67 161.363
R24023 XThR.Tn[0] XThR.Tn[0].n62 161.363
R24024 XThR.Tn[0] XThR.Tn[0].n57 161.363
R24025 XThR.Tn[0] XThR.Tn[0].n52 161.363
R24026 XThR.Tn[0] XThR.Tn[0].n47 161.363
R24027 XThR.Tn[0] XThR.Tn[0].n42 161.363
R24028 XThR.Tn[0] XThR.Tn[0].n37 161.363
R24029 XThR.Tn[0] XThR.Tn[0].n32 161.363
R24030 XThR.Tn[0] XThR.Tn[0].n27 161.363
R24031 XThR.Tn[0] XThR.Tn[0].n22 161.363
R24032 XThR.Tn[0] XThR.Tn[0].n17 161.363
R24033 XThR.Tn[0] XThR.Tn[0].n12 161.363
R24034 XThR.Tn[0] XThR.Tn[0].n10 161.363
R24035 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R24036 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R24037 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R24038 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R24039 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R24040 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R24041 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R24042 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R24043 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R24044 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R24045 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R24046 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R24047 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R24048 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R24049 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R24050 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R24051 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R24052 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R24053 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R24054 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R24055 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R24056 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R24057 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R24058 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R24059 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R24060 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R24061 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R24062 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R24063 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R24064 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R24065 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R24066 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R24067 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R24068 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R24069 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R24070 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R24071 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R24072 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R24073 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R24074 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R24075 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R24076 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R24077 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R24078 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R24079 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R24080 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R24081 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R24082 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R24083 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R24084 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R24085 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R24086 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R24087 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R24088 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R24089 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R24090 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R24091 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R24092 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R24093 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R24094 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R24095 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R24096 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R24097 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R24098 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R24099 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R24100 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R24101 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R24102 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R24103 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R24104 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R24105 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R24106 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R24107 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R24108 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R24109 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R24110 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R24111 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R24112 XThR.Tn[0].n7 XThR.Tn[0].n5 135.249
R24113 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R24114 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R24115 XThR.Tn[0].n7 XThR.Tn[0].n6 98.982
R24116 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R24117 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R24118 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R24119 XThR.Tn[0].n1 XThR.Tn[0].t4 26.5955
R24120 XThR.Tn[0].n1 XThR.Tn[0].t3 26.5955
R24121 XThR.Tn[0].n0 XThR.Tn[0].t5 26.5955
R24122 XThR.Tn[0].n0 XThR.Tn[0].t6 26.5955
R24123 XThR.Tn[0].n3 XThR.Tn[0].t8 24.9236
R24124 XThR.Tn[0].n3 XThR.Tn[0].t9 24.9236
R24125 XThR.Tn[0].n4 XThR.Tn[0].t7 24.9236
R24126 XThR.Tn[0].n4 XThR.Tn[0].t10 24.9236
R24127 XThR.Tn[0].n5 XThR.Tn[0].t11 24.9236
R24128 XThR.Tn[0].n5 XThR.Tn[0].t2 24.9236
R24129 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R24130 XThR.Tn[0].n6 XThR.Tn[0].t1 24.9236
R24131 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R24132 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R24133 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R24134 XThR.Tn[0] XThR.Tn[0].n11 5.4407
R24135 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R24136 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R24137 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R24138 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R24139 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R24140 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R24141 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R24142 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R24143 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R24144 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R24145 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R24146 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R24147 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R24148 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R24149 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R24150 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R24151 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R24152 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R24153 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R24154 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R24155 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R24156 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R24157 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R24158 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R24159 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R24160 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R24161 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R24162 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R24163 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R24164 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R24165 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R24166 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R24167 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R24168 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R24169 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R24170 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R24171 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R24172 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R24173 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R24174 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R24175 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R24176 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R24177 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R24178 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R24179 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R24180 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R24181 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R24182 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R24183 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R24184 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R24185 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R24186 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R24187 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R24188 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R24189 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R24190 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R24191 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R24192 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R24193 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R24194 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R24195 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R24196 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R24197 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R24198 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R24199 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R24200 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R24201 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R24202 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R24203 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R24204 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R24205 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R24206 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R24207 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R24208 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R24209 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R24210 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R24211 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R24212 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R24213 XThR.Tn[0] XThR.Tn[0].n87 0.038
R24214 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R24215 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R24216 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R24217 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R24218 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R24219 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R24220 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R24221 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R24222 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R24223 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R24224 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R24225 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R24226 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R24227 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R24228 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R24229 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R24230 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R24231 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R24232 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R24233 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R24234 XThR.Tn[8].n87 XThR.Tn[8].n85 202.095
R24235 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R24236 XThR.Tn[8] XThR.Tn[8].n78 161.363
R24237 XThR.Tn[8] XThR.Tn[8].n73 161.363
R24238 XThR.Tn[8] XThR.Tn[8].n68 161.363
R24239 XThR.Tn[8] XThR.Tn[8].n63 161.363
R24240 XThR.Tn[8] XThR.Tn[8].n58 161.363
R24241 XThR.Tn[8] XThR.Tn[8].n53 161.363
R24242 XThR.Tn[8] XThR.Tn[8].n48 161.363
R24243 XThR.Tn[8] XThR.Tn[8].n43 161.363
R24244 XThR.Tn[8] XThR.Tn[8].n38 161.363
R24245 XThR.Tn[8] XThR.Tn[8].n33 161.363
R24246 XThR.Tn[8] XThR.Tn[8].n28 161.363
R24247 XThR.Tn[8] XThR.Tn[8].n23 161.363
R24248 XThR.Tn[8] XThR.Tn[8].n18 161.363
R24249 XThR.Tn[8] XThR.Tn[8].n13 161.363
R24250 XThR.Tn[8] XThR.Tn[8].n8 161.363
R24251 XThR.Tn[8] XThR.Tn[8].n6 161.363
R24252 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R24253 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R24254 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R24255 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R24256 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R24257 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R24258 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R24259 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R24260 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R24261 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R24262 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R24263 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R24264 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R24265 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R24266 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R24267 XThR.Tn[8].n78 XThR.Tn[8].t23 161.106
R24268 XThR.Tn[8].n73 XThR.Tn[8].t29 161.106
R24269 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R24270 XThR.Tn[8].n63 XThR.Tn[8].t57 161.106
R24271 XThR.Tn[8].n58 XThR.Tn[8].t21 161.106
R24272 XThR.Tn[8].n53 XThR.Tn[8].t46 161.106
R24273 XThR.Tn[8].n48 XThR.Tn[8].t27 161.106
R24274 XThR.Tn[8].n43 XThR.Tn[8].t69 161.106
R24275 XThR.Tn[8].n38 XThR.Tn[8].t56 161.106
R24276 XThR.Tn[8].n33 XThR.Tn[8].t61 161.106
R24277 XThR.Tn[8].n28 XThR.Tn[8].t44 161.106
R24278 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R24279 XThR.Tn[8].n18 XThR.Tn[8].t43 161.106
R24280 XThR.Tn[8].n13 XThR.Tn[8].t26 161.106
R24281 XThR.Tn[8].n8 XThR.Tn[8].t49 161.106
R24282 XThR.Tn[8].n6 XThR.Tn[8].t33 161.106
R24283 XThR.Tn[8].n79 XThR.Tn[8].t19 159.978
R24284 XThR.Tn[8].n74 XThR.Tn[8].t25 159.978
R24285 XThR.Tn[8].n69 XThR.Tn[8].t67 159.978
R24286 XThR.Tn[8].n64 XThR.Tn[8].t54 159.978
R24287 XThR.Tn[8].n59 XThR.Tn[8].t16 159.978
R24288 XThR.Tn[8].n54 XThR.Tn[8].t42 159.978
R24289 XThR.Tn[8].n49 XThR.Tn[8].t24 159.978
R24290 XThR.Tn[8].n44 XThR.Tn[8].t64 159.978
R24291 XThR.Tn[8].n39 XThR.Tn[8].t51 159.978
R24292 XThR.Tn[8].n34 XThR.Tn[8].t58 159.978
R24293 XThR.Tn[8].n29 XThR.Tn[8].t41 159.978
R24294 XThR.Tn[8].n24 XThR.Tn[8].t66 159.978
R24295 XThR.Tn[8].n19 XThR.Tn[8].t40 159.978
R24296 XThR.Tn[8].n14 XThR.Tn[8].t22 159.978
R24297 XThR.Tn[8].n9 XThR.Tn[8].t45 159.978
R24298 XThR.Tn[8].n78 XThR.Tn[8].t73 145.038
R24299 XThR.Tn[8].n73 XThR.Tn[8].t35 145.038
R24300 XThR.Tn[8].n68 XThR.Tn[8].t15 145.038
R24301 XThR.Tn[8].n63 XThR.Tn[8].t62 145.038
R24302 XThR.Tn[8].n58 XThR.Tn[8].t30 145.038
R24303 XThR.Tn[8].n53 XThR.Tn[8].t72 145.038
R24304 XThR.Tn[8].n48 XThR.Tn[8].t17 145.038
R24305 XThR.Tn[8].n43 XThR.Tn[8].t63 145.038
R24306 XThR.Tn[8].n38 XThR.Tn[8].t60 145.038
R24307 XThR.Tn[8].n33 XThR.Tn[8].t28 145.038
R24308 XThR.Tn[8].n28 XThR.Tn[8].t52 145.038
R24309 XThR.Tn[8].n23 XThR.Tn[8].t12 145.038
R24310 XThR.Tn[8].n18 XThR.Tn[8].t50 145.038
R24311 XThR.Tn[8].n13 XThR.Tn[8].t34 145.038
R24312 XThR.Tn[8].n8 XThR.Tn[8].t59 145.038
R24313 XThR.Tn[8].n6 XThR.Tn[8].t39 145.038
R24314 XThR.Tn[8].n79 XThR.Tn[8].t32 143.911
R24315 XThR.Tn[8].n74 XThR.Tn[8].t55 143.911
R24316 XThR.Tn[8].n69 XThR.Tn[8].t37 143.911
R24317 XThR.Tn[8].n64 XThR.Tn[8].t18 143.911
R24318 XThR.Tn[8].n59 XThR.Tn[8].t48 143.911
R24319 XThR.Tn[8].n54 XThR.Tn[8].t31 143.911
R24320 XThR.Tn[8].n49 XThR.Tn[8].t38 143.911
R24321 XThR.Tn[8].n44 XThR.Tn[8].t20 143.911
R24322 XThR.Tn[8].n39 XThR.Tn[8].t14 143.911
R24323 XThR.Tn[8].n34 XThR.Tn[8].t47 143.911
R24324 XThR.Tn[8].n29 XThR.Tn[8].t68 143.911
R24325 XThR.Tn[8].n24 XThR.Tn[8].t36 143.911
R24326 XThR.Tn[8].n19 XThR.Tn[8].t65 143.911
R24327 XThR.Tn[8].n14 XThR.Tn[8].t53 143.911
R24328 XThR.Tn[8].n9 XThR.Tn[8].t13 143.911
R24329 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R24330 XThR.Tn[8].n85 XThR.Tn[8].t3 26.5955
R24331 XThR.Tn[8].n85 XThR.Tn[8].t10 26.5955
R24332 XThR.Tn[8].n0 XThR.Tn[8].t6 26.5955
R24333 XThR.Tn[8].n0 XThR.Tn[8].t4 26.5955
R24334 XThR.Tn[8].n1 XThR.Tn[8].t7 26.5955
R24335 XThR.Tn[8].n1 XThR.Tn[8].t5 26.5955
R24336 XThR.Tn[8].n86 XThR.Tn[8].t9 26.5955
R24337 XThR.Tn[8].n86 XThR.Tn[8].t0 26.5955
R24338 XThR.Tn[8].n4 XThR.Tn[8].t1 24.9236
R24339 XThR.Tn[8].n4 XThR.Tn[8].t2 24.9236
R24340 XThR.Tn[8].n3 XThR.Tn[8].t11 24.9236
R24341 XThR.Tn[8].n3 XThR.Tn[8].t8 24.9236
R24342 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R24343 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R24344 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R24345 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R24346 XThR.Tn[8] XThR.Tn[8].n7 5.4407
R24347 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R24348 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R24349 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R24350 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R24351 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R24352 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R24353 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R24354 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R24355 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R24356 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R24357 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R24358 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R24359 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R24360 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R24361 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R24362 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R24363 XThR.Tn[8].n12 XThR.Tn[8] 2.52282
R24364 XThR.Tn[8].n17 XThR.Tn[8] 2.52282
R24365 XThR.Tn[8].n22 XThR.Tn[8] 2.52282
R24366 XThR.Tn[8].n27 XThR.Tn[8] 2.52282
R24367 XThR.Tn[8].n32 XThR.Tn[8] 2.52282
R24368 XThR.Tn[8].n37 XThR.Tn[8] 2.52282
R24369 XThR.Tn[8].n42 XThR.Tn[8] 2.52282
R24370 XThR.Tn[8].n47 XThR.Tn[8] 2.52282
R24371 XThR.Tn[8].n52 XThR.Tn[8] 2.52282
R24372 XThR.Tn[8].n57 XThR.Tn[8] 2.52282
R24373 XThR.Tn[8].n62 XThR.Tn[8] 2.52282
R24374 XThR.Tn[8].n67 XThR.Tn[8] 2.52282
R24375 XThR.Tn[8].n72 XThR.Tn[8] 2.52282
R24376 XThR.Tn[8].n77 XThR.Tn[8] 2.52282
R24377 XThR.Tn[8].n82 XThR.Tn[8] 2.52282
R24378 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R24379 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R24380 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R24381 XThR.Tn[8].n80 XThR.Tn[8] 1.08677
R24382 XThR.Tn[8].n75 XThR.Tn[8] 1.08677
R24383 XThR.Tn[8].n70 XThR.Tn[8] 1.08677
R24384 XThR.Tn[8].n65 XThR.Tn[8] 1.08677
R24385 XThR.Tn[8].n60 XThR.Tn[8] 1.08677
R24386 XThR.Tn[8].n55 XThR.Tn[8] 1.08677
R24387 XThR.Tn[8].n50 XThR.Tn[8] 1.08677
R24388 XThR.Tn[8].n45 XThR.Tn[8] 1.08677
R24389 XThR.Tn[8].n40 XThR.Tn[8] 1.08677
R24390 XThR.Tn[8].n35 XThR.Tn[8] 1.08677
R24391 XThR.Tn[8].n30 XThR.Tn[8] 1.08677
R24392 XThR.Tn[8].n25 XThR.Tn[8] 1.08677
R24393 XThR.Tn[8].n20 XThR.Tn[8] 1.08677
R24394 XThR.Tn[8].n15 XThR.Tn[8] 1.08677
R24395 XThR.Tn[8].n10 XThR.Tn[8] 1.08677
R24396 XThR.Tn[8] XThR.Tn[8].n12 0.839786
R24397 XThR.Tn[8] XThR.Tn[8].n17 0.839786
R24398 XThR.Tn[8] XThR.Tn[8].n22 0.839786
R24399 XThR.Tn[8] XThR.Tn[8].n27 0.839786
R24400 XThR.Tn[8] XThR.Tn[8].n32 0.839786
R24401 XThR.Tn[8] XThR.Tn[8].n37 0.839786
R24402 XThR.Tn[8] XThR.Tn[8].n42 0.839786
R24403 XThR.Tn[8] XThR.Tn[8].n47 0.839786
R24404 XThR.Tn[8] XThR.Tn[8].n52 0.839786
R24405 XThR.Tn[8] XThR.Tn[8].n57 0.839786
R24406 XThR.Tn[8] XThR.Tn[8].n62 0.839786
R24407 XThR.Tn[8] XThR.Tn[8].n67 0.839786
R24408 XThR.Tn[8] XThR.Tn[8].n72 0.839786
R24409 XThR.Tn[8] XThR.Tn[8].n77 0.839786
R24410 XThR.Tn[8] XThR.Tn[8].n82 0.839786
R24411 XThR.Tn[8].n7 XThR.Tn[8] 0.499542
R24412 XThR.Tn[8].n81 XThR.Tn[8] 0.063
R24413 XThR.Tn[8].n76 XThR.Tn[8] 0.063
R24414 XThR.Tn[8].n71 XThR.Tn[8] 0.063
R24415 XThR.Tn[8].n66 XThR.Tn[8] 0.063
R24416 XThR.Tn[8].n61 XThR.Tn[8] 0.063
R24417 XThR.Tn[8].n56 XThR.Tn[8] 0.063
R24418 XThR.Tn[8].n51 XThR.Tn[8] 0.063
R24419 XThR.Tn[8].n46 XThR.Tn[8] 0.063
R24420 XThR.Tn[8].n41 XThR.Tn[8] 0.063
R24421 XThR.Tn[8].n36 XThR.Tn[8] 0.063
R24422 XThR.Tn[8].n31 XThR.Tn[8] 0.063
R24423 XThR.Tn[8].n26 XThR.Tn[8] 0.063
R24424 XThR.Tn[8].n21 XThR.Tn[8] 0.063
R24425 XThR.Tn[8].n16 XThR.Tn[8] 0.063
R24426 XThR.Tn[8].n11 XThR.Tn[8] 0.063
R24427 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R24428 XThR.Tn[8] XThR.Tn[8].n83 0.038
R24429 XThR.Tn[8].n7 XThR.Tn[8] 0.0143889
R24430 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00771154
R24431 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00771154
R24432 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00771154
R24433 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00771154
R24434 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00771154
R24435 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00771154
R24436 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00771154
R24437 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00771154
R24438 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00771154
R24439 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00771154
R24440 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00771154
R24441 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00771154
R24442 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00771154
R24443 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00771154
R24444 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00771154
R24445 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R24446 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R24447 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R24448 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R24449 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R24450 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R24451 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R24452 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R24453 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R24454 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R24455 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R24456 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R24457 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R24458 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R24459 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R24460 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R24461 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R24462 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R24463 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R24464 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R24465 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R24466 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R24467 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R24468 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R24469 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R24470 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R24471 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R24472 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R24473 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R24474 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R24475 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R24476 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R24477 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R24478 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R24479 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R24480 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R24481 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R24482 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R24483 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R24484 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R24485 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R24486 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R24487 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R24488 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R24489 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R24490 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R24491 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R24492 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R24493 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R24494 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R24495 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R24496 data[4].n3 data[4].t0 231.835
R24497 data[4].n0 data[4].t3 230.155
R24498 data[4].n0 data[4].t1 157.856
R24499 data[4].n3 data[4].t2 157.07
R24500 data[4].n1 data[4].n0 152
R24501 data[4].n4 data[4].n3 152
R24502 data[4].n2 data[4].n1 25.6681
R24503 data[4].n4 data[4].n2 10.7642
R24504 data[4].n2 data[4] 2.763
R24505 data[4].n1 data[4] 2.10199
R24506 data[4] data[4].n4 2.01193
R24507 XThR.Tn[13].n87 XThR.Tn[13].n86 256.104
R24508 XThR.Tn[13].n2 XThR.Tn[13].n1 243.68
R24509 XThR.Tn[13].n5 XThR.Tn[13].n3 241.847
R24510 XThR.Tn[13].n2 XThR.Tn[13].n0 205.28
R24511 XThR.Tn[13].n87 XThR.Tn[13].n85 202.094
R24512 XThR.Tn[13].n5 XThR.Tn[13].n4 185
R24513 XThR.Tn[13] XThR.Tn[13].n78 161.363
R24514 XThR.Tn[13] XThR.Tn[13].n73 161.363
R24515 XThR.Tn[13] XThR.Tn[13].n68 161.363
R24516 XThR.Tn[13] XThR.Tn[13].n63 161.363
R24517 XThR.Tn[13] XThR.Tn[13].n58 161.363
R24518 XThR.Tn[13] XThR.Tn[13].n53 161.363
R24519 XThR.Tn[13] XThR.Tn[13].n48 161.363
R24520 XThR.Tn[13] XThR.Tn[13].n43 161.363
R24521 XThR.Tn[13] XThR.Tn[13].n38 161.363
R24522 XThR.Tn[13] XThR.Tn[13].n33 161.363
R24523 XThR.Tn[13] XThR.Tn[13].n28 161.363
R24524 XThR.Tn[13] XThR.Tn[13].n23 161.363
R24525 XThR.Tn[13] XThR.Tn[13].n18 161.363
R24526 XThR.Tn[13] XThR.Tn[13].n13 161.363
R24527 XThR.Tn[13] XThR.Tn[13].n8 161.363
R24528 XThR.Tn[13] XThR.Tn[13].n6 161.363
R24529 XThR.Tn[13].n80 XThR.Tn[13].n79 161.3
R24530 XThR.Tn[13].n75 XThR.Tn[13].n74 161.3
R24531 XThR.Tn[13].n70 XThR.Tn[13].n69 161.3
R24532 XThR.Tn[13].n65 XThR.Tn[13].n64 161.3
R24533 XThR.Tn[13].n60 XThR.Tn[13].n59 161.3
R24534 XThR.Tn[13].n55 XThR.Tn[13].n54 161.3
R24535 XThR.Tn[13].n50 XThR.Tn[13].n49 161.3
R24536 XThR.Tn[13].n45 XThR.Tn[13].n44 161.3
R24537 XThR.Tn[13].n40 XThR.Tn[13].n39 161.3
R24538 XThR.Tn[13].n35 XThR.Tn[13].n34 161.3
R24539 XThR.Tn[13].n30 XThR.Tn[13].n29 161.3
R24540 XThR.Tn[13].n25 XThR.Tn[13].n24 161.3
R24541 XThR.Tn[13].n20 XThR.Tn[13].n19 161.3
R24542 XThR.Tn[13].n15 XThR.Tn[13].n14 161.3
R24543 XThR.Tn[13].n10 XThR.Tn[13].n9 161.3
R24544 XThR.Tn[13].n78 XThR.Tn[13].t56 161.106
R24545 XThR.Tn[13].n73 XThR.Tn[13].t62 161.106
R24546 XThR.Tn[13].n68 XThR.Tn[13].t40 161.106
R24547 XThR.Tn[13].n63 XThR.Tn[13].t27 161.106
R24548 XThR.Tn[13].n58 XThR.Tn[13].t55 161.106
R24549 XThR.Tn[13].n53 XThR.Tn[13].t17 161.106
R24550 XThR.Tn[13].n48 XThR.Tn[13].t59 161.106
R24551 XThR.Tn[13].n43 XThR.Tn[13].t38 161.106
R24552 XThR.Tn[13].n38 XThR.Tn[13].t25 161.106
R24553 XThR.Tn[13].n33 XThR.Tn[13].t30 161.106
R24554 XThR.Tn[13].n28 XThR.Tn[13].t16 161.106
R24555 XThR.Tn[13].n23 XThR.Tn[13].t39 161.106
R24556 XThR.Tn[13].n18 XThR.Tn[13].t14 161.106
R24557 XThR.Tn[13].n13 XThR.Tn[13].t57 161.106
R24558 XThR.Tn[13].n8 XThR.Tn[13].t21 161.106
R24559 XThR.Tn[13].n6 XThR.Tn[13].t64 161.106
R24560 XThR.Tn[13].n79 XThR.Tn[13].t47 159.978
R24561 XThR.Tn[13].n74 XThR.Tn[13].t54 159.978
R24562 XThR.Tn[13].n69 XThR.Tn[13].t36 159.978
R24563 XThR.Tn[13].n64 XThR.Tn[13].t20 159.978
R24564 XThR.Tn[13].n59 XThR.Tn[13].t45 159.978
R24565 XThR.Tn[13].n54 XThR.Tn[13].t73 159.978
R24566 XThR.Tn[13].n49 XThR.Tn[13].t53 159.978
R24567 XThR.Tn[13].n44 XThR.Tn[13].t33 159.978
R24568 XThR.Tn[13].n39 XThR.Tn[13].t18 159.978
R24569 XThR.Tn[13].n34 XThR.Tn[13].t26 159.978
R24570 XThR.Tn[13].n29 XThR.Tn[13].t71 159.978
R24571 XThR.Tn[13].n24 XThR.Tn[13].t35 159.978
R24572 XThR.Tn[13].n19 XThR.Tn[13].t70 159.978
R24573 XThR.Tn[13].n14 XThR.Tn[13].t52 159.978
R24574 XThR.Tn[13].n9 XThR.Tn[13].t12 159.978
R24575 XThR.Tn[13].n78 XThR.Tn[13].t42 145.038
R24576 XThR.Tn[13].n73 XThR.Tn[13].t69 145.038
R24577 XThR.Tn[13].n68 XThR.Tn[13].t50 145.038
R24578 XThR.Tn[13].n63 XThR.Tn[13].t31 145.038
R24579 XThR.Tn[13].n58 XThR.Tn[13].t63 145.038
R24580 XThR.Tn[13].n53 XThR.Tn[13].t41 145.038
R24581 XThR.Tn[13].n48 XThR.Tn[13].t51 145.038
R24582 XThR.Tn[13].n43 XThR.Tn[13].t32 145.038
R24583 XThR.Tn[13].n38 XThR.Tn[13].t29 145.038
R24584 XThR.Tn[13].n33 XThR.Tn[13].t60 145.038
R24585 XThR.Tn[13].n28 XThR.Tn[13].t24 145.038
R24586 XThR.Tn[13].n23 XThR.Tn[13].t49 145.038
R24587 XThR.Tn[13].n18 XThR.Tn[13].t22 145.038
R24588 XThR.Tn[13].n13 XThR.Tn[13].t65 145.038
R24589 XThR.Tn[13].n8 XThR.Tn[13].t28 145.038
R24590 XThR.Tn[13].n6 XThR.Tn[13].t72 145.038
R24591 XThR.Tn[13].n79 XThR.Tn[13].t61 143.911
R24592 XThR.Tn[13].n74 XThR.Tn[13].t23 143.911
R24593 XThR.Tn[13].n69 XThR.Tn[13].t67 143.911
R24594 XThR.Tn[13].n64 XThR.Tn[13].t46 143.911
R24595 XThR.Tn[13].n59 XThR.Tn[13].t15 143.911
R24596 XThR.Tn[13].n54 XThR.Tn[13].t58 143.911
R24597 XThR.Tn[13].n49 XThR.Tn[13].t68 143.911
R24598 XThR.Tn[13].n44 XThR.Tn[13].t48 143.911
R24599 XThR.Tn[13].n39 XThR.Tn[13].t43 143.911
R24600 XThR.Tn[13].n34 XThR.Tn[13].t13 143.911
R24601 XThR.Tn[13].n29 XThR.Tn[13].t37 143.911
R24602 XThR.Tn[13].n24 XThR.Tn[13].t66 143.911
R24603 XThR.Tn[13].n19 XThR.Tn[13].t34 143.911
R24604 XThR.Tn[13].n14 XThR.Tn[13].t19 143.911
R24605 XThR.Tn[13].n9 XThR.Tn[13].t44 143.911
R24606 XThR.Tn[13] XThR.Tn[13].n2 35.7652
R24607 XThR.Tn[13].n85 XThR.Tn[13].t6 26.5955
R24608 XThR.Tn[13].n85 XThR.Tn[13].t4 26.5955
R24609 XThR.Tn[13].n86 XThR.Tn[13].t7 26.5955
R24610 XThR.Tn[13].n86 XThR.Tn[13].t5 26.5955
R24611 XThR.Tn[13].n0 XThR.Tn[13].t2 26.5955
R24612 XThR.Tn[13].n0 XThR.Tn[13].t0 26.5955
R24613 XThR.Tn[13].n1 XThR.Tn[13].t1 26.5955
R24614 XThR.Tn[13].n1 XThR.Tn[13].t3 26.5955
R24615 XThR.Tn[13].n4 XThR.Tn[13].t10 24.9236
R24616 XThR.Tn[13].n4 XThR.Tn[13].t8 24.9236
R24617 XThR.Tn[13].n3 XThR.Tn[13].t11 24.9236
R24618 XThR.Tn[13].n3 XThR.Tn[13].t9 24.9236
R24619 XThR.Tn[13] XThR.Tn[13].n5 22.9615
R24620 XThR.Tn[13].n88 XThR.Tn[13].n87 13.5534
R24621 XThR.Tn[13].n84 XThR.Tn[13] 8.8494
R24622 XThR.Tn[13] XThR.Tn[13].n7 5.4407
R24623 XThR.Tn[13].n12 XThR.Tn[13].n11 4.5005
R24624 XThR.Tn[13].n17 XThR.Tn[13].n16 4.5005
R24625 XThR.Tn[13].n22 XThR.Tn[13].n21 4.5005
R24626 XThR.Tn[13].n27 XThR.Tn[13].n26 4.5005
R24627 XThR.Tn[13].n32 XThR.Tn[13].n31 4.5005
R24628 XThR.Tn[13].n37 XThR.Tn[13].n36 4.5005
R24629 XThR.Tn[13].n42 XThR.Tn[13].n41 4.5005
R24630 XThR.Tn[13].n47 XThR.Tn[13].n46 4.5005
R24631 XThR.Tn[13].n52 XThR.Tn[13].n51 4.5005
R24632 XThR.Tn[13].n57 XThR.Tn[13].n56 4.5005
R24633 XThR.Tn[13].n62 XThR.Tn[13].n61 4.5005
R24634 XThR.Tn[13].n67 XThR.Tn[13].n66 4.5005
R24635 XThR.Tn[13].n72 XThR.Tn[13].n71 4.5005
R24636 XThR.Tn[13].n77 XThR.Tn[13].n76 4.5005
R24637 XThR.Tn[13].n82 XThR.Tn[13].n81 4.5005
R24638 XThR.Tn[13].n83 XThR.Tn[13] 3.70586
R24639 XThR.Tn[13].n88 XThR.Tn[13].n84 2.99115
R24640 XThR.Tn[13].n88 XThR.Tn[13] 2.87153
R24641 XThR.Tn[13].n12 XThR.Tn[13] 2.52282
R24642 XThR.Tn[13].n17 XThR.Tn[13] 2.52282
R24643 XThR.Tn[13].n22 XThR.Tn[13] 2.52282
R24644 XThR.Tn[13].n27 XThR.Tn[13] 2.52282
R24645 XThR.Tn[13].n32 XThR.Tn[13] 2.52282
R24646 XThR.Tn[13].n37 XThR.Tn[13] 2.52282
R24647 XThR.Tn[13].n42 XThR.Tn[13] 2.52282
R24648 XThR.Tn[13].n47 XThR.Tn[13] 2.52282
R24649 XThR.Tn[13].n52 XThR.Tn[13] 2.52282
R24650 XThR.Tn[13].n57 XThR.Tn[13] 2.52282
R24651 XThR.Tn[13].n62 XThR.Tn[13] 2.52282
R24652 XThR.Tn[13].n67 XThR.Tn[13] 2.52282
R24653 XThR.Tn[13].n72 XThR.Tn[13] 2.52282
R24654 XThR.Tn[13].n77 XThR.Tn[13] 2.52282
R24655 XThR.Tn[13].n82 XThR.Tn[13] 2.52282
R24656 XThR.Tn[13].n84 XThR.Tn[13] 2.2734
R24657 XThR.Tn[13] XThR.Tn[13].n88 1.50638
R24658 XThR.Tn[13].n80 XThR.Tn[13] 1.08677
R24659 XThR.Tn[13].n75 XThR.Tn[13] 1.08677
R24660 XThR.Tn[13].n70 XThR.Tn[13] 1.08677
R24661 XThR.Tn[13].n65 XThR.Tn[13] 1.08677
R24662 XThR.Tn[13].n60 XThR.Tn[13] 1.08677
R24663 XThR.Tn[13].n55 XThR.Tn[13] 1.08677
R24664 XThR.Tn[13].n50 XThR.Tn[13] 1.08677
R24665 XThR.Tn[13].n45 XThR.Tn[13] 1.08677
R24666 XThR.Tn[13].n40 XThR.Tn[13] 1.08677
R24667 XThR.Tn[13].n35 XThR.Tn[13] 1.08677
R24668 XThR.Tn[13].n30 XThR.Tn[13] 1.08677
R24669 XThR.Tn[13].n25 XThR.Tn[13] 1.08677
R24670 XThR.Tn[13].n20 XThR.Tn[13] 1.08677
R24671 XThR.Tn[13].n15 XThR.Tn[13] 1.08677
R24672 XThR.Tn[13].n10 XThR.Tn[13] 1.08677
R24673 XThR.Tn[13] XThR.Tn[13].n12 0.839786
R24674 XThR.Tn[13] XThR.Tn[13].n17 0.839786
R24675 XThR.Tn[13] XThR.Tn[13].n22 0.839786
R24676 XThR.Tn[13] XThR.Tn[13].n27 0.839786
R24677 XThR.Tn[13] XThR.Tn[13].n32 0.839786
R24678 XThR.Tn[13] XThR.Tn[13].n37 0.839786
R24679 XThR.Tn[13] XThR.Tn[13].n42 0.839786
R24680 XThR.Tn[13] XThR.Tn[13].n47 0.839786
R24681 XThR.Tn[13] XThR.Tn[13].n52 0.839786
R24682 XThR.Tn[13] XThR.Tn[13].n57 0.839786
R24683 XThR.Tn[13] XThR.Tn[13].n62 0.839786
R24684 XThR.Tn[13] XThR.Tn[13].n67 0.839786
R24685 XThR.Tn[13] XThR.Tn[13].n72 0.839786
R24686 XThR.Tn[13] XThR.Tn[13].n77 0.839786
R24687 XThR.Tn[13] XThR.Tn[13].n82 0.839786
R24688 XThR.Tn[13].n7 XThR.Tn[13] 0.499542
R24689 XThR.Tn[13].n81 XThR.Tn[13] 0.063
R24690 XThR.Tn[13].n76 XThR.Tn[13] 0.063
R24691 XThR.Tn[13].n71 XThR.Tn[13] 0.063
R24692 XThR.Tn[13].n66 XThR.Tn[13] 0.063
R24693 XThR.Tn[13].n61 XThR.Tn[13] 0.063
R24694 XThR.Tn[13].n56 XThR.Tn[13] 0.063
R24695 XThR.Tn[13].n51 XThR.Tn[13] 0.063
R24696 XThR.Tn[13].n46 XThR.Tn[13] 0.063
R24697 XThR.Tn[13].n41 XThR.Tn[13] 0.063
R24698 XThR.Tn[13].n36 XThR.Tn[13] 0.063
R24699 XThR.Tn[13].n31 XThR.Tn[13] 0.063
R24700 XThR.Tn[13].n26 XThR.Tn[13] 0.063
R24701 XThR.Tn[13].n21 XThR.Tn[13] 0.063
R24702 XThR.Tn[13].n16 XThR.Tn[13] 0.063
R24703 XThR.Tn[13].n11 XThR.Tn[13] 0.063
R24704 XThR.Tn[13].n83 XThR.Tn[13] 0.0540714
R24705 XThR.Tn[13] XThR.Tn[13].n83 0.038
R24706 XThR.Tn[13].n7 XThR.Tn[13] 0.0143889
R24707 XThR.Tn[13].n81 XThR.Tn[13].n80 0.00771154
R24708 XThR.Tn[13].n76 XThR.Tn[13].n75 0.00771154
R24709 XThR.Tn[13].n71 XThR.Tn[13].n70 0.00771154
R24710 XThR.Tn[13].n66 XThR.Tn[13].n65 0.00771154
R24711 XThR.Tn[13].n61 XThR.Tn[13].n60 0.00771154
R24712 XThR.Tn[13].n56 XThR.Tn[13].n55 0.00771154
R24713 XThR.Tn[13].n51 XThR.Tn[13].n50 0.00771154
R24714 XThR.Tn[13].n46 XThR.Tn[13].n45 0.00771154
R24715 XThR.Tn[13].n41 XThR.Tn[13].n40 0.00771154
R24716 XThR.Tn[13].n36 XThR.Tn[13].n35 0.00771154
R24717 XThR.Tn[13].n31 XThR.Tn[13].n30 0.00771154
R24718 XThR.Tn[13].n26 XThR.Tn[13].n25 0.00771154
R24719 XThR.Tn[13].n21 XThR.Tn[13].n20 0.00771154
R24720 XThR.Tn[13].n16 XThR.Tn[13].n15 0.00771154
R24721 XThR.Tn[13].n11 XThR.Tn[13].n10 0.00771154
R24722 data[0].n1 data[0].t0 230.155
R24723 data[0].n0 data[0].t2 228.463
R24724 data[0].n1 data[0].t1 157.856
R24725 data[0].n0 data[0].t3 157.07
R24726 data[0].n2 data[0].n1 152.768
R24727 data[0].n4 data[0].n0 152.256
R24728 data[0].n3 data[0].n2 24.1398
R24729 data[0].n4 data[0].n3 9.48418
R24730 data[0] data[0].n4 6.1445
R24731 data[0].n2 data[0] 5.6325
R24732 data[0].n3 data[0] 2.638
R24733 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R24734 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R24735 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R24736 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R24737 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R24738 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R24739 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R24740 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R24741 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24742 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24743 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24744 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24745 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24746 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24747 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24748 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24749 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24750 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24751 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24752 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24753 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24754 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24755 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24756 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24757 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24758 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24759 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24760 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24761 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24762 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24763 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24764 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24765 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24766 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24767 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24768 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24769 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24770 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24771 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24772 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24773 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24774 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24775 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24776 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24777 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24778 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24779 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24780 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24781 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24782 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24783 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24784 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24785 data[6].n0 data[6].t0 230.576
R24786 data[6].n0 data[6].t1 158.275
R24787 data[6].n1 data[6].n0 152
R24788 data[6].n1 data[6] 11.9995
R24789 data[6] data[6].n1 6.66717
R24790 data[1].n4 data[1].t2 230.576
R24791 data[1].n1 data[1].t0 230.363
R24792 data[1].n0 data[1].t4 229.369
R24793 data[1].n4 data[1].t5 158.275
R24794 data[1].n1 data[1].t3 158.064
R24795 data[1].n0 data[1].t1 157.07
R24796 data[1].n2 data[1].n1 153.28
R24797 data[1].n7 data[1].n0 153.147
R24798 data[1].n5 data[1].n4 152
R24799 data[1].n7 data[1].n6 16.3874
R24800 data[1].n6 data[1].n5 14.9641
R24801 data[1].n3 data[1].n2 9.3005
R24802 data[1].n6 data[1].n3 6.49639
R24803 data[1] data[1].n7 3.24826
R24804 data[1].n2 data[1] 2.92621
R24805 data[1].n3 data[1] 2.15819
R24806 data[1].n5 data[1] 2.13383
R24807 data[2].n0 data[2].t0 230.576
R24808 data[2].n0 data[2].t1 158.275
R24809 data[2].n1 data[2].n0 152
R24810 data[2].n1 data[2] 12.7714
R24811 data[2] data[2].n1 2.13383
R24812 data[5].n4 data[5].t2 230.576
R24813 data[5].n1 data[5].t0 230.363
R24814 data[5].n0 data[5].t1 229.369
R24815 data[5].n4 data[5].t5 158.275
R24816 data[5].n1 data[5].t3 158.064
R24817 data[5].n0 data[5].t4 157.07
R24818 data[5].n2 data[5].n1 152.256
R24819 data[5].n7 data[5].n0 152.238
R24820 data[5].n5 data[5].n4 152
R24821 data[5].n7 data[5].n6 16.3874
R24822 data[5].n6 data[5].n5 14.6005
R24823 data[5].n3 data[5].n2 9.3005
R24824 data[5].n5 data[5] 6.66717
R24825 data[5].n6 data[5].n3 6.49639
R24826 data[5].n2 data[5] 6.1445
R24827 data[5] data[5].n7 5.68939
R24828 data[5].n3 data[5] 2.28319
R24829 bias[1].n0 bias[1].t1 81.1889
R24830 bias[1].n2 bias[1].t0 81.1889
R24831 bias[1].n1 bias[1] 9.32819
R24832 bias[1].n1 bias[1].n0 1.06523
R24833 bias[1].n2 bias[1].n1 0.895589
R24834 bias[1] bias[1].n2 0.301839
R24835 bias[1].n0 bias[1] 0.221482
R24836 data[3].n0 data[3].t1 230.576
R24837 data[3].n0 data[3].t0 158.275
R24838 data[3].n1 data[3].n0 153.553
R24839 data[3].n1 data[3] 11.6078
R24840 data[3] data[3].n1 2.90959
R24841 data[7].n0 data[7].t0 230.576
R24842 data[7].n0 data[7].t1 158.275
R24843 data[7].n1 data[7].n0 152
R24844 data[7].n1 data[7] 11.9995
R24845 data[7] data[7].n1 6.66717
R24846 bias[2].n0 bias[2].t1 136.779
R24847 bias[2].n2 bias[2].t0 136.779
R24848 bias[2].n1 bias[2] 7.84903
R24849 bias[2].n1 bias[2].n0 1.2438
R24850 bias[2].n2 bias[2].n1 0.717018
R24851 bias[2] bias[2].n2 0.301839
R24852 bias[2].n0 bias[2] 0.221482
R24853 bias[0].n0 bias[0].t0 57.5124
R24854 bias[0].n2 bias[0].t1 57.5124
R24855 bias[0].n1 bias[0] 11.1563
R24856 bias[0].n2 bias[0].n1 1.10095
R24857 bias[0].n1 bias[0].n0 0.859875
R24858 bias[0] bias[0].n2 0.301839
R24859 bias[0].n0 bias[0] 0.221482
C0 XA.XIR[13].XIC[3].icell.Ien Vbias 0.19151f
C1 XA.XIR[8].XIC[1].icell.Ien VPWR 0.21079f
C2 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04035f
C3 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01768f
C4 XA.XIR[3].XIC[3].icell.Ien VPWR 0.21079f
C5 XA.XIR[6].XIC[8].icell.PUM VPWR 0.01079f
C6 XThC.Tn[4] XThR.Tn[9] 0.39123f
C7 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02601f
C8 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.04573f
C9 XThC.Tn[0] XThR.Tn[8] 0.39119f
C10 XA.XIR[15].XIC[9].icell.Ien VPWR 0.3396f
C11 XThR.XTB7.A XThR.Tn[4] 0.02736f
C12 XA.XIR[11].XIC[6].icell.Ien Vbias 0.19151f
C13 XA.XIR[0].XIC[9].icell.Ien Iout 0.06712f
C14 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.14207f
C15 XThC.XTBN.Y a_9827_9569# 0.22873f
C16 XThR.XTB7.A a_n1049_7493# 0.0127f
C17 XA.XIR[4].XIC[12].icell.Ien VPWR 0.21079f
C18 XA.XIR[10].XIC[8].icell.Ien Vbias 0.19151f
C19 XA.XIR[3].XIC[1].icell.PDM VPWR 0.01373f
C20 XA.XIR[8].XIC[3].icell.PDM VPWR 0.01373f
C21 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C22 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.14207f
C23 XA.XIR[2].XIC[7].icell.PDM VPWR 0.01373f
C24 XA.XIR[13].XIC[4].icell.PUM VPWR 0.01079f
C25 XA.XIR[7].XIC[12].icell.Ien Iout 0.06763f
C26 XA.XIR[8].XIC[6].icell.Ien VPWR 0.21079f
C27 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C28 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04035f
C29 XA.XIR[11].XIC[7].icell.PUM VPWR 0.01079f
C30 XA.XIR[2].XIC[10].icell.Ien Vbias 0.19151f
C31 XA.XIR[10].XIC[11].icell.Ien Iout 0.06763f
C32 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C33 XA.XIR[9].XIC_15.icell.Ien VPWR 0.2801f
C34 XA.XIR[3].XIC[1].icell.Ien Iout 0.06763f
C35 XA.XIR[1].XIC[12].icell.Ien Vbias 0.19162f
C36 XA.XIR[10].XIC[9].icell.PUM VPWR 0.01079f
C37 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C38 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C39 XThR.XTB7.B XThR.XTBN.A 0.35142f
C40 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01687f
C41 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C42 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.14207f
C43 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C44 XA.XIR[0].XIC[8].icell.Ien VPWR 0.21227f
C45 XThR.XTB7.B XThR.Tn[6] 0.04822f
C46 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04035f
C47 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C48 XA.XIR[12].XIC[10].icell.Ien VPWR 0.21079f
C49 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.02965f
C50 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04035f
C51 XA.XIR[7].XIC[11].icell.Ien VPWR 0.21079f
C52 XA.XIR[2].XIC[11].icell.PUM VPWR 0.01079f
C53 XThC.Tn[12] XThR.Tn[7] 0.39123f
C54 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C55 XA.XIR[1].XIC[13].icell.PUM VPWR 0.01079f
C56 XA.XIR[7].XIC[6].icell.PDM Vbias 0.03922f
C57 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04035f
C58 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02601f
C59 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C60 XThC.XTB7.B XThC.Tn[10] 0.06229f
C61 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.1155f
C62 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C63 XA.XIR[15].XIC[4].icell.PDM Vbias 0.03922f
C64 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C65 XA.XIR[6].XIC[13].icell.PDM Vbias 0.03922f
C66 XA.XIR[15].XIC[13].icell.PUM VPWR 0.01079f
C67 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.14207f
C68 XA.XIR[3].XIC[0].icell.Ien VPWR 0.21079f
C69 XThR.Tn[8] VPWR 10.5606f
C70 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C71 XA.XIR[13].XIC[13].icell.Ien Iout 0.06763f
C72 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02601f
C73 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.04573f
C74 XA.XIR[14].XIC[10].icell.PDM Vbias 0.03922f
C75 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02601f
C76 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C77 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08254f
C78 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C79 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C80 XThR.XTB3.Y data[4] 0.03253f
C81 XA.XIR[11].XIC[1].icell.Ien VPWR 0.21079f
C82 bias[0] Vbias 0.82324f
C83 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.14207f
C84 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04035f
C85 XA.XIR[9].XIC[2].icell.PDM Vbias 0.03922f
C86 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.04261f
C87 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.04627f
C88 XA.XIR[7].XIC[7].icell.PDM VPWR 0.01373f
C89 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C90 a_3773_9615# XThC.Tn[1] 0.26251f
C91 XA.XIR[12].XIC[13].icell.Ien Vbias 0.19151f
C92 XThR.Tn[14] a_n997_715# 0.1927f
C93 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.14207f
C94 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01714f
C95 XA.XIR[3].XIC[9].icell.Ien Iout 0.06763f
C96 XA.XIR[6].XIC[14].icell.PDM VPWR 0.01349f
C97 XThR.Tn[11] a_n997_2667# 0.19413f
C98 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.04573f
C99 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.14207f
C100 XThC.Tn[11] XThR.Tn[3] 0.39123f
C101 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C102 XA.XIR[2].XIC[2].icell.Ien Iout 0.06763f
C103 XA.XIR[15].XIC[14].icell.Ien VPWR 0.33336f
C104 XA.XIR[1].XIC[7].icell.PDM Vbias 0.03922f
C105 XA.XIR[1].XIC[4].icell.Ien Iout 0.06763f
C106 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01545f
C107 XA.XIR[6].XIC[12].icell.Ien Vbias 0.19151f
C108 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.14207f
C109 XA.XIR[9].XIC[3].icell.PDM VPWR 0.01373f
C110 XA.XIR[4].XIC[7].icell.PDM Vbias 0.03922f
C111 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.04573f
C112 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C113 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C114 XA.XIR[8].XIC[12].icell.Ien Iout 0.06763f
C115 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02602f
C116 XThC.Tn[14] XThR.Tn[0] 0.39146f
C117 XA.XIR[3].XIC_15.icell.PDM Vbias 0.03927f
C118 XThC.XTB4.Y a_8963_9569# 0.07199f
C119 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C120 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C121 XA.XIR[14].XIC[6].icell.Ien Vbias 0.19151f
C122 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C123 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C124 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02601f
C125 XA.XIR[13].XIC[8].icell.Ien Vbias 0.19151f
C126 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04035f
C127 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C128 XA.XIR[3].XIC[8].icell.Ien VPWR 0.21079f
C129 XA.XIR[1].XIC[8].icell.PDM VPWR 0.01373f
C130 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C131 XA.XIR[6].XIC[13].icell.PUM VPWR 0.01079f
C132 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C133 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C134 XA.XIR[0].XIC[14].icell.Ien Iout 0.06712f
C135 XA.XIR[4].XIC[8].icell.PDM VPWR 0.01373f
C136 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C137 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04035f
C138 XA.XIR[15].XIC[11].icell.PUM VPWR 0.01079f
C139 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C140 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C141 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C142 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02601f
C143 XA.XIR[1].XIC[3].icell.Ien VPWR 0.21079f
C144 XA.XIR[14].XIC[7].icell.PUM VPWR 0.01079f
C145 XThC.XTB7.Y a_6243_10571# 0.01283f
C146 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C147 XA.XIR[13].XIC[11].icell.Ien Iout 0.06763f
C148 a_n1049_7493# XThR.Tn[2] 0.26564f
C149 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C150 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C151 XThR.XTBN.Y XThR.Tn[6] 0.59879f
C152 XA.XIR[12].XIC_15.icell.Ien VPWR 0.2801f
C153 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04035f
C154 XA.XIR[13].XIC[9].icell.PUM VPWR 0.01079f
C155 XA.XIR[8].XIC[11].icell.Ien VPWR 0.21079f
C156 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C157 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C158 VPWR data[4] 0.53035f
C159 XA.XIR[2].XIC_15.icell.Ien Vbias 0.19187f
C160 XThC.Tn[13] XThR.Tn[2] 0.39125f
C161 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C162 XA.XIR[12].XIC[11].icell.Ien Vbias 0.19151f
C163 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C164 a_n997_3755# VPWR 0.01462f
C165 XThR.XTB2.Y VPWR 0.99107f
C166 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04035f
C167 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.04573f
C168 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02601f
C169 XA.XIR[15].XIC[12].icell.Ien VPWR 0.3396f
C170 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C171 XA.XIR[0].XIC[13].icell.Ien VPWR 0.21044f
C172 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C173 XA.XIR[6].XIC[4].icell.Ien Iout 0.06763f
C174 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02601f
C175 XThR.XTBN.A XThR.Tn[10] 0.12147f
C176 XA.XIR[10].XIC[1].icell.PDM Vbias 0.03922f
C177 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.04574f
C178 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.14207f
C179 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.14207f
C180 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.1155f
C181 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02601f
C182 data[6] data[7] 0.04128f
C183 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04035f
C184 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02602f
C185 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.0176f
C186 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02601f
C187 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C188 a_n1049_5611# VPWR 0.71932f
C189 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.14207f
C190 XA.XIR[5].XIC[5].icell.Ien Vbias 0.19151f
C191 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C192 XThC.Tn[9] XThR.Tn[6] 0.39123f
C193 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C194 XA.XIR[14].XIC[1].icell.Ien VPWR 0.21134f
C195 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C196 XA.XIR[10].XIC[2].icell.PDM VPWR 0.01373f
C197 XThC.Tn[11] XThR.Tn[11] 0.39123f
C198 XA.XIR[11].XIC[3].icell.Ien Iout 0.06763f
C199 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C200 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.04573f
C201 XThR.XTBN.Y XThR.Tn[4] 0.60348f
C202 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C203 XThC.Tn[1] XThR.Tn[7] 0.39123f
C204 XA.XIR[6].XIC[3].icell.Ien VPWR 0.21079f
C205 XThR.Tn[5] Vbias 1.38578f
C206 XA.XIR[10].XIC[5].icell.Ien Iout 0.06763f
C207 XThR.XTBN.Y a_n1049_7493# 0.08456f
C208 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C209 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C210 XA.XIR[0].XIC[9].icell.PDM Vbias 0.03922f
C211 XA.XIR[5].XIC[6].icell.PUM VPWR 0.01079f
C212 XThC.XTB7.B a_7651_9569# 0.01152f
C213 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C214 XA.XIR[3].XIC[14].icell.Ien Iout 0.06763f
C215 XThC.XTB5.Y XThC.Tn[12] 0.32158f
C216 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.03366f
C217 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.14207f
C218 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C219 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C220 XA.XIR[2].XIC[7].icell.Ien Iout 0.06763f
C221 XThC.Tn[14] XThR.Tn[1] 0.39129f
C222 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.04573f
C223 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C224 XA.XIR[1].XIC[9].icell.Ien Iout 0.06763f
C225 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C226 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02601f
C227 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C228 XA.XIR[2].XIC[1].icell.Ien VPWR 0.21079f
C229 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.13138f
C230 XA.XIR[0].XIC[10].icell.PDM VPWR 0.01334f
C231 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C232 XA.XIR[11].XIC[2].icell.Ien VPWR 0.21079f
C233 XA.XIR[15].XIC[10].icell.Ien VPWR 0.3396f
C234 XThC.Tn[14] XThR.Tn[12] 0.39123f
C235 XThC.XTB7.A VPWR 0.87269f
C236 XA.XIR[10].XIC[4].icell.Ien VPWR 0.21079f
C237 XThC.Tn[0] XThR.Tn[3] 0.39121f
C238 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.04573f
C239 XThR.XTBN.A a_n997_1803# 0.09118f
C240 XThC.Tn[9] XThR.Tn[4] 0.39123f
C241 XThC.XTBN.Y XThC.Tn[12] 0.45161f
C242 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C243 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04035f
C244 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C245 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02601f
C246 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04035f
C247 XA.XIR[3].XIC[13].icell.Ien VPWR 0.21079f
C248 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C249 XA.XIR[2].XIC[6].icell.Ien VPWR 0.21079f
C250 XThC.Tn[3] XThR.Tn[0] 0.39147f
C251 XThC.Tn[13] XThR.Tn[10] 0.39123f
C252 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C253 XThC.Tn[5] XThR.Tn[5] 0.39123f
C254 a_n997_715# VPWR 0.02818f
C255 XA.XIR[1].XIC[8].icell.Ien VPWR 0.21079f
C256 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.36378f
C257 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.14207f
C258 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.03366f
C259 XA.XIR[6].XIC[0].icell.PDM Vbias 0.03915f
C260 XA.XIR[15].XIC[13].icell.Ien Vbias 0.15955f
C261 XA.XIR[5].XIC[7].icell.PDM Vbias 0.03922f
C262 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02601f
C263 XA.XIR[13].XIC[1].icell.PDM Vbias 0.03922f
C264 XA.XIR[15].XIC[0].icell.PUM VPWR 0.01079f
C265 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C266 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.14207f
C267 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02601f
C268 XA.XIR[12].XIC[6].icell.PDM Vbias 0.03922f
C269 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C270 a_5949_9615# VPWR 0.7053f
C271 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.04573f
C272 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.04573f
C273 XA.XIR[6].XIC[1].icell.PDM VPWR 0.01373f
C274 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C275 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04035f
C276 XA.XIR[6].XIC[9].icell.Ien Iout 0.06763f
C277 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C278 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.04629f
C279 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.14207f
C280 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.14207f
C281 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C282 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C283 XA.XIR[5].XIC[8].icell.PDM VPWR 0.01373f
C284 Vbias Iout 73.9689f
C285 XThC.Tn[2] XThR.Tn[2] 0.39125f
C286 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C287 XA.XIR[13].XIC[2].icell.PDM VPWR 0.01373f
C288 XThC.Tn[11] XThR.Tn[14] 0.39123f
C289 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.04576f
C290 XA.XIR[14].XIC[3].icell.Ien Iout 0.06763f
C291 XThC.XTB5.A VPWR 0.82807f
C292 XThR.Tn[3] VPWR 9.69701f
C293 XThC.XTB6.Y Vbias 0.01779f
C294 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C295 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C296 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C297 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C298 XA.XIR[12].XIC[7].icell.PDM VPWR 0.01373f
C299 XA.XIR[5].XIC[10].icell.Ien Vbias 0.19151f
C300 XA.XIR[13].XIC[5].icell.Ien Iout 0.06763f
C301 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C302 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C303 XA.XIR[3].XIC[2].icell.PDM Vbias 0.03922f
C304 XA.XIR[8].XIC[4].icell.PDM Vbias 0.03922f
C305 XThR.XTB7.Y VPWR 1.14813f
C306 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.04573f
C307 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.13184f
C308 XA.XIR[2].XIC[8].icell.PDM Vbias 0.03922f
C309 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C310 XA.XIR[11].XIC[8].icell.Ien Iout 0.06763f
C311 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C312 XA.XIR[15].XIC_15.icell.Ien VPWR 0.39202f
C313 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04035f
C314 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C315 XA.XIR[12].XIC[5].icell.Ien Vbias 0.19151f
C316 XA.XIR[6].XIC[8].icell.Ien VPWR 0.21079f
C317 XThC.Tn[7] XThR.Tn[6] 0.39123f
C318 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.04573f
C319 XA.XIR[5].XIC[11].icell.PUM VPWR 0.01079f
C320 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.04573f
C321 XThC.XTBN.A XThC.Tn[9] 0.12399f
C322 XThC.XTBN.Y a_10915_9569# 0.21503f
C323 XA.XIR[8].XIC[5].icell.PDM VPWR 0.01373f
C324 XThC.Tn[0] XThR.Tn[11] 0.39119f
C325 XA.XIR[3].XIC[3].icell.PDM VPWR 0.01373f
C326 XA.XIR[15].XIC[11].icell.Ien Vbias 0.15955f
C327 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C328 XA.XIR[14].XIC[2].icell.Ien VPWR 0.21134f
C329 XThC.XTB4.Y Vbias 0.01643f
C330 XThC.XTB7.A XThC.XTB7.B 0.35844f
C331 XA.XIR[2].XIC[9].icell.PDM VPWR 0.01373f
C332 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C333 XA.XIR[13].XIC[4].icell.Ien VPWR 0.21079f
C334 XA.XIR[2].XIC[12].icell.Ien Iout 0.06763f
C335 XA.XIR[12].XIC[6].icell.PUM VPWR 0.01079f
C336 XA.XIR[1].XIC[14].icell.Ien Iout 0.06763f
C337 XThC.Tn[5] Iout 0.02219f
C338 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.04573f
C339 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02601f
C340 VPWR data[0] 0.52929f
C341 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01768f
C342 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21445f
C343 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C344 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C345 XA.XIR[11].XIC[7].icell.Ien VPWR 0.21079f
C346 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04035f
C347 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C348 XThC.XTB6.Y XThC.Tn[5] 0.20249f
C349 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.02965f
C350 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C351 XA.XIR[10].XIC[9].icell.Ien VPWR 0.21079f
C352 XThC.Tn[13] XThR.Tn[13] 0.39123f
C353 XA.XIR[12].XIC[1].icell.Ien Iout 0.06763f
C354 XThC.Tn[3] XThR.Tn[1] 0.39128f
C355 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C356 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.04573f
C357 a_n997_2667# VPWR 0.01739f
C358 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.36378f
C359 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C360 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04035f
C361 XA.XIR[5].XIC[2].icell.Ien Iout 0.06763f
C362 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.04573f
C363 XThC.Tn[3] XThR.Tn[12] 0.39123f
C364 XThC.Tn[12] XThR.Tn[8] 0.39123f
C365 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.40495f
C366 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04035f
C367 XA.XIR[2].XIC[11].icell.Ien VPWR 0.21079f
C368 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.04573f
C369 XThC.XTBN.Y XThC.Tn[1] 0.4915f
C370 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04035f
C371 XA.XIR[1].XIC[13].icell.Ien VPWR 0.21079f
C372 XA.XIR[7].XIC[8].icell.PDM Vbias 0.03922f
C373 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.14207f
C374 XA.XIR[9].XIC[1].icell.Ien Vbias 0.19151f
C375 XThC.Tn[7] XThR.Tn[4] 0.39123f
C376 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C377 XA.XIR[4].XIC[3].icell.Ien Vbias 0.19151f
C378 XA.XIR[15].XIC[6].icell.PDM Vbias 0.03922f
C379 XA.XIR[6].XIC_15.icell.PDM Vbias 0.03927f
C380 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.03758f
C381 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C382 XThC.Tn[2] XThR.Tn[10] 0.39123f
C383 XA.XIR[12].XIC[0].icell.Ien VPWR 0.21079f
C384 XThC.XTB6.Y a_10051_9569# 0.07626f
C385 XThR.Tn[11] VPWR 10.6372f
C386 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.14207f
C387 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04035f
C388 XA.XIR[9].XIC[4].icell.PDM Vbias 0.03922f
C389 XA.XIR[7].XIC[9].icell.PDM VPWR 0.01373f
C390 XThC.XTB2.Y Vbias 0.01483f
C391 XThC.XTB5.A XThC.XTB7.B 0.30355f
C392 XA.XIR[9].XIC[2].icell.PUM VPWR 0.01079f
C393 XA.XIR[9].XIC[6].icell.Ien Vbias 0.19151f
C394 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01714f
C395 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C396 XA.XIR[4].XIC[4].icell.PUM VPWR 0.01079f
C397 XA.XIR[6].XIC[14].icell.Ien Iout 0.06763f
C398 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.14207f
C399 XA.XIR[10].XIC[13].icell.PUM VPWR 0.01079f
C400 XA.XIR[1].XIC[9].icell.PDM Vbias 0.03922f
C401 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C402 XA.XIR[14].XIC[8].icell.Ien Iout 0.06763f
C403 XA.XIR[9].XIC[5].icell.PDM VPWR 0.01373f
C404 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C405 XA.XIR[5].XIC_15.icell.Ien Vbias 0.19187f
C406 XA.XIR[7].XIC[2].icell.Ien Vbias 0.19151f
C407 XA.XIR[4].XIC[9].icell.PDM Vbias 0.03922f
C408 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.04573f
C409 XA.XIR[9].XIC[7].icell.PUM VPWR 0.01079f
C410 XThR.XTBN.A a_n997_3979# 0.02087f
C411 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.04573f
C412 XA.XIR[12].XIC_15.icell.PDM Vbias 0.03927f
C413 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C414 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C415 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C416 XThC.Tn[0] XThR.Tn[14] 0.39118f
C417 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04035f
C418 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02601f
C419 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C420 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.04573f
C421 XA.XIR[1].XIC[10].icell.PDM VPWR 0.01373f
C422 XA.XIR[6].XIC[13].icell.Ien VPWR 0.21079f
C423 XA.XIR[10].XIC[14].icell.Ien VPWR 0.20455f
C424 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02601f
C425 XA.XIR[4].XIC[10].icell.PDM VPWR 0.01373f
C426 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.0176f
C427 XA.XIR[7].XIC[3].icell.PUM VPWR 0.01079f
C428 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04035f
C429 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02602f
C430 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02601f
C431 XThR.Tn[9] Vbias 1.38584f
C432 XThC.XTB7.B data[0] 0.0138f
C433 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01768f
C434 XA.XIR[14].XIC[7].icell.Ien VPWR 0.21134f
C435 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C436 XA.XIR[13].XIC[9].icell.Ien VPWR 0.21079f
C437 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04035f
C438 XThC.Tn[11] VPWR 7.99883f
C439 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.04261f
C440 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C441 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01687f
C442 XThC.XTBN.A XThC.Tn[7] 0.01451f
C443 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.03366f
C444 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.14207f
C445 XThR.XTB6.A data[5] 0.37233f
C446 XA.XIR[15].XIC[0].icell.Ien Vbias 0.15953f
C447 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04035f
C448 XThR.XTBN.A XThR.Tn[7] 0.01439f
C449 XThR.XTBN.A a_n997_2891# 0.01719f
C450 XA.XIR[10].XIC[11].icell.PUM VPWR 0.01079f
C451 XThR.Tn[6] XThR.Tn[7] 0.10592f
C452 VPWR bias[2] 1.67895f
C453 XA.XIR[10].XIC[3].icell.PDM Vbias 0.03922f
C454 XThC.Tn[4] Vbias 0.33409f
C455 XA.XIR[5].XIC[7].icell.Ien Iout 0.06763f
C456 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.04573f
C457 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04023f
C458 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04035f
C459 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C460 XThC.Tn[2] XThR.Tn[13] 0.39123f
C461 XA.XIR[15].XIC[1].icell.PUM VPWR 0.01079f
C462 XA.XIR[5].XIC[1].icell.Ien VPWR 0.21079f
C463 XA.XIR[15].XIC[5].icell.Ien Vbias 0.15955f
C464 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.14207f
C465 XThR.Tn[14] VPWR 10.8855f
C466 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.04575f
C467 XA.XIR[11].XIC[0].icell.PDM VPWR 0.01373f
C468 XA.XIR[4].XIC[8].icell.Ien Vbias 0.19151f
C469 XThC.Tn[5] XThR.Tn[9] 0.39123f
C470 XA.XIR[12].XIC[2].icell.Ien Iout 0.06763f
C471 XThC.Tn[1] XThR.Tn[8] 0.39123f
C472 XA.XIR[10].XIC[4].icell.PDM VPWR 0.01373f
C473 XA.XIR[10].XIC[12].icell.Ien VPWR 0.21079f
C474 XThR.XTB2.Y a_n1335_8107# 0.01006f
C475 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C476 XA.XIR[8].XIC[2].icell.Ien Vbias 0.19151f
C477 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02601f
C478 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.04573f
C479 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C480 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.14207f
C481 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C482 XA.XIR[13].XIC[13].icell.PUM VPWR 0.01079f
C483 XA.XIR[0].XIC[11].icell.PDM Vbias 0.03922f
C484 XA.XIR[15].XIC[6].icell.PUM VPWR 0.01079f
C485 XA.XIR[5].XIC[6].icell.Ien VPWR 0.21079f
C486 XThC.XTB7.B a_8739_9569# 0.0168f
C487 XA.XIR[9].XIC[11].icell.Ien Vbias 0.19151f
C488 XA.XIR[4].XIC[9].icell.PUM VPWR 0.01079f
C489 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.04573f
C490 XA.XIR[12].XIC[14].icell.PDM Vbias 0.03922f
C491 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.04573f
C492 XA.XIR[0].XIC[4].icell.Ien Vbias 0.19186f
C493 XA.XIR[8].XIC[3].icell.PUM VPWR 0.01079f
C494 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.14207f
C495 XA.XIR[15].XIC_15.icell.PDM Vbias 0.03927f
C496 XThC.Tn[4] XThC.Tn[5] 0.31866f
C497 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.34325f
C498 XThR.XTB2.Y a_n1049_7787# 0.2342f
C499 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02601f
C500 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.13138f
C501 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01653f
C502 XA.XIR[7].XIC[7].icell.Ien Vbias 0.19151f
C503 XA.XIR[13].XIC[14].icell.Ien VPWR 0.20455f
C504 XA.XIR[9].XIC[12].icell.PUM VPWR 0.01079f
C505 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.04261f
C506 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02602f
C507 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.14207f
C508 XA.XIR[0].XIC[5].icell.PUM VPWR 0.01038f
C509 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C510 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C511 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04035f
C512 XThR.Tn[0] Iout 1.10107f
C513 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C514 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C515 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04035f
C516 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C517 XThC.Tn[13] XThR.Tn[7] 0.39123f
C518 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C519 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.04573f
C520 XThC.XTB7.B XThC.Tn[11] 0.03651f
C521 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.04573f
C522 XA.XIR[7].XIC[8].icell.PUM VPWR 0.01079f
C523 data[2] data[3] 0.04128f
C524 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C525 XA.XIR[10].XIC[10].icell.Ien VPWR 0.21079f
C526 XA.XIR[6].XIC[2].icell.PDM Vbias 0.03922f
C527 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C528 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.14207f
C529 XA.XIR[5].XIC[9].icell.PDM Vbias 0.03922f
C530 XA.XIR[13].XIC[11].icell.PUM VPWR 0.01079f
C531 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.04036f
C532 a_3773_9615# XThC.Tn[2] 0.01043f
C533 XA.XIR[9].XIC[3].icell.Ien Iout 0.06763f
C534 XA.XIR[13].XIC[3].icell.PDM Vbias 0.03922f
C535 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C536 XThR.XTB3.Y VPWR 1.08016f
C537 XA.XIR[12].XIC[8].icell.PDM Vbias 0.03922f
C538 XThC.Tn[12] XThR.Tn[3] 0.39123f
C539 XThR.XTB5.A XThR.XTB6.A 1.80461f
C540 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08254f
C541 XThC.Tn[0] VPWR 7.09956f
C542 XA.XIR[6].XIC[3].icell.PDM VPWR 0.01373f
C543 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.04036f
C544 XA.XIR[14].XIC[0].icell.PDM VPWR 0.01373f
C545 XA.XIR[5].XIC[10].icell.PDM VPWR 0.01373f
C546 XA.XIR[5].XIC[12].icell.Ien Iout 0.06763f
C547 XThC.Tn[8] XThR.Tn[5] 0.39123f
C548 XA.XIR[13].XIC[4].icell.PDM VPWR 0.01373f
C549 XA.XIR[10].XIC[13].icell.Ien Vbias 0.19151f
C550 XA.XIR[3].XIC[4].icell.Ien Vbias 0.19151f
C551 XA.XIR[13].XIC[12].icell.Ien VPWR 0.21079f
C552 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02601f
C553 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.04573f
C554 XA.XIR[12].XIC[9].icell.PDM VPWR 0.01373f
C555 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C556 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C557 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C558 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.04573f
C559 XA.XIR[9].XIC[2].icell.Ien VPWR 0.21079f
C560 XA.XIR[12].XIC[13].icell.PDM Vbias 0.03922f
C561 XA.XIR[3].XIC[4].icell.PDM Vbias 0.03922f
C562 XA.XIR[4].XIC[13].icell.Ien Vbias 0.19151f
C563 XA.XIR[8].XIC[6].icell.PDM Vbias 0.03922f
C564 XA.XIR[12].XIC[7].icell.Ien Iout 0.06763f
C565 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C566 XA.XIR[2].XIC[10].icell.PDM Vbias 0.03922f
C567 XA.XIR[8].XIC[7].icell.Ien Vbias 0.19151f
C568 XA.XIR[15].XIC[14].icell.PDM Vbias 0.03922f
C569 XA.XIR[3].XIC[5].icell.PUM VPWR 0.01079f
C570 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04035f
C571 XA.XIR[5].XIC[11].icell.Ien VPWR 0.21079f
C572 XA.XIR[3].XIC[5].icell.PDM VPWR 0.01373f
C573 XA.XIR[8].XIC[7].icell.PDM VPWR 0.01373f
C574 XA.XIR[4].XIC[14].icell.PUM VPWR 0.01079f
C575 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C576 XThR.XTB7.B data[6] 0.07481f
C577 XA.XIR[2].XIC[11].icell.PDM VPWR 0.01373f
C578 XA.XIR[0].XIC[9].icell.Ien Vbias 0.19186f
C579 XThC.Tn[14] XThR.Tn[2] 0.39126f
C580 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C581 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04035f
C582 XA.XIR[8].XIC[8].icell.PUM VPWR 0.01079f
C583 XA.XIR[1].XIC[0].icell.Ien Iout 0.06763f
C584 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C585 XA.XIR[12].XIC[6].icell.Ien VPWR 0.21079f
C586 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.04574f
C587 XA.XIR[10].XIC_15.icell.Ien VPWR 0.2801f
C588 XA.XIR[4].XIC[0].icell.Ien Iout 0.06763f
C589 XThR.XTB6.Y a_n997_1579# 0.07626f
C590 XThR.Tn[1] Iout 1.10105f
C591 XA.XIR[7].XIC[12].icell.Ien Vbias 0.19151f
C592 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.04573f
C593 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C594 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C595 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.14207f
C596 XThR.Tn[12] Iout 1.10102f
C597 XA.XIR[0].XIC[10].icell.PUM VPWR 0.01038f
C598 XA.XIR[10].XIC[11].icell.Ien Vbias 0.19151f
C599 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C600 XA.XIR[13].XIC[10].icell.Ien VPWR 0.21079f
C601 XA.XIR[3].XIC[1].icell.Ien Vbias 0.19151f
C602 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04035f
C603 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C604 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04035f
C605 XA.XIR[15].XIC[2].icell.Ien Iout 0.07153f
C606 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C607 XThC.Tn[10] XThR.Tn[6] 0.39123f
C608 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04035f
C609 XA.XIR[7].XIC[13].icell.PUM VPWR 0.01079f
C610 XA.XIR[4].XIC[5].icell.Ien Iout 0.06763f
C611 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C612 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.1155f
C613 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.04036f
C614 XThC.Tn[12] XThR.Tn[11] 0.39123f
C615 XA.XIR[7].XIC[10].icell.PDM Vbias 0.03922f
C616 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C617 XThC.Tn[2] XThR.Tn[7] 0.39123f
C618 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04023f
C619 XA.XIR[15].XIC[8].icell.PDM Vbias 0.03922f
C620 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.14207f
C621 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08254f
C622 XA.XIR[3].XIC[2].icell.PUM VPWR 0.01079f
C623 XThC.Tn[8] Iout 0.02193f
C624 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C625 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.14207f
C626 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C627 XThC.XTB6.Y XThC.Tn[8] 0.02463f
C628 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C629 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.04573f
C630 XA.XIR[9].XIC[8].icell.Ien Iout 0.06763f
C631 XA.XIR[9].XIC[6].icell.PDM Vbias 0.03922f
C632 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04023f
C633 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C634 XA.XIR[13].XIC[13].icell.Ien Vbias 0.19151f
C635 XA.XIR[7].XIC[11].icell.PDM VPWR 0.01373f
C636 XThR.XTB7.Y a_n1319_5317# 0.01283f
C637 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.14207f
C638 XA.XIR[12].XIC[12].icell.PDM Vbias 0.03922f
C639 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02601f
C640 XA.XIR[4].XIC[4].icell.Ien VPWR 0.21079f
C641 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01714f
C642 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C643 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02602f
C644 XA.XIR[7].XIC[4].icell.Ien Iout 0.06763f
C645 XA.XIR[15].XIC[13].icell.PDM Vbias 0.03922f
C646 XA.XIR[3].XIC[9].icell.Ien Vbias 0.19151f
C647 XA.XIR[1].XIC[11].icell.PDM Vbias 0.03922f
C648 XThC.Tn[1] XThR.Tn[3] 0.39123f
C649 XA.XIR[9].XIC[7].icell.PDM VPWR 0.01373f
C650 XThC.XTBN.Y XThC.Tn[13] 0.40384f
C651 XThC.Tn[10] XThR.Tn[4] 0.39123f
C652 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C653 XA.XIR[4].XIC[11].icell.PDM Vbias 0.03922f
C654 XA.XIR[2].XIC[2].icell.Ien Vbias 0.19151f
C655 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C656 XThC.XTB6.A data[1] 0.37233f
C657 XA.XIR[9].XIC[7].icell.Ien VPWR 0.21079f
C658 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C659 XA.XIR[1].XIC[4].icell.Ien Vbias 0.19162f
C660 XThC.XTB4.Y XThC.Tn[8] 0.01307f
C661 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C662 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C663 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.14207f
C664 XThC.Tn[4] XThR.Tn[0] 0.39146f
C665 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C666 XThC.Tn[14] XThR.Tn[10] 0.39123f
C667 XA.XIR[8].XIC[12].icell.Ien Vbias 0.19151f
C668 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04035f
C669 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02601f
C670 XThC.Tn[6] XThR.Tn[5] 0.39123f
C671 XA.XIR[3].XIC[10].icell.PUM VPWR 0.01079f
C672 XA.XIR[1].XIC[12].icell.PDM VPWR 0.01373f
C673 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C674 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C675 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.04627f
C676 XThC.Tn[11] XThC.Tn[12] 0.12311f
C677 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C678 XA.XIR[2].XIC[3].icell.PUM VPWR 0.01079f
C679 XA.XIR[7].XIC[3].icell.Ien VPWR 0.21079f
C680 XA.XIR[4].XIC[12].icell.PDM VPWR 0.01373f
C681 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04035f
C682 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C683 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C684 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C685 XThC.XTB7.B VPWR 1.33382f
C686 XA.XIR[13].XIC_15.icell.Ien VPWR 0.2801f
C687 XA.XIR[1].XIC[5].icell.PUM VPWR 0.01079f
C688 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C689 XA.XIR[0].XIC[14].icell.Ien Vbias 0.19186f
C690 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C691 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04035f
C692 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04035f
C693 XA.XIR[8].XIC[13].icell.PUM VPWR 0.01079f
C694 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C695 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.04626f
C696 XA.XIR[13].XIC[11].icell.Ien Vbias 0.19151f
C697 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C698 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.14207f
C699 XThR.XTBN.A XThR.Tn[8] 0.1369f
C700 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02601f
C701 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.14207f
C702 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04035f
C703 XThC.Tn[3] XThR.Tn[2] 0.39125f
C704 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.04036f
C705 XA.XIR[11].XIC[1].icell.PDM Vbias 0.03922f
C706 XThC.XTB7.Y a_6243_9615# 0.27822f
C707 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01693f
C708 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.1155f
C709 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.14207f
C710 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.14207f
C711 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.0404f
C712 XThC.Tn[12] XThR.Tn[14] 0.39123f
C713 XA.XIR[10].XIC[5].icell.PDM Vbias 0.03922f
C714 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02601f
C715 XA.XIR[15].XIC[7].icell.Ien Iout 0.07153f
C716 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C717 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04035f
C718 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.04573f
C719 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.14207f
C720 XA.XIR[4].XIC[10].icell.Ien Iout 0.06763f
C721 XA.XIR[6].XIC[4].icell.Ien Vbias 0.19151f
C722 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C723 XA.XIR[15].XIC[1].icell.Ien VPWR 0.3396f
C724 XA.XIR[0].XIC[1].icell.Ien Iout 0.06712f
C725 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.13194f
C726 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.04573f
C727 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C728 XA.XIR[12].XIC[11].icell.PDM Vbias 0.03922f
C729 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C730 XA.XIR[8].XIC[4].icell.Ien Iout 0.06763f
C731 XA.XIR[11].XIC[2].icell.PDM VPWR 0.01373f
C732 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C733 XA.XIR[10].XIC[6].icell.PDM VPWR 0.01373f
C734 XA.XIR[15].XIC[12].icell.PDM Vbias 0.03922f
C735 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02602f
C736 XThC.XTBN.A XThC.Tn[10] 0.12208f
C737 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13586f
C738 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C739 XA.XIR[9].XIC[13].icell.Ien Iout 0.06763f
C740 XThC.Tn[1] XThR.Tn[11] 0.39123f
C741 XA.XIR[6].XIC[5].icell.PUM VPWR 0.01079f
C742 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02601f
C743 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C744 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C745 XA.XIR[0].XIC[13].icell.PDM Vbias 0.03922f
C746 XA.XIR[11].XIC[3].icell.Ien Vbias 0.19151f
C747 XA.XIR[15].XIC[6].icell.Ien VPWR 0.3396f
C748 XA.XIR[0].XIC[6].icell.Ien Iout 0.06712f
C749 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.04573f
C750 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.14207f
C751 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.0279f
C752 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C753 XA.XIR[10].XIC[5].icell.Ien Vbias 0.19151f
C754 XA.XIR[4].XIC[9].icell.Ien VPWR 0.21079f
C755 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.04574f
C756 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C757 XThC.Tn[6] Iout 0.02211f
C758 XA.XIR[0].XIC[0].icell.Ien VPWR 0.21044f
C759 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C760 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.04573f
C761 XA.XIR[7].XIC[9].icell.Ien Iout 0.06763f
C762 XA.XIR[8].XIC[3].icell.Ien VPWR 0.21079f
C763 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C764 XThC.XTB6.Y XThC.Tn[6] 0.01038f
C765 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02601f
C766 XA.XIR[3].XIC[14].icell.Ien Vbias 0.19151f
C767 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C768 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C769 XThC.Tn[14] XThR.Tn[13] 0.39123f
C770 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02601f
C771 XThC.Tn[4] XThR.Tn[1] 0.39128f
C772 XA.XIR[0].XIC[14].icell.PDM VPWR 0.0131f
C773 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C774 XA.XIR[11].XIC[4].icell.PUM VPWR 0.01079f
C775 XA.XIR[2].XIC[7].icell.Ien Vbias 0.19151f
C776 XThC.Tn[8] XThR.Tn[9] 0.39123f
C777 XA.XIR[9].XIC[12].icell.Ien VPWR 0.21079f
C778 XA.XIR[10].XIC[6].icell.PUM VPWR 0.01079f
C779 XA.XIR[1].XIC[9].icell.Ien Vbias 0.19162f
C780 XThR.XTBN.A data[4] 0.02581f
C781 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C782 XThC.Tn[4] XThR.Tn[12] 0.39123f
C783 XThC.Tn[13] XThR.Tn[8] 0.39123f
C784 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.14207f
C785 XA.XIR[2].XIC[0].icell.Ien Iout 0.06763f
C786 XA.XIR[0].XIC[5].icell.Ien VPWR 0.21065f
C787 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C788 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04035f
C789 XThR.XTBN.A a_n997_3755# 0.01939f
C790 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C791 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01768f
C792 XThC.XTBN.Y XThC.Tn[2] 0.49f
C793 XA.XIR[10].XIC[1].icell.Ien Iout 0.06763f
C794 XThR.XTB7.A XThR.Tn[5] 0.02751f
C795 XA.XIR[2].XIC[8].icell.PUM VPWR 0.01079f
C796 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C797 XA.XIR[7].XIC[8].icell.Ien VPWR 0.21079f
C798 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.36378f
C799 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C800 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C801 XA.XIR[1].XIC[10].icell.PUM VPWR 0.01079f
C802 XA.XIR[0].XIC[0].icell.PUM VPWR 0.01038f
C803 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02601f
C804 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.0404f
C805 XThC.Tn[3] XThR.Tn[10] 0.39123f
C806 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04035f
C807 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02601f
C808 XThC.XTB3.Y XThC.Tn[10] 0.29566f
C809 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.04573f
C810 XA.XIR[6].XIC[4].icell.PDM Vbias 0.03922f
C811 XA.XIR[14].XIC[1].icell.PDM Vbias 0.03922f
C812 XA.XIR[5].XIC[11].icell.PDM Vbias 0.03922f
C813 XThR.XTB7.A data[5] 0.06538f
C814 a_n1049_8581# VPWR 0.72063f
C815 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C816 XA.XIR[13].XIC[5].icell.PDM Vbias 0.03922f
C817 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04035f
C818 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.14207f
C819 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C820 XA.XIR[12].XIC[10].icell.PDM Vbias 0.03922f
C821 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.04573f
C822 XA.XIR[11].XIC[13].icell.Ien Iout 0.06763f
C823 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C824 XA.XIR[10].XIC[0].icell.Ien VPWR 0.21079f
C825 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C826 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.04573f
C827 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C828 XA.XIR[3].XIC[6].icell.Ien Iout 0.06763f
C829 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C830 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.14207f
C831 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.14207f
C832 XA.XIR[6].XIC[5].icell.PDM VPWR 0.01373f
C833 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.04573f
C834 XA.XIR[15].XIC[11].icell.PDM Vbias 0.03922f
C835 XA.XIR[14].XIC[2].icell.PDM VPWR 0.01373f
C836 XA.XIR[5].XIC[12].icell.PDM VPWR 0.01373f
C837 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C838 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.14207f
C839 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C840 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.04573f
C841 XA.XIR[13].XIC[6].icell.PDM VPWR 0.01373f
C842 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C843 XA.XIR[6].XIC[9].icell.Ien Vbias 0.19151f
C844 XA.XIR[4].XIC_15.icell.Ien Iout 0.0694f
C845 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.14207f
C846 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.04573f
C847 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C848 XThC.Tn[1] XThR.Tn[14] 0.39123f
C849 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C850 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02601f
C851 XA.XIR[8].XIC[9].icell.Ien Iout 0.06763f
C852 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01244f
C853 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C854 XA.XIR[3].XIC[6].icell.PDM Vbias 0.03922f
C855 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02803f
C856 XA.XIR[8].XIC[8].icell.PDM Vbias 0.03922f
C857 XThR.XTB2.Y a_n1049_7493# 0.02133f
C858 XA.XIR[14].XIC[3].icell.Ien Vbias 0.19151f
C859 XA.XIR[2].XIC[12].icell.PDM Vbias 0.03922f
C860 XA.XIR[13].XIC[5].icell.Ien Vbias 0.19151f
C861 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C862 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C863 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.13181f
C864 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04035f
C865 XA.XIR[3].XIC[5].icell.Ien VPWR 0.21079f
C866 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.04573f
C867 XA.XIR[6].XIC[10].icell.PUM VPWR 0.01079f
C868 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C869 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.04573f
C870 XA.XIR[0].XIC[11].icell.Ien Iout 0.06712f
C871 XA.XIR[11].XIC[8].icell.Ien Vbias 0.19151f
C872 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02601f
C873 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13586f
C874 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C875 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C876 XThC.Tn[12] VPWR 7.97657f
C877 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.04629f
C878 XA.XIR[3].XIC[7].icell.PDM VPWR 0.01373f
C879 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C880 XA.XIR[4].XIC[14].icell.Ien VPWR 0.20455f
C881 XA.XIR[14].XIC[4].icell.PUM VPWR 0.01079f
C882 XA.XIR[8].XIC[9].icell.PDM VPWR 0.01373f
C883 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C884 XA.XIR[2].XIC[13].icell.PDM VPWR 0.01373f
C885 XThC.XTBN.A a_7651_9569# 0.02087f
C886 XA.XIR[13].XIC[6].icell.PUM VPWR 0.01079f
C887 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.04575f
C888 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04035f
C889 XA.XIR[7].XIC[14].icell.Ien Iout 0.06763f
C890 XA.XIR[8].XIC[8].icell.Ien VPWR 0.21079f
C891 XThR.XTB6.Y a_n1049_5611# 0.26831f
C892 XA.XIR[11].XIC[11].icell.Ien Iout 0.06763f
C893 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C894 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07604f
C895 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C896 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C897 XA.XIR[2].XIC[12].icell.Ien Vbias 0.19151f
C898 XA.XIR[11].XIC[9].icell.PUM VPWR 0.01079f
C899 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.40931f
C900 XA.XIR[13].XIC[1].icell.Ien Iout 0.06763f
C901 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04035f
C902 XA.XIR[1].XIC[14].icell.Ien Vbias 0.19162f
C903 XThC.Tn[5] Vbias 0.32211f
C904 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.36378f
C905 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.14207f
C906 XA.XIR[0].XIC[10].icell.Ien VPWR 0.21044f
C907 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C908 XThC.Tn[3] XThR.Tn[13] 0.39123f
C909 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04035f
C910 XA.XIR[12].XIC[1].icell.Ien Vbias 0.19151f
C911 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.04573f
C912 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04035f
C913 XA.XIR[2].XIC[13].icell.PUM VPWR 0.01079f
C914 XA.XIR[7].XIC[13].icell.Ien VPWR 0.21079f
C915 XThC.Tn[6] XThR.Tn[9] 0.39123f
C916 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02601f
C917 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.14207f
C918 XThC.Tn[2] XThR.Tn[8] 0.39123f
C919 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01768f
C920 XA.XIR[5].XIC[2].icell.Ien Vbias 0.19151f
C921 XA.XIR[7].XIC[12].icell.PDM Vbias 0.03922f
C922 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.04573f
C923 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C924 XA.XIR[14].XIC[13].icell.Ien Iout 0.06763f
C925 XA.XIR[15].XIC[10].icell.PDM Vbias 0.03922f
C926 XA.XIR[13].XIC[0].icell.Ien VPWR 0.21079f
C927 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C928 XThC.XTBN.Y a_2979_9615# 0.0607f
C929 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C930 XA.XIR[12].XIC[2].icell.PUM VPWR 0.01079f
C931 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C932 XA.XIR[1].XIC[1].icell.Ien Iout 0.06763f
C933 XA.XIR[10].XIC[2].icell.Ien Iout 0.06763f
C934 XA.XIR[9].XIC[8].icell.PDM Vbias 0.03922f
C935 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.14207f
C936 XThR.XTB5.A XThR.XTB7.A 0.07862f
C937 XA.XIR[0].XIC[0].icell.PDM Vbias 0.03917f
C938 XA.XIR[5].XIC[3].icell.PUM VPWR 0.01079f
C939 a_9827_9569# XThC.Tn[12] 0.20217f
C940 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C941 XA.XIR[7].XIC[13].icell.PDM VPWR 0.01373f
C942 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.04573f
C943 XThC.Tn[0] XThC.Tn[1] 0.88261f
C944 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.14207f
C945 XA.XIR[3].XIC[11].icell.Ien Iout 0.06763f
C946 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.04573f
C947 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.14207f
C948 XA.XIR[2].XIC[4].icell.Ien Iout 0.06763f
C949 a_n1049_7787# VPWR 0.72275f
C950 XA.XIR[1].XIC[13].icell.PDM Vbias 0.03922f
C951 XA.XIR[1].XIC[6].icell.Ien Iout 0.06763f
C952 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13586f
C953 XA.XIR[6].XIC[14].icell.Ien Vbias 0.19151f
C954 XA.XIR[9].XIC[9].icell.PDM VPWR 0.01373f
C955 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02602f
C956 XA.XIR[0].XIC[1].icell.PDM VPWR 0.01334f
C957 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C958 XA.XIR[4].XIC[13].icell.PDM Vbias 0.03922f
C959 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C960 XA.XIR[8].XIC[14].icell.Ien Iout 0.06763f
C961 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.04573f
C962 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02601f
C963 XThC.Tn[14] XThR.Tn[7] 0.39123f
C964 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C965 XThC.XTB5.A a_7331_10587# 0.01243f
C966 XA.XIR[14].XIC[8].icell.Ien Vbias 0.19151f
C967 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C968 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04035f
C969 XThR.XTBN.Y XThR.Tn[5] 0.5991f
C970 XA.XIR[3].XIC[10].icell.Ien VPWR 0.21079f
C971 XA.XIR[1].XIC[14].icell.PDM VPWR 0.01349f
C972 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01768f
C973 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C974 XA.XIR[10].XIC[14].icell.PDM VPWR 0.01349f
C975 XThR.XTBN.A a_n997_2667# 0.01679f
C976 XThR.Tn[3] XThR.Tn[4] 0.10942f
C977 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02601f
C978 XA.XIR[2].XIC[3].icell.Ien VPWR 0.21079f
C979 XA.XIR[4].XIC[14].icell.PDM VPWR 0.01349f
C980 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.01601f
C981 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04035f
C982 XA.XIR[14].XIC[11].icell.Ien Iout 0.06763f
C983 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07604f
C984 XA.XIR[1].XIC[5].icell.Ien VPWR 0.21079f
C985 XA.XIR[14].XIC[9].icell.PUM VPWR 0.01079f
C986 XA.XIR[6].XIC[1].icell.Ien Iout 0.06763f
C987 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.04036f
C988 XA.XIR[8].XIC[13].icell.Ien VPWR 0.21079f
C989 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C990 XThC.Tn[13] XThR.Tn[3] 0.39123f
C991 XThR.Tn[2] Iout 1.10104f
C992 XThC.XTB7.A XThC.XTBN.A 0.197f
C993 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02602f
C994 XThC.XTB1.Y a_7651_9569# 0.06353f
C995 XThC.Tn[1] VPWR 7.02414f
C996 XA.XIR[1].XIC[0].icell.PUM VPWR 0.01079f
C997 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02601f
C998 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C999 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04035f
C1000 XA.XIR[4].XIC[0].icell.PUM VPWR 0.01079f
C1001 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C1002 XThR.XTBN.A XThR.Tn[11] 0.11968f
C1003 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02601f
C1004 XThC.Tn[9] XThR.Tn[5] 0.39123f
C1005 XA.XIR[11].XIC[3].icell.PDM Vbias 0.03922f
C1006 XA.XIR[0].XIC_15.icell.Ien VPWR 0.27821f
C1007 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.04573f
C1008 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02801f
C1009 XA.XIR[6].XIC[6].icell.Ien Iout 0.06763f
C1010 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04035f
C1011 XA.XIR[10].XIC[7].icell.PDM Vbias 0.03922f
C1012 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.14207f
C1013 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.14207f
C1014 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.14207f
C1015 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02601f
C1016 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C1017 XA.XIR[6].XIC[0].icell.Ien VPWR 0.21079f
C1018 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C1019 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04035f
C1020 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C1021 XThR.XTB5.A XThR.XTB7.B 0.30355f
C1022 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.27178f
C1023 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.02965f
C1024 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.14207f
C1025 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02601f
C1026 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.04573f
C1027 a_6243_9615# XThC.Tn[6] 0.26385f
C1028 XA.XIR[5].XIC[7].icell.Ien Vbias 0.19151f
C1029 XA.XIR[13].XIC[2].icell.Ien Iout 0.06763f
C1030 XA.XIR[11].XIC[4].icell.PDM VPWR 0.01373f
C1031 XA.XIR[10].XIC[8].icell.PDM VPWR 0.01373f
C1032 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12344f
C1033 XA.XIR[11].XIC[5].icell.Ien Iout 0.06763f
C1034 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C1035 XA.XIR[10].XIC[7].icell.Ien Iout 0.06763f
C1036 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C1037 XA.XIR[6].XIC[5].icell.Ien VPWR 0.21079f
C1038 XA.XIR[12].XIC[2].icell.Ien Vbias 0.19151f
C1039 XA.XIR[0].XIC_15.icell.PDM Vbias 0.03927f
C1040 XA.XIR[5].XIC[8].icell.PUM VPWR 0.01079f
C1041 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02602f
C1042 XThC.XTB7.Y Vbias 0.0196f
C1043 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02601f
C1044 bias[2] bias[1] 0.67657f
C1045 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.04573f
C1046 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02601f
C1047 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C1048 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.14207f
C1049 XA.XIR[2].XIC[0].icell.PDM VPWR 0.01373f
C1050 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02601f
C1051 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.04573f
C1052 XThC.XTB5.A XThC.XTBN.A 0.06305f
C1053 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01687f
C1054 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02601f
C1055 XA.XIR[2].XIC[9].icell.Ien Iout 0.06763f
C1056 XA.XIR[10].XIC[13].icell.PDM VPWR 0.01373f
C1057 XThC.XTB7.A XThC.Tn[2] 0.1255f
C1058 XA.XIR[1].XIC[11].icell.Ien Iout 0.06763f
C1059 XA.XIR[12].XIC[3].icell.PUM VPWR 0.01079f
C1060 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C1061 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.04575f
C1062 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C1063 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04035f
C1064 XA.XIR[11].XIC[4].icell.Ien VPWR 0.21079f
C1065 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02601f
C1066 XA.XIR[13].XIC[14].icell.PDM VPWR 0.01349f
C1067 XA.XIR[10].XIC[6].icell.Ien VPWR 0.21079f
C1068 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.14207f
C1069 XThC.Tn[11] XThR.Tn[6] 0.39123f
C1070 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C1071 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C1072 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C1073 XA.XIR[3].XIC_15.icell.Ien VPWR 0.2801f
C1074 XThC.Tn[13] XThR.Tn[11] 0.39123f
C1075 XThR.Tn[10] Iout 1.10102f
C1076 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C1077 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.40971f
C1078 XThR.Tn[0] Vbias 1.38698f
C1079 XA.XIR[2].XIC[8].icell.Ien VPWR 0.21079f
C1080 XThC.Tn[3] XThR.Tn[7] 0.39123f
C1081 XThC.Tn[9] Iout 0.02193f
C1082 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.40905f
C1083 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C1084 XA.XIR[1].XIC[10].icell.Ien VPWR 0.21079f
C1085 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04035f
C1086 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.14207f
C1087 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02601f
C1088 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C1089 XA.XIR[6].XIC[6].icell.PDM Vbias 0.03922f
C1090 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C1091 XThC.XTBN.A data[0] 0.02545f
C1092 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C1093 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02803f
C1094 XA.XIR[14].XIC[3].icell.PDM Vbias 0.03922f
C1095 XA.XIR[5].XIC[13].icell.PDM Vbias 0.03922f
C1096 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.04573f
C1097 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.04573f
C1098 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1099 XA.XIR[13].XIC[7].icell.PDM Vbias 0.03922f
C1100 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02601f
C1101 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C1102 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.14207f
C1103 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04035f
C1104 XThR.XTB7.B XThR.Tn[9] 0.0565f
C1105 XA.XIR[7].XIC[0].icell.PDM VPWR 0.01373f
C1106 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C1107 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C1108 XA.XIR[9].XIC[3].icell.Ien Vbias 0.19151f
C1109 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02601f
C1110 XA.XIR[6].XIC[7].icell.PDM VPWR 0.01373f
C1111 XThC.Tn[2] XThR.Tn[3] 0.39123f
C1112 XA.XIR[6].XIC[11].icell.Ien Iout 0.06763f
C1113 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.14207f
C1114 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.14207f
C1115 XA.XIR[5].XIC[14].icell.PDM VPWR 0.01349f
C1116 XA.XIR[14].XIC[4].icell.PDM VPWR 0.01373f
C1117 XThC.XTBN.Y XThC.Tn[14] 0.42542f
C1118 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.04573f
C1119 XThC.Tn[11] XThR.Tn[4] 0.39123f
C1120 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.04574f
C1121 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C1122 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C1123 XA.XIR[13].XIC[8].icell.PDM VPWR 0.01373f
C1124 XA.XIR[1].XIC[0].icell.PDM Vbias 0.03915f
C1125 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C1126 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.04261f
C1127 XA.XIR[14].XIC[5].icell.Ien Iout 0.06763f
C1128 XThC.XTB7.Y a_10051_9569# 0.013f
C1129 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.14207f
C1130 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C1131 XA.XIR[4].XIC[0].icell.PDM Vbias 0.03915f
C1132 XThC.Tn[5] XThR.Tn[0] 0.39148f
C1133 XA.XIR[5].XIC[12].icell.Ien Vbias 0.19151f
C1134 XA.XIR[13].XIC[7].icell.Ien Iout 0.06763f
C1135 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.14207f
C1136 XThC.Tn[7] XThR.Tn[5] 0.39123f
C1137 XA.XIR[9].XIC[4].icell.PUM VPWR 0.01079f
C1138 XA.XIR[3].XIC[8].icell.PDM Vbias 0.03922f
C1139 XA.XIR[8].XIC[10].icell.PDM Vbias 0.03922f
C1140 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08254f
C1141 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C1142 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02601f
C1143 XA.XIR[2].XIC[14].icell.PDM Vbias 0.03922f
C1144 XA.XIR[10].XIC[12].icell.PDM VPWR 0.01373f
C1145 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C1146 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02601f
C1147 XA.XIR[1].XIC[1].icell.PDM VPWR 0.01373f
C1148 XA.XIR[12].XIC[7].icell.Ien Vbias 0.19151f
C1149 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.04573f
C1150 XA.XIR[6].XIC[10].icell.Ien VPWR 0.21079f
C1151 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.14207f
C1152 XA.XIR[5].XIC[13].icell.PUM VPWR 0.01079f
C1153 XA.XIR[4].XIC[1].icell.PDM VPWR 0.01373f
C1154 XA.XIR[13].XIC[13].icell.PDM VPWR 0.01373f
C1155 XThC.XTB3.Y data[0] 0.03253f
C1156 XA.XIR[3].XIC[9].icell.PDM VPWR 0.01373f
C1157 XA.XIR[8].XIC[11].icell.PDM VPWR 0.01373f
C1158 XA.XIR[14].XIC[4].icell.Ien VPWR 0.21134f
C1159 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C1160 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07604f
C1161 XThC.XTBN.A a_8739_9569# 0.01719f
C1162 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.0404f
C1163 XA.XIR[13].XIC[6].icell.Ien VPWR 0.21079f
C1164 XA.XIR[2].XIC[14].icell.Ien Iout 0.06763f
C1165 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C1166 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04035f
C1167 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C1168 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01768f
C1169 XA.XIR[12].XIC[8].icell.PUM VPWR 0.01079f
C1170 XThC.Tn[4] XThR.Tn[2] 0.39125f
C1171 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01687f
C1172 XA.XIR[14].XIC[0].icell.Ien Iout 0.06763f
C1173 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C1174 XA.XIR[11].XIC[9].icell.Ien VPWR 0.21079f
C1175 XThC.Tn[13] XThR.Tn[14] 0.39123f
C1176 XA.XIR[1].XIC[0].icell.Ien Vbias 0.1916f
C1177 XThR.Tn[13] Iout 1.10105f
C1178 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01687f
C1179 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C1180 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C1181 XA.XIR[4].XIC[0].icell.Ien Vbias 0.19149f
C1182 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C1183 XThR.Tn[1] Vbias 1.38583f
C1184 a_7875_9569# XThC.Tn[9] 0.19271f
C1185 XThC.XTB2.Y XThC.Tn[9] 0.292f
C1186 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.04036f
C1187 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C1188 XA.XIR[2].XIC[0].icell.PUM VPWR 0.01079f
C1189 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C1190 XA.XIR[5].XIC[4].icell.Ien Iout 0.06763f
C1191 XThR.Tn[12] Vbias 1.38583f
C1192 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04035f
C1193 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C1194 XA.XIR[2].XIC[13].icell.Ien VPWR 0.21079f
C1195 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02601f
C1196 XThC.Tn[0] XThR.Tn[6] 0.3912f
C1197 XThR.XTBN.Y XThR.Tn[9] 0.48046f
C1198 XA.XIR[1].XIC[1].icell.PUM VPWR 0.01079f
C1199 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08254f
C1200 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C1201 XA.XIR[15].XIC[2].icell.Ien Vbias 0.15955f
C1202 XA.XIR[1].XIC_15.icell.Ien VPWR 0.2801f
C1203 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C1204 XThC.XTBN.A XThC.Tn[11] 0.11997f
C1205 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.14207f
C1206 XA.XIR[7].XIC[14].icell.PDM Vbias 0.03922f
C1207 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.14207f
C1208 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02602f
C1209 XA.XIR[4].XIC[1].icell.PUM VPWR 0.01079f
C1210 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C1211 XA.XIR[4].XIC[5].icell.Ien Vbias 0.19151f
C1212 XThC.Tn[2] XThR.Tn[11] 0.39123f
C1213 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.3624f
C1214 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02601f
C1215 XThC.XTBN.Y a_4067_9615# 0.08456f
C1216 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C1217 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13586f
C1218 VPWR bias[1] 1.65687f
C1219 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.02965f
C1220 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C1221 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.14207f
C1222 XThC.Tn[7] Iout 0.02244f
C1223 XThC.Tn[8] Vbias 0.31312f
C1224 XA.XIR[9].XIC[10].icell.PDM Vbias 0.03922f
C1225 XThC.XTB1.Y data[0] 0.06453f
C1226 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C1227 XA.XIR[15].XIC[3].icell.PUM VPWR 0.01079f
C1228 XA.XIR[0].XIC[2].icell.PDM Vbias 0.03922f
C1229 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07604f
C1230 XA.XIR[5].XIC[3].icell.Ien VPWR 0.21079f
C1231 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C1232 XThC.XTB3.Y a_8739_9569# 0.07285f
C1233 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C1234 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02601f
C1235 XThC.XTB6.Y XThC.Tn[7] 0.01474f
C1236 XA.XIR[9].XIC[8].icell.Ien Vbias 0.19151f
C1237 XA.XIR[4].XIC[6].icell.PUM VPWR 0.01079f
C1238 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1239 XThR.Tn[9] XThR.Tn[10] 0.11751f
C1240 XA.XIR[11].XIC[13].icell.PUM VPWR 0.01079f
C1241 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.14207f
C1242 XThC.Tn[5] XThR.Tn[1] 0.39128f
C1243 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.04627f
C1244 XA.XIR[10].XIC[11].icell.PDM VPWR 0.01373f
C1245 XThC.Tn[9] XThR.Tn[9] 0.39123f
C1246 XA.XIR[1].XIC_15.icell.PDM Vbias 0.03927f
C1247 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C1248 XA.XIR[9].XIC[11].icell.PDM VPWR 0.01373f
C1249 XThC.Tn[5] XThR.Tn[12] 0.39123f
C1250 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.04573f
C1251 XThC.Tn[14] XThR.Tn[8] 0.39123f
C1252 XA.XIR[13].XIC[12].icell.PDM VPWR 0.01373f
C1253 XA.XIR[0].XIC[3].icell.PDM VPWR 0.01334f
C1254 XA.XIR[4].XIC_15.icell.PDM Vbias 0.03927f
C1255 XA.XIR[7].XIC[4].icell.Ien Vbias 0.19151f
C1256 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C1257 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C1258 XThC.XTB6.Y a_5949_10571# 0.01283f
C1259 XA.XIR[9].XIC[9].icell.PUM VPWR 0.01079f
C1260 XThR.XTB3.Y a_n1049_7493# 0.23056f
C1261 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C1262 XThC.Tn[0] XThR.Tn[4] 0.39119f
C1263 XThC.XTBN.Y XThC.Tn[3] 0.48737f
C1264 XThR.XTBN.A VPWR 0.90745f
C1265 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C1266 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C1267 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C1268 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02601f
C1269 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.14207f
C1270 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02601f
C1271 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C1272 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.04573f
C1273 XThR.XTB5.Y a_n1049_6405# 0.24821f
C1274 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04035f
C1275 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04035f
C1276 XThR.Tn[6] VPWR 9.6234f
C1277 XA.XIR[11].XIC[14].icell.Ien VPWR 0.20455f
C1278 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C1279 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C1280 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1281 XThC.XTB4.Y XThC.Tn[7] 0.01805f
C1282 XA.XIR[6].XIC_15.icell.Ien VPWR 0.2801f
C1283 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01445f
C1284 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02601f
C1285 XThC.Tn[4] XThR.Tn[10] 0.39123f
C1286 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.14207f
C1287 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02601f
C1288 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C1289 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1290 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01768f
C1291 XA.XIR[7].XIC[5].icell.PUM VPWR 0.01079f
C1292 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.04261f
C1293 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C1294 XA.XIR[14].XIC[9].icell.Ien VPWR 0.21134f
C1295 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C1296 a_4861_9615# XThC.Tn[3] 0.26251f
C1297 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C1298 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.02965f
C1299 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.40895f
C1300 XA.XIR[5].XIC[0].icell.PDM Vbias 0.03915f
C1301 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.36378f
C1302 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.14207f
C1303 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C1304 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C1305 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C1306 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1307 XA.XIR[11].XIC[11].icell.PUM VPWR 0.01079f
C1308 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C1309 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04035f
C1310 XA.XIR[11].XIC[5].icell.PDM Vbias 0.03922f
C1311 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02602f
C1312 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04035f
C1313 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C1314 XA.XIR[10].XIC[9].icell.PDM Vbias 0.03922f
C1315 XA.XIR[5].XIC[1].icell.PDM VPWR 0.01373f
C1316 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02601f
C1317 XThC.Tn[2] XThR.Tn[14] 0.39123f
C1318 XA.XIR[5].XIC[9].icell.Ien Iout 0.06763f
C1319 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.04573f
C1320 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04035f
C1321 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02601f
C1322 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C1323 XThR.Tn[4] VPWR 9.6653f
C1324 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.04574f
C1325 XA.XIR[15].XIC[7].icell.Ien Vbias 0.15955f
C1326 XA.XIR[12].XIC[0].icell.PDM VPWR 0.01373f
C1327 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13586f
C1328 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C1329 a_n1049_7493# VPWR 0.7213f
C1330 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C1331 XA.XIR[11].XIC[6].icell.PDM VPWR 0.01373f
C1332 XA.XIR[11].XIC[12].icell.Ien VPWR 0.21079f
C1333 XA.XIR[4].XIC[10].icell.Ien Vbias 0.19151f
C1334 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C1335 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C1336 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02601f
C1337 XA.XIR[12].XIC[4].icell.Ien Iout 0.06763f
C1338 XA.XIR[10].XIC[10].icell.PDM VPWR 0.01373f
C1339 XA.XIR[0].XIC[1].icell.Ien Vbias 0.19186f
C1340 XA.XIR[2].XIC[1].icell.PDM Vbias 0.03922f
C1341 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.14207f
C1342 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C1343 XThR.XTB6.Y VPWR 1.05562f
C1344 XA.XIR[8].XIC[4].icell.Ien Vbias 0.19151f
C1345 XA.XIR[14].XIC[13].icell.PUM VPWR 0.01079f
C1346 XThC.Tn[13] VPWR 8.02161f
C1347 XA.XIR[13].XIC[11].icell.PDM VPWR 0.01373f
C1348 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.14207f
C1349 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C1350 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C1351 XA.XIR[15].XIC[8].icell.PUM VPWR 0.01079f
C1352 XA.XIR[5].XIC[8].icell.Ien VPWR 0.21079f
C1353 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.13345f
C1354 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.04573f
C1355 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C1356 XA.XIR[9].XIC[13].icell.Ien Vbias 0.19151f
C1357 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C1358 XA.XIR[4].XIC[11].icell.PUM VPWR 0.01079f
C1359 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C1360 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.04573f
C1361 XA.XIR[0].XIC[2].icell.PUM VPWR 0.01038f
C1362 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C1363 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02601f
C1364 XA.XIR[2].XIC[2].icell.PDM VPWR 0.01373f
C1365 XA.XIR[0].XIC[6].icell.Ien Vbias 0.19186f
C1366 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C1367 XA.XIR[8].XIC[5].icell.PUM VPWR 0.01079f
C1368 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02601f
C1369 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02601f
C1370 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C1371 XA.XIR[12].XIC[3].icell.Ien VPWR 0.21079f
C1372 XThC.Tn[6] Vbias 0.32012f
C1373 XA.XIR[14].XIC[14].icell.Ien VPWR 0.2051f
C1374 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02803f
C1375 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C1376 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04035f
C1377 XA.XIR[7].XIC[9].icell.Ien Vbias 0.19151f
C1378 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02601f
C1379 XThC.Tn[4] XThR.Tn[13] 0.39123f
C1380 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02601f
C1381 XA.XIR[9].XIC[14].icell.PUM VPWR 0.01079f
C1382 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C1383 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.14207f
C1384 XThC.XTB2.Y a_3773_9615# 0.2342f
C1385 XA.XIR[0].XIC[7].icell.PUM VPWR 0.01038f
C1386 XThR.Tn[7] Iout 1.10104f
C1387 XThC.Tn[7] XThR.Tn[9] 0.39123f
C1388 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C1389 XThC.Tn[3] XThR.Tn[8] 0.39123f
C1390 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0404f
C1391 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.04573f
C1392 XA.XIR[2].XIC[0].icell.Ien Vbias 0.19149f
C1393 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C1394 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.14207f
C1395 XA.XIR[4].XIC[2].icell.Ien Iout 0.06763f
C1396 XA.XIR[7].XIC[10].icell.PUM VPWR 0.01079f
C1397 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C1398 XA.XIR[11].XIC[10].icell.Ien VPWR 0.21079f
C1399 XA.XIR[7].XIC[1].icell.PDM Vbias 0.03922f
C1400 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04035f
C1401 XA.XIR[10].XIC[1].icell.Ien Vbias 0.19151f
C1402 XA.XIR[6].XIC[8].icell.PDM Vbias 0.03922f
C1403 XA.XIR[14].XIC[11].icell.PUM VPWR 0.01079f
C1404 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.14207f
C1405 XThC.XTBN.A VPWR 0.88816f
C1406 XA.XIR[5].XIC_15.icell.PDM Vbias 0.03927f
C1407 XA.XIR[14].XIC[5].icell.PDM Vbias 0.03922f
C1408 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.14207f
C1409 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C1410 XA.XIR[2].XIC[1].icell.PUM VPWR 0.01079f
C1411 XA.XIR[13].XIC[9].icell.PDM Vbias 0.03922f
C1412 XA.XIR[9].XIC[5].icell.Ien Iout 0.06763f
C1413 XA.XIR[11].XIC[0].icell.Ien VPWR 0.21079f
C1414 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C1415 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08254f
C1416 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02601f
C1417 XThC.Tn[5] XThC.Tn[6] 0.14628f
C1418 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04035f
C1419 XA.XIR[7].XIC[2].icell.PDM VPWR 0.01373f
C1420 XA.XIR[10].XIC[2].icell.PUM VPWR 0.01079f
C1421 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C1422 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.14207f
C1423 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.36378f
C1424 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13586f
C1425 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C1426 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01714f
C1427 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C1428 XA.XIR[6].XIC[9].icell.PDM VPWR 0.01373f
C1429 XA.XIR[11].XIC[13].icell.Ien Vbias 0.19151f
C1430 XA.XIR[14].XIC[6].icell.PDM VPWR 0.01373f
C1431 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C1432 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C1433 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1434 XA.XIR[5].XIC[14].icell.Ien Iout 0.06763f
C1435 XA.XIR[14].XIC[12].icell.Ien VPWR 0.21134f
C1436 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.04573f
C1437 XA.XIR[3].XIC[6].icell.Ien Vbias 0.19151f
C1438 XA.XIR[13].XIC[10].icell.PDM VPWR 0.01373f
C1439 XA.XIR[1].XIC[2].icell.PDM Vbias 0.03922f
C1440 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C1441 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02601f
C1442 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.04625f
C1443 XThC.XTB7.Y XThC.Tn[8] 0.07809f
C1444 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C1445 XA.XIR[4].XIC[2].icell.PDM Vbias 0.03922f
C1446 XA.XIR[9].XIC[4].icell.Ien VPWR 0.21079f
C1447 XThR.Tn[0] XThR.Tn[1] 0.26294f
C1448 XA.XIR[8].XIC[12].icell.PDM Vbias 0.03922f
C1449 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.04576f
C1450 XA.XIR[4].XIC_15.icell.Ien Vbias 0.19187f
C1451 XA.XIR[3].XIC[10].icell.PDM Vbias 0.03922f
C1452 XA.XIR[12].XIC[9].icell.Ien Iout 0.06763f
C1453 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C1454 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.1323f
C1455 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.14207f
C1456 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C1457 XA.XIR[8].XIC[9].icell.Ien Vbias 0.19151f
C1458 XA.XIR[3].XIC[7].icell.PUM VPWR 0.01079f
C1459 XA.XIR[1].XIC[3].icell.PDM VPWR 0.01373f
C1460 XA.XIR[9].XIC[0].icell.Ien Iout 0.06763f
C1461 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02601f
C1462 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.04573f
C1463 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C1464 XA.XIR[4].XIC[3].icell.PDM VPWR 0.01373f
C1465 XA.XIR[5].XIC[13].icell.Ien VPWR 0.21079f
C1466 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C1467 XThC.XTB3.Y VPWR 1.07064f
C1468 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02601f
C1469 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.0176f
C1470 XA.XIR[3].XIC[11].icell.PDM VPWR 0.01373f
C1471 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C1472 XThC.XTB1.Y XThC.Tn[0] 0.1842f
C1473 XA.XIR[8].XIC[13].icell.PDM VPWR 0.01373f
C1474 XThC.Tn[14] XThR.Tn[3] 0.39123f
C1475 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.04573f
C1476 XThC.XTBN.A a_9827_9569# 0.09118f
C1477 XThC.Tn[2] VPWR 7.06853f
C1478 XA.XIR[0].XIC[11].icell.Ien Vbias 0.19186f
C1479 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04035f
C1480 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04035f
C1481 XA.XIR[8].XIC[10].icell.PUM VPWR 0.01079f
C1482 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C1483 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07604f
C1484 XA.XIR[11].XIC_15.icell.Ien VPWR 0.2801f
C1485 XA.XIR[12].XIC[8].icell.Ien VPWR 0.21079f
C1486 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C1487 XThC.Tn[8] XThR.Tn[0] 0.39143f
C1488 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.36378f
C1489 XThC.Tn[10] XThR.Tn[5] 0.39123f
C1490 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C1491 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C1492 XA.XIR[7].XIC[14].icell.Ien Vbias 0.19151f
C1493 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C1494 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C1495 XA.XIR[11].XIC[11].icell.Ien Vbias 0.19151f
C1496 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.04573f
C1497 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.14207f
C1498 XA.XIR[14].XIC[10].icell.Ien VPWR 0.21134f
C1499 XThC.XTB5.Y a_5155_9615# 0.24821f
C1500 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C1501 XA.XIR[0].XIC[12].icell.PUM VPWR 0.01038f
C1502 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C1503 XA.XIR[13].XIC[1].icell.Ien Vbias 0.19151f
C1504 XThC.XTB7.A a_4067_9615# 0.0127f
C1505 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C1506 XA.XIR[15].XIC[4].icell.Ien Iout 0.07153f
C1507 XThC.XTBN.A XThC.XTB7.B 0.35142f
C1508 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04023f
C1509 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1510 XA.XIR[4].XIC[7].icell.Ien Iout 0.06763f
C1511 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.04573f
C1512 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01768f
C1513 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.14207f
C1514 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.04573f
C1515 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08285f
C1516 XA.XIR[4].XIC[1].icell.Ien VPWR 0.21079f
C1517 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C1518 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.04573f
C1519 XA.XIR[13].XIC[2].icell.PUM VPWR 0.01079f
C1520 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.14207f
C1521 XThC.XTBN.Y a_5155_9615# 0.07602f
C1522 XA.XIR[7].XIC[1].icell.Ien Iout 0.06763f
C1523 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.14207f
C1524 XA.XIR[14].XIC[13].icell.Ien Vbias 0.19151f
C1525 XA.XIR[9].XIC[10].icell.Ien Iout 0.06763f
C1526 XA.XIR[9].XIC[12].icell.PDM Vbias 0.03922f
C1527 XThC.XTB1.Y VPWR 1.11809f
C1528 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C1529 XA.XIR[12].XIC[14].icell.Ien Iout 0.06763f
C1530 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02601f
C1531 XA.XIR[15].XIC[3].icell.Ien VPWR 0.3396f
C1532 XA.XIR[0].XIC[4].icell.PDM Vbias 0.03922f
C1533 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C1534 XA.XIR[0].XIC[3].icell.Ien Iout 0.06712f
C1535 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.14207f
C1536 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02601f
C1537 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02601f
C1538 XA.XIR[1].XIC[1].icell.Ien Vbias 0.19162f
C1539 XThC.XTB7.A XThC.Tn[3] 0.0337f
C1540 XA.XIR[10].XIC[2].icell.Ien Vbias 0.19151f
C1541 XA.XIR[4].XIC[6].icell.Ien VPWR 0.21079f
C1542 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.14207f
C1543 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01244f
C1544 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C1545 XA.XIR[7].XIC[6].icell.Ien Iout 0.06763f
C1546 a_2979_9615# XThC.Tn[0] 0.27729f
C1547 XA.XIR[3].XIC[11].icell.Ien Vbias 0.19151f
C1548 XA.XIR[9].XIC[13].icell.PDM VPWR 0.01373f
C1549 XThC.Tn[12] XThR.Tn[6] 0.39123f
C1550 XA.XIR[0].XIC[5].icell.PDM VPWR 0.01462f
C1551 XA.XIR[7].XIC[0].icell.Ien VPWR 0.21079f
C1552 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.04573f
C1553 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C1554 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C1555 XA.XIR[2].XIC[4].icell.Ien Vbias 0.19151f
C1556 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C1557 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C1558 XA.XIR[1].XIC[2].icell.PUM VPWR 0.01079f
C1559 XA.XIR[9].XIC[9].icell.Ien VPWR 0.21079f
C1560 XA.XIR[10].XIC[3].icell.PUM VPWR 0.01079f
C1561 XA.XIR[1].XIC[6].icell.Ien Vbias 0.19162f
C1562 XThC.Tn[14] XThR.Tn[11] 0.39123f
C1563 XA.XIR[0].XIC[2].icell.Ien VPWR 0.21044f
C1564 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C1565 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.14207f
C1566 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C1567 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04035f
C1568 XThC.Tn[4] XThR.Tn[7] 0.39123f
C1569 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C1570 XA.XIR[11].XIC[14].icell.PDM VPWR 0.01349f
C1571 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04035f
C1572 XA.XIR[8].XIC[14].icell.Ien Vbias 0.19151f
C1573 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04035f
C1574 XA.XIR[3].XIC[12].icell.PUM VPWR 0.01079f
C1575 XThC.Tn[10] Iout 0.02225f
C1576 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02602f
C1577 XThC.XTB7.Y XThC.Tn[6] 0.2182f
C1578 XThC.XTB6.Y XThC.Tn[10] 0.02478f
C1579 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C1580 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07604f
C1581 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02601f
C1582 XA.XIR[14].XIC_15.icell.Ien VPWR 0.28041f
C1583 XA.XIR[7].XIC[5].icell.Ien VPWR 0.21079f
C1584 XA.XIR[2].XIC[5].icell.PUM VPWR 0.01079f
C1585 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.04573f
C1586 XA.XIR[1].XIC[7].icell.PUM VPWR 0.01079f
C1587 XThC.Tn[8] XThR.Tn[1] 0.39128f
C1588 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.14207f
C1589 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.14207f
C1590 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01768f
C1591 XA.XIR[14].XIC[11].icell.Ien Vbias 0.19151f
C1592 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C1593 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C1594 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02601f
C1595 XThC.Tn[8] XThR.Tn[12] 0.39123f
C1596 XA.XIR[5].XIC[2].icell.PDM Vbias 0.03922f
C1597 XA.XIR[12].XIC[12].icell.Ien Iout 0.06763f
C1598 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C1599 XA.XIR[6].XIC[1].icell.Ien Vbias 0.19151f
C1600 XThC.Tn[3] XThR.Tn[3] 0.39123f
C1601 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C1602 XA.XIR[12].XIC[1].icell.PDM Vbias 0.03922f
C1603 XThC.Tn[12] XThR.Tn[4] 0.39123f
C1604 XA.XIR[14].XIC[0].icell.PUM VPWR 0.01079f
C1605 XA.XIR[8].XIC[1].icell.Ien Iout 0.06763f
C1606 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04023f
C1607 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1608 XThR.Tn[2] Vbias 1.38579f
C1609 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.14207f
C1610 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.04573f
C1611 a_2979_9615# VPWR 0.70527f
C1612 XA.XIR[11].XIC[7].icell.PDM Vbias 0.03922f
C1613 XA.XIR[3].XIC[3].icell.Ien Iout 0.06763f
C1614 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.14207f
C1615 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.14207f
C1616 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.14207f
C1617 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04035f
C1618 XThC.XTB4.Y XThC.Tn[10] 0.01405f
C1619 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.04573f
C1620 XA.XIR[5].XIC[3].icell.PDM VPWR 0.01373f
C1621 XA.XIR[15].XIC[9].icell.Ien Iout 0.07153f
C1622 XThC.XTB4.Y a_4861_9615# 0.23756f
C1623 XThC.Tn[6] XThR.Tn[0] 0.3915f
C1624 XA.XIR[6].XIC[2].icell.PUM VPWR 0.01079f
C1625 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.04036f
C1626 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02601f
C1627 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C1628 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.14207f
C1629 XA.XIR[4].XIC[12].icell.Ien Iout 0.06763f
C1630 XA.XIR[6].XIC[6].icell.Ien Vbias 0.19151f
C1631 XThC.Tn[12] XThC.Tn[13] 0.17915f
C1632 XA.XIR[12].XIC[2].icell.PDM VPWR 0.01373f
C1633 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C1634 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02601f
C1635 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C1636 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.04573f
C1637 XA.XIR[8].XIC[6].icell.Ien Iout 0.06763f
C1638 XA.XIR[11].XIC[8].icell.PDM VPWR 0.01373f
C1639 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02602f
C1640 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02601f
C1641 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C1642 XA.XIR[2].XIC[3].icell.PDM Vbias 0.03922f
C1643 XA.XIR[13].XIC[2].icell.Ien Vbias 0.19151f
C1644 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.04575f
C1645 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04035f
C1646 XA.XIR[3].XIC[2].icell.Ien VPWR 0.21079f
C1647 XA.XIR[9].XIC_15.icell.Ien Iout 0.0694f
C1648 XA.XIR[6].XIC[7].icell.PUM VPWR 0.01079f
C1649 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.04573f
C1650 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C1651 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02601f
C1652 XA.XIR[15].XIC[8].icell.Ien VPWR 0.3396f
C1653 XA.XIR[11].XIC[5].icell.Ien Vbias 0.19151f
C1654 XA.XIR[0].XIC[8].icell.Ien Iout 0.06712f
C1655 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.14207f
C1656 XThC.XTBN.Y a_7875_9569# 0.229f
C1657 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.14207f
C1658 XA.XIR[10].XIC[7].icell.Ien Vbias 0.19151f
C1659 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C1660 XA.XIR[4].XIC[11].icell.Ien VPWR 0.21079f
C1661 XA.XIR[8].XIC[0].icell.PDM VPWR 0.01373f
C1662 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C1663 XThC.Tn[5] XThR.Tn[2] 0.39125f
C1664 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C1665 XA.XIR[12].XIC[10].icell.Ien Iout 0.06763f
C1666 XA.XIR[11].XIC[13].icell.PDM VPWR 0.01373f
C1667 XA.XIR[2].XIC[4].icell.PDM VPWR 0.01373f
C1668 XA.XIR[13].XIC[3].icell.PUM VPWR 0.01079f
C1669 XA.XIR[7].XIC[11].icell.Ien Iout 0.06763f
C1670 XA.XIR[8].XIC[5].icell.Ien VPWR 0.21079f
C1671 XThC.Tn[14] XThR.Tn[14] 0.39123f
C1672 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C1673 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.04573f
C1674 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C1675 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C1676 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C1677 XA.XIR[14].XIC[14].icell.PDM VPWR 0.01349f
C1678 XA.XIR[11].XIC[6].icell.PUM VPWR 0.01079f
C1679 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04035f
C1680 XA.XIR[2].XIC[9].icell.Ien Vbias 0.19151f
C1681 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C1682 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C1683 XThR.Tn[8] Iout 1.10104f
C1684 XA.XIR[9].XIC[14].icell.Ien VPWR 0.20455f
C1685 XA.XIR[3].XIC[0].icell.Ien Iout 0.06763f
C1686 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C1687 XA.XIR[10].XIC[8].icell.PUM VPWR 0.01079f
C1688 XA.XIR[1].XIC[11].icell.Ien Vbias 0.19162f
C1689 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02601f
C1690 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.14207f
C1691 XA.XIR[0].XIC[7].icell.Ien VPWR 0.21044f
C1692 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C1693 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C1694 XA.XIR[11].XIC[1].icell.Ien Iout 0.06763f
C1695 XThC.Tn[1] XThR.Tn[6] 0.39123f
C1696 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04035f
C1697 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.04261f
C1698 data[5] data[4] 0.64735f
C1699 XThC.XTBN.A XThC.Tn[12] 0.22871f
C1700 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.36378f
C1701 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C1702 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04035f
C1703 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02601f
C1704 XThR.Tn[5] a_n1049_5611# 0.27042f
C1705 XA.XIR[2].XIC[10].icell.PUM VPWR 0.01079f
C1706 XA.XIR[7].XIC[10].icell.Ien VPWR 0.21079f
C1707 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C1708 XThC.Tn[3] XThR.Tn[11] 0.39123f
C1709 XThR.XTB2.Y data[5] 0.017f
C1710 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.40895f
C1711 XA.XIR[1].XIC[12].icell.PUM VPWR 0.01079f
C1712 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04035f
C1713 XA.XIR[7].XIC[3].icell.PDM Vbias 0.03922f
C1714 XThR.Tn[10] Vbias 1.38583f
C1715 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.04573f
C1716 XA.XIR[15].XIC[14].icell.Ien Iout 0.07153f
C1717 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.04573f
C1718 XA.XIR[6].XIC[10].icell.PDM Vbias 0.03922f
C1719 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C1720 XA.XIR[15].XIC[1].icell.PDM Vbias 0.03922f
C1721 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C1722 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C1723 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.14207f
C1724 XThC.Tn[9] Vbias 0.31367f
C1725 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.04573f
C1726 XA.XIR[8].XIC[0].icell.Ien VPWR 0.21079f
C1727 XA.XIR[14].XIC[7].icell.PDM Vbias 0.03922f
C1728 XThC.XTB5.Y XThC.Tn[4] 0.20108f
C1729 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.04573f
C1730 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C1731 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.14207f
C1732 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04035f
C1733 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02601f
C1734 XA.XIR[7].XIC[4].icell.PDM VPWR 0.01373f
C1735 XThC.Tn[6] XThR.Tn[1] 0.39128f
C1736 XThC.Tn[10] XThR.Tn[9] 0.39123f
C1737 XThR.XTB6.A XThR.XTB7.A 0.44014f
C1738 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C1739 XA.XIR[3].XIC[8].icell.Ien Iout 0.06763f
C1740 XA.XIR[6].XIC[11].icell.PDM VPWR 0.01373f
C1741 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.14207f
C1742 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01714f
C1743 XThC.Tn[6] XThR.Tn[12] 0.39123f
C1744 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.14207f
C1745 XA.XIR[14].XIC[8].icell.PDM VPWR 0.01373f
C1746 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02601f
C1747 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C1748 XThR.XTB5.Y a_n997_1803# 0.06458f
C1749 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C1750 XThC.XTBN.Y XThC.Tn[4] 0.4886f
C1751 XA.XIR[1].XIC[4].icell.PDM Vbias 0.03922f
C1752 XA.XIR[6].XIC[11].icell.Ien Vbias 0.19151f
C1753 XA.XIR[1].XIC[3].icell.Ien Iout 0.06763f
C1754 XThC.Tn[1] XThR.Tn[4] 0.39123f
C1755 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.14207f
C1756 XA.XIR[9].XIC[0].icell.PDM VPWR 0.01373f
C1757 XA.XIR[12].XIC_15.icell.Ien Iout 0.0694f
C1758 XA.XIR[4].XIC[4].icell.PDM Vbias 0.03922f
C1759 XA.XIR[8].XIC[11].icell.Ien Iout 0.06763f
C1760 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08254f
C1761 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02601f
C1762 XA.XIR[8].XIC[14].icell.PDM Vbias 0.03922f
C1763 XA.XIR[3].XIC[12].icell.PDM Vbias 0.03922f
C1764 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.04573f
C1765 XThC.Tn[5] XThR.Tn[10] 0.39123f
C1766 XA.XIR[14].XIC[5].icell.Ien Vbias 0.19151f
C1767 XA.XIR[11].XIC[12].icell.PDM VPWR 0.01373f
C1768 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.04573f
C1769 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C1770 XA.XIR[13].XIC[7].icell.Ien Vbias 0.19151f
C1771 XA.XIR[3].XIC[7].icell.Ien VPWR 0.21079f
C1772 XA.XIR[1].XIC[5].icell.PDM VPWR 0.01373f
C1773 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C1774 XA.XIR[14].XIC[13].icell.PDM VPWR 0.01373f
C1775 XA.XIR[6].XIC[12].icell.PUM VPWR 0.01079f
C1776 XA.XIR[15].XIC[12].icell.Ien Iout 0.07153f
C1777 XA.XIR[0].XIC[13].icell.Ien Iout 0.06712f
C1778 XA.XIR[4].XIC[5].icell.PDM VPWR 0.01373f
C1779 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04035f
C1780 XA.XIR[3].XIC[13].icell.PDM VPWR 0.01373f
C1781 XA.XIR[1].XIC[2].icell.Ien VPWR 0.21079f
C1782 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07604f
C1783 XA.XIR[14].XIC[6].icell.PUM VPWR 0.01079f
C1784 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C1785 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.04574f
C1786 XA.XIR[13].XIC[8].icell.PUM VPWR 0.01079f
C1787 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04035f
C1788 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04035f
C1789 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C1790 XA.XIR[8].XIC[10].icell.Ien VPWR 0.21079f
C1791 XA.XIR[14].XIC[1].icell.Ien Iout 0.06763f
C1792 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01687f
C1793 XA.XIR[2].XIC[14].icell.Ien Vbias 0.19151f
C1794 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.36378f
C1795 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C1796 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C1797 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04035f
C1798 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02601f
C1799 XA.XIR[14].XIC[0].icell.Ien Vbias 0.19149f
C1800 XThC.Tn[3] XThR.Tn[14] 0.39123f
C1801 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13586f
C1802 XA.XIR[0].XIC[12].icell.Ien VPWR 0.21288f
C1803 XA.XIR[6].XIC[3].icell.Ien Iout 0.06763f
C1804 XThR.Tn[13] Vbias 1.38584f
C1805 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.04573f
C1806 XThC.XTB7.A a_5155_9615# 0.02287f
C1807 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C1808 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C1809 XThR.XTB5.A data[4] 0.14415f
C1810 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04039f
C1811 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01768f
C1812 XA.XIR[7].XIC_15.icell.Ien VPWR 0.2801f
C1813 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.14207f
C1814 XA.XIR[5].XIC[0].icell.Ien VPWR 0.21079f
C1815 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C1816 XThR.XTB7.B XThR.XTB6.A 1.47641f
C1817 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C1818 XA.XIR[5].XIC[4].icell.Ien Vbias 0.19151f
C1819 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C1820 XA.XIR[14].XIC[1].icell.PUM VPWR 0.01079f
C1821 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C1822 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.13138f
C1823 XThC.Tn[14] VPWR 7.97621f
C1824 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02601f
C1825 XThC.XTBN.Y a_6243_9615# 0.07767f
C1826 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.02965f
C1827 XA.XIR[2].XIC[1].icell.Ien Iout 0.06763f
C1828 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C1829 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C1830 XA.XIR[11].XIC[2].icell.Ien Iout 0.06763f
C1831 XA.XIR[15].XIC[10].icell.Ien Iout 0.07153f
C1832 XThR.Tn[8] XThR.Tn[9] 0.09761f
C1833 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C1834 XA.XIR[10].XIC[4].icell.Ien Iout 0.06763f
C1835 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08254f
C1836 XA.XIR[6].XIC[2].icell.Ien VPWR 0.21079f
C1837 XA.XIR[9].XIC[14].icell.PDM Vbias 0.03922f
C1838 XA.XIR[0].XIC[6].icell.PDM Vbias 0.03922f
C1839 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01459f
C1840 XA.XIR[5].XIC[5].icell.PUM VPWR 0.01079f
C1841 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C1842 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1843 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01244f
C1844 XA.XIR[3].XIC[13].icell.Ien Iout 0.06763f
C1845 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01544f
C1846 XA.XIR[11].XIC[11].icell.PDM VPWR 0.01373f
C1847 XThC.Tn[7] Vbias 0.33095f
C1848 VPWR data[6] 0.21222f
C1849 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.14207f
C1850 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C1851 XA.XIR[2].XIC[6].icell.Ien Iout 0.06763f
C1852 XA.XIR[14].XIC[12].icell.PDM VPWR 0.01373f
C1853 XThC.Tn[5] XThR.Tn[13] 0.39123f
C1854 XA.XIR[1].XIC[8].icell.Ien Iout 0.06763f
C1855 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07604f
C1856 XA.XIR[0].XIC[7].icell.PDM VPWR 0.01334f
C1857 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C1858 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C1859 XThC.Tn[4] XThR.Tn[8] 0.39123f
C1860 XA.XIR[10].XIC[3].icell.Ien VPWR 0.21079f
C1861 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C1862 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C1863 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C1864 bias[2] bias[0] 0.04602f
C1865 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04035f
C1866 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04023f
C1867 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04035f
C1868 XA.XIR[3].XIC[12].icell.Ien VPWR 0.21079f
C1869 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C1870 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C1871 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C1872 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C1873 XA.XIR[2].XIC[5].icell.Ien VPWR 0.21079f
C1874 XA.XIR[9].XIC[0].icell.PUM VPWR 0.01079f
C1875 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C1876 XA.XIR[1].XIC[7].icell.Ien VPWR 0.21079f
C1877 XThC.XTB6.Y a_5949_9615# 0.26831f
C1878 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.14207f
C1879 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.04628f
C1880 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C1881 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.03819f
C1882 a_3773_9615# Vbias 0.0139f
C1883 XThC.Tn[1] XThC.Tn[2] 0.71416f
C1884 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C1885 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02601f
C1886 XThR.Tn[3] Iout 1.10104f
C1887 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.14207f
C1888 XA.XIR[8].XIC_15.icell.Ien VPWR 0.2801f
C1889 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02602f
C1890 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02601f
C1891 XThR.XTB7.A a_n1049_5317# 0.02018f
C1892 XA.XIR[5].XIC[4].icell.PDM Vbias 0.03922f
C1893 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C1894 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C1895 XA.XIR[12].XIC[3].icell.PDM Vbias 0.03922f
C1896 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.02965f
C1897 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C1898 a_4067_9615# VPWR 0.70663f
C1899 XA.XIR[11].XIC[9].icell.PDM Vbias 0.03922f
C1900 a_n997_3755# XThR.Tn[9] 0.19352f
C1901 XThR.XTB2.Y XThR.Tn[9] 0.292f
C1902 XA.XIR[15].XIC_15.icell.Ien Iout 0.07331f
C1903 XA.XIR[6].XIC[8].icell.Ien Iout 0.06763f
C1904 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04035f
C1905 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.14207f
C1906 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C1907 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.14207f
C1908 XA.XIR[5].XIC[5].icell.PDM VPWR 0.01373f
C1909 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.04573f
C1910 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C1911 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.1155f
C1912 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02601f
C1913 XA.XIR[14].XIC[2].icell.Ien Iout 0.06763f
C1914 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C1915 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C1916 XA.XIR[12].XIC[4].icell.PDM VPWR 0.01373f
C1917 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C1918 XA.XIR[5].XIC[9].icell.Ien Vbias 0.19151f
C1919 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C1920 XA.XIR[13].XIC[4].icell.Ien Iout 0.06763f
C1921 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.04573f
C1922 XA.XIR[11].XIC[10].icell.PDM VPWR 0.01373f
C1923 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C1924 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C1925 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C1926 XA.XIR[8].XIC[1].icell.PDM Vbias 0.03922f
C1927 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C1928 XA.XIR[2].XIC[5].icell.PDM Vbias 0.03922f
C1929 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C1930 XA.XIR[11].XIC[7].icell.Ien Iout 0.06763f
C1931 XA.XIR[14].XIC[11].icell.PDM VPWR 0.01373f
C1932 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04035f
C1933 XA.XIR[10].XIC[9].icell.Ien Iout 0.06763f
C1934 XA.XIR[12].XIC[4].icell.Ien Vbias 0.19151f
C1935 XA.XIR[6].XIC[7].icell.Ien VPWR 0.21079f
C1936 XThC.XTB1.Y XThC.Tn[1] 0.01068f
C1937 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C1938 XThR.XTB7.A a_n1049_6405# 0.02287f
C1939 XThC.Tn[3] VPWR 7.02568f
C1940 XA.XIR[5].XIC[10].icell.PUM VPWR 0.01079f
C1941 XThC.XTBN.Y a_8963_9569# 0.22784f
C1942 XThC.XTB7.A data[1] 0.06544f
C1943 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02601f
C1944 XA.XIR[3].XIC[0].icell.PDM VPWR 0.01373f
C1945 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C1946 XA.XIR[8].XIC[2].icell.PDM VPWR 0.01373f
C1947 XA.XIR[12].XIC[14].icell.PUM VPWR 0.01079f
C1948 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C1949 XThC.Tn[9] XThR.Tn[0] 0.39143f
C1950 XA.XIR[2].XIC[6].icell.PDM VPWR 0.01373f
C1951 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13586f
C1952 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C1953 XThC.Tn[11] XThR.Tn[5] 0.39123f
C1954 XThR.Tn[1] XThR.Tn[2] 0.14437f
C1955 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.04573f
C1956 XA.XIR[13].XIC[3].icell.Ien VPWR 0.21079f
C1957 XA.XIR[2].XIC[11].icell.Ien Iout 0.06763f
C1958 XThR.XTB1.Y a_n997_3979# 0.06353f
C1959 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C1960 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.04574f
C1961 XA.XIR[12].XIC[5].icell.PUM VPWR 0.01079f
C1962 XA.XIR[1].XIC[13].icell.Ien Iout 0.06763f
C1963 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C1964 XA.XIR[11].XIC[6].icell.Ien VPWR 0.21079f
C1965 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.40907f
C1966 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04035f
C1967 XA.XIR[10].XIC[8].icell.Ien VPWR 0.21079f
C1968 XA.XIR[12].XIC[0].icell.Ien Iout 0.06763f
C1969 XThR.Tn[11] Iout 1.10104f
C1970 XThR.XTB7.B a_n1049_5317# 0.01743f
C1971 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02602f
C1972 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04035f
C1973 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C1974 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C1975 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04035f
C1976 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.14207f
C1977 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.03366f
C1978 XA.XIR[2].XIC[10].icell.Ien VPWR 0.21079f
C1979 XThR.Tn[7] Vbias 1.38578f
C1980 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C1981 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C1982 XThC.Tn[8] XThR.Tn[2] 0.39125f
C1983 XA.XIR[1].XIC[12].icell.Ien VPWR 0.21079f
C1984 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04035f
C1985 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.14207f
C1986 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C1987 XA.XIR[7].XIC[5].icell.PDM Vbias 0.03922f
C1988 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02792f
C1989 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C1990 XA.XIR[4].XIC[2].icell.Ien Vbias 0.19151f
C1991 XA.XIR[6].XIC[12].icell.PDM Vbias 0.03922f
C1992 XA.XIR[15].XIC[3].icell.PDM Vbias 0.03922f
C1993 XA.XIR[14].XIC[9].icell.PDM Vbias 0.03922f
C1994 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C1995 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.04573f
C1996 XThC.XTB5.A data[1] 0.11102f
C1997 XThC.XTB7.A XThC.Tn[4] 0.02779f
C1998 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C1999 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02601f
C2000 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.14207f
C2001 XA.XIR[9].XIC[1].icell.PDM Vbias 0.03922f
C2002 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04035f
C2003 XA.XIR[12].XIC[12].icell.PUM VPWR 0.01079f
C2004 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.36378f
C2005 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C2006 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C2007 XA.XIR[7].XIC[6].icell.PDM VPWR 0.01373f
C2008 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C2009 XA.XIR[9].XIC[5].icell.Ien Vbias 0.19151f
C2010 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C2011 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01714f
C2012 XA.XIR[4].XIC[3].icell.PUM VPWR 0.01079f
C2013 XA.XIR[6].XIC[13].icell.PDM VPWR 0.01373f
C2014 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C2015 XA.XIR[6].XIC[13].icell.Ien Iout 0.06763f
C2016 XA.XIR[10].XIC[14].icell.Ien Iout 0.06763f
C2017 XThC.Tn[13] XThR.Tn[6] 0.39123f
C2018 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.04573f
C2019 VPWR data[2] 0.21031f
C2020 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C2021 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.14207f
C2022 XA.XIR[14].XIC[10].icell.PDM VPWR 0.01373f
C2023 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C2024 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C2025 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02601f
C2026 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C2027 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C2028 XA.XIR[1].XIC[6].icell.PDM Vbias 0.03922f
C2029 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01244f
C2030 VPWR bias[0] 2.91967f
C2031 XA.XIR[9].XIC[2].icell.PDM VPWR 0.01373f
C2032 XA.XIR[14].XIC[7].icell.Ien Iout 0.06763f
C2033 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C2034 XA.XIR[4].XIC[6].icell.PDM Vbias 0.03922f
C2035 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.04573f
C2036 XThC.Tn[5] XThR.Tn[7] 0.39123f
C2037 XA.XIR[5].XIC[14].icell.Ien Vbias 0.19151f
C2038 XA.XIR[13].XIC[9].icell.Ien Iout 0.06763f
C2039 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08254f
C2040 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C2041 XThC.Tn[11] Iout 0.02285f
C2042 XA.XIR[9].XIC[6].icell.PUM VPWR 0.01079f
C2043 XA.XIR[12].XIC[13].icell.Ien VPWR 0.21079f
C2044 XA.XIR[3].XIC[14].icell.PDM Vbias 0.03922f
C2045 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02601f
C2046 XThC.XTB7.Y XThC.Tn[7] 0.08399f
C2047 XThC.XTB6.Y XThC.Tn[11] 0.02473f
C2048 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04035f
C2049 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C2050 XA.XIR[1].XIC[7].icell.PDM VPWR 0.01373f
C2051 XA.XIR[6].XIC[12].icell.Ien VPWR 0.21079f
C2052 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C2053 XA.XIR[12].XIC[9].icell.Ien Vbias 0.19151f
C2054 XThC.Tn[9] XThR.Tn[1] 0.39128f
C2055 data[1] data[0] 0.64735f
C2056 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01768f
C2057 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C2058 XA.XIR[4].XIC[7].icell.PDM VPWR 0.01373f
C2059 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04035f
C2060 XThC.Tn[9] XThR.Tn[12] 0.39123f
C2061 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07604f
C2062 XA.XIR[9].XIC[0].icell.Ien Vbias 0.19149f
C2063 XA.XIR[14].XIC[6].icell.Ien VPWR 0.21134f
C2064 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.04573f
C2065 XThR.XTBN.Y a_n1049_5317# 0.07731f
C2066 XA.XIR[13].XIC[8].icell.Ien VPWR 0.21079f
C2067 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04035f
C2068 XThC.Tn[4] XThR.Tn[3] 0.39123f
C2069 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.04629f
C2070 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C2071 XA.XIR[5].XIC[1].icell.Ien Iout 0.06763f
C2072 XA.XIR[12].XIC[10].icell.PUM VPWR 0.01079f
C2073 XThC.Tn[13] XThR.Tn[4] 0.39123f
C2074 XThR.Tn[14] Iout 1.10103f
C2075 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.04261f
C2076 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C2077 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C2078 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.04575f
C2079 XThC.XTB4.Y XThC.Tn[11] 0.30457f
C2080 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C2081 XThC.Tn[8] XThR.Tn[10] 0.39123f
C2082 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C2083 XThC.Tn[0] XThR.Tn[5] 0.39119f
C2084 XA.XIR[10].XIC[12].icell.Ien Iout 0.06763f
C2085 XA.XIR[9].XIC[1].icell.PUM VPWR 0.01079f
C2086 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04035f
C2087 XThC.Tn[7] XThR.Tn[0] 0.39143f
C2088 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C2089 XThC.Tn[8] XThC.Tn[9] 0.0619f
C2090 XA.XIR[3].XIC[0].icell.PUM VPWR 0.01079f
C2091 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C2092 XA.XIR[10].XIC[0].icell.PDM Vbias 0.03915f
C2093 XThC.XTB7.A a_6243_9615# 0.02018f
C2094 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.36378f
C2095 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.04573f
C2096 XA.XIR[5].XIC[6].icell.Ien Iout 0.06763f
C2097 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04035f
C2098 XA.XIR[2].XIC_15.icell.Ien VPWR 0.2801f
C2099 XA.XIR[12].XIC[11].icell.Ien VPWR 0.21079f
C2100 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C2101 XA.XIR[15].XIC[4].icell.Ien Vbias 0.15955f
C2102 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.14207f
C2103 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.04573f
C2104 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02601f
C2105 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C2106 XA.XIR[4].XIC[7].icell.Ien Vbias 0.19151f
C2107 XA.XIR[10].XIC[1].icell.PDM VPWR 0.01373f
C2108 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.02965f
C2109 XA.XIR[15].XIC[14].icell.PUM VPWR 0.01079f
C2110 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.04573f
C2111 XThR.Tn[12] a_n997_1803# 0.18719f
C2112 XThR.XTBN.Y a_n1049_6405# 0.07602f
C2113 XThC.XTB7.B data[2] 0.07481f
C2114 XA.XIR[13].XIC[14].icell.Ien Iout 0.06763f
C2115 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.14207f
C2116 XThC.Tn[6] XThR.Tn[2] 0.39125f
C2117 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02601f
C2118 XA.XIR[7].XIC[1].icell.Ien Vbias 0.19151f
C2119 XA.XIR[0].XIC[8].icell.PDM Vbias 0.03922f
C2120 XA.XIR[15].XIC[5].icell.PUM VPWR 0.01079f
C2121 XA.XIR[5].XIC[5].icell.Ien VPWR 0.21079f
C2122 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.1155f
C2123 XThC.XTB5.Y Vbias 0.01606f
C2124 XA.XIR[9].XIC[10].icell.Ien Vbias 0.19151f
C2125 XA.XIR[4].XIC[8].icell.PUM VPWR 0.01079f
C2126 XA.XIR[12].XIC[14].icell.Ien Vbias 0.19151f
C2127 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C2128 XA.XIR[0].XIC[3].icell.Ien Vbias 0.19186f
C2129 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.04573f
C2130 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02601f
C2131 XThR.XTB4.Y a_n1049_6405# 0.01546f
C2132 XThR.Tn[5] VPWR 9.66314f
C2133 XA.XIR[10].XIC[10].icell.Ien Iout 0.06763f
C2134 XA.XIR[7].XIC[2].icell.PUM VPWR 0.01079f
C2135 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.04573f
C2136 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.14207f
C2137 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01653f
C2138 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C2139 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C2140 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C2141 XA.XIR[7].XIC[6].icell.Ien Vbias 0.19151f
C2142 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02601f
C2143 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.04573f
C2144 XThC.Tn[2] XThR.Tn[6] 0.39123f
C2145 XA.XIR[9].XIC[11].icell.PUM VPWR 0.01079f
C2146 XThR.Tn[12] XThR.Tn[13] 0.1027f
C2147 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C2148 XThC.XTBN.Y Vbias 0.16653f
C2149 XA.XIR[0].XIC[4].icell.PUM VPWR 0.01038f
C2150 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04035f
C2151 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C2152 XThC.Tn[4] XThR.Tn[11] 0.39123f
C2153 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04035f
C2154 VPWR data[5] 0.44032f
C2155 XThC.Tn[0] Iout 0.02199f
C2156 XA.XIR[7].XIC[7].icell.PUM VPWR 0.01079f
C2157 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02601f
C2158 XThC.Tn[10] Vbias 0.32711f
C2159 XA.XIR[15].XIC[12].icell.PUM VPWR 0.01079f
C2160 XThC.XTB5.Y XThC.Tn[5] 0.01168f
C2161 a_10915_9569# XThC.Tn[14] 0.20879f
C2162 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.40991f
C2163 XThC.Tn[8] XThR.Tn[13] 0.39123f
C2164 XA.XIR[13].XIC[12].icell.Ien Iout 0.06763f
C2165 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.03823f
C2166 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.03366f
C2167 XA.XIR[5].XIC[6].icell.PDM Vbias 0.03922f
C2168 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.14207f
C2169 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C2170 XThC.Tn[7] XThR.Tn[1] 0.39128f
C2171 XThC.Tn[11] XThR.Tn[9] 0.39123f
C2172 XA.XIR[9].XIC[2].icell.Ien Iout 0.06763f
C2173 XA.XIR[13].XIC[0].icell.PDM Vbias 0.03915f
C2174 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C2175 XThC.Tn[7] XThR.Tn[12] 0.39123f
C2176 XA.XIR[12].XIC[5].icell.PDM Vbias 0.03922f
C2177 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02602f
C2178 XA.XIR[12].XIC[12].icell.Ien Vbias 0.19151f
C2179 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02601f
C2180 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04023f
C2181 a_5155_9615# VPWR 0.7051f
C2182 XA.XIR[6].XIC[0].icell.PDM VPWR 0.01373f
C2183 XThC.Tn[2] XThR.Tn[4] 0.39123f
C2184 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02601f
C2185 XThC.XTBN.Y XThC.Tn[5] 0.4867f
C2186 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04035f
C2187 XA.XIR[15].XIC[13].icell.Ien VPWR 0.3396f
C2188 XA.XIR[5].XIC[7].icell.PDM VPWR 0.01373f
C2189 XA.XIR[8].XIC[1].icell.Ien Vbias 0.19151f
C2190 XA.XIR[5].XIC[11].icell.Ien Iout 0.06763f
C2191 XA.XIR[3].XIC[3].icell.Ien Vbias 0.19151f
C2192 XA.XIR[13].XIC[1].icell.PDM VPWR 0.01373f
C2193 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C2194 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.04573f
C2195 XThR.XTB7.B XThR.XTB7.A 0.35833f
C2196 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C2197 XThC.Tn[6] XThR.Tn[10] 0.39123f
C2198 XA.XIR[15].XIC[9].icell.Ien Vbias 0.15955f
C2199 XA.XIR[12].XIC[6].icell.PDM VPWR 0.01373f
C2200 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02601f
C2201 XThC.Tn[7] XThC.Tn[8] 0.06603f
C2202 XA.XIR[3].XIC[1].icell.PDM Vbias 0.03922f
C2203 XA.XIR[4].XIC[12].icell.Ien Vbias 0.19151f
C2204 XA.XIR[12].XIC[6].icell.Ien Iout 0.06763f
C2205 XA.XIR[8].XIC[3].icell.PDM Vbias 0.03922f
C2206 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.04573f
C2207 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C2208 XA.XIR[2].XIC[7].icell.PDM Vbias 0.03922f
C2209 XA.XIR[10].XIC_15.icell.Ien Iout 0.0694f
C2210 XA.XIR[8].XIC[2].icell.PUM VPWR 0.01079f
C2211 VPWR Iout 66.3711f
C2212 XA.XIR[8].XIC[6].icell.Ien Vbias 0.19151f
C2213 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04035f
C2214 XA.XIR[3].XIC[4].icell.PUM VPWR 0.01079f
C2215 XThC.XTB6.Y VPWR 1.03166f
C2216 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C2217 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.13138f
C2218 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C2219 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02602f
C2220 XA.XIR[15].XIC[10].icell.PUM VPWR 0.01079f
C2221 XA.XIR[5].XIC[10].icell.Ien VPWR 0.21079f
C2222 XThC.XTBN.Y a_10051_9569# 0.23006f
C2223 XA.XIR[13].XIC[10].icell.Ien Iout 0.06763f
C2224 XThR.XTB7.A XThR.Tn[2] 0.12549f
C2225 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C2226 XA.XIR[9].XIC_15.icell.Ien Vbias 0.19187f
C2227 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C2228 XA.XIR[4].XIC[13].icell.PUM VPWR 0.01079f
C2229 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02601f
C2230 XA.XIR[3].XIC[2].icell.PDM VPWR 0.01373f
C2231 XA.XIR[8].XIC[4].icell.PDM VPWR 0.01373f
C2232 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.14207f
C2233 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.14207f
C2234 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02601f
C2235 XA.XIR[2].XIC[8].icell.PDM VPWR 0.01373f
C2236 XA.XIR[0].XIC[8].icell.Ien Vbias 0.19186f
C2237 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.14207f
C2238 XA.XIR[8].XIC[7].icell.PUM VPWR 0.01079f
C2239 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.0279f
C2240 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C2241 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C2242 XA.XIR[12].XIC[5].icell.Ien VPWR 0.21079f
C2243 XThC.Tn[4] XThR.Tn[14] 0.39123f
C2244 XA.XIR[12].XIC[10].icell.Ien Vbias 0.19151f
C2245 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.04573f
C2246 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C2247 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04035f
C2248 XA.XIR[7].XIC[11].icell.Ien Vbias 0.19151f
C2249 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02601f
C2250 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.0176f
C2251 XA.XIR[15].XIC[11].icell.Ien VPWR 0.3396f
C2252 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.14207f
C2253 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02601f
C2254 XThC.XTB4.Y VPWR 0.91479f
C2255 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C2256 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.04575f
C2257 XA.XIR[0].XIC[9].icell.PUM VPWR 0.01038f
C2258 XA.XIR[3].XIC[0].icell.Ien Vbias 0.19149f
C2259 XThR.Tn[8] Vbias 1.38578f
C2260 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04035f
C2261 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C2262 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C2263 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04035f
C2264 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C2265 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.03916f
C2266 XA.XIR[7].XIC[12].icell.PUM VPWR 0.01079f
C2267 XA.XIR[4].XIC[4].icell.Ien Iout 0.06763f
C2268 XThR.XTB5.A VPWR 0.83253f
C2269 XA.XIR[11].XIC[1].icell.Ien Vbias 0.19151f
C2270 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.04036f
C2271 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C2272 XA.XIR[7].XIC[7].icell.PDM Vbias 0.03922f
C2273 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04035f
C2274 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08254f
C2275 XA.XIR[6].XIC[14].icell.PDM Vbias 0.03922f
C2276 XA.XIR[15].XIC[5].icell.PDM Vbias 0.03922f
C2277 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C2278 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02601f
C2279 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.14207f
C2280 XA.XIR[3].XIC[1].icell.PUM VPWR 0.01079f
C2281 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02601f
C2282 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.14207f
C2283 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02601f
C2284 XA.XIR[15].XIC[14].icell.Ien Vbias 0.15955f
C2285 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C2286 XA.XIR[9].XIC[7].icell.Ien Iout 0.06763f
C2287 XA.XIR[11].XIC[2].icell.PUM VPWR 0.01079f
C2288 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C2289 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04035f
C2290 XA.XIR[9].XIC[3].icell.PDM Vbias 0.03922f
C2291 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.36378f
C2292 XA.XIR[7].XIC[8].icell.PDM VPWR 0.01373f
C2293 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.04573f
C2294 XA.XIR[9].XIC[1].icell.Ien VPWR 0.21079f
C2295 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.14207f
C2296 XThC.Tn[6] XThR.Tn[13] 0.39123f
C2297 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01714f
C2298 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07604f
C2299 XA.XIR[4].XIC[3].icell.Ien VPWR 0.21079f
C2300 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.04261f
C2301 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C2302 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C2303 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C2304 XThC.Tn[0] XThR.Tn[9] 0.39118f
C2305 XA.XIR[7].XIC[3].icell.Ien Iout 0.06763f
C2306 XA.XIR[3].XIC[8].icell.Ien Vbias 0.19151f
C2307 XThC.Tn[5] XThR.Tn[8] 0.39123f
C2308 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C2309 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C2310 XA.XIR[1].XIC[8].icell.PDM Vbias 0.03922f
C2311 XA.XIR[13].XIC_15.icell.Ien Iout 0.0694f
C2312 XA.XIR[9].XIC[4].icell.PDM VPWR 0.01373f
C2313 XThC.XTB2.Y VPWR 0.97672f
C2314 XA.XIR[4].XIC[8].icell.PDM Vbias 0.03922f
C2315 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.04573f
C2316 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.04574f
C2317 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C2318 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C2319 XA.XIR[9].XIC[6].icell.Ien VPWR 0.21079f
C2320 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.13138f
C2321 XA.XIR[1].XIC[3].icell.Ien Vbias 0.19162f
C2322 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.04261f
C2323 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.14207f
C2324 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C2325 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C2326 XA.XIR[12].XIC_15.icell.Ien Vbias 0.19187f
C2327 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02601f
C2328 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04035f
C2329 XA.XIR[8].XIC[11].icell.Ien Vbias 0.19151f
C2330 XA.XIR[3].XIC[9].icell.PUM VPWR 0.01079f
C2331 XA.XIR[1].XIC[9].icell.PDM VPWR 0.01373f
C2332 XThC.XTB3.Y XThC.Tn[2] 0.18399f
C2333 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02803f
C2334 VPWR data[1] 0.44103f
C2335 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C2336 XA.XIR[7].XIC[2].icell.Ien VPWR 0.21079f
C2337 XA.XIR[4].XIC[9].icell.PDM VPWR 0.01373f
C2338 XA.XIR[5].XIC_15.icell.Ien VPWR 0.2801f
C2339 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02601f
C2340 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C2341 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04035f
C2342 XThC.Tn[6] XThC.Tn[7] 0.09739f
C2343 XA.XIR[1].XIC[4].icell.PUM VPWR 0.01079f
C2344 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C2345 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C2346 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07604f
C2347 XA.XIR[15].XIC[12].icell.Ien Vbias 0.15955f
C2348 XA.XIR[0].XIC[13].icell.Ien Vbias 0.19186f
C2349 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02601f
C2350 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.0176f
C2351 XThR.XTB1.Y data[4] 0.06453f
C2352 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C2353 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04035f
C2354 XA.XIR[8].XIC[12].icell.PUM VPWR 0.01079f
C2355 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C2356 XA.XIR[15].XIC[1].icell.Ien Iout 0.07153f
C2357 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.02965f
C2358 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C2359 XThC.Tn[8] XThR.Tn[7] 0.39123f
C2360 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04035f
C2361 XThC.XTB7.Y XThC.Tn[10] 0.07427f
C2362 XThR.Tn[9] VPWR 10.6021f
C2363 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C2364 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04035f
C2365 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.1155f
C2366 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C2367 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.14207f
C2368 XA.XIR[14].XIC[1].icell.Ien Vbias 0.19151f
C2369 XA.XIR[0].XIC[14].icell.PUM VPWR 0.01038f
C2370 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.14207f
C2371 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.14207f
C2372 XA.XIR[10].XIC[2].icell.PDM Vbias 0.03922f
C2373 XA.XIR[15].XIC[6].icell.Ien Iout 0.07153f
C2374 XA.XIR[12].XIC[0].icell.PUM VPWR 0.01079f
C2375 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C2376 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04035f
C2377 XA.XIR[4].XIC[9].icell.Ien Iout 0.06763f
C2378 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04023f
C2379 XA.XIR[6].XIC[3].icell.Ien Vbias 0.19151f
C2380 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.14207f
C2381 XA.XIR[15].XIC[0].icell.Ien VPWR 0.3396f
C2382 XA.XIR[0].XIC[0].icell.Ien Iout 0.06712f
C2383 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.04573f
C2384 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C2385 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C2386 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C2387 XA.XIR[14].XIC[2].icell.PUM VPWR 0.01079f
C2388 XA.XIR[8].XIC[3].icell.Ien Iout 0.06763f
C2389 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02601f
C2390 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.14207f
C2391 XA.XIR[10].XIC[3].icell.PDM VPWR 0.01373f
C2392 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C2393 XThC.Tn[4] VPWR 7.06697f
C2394 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.14207f
C2395 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C2396 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C2397 XA.XIR[9].XIC[12].icell.Ien Iout 0.06763f
C2398 XA.XIR[6].XIC[4].icell.PUM VPWR 0.01079f
C2399 XThR.XTBN.Y XThR.Tn[2] 0.61889f
C2400 XA.XIR[2].XIC[1].icell.Ien Vbias 0.19151f
C2401 XThC.Tn[10] XThR.Tn[0] 0.39146f
C2402 XA.XIR[15].XIC[5].icell.Ien VPWR 0.3396f
C2403 XA.XIR[0].XIC[10].icell.PDM Vbias 0.03922f
C2404 XThC.Tn[12] XThR.Tn[5] 0.39123f
C2405 XA.XIR[0].XIC[5].icell.Ien Iout 0.06712f
C2406 XA.XIR[11].XIC[2].icell.Ien Vbias 0.19151f
C2407 XA.XIR[15].XIC[10].icell.Ien Vbias 0.15955f
C2408 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.14207f
C2409 XThR.XTB7.B XThR.Tn[10] 0.06102f
C2410 XThC.XTB7.B a_7875_9569# 0.01174f
C2411 XThC.XTB7.A Vbias 0.0148f
C2412 XA.XIR[4].XIC[8].icell.Ien VPWR 0.21079f
C2413 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C2414 XA.XIR[10].XIC[4].icell.Ien Vbias 0.19151f
C2415 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C2416 a_8963_9569# XThC.Tn[11] 0.1927f
C2417 XA.XIR[8].XIC[2].icell.Ien VPWR 0.21079f
C2418 XA.XIR[7].XIC[8].icell.Ien Iout 0.06763f
C2419 XA.XIR[3].XIC[13].icell.Ien Vbias 0.19151f
C2420 XA.XIR[10].XIC[14].icell.PUM VPWR 0.01079f
C2421 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C2422 XA.XIR[2].XIC[2].icell.PUM VPWR 0.01079f
C2423 XA.XIR[0].XIC[11].icell.PDM VPWR 0.01334f
C2424 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.14207f
C2425 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.04627f
C2426 XA.XIR[11].XIC[3].icell.PUM VPWR 0.01079f
C2427 XA.XIR[2].XIC[6].icell.Ien Vbias 0.19151f
C2428 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C2429 XA.XIR[9].XIC[11].icell.Ien VPWR 0.21079f
C2430 XA.XIR[10].XIC[5].icell.PUM VPWR 0.01079f
C2431 XA.XIR[1].XIC[8].icell.Ien Vbias 0.19162f
C2432 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C2433 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C2434 XA.XIR[12].XIC[14].icell.PDM VPWR 0.01349f
C2435 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02602f
C2436 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.14207f
C2437 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C2438 XA.XIR[0].XIC[4].icell.Ien VPWR 0.21056f
C2439 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04035f
C2440 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04035f
C2441 XThC.Tn[9] XThR.Tn[2] 0.39125f
C2442 XA.XIR[3].XIC[14].icell.PUM VPWR 0.01079f
C2443 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02601f
C2444 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C2445 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07945f
C2446 XA.XIR[10].XIC[0].icell.Ien Iout 0.06763f
C2447 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C2448 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.04573f
C2449 XA.XIR[7].XIC[7].icell.Ien VPWR 0.21079f
C2450 XA.XIR[2].XIC[7].icell.PUM VPWR 0.01079f
C2451 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04035f
C2452 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C2453 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01256f
C2454 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C2455 XA.XIR[1].XIC[9].icell.PUM VPWR 0.01079f
C2456 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C2457 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02601f
C2458 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C2459 XA.XIR[6].XIC[1].icell.PDM Vbias 0.03922f
C2460 XThC.XTB7.A XThC.Tn[5] 0.02777f
C2461 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.40914f
C2462 XA.XIR[5].XIC[8].icell.PDM Vbias 0.03922f
C2463 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C2464 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C2465 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.04036f
C2466 XA.XIR[13].XIC[2].icell.PDM Vbias 0.03922f
C2467 XThR.Tn[3] Vbias 1.38579f
C2468 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.14207f
C2469 XThC.Tn[14] XThR.Tn[6] 0.39123f
C2470 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.04573f
C2471 XA.XIR[12].XIC[7].icell.PDM Vbias 0.03922f
C2472 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.14207f
C2473 a_6243_9615# VPWR 0.7055f
C2474 XA.XIR[3].XIC[5].icell.Ien Iout 0.06763f
C2475 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.02965f
C2476 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.14207f
C2477 XA.XIR[6].XIC[2].icell.PDM VPWR 0.01373f
C2478 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.04573f
C2479 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04035f
C2480 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.14207f
C2481 XA.XIR[10].XIC[12].icell.PUM VPWR 0.01079f
C2482 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C2483 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C2484 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02601f
C2485 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.14207f
C2486 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C2487 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02601f
C2488 XA.XIR[5].XIC[9].icell.PDM VPWR 0.01373f
C2489 XThC.Tn[6] XThR.Tn[7] 0.39123f
C2490 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C2491 XA.XIR[15].XIC_15.icell.Ien Vbias 0.15958f
C2492 XThC.Tn[12] Iout 0.02212f
C2493 XA.XIR[13].XIC[3].icell.PDM VPWR 0.01373f
C2494 XA.XIR[4].XIC[14].icell.Ien Iout 0.06763f
C2495 XA.XIR[6].XIC[8].icell.Ien Vbias 0.19151f
C2496 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.14207f
C2497 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.02805f
C2498 XThR.XTBN.Y XThR.Tn[10] 0.46534f
C2499 XThC.XTB5.Y XThC.Tn[8] 0.0173f
C2500 XA.XIR[12].XIC[8].icell.PDM VPWR 0.01373f
C2501 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C2502 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02601f
C2503 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C2504 XThC.XTB6.Y XThC.Tn[12] 0.0253f
C2505 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C2506 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C2507 XA.XIR[8].XIC[8].icell.Ien Iout 0.06763f
C2508 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.04573f
C2509 XA.XIR[8].XIC[5].icell.PDM Vbias 0.03922f
C2510 XA.XIR[3].XIC[3].icell.PDM Vbias 0.03922f
C2511 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C2512 XA.XIR[14].XIC[2].icell.Ien Vbias 0.19151f
C2513 XThC.Tn[10] XThR.Tn[1] 0.39128f
C2514 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.04574f
C2515 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02601f
C2516 a_5949_9615# XThC.Tn[5] 0.26251f
C2517 XA.XIR[2].XIC[9].icell.PDM Vbias 0.03922f
C2518 XA.XIR[13].XIC[4].icell.Ien Vbias 0.19151f
C2519 XA.XIR[10].XIC[13].icell.Ien VPWR 0.21079f
C2520 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04035f
C2521 XA.XIR[3].XIC[4].icell.Ien VPWR 0.21079f
C2522 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.0176f
C2523 XThC.Tn[10] XThR.Tn[12] 0.39123f
C2524 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C2525 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02601f
C2526 XA.XIR[6].XIC[9].icell.PUM VPWR 0.01079f
C2527 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C2528 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C2529 XA.XIR[0].XIC[10].icell.Ien Iout 0.06712f
C2530 XA.XIR[11].XIC[7].icell.Ien Vbias 0.19151f
C2531 XA.XIR[13].XIC[14].icell.PUM VPWR 0.01079f
C2532 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.14207f
C2533 XThC.XTBN.Y XThC.Tn[8] 0.40735f
C2534 XThC.Tn[5] XThR.Tn[3] 0.39123f
C2535 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C2536 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C2537 XA.XIR[4].XIC[13].icell.Ien VPWR 0.21079f
C2538 XA.XIR[10].XIC[9].icell.Ien Vbias 0.19151f
C2539 XA.XIR[8].XIC[6].icell.PDM VPWR 0.01373f
C2540 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.03888f
C2541 XThC.XTB1.Y a_2979_9615# 0.21263f
C2542 XA.XIR[3].XIC[4].icell.PDM VPWR 0.01373f
C2543 XA.XIR[12].XIC[13].icell.PDM VPWR 0.01373f
C2544 XThC.Tn[14] XThR.Tn[4] 0.39123f
C2545 XA.XIR[14].XIC[3].icell.PUM VPWR 0.01079f
C2546 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.03823f
C2547 XA.XIR[2].XIC[10].icell.PDM VPWR 0.01373f
C2548 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C2549 XA.XIR[13].XIC[5].icell.PUM VPWR 0.01079f
C2550 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04035f
C2551 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02602f
C2552 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C2553 XA.XIR[7].XIC[13].icell.Ien Iout 0.06763f
C2554 XA.XIR[8].XIC[7].icell.Ien VPWR 0.21079f
C2555 XA.XIR[15].XIC[14].icell.PDM VPWR 0.0169f
C2556 XThC.Tn[9] XThR.Tn[10] 0.39123f
C2557 XThC.Tn[1] XThR.Tn[5] 0.39123f
C2558 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C2559 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02601f
C2560 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.14207f
C2561 XA.XIR[11].XIC[8].icell.PUM VPWR 0.01079f
C2562 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C2563 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C2564 XA.XIR[2].XIC[11].icell.Ien Vbias 0.19151f
C2565 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02601f
C2566 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04035f
C2567 XA.XIR[13].XIC[0].icell.Ien Iout 0.06763f
C2568 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.36378f
C2569 XA.XIR[10].XIC[10].icell.PUM VPWR 0.01079f
C2570 XThC.Tn[13] XThC.Tn[14] 0.3543f
C2571 XA.XIR[1].XIC[13].icell.Ien Vbias 0.19162f
C2572 XA.XIR[0].XIC[9].icell.Ien VPWR 0.21193f
C2573 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.14207f
C2574 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01687f
C2575 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02601f
C2576 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C2577 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04035f
C2578 XA.XIR[12].XIC[0].icell.Ien Vbias 0.19149f
C2579 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04035f
C2580 XThR.XTBN.Y a_n997_1803# 0.22873f
C2581 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04035f
C2582 XA.XIR[2].XIC[12].icell.PUM VPWR 0.01079f
C2583 XA.XIR[7].XIC[12].icell.Ien VPWR 0.21079f
C2584 XThR.Tn[11] Vbias 1.38584f
C2585 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C2586 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.14207f
C2587 XThR.XTB6.A data[4] 0.48493f
C2588 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.04573f
C2589 XA.XIR[1].XIC[14].icell.PUM VPWR 0.01079f
C2590 XA.XIR[7].XIC[9].icell.PDM Vbias 0.03922f
C2591 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04035f
C2592 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C2593 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.04573f
C2594 XA.XIR[10].XIC[11].icell.Ien VPWR 0.21079f
C2595 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C2596 XA.XIR[15].XIC[7].icell.PDM Vbias 0.03922f
C2597 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C2598 XThC.Tn[7] XThR.Tn[2] 0.39125f
C2599 XA.XIR[3].XIC[1].icell.Ien VPWR 0.21079f
C2600 XThC.XTB7.B a_6243_9615# 0.01743f
C2601 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02601f
C2602 XA.XIR[12].XIC[1].icell.PUM VPWR 0.01079f
C2603 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C2604 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C2605 XA.XIR[13].XIC[12].icell.PUM VPWR 0.01079f
C2606 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02601f
C2607 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.04036f
C2608 XA.XIR[9].XIC[5].icell.PDM Vbias 0.03922f
C2609 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.14207f
C2610 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02804f
C2611 XA.XIR[7].XIC[10].icell.PDM VPWR 0.01373f
C2612 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C2613 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.13138f
C2614 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C2615 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02601f
C2616 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C2617 XA.XIR[3].XIC[10].icell.Ien Iout 0.06763f
C2618 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C2619 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C2620 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01714f
C2621 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.14207f
C2622 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C2623 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.14207f
C2624 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C2625 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.14207f
C2626 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C2627 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C2628 XA.XIR[2].XIC[3].icell.Ien Iout 0.06763f
C2629 XThC.Tn[3] XThR.Tn[6] 0.39123f
C2630 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02601f
C2631 XA.XIR[1].XIC[10].icell.PDM Vbias 0.03922f
C2632 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C2633 XA.XIR[1].XIC[5].icell.Ien Iout 0.06763f
C2634 XA.XIR[6].XIC[13].icell.Ien Vbias 0.19151f
C2635 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.14207f
C2636 XA.XIR[9].XIC[6].icell.PDM VPWR 0.01373f
C2637 XA.XIR[10].XIC[14].icell.Ien Vbias 0.19151f
C2638 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C2639 XA.XIR[13].XIC[13].icell.Ien VPWR 0.21079f
C2640 XA.XIR[4].XIC[10].icell.PDM Vbias 0.03922f
C2641 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02601f
C2642 XA.XIR[12].XIC[12].icell.PDM VPWR 0.01373f
C2643 XThC.Tn[5] XThR.Tn[11] 0.39123f
C2644 XA.XIR[8].XIC[13].icell.Ien Iout 0.06763f
C2645 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C2646 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C2647 XA.XIR[14].XIC[7].icell.Ien Vbias 0.19151f
C2648 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.04623f
C2649 XThC.Tn[1] Iout 0.0226f
C2650 XA.XIR[13].XIC[9].icell.Ien Vbias 0.19151f
C2651 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01714f
C2652 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04035f
C2653 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.04573f
C2654 XThC.Tn[11] Vbias 0.3277f
C2655 XA.XIR[1].XIC[11].icell.PDM VPWR 0.01373f
C2656 XA.XIR[3].XIC[9].icell.Ien VPWR 0.21079f
C2657 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.04575f
C2658 XA.XIR[6].XIC[14].icell.PUM VPWR 0.01079f
C2659 XThC.Tn[9] XThR.Tn[13] 0.39123f
C2660 XA.XIR[4].XIC[11].icell.PDM VPWR 0.01373f
C2661 XA.XIR[2].XIC[2].icell.Ien VPWR 0.21079f
C2662 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C2663 XA.XIR[0].XIC_15.icell.Ien Iout 0.06774f
C2664 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C2665 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04035f
C2666 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02601f
C2667 XA.XIR[1].XIC[4].icell.Ien VPWR 0.21079f
C2668 XA.XIR[14].XIC[8].icell.PUM VPWR 0.01079f
C2669 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.04573f
C2670 XThC.Tn[12] XThR.Tn[9] 0.39123f
C2671 XA.XIR[6].XIC[0].icell.Ien Iout 0.06763f
C2672 XThC.Tn[8] XThR.Tn[8] 0.39123f
C2673 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04035f
C2674 XA.XIR[13].XIC[10].icell.PUM VPWR 0.01079f
C2675 XA.XIR[8].XIC[12].icell.Ien VPWR 0.21079f
C2676 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.02965f
C2677 bias[1] bias[0] 0.6046f
C2678 bias[2] Vbias 0.4026f
C2679 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04035f
C2680 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.04573f
C2681 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C2682 XThC.XTBN.Y XThC.Tn[6] 0.48987f
C2683 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C2684 XThR.XTB7.B a_n997_3979# 0.01152f
C2685 XThC.Tn[3] XThR.Tn[4] 0.39123f
C2686 XA.XIR[5].XIC[1].icell.Ien Vbias 0.19151f
C2687 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C2688 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04035f
C2689 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C2690 XThR.Tn[14] Vbias 1.38585f
C2691 XA.XIR[11].XIC[0].icell.PDM Vbias 0.03915f
C2692 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C2693 XA.XIR[0].XIC[14].icell.Ien VPWR 0.2042f
C2694 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C2695 XA.XIR[6].XIC[5].icell.Ien Iout 0.06763f
C2696 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.14207f
C2697 XThC.Tn[7] XThR.Tn[10] 0.39123f
C2698 XA.XIR[10].XIC[4].icell.PDM Vbias 0.03922f
C2699 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.14207f
C2700 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C2701 XA.XIR[10].XIC[12].icell.Ien Vbias 0.19151f
C2702 XA.XIR[13].XIC[11].icell.Ien VPWR 0.21079f
C2703 a_7651_9569# XThC.Tn[8] 0.1927f
C2704 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04035f
C2705 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02601f
C2706 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.14207f
C2707 XA.XIR[5].XIC[2].icell.PUM VPWR 0.01079f
C2708 XA.XIR[5].XIC[6].icell.Ien Vbias 0.19151f
C2709 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13586f
C2710 XA.XIR[11].XIC[1].icell.PDM VPWR 0.01373f
C2711 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C2712 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.04573f
C2713 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02601f
C2714 XA.XIR[10].XIC[5].icell.PDM VPWR 0.01373f
C2715 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C2716 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.04573f
C2717 XA.XIR[11].XIC[4].icell.Ien Iout 0.06763f
C2718 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02602f
C2719 XThR.XTB7.B XThR.Tn[7] 0.07415f
C2720 XA.XIR[6].XIC[4].icell.Ien VPWR 0.21079f
C2721 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.04573f
C2722 XA.XIR[10].XIC[6].icell.Ien Iout 0.06763f
C2723 XThR.XTB7.B a_n997_2891# 0.0168f
C2724 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02601f
C2725 XA.XIR[0].XIC[12].icell.PDM Vbias 0.03922f
C2726 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.04573f
C2727 XA.XIR[5].XIC[7].icell.PUM VPWR 0.01079f
C2728 XA.XIR[12].XIC[11].icell.PDM VPWR 0.01373f
C2729 XThC.XTB7.B a_8963_9569# 0.02071f
C2730 XA.XIR[13].XIC[14].icell.Ien Vbias 0.19151f
C2731 XA.XIR[3].XIC_15.icell.Ien Iout 0.0694f
C2732 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C2733 XThC.Tn[5] XThR.Tn[14] 0.39123f
C2734 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.14207f
C2735 XThC.XTB6.A XThC.XTB7.A 0.44014f
C2736 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01714f
C2737 XA.XIR[2].XIC[8].icell.Ien Iout 0.06763f
C2738 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C2739 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C2740 XA.XIR[1].XIC[10].icell.Ien Iout 0.06763f
C2741 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C2742 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.04573f
C2743 XA.XIR[0].XIC[13].icell.PDM VPWR 0.01334f
C2744 XA.XIR[11].XIC[3].icell.Ien VPWR 0.21079f
C2745 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C2746 XThC.XTB2.Y XThC.Tn[1] 0.18085f
C2747 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C2748 XA.XIR[10].XIC[5].icell.Ien VPWR 0.21079f
C2749 XA.XIR[10].XIC[10].icell.Ien Vbias 0.19151f
C2750 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C2751 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.04573f
C2752 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C2753 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C2754 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04035f
C2755 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04035f
C2756 XA.XIR[3].XIC[14].icell.Ien VPWR 0.20455f
C2757 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02601f
C2758 XThR.XTBN.Y a_n997_3979# 0.23021f
C2759 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C2760 XA.XIR[2].XIC[7].icell.Ien VPWR 0.21079f
C2761 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04023f
C2762 XA.XIR[1].XIC[9].icell.Ien VPWR 0.21079f
C2763 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C2764 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02601f
C2765 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.14207f
C2766 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C2767 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02601f
C2768 XThC.Tn[0] Vbias 0.23747f
C2769 XA.XIR[6].XIC[3].icell.PDM Vbias 0.03922f
C2770 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C2771 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C2772 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.04573f
C2773 XThC.XTB3.Y a_4067_9615# 0.23056f
C2774 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C2775 XA.XIR[14].XIC[0].icell.PDM Vbias 0.03915f
C2776 XA.XIR[5].XIC[10].icell.PDM Vbias 0.03922f
C2777 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C2778 a_4067_9615# XThC.Tn[2] 0.27296f
C2779 XThC.Tn[7] XThR.Tn[13] 0.39123f
C2780 XA.XIR[13].XIC[4].icell.PDM Vbias 0.03922f
C2781 XA.XIR[13].XIC[12].icell.Ien Vbias 0.19151f
C2782 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.14207f
C2783 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02601f
C2784 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.0404f
C2785 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.04573f
C2786 XThC.Tn[1] XThR.Tn[9] 0.39123f
C2787 XA.XIR[12].XIC[9].icell.PDM Vbias 0.03922f
C2788 XThC.XTB5.A XThC.XTB6.A 1.80461f
C2789 XA.XIR[9].XIC[2].icell.Ien Vbias 0.19151f
C2790 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C2791 XThC.Tn[6] XThR.Tn[8] 0.39123f
C2792 XA.XIR[6].XIC[4].icell.PDM VPWR 0.01373f
C2793 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04023f
C2794 XA.XIR[6].XIC[10].icell.Ien Iout 0.06763f
C2795 XThR.XTB7.A a_n1049_6699# 0.02294f
C2796 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.14207f
C2797 XA.XIR[14].XIC[1].icell.PDM VPWR 0.01373f
C2798 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.14207f
C2799 XThR.XTB5.Y VPWR 1.02746f
C2800 XA.XIR[5].XIC[11].icell.PDM VPWR 0.01373f
C2801 XThR.XTBN.Y XThR.Tn[7] 0.89976f
C2802 XThR.XTBN.Y a_n997_2891# 0.22804f
C2803 XA.XIR[13].XIC[5].icell.PDM VPWR 0.01373f
C2804 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02602f
C2805 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C2806 XA.XIR[14].XIC[4].icell.Ien Iout 0.06763f
C2807 XA.XIR[12].XIC[10].icell.PDM VPWR 0.01373f
C2808 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02601f
C2809 XA.XIR[5].XIC[11].icell.Ien Vbias 0.19151f
C2810 XA.XIR[13].XIC[6].icell.Ien Iout 0.06763f
C2811 XA.XIR[9].XIC[3].icell.PUM VPWR 0.01079f
C2812 XThC.XTB3.Y XThC.Tn[3] 0.01335f
C2813 XA.XIR[8].XIC[7].icell.PDM Vbias 0.03922f
C2814 XA.XIR[3].XIC[5].icell.PDM Vbias 0.03922f
C2815 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01714f
C2816 XThC.Tn[2] XThC.Tn[3] 0.59595f
C2817 XThR.Tn[5] XThR.Tn[6] 0.10623f
C2818 XA.XIR[2].XIC[11].icell.PDM Vbias 0.03922f
C2819 XA.XIR[11].XIC[9].icell.Ien Iout 0.06763f
C2820 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C2821 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04035f
C2822 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02601f
C2823 XA.XIR[12].XIC[6].icell.Ien Vbias 0.19151f
C2824 XA.XIR[6].XIC[9].icell.Ien VPWR 0.21079f
C2825 XA.XIR[10].XIC_15.icell.Ien Vbias 0.19187f
C2826 VPWR Vbias 0.1158p
C2827 XA.XIR[5].XIC[12].icell.PUM VPWR 0.01079f
C2828 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.04575f
C2829 XThR.XTBN.A data[5] 0.0148f
C2830 XThR.Tn[10] a_n997_2891# 0.1927f
C2831 XThC.XTB6.A data[0] 0.48493f
C2832 XA.XIR[3].XIC[6].icell.PDM VPWR 0.01373f
C2833 XA.XIR[14].XIC[3].icell.Ien VPWR 0.21134f
C2834 XA.XIR[8].XIC[8].icell.PDM VPWR 0.01373f
C2835 XThC.Tn[9] XThR.Tn[7] 0.39123f
C2836 XA.XIR[2].XIC[12].icell.PDM VPWR 0.01373f
C2837 XA.XIR[13].XIC[5].icell.Ien VPWR 0.21079f
C2838 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C2839 XA.XIR[2].XIC[13].icell.Ien Iout 0.06763f
C2840 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04035f
C2841 XThR.XTB1.Y VPWR 1.13493f
C2842 XA.XIR[13].XIC[10].icell.Ien Vbias 0.19151f
C2843 XThC.XTB2.Y a_3523_10575# 0.01006f
C2844 XThC.XTB7.Y XThC.Tn[11] 0.07422f
C2845 XA.XIR[12].XIC[7].icell.PUM VPWR 0.01079f
C2846 XA.XIR[1].XIC_15.icell.Ien Iout 0.0694f
C2847 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C2848 XThR.XTB6.Y a_n1319_5611# 0.01283f
C2849 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C2850 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02601f
C2851 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.04036f
C2852 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.0176f
C2853 XA.XIR[11].XIC[8].icell.Ien VPWR 0.21079f
C2854 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02601f
C2855 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C2856 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.04573f
C2857 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02804f
C2858 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C2859 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02601f
C2860 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02601f
C2861 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04035f
C2862 XA.XIR[5].XIC[3].icell.Ien Iout 0.06763f
C2863 XThR.Tn[4] XThR.Tn[5] 0.11363f
C2864 XThC.Tn[8] XThR.Tn[3] 0.39123f
C2865 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04035f
C2866 XA.XIR[2].XIC[12].icell.Ien VPWR 0.21079f
C2867 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C2868 XA.XIR[10].XIC[0].icell.PUM VPWR 0.01079f
C2869 XA.XIR[1].XIC[14].icell.Ien VPWR 0.20455f
C2870 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.04261f
C2871 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.14207f
C2872 XThC.Tn[5] VPWR 7.01912f
C2873 XA.XIR[7].XIC[11].icell.PDM Vbias 0.03922f
C2874 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04023f
C2875 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02601f
C2876 XA.XIR[15].XIC[9].icell.PDM Vbias 0.03922f
C2877 XA.XIR[4].XIC[4].icell.Ien Vbias 0.19151f
C2878 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C2879 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.13413f
C2880 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C2881 XThC.Tn[11] XThR.Tn[0] 0.39146f
C2882 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.04573f
C2883 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.04573f
C2884 XThC.Tn[13] XThR.Tn[5] 0.39123f
C2885 XA.XIR[12].XIC[1].icell.Ien VPWR 0.21079f
C2886 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.04573f
C2887 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C2888 XA.XIR[9].XIC[7].icell.PDM Vbias 0.03922f
C2889 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.14207f
C2890 XThR.XTBN.Y a_n997_1579# 0.23006f
C2891 XA.XIR[5].XIC[2].icell.Ien VPWR 0.21079f
C2892 XA.XIR[7].XIC[12].icell.PDM VPWR 0.01373f
C2893 XThR.XTB7.Y a_n1049_5317# 0.27822f
C2894 XA.XIR[9].XIC[7].icell.Ien Vbias 0.19151f
C2895 XA.XIR[11].XIC[14].icell.Ien Iout 0.06763f
C2896 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.04573f
C2897 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C2898 XThR.Tn[6] Iout 1.10102f
C2899 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01714f
C2900 XA.XIR[4].XIC[5].icell.PUM VPWR 0.01079f
C2901 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C2902 XA.XIR[6].XIC_15.icell.Ien Iout 0.0694f
C2903 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02601f
C2904 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02601f
C2905 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C2906 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.14207f
C2907 XA.XIR[1].XIC[12].icell.PDM Vbias 0.03922f
C2908 XThC.Tn[8] data[0] 0.01744f
C2909 XA.XIR[9].XIC[8].icell.PDM VPWR 0.01373f
C2910 XA.XIR[14].XIC[9].icell.Ien Iout 0.06763f
C2911 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C2912 XA.XIR[0].XIC[0].icell.PDM VPWR 0.01334f
C2913 XA.XIR[7].XIC[3].icell.Ien Vbias 0.19151f
C2914 XA.XIR[4].XIC[12].icell.PDM Vbias 0.03922f
C2915 XA.XIR[9].XIC[8].icell.PUM VPWR 0.01079f
C2916 XThC.Tn[10] XThR.Tn[2] 0.39125f
C2917 XThC.XTB7.B Vbias 0.11961f
C2918 XA.XIR[13].XIC_15.icell.Ien Vbias 0.19187f
C2919 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.14207f
C2920 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C2921 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04035f
C2922 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C2923 XThR.Tn[11] XThR.Tn[12] 0.15424f
C2924 XA.XIR[1].XIC[13].icell.PDM VPWR 0.01373f
C2925 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.04573f
C2926 XA.XIR[6].XIC[14].icell.Ien VPWR 0.20455f
C2927 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04035f
C2928 XA.XIR[4].XIC[13].icell.PDM VPWR 0.01373f
C2929 XA.XIR[7].XIC[4].icell.PUM VPWR 0.01079f
C2930 XThC.XTB7.A XThC.Tn[6] 0.10502f
C2931 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04035f
C2932 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.0176f
C2933 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02601f
C2934 XA.XIR[14].XIC[8].icell.Ien VPWR 0.21134f
C2935 XThR.XTB5.A XThR.XTBN.A 0.06303f
C2936 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.04261f
C2937 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04035f
C2938 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C2939 XThR.Tn[4] Iout 1.10104f
C2940 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02601f
C2941 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C2942 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.04574f
C2943 XThC.Tn[8] XThR.Tn[11] 0.39123f
C2944 XA.XIR[11].XIC[12].icell.Ien Iout 0.06763f
C2945 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.40998f
C2946 XA.XIR[15].XIC[1].icell.Ien Vbias 0.15955f
C2947 XThR.XTBN.Y a_n1049_6699# 0.07601f
C2948 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C2949 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04035f
C2950 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C2951 XThC.Tn[7] XThR.Tn[7] 0.39123f
C2952 XA.XIR[11].XIC[2].icell.PDM Vbias 0.03922f
C2953 XA.XIR[13].XIC[0].icell.PUM VPWR 0.01079f
C2954 XThC.Tn[13] Iout 0.02211f
C2955 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04035f
C2956 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C2957 XA.XIR[10].XIC[6].icell.PDM Vbias 0.03922f
C2958 XA.XIR[5].XIC[8].icell.Ien Iout 0.06763f
C2959 XThC.XTB6.Y XThC.Tn[13] 0.32317f
C2960 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.02965f
C2961 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04035f
C2962 XThR.XTB7.A data[4] 0.8689f
C2963 XA.XIR[15].XIC[2].icell.PUM VPWR 0.01079f
C2964 XThC.Tn[11] XThR.Tn[1] 0.39128f
C2965 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.04573f
C2966 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C2967 XA.XIR[15].XIC[6].icell.Ien Vbias 0.15955f
C2968 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.14207f
C2969 XThR.XTB4.Y a_n1049_6699# 0.23756f
C2970 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C2971 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C2972 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C2973 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C2974 XA.XIR[11].XIC[3].icell.PDM VPWR 0.01373f
C2975 XA.XIR[4].XIC[9].icell.Ien Vbias 0.19151f
C2976 XThC.Tn[11] XThR.Tn[12] 0.39123f
C2977 XA.XIR[12].XIC[3].icell.Ien Iout 0.06763f
C2978 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C2979 XA.XIR[0].XIC[0].icell.Ien Vbias 0.1919f
C2980 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.04573f
C2981 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C2982 XThR.XTB7.B XThR.Tn[8] 0.05091f
C2983 XA.XIR[10].XIC[7].icell.PDM VPWR 0.01373f
C2984 XA.XIR[14].XIC[14].icell.Ien Iout 0.06763f
C2985 XA.XIR[8].XIC[3].icell.Ien Vbias 0.19151f
C2986 XThC.XTBN.Y XThC.Tn[9] 0.39482f
C2987 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02601f
C2988 XThC.Tn[6] XThR.Tn[3] 0.39123f
C2989 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C2990 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.14207f
C2991 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08212f
C2992 XA.XIR[15].XIC[7].icell.PUM VPWR 0.01079f
C2993 XA.XIR[0].XIC[14].icell.PDM Vbias 0.03922f
C2994 XA.XIR[5].XIC[7].icell.Ien VPWR 0.21079f
C2995 XThR.XTB7.A a_n1049_5611# 0.01824f
C2996 XThC.Tn[0] XThR.Tn[0] 0.39682f
C2997 XA.XIR[9].XIC[12].icell.Ien Vbias 0.19151f
C2998 XThC.Tn[10] XThR.Tn[10] 0.39123f
C2999 XA.XIR[4].XIC[10].icell.PUM VPWR 0.01079f
C3000 XThC.Tn[2] XThR.Tn[5] 0.39123f
C3001 XA.XIR[0].XIC[1].icell.PUM VPWR 0.01038f
C3002 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02601f
C3003 XA.XIR[0].XIC[5].icell.Ien Vbias 0.19186f
C3004 XThC.Tn[9] XThC.Tn[10] 0.0671f
C3005 XA.XIR[11].XIC[10].icell.Ien Iout 0.06763f
C3006 XA.XIR[8].XIC[4].icell.PUM VPWR 0.01079f
C3007 XThR.Tn[13] a_n997_1579# 0.19413f
C3008 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04035f
C3009 XA.XIR[12].XIC[2].icell.Ien VPWR 0.21079f
C3010 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07467f
C3011 XThC.XTB7.Y VPWR 1.07719f
C3012 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C3013 XA.XIR[7].XIC[8].icell.Ien Vbias 0.19151f
C3014 XA.XIR[9].XIC[13].icell.PUM VPWR 0.01079f
C3015 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C3016 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.14207f
C3017 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C3018 XA.XIR[0].XIC[6].icell.PUM VPWR 0.01038f
C3019 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C3020 XThR.XTBN.A XThR.Tn[9] 0.12398f
C3021 XA.XIR[11].XIC[0].icell.Ien Iout 0.06763f
C3022 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C3023 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C3024 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3025 XA.XIR[7].XIC[9].icell.PUM VPWR 0.01079f
C3026 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02602f
C3027 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C3028 XThR.XTB6.A VPWR 0.6882f
C3029 XThC.Tn[8] XThR.Tn[14] 0.39123f
C3030 XA.XIR[10].XIC[0].icell.Ien Vbias 0.19149f
C3031 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04035f
C3032 XA.XIR[14].XIC[12].icell.Ien Iout 0.06763f
C3033 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C3034 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C3035 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.40995f
C3036 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C3037 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02601f
C3038 XA.XIR[6].XIC[5].icell.PDM Vbias 0.03922f
C3039 XThR.XTB1.Y a_n1049_8581# 0.21263f
C3040 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.04261f
C3041 XA.XIR[14].XIC[2].icell.PDM Vbias 0.03922f
C3042 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.04628f
C3043 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.14207f
C3044 XA.XIR[5].XIC[12].icell.PDM Vbias 0.03922f
C3045 XA.XIR[6].XIC[0].icell.PUM VPWR 0.01079f
C3046 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C3047 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C3048 XThR.XTB7.B data[4] 0.01382f
C3049 XA.XIR[13].XIC[6].icell.PDM Vbias 0.03922f
C3050 XA.XIR[9].XIC[4].icell.Ien Iout 0.06763f
C3051 XThR.Tn[0] VPWR 9.73945f
C3052 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C3053 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04035f
C3054 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C3055 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.02965f
C3056 XThR.XTB7.B a_n997_3755# 0.01174f
C3057 XA.XIR[10].XIC[1].icell.PUM VPWR 0.01079f
C3058 XThC.Tn[4] XThR.Tn[6] 0.39123f
C3059 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C3060 XA.XIR[6].XIC[6].icell.PDM VPWR 0.01373f
C3061 XThR.XTBN.Y XThR.Tn[8] 0.47809f
C3062 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C3063 XA.XIR[5].XIC[13].icell.PDM VPWR 0.01373f
C3064 XA.XIR[14].XIC[3].icell.PDM VPWR 0.01373f
C3065 XA.XIR[5].XIC[13].icell.Ien Iout 0.06763f
C3066 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.04573f
C3067 XThC.Tn[6] XThR.Tn[11] 0.39123f
C3068 XA.XIR[3].XIC[5].icell.Ien Vbias 0.19151f
C3069 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C3070 XA.XIR[13].XIC[7].icell.PDM VPWR 0.01373f
C3071 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C3072 XThC.Tn[2] Iout 0.02214f
C3073 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C3074 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C3075 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C3076 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02601f
C3077 XThC.Tn[12] Vbias 0.32228f
C3078 XA.XIR[9].XIC[3].icell.Ien VPWR 0.21079f
C3079 XA.XIR[11].XIC_15.icell.Ien Iout 0.0694f
C3080 XA.XIR[3].XIC[7].icell.PDM Vbias 0.03922f
C3081 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C3082 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.04575f
C3083 XA.XIR[8].XIC[9].icell.PDM Vbias 0.03922f
C3084 XA.XIR[4].XIC[14].icell.Ien Vbias 0.19151f
C3085 XA.XIR[12].XIC[8].icell.Ien Iout 0.06763f
C3086 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C3087 VPWR data[7] 0.21201f
C3088 XA.XIR[2].XIC[13].icell.PDM Vbias 0.03922f
C3089 XThC.Tn[10] XThR.Tn[13] 0.39123f
C3090 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.04573f
C3091 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02601f
C3092 XA.XIR[8].XIC[8].icell.Ien Vbias 0.19151f
C3093 XThC.Tn[0] XThR.Tn[1] 0.39127f
C3094 XA.XIR[3].XIC[6].icell.PUM VPWR 0.01079f
C3095 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02602f
C3096 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04035f
C3097 XA.XIR[1].XIC[0].icell.PDM VPWR 0.01373f
C3098 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02601f
C3099 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C3100 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C3101 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C3102 XA.XIR[10].XIC_15.icell.PDM Vbias 0.03927f
C3103 XThC.Tn[13] XThR.Tn[9] 0.39123f
C3104 XA.XIR[14].XIC[10].icell.Ien Iout 0.06763f
C3105 XThR.XTB7.A XThR.Tn[3] 0.0306f
C3106 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C3107 XA.XIR[5].XIC[12].icell.Ien VPWR 0.21079f
C3108 XA.XIR[4].XIC[0].icell.PDM VPWR 0.01373f
C3109 XThC.Tn[0] XThR.Tn[12] 0.39118f
C3110 XThC.Tn[9] XThR.Tn[8] 0.39123f
C3111 XThC.XTB6.A VPWR 0.68179f
C3112 XA.XIR[3].XIC[8].icell.PDM VPWR 0.01373f
C3113 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C3114 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01768f
C3115 XA.XIR[8].XIC[10].icell.PDM VPWR 0.01373f
C3116 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C3117 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C3118 XThC.XTBN.A a_7875_9569# 0.01939f
C3119 XA.XIR[2].XIC[14].icell.PDM VPWR 0.01349f
C3120 XA.XIR[0].XIC[10].icell.Ien Vbias 0.19186f
C3121 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C3122 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C3123 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C3124 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04035f
C3125 XThC.XTBN.Y XThC.Tn[7] 0.85468f
C3126 XThC.Tn[4] XThR.Tn[4] 0.39123f
C3127 XA.XIR[8].XIC[9].icell.PUM VPWR 0.01079f
C3128 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C3129 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C3130 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C3131 XA.XIR[12].XIC[7].icell.Ien VPWR 0.21079f
C3132 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3133 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.04573f
C3134 XA.XIR[4].XIC[1].icell.Ien Iout 0.06763f
C3135 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C3136 XA.XIR[7].XIC[13].icell.Ien Vbias 0.19151f
C3137 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.04574f
C3138 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3139 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.14207f
C3140 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.14207f
C3141 XA.XIR[0].XIC[11].icell.PUM VPWR 0.01038f
C3142 XThC.XTBN.A data[1] 0.01444f
C3143 XA.XIR[13].XIC[0].icell.Ien Vbias 0.19149f
C3144 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C3145 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04035f
C3146 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.40988f
C3147 XA.XIR[15].XIC[3].icell.Ien Iout 0.07153f
C3148 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C3149 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04035f
C3150 XThR.XTBN.Y a_n997_3755# 0.229f
C3151 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C3152 XA.XIR[7].XIC[14].icell.PUM VPWR 0.01079f
C3153 XA.XIR[4].XIC[6].icell.Ien Iout 0.06763f
C3154 XA.XIR[1].XIC[0].icell.Ien VPWR 0.21079f
C3155 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C3156 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.14207f
C3157 XA.XIR[7].XIC[13].icell.PDM Vbias 0.03922f
C3158 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C3159 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C3160 XA.XIR[4].XIC[0].icell.Ien VPWR 0.21079f
C3161 XThR.Tn[1] VPWR 9.7268f
C3162 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02601f
C3163 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C3164 XA.XIR[13].XIC[1].icell.PUM VPWR 0.01079f
C3165 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.14207f
C3166 XThC.XTBN.Y a_3773_9615# 0.08456f
C3167 XA.XIR[7].XIC[0].icell.Ien Iout 0.06763f
C3168 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.14207f
C3169 XThR.Tn[12] VPWR 10.6247f
C3170 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C3171 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C3172 XA.XIR[9].XIC[9].icell.Ien Iout 0.06763f
C3173 XThR.XTBN.Y a_n1049_5611# 0.0768f
C3174 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C3175 a_10915_9569# Vbias 0.01383f
C3176 XA.XIR[9].XIC[9].icell.PDM Vbias 0.03922f
C3177 XThC.Tn[6] XThR.Tn[14] 0.39123f
C3178 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C3179 XA.XIR[15].XIC[2].icell.Ien VPWR 0.3396f
C3180 XA.XIR[0].XIC[1].icell.PDM Vbias 0.03922f
C3181 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C3182 XA.XIR[0].XIC[2].icell.Ien Iout 0.06712f
C3183 XA.XIR[7].XIC[14].icell.PDM VPWR 0.01349f
C3184 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C3185 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.14207f
C3186 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C3187 XA.XIR[4].XIC[5].icell.Ien VPWR 0.21079f
C3188 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.04573f
C3189 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C3190 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C3191 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C3192 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02601f
C3193 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C3194 XA.XIR[14].XIC_15.icell.Ien Iout 0.0694f
C3195 XA.XIR[7].XIC[5].icell.Ien Iout 0.06763f
C3196 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08254f
C3197 XA.XIR[3].XIC[10].icell.Ien Vbias 0.19151f
C3198 XA.XIR[1].XIC[14].icell.PDM Vbias 0.03922f
C3199 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C3200 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02602f
C3201 XA.XIR[10].XIC[14].icell.PDM Vbias 0.03922f
C3202 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.04573f
C3203 XThC.Tn[8] VPWR 7.96808f
C3204 XA.XIR[9].XIC[10].icell.PDM VPWR 0.01373f
C3205 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02601f
C3206 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08254f
C3207 XA.XIR[0].XIC[2].icell.PDM VPWR 0.01334f
C3208 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C3209 XA.XIR[4].XIC[14].icell.PDM Vbias 0.03922f
C3210 XA.XIR[2].XIC[3].icell.Ien Vbias 0.19151f
C3211 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.14207f
C3212 XA.XIR[13].XIC_15.icell.PDM Vbias 0.03927f
C3213 XA.XIR[9].XIC[8].icell.Ien VPWR 0.21079f
C3214 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C3215 XA.XIR[1].XIC[5].icell.Ien Vbias 0.19162f
C3216 XA.XIR[7].XIC[0].icell.PUM VPWR 0.01079f
C3217 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C3218 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C3219 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.14207f
C3220 XThC.XTB6.A XThC.XTB7.B 1.47641f
C3221 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.04573f
C3222 XThR.XTB5.Y a_n1319_6405# 0.01188f
C3223 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04035f
C3224 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C3225 XA.XIR[8].XIC[13].icell.Ien Vbias 0.19151f
C3226 a_n1049_5317# VPWR 0.72143f
C3227 XA.XIR[3].XIC[11].icell.PUM VPWR 0.01079f
C3228 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07604f
C3229 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C3230 XThC.Tn[1] Vbias 0.32784f
C3231 XA.XIR[7].XIC[4].icell.Ien VPWR 0.21079f
C3232 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07604f
C3233 XA.XIR[2].XIC[4].icell.PUM VPWR 0.01079f
C3234 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C3235 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C3236 XThR.Tn[2] XThR.Tn[3] 0.14493f
C3237 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C3238 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3239 XA.XIR[1].XIC[6].icell.PUM VPWR 0.01079f
C3240 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C3241 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.14207f
C3242 XA.XIR[0].XIC_15.icell.Ien Vbias 0.19223f
C3243 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04023f
C3244 XA.XIR[8].XIC[14].icell.PUM VPWR 0.01079f
C3245 XThC.Tn[2] XThR.Tn[9] 0.39123f
C3246 XThR.XTBN.Y a_n997_715# 0.21503f
C3247 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.04573f
C3248 XA.XIR[6].XIC[0].icell.Ien Vbias 0.19149f
C3249 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.14207f
C3250 XThC.Tn[7] XThR.Tn[8] 0.39123f
C3251 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C3252 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C3253 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C3254 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.04629f
C3255 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04035f
C3256 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.14207f
C3257 XA.XIR[3].XIC[2].icell.Ien Iout 0.06763f
C3258 XA.XIR[11].XIC[4].icell.PDM Vbias 0.03922f
C3259 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01602f
C3260 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.14207f
C3261 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.04575f
C3262 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C3263 XThR.XTB7.B a_n997_2667# 0.02071f
C3264 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.14207f
C3265 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04035f
C3266 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.04573f
C3267 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02601f
C3268 XA.XIR[10].XIC[8].icell.PDM Vbias 0.03922f
C3269 XA.XIR[5].XIC[0].icell.PDM VPWR 0.01373f
C3270 XA.XIR[15].XIC[8].icell.Ien Iout 0.07153f
C3271 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C3272 XA.XIR[6].XIC[1].icell.PUM VPWR 0.01079f
C3273 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04035f
C3274 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.04573f
C3275 a_n1049_6405# VPWR 0.72203f
C3276 XA.XIR[6].XIC[5].icell.Ien Vbias 0.19151f
C3277 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C3278 XA.XIR[4].XIC[11].icell.Ien Iout 0.06763f
C3279 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.14207f
C3280 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.0125f
C3281 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02601f
C3282 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C3283 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.04573f
C3284 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C3285 XA.XIR[8].XIC[5].icell.Ien Iout 0.06763f
C3286 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C3287 XA.XIR[11].XIC[5].icell.PDM VPWR 0.01373f
C3288 XA.XIR[10].XIC[9].icell.PDM VPWR 0.01373f
C3289 VPWR data[3] 0.20846f
C3290 XA.XIR[2].XIC[0].icell.PDM Vbias 0.03915f
C3291 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C3292 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.04573f
C3293 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.04573f
C3294 XThR.XTBN.Y XThR.Tn[3] 0.625f
C3295 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C3296 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01244f
C3297 XA.XIR[9].XIC[14].icell.Ien Iout 0.06763f
C3298 XA.XIR[10].XIC[13].icell.PDM Vbias 0.03922f
C3299 a_n1049_8581# XThR.Tn[0] 0.2685f
C3300 XA.XIR[6].XIC[6].icell.PUM VPWR 0.01079f
C3301 XThR.XTB7.B XThR.Tn[11] 0.03888f
C3302 XThC.Tn[10] XThR.Tn[7] 0.39123f
C3303 XA.XIR[15].XIC[7].icell.Ien VPWR 0.3396f
C3304 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C3305 XA.XIR[0].XIC[7].icell.Ien Iout 0.06712f
C3306 XA.XIR[11].XIC[4].icell.Ien Vbias 0.19151f
C3307 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.04574f
C3308 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.14207f
C3309 XA.XIR[13].XIC[14].icell.PDM Vbias 0.03922f
C3310 XThC.XTB7.B XThC.Tn[8] 0.0473f
C3311 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.04573f
C3312 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.40895f
C3313 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C3314 XA.XIR[4].XIC[10].icell.Ien VPWR 0.21079f
C3315 XThC.XTB7.Y XThC.Tn[12] 0.07091f
C3316 XA.XIR[10].XIC[6].icell.Ien Vbias 0.19151f
C3317 XA.XIR[0].XIC[1].icell.Ien VPWR 0.21044f
C3318 XA.XIR[2].XIC[1].icell.PDM VPWR 0.01373f
C3319 XA.XIR[11].XIC[14].icell.PUM VPWR 0.01079f
C3320 XA.XIR[7].XIC[10].icell.Ien Iout 0.06763f
C3321 XA.XIR[8].XIC[4].icell.Ien VPWR 0.21079f
C3322 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C3323 XA.XIR[3].XIC_15.icell.Ien Vbias 0.19187f
C3324 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C3325 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C3326 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C3327 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04035f
C3328 XA.XIR[11].XIC[5].icell.PUM VPWR 0.01079f
C3329 XA.XIR[2].XIC[8].icell.Ien Vbias 0.19151f
C3330 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.04573f
C3331 XA.XIR[8].XIC[0].icell.Ien Iout 0.06763f
C3332 XA.XIR[9].XIC[13].icell.Ien VPWR 0.21079f
C3333 XA.XIR[1].XIC[10].icell.Ien Vbias 0.19162f
C3334 XA.XIR[10].XIC[7].icell.PUM VPWR 0.01079f
C3335 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C3336 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.04573f
C3337 XThC.Tn[9] XThR.Tn[3] 0.39123f
C3338 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.14207f
C3339 XA.XIR[0].XIC[6].icell.Ien VPWR 0.21048f
C3340 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C3341 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3342 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.04573f
C3343 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C3344 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.0176f
C3345 XThC.Tn[6] VPWR 7.0553f
C3346 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C3347 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.14207f
C3348 XA.XIR[7].XIC[9].icell.Ien VPWR 0.21079f
C3349 XA.XIR[2].XIC[9].icell.PUM VPWR 0.01079f
C3350 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.14207f
C3351 XThC.Tn[12] XThR.Tn[0] 0.39146f
C3352 XA.XIR[1].XIC[11].icell.PUM VPWR 0.01079f
C3353 XThC.Tn[14] XThR.Tn[5] 0.39123f
C3354 XA.XIR[7].XIC[0].icell.PDM Vbias 0.03915f
C3355 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04035f
C3356 XThR.XTBN.Y a_n997_2667# 0.22784f
C3357 XA.XIR[6].XIC[7].icell.PDM Vbias 0.03922f
C3358 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C3359 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C3360 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08254f
C3361 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C3362 XA.XIR[14].XIC[4].icell.PDM Vbias 0.03922f
C3363 XA.XIR[5].XIC[14].icell.PDM Vbias 0.03922f
C3364 XThR.Tn[8] a_n997_3979# 0.1927f
C3365 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C3366 XA.XIR[2].XIC[0].icell.Ien VPWR 0.21079f
C3367 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.04573f
C3368 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02601f
C3369 XA.XIR[13].XIC[8].icell.PDM Vbias 0.03922f
C3370 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.14207f
C3371 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04035f
C3372 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02602f
C3373 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01542f
C3374 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.04573f
C3375 XA.XIR[7].XIC[1].icell.PDM VPWR 0.01373f
C3376 XA.XIR[10].XIC[1].icell.Ien VPWR 0.21079f
C3377 XA.XIR[11].XIC[12].icell.PUM VPWR 0.01079f
C3378 XThR.XTB4.Y a_n997_2667# 0.07199f
C3379 XA.XIR[3].XIC[7].icell.Ien Iout 0.06763f
C3380 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02601f
C3381 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.14207f
C3382 XA.XIR[6].XIC[8].icell.PDM VPWR 0.01373f
C3383 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.14207f
C3384 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.14207f
C3385 XA.XIR[14].XIC[5].icell.PDM VPWR 0.01373f
C3386 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07604f
C3387 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.04573f
C3388 XA.XIR[10].XIC[12].icell.PDM Vbias 0.03922f
C3389 XThR.XTBN.Y XThR.Tn[11] 0.52265f
C3390 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C3391 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C3392 XA.XIR[1].XIC[1].icell.PDM Vbias 0.03922f
C3393 XThC.Tn[11] XThR.Tn[2] 0.39125f
C3394 XA.XIR[13].XIC[9].icell.PDM VPWR 0.01373f
C3395 XA.XIR[6].XIC[10].icell.Ien Vbias 0.19151f
C3396 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.14207f
C3397 XA.XIR[1].XIC[2].icell.Ien Iout 0.06763f
C3398 XThC.XTB7.Y a_10915_9569# 0.06874f
C3399 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C3400 XA.XIR[13].XIC[13].icell.PDM Vbias 0.03922f
C3401 XA.XIR[4].XIC[1].icell.PDM Vbias 0.03922f
C3402 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3403 XA.XIR[8].XIC[10].icell.Ien Iout 0.06763f
C3404 data[5] data[6] 0.01513f
C3405 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.04573f
C3406 XA.XIR[3].XIC[9].icell.PDM Vbias 0.03922f
C3407 XA.XIR[14].XIC[4].icell.Ien Vbias 0.19151f
C3408 XA.XIR[8].XIC[11].icell.PDM Vbias 0.03922f
C3409 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C3410 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C3411 XA.XIR[11].XIC[13].icell.Ien VPWR 0.21079f
C3412 XThR.Tn[7] XThR.Tn[8] 0.114f
C3413 XA.XIR[2].XIC_15.icell.PDM Vbias 0.03927f
C3414 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C3415 XA.XIR[13].XIC[6].icell.Ien Vbias 0.19151f
C3416 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C3417 XA.XIR[3].XIC[6].icell.Ien VPWR 0.21079f
C3418 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.14207f
C3419 XA.XIR[1].XIC[2].icell.PDM VPWR 0.01373f
C3420 XA.XIR[6].XIC[11].icell.PUM VPWR 0.01079f
C3421 XA.XIR[14].XIC[14].icell.PUM VPWR 0.01079f
C3422 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.04573f
C3423 XA.XIR[4].XIC[2].icell.PDM VPWR 0.01373f
C3424 XA.XIR[0].XIC[12].icell.Ien Iout 0.06712f
C3425 XA.XIR[11].XIC[9].icell.Ien Vbias 0.19151f
C3426 XThR.Tn[10] XThR.Tn[11] 0.09883f
C3427 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C3428 XA.XIR[4].XIC_15.icell.Ien VPWR 0.2801f
C3429 XA.XIR[3].XIC[10].icell.PDM VPWR 0.01373f
C3430 XA.XIR[8].XIC[12].icell.PDM VPWR 0.01373f
C3431 XA.XIR[14].XIC[5].icell.PUM VPWR 0.01079f
C3432 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C3433 XThC.Tn[9] XThR.Tn[11] 0.39123f
C3434 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3435 XThC.XTBN.A a_8963_9569# 0.01679f
C3436 XA.XIR[13].XIC[7].icell.PUM VPWR 0.01079f
C3437 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04035f
C3438 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04035f
C3439 XA.XIR[7].XIC_15.icell.Ien Iout 0.0694f
C3440 XA.XIR[8].XIC[9].icell.Ien VPWR 0.21079f
C3441 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02601f
C3442 XA.XIR[5].XIC[0].icell.Ien Iout 0.06763f
C3443 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C3444 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C3445 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C3446 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.02965f
C3447 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C3448 XA.XIR[2].XIC[13].icell.Ien Vbias 0.19151f
C3449 XThC.Tn[14] Iout 0.02232f
C3450 XA.XIR[11].XIC[10].icell.PUM VPWR 0.01079f
C3451 XThC.XTB7.B XThC.Tn[6] 0.04236f
C3452 XThC.XTB5.Y XThC.Tn[10] 0.01755f
C3453 XA.XIR[1].XIC_15.icell.Ien Vbias 0.19199f
C3454 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.04573f
C3455 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.14207f
C3456 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C3457 XA.XIR[0].XIC[11].icell.Ien VPWR 0.2115f
C3458 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.03366f
C3459 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.1155f
C3460 XA.XIR[6].XIC[2].icell.Ien Iout 0.06763f
C3461 XThC.Tn[12] XThR.Tn[1] 0.39128f
C3462 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04023f
C3463 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C3464 bias[1] Vbias 0.68866f
C3465 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C3466 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.04575f
C3467 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.04036f
C3468 XA.XIR[11].XIC[0].icell.PUM VPWR 0.01079f
C3469 XA.XIR[7].XIC[14].icell.Ien VPWR 0.20455f
C3470 XA.XIR[2].XIC[14].icell.PUM VPWR 0.01079f
C3471 XThC.Tn[12] XThR.Tn[12] 0.39123f
C3472 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C3473 XThR.XTB7.A VPWR 0.88654f
C3474 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.14207f
C3475 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.14207f
C3476 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.03822f
C3477 XA.XIR[5].XIC[3].icell.Ien Vbias 0.19151f
C3478 XA.XIR[7].XIC_15.icell.PDM Vbias 0.03927f
C3479 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.0176f
C3480 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02602f
C3481 XA.XIR[11].XIC[11].icell.Ien VPWR 0.21079f
C3482 XThC.XTBN.Y XThC.Tn[10] 0.44415f
C3483 XThC.Tn[7] XThR.Tn[3] 0.39123f
C3484 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C3485 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02601f
C3486 XA.XIR[13].XIC[1].icell.Ien VPWR 0.21079f
C3487 XThC.XTBN.Y a_4861_9615# 0.07601f
C3488 XA.XIR[14].XIC[12].icell.PUM VPWR 0.01079f
C3489 XA.XIR[10].XIC[11].icell.PDM Vbias 0.03922f
C3490 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.0279f
C3491 XThC.Tn[1] XThR.Tn[0] 0.39146f
C3492 XThC.Tn[11] XThR.Tn[10] 0.39123f
C3493 XThC.Tn[3] XThR.Tn[5] 0.39123f
C3494 XA.XIR[10].XIC[3].icell.Ien Iout 0.06763f
C3495 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C3496 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C3497 XThC.XTB5.Y a_5155_10571# 0.01188f
C3498 XA.XIR[9].XIC[11].icell.PDM Vbias 0.03922f
C3499 XA.XIR[13].XIC[12].icell.PDM Vbias 0.03922f
C3500 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.04573f
C3501 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C3502 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C3503 XA.XIR[0].XIC[3].icell.PDM Vbias 0.03922f
C3504 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3505 XA.XIR[5].XIC[4].icell.PUM VPWR 0.01079f
C3506 XA.XIR[3].XIC[12].icell.Ien Iout 0.06763f
C3507 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13586f
C3508 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02601f
C3509 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.14207f
C3510 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.04573f
C3511 XA.XIR[2].XIC[5].icell.Ien Iout 0.06763f
C3512 XA.XIR[11].XIC[14].icell.Ien Vbias 0.19151f
C3513 XThR.Tn[6] Vbias 1.38578f
C3514 XA.XIR[14].XIC[13].icell.Ien VPWR 0.21134f
C3515 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C3516 XA.XIR[6].XIC_15.icell.Ien Vbias 0.19187f
C3517 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.04261f
C3518 XA.XIR[1].XIC[7].icell.Ien Iout 0.06763f
C3519 XA.XIR[9].XIC[12].icell.PDM VPWR 0.01373f
C3520 XA.XIR[0].XIC[4].icell.PDM VPWR 0.01337f
C3521 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C3522 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C3523 XA.XIR[8].XIC_15.icell.Ien Iout 0.0694f
C3524 XA.XIR[1].XIC[1].icell.Ien VPWR 0.21079f
C3525 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C3526 XA.XIR[10].XIC[2].icell.Ien VPWR 0.21079f
C3527 XA.XIR[14].XIC[9].icell.Ien Vbias 0.19151f
C3528 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.04573f
C3529 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C3530 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.04574f
C3531 XThC.Tn[0] XThR.Tn[2] 0.39123f
C3532 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.04573f
C3533 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04035f
C3534 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04035f
C3535 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C3536 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04035f
C3537 XA.XIR[3].XIC[11].icell.Ien VPWR 0.21079f
C3538 XThC.Tn[9] XThR.Tn[14] 0.39123f
C3539 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.14207f
C3540 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.0176f
C3541 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02601f
C3542 XA.XIR[2].XIC[4].icell.Ien VPWR 0.21079f
C3543 XThR.Tn[1] a_n1049_7787# 0.26879f
C3544 XA.XIR[1].XIC[6].icell.Ien VPWR 0.21079f
C3545 XA.XIR[14].XIC[10].icell.PUM VPWR 0.01079f
C3546 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C3547 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C3548 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C3549 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C3550 XA.XIR[8].XIC[14].icell.Ien VPWR 0.20455f
C3551 XA.XIR[5].XIC[1].icell.PDM Vbias 0.03922f
C3552 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.40907f
C3553 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.04f
C3554 XThC.Tn[5] XThR.Tn[6] 0.39123f
C3555 XThR.XTB7.B VPWR 1.67902f
C3556 XThR.Tn[4] Vbias 1.38578f
C3557 XA.XIR[12].XIC[0].icell.PDM Vbias 0.03915f
C3558 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C3559 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C3560 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.04036f
C3561 XThC.Tn[7] XThR.Tn[11] 0.39123f
C3562 XA.XIR[11].XIC[6].icell.PDM Vbias 0.03922f
C3563 XA.XIR[11].XIC[12].icell.Ien Vbias 0.19151f
C3564 XA.XIR[6].XIC[7].icell.Ien Iout 0.06763f
C3565 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04035f
C3566 XA.XIR[14].XIC[11].icell.Ien VPWR 0.21134f
C3567 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.14207f
C3568 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.14207f
C3569 XA.XIR[10].XIC[10].icell.PDM Vbias 0.03922f
C3570 XA.XIR[5].XIC[2].icell.PDM VPWR 0.01373f
C3571 XThC.Tn[3] Iout 0.02217f
C3572 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02601f
C3573 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C3574 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04035f
C3575 XA.XIR[6].XIC[1].icell.Ien VPWR 0.21079f
C3576 XThC.Tn[13] Vbias 0.32423f
C3577 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.04573f
C3578 XA.XIR[13].XIC[11].icell.PDM Vbias 0.03922f
C3579 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.14207f
C3580 XA.XIR[12].XIC[1].icell.PDM VPWR 0.01373f
C3581 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C3582 XA.XIR[5].XIC[8].icell.Ien Vbias 0.19151f
C3583 XThC.Tn[11] XThR.Tn[13] 0.39123f
C3584 XA.XIR[13].XIC[3].icell.Ien Iout 0.06763f
C3585 XThR.Tn[2] VPWR 9.68084f
C3586 XA.XIR[11].XIC[7].icell.PDM VPWR 0.01373f
C3587 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C3588 XThC.Tn[1] XThR.Tn[1] 0.39128f
C3589 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C3590 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.14207f
C3591 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C3592 XThC.Tn[14] XThR.Tn[9] 0.39123f
C3593 XA.XIR[2].XIC[2].icell.PDM Vbias 0.03922f
C3594 XThC.Tn[1] XThR.Tn[12] 0.39123f
C3595 XA.XIR[11].XIC[6].icell.Ien Iout 0.06763f
C3596 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02601f
C3597 XThC.Tn[10] XThR.Tn[8] 0.39123f
C3598 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C3599 XA.XIR[10].XIC[8].icell.Ien Iout 0.06763f
C3600 XA.XIR[12].XIC[3].icell.Ien Vbias 0.19151f
C3601 XA.XIR[6].XIC[6].icell.Ien VPWR 0.21079f
C3602 XA.XIR[14].XIC[14].icell.Ien Vbias 0.19151f
C3603 XA.XIR[5].XIC[9].icell.PUM VPWR 0.01079f
C3604 XThC.XTBN.Y a_7651_9569# 0.23021f
C3605 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C3606 XThC.Tn[5] XThR.Tn[4] 0.39123f
C3607 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C3608 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.13934f
C3609 XThC.XTB4.Y XThC.Tn[3] 0.1917f
C3610 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.14207f
C3611 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.14207f
C3612 XThC.Tn[0] XThR.Tn[10] 0.39118f
C3613 XA.XIR[2].XIC[3].icell.PDM VPWR 0.01373f
C3614 XA.XIR[13].XIC[2].icell.Ien VPWR 0.21079f
C3615 XA.XIR[2].XIC[10].icell.Ien Iout 0.06763f
C3616 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C3617 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.04573f
C3618 XThR.Tn[13] XThR.Tn[14] 0.19422f
C3619 XA.XIR[1].XIC[12].icell.Ien Iout 0.06763f
C3620 XA.XIR[12].XIC[4].icell.PUM VPWR 0.01079f
C3621 XA.XIR[11].XIC[5].icell.Ien VPWR 0.21079f
C3622 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04035f
C3623 XA.XIR[11].XIC[10].icell.Ien Vbias 0.19151f
C3624 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.14207f
C3625 XA.XIR[10].XIC[7].icell.Ien VPWR 0.21079f
C3626 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C3627 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C3628 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C3629 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.36378f
C3630 XThC.XTB2.Y a_4067_9615# 0.02133f
C3631 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C3632 XThC.XTBN.A Vbias 0.01693f
C3633 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02601f
C3634 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C3635 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C3636 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04035f
C3637 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3638 XThR.XTBN.Y VPWR 4.58541f
C3639 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.0404f
C3640 XA.XIR[2].XIC[9].icell.Ien VPWR 0.21079f
C3641 XA.XIR[11].XIC[0].icell.Ien Vbias 0.19149f
C3642 XA.XIR[1].XIC[11].icell.Ien VPWR 0.21079f
C3643 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C3644 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.14207f
C3645 XA.XIR[7].XIC[2].icell.PDM Vbias 0.03922f
C3646 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04035f
C3647 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C3648 XA.XIR[6].XIC[9].icell.PDM Vbias 0.03922f
C3649 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.04573f
C3650 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C3651 XA.XIR[15].XIC[0].icell.PDM Vbias 0.03915f
C3652 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02601f
C3653 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C3654 XThC.Tn[7] XThR.Tn[14] 0.39123f
C3655 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.14207f
C3656 XA.XIR[14].XIC[6].icell.PDM Vbias 0.03922f
C3657 XA.XIR[14].XIC[12].icell.Ien Vbias 0.19151f
C3658 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02601f
C3659 a_10051_9569# XThC.Tn[13] 0.1927f
C3660 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C3661 XThR.XTB4.Y VPWR 0.92877f
C3662 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04023f
C3663 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C3664 XA.XIR[12].XIC[13].icell.Ien Iout 0.06763f
C3665 XA.XIR[13].XIC[10].icell.PDM Vbias 0.03922f
C3666 XA.XIR[11].XIC[1].icell.PUM VPWR 0.01079f
C3667 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.14207f
C3668 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04035f
C3669 XThR.Tn[10] VPWR 10.5778f
C3670 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13586f
C3671 XA.XIR[7].XIC[3].icell.PDM VPWR 0.01373f
C3672 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01542f
C3673 XA.XIR[9].XIC[4].icell.Ien Vbias 0.19151f
C3674 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01714f
C3675 XA.XIR[6].XIC[10].icell.PDM VPWR 0.01373f
C3676 XA.XIR[6].XIC[12].icell.Ien Iout 0.06763f
C3677 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C3678 XThC.Tn[9] VPWR 7.96526f
C3679 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02602f
C3680 XThR.XTB5.A a_n1335_4229# 0.01243f
C3681 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.14207f
C3682 XA.XIR[14].XIC[7].icell.PDM VPWR 0.01373f
C3683 XA.XIR[1].XIC[3].icell.PDM Vbias 0.03922f
C3684 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02601f
C3685 XA.XIR[14].XIC[6].icell.Ien Iout 0.06763f
C3686 XA.XIR[4].XIC[3].icell.PDM Vbias 0.03922f
C3687 XA.XIR[5].XIC[13].icell.Ien Vbias 0.19151f
C3688 XA.XIR[13].XIC[8].icell.Ien Iout 0.06763f
C3689 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C3690 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C3691 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C3692 XA.XIR[9].XIC[5].icell.PUM VPWR 0.01079f
C3693 XThC.XTB3.Y Vbias 0.01224f
C3694 XA.XIR[8].XIC[13].icell.PDM Vbias 0.03922f
C3695 XA.XIR[3].XIC[11].icell.PDM Vbias 0.03922f
C3696 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C3697 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C3698 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C3699 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02601f
C3700 XThC.Tn[2] Vbias 0.32256f
C3701 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.04573f
C3702 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C3703 XA.XIR[11].XIC_15.icell.PDM Vbias 0.03927f
C3704 XA.XIR[1].XIC[4].icell.PDM VPWR 0.01373f
C3705 XA.XIR[11].XIC_15.icell.Ien Vbias 0.19187f
C3706 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C3707 XThC.Tn[0] XThR.Tn[13] 0.39121f
C3708 XA.XIR[12].XIC[8].icell.Ien Vbias 0.19151f
C3709 XA.XIR[6].XIC[11].icell.Ien VPWR 0.21079f
C3710 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C3711 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C3712 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.04574f
C3713 XA.XIR[4].XIC[4].icell.PDM VPWR 0.01373f
C3714 XA.XIR[5].XIC[14].icell.PUM VPWR 0.01079f
C3715 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04035f
C3716 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C3717 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C3718 XThC.Tn[3] XThR.Tn[9] 0.39123f
C3719 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C3720 XA.XIR[8].XIC[14].icell.PDM VPWR 0.01349f
C3721 XA.XIR[3].XIC[12].icell.PDM VPWR 0.01373f
C3722 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C3723 XA.XIR[14].XIC[5].icell.Ien VPWR 0.21134f
C3724 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C3725 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.14207f
C3726 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.04628f
C3727 XA.XIR[14].XIC[10].icell.Ien Vbias 0.19151f
C3728 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C3729 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02602f
C3730 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04035f
C3731 XA.XIR[2].XIC_15.icell.Ien Iout 0.0694f
C3732 XA.XIR[13].XIC[7].icell.Ien VPWR 0.21079f
C3733 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04035f
C3734 XThR.XTB6.A XThR.XTBN.A 0.0512f
C3735 XA.XIR[12].XIC[11].icell.Ien Iout 0.06763f
C3736 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3737 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.0176f
C3738 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02601f
C3739 XA.XIR[12].XIC[9].icell.PUM VPWR 0.01079f
C3740 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C3741 XThR.XTB7.Y a_n997_1579# 0.013f
C3742 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02601f
C3743 a_n997_1803# VPWR 0.02096f
C3744 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02792f
C3745 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.04261f
C3746 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01244f
C3747 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.0404f
C3748 XA.XIR[4].XIC[1].icell.Ien Vbias 0.19151f
C3749 XA.XIR[8].XIC[0].icell.PUM VPWR 0.01079f
C3750 XThC.XTB7.A a_4861_9615# 0.02294f
C3751 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02601f
C3752 XThC.Tn[3] XThC.Tn[4] 0.45991f
C3753 XA.XIR[5].XIC[5].icell.Ien Iout 0.06763f
C3754 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C3755 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02601f
C3756 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.04036f
C3757 XA.XIR[2].XIC[14].icell.Ien VPWR 0.20455f
C3758 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C3759 XThC.XTB1.Y Vbias 0.01575f
C3760 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C3761 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02601f
C3762 XA.XIR[15].XIC[3].icell.Ien Vbias 0.15955f
C3763 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.14207f
C3764 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C3765 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C3766 XA.XIR[14].XIC[0].icell.Ien VPWR 0.21134f
C3767 XA.XIR[4].XIC[2].icell.PUM VPWR 0.01079f
C3768 XA.XIR[4].XIC[6].icell.Ien Vbias 0.19151f
C3769 XThR.Tn[13] VPWR 10.6686f
C3770 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C3771 XThR.Tn[5] Iout 1.10104f
C3772 data[1] data[2] 0.01393f
C3773 XThR.Tn[8] data[4] 0.01643f
C3774 XThC.XTBN.Y a_5949_9615# 0.07703f
C3775 XThC.Tn[11] XThR.Tn[7] 0.39123f
C3776 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.04573f
C3777 XThC.XTB7.B XThC.Tn[9] 0.05138f
C3778 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C3779 XThR.XTBN.A data[7] 0.07741f
C3780 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C3781 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C3782 XThC.XTB7.Y XThC.Tn[13] 0.10845f
C3783 XA.XIR[9].XIC[13].icell.PDM Vbias 0.03922f
C3784 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.14207f
C3785 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C3786 XA.XIR[0].XIC[5].icell.PDM Vbias 0.03922f
C3787 XA.XIR[7].XIC[0].icell.Ien Vbias 0.19149f
C3788 XA.XIR[15].XIC[4].icell.PUM VPWR 0.01079f
C3789 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.14207f
C3790 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02601f
C3791 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.04573f
C3792 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02601f
C3793 XA.XIR[5].XIC[4].icell.Ien VPWR 0.21079f
C3794 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C3795 XA.XIR[9].XIC[9].icell.Ien Vbias 0.19151f
C3796 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C3797 XThR.Tn[3] a_n1049_6699# 0.27008f
C3798 XA.XIR[4].XIC[7].icell.PUM VPWR 0.01079f
C3799 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13586f
C3800 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C3801 XA.XIR[0].XIC[2].icell.Ien Vbias 0.19186f
C3802 XA.XIR[11].XIC[14].icell.PDM Vbias 0.03922f
C3803 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02601f
C3804 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C3805 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C3806 XA.XIR[9].XIC[14].icell.PDM VPWR 0.01349f
C3807 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C3808 XA.XIR[0].XIC[6].icell.PDM VPWR 0.0134f
C3809 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C3810 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C3811 XA.XIR[7].XIC[1].icell.PUM VPWR 0.01079f
C3812 XThC.Tn[10] XThR.Tn[3] 0.39123f
C3813 XA.XIR[14].XIC_15.icell.PDM Vbias 0.03927f
C3814 XA.XIR[14].XIC_15.icell.Ien Vbias 0.19187f
C3815 XA.XIR[7].XIC[5].icell.Ien Vbias 0.19151f
C3816 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.13232f
C3817 XA.XIR[9].XIC[10].icell.PUM VPWR 0.01079f
C3818 XThC.Tn[7] VPWR 7.39928f
C3819 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C3820 XA.XIR[0].XIC[3].icell.PUM VPWR 0.01038f
C3821 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04035f
C3822 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04035f
C3823 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.04036f
C3824 XThC.Tn[13] XThR.Tn[0] 0.39146f
C3825 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C3826 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C3827 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C3828 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02601f
C3829 XA.XIR[7].XIC[6].icell.PUM VPWR 0.01079f
C3830 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.0176f
C3831 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.04573f
C3832 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C3833 XA.XIR[15].XIC[13].icell.Ien Iout 0.07153f
C3834 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C3835 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02803f
C3836 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C3837 a_2979_9615# Vbias 0.01329f
C3838 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01263f
C3839 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.4095f
C3840 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02601f
C3841 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C3842 XA.XIR[5].XIC[3].icell.PDM Vbias 0.03922f
C3843 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04035f
C3844 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.14207f
C3845 XThR.XTB5.A data[5] 0.11096f
C3846 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.04573f
C3847 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C3848 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02601f
C3849 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C3850 XA.XIR[5].XIC[0].icell.PUM VPWR 0.01079f
C3851 XThR.XTBN.A XThR.Tn[12] 0.22096f
C3852 XA.XIR[12].XIC[2].icell.PDM Vbias 0.03922f
C3853 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C3854 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.04573f
C3855 a_3773_9615# VPWR 0.70508f
C3856 XA.XIR[11].XIC[8].icell.PDM Vbias 0.03922f
C3857 XThR.XTB2.Y a_n997_3755# 0.06476f
C3858 XThC.Tn[12] XThR.Tn[2] 0.39125f
C3859 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C3860 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04035f
C3861 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C3862 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.02965f
C3863 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C3864 XA.XIR[5].XIC[4].icell.PDM VPWR 0.01373f
C3865 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C3866 XA.XIR[5].XIC[10].icell.Ien Iout 0.06763f
C3867 XThC.XTB4.Y a_5155_9615# 0.01546f
C3868 XThR.XTBN.Y a_n1049_8581# 0.0607f
C3869 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13586f
C3870 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C3871 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04023f
C3872 XA.XIR[3].XIC[2].icell.Ien Vbias 0.19151f
C3873 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.13192f
C3874 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C3875 XA.XIR[12].XIC[3].icell.PDM VPWR 0.01373f
C3876 XA.XIR[15].XIC[8].icell.Ien Vbias 0.15955f
C3877 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C3878 XA.XIR[11].XIC[9].icell.PDM VPWR 0.01373f
C3879 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02601f
C3880 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C3881 XA.XIR[8].XIC[0].icell.PDM Vbias 0.03915f
C3882 XA.XIR[4].XIC[11].icell.Ien Vbias 0.19151f
C3883 XA.XIR[12].XIC[5].icell.Ien Iout 0.06763f
C3884 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.04573f
C3885 XA.XIR[11].XIC[13].icell.PDM Vbias 0.03922f
C3886 XA.XIR[2].XIC[4].icell.PDM Vbias 0.03922f
C3887 XThC.Tn[8] XThR.Tn[6] 0.39123f
C3888 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.04573f
C3889 XA.XIR[8].XIC[5].icell.Ien Vbias 0.19151f
C3890 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04035f
C3891 XA.XIR[3].XIC[3].icell.PUM VPWR 0.01079f
C3892 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.04629f
C3893 XA.XIR[15].XIC[11].icell.Ien Iout 0.07153f
C3894 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13586f
C3895 XA.XIR[14].XIC[14].icell.PDM Vbias 0.03922f
C3896 XThR.XTB3.Y a_n997_2891# 0.07285f
C3897 XThC.Tn[10] XThR.Tn[11] 0.39123f
C3898 XA.XIR[15].XIC[9].icell.PUM VPWR 0.01079f
C3899 XA.XIR[5].XIC[9].icell.Ien VPWR 0.21079f
C3900 XThC.XTBN.Y a_8739_9569# 0.22804f
C3901 XA.XIR[9].XIC[14].icell.Ien Vbias 0.19151f
C3902 XThC.Tn[0] XThR.Tn[7] 0.39119f
C3903 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.14207f
C3904 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.04573f
C3905 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C3906 XA.XIR[4].XIC[12].icell.PUM VPWR 0.01079f
C3907 XA.XIR[8].XIC[1].icell.PDM VPWR 0.01373f
C3908 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C3909 a_n1049_5317# XThR.Tn[6] 0.26047f
C3910 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.14207f
C3911 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.14207f
C3912 XA.XIR[0].XIC[7].icell.Ien Vbias 0.19186f
C3913 XA.XIR[2].XIC[5].icell.PDM VPWR 0.01373f
C3914 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C3915 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C3916 XThC.XTB7.B XThC.Tn[7] 0.07144f
C3917 XA.XIR[8].XIC[6].icell.PUM VPWR 0.01079f
C3918 XThC.XTB5.Y XThC.Tn[11] 0.02112f
C3919 XA.XIR[12].XIC[4].icell.Ien VPWR 0.21079f
C3920 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C3921 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C3922 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C3923 a_8739_9569# XThC.Tn[10] 0.21014f
C3924 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C3925 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04035f
C3926 a_n997_3979# VPWR 0.01765f
C3927 XA.XIR[7].XIC[10].icell.Ien Vbias 0.19151f
C3928 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.04575f
C3929 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.03942f
C3930 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01768f
C3931 XThC.Tn[13] XThR.Tn[1] 0.39128f
C3932 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.14207f
C3933 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01687f
C3934 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.04573f
C3935 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C3936 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C3937 XA.XIR[0].XIC[8].icell.PUM VPWR 0.01039f
C3938 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C3939 XThC.Tn[13] XThR.Tn[12] 0.39123f
C3940 XA.XIR[8].XIC[0].icell.Ien Vbias 0.19149f
C3941 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04035f
C3942 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C3943 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04035f
C3944 XThC.XTB6.A XThC.XTBN.A 0.0513f
C3945 XA.XIR[9].XIC[1].icell.Ien Iout 0.06763f
C3946 XThC.XTBN.Y XThC.Tn[11] 0.39675f
C3947 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02602f
C3948 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.04573f
C3949 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04035f
C3950 XThC.Tn[8] XThR.Tn[4] 0.39123f
C3951 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.40932f
C3952 XA.XIR[7].XIC[11].icell.PUM VPWR 0.01079f
C3953 XA.XIR[4].XIC[3].icell.Ien Iout 0.06763f
C3954 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02601f
C3955 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04035f
C3956 XA.XIR[7].XIC[4].icell.PDM Vbias 0.03922f
C3957 XThC.Tn[2] XThR.Tn[0] 0.39148f
C3958 XThC.Tn[12] XThR.Tn[10] 0.39123f
C3959 XA.XIR[15].XIC[2].icell.PDM Vbias 0.03922f
C3960 XA.XIR[6].XIC[11].icell.PDM Vbias 0.03922f
C3961 XThC.Tn[4] XThR.Tn[5] 0.39123f
C3962 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.14207f
C3963 XA.XIR[8].XIC[1].icell.PUM VPWR 0.01079f
C3964 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.14207f
C3965 XA.XIR[14].XIC[8].icell.PDM Vbias 0.03922f
C3966 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C3967 XThC.Tn[10] XThC.Tn[11] 0.07237f
C3968 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02601f
C3969 XA.XIR[9].XIC[6].icell.Ien Iout 0.06763f
C3970 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.02965f
C3971 XThR.Tn[7] VPWR 10.0243f
C3972 a_n997_2891# VPWR 0.01421f
C3973 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04035f
C3974 XA.XIR[9].XIC[0].icell.PDM Vbias 0.03915f
C3975 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.04573f
C3976 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C3977 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C3978 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.04573f
C3979 XA.XIR[7].XIC[5].icell.PDM VPWR 0.01373f
C3980 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.14207f
C3981 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C3982 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01714f
C3983 XA.XIR[4].XIC[2].icell.Ien VPWR 0.21079f
C3984 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C3985 XA.XIR[6].XIC[12].icell.PDM VPWR 0.01373f
C3986 XThR.XTB6.Y a_n1049_5317# 0.01199f
C3987 XA.XIR[11].XIC[12].icell.PDM Vbias 0.03922f
C3988 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.04573f
C3989 XA.XIR[14].XIC[9].icell.PDM VPWR 0.01373f
C3990 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C3991 XA.XIR[5].XIC_15.icell.Ien Iout 0.0694f
C3992 XA.XIR[7].XIC[2].icell.Ien Iout 0.06763f
C3993 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.04573f
C3994 XA.XIR[3].XIC[7].icell.Ien Vbias 0.19151f
C3995 XA.XIR[1].XIC[5].icell.PDM Vbias 0.03922f
C3996 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C3997 XA.XIR[14].XIC[13].icell.PDM Vbias 0.03922f
C3998 XA.XIR[9].XIC[1].icell.PDM VPWR 0.01373f
C3999 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02601f
C4000 XThC.Tn[1] XThR.Tn[2] 0.39125f
C4001 XA.XIR[4].XIC[5].icell.PDM Vbias 0.03922f
C4002 XA.XIR[9].XIC[5].icell.Ien VPWR 0.21079f
C4003 XA.XIR[1].XIC[2].icell.Ien Vbias 0.19162f
C4004 XThC.Tn[10] XThR.Tn[14] 0.39123f
C4005 XA.XIR[8].XIC_15.icell.PDM Vbias 0.03927f
C4006 XA.XIR[3].XIC[13].icell.PDM Vbias 0.03922f
C4007 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C4008 XThR.XTBN.Y a_n1049_7787# 0.08456f
C4009 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C4010 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02601f
C4011 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C4012 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.0404f
C4013 XA.XIR[8].XIC[10].icell.Ien Vbias 0.19151f
C4014 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C4015 XA.XIR[3].XIC[8].icell.PUM VPWR 0.01079f
C4016 XA.XIR[1].XIC[6].icell.PDM VPWR 0.01373f
C4017 XThR.Tn[9] Iout 1.10103f
C4018 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02601f
C4019 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C4020 a_n1049_6405# XThR.Tn[4] 0.26564f
C4021 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C4022 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.14207f
C4023 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01687f
C4024 a_5155_9615# XThC.Tn[4] 0.27224f
C4025 XA.XIR[4].XIC[6].icell.PDM VPWR 0.01373f
C4026 XA.XIR[5].XIC[14].icell.Ien VPWR 0.20455f
C4027 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04035f
C4028 XA.XIR[1].XIC[3].icell.PUM VPWR 0.01079f
C4029 XA.XIR[3].XIC[14].icell.PDM VPWR 0.01349f
C4030 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C4031 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C4032 XThC.Tn[6] XThR.Tn[6] 0.39123f
C4033 XThC.XTBN.A XThC.Tn[8] 0.13691f
C4034 XA.XIR[0].XIC[12].icell.Ien Vbias 0.19186f
C4035 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01768f
C4036 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04035f
C4037 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04035f
C4038 XA.XIR[8].XIC[11].icell.PUM VPWR 0.01079f
C4039 XA.XIR[15].XIC[0].icell.Ien Iout 0.07153f
C4040 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C4041 XA.XIR[12].XIC[9].icell.Ien VPWR 0.21079f
C4042 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01687f
C4043 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02602f
C4044 XA.XIR[7].XIC_15.icell.Ien Vbias 0.19187f
C4045 XA.XIR[5].XIC[0].icell.Ien Vbias 0.19149f
C4046 XA.XIR[9].XIC[0].icell.Ien VPWR 0.21079f
C4047 XThC.Tn[4] Iout 0.02297f
C4048 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C4049 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.14207f
C4050 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02601f
C4051 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04035f
C4052 XA.XIR[0].XIC[13].icell.PUM VPWR 0.01038f
C4053 XThC.Tn[14] Vbias 0.33142f
C4054 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02601f
C4055 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.14207f
C4056 XThC.XTB7.A a_5949_9615# 0.01824f
C4057 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.04573f
C4058 XA.XIR[15].XIC[5].icell.Ien Iout 0.07153f
C4059 XThC.Tn[12] XThR.Tn[13] 0.39123f
C4060 XThC.Tn[2] XThR.Tn[1] 0.39128f
C4061 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04035f
C4062 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C4063 XA.XIR[6].XIC[2].icell.Ien Vbias 0.19151f
C4064 XA.XIR[4].XIC[8].icell.Ien Iout 0.06763f
C4065 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02601f
C4066 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.14207f
C4067 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.0176f
C4068 XA.XIR[5].XIC[1].icell.PUM VPWR 0.01079f
C4069 XThC.XTB2.Y a_7875_9569# 0.06476f
C4070 XThC.Tn[2] XThR.Tn[12] 0.39123f
C4071 XThC.XTB5.A XThC.XTB7.A 0.07824f
C4072 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C4073 a_n997_1579# VPWR 0.02465f
C4074 XThC.Tn[11] XThR.Tn[8] 0.39123f
C4075 XA.XIR[8].XIC[2].icell.Ien Iout 0.06763f
C4076 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C4077 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.04573f
C4078 XA.XIR[11].XIC[11].icell.PDM Vbias 0.03922f
C4079 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C4080 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.14207f
C4081 XThC.XTBN.Y XThC.Tn[0] 0.45269f
C4082 XA.XIR[10].XIC[0].icell.PDM VPWR 0.01373f
C4083 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C4084 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.04261f
C4085 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.14207f
C4086 XThC.Tn[6] XThR.Tn[4] 0.39123f
C4087 XA.XIR[9].XIC[11].icell.Ien Iout 0.06763f
C4088 XA.XIR[14].XIC[12].icell.PDM Vbias 0.03922f
C4089 XA.XIR[6].XIC[3].icell.PUM VPWR 0.01079f
C4090 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C4091 XA.XIR[9].XIC_15.icell.PDM Vbias 0.03927f
C4092 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C4093 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.04573f
C4094 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C4095 XA.XIR[15].XIC[4].icell.Ien VPWR 0.3396f
C4096 XA.XIR[0].XIC[7].icell.PDM Vbias 0.03922f
C4097 XThC.XTB2.Y data[1] 0.017f
C4098 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02601f
C4099 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.04573f
C4100 XA.XIR[0].XIC[4].icell.Ien Iout 0.06712f
C4101 XThC.Tn[1] XThR.Tn[10] 0.39123f
C4102 XA.XIR[12].XIC[13].icell.PUM VPWR 0.01079f
C4103 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.14207f
C4104 XA.XIR[10].XIC[3].icell.Ien Vbias 0.19151f
C4105 XA.XIR[4].XIC[7].icell.Ien VPWR 0.21079f
C4106 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02601f
C4107 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.14207f
C4108 XThR.XTB7.Y a_n997_715# 0.06874f
C4109 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02803f
C4110 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.04575f
C4111 XA.XIR[7].XIC[7].icell.Ien Iout 0.06763f
C4112 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02601f
C4113 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.04573f
C4114 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02601f
C4115 XA.XIR[3].XIC[12].icell.Ien Vbias 0.19151f
C4116 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C4117 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C4118 XA.XIR[7].XIC[1].icell.Ien VPWR 0.21079f
C4119 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01653f
C4120 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.14207f
C4121 XA.XIR[2].XIC[5].icell.Ien Vbias 0.19151f
C4122 XThC.XTB5.Y VPWR 1.01219f
C4123 XThC.XTBN.A data[3] 0.07741f
C4124 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02601f
C4125 XA.XIR[9].XIC[10].icell.Ien VPWR 0.21079f
C4126 XA.XIR[1].XIC[7].icell.Ien Vbias 0.19162f
C4127 XThC.XTB7.A data[0] 0.86893f
C4128 XA.XIR[10].XIC[4].icell.PUM VPWR 0.01079f
C4129 XA.XIR[12].XIC[14].icell.Ien VPWR 0.20455f
C4130 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C4131 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.14207f
C4132 XA.XIR[0].XIC[3].icell.Ien VPWR 0.21044f
C4133 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04035f
C4134 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04035f
C4135 XA.XIR[8].XIC_15.icell.Ien Vbias 0.19187f
C4136 XA.XIR[3].XIC[13].icell.PUM VPWR 0.01079f
C4137 XA.XIR[2].XIC[6].icell.PUM VPWR 0.01079f
C4138 XA.XIR[7].XIC[6].icell.Ien VPWR 0.21079f
C4139 XThC.XTBN.Y VPWR 4.08404f
C4140 XA.XIR[1].XIC[8].icell.PUM VPWR 0.01079f
C4141 XThC.XTB6.Y a_6243_9615# 0.01199f
C4142 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.04573f
C4143 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C4144 a_n1049_6699# VPWR 0.72212f
C4145 XThR.XTB7.A XThR.XTBN.A 0.19736f
C4146 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C4147 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02601f
C4148 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.0176f
C4149 XA.XIR[5].XIC[5].icell.PDM Vbias 0.03922f
C4150 XThR.XTB7.A XThR.Tn[6] 0.10551f
C4151 XA.XIR[12].XIC[11].icell.PUM VPWR 0.01079f
C4152 XThC.XTB1.Y XThC.Tn[8] 0.29214f
C4153 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.14207f
C4154 XThC.Tn[10] VPWR 7.96973f
C4155 XA.XIR[12].XIC[4].icell.PDM Vbias 0.03922f
C4156 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.04574f
C4157 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.04573f
C4158 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13586f
C4159 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.04573f
C4160 XA.XIR[10].XIC[13].icell.Ien Iout 0.06763f
C4161 XA.XIR[11].XIC[10].icell.PDM Vbias 0.03922f
C4162 a_4861_9615# VPWR 0.70519f
C4163 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.14207f
C4164 XA.XIR[3].XIC[4].icell.Ien Iout 0.06763f
C4165 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.14207f
C4166 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08254f
C4167 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04035f
C4168 XA.XIR[5].XIC[6].icell.PDM VPWR 0.01373f
C4169 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.04573f
C4170 XA.XIR[14].XIC[11].icell.PDM Vbias 0.03922f
C4171 XA.XIR[13].XIC[0].icell.PDM VPWR 0.01373f
C4172 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.14207f
C4173 XA.XIR[4].XIC[13].icell.Ien Iout 0.06763f
C4174 XA.XIR[6].XIC[7].icell.Ien Vbias 0.19151f
C4175 XThC.XTB5.A data[0] 0.14415f
C4176 XThC.XTB5.Y a_9827_9569# 0.06458f
C4177 XA.XIR[12].XIC[5].icell.PDM VPWR 0.01373f
C4178 XThC.Tn[3] Vbias 0.33184f
C4179 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C4180 XA.XIR[12].XIC[12].icell.Ien VPWR 0.21079f
C4181 XA.XIR[8].XIC[7].icell.Ien Iout 0.06763f
C4182 XA.XIR[3].XIC[0].icell.PDM Vbias 0.03915f
C4183 XA.XIR[8].XIC[2].icell.PDM Vbias 0.03922f
C4184 XThC.Tn[1] XThR.Tn[13] 0.39123f
C4185 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02601f
C4186 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.04573f
C4187 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C4188 XA.XIR[2].XIC[6].icell.PDM Vbias 0.03922f
C4189 data[7] VGND 0.49949f
C4190 data[6] VGND 0.47974f
C4191 data[4] VGND 0.59315f
C4192 data[5] VGND 1.17814f
C4193 Iout VGND 0.32144p
C4194 data[3] VGND 0.49963f
C4195 data[2] VGND 0.48064f
C4196 data[0] VGND 0.59271f
C4197 data[1] VGND 1.17844f
C4198 Vbias VGND 0.17693p
C4199 bias[0] VGND 1.39569f
C4200 bias[1] VGND 0.46888f
C4201 bias[2] VGND 0.40015f
C4202 VPWR VGND 0.42118p
C4203 a_n997_715# VGND 0.5638f
C4204 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C4205 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C4206 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64463f
C4207 XA.XIR[15].XIC_15.icell.Ien VGND 0.44415f
C4208 XA.XIR[15].XIC[14].icell.Ien VGND 0.44309f
C4209 XA.XIR[15].XIC[13].icell.Ien VGND 0.44309f
C4210 XA.XIR[15].XIC[12].icell.Ien VGND 0.44309f
C4211 XA.XIR[15].XIC[11].icell.Ien VGND 0.44309f
C4212 XA.XIR[15].XIC[10].icell.Ien VGND 0.44309f
C4213 XA.XIR[15].XIC[9].icell.Ien VGND 0.44309f
C4214 XA.XIR[15].XIC[8].icell.Ien VGND 0.44309f
C4215 XA.XIR[15].XIC[7].icell.Ien VGND 0.44309f
C4216 XA.XIR[15].XIC[6].icell.Ien VGND 0.44309f
C4217 XA.XIR[15].XIC[5].icell.Ien VGND 0.44309f
C4218 XA.XIR[15].XIC[4].icell.Ien VGND 0.44309f
C4219 XA.XIR[15].XIC[3].icell.Ien VGND 0.44309f
C4220 XA.XIR[15].XIC[2].icell.Ien VGND 0.44309f
C4221 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70493f
C4222 XA.XIR[15].XIC[1].icell.Ien VGND 0.44309f
C4223 XA.XIR[15].XIC[0].icell.Ien VGND 0.44311f
C4224 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01013f
C4225 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.6116f
C4226 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C4227 XA.XIR[15].XIC_15.icell.PDM VGND 0.18773f
C4228 XA.XIR[15].XIC[14].icell.PDM VGND 0.18726f
C4229 XA.XIR[15].XIC[13].icell.PDM VGND 0.18726f
C4230 XA.XIR[15].XIC[12].icell.PDM VGND 0.18726f
C4231 XA.XIR[15].XIC[11].icell.PDM VGND 0.18726f
C4232 XA.XIR[15].XIC[10].icell.PDM VGND 0.18726f
C4233 XA.XIR[15].XIC[9].icell.PDM VGND 0.18726f
C4234 XA.XIR[15].XIC[8].icell.PDM VGND 0.18726f
C4235 XA.XIR[15].XIC[7].icell.PDM VGND 0.18726f
C4236 XA.XIR[15].XIC[6].icell.PDM VGND 0.18726f
C4237 XA.XIR[15].XIC[5].icell.PDM VGND 0.18726f
C4238 XA.XIR[15].XIC[4].icell.PDM VGND 0.18726f
C4239 XA.XIR[15].XIC[3].icell.PDM VGND 0.18726f
C4240 XA.XIR[15].XIC[2].icell.PDM VGND 0.18726f
C4241 XA.XIR[15].XIC[1].icell.PDM VGND 0.18726f
C4242 XA.XIR[15].XIC[0].icell.PDM VGND 0.18734f
C4243 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C4244 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C4245 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C4246 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60749f
C4247 XA.XIR[14].XIC_15.icell.Ien VGND 0.37186f
C4248 XA.XIR[14].XIC[14].icell.Ien VGND 0.37133f
C4249 XA.XIR[14].XIC[13].icell.Ien VGND 0.37133f
C4250 XA.XIR[14].XIC[12].icell.Ien VGND 0.37133f
C4251 XA.XIR[14].XIC[11].icell.Ien VGND 0.37133f
C4252 XA.XIR[14].XIC[10].icell.Ien VGND 0.37133f
C4253 XA.XIR[14].XIC[9].icell.Ien VGND 0.37133f
C4254 XA.XIR[14].XIC[8].icell.Ien VGND 0.37133f
C4255 XA.XIR[14].XIC[7].icell.Ien VGND 0.37133f
C4256 XA.XIR[14].XIC[6].icell.Ien VGND 0.37133f
C4257 XA.XIR[14].XIC[5].icell.Ien VGND 0.37133f
C4258 XA.XIR[14].XIC[4].icell.Ien VGND 0.37133f
C4259 XA.XIR[14].XIC[3].icell.Ien VGND 0.37133f
C4260 XA.XIR[14].XIC[2].icell.Ien VGND 0.37133f
C4261 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.80471f
C4262 XThR.Tn[14] VGND 13.61789f
C4263 XA.XIR[14].XIC[1].icell.Ien VGND 0.37133f
C4264 a_n997_1579# VGND 0.54776f
C4265 XA.XIR[14].XIC[0].icell.Ien VGND 0.37135f
C4266 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01013f
C4267 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.5751f
C4268 a_n997_1803# VGND 0.53619f
C4269 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C4270 XA.XIR[14].XIC_15.icell.PDM VGND 0.18849f
C4271 XA.XIR[14].XIC[14].icell.PDM VGND 0.18803f
C4272 XA.XIR[14].XIC[13].icell.PDM VGND 0.18803f
C4273 XA.XIR[14].XIC[12].icell.PDM VGND 0.18803f
C4274 XA.XIR[14].XIC[11].icell.PDM VGND 0.18803f
C4275 XA.XIR[14].XIC[10].icell.PDM VGND 0.18803f
C4276 XA.XIR[14].XIC[9].icell.PDM VGND 0.18803f
C4277 XA.XIR[14].XIC[8].icell.PDM VGND 0.18803f
C4278 XA.XIR[14].XIC[7].icell.PDM VGND 0.18803f
C4279 XA.XIR[14].XIC[6].icell.PDM VGND 0.18803f
C4280 XA.XIR[14].XIC[5].icell.PDM VGND 0.18803f
C4281 XA.XIR[14].XIC[4].icell.PDM VGND 0.18803f
C4282 XA.XIR[14].XIC[3].icell.PDM VGND 0.18803f
C4283 XA.XIR[14].XIC[2].icell.PDM VGND 0.18803f
C4284 XA.XIR[14].XIC[1].icell.PDM VGND 0.18803f
C4285 XA.XIR[14].XIC[0].icell.PDM VGND 0.1881f
C4286 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C4287 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C4288 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C4289 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60749f
C4290 XA.XIR[13].XIC_15.icell.Ien VGND 0.37186f
C4291 XA.XIR[13].XIC[14].icell.Ien VGND 0.37133f
C4292 XA.XIR[13].XIC[13].icell.Ien VGND 0.37133f
C4293 XA.XIR[13].XIC[12].icell.Ien VGND 0.37133f
C4294 XA.XIR[13].XIC[11].icell.Ien VGND 0.37133f
C4295 XA.XIR[13].XIC[10].icell.Ien VGND 0.37133f
C4296 XA.XIR[13].XIC[9].icell.Ien VGND 0.37133f
C4297 XA.XIR[13].XIC[8].icell.Ien VGND 0.37133f
C4298 XA.XIR[13].XIC[7].icell.Ien VGND 0.37133f
C4299 XA.XIR[13].XIC[6].icell.Ien VGND 0.37133f
C4300 XA.XIR[13].XIC[5].icell.Ien VGND 0.37133f
C4301 XA.XIR[13].XIC[4].icell.Ien VGND 0.37133f
C4302 XA.XIR[13].XIC[3].icell.Ien VGND 0.37133f
C4303 XA.XIR[13].XIC[2].icell.Ien VGND 0.37133f
C4304 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.80475f
C4305 XThR.Tn[13] VGND 13.49599f
C4306 XA.XIR[13].XIC[1].icell.Ien VGND 0.37133f
C4307 XA.XIR[13].XIC[0].icell.Ien VGND 0.37135f
C4308 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01013f
C4309 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57422f
C4310 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C4311 XA.XIR[13].XIC_15.icell.PDM VGND 0.18849f
C4312 XA.XIR[13].XIC[14].icell.PDM VGND 0.18803f
C4313 XA.XIR[13].XIC[13].icell.PDM VGND 0.18803f
C4314 XA.XIR[13].XIC[12].icell.PDM VGND 0.18803f
C4315 XA.XIR[13].XIC[11].icell.PDM VGND 0.18803f
C4316 XA.XIR[13].XIC[10].icell.PDM VGND 0.18803f
C4317 XA.XIR[13].XIC[9].icell.PDM VGND 0.18803f
C4318 XA.XIR[13].XIC[8].icell.PDM VGND 0.18803f
C4319 XA.XIR[13].XIC[7].icell.PDM VGND 0.18803f
C4320 XA.XIR[13].XIC[6].icell.PDM VGND 0.18803f
C4321 XA.XIR[13].XIC[5].icell.PDM VGND 0.18803f
C4322 XA.XIR[13].XIC[4].icell.PDM VGND 0.18803f
C4323 XA.XIR[13].XIC[3].icell.PDM VGND 0.18803f
C4324 XA.XIR[13].XIC[2].icell.PDM VGND 0.18803f
C4325 XA.XIR[13].XIC[1].icell.PDM VGND 0.18803f
C4326 XA.XIR[13].XIC[0].icell.PDM VGND 0.1881f
C4327 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C4328 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C4329 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C4330 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60749f
C4331 XA.XIR[12].XIC_15.icell.Ien VGND 0.37186f
C4332 XA.XIR[12].XIC[14].icell.Ien VGND 0.37133f
C4333 XA.XIR[12].XIC[13].icell.Ien VGND 0.37133f
C4334 XA.XIR[12].XIC[12].icell.Ien VGND 0.37133f
C4335 XA.XIR[12].XIC[11].icell.Ien VGND 0.37133f
C4336 XA.XIR[12].XIC[10].icell.Ien VGND 0.37133f
C4337 XA.XIR[12].XIC[9].icell.Ien VGND 0.37133f
C4338 XA.XIR[12].XIC[8].icell.Ien VGND 0.37133f
C4339 XA.XIR[12].XIC[7].icell.Ien VGND 0.37133f
C4340 XA.XIR[12].XIC[6].icell.Ien VGND 0.37133f
C4341 XA.XIR[12].XIC[5].icell.Ien VGND 0.37133f
C4342 XA.XIR[12].XIC[4].icell.Ien VGND 0.37133f
C4343 XA.XIR[12].XIC[3].icell.Ien VGND 0.37133f
C4344 XA.XIR[12].XIC[2].icell.Ien VGND 0.37133f
C4345 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80341f
C4346 XThR.Tn[12] VGND 13.34864f
C4347 XA.XIR[12].XIC[1].icell.Ien VGND 0.37133f
C4348 XA.XIR[12].XIC[0].icell.Ien VGND 0.37135f
C4349 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01013f
C4350 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.5728f
C4351 a_n997_2667# VGND 0.5457f
C4352 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C4353 XA.XIR[12].XIC_15.icell.PDM VGND 0.18849f
C4354 XA.XIR[12].XIC[14].icell.PDM VGND 0.18803f
C4355 XA.XIR[12].XIC[13].icell.PDM VGND 0.18803f
C4356 XA.XIR[12].XIC[12].icell.PDM VGND 0.18803f
C4357 XA.XIR[12].XIC[11].icell.PDM VGND 0.18803f
C4358 XA.XIR[12].XIC[10].icell.PDM VGND 0.18803f
C4359 XA.XIR[12].XIC[9].icell.PDM VGND 0.18803f
C4360 XA.XIR[12].XIC[8].icell.PDM VGND 0.18803f
C4361 XA.XIR[12].XIC[7].icell.PDM VGND 0.18803f
C4362 XA.XIR[12].XIC[6].icell.PDM VGND 0.18803f
C4363 XA.XIR[12].XIC[5].icell.PDM VGND 0.18803f
C4364 XA.XIR[12].XIC[4].icell.PDM VGND 0.18803f
C4365 XA.XIR[12].XIC[3].icell.PDM VGND 0.18803f
C4366 XA.XIR[12].XIC[2].icell.PDM VGND 0.18803f
C4367 XA.XIR[12].XIC[1].icell.PDM VGND 0.18803f
C4368 XA.XIR[12].XIC[0].icell.PDM VGND 0.1881f
C4369 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C4370 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C4371 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C4372 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60749f
C4373 XA.XIR[11].XIC_15.icell.Ien VGND 0.37186f
C4374 XA.XIR[11].XIC[14].icell.Ien VGND 0.37133f
C4375 XA.XIR[11].XIC[13].icell.Ien VGND 0.37133f
C4376 XA.XIR[11].XIC[12].icell.Ien VGND 0.37133f
C4377 XA.XIR[11].XIC[11].icell.Ien VGND 0.37133f
C4378 XA.XIR[11].XIC[10].icell.Ien VGND 0.37133f
C4379 XA.XIR[11].XIC[9].icell.Ien VGND 0.37133f
C4380 XA.XIR[11].XIC[8].icell.Ien VGND 0.37133f
C4381 XA.XIR[11].XIC[7].icell.Ien VGND 0.37133f
C4382 XA.XIR[11].XIC[6].icell.Ien VGND 0.37133f
C4383 XA.XIR[11].XIC[5].icell.Ien VGND 0.37133f
C4384 XA.XIR[11].XIC[4].icell.Ien VGND 0.37133f
C4385 XA.XIR[11].XIC[3].icell.Ien VGND 0.37133f
C4386 XA.XIR[11].XIC[2].icell.Ien VGND 0.37133f
C4387 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.80576f
C4388 XThR.Tn[11] VGND 13.40885f
C4389 XA.XIR[11].XIC[1].icell.Ien VGND 0.37133f
C4390 a_n997_2891# VGND 0.54795f
C4391 XA.XIR[11].XIC[0].icell.Ien VGND 0.37135f
C4392 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01013f
C4393 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57294f
C4394 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C4395 XA.XIR[11].XIC_15.icell.PDM VGND 0.18849f
C4396 XA.XIR[11].XIC[14].icell.PDM VGND 0.18803f
C4397 XA.XIR[11].XIC[13].icell.PDM VGND 0.18803f
C4398 XA.XIR[11].XIC[12].icell.PDM VGND 0.18803f
C4399 XA.XIR[11].XIC[11].icell.PDM VGND 0.18803f
C4400 XA.XIR[11].XIC[10].icell.PDM VGND 0.18803f
C4401 XA.XIR[11].XIC[9].icell.PDM VGND 0.18803f
C4402 XA.XIR[11].XIC[8].icell.PDM VGND 0.18803f
C4403 XA.XIR[11].XIC[7].icell.PDM VGND 0.18803f
C4404 XA.XIR[11].XIC[6].icell.PDM VGND 0.18803f
C4405 XA.XIR[11].XIC[5].icell.PDM VGND 0.18803f
C4406 XA.XIR[11].XIC[4].icell.PDM VGND 0.18803f
C4407 XA.XIR[11].XIC[3].icell.PDM VGND 0.18803f
C4408 XA.XIR[11].XIC[2].icell.PDM VGND 0.18803f
C4409 XA.XIR[11].XIC[1].icell.PDM VGND 0.18803f
C4410 XA.XIR[11].XIC[0].icell.PDM VGND 0.1881f
C4411 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C4412 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C4413 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C4414 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60749f
C4415 XA.XIR[10].XIC_15.icell.Ien VGND 0.37186f
C4416 XA.XIR[10].XIC[14].icell.Ien VGND 0.37133f
C4417 XA.XIR[10].XIC[13].icell.Ien VGND 0.37133f
C4418 XA.XIR[10].XIC[12].icell.Ien VGND 0.37133f
C4419 XA.XIR[10].XIC[11].icell.Ien VGND 0.37133f
C4420 XA.XIR[10].XIC[10].icell.Ien VGND 0.37133f
C4421 XA.XIR[10].XIC[9].icell.Ien VGND 0.37133f
C4422 XA.XIR[10].XIC[8].icell.Ien VGND 0.37133f
C4423 XA.XIR[10].XIC[7].icell.Ien VGND 0.37133f
C4424 XA.XIR[10].XIC[6].icell.Ien VGND 0.37133f
C4425 XA.XIR[10].XIC[5].icell.Ien VGND 0.37133f
C4426 XA.XIR[10].XIC[4].icell.Ien VGND 0.37133f
C4427 XA.XIR[10].XIC[3].icell.Ien VGND 0.37133f
C4428 XA.XIR[10].XIC[2].icell.Ien VGND 0.37133f
C4429 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80459f
C4430 XThR.Tn[10] VGND 13.3903f
C4431 XA.XIR[10].XIC[1].icell.Ien VGND 0.37133f
C4432 XA.XIR[10].XIC[0].icell.Ien VGND 0.37135f
C4433 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01013f
C4434 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57422f
C4435 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C4436 XA.XIR[10].XIC_15.icell.PDM VGND 0.18849f
C4437 XA.XIR[10].XIC[14].icell.PDM VGND 0.18803f
C4438 XA.XIR[10].XIC[13].icell.PDM VGND 0.18803f
C4439 XA.XIR[10].XIC[12].icell.PDM VGND 0.18803f
C4440 XA.XIR[10].XIC[11].icell.PDM VGND 0.18803f
C4441 XA.XIR[10].XIC[10].icell.PDM VGND 0.18803f
C4442 XA.XIR[10].XIC[9].icell.PDM VGND 0.18803f
C4443 XA.XIR[10].XIC[8].icell.PDM VGND 0.18803f
C4444 XA.XIR[10].XIC[7].icell.PDM VGND 0.18803f
C4445 XA.XIR[10].XIC[6].icell.PDM VGND 0.18803f
C4446 XA.XIR[10].XIC[5].icell.PDM VGND 0.18803f
C4447 XA.XIR[10].XIC[4].icell.PDM VGND 0.18803f
C4448 XA.XIR[10].XIC[3].icell.PDM VGND 0.18803f
C4449 XA.XIR[10].XIC[2].icell.PDM VGND 0.18803f
C4450 XA.XIR[10].XIC[1].icell.PDM VGND 0.18803f
C4451 XA.XIR[10].XIC[0].icell.PDM VGND 0.1881f
C4452 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C4453 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C4454 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C4455 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60749f
C4456 XA.XIR[9].XIC_15.icell.Ien VGND 0.37186f
C4457 XA.XIR[9].XIC[14].icell.Ien VGND 0.37133f
C4458 XA.XIR[9].XIC[13].icell.Ien VGND 0.37133f
C4459 XA.XIR[9].XIC[12].icell.Ien VGND 0.37133f
C4460 XA.XIR[9].XIC[11].icell.Ien VGND 0.37133f
C4461 XA.XIR[9].XIC[10].icell.Ien VGND 0.37133f
C4462 XA.XIR[9].XIC[9].icell.Ien VGND 0.37133f
C4463 XA.XIR[9].XIC[8].icell.Ien VGND 0.37133f
C4464 XA.XIR[9].XIC[7].icell.Ien VGND 0.37133f
C4465 XA.XIR[9].XIC[6].icell.Ien VGND 0.37133f
C4466 XA.XIR[9].XIC[5].icell.Ien VGND 0.37133f
C4467 XA.XIR[9].XIC[4].icell.Ien VGND 0.37133f
C4468 XA.XIR[9].XIC[3].icell.Ien VGND 0.37133f
C4469 XA.XIR[9].XIC[2].icell.Ien VGND 0.37133f
C4470 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.80646f
C4471 XA.XIR[9].XIC[1].icell.Ien VGND 0.37133f
C4472 XThR.Tn[9] VGND 13.39284f
C4473 a_n997_3755# VGND 0.54861f
C4474 XA.XIR[9].XIC[0].icell.Ien VGND 0.37135f
C4475 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01013f
C4476 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.5732f
C4477 a_n997_3979# VGND 0.54721f
C4478 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C4479 XA.XIR[9].XIC_15.icell.PDM VGND 0.18849f
C4480 XA.XIR[9].XIC[14].icell.PDM VGND 0.18803f
C4481 XA.XIR[9].XIC[13].icell.PDM VGND 0.18803f
C4482 XA.XIR[9].XIC[12].icell.PDM VGND 0.18803f
C4483 XA.XIR[9].XIC[11].icell.PDM VGND 0.18803f
C4484 XA.XIR[9].XIC[10].icell.PDM VGND 0.18803f
C4485 XA.XIR[9].XIC[9].icell.PDM VGND 0.18803f
C4486 XA.XIR[9].XIC[8].icell.PDM VGND 0.18803f
C4487 XA.XIR[9].XIC[7].icell.PDM VGND 0.18803f
C4488 XA.XIR[9].XIC[6].icell.PDM VGND 0.18803f
C4489 XA.XIR[9].XIC[5].icell.PDM VGND 0.18803f
C4490 XA.XIR[9].XIC[4].icell.PDM VGND 0.18803f
C4491 XA.XIR[9].XIC[3].icell.PDM VGND 0.18803f
C4492 XA.XIR[9].XIC[2].icell.PDM VGND 0.18803f
C4493 XA.XIR[9].XIC[1].icell.PDM VGND 0.18803f
C4494 XA.XIR[9].XIC[0].icell.PDM VGND 0.1881f
C4495 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C4496 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C4497 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C4498 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60749f
C4499 XA.XIR[8].XIC_15.icell.Ien VGND 0.37186f
C4500 XA.XIR[8].XIC[14].icell.Ien VGND 0.37133f
C4501 XA.XIR[8].XIC[13].icell.Ien VGND 0.37133f
C4502 XA.XIR[8].XIC[12].icell.Ien VGND 0.37133f
C4503 XA.XIR[8].XIC[11].icell.Ien VGND 0.37133f
C4504 XA.XIR[8].XIC[10].icell.Ien VGND 0.37133f
C4505 XA.XIR[8].XIC[9].icell.Ien VGND 0.37133f
C4506 XA.XIR[8].XIC[8].icell.Ien VGND 0.37133f
C4507 XA.XIR[8].XIC[7].icell.Ien VGND 0.37133f
C4508 XA.XIR[8].XIC[6].icell.Ien VGND 0.37133f
C4509 XA.XIR[8].XIC[5].icell.Ien VGND 0.37133f
C4510 XA.XIR[8].XIC[4].icell.Ien VGND 0.37133f
C4511 XA.XIR[8].XIC[3].icell.Ien VGND 0.37133f
C4512 XA.XIR[8].XIC[2].icell.Ien VGND 0.37133f
C4513 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80378f
C4514 XA.XIR[8].XIC[1].icell.Ien VGND 0.37133f
C4515 XThR.Tn[8] VGND 13.37547f
C4516 XA.XIR[8].XIC[0].icell.Ien VGND 0.37135f
C4517 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01013f
C4518 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57308f
C4519 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C4520 XA.XIR[8].XIC_15.icell.PDM VGND 0.18849f
C4521 XA.XIR[8].XIC[14].icell.PDM VGND 0.18803f
C4522 XA.XIR[8].XIC[13].icell.PDM VGND 0.18803f
C4523 XA.XIR[8].XIC[12].icell.PDM VGND 0.18803f
C4524 XA.XIR[8].XIC[11].icell.PDM VGND 0.18803f
C4525 XA.XIR[8].XIC[10].icell.PDM VGND 0.18803f
C4526 XA.XIR[8].XIC[9].icell.PDM VGND 0.18803f
C4527 XA.XIR[8].XIC[8].icell.PDM VGND 0.18803f
C4528 XA.XIR[8].XIC[7].icell.PDM VGND 0.18803f
C4529 XA.XIR[8].XIC[6].icell.PDM VGND 0.18803f
C4530 XA.XIR[8].XIC[5].icell.PDM VGND 0.18803f
C4531 XA.XIR[8].XIC[4].icell.PDM VGND 0.18803f
C4532 XA.XIR[8].XIC[3].icell.PDM VGND 0.18803f
C4533 XA.XIR[8].XIC[2].icell.PDM VGND 0.18803f
C4534 XA.XIR[8].XIC[1].icell.PDM VGND 0.18803f
C4535 XA.XIR[8].XIC[0].icell.PDM VGND 0.1881f
C4536 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C4537 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C4538 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C4539 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60749f
C4540 XA.XIR[7].XIC_15.icell.Ien VGND 0.37186f
C4541 XA.XIR[7].XIC[14].icell.Ien VGND 0.37133f
C4542 XA.XIR[7].XIC[13].icell.Ien VGND 0.37133f
C4543 XA.XIR[7].XIC[12].icell.Ien VGND 0.37133f
C4544 XA.XIR[7].XIC[11].icell.Ien VGND 0.37133f
C4545 XA.XIR[7].XIC[10].icell.Ien VGND 0.37133f
C4546 XA.XIR[7].XIC[9].icell.Ien VGND 0.37133f
C4547 XA.XIR[7].XIC[8].icell.Ien VGND 0.37133f
C4548 XA.XIR[7].XIC[7].icell.Ien VGND 0.37133f
C4549 XA.XIR[7].XIC[6].icell.Ien VGND 0.37133f
C4550 XA.XIR[7].XIC[5].icell.Ien VGND 0.37133f
C4551 XA.XIR[7].XIC[4].icell.Ien VGND 0.37133f
C4552 XA.XIR[7].XIC[3].icell.Ien VGND 0.37133f
C4553 XA.XIR[7].XIC[2].icell.Ien VGND 0.37133f
C4554 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80409f
C4555 XA.XIR[7].XIC[1].icell.Ien VGND 0.37133f
C4556 XA.XIR[7].XIC[0].icell.Ien VGND 0.37135f
C4557 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01013f
C4558 XThR.Tn[7] VGND 13.8085f
C4559 XThR.XTBN.A VGND 1.22812f
C4560 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57516f
C4561 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C4562 XA.XIR[7].XIC_15.icell.PDM VGND 0.18849f
C4563 XA.XIR[7].XIC[14].icell.PDM VGND 0.18803f
C4564 XA.XIR[7].XIC[13].icell.PDM VGND 0.18803f
C4565 XA.XIR[7].XIC[12].icell.PDM VGND 0.18803f
C4566 XA.XIR[7].XIC[11].icell.PDM VGND 0.18803f
C4567 XA.XIR[7].XIC[10].icell.PDM VGND 0.18803f
C4568 XA.XIR[7].XIC[9].icell.PDM VGND 0.18803f
C4569 XA.XIR[7].XIC[8].icell.PDM VGND 0.18803f
C4570 XA.XIR[7].XIC[7].icell.PDM VGND 0.18803f
C4571 XA.XIR[7].XIC[6].icell.PDM VGND 0.18803f
C4572 XA.XIR[7].XIC[5].icell.PDM VGND 0.18803f
C4573 XA.XIR[7].XIC[4].icell.PDM VGND 0.18803f
C4574 XA.XIR[7].XIC[3].icell.PDM VGND 0.18803f
C4575 XA.XIR[7].XIC[2].icell.PDM VGND 0.18803f
C4576 XA.XIR[7].XIC[1].icell.PDM VGND 0.18803f
C4577 XA.XIR[7].XIC[0].icell.PDM VGND 0.1881f
C4578 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C4579 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C4580 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C4581 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60749f
C4582 XA.XIR[6].XIC_15.icell.Ien VGND 0.37186f
C4583 XA.XIR[6].XIC[14].icell.Ien VGND 0.37133f
C4584 XA.XIR[6].XIC[13].icell.Ien VGND 0.37133f
C4585 XA.XIR[6].XIC[12].icell.Ien VGND 0.37133f
C4586 XA.XIR[6].XIC[11].icell.Ien VGND 0.37133f
C4587 XA.XIR[6].XIC[10].icell.Ien VGND 0.37133f
C4588 XA.XIR[6].XIC[9].icell.Ien VGND 0.37133f
C4589 XA.XIR[6].XIC[8].icell.Ien VGND 0.37133f
C4590 XA.XIR[6].XIC[7].icell.Ien VGND 0.37133f
C4591 XA.XIR[6].XIC[6].icell.Ien VGND 0.37133f
C4592 XA.XIR[6].XIC[5].icell.Ien VGND 0.37133f
C4593 XA.XIR[6].XIC[4].icell.Ien VGND 0.37133f
C4594 XA.XIR[6].XIC[3].icell.Ien VGND 0.37133f
C4595 XA.XIR[6].XIC[2].icell.Ien VGND 0.37133f
C4596 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80504f
C4597 XA.XIR[6].XIC[1].icell.Ien VGND 0.37133f
C4598 XA.XIR[6].XIC[0].icell.Ien VGND 0.37135f
C4599 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01013f
C4600 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57422f
C4601 XThR.Tn[6] VGND 13.43458f
C4602 a_n1049_5317# VGND 0.02283f
C4603 XThR.XTB7.Y VGND 1.36131f
C4604 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C4605 XA.XIR[6].XIC_15.icell.PDM VGND 0.18849f
C4606 XA.XIR[6].XIC[14].icell.PDM VGND 0.18803f
C4607 XA.XIR[6].XIC[13].icell.PDM VGND 0.18803f
C4608 XA.XIR[6].XIC[12].icell.PDM VGND 0.18803f
C4609 XA.XIR[6].XIC[11].icell.PDM VGND 0.18803f
C4610 XA.XIR[6].XIC[10].icell.PDM VGND 0.18803f
C4611 XA.XIR[6].XIC[9].icell.PDM VGND 0.18803f
C4612 XA.XIR[6].XIC[8].icell.PDM VGND 0.18803f
C4613 XA.XIR[6].XIC[7].icell.PDM VGND 0.18803f
C4614 XA.XIR[6].XIC[6].icell.PDM VGND 0.18803f
C4615 XA.XIR[6].XIC[5].icell.PDM VGND 0.18803f
C4616 XA.XIR[6].XIC[4].icell.PDM VGND 0.18803f
C4617 XA.XIR[6].XIC[3].icell.PDM VGND 0.18803f
C4618 XA.XIR[6].XIC[2].icell.PDM VGND 0.18803f
C4619 XA.XIR[6].XIC[1].icell.PDM VGND 0.18803f
C4620 XA.XIR[6].XIC[0].icell.PDM VGND 0.1881f
C4621 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C4622 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C4623 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C4624 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60749f
C4625 XA.XIR[5].XIC_15.icell.Ien VGND 0.37186f
C4626 XA.XIR[5].XIC[14].icell.Ien VGND 0.37133f
C4627 XA.XIR[5].XIC[13].icell.Ien VGND 0.37133f
C4628 XA.XIR[5].XIC[12].icell.Ien VGND 0.37133f
C4629 XA.XIR[5].XIC[11].icell.Ien VGND 0.37133f
C4630 XA.XIR[5].XIC[10].icell.Ien VGND 0.37133f
C4631 XA.XIR[5].XIC[9].icell.Ien VGND 0.37133f
C4632 XA.XIR[5].XIC[8].icell.Ien VGND 0.37133f
C4633 XA.XIR[5].XIC[7].icell.Ien VGND 0.37133f
C4634 XA.XIR[5].XIC[6].icell.Ien VGND 0.37133f
C4635 XA.XIR[5].XIC[5].icell.Ien VGND 0.37133f
C4636 XA.XIR[5].XIC[4].icell.Ien VGND 0.37133f
C4637 XA.XIR[5].XIC[3].icell.Ien VGND 0.37133f
C4638 XA.XIR[5].XIC[2].icell.Ien VGND 0.37133f
C4639 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80373f
C4640 XA.XIR[5].XIC[1].icell.Ien VGND 0.37133f
C4641 a_n1049_5611# VGND 0.02888f
C4642 XA.XIR[5].XIC[0].icell.Ien VGND 0.37135f
C4643 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01013f
C4644 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57288f
C4645 XThR.Tn[5] VGND 13.45136f
C4646 XThR.XTB6.Y VGND 1.38207f
C4647 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C4648 XA.XIR[5].XIC_15.icell.PDM VGND 0.18849f
C4649 XA.XIR[5].XIC[14].icell.PDM VGND 0.18803f
C4650 XA.XIR[5].XIC[13].icell.PDM VGND 0.18803f
C4651 XA.XIR[5].XIC[12].icell.PDM VGND 0.18803f
C4652 XA.XIR[5].XIC[11].icell.PDM VGND 0.18803f
C4653 XA.XIR[5].XIC[10].icell.PDM VGND 0.18803f
C4654 XA.XIR[5].XIC[9].icell.PDM VGND 0.18803f
C4655 XA.XIR[5].XIC[8].icell.PDM VGND 0.18803f
C4656 XA.XIR[5].XIC[7].icell.PDM VGND 0.18803f
C4657 XA.XIR[5].XIC[6].icell.PDM VGND 0.18803f
C4658 XA.XIR[5].XIC[5].icell.PDM VGND 0.18803f
C4659 XA.XIR[5].XIC[4].icell.PDM VGND 0.18803f
C4660 XA.XIR[5].XIC[3].icell.PDM VGND 0.18803f
C4661 XA.XIR[5].XIC[2].icell.PDM VGND 0.18803f
C4662 XA.XIR[5].XIC[1].icell.PDM VGND 0.18803f
C4663 XA.XIR[5].XIC[0].icell.PDM VGND 0.1881f
C4664 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C4665 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C4666 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C4667 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60749f
C4668 XA.XIR[4].XIC_15.icell.Ien VGND 0.37186f
C4669 XA.XIR[4].XIC[14].icell.Ien VGND 0.37133f
C4670 XA.XIR[4].XIC[13].icell.Ien VGND 0.37133f
C4671 XA.XIR[4].XIC[12].icell.Ien VGND 0.37133f
C4672 XA.XIR[4].XIC[11].icell.Ien VGND 0.37133f
C4673 XA.XIR[4].XIC[10].icell.Ien VGND 0.37133f
C4674 XA.XIR[4].XIC[9].icell.Ien VGND 0.37133f
C4675 XA.XIR[4].XIC[8].icell.Ien VGND 0.37133f
C4676 XA.XIR[4].XIC[7].icell.Ien VGND 0.37133f
C4677 XA.XIR[4].XIC[6].icell.Ien VGND 0.37133f
C4678 XA.XIR[4].XIC[5].icell.Ien VGND 0.37133f
C4679 XA.XIR[4].XIC[4].icell.Ien VGND 0.37133f
C4680 XA.XIR[4].XIC[3].icell.Ien VGND 0.37133f
C4681 XA.XIR[4].XIC[2].icell.Ien VGND 0.37133f
C4682 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.80546f
C4683 XA.XIR[4].XIC[1].icell.Ien VGND 0.37133f
C4684 XA.XIR[4].XIC[0].icell.Ien VGND 0.37135f
C4685 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01013f
C4686 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57333f
C4687 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C4688 XA.XIR[4].XIC_15.icell.PDM VGND 0.18849f
C4689 XA.XIR[4].XIC[14].icell.PDM VGND 0.18803f
C4690 XA.XIR[4].XIC[13].icell.PDM VGND 0.18803f
C4691 XA.XIR[4].XIC[12].icell.PDM VGND 0.18803f
C4692 XA.XIR[4].XIC[11].icell.PDM VGND 0.18803f
C4693 XA.XIR[4].XIC[10].icell.PDM VGND 0.18803f
C4694 XA.XIR[4].XIC[9].icell.PDM VGND 0.18803f
C4695 XA.XIR[4].XIC[8].icell.PDM VGND 0.18803f
C4696 XA.XIR[4].XIC[7].icell.PDM VGND 0.18803f
C4697 XA.XIR[4].XIC[6].icell.PDM VGND 0.18803f
C4698 XA.XIR[4].XIC[5].icell.PDM VGND 0.18803f
C4699 XA.XIR[4].XIC[4].icell.PDM VGND 0.18803f
C4700 XA.XIR[4].XIC[3].icell.PDM VGND 0.18803f
C4701 XA.XIR[4].XIC[2].icell.PDM VGND 0.18803f
C4702 XA.XIR[4].XIC[1].icell.PDM VGND 0.18803f
C4703 XA.XIR[4].XIC[0].icell.PDM VGND 0.1881f
C4704 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C4705 XThR.Tn[4] VGND 13.51876f
C4706 a_n1049_6405# VGND 0.02935f
C4707 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C4708 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C4709 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60749f
C4710 XA.XIR[3].XIC_15.icell.Ien VGND 0.37186f
C4711 XA.XIR[3].XIC[14].icell.Ien VGND 0.37133f
C4712 XA.XIR[3].XIC[13].icell.Ien VGND 0.37133f
C4713 XA.XIR[3].XIC[12].icell.Ien VGND 0.37133f
C4714 XA.XIR[3].XIC[11].icell.Ien VGND 0.37133f
C4715 XA.XIR[3].XIC[10].icell.Ien VGND 0.37133f
C4716 XA.XIR[3].XIC[9].icell.Ien VGND 0.37133f
C4717 XA.XIR[3].XIC[8].icell.Ien VGND 0.37133f
C4718 XA.XIR[3].XIC[7].icell.Ien VGND 0.37133f
C4719 XA.XIR[3].XIC[6].icell.Ien VGND 0.37133f
C4720 XA.XIR[3].XIC[5].icell.Ien VGND 0.37133f
C4721 XA.XIR[3].XIC[4].icell.Ien VGND 0.37133f
C4722 XA.XIR[3].XIC[3].icell.Ien VGND 0.37133f
C4723 XA.XIR[3].XIC[2].icell.Ien VGND 0.37133f
C4724 XThR.XTB5.Y VGND 1.32752f
C4725 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80386f
C4726 XA.XIR[3].XIC[1].icell.Ien VGND 0.37133f
C4727 XA.XIR[3].XIC[0].icell.Ien VGND 0.37135f
C4728 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01013f
C4729 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57422f
C4730 a_n1049_6699# VGND 0.02979f
C4731 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C4732 XA.XIR[3].XIC_15.icell.PDM VGND 0.18849f
C4733 XA.XIR[3].XIC[14].icell.PDM VGND 0.18803f
C4734 XA.XIR[3].XIC[13].icell.PDM VGND 0.18803f
C4735 XA.XIR[3].XIC[12].icell.PDM VGND 0.18803f
C4736 XA.XIR[3].XIC[11].icell.PDM VGND 0.18803f
C4737 XA.XIR[3].XIC[10].icell.PDM VGND 0.18803f
C4738 XA.XIR[3].XIC[9].icell.PDM VGND 0.18803f
C4739 XA.XIR[3].XIC[8].icell.PDM VGND 0.18803f
C4740 XA.XIR[3].XIC[7].icell.PDM VGND 0.18803f
C4741 XA.XIR[3].XIC[6].icell.PDM VGND 0.18803f
C4742 XA.XIR[3].XIC[5].icell.PDM VGND 0.18803f
C4743 XA.XIR[3].XIC[4].icell.PDM VGND 0.18803f
C4744 XA.XIR[3].XIC[3].icell.PDM VGND 0.18803f
C4745 XA.XIR[3].XIC[2].icell.PDM VGND 0.18803f
C4746 XA.XIR[3].XIC[1].icell.PDM VGND 0.18803f
C4747 XA.XIR[3].XIC[0].icell.PDM VGND 0.1881f
C4748 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C4749 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C4750 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C4751 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60749f
C4752 XA.XIR[2].XIC_15.icell.Ien VGND 0.37186f
C4753 XA.XIR[2].XIC[14].icell.Ien VGND 0.3714f
C4754 XA.XIR[2].XIC[13].icell.Ien VGND 0.3714f
C4755 XA.XIR[2].XIC[12].icell.Ien VGND 0.3714f
C4756 XA.XIR[2].XIC[11].icell.Ien VGND 0.3714f
C4757 XA.XIR[2].XIC[10].icell.Ien VGND 0.3714f
C4758 XA.XIR[2].XIC[9].icell.Ien VGND 0.3714f
C4759 XA.XIR[2].XIC[8].icell.Ien VGND 0.3714f
C4760 XA.XIR[2].XIC[7].icell.Ien VGND 0.3714f
C4761 XA.XIR[2].XIC[6].icell.Ien VGND 0.3714f
C4762 XA.XIR[2].XIC[5].icell.Ien VGND 0.3714f
C4763 XA.XIR[2].XIC[4].icell.Ien VGND 0.3714f
C4764 XA.XIR[2].XIC[3].icell.Ien VGND 0.3714f
C4765 XA.XIR[2].XIC[2].icell.Ien VGND 0.3714f
C4766 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80601f
C4767 XA.XIR[2].XIC[1].icell.Ien VGND 0.3714f
C4768 XThR.Tn[3] VGND 13.46766f
C4769 XThR.XTB4.Y VGND 1.48813f
C4770 XA.XIR[2].XIC[0].icell.Ien VGND 0.37142f
C4771 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01013f
C4772 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57552f
C4773 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C4774 XA.XIR[2].XIC_15.icell.PDM VGND 0.18849f
C4775 XA.XIR[2].XIC[14].icell.PDM VGND 0.1883f
C4776 XA.XIR[2].XIC[13].icell.PDM VGND 0.1883f
C4777 XA.XIR[2].XIC[12].icell.PDM VGND 0.1883f
C4778 XA.XIR[2].XIC[11].icell.PDM VGND 0.1883f
C4779 XA.XIR[2].XIC[10].icell.PDM VGND 0.1883f
C4780 XA.XIR[2].XIC[9].icell.PDM VGND 0.1883f
C4781 XA.XIR[2].XIC[8].icell.PDM VGND 0.1883f
C4782 XA.XIR[2].XIC[7].icell.PDM VGND 0.1883f
C4783 XA.XIR[2].XIC[6].icell.PDM VGND 0.1883f
C4784 XA.XIR[2].XIC[5].icell.PDM VGND 0.1883f
C4785 XA.XIR[2].XIC[4].icell.PDM VGND 0.1883f
C4786 XA.XIR[2].XIC[3].icell.PDM VGND 0.1883f
C4787 XA.XIR[2].XIC[2].icell.PDM VGND 0.1883f
C4788 XA.XIR[2].XIC[1].icell.PDM VGND 0.1883f
C4789 XA.XIR[2].XIC[0].icell.PDM VGND 0.18837f
C4790 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C4791 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C4792 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C4793 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60749f
C4794 XA.XIR[1].XIC_15.icell.Ien VGND 0.37186f
C4795 XA.XIR[1].XIC[14].icell.Ien VGND 0.37167f
C4796 XA.XIR[1].XIC[13].icell.Ien VGND 0.37167f
C4797 XA.XIR[1].XIC[12].icell.Ien VGND 0.37167f
C4798 XA.XIR[1].XIC[11].icell.Ien VGND 0.37167f
C4799 XA.XIR[1].XIC[10].icell.Ien VGND 0.37167f
C4800 XA.XIR[1].XIC[9].icell.Ien VGND 0.37167f
C4801 XA.XIR[1].XIC[8].icell.Ien VGND 0.37167f
C4802 XA.XIR[1].XIC[7].icell.Ien VGND 0.37167f
C4803 XA.XIR[1].XIC[6].icell.Ien VGND 0.37167f
C4804 XA.XIR[1].XIC[5].icell.Ien VGND 0.37167f
C4805 XA.XIR[1].XIC[4].icell.Ien VGND 0.37167f
C4806 XA.XIR[1].XIC[3].icell.Ien VGND 0.37167f
C4807 XA.XIR[1].XIC[2].icell.Ien VGND 0.37167f
C4808 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80386f
C4809 XA.XIR[1].XIC[1].icell.Ien VGND 0.37167f
C4810 XThR.Tn[2] VGND 13.52038f
C4811 a_n1049_7493# VGND 0.02484f
C4812 XThR.XTB3.Y VGND 1.24034f
C4813 XThR.XTB7.A VGND 1.95524f
C4814 XA.XIR[1].XIC[0].icell.Ien VGND 0.37169f
C4815 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01013f
C4816 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57375f
C4817 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C4818 XA.XIR[1].XIC_15.icell.PDM VGND 0.18849f
C4819 XA.XIR[1].XIC[14].icell.PDM VGND 0.18855f
C4820 XA.XIR[1].XIC[13].icell.PDM VGND 0.18855f
C4821 XA.XIR[1].XIC[12].icell.PDM VGND 0.18855f
C4822 XA.XIR[1].XIC[11].icell.PDM VGND 0.18855f
C4823 XA.XIR[1].XIC[10].icell.PDM VGND 0.18855f
C4824 XA.XIR[1].XIC[9].icell.PDM VGND 0.18855f
C4825 XA.XIR[1].XIC[8].icell.PDM VGND 0.18855f
C4826 XA.XIR[1].XIC[7].icell.PDM VGND 0.18855f
C4827 XA.XIR[1].XIC[6].icell.PDM VGND 0.18855f
C4828 XA.XIR[1].XIC[5].icell.PDM VGND 0.18855f
C4829 XA.XIR[1].XIC[4].icell.PDM VGND 0.18855f
C4830 XA.XIR[1].XIC[3].icell.PDM VGND 0.18855f
C4831 XA.XIR[1].XIC[2].icell.PDM VGND 0.18855f
C4832 XA.XIR[1].XIC[1].icell.PDM VGND 0.18855f
C4833 XA.XIR[1].XIC[0].icell.PDM VGND 0.18862f
C4834 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C4835 a_n1049_7787# VGND 0.03396f
C4836 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87401f
C4837 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C4838 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61803f
C4839 XA.XIR[0].XIC_15.icell.Ien VGND 0.3793f
C4840 XA.XIR[0].XIC[14].icell.Ien VGND 0.3898f
C4841 XA.XIR[0].XIC[13].icell.Ien VGND 0.38977f
C4842 XA.XIR[0].XIC[12].icell.Ien VGND 0.3864f
C4843 XA.XIR[0].XIC[11].icell.Ien VGND 0.38713f
C4844 XA.XIR[0].XIC[10].icell.Ien VGND 0.38848f
C4845 XA.XIR[0].XIC[9].icell.Ien VGND 0.38677f
C4846 XA.XIR[0].XIC[8].icell.Ien VGND 0.38726f
C4847 XA.XIR[0].XIC[7].icell.Ien VGND 0.38752f
C4848 XA.XIR[0].XIC[6].icell.Ien VGND 0.3875f
C4849 XA.XIR[0].XIC[5].icell.Ien VGND 0.38643f
C4850 XA.XIR[0].XIC[4].icell.Ien VGND 0.38645f
C4851 XA.XIR[0].XIC[3].icell.Ien VGND 0.38768f
C4852 XA.XIR[0].XIC[2].icell.Ien VGND 0.38976f
C4853 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83f
C4854 XA.XIR[0].XIC[1].icell.Ien VGND 0.39004f
C4855 XA.XIR[0].XIC[0].icell.Ien VGND 0.38887f
C4856 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01013f
C4857 XThR.Tn[1] VGND 13.52625f
C4858 XThR.XTB2.Y VGND 1.47429f
C4859 XThR.XTB6.A VGND 0.95405f
C4860 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58593f
C4861 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.25235f
C4862 XA.XIR[0].XIC_15.icell.PDM VGND 0.20832f
C4863 XA.XIR[0].XIC[14].icell.PDM VGND 0.24785f
C4864 XA.XIR[0].XIC[13].icell.PDM VGND 0.24797f
C4865 XA.XIR[0].XIC[12].icell.PDM VGND 0.24357f
C4866 XA.XIR[0].XIC[11].icell.PDM VGND 0.24401f
C4867 XA.XIR[0].XIC[10].icell.PDM VGND 0.24391f
C4868 XA.XIR[0].XIC[9].icell.PDM VGND 0.24364f
C4869 XA.XIR[0].XIC[8].icell.PDM VGND 0.24363f
C4870 XA.XIR[0].XIC[7].icell.PDM VGND 0.24632f
C4871 XA.XIR[0].XIC[6].icell.PDM VGND 0.24369f
C4872 XA.XIR[0].XIC[5].icell.PDM VGND 0.24528f
C4873 XA.XIR[0].XIC[4].icell.PDM VGND 0.24366f
C4874 XA.XIR[0].XIC[3].icell.PDM VGND 0.24652f
C4875 XA.XIR[0].XIC[2].icell.PDM VGND 0.24787f
C4876 XA.XIR[0].XIC[1].icell.PDM VGND 0.24823f
C4877 XA.XIR[0].XIC[0].icell.PDM VGND 0.24704f
C4878 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.25065f
C4879 XThR.Tn[0] VGND 13.85341f
C4880 a_n1049_8581# VGND 0.0432f
C4881 XThR.XTBN.Y VGND 7.75072f
C4882 XThR.XTB1.Y VGND 1.8088f
C4883 XThR.XTB7.B VGND 2.60658f
C4884 XThR.XTB5.A VGND 1.75667f
C4885 XThC.Tn[14] VGND 6.00623f
C4886 XThC.Tn[13] VGND 5.60193f
C4887 XThC.Tn[12] VGND 5.57147f
C4888 XThC.Tn[11] VGND 6.15635f
C4889 XThC.Tn[10] VGND 5.26243f
C4890 XThC.Tn[9] VGND 5.77617f
C4891 XThC.Tn[8] VGND 4.97998f
C4892 a_10915_9569# VGND 0.57433f
C4893 a_10051_9569# VGND 0.56318f
C4894 a_9827_9569# VGND 0.55231f
C4895 a_8963_9569# VGND 0.56097f
C4896 a_8739_9569# VGND 0.55929f
C4897 a_7875_9569# VGND 0.56085f
C4898 a_7651_9569# VGND 0.5637f
C4899 XThC.Tn[7] VGND 5.70917f
C4900 XThC.Tn[6] VGND 5.91047f
C4901 XThC.Tn[5] VGND 6.0719f
C4902 XThC.Tn[4] VGND 6.05697f
C4903 XThC.Tn[3] VGND 6.69514f
C4904 XThC.Tn[2] VGND 6.2357f
C4905 XThC.Tn[1] VGND 6.43885f
C4906 XThC.Tn[0] VGND 7.38918f
C4907 a_6243_9615# VGND 0.03813f
C4908 a_5949_9615# VGND 0.04241f
C4909 a_5155_9615# VGND 0.04331f
C4910 a_4861_9615# VGND 0.04637f
C4911 a_4067_9615# VGND 0.04009f
C4912 a_3773_9615# VGND 0.04579f
C4913 a_2979_9615# VGND 0.05579f
C4914 XThC.XTBN.Y VGND 9.62582f
C4915 XThC.XTB7.Y VGND 1.36148f
C4916 XThC.XTB6.Y VGND 1.38096f
C4917 XThC.XTB7.B VGND 2.86322f
C4918 XThC.XTB5.Y VGND 1.32715f
C4919 XThC.XTBN.A VGND 1.22509f
C4920 XThC.XTB4.Y VGND 1.69459f
C4921 XThC.XTB3.Y VGND 1.96884f
C4922 XThC.XTB7.A VGND 1.95016f
C4923 XThC.XTB6.A VGND 0.95488f
C4924 XThC.XTB2.Y VGND 1.47578f
C4925 XThC.XTB1.Y VGND 1.77909f
C4926 XThC.XTB5.A VGND 1.76008f
C4927 bias[0].t0 VGND 0.86609f
C4928 bias[0].n0 VGND 0.31538f
C4929 bias[0].n1 VGND 0.22269f
C4930 bias[0].t1 VGND 0.86609f
C4931 bias[0].n2 VGND 0.33687f
C4932 XThR.XTB1.Y.t1 VGND 0.03165f
C4933 XThR.XTB1.Y.t8 VGND 0.02512f
C4934 XThR.XTB1.Y.t15 VGND 0.0148f
C4935 XThR.XTB1.Y.t14 VGND 0.02512f
C4936 XThR.XTB1.Y.t7 VGND 0.0148f
C4937 XThR.XTB1.Y.t10 VGND 0.02512f
C4938 XThR.XTB1.Y.t18 VGND 0.0148f
C4939 XThR.XTB1.Y.n1 VGND 0.04215f
C4940 XThR.XTB1.Y.n2 VGND 0.04452f
C4941 XThR.XTB1.Y.n3 VGND 0.01831f
C4942 XThR.XTB1.Y.n4 VGND 0.03623f
C4943 XThR.XTB1.Y.t13 VGND 0.02512f
C4944 XThR.XTB1.Y.t4 VGND 0.0148f
C4945 XThR.XTB1.Y.n5 VGND 0.03386f
C4946 XThR.XTB1.Y.n6 VGND 0.01658f
C4947 XThR.XTB1.Y.n7 VGND 0.01376f
C4948 XThR.XTB1.Y.t6 VGND 0.02512f
C4949 XThR.XTB1.Y.t11 VGND 0.0148f
C4950 XThR.XTB1.Y.n8 VGND 0.0154f
C4951 XThR.XTB1.Y.t12 VGND 0.02512f
C4952 XThR.XTB1.Y.t16 VGND 0.0148f
C4953 XThR.XTB1.Y.n9 VGND 0.0307f
C4954 XThR.XTB1.Y.t17 VGND 0.02512f
C4955 XThR.XTB1.Y.t5 VGND 0.0148f
C4956 XThR.XTB1.Y.n10 VGND 0.03307f
C4957 XThR.XTB1.Y.n11 VGND 0.01868f
C4958 XThR.XTB1.Y.n12 VGND 0.03092f
C4959 XThR.XTB1.Y.n13 VGND 0.01603f
C4960 XThR.XTB1.Y.n14 VGND 0.01461f
C4961 XThR.XTB1.Y.n15 VGND 0.03307f
C4962 XThR.XTB1.Y.t3 VGND 0.02512f
C4963 XThR.XTB1.Y.t9 VGND 0.0148f
C4964 XThR.XTB1.Y.n16 VGND 0.02991f
C4965 XThR.XTB1.Y.n17 VGND 0.01658f
C4966 XThR.XTB1.Y.n18 VGND 0.02412f
C4967 XThR.XTB1.Y.n19 VGND 0.75219f
C4968 XThR.XTB1.Y.t0 VGND 0.01615f
C4969 XThR.XTB1.Y.t2 VGND 0.01615f
C4970 XThR.XTB1.Y.n20 VGND 0.03467f
C4971 XThR.XTB1.Y.n21 VGND 0.08068f
C4972 XThR.XTB1.Y.n22 VGND 0.01689f
C4973 XThR.Tn[13].t2 VGND 0.02271f
C4974 XThR.Tn[13].t0 VGND 0.02271f
C4975 XThR.Tn[13].n0 VGND 0.05049f
C4976 XThR.Tn[13].t1 VGND 0.02271f
C4977 XThR.Tn[13].t3 VGND 0.02271f
C4978 XThR.Tn[13].n1 VGND 0.06896f
C4979 XThR.Tn[13].n2 VGND 0.22956f
C4980 XThR.Tn[13].t11 VGND 0.01476f
C4981 XThR.Tn[13].t9 VGND 0.01476f
C4982 XThR.Tn[13].n3 VGND 0.03682f
C4983 XThR.Tn[13].t10 VGND 0.01476f
C4984 XThR.Tn[13].t8 VGND 0.01476f
C4985 XThR.Tn[13].n4 VGND 0.02953f
C4986 XThR.Tn[13].n5 VGND 0.07427f
C4987 XThR.Tn[13].t72 VGND 0.01775f
C4988 XThR.Tn[13].t64 VGND 0.01944f
C4989 XThR.Tn[13].n6 VGND 0.04746f
C4990 XThR.Tn[13].n7 VGND 0.07376f
C4991 XThR.Tn[13].t28 VGND 0.01775f
C4992 XThR.Tn[13].t21 VGND 0.01944f
C4993 XThR.Tn[13].n8 VGND 0.04746f
C4994 XThR.Tn[13].t44 VGND 0.01769f
C4995 XThR.Tn[13].t12 VGND 0.01937f
C4996 XThR.Tn[13].n9 VGND 0.04938f
C4997 XThR.Tn[13].n10 VGND 0.03469f
C4998 XThR.Tn[13].n12 VGND 0.11133f
C4999 XThR.Tn[13].t65 VGND 0.01775f
C5000 XThR.Tn[13].t57 VGND 0.01944f
C5001 XThR.Tn[13].n13 VGND 0.04746f
C5002 XThR.Tn[13].t19 VGND 0.01769f
C5003 XThR.Tn[13].t52 VGND 0.01937f
C5004 XThR.Tn[13].n14 VGND 0.04938f
C5005 XThR.Tn[13].n15 VGND 0.03469f
C5006 XThR.Tn[13].n17 VGND 0.11133f
C5007 XThR.Tn[13].t22 VGND 0.01775f
C5008 XThR.Tn[13].t14 VGND 0.01944f
C5009 XThR.Tn[13].n18 VGND 0.04746f
C5010 XThR.Tn[13].t34 VGND 0.01769f
C5011 XThR.Tn[13].t70 VGND 0.01937f
C5012 XThR.Tn[13].n19 VGND 0.04938f
C5013 XThR.Tn[13].n20 VGND 0.03469f
C5014 XThR.Tn[13].n22 VGND 0.11133f
C5015 XThR.Tn[13].t49 VGND 0.01775f
C5016 XThR.Tn[13].t39 VGND 0.01944f
C5017 XThR.Tn[13].n23 VGND 0.04746f
C5018 XThR.Tn[13].t66 VGND 0.01769f
C5019 XThR.Tn[13].t35 VGND 0.01937f
C5020 XThR.Tn[13].n24 VGND 0.04938f
C5021 XThR.Tn[13].n25 VGND 0.03469f
C5022 XThR.Tn[13].n27 VGND 0.11133f
C5023 XThR.Tn[13].t24 VGND 0.01775f
C5024 XThR.Tn[13].t16 VGND 0.01944f
C5025 XThR.Tn[13].n28 VGND 0.04746f
C5026 XThR.Tn[13].t37 VGND 0.01769f
C5027 XThR.Tn[13].t71 VGND 0.01937f
C5028 XThR.Tn[13].n29 VGND 0.04938f
C5029 XThR.Tn[13].n30 VGND 0.03469f
C5030 XThR.Tn[13].n32 VGND 0.11133f
C5031 XThR.Tn[13].t60 VGND 0.01775f
C5032 XThR.Tn[13].t30 VGND 0.01944f
C5033 XThR.Tn[13].n33 VGND 0.04746f
C5034 XThR.Tn[13].t13 VGND 0.01769f
C5035 XThR.Tn[13].t26 VGND 0.01937f
C5036 XThR.Tn[13].n34 VGND 0.04938f
C5037 XThR.Tn[13].n35 VGND 0.03469f
C5038 XThR.Tn[13].n37 VGND 0.11133f
C5039 XThR.Tn[13].t29 VGND 0.01775f
C5040 XThR.Tn[13].t25 VGND 0.01944f
C5041 XThR.Tn[13].n38 VGND 0.04746f
C5042 XThR.Tn[13].t43 VGND 0.01769f
C5043 XThR.Tn[13].t18 VGND 0.01937f
C5044 XThR.Tn[13].n39 VGND 0.04938f
C5045 XThR.Tn[13].n40 VGND 0.03469f
C5046 XThR.Tn[13].n42 VGND 0.11133f
C5047 XThR.Tn[13].t32 VGND 0.01775f
C5048 XThR.Tn[13].t38 VGND 0.01944f
C5049 XThR.Tn[13].n43 VGND 0.04746f
C5050 XThR.Tn[13].t48 VGND 0.01769f
C5051 XThR.Tn[13].t33 VGND 0.01937f
C5052 XThR.Tn[13].n44 VGND 0.04938f
C5053 XThR.Tn[13].n45 VGND 0.03469f
C5054 XThR.Tn[13].n47 VGND 0.11133f
C5055 XThR.Tn[13].t51 VGND 0.01775f
C5056 XThR.Tn[13].t59 VGND 0.01944f
C5057 XThR.Tn[13].n48 VGND 0.04746f
C5058 XThR.Tn[13].t68 VGND 0.01769f
C5059 XThR.Tn[13].t53 VGND 0.01937f
C5060 XThR.Tn[13].n49 VGND 0.04938f
C5061 XThR.Tn[13].n50 VGND 0.03469f
C5062 XThR.Tn[13].n52 VGND 0.11133f
C5063 XThR.Tn[13].t41 VGND 0.01775f
C5064 XThR.Tn[13].t17 VGND 0.01944f
C5065 XThR.Tn[13].n53 VGND 0.04746f
C5066 XThR.Tn[13].t58 VGND 0.01769f
C5067 XThR.Tn[13].t73 VGND 0.01937f
C5068 XThR.Tn[13].n54 VGND 0.04938f
C5069 XThR.Tn[13].n55 VGND 0.03469f
C5070 XThR.Tn[13].n57 VGND 0.11133f
C5071 XThR.Tn[13].t63 VGND 0.01775f
C5072 XThR.Tn[13].t55 VGND 0.01944f
C5073 XThR.Tn[13].n58 VGND 0.04746f
C5074 XThR.Tn[13].t15 VGND 0.01769f
C5075 XThR.Tn[13].t45 VGND 0.01937f
C5076 XThR.Tn[13].n59 VGND 0.04938f
C5077 XThR.Tn[13].n60 VGND 0.03469f
C5078 XThR.Tn[13].n62 VGND 0.11133f
C5079 XThR.Tn[13].t31 VGND 0.01775f
C5080 XThR.Tn[13].t27 VGND 0.01944f
C5081 XThR.Tn[13].n63 VGND 0.04746f
C5082 XThR.Tn[13].t46 VGND 0.01769f
C5083 XThR.Tn[13].t20 VGND 0.01937f
C5084 XThR.Tn[13].n64 VGND 0.04938f
C5085 XThR.Tn[13].n65 VGND 0.03469f
C5086 XThR.Tn[13].n67 VGND 0.11133f
C5087 XThR.Tn[13].t50 VGND 0.01775f
C5088 XThR.Tn[13].t40 VGND 0.01944f
C5089 XThR.Tn[13].n68 VGND 0.04746f
C5090 XThR.Tn[13].t67 VGND 0.01769f
C5091 XThR.Tn[13].t36 VGND 0.01937f
C5092 XThR.Tn[13].n69 VGND 0.04938f
C5093 XThR.Tn[13].n70 VGND 0.03469f
C5094 XThR.Tn[13].n72 VGND 0.11133f
C5095 XThR.Tn[13].t69 VGND 0.01775f
C5096 XThR.Tn[13].t62 VGND 0.01944f
C5097 XThR.Tn[13].n73 VGND 0.04746f
C5098 XThR.Tn[13].t23 VGND 0.01769f
C5099 XThR.Tn[13].t54 VGND 0.01937f
C5100 XThR.Tn[13].n74 VGND 0.04938f
C5101 XThR.Tn[13].n75 VGND 0.03469f
C5102 XThR.Tn[13].n77 VGND 0.11133f
C5103 XThR.Tn[13].t42 VGND 0.01775f
C5104 XThR.Tn[13].t56 VGND 0.01944f
C5105 XThR.Tn[13].n78 VGND 0.04746f
C5106 XThR.Tn[13].t61 VGND 0.01769f
C5107 XThR.Tn[13].t47 VGND 0.01937f
C5108 XThR.Tn[13].n79 VGND 0.04938f
C5109 XThR.Tn[13].n80 VGND 0.03469f
C5110 XThR.Tn[13].n82 VGND 0.11133f
C5111 XThR.Tn[13].n83 VGND 0.10118f
C5112 XThR.Tn[13].n84 VGND 0.39667f
C5113 XThR.Tn[13].t6 VGND 0.02271f
C5114 XThR.Tn[13].t4 VGND 0.02271f
C5115 XThR.Tn[13].n85 VGND 0.04907f
C5116 XThR.Tn[13].t7 VGND 0.02271f
C5117 XThR.Tn[13].t5 VGND 0.02271f
C5118 XThR.Tn[13].n86 VGND 0.07469f
C5119 XThR.Tn[13].n87 VGND 0.20738f
C5120 XThR.Tn[13].n88 VGND 0.02777f
C5121 XThC.XTB3.Y.t1 VGND 0.06296f
C5122 XThC.XTB3.Y.n0 VGND 0.04069f
C5123 XThC.XTB3.Y.n1 VGND 0.05192f
C5124 XThC.XTB3.Y.t2 VGND 0.03159f
C5125 XThC.XTB3.Y.t0 VGND 0.03159f
C5126 XThC.XTB3.Y.n2 VGND 0.06782f
C5127 XThC.XTB3.Y.t10 VGND 0.04914f
C5128 XThC.XTB3.Y.t17 VGND 0.02896f
C5129 XThC.XTB3.Y.n3 VGND 0.05852f
C5130 XThC.XTB3.Y.t14 VGND 0.04914f
C5131 XThC.XTB3.Y.t5 VGND 0.02896f
C5132 XThC.XTB3.Y.n4 VGND 0.03012f
C5133 XThC.XTB3.Y.t15 VGND 0.04914f
C5134 XThC.XTB3.Y.t6 VGND 0.02896f
C5135 XThC.XTB3.Y.n5 VGND 0.06469f
C5136 XThC.XTB3.Y.t3 VGND 0.04914f
C5137 XThC.XTB3.Y.t9 VGND 0.02896f
C5138 XThC.XTB3.Y.n6 VGND 0.06006f
C5139 XThC.XTB3.Y.n7 VGND 0.03654f
C5140 XThC.XTB3.Y.n8 VGND 0.06049f
C5141 XThC.XTB3.Y.n9 VGND 0.0234f
C5142 XThC.XTB3.Y.n10 VGND 0.02857f
C5143 XThC.XTB3.Y.n11 VGND 0.06469f
C5144 XThC.XTB3.Y.n12 VGND 0.03243f
C5145 XThC.XTB3.Y.n13 VGND 0.05514f
C5146 XThC.XTB3.Y.t16 VGND 0.04914f
C5147 XThC.XTB3.Y.t7 VGND 0.02896f
C5148 XThC.XTB3.Y.n14 VGND 0.06624f
C5149 XThC.XTB3.Y.t4 VGND 0.04914f
C5150 XThC.XTB3.Y.t13 VGND 0.02896f
C5151 XThC.XTB3.Y.t12 VGND 0.04914f
C5152 XThC.XTB3.Y.t18 VGND 0.02896f
C5153 XThC.XTB3.Y.t11 VGND 0.04914f
C5154 XThC.XTB3.Y.t8 VGND 0.02896f
C5155 XThC.XTB3.Y.n15 VGND 0.08245f
C5156 XThC.XTB3.Y.n16 VGND 0.08709f
C5157 XThC.XTB3.Y.n17 VGND 0.03356f
C5158 XThC.XTB3.Y.n18 VGND 0.07087f
C5159 XThC.XTB3.Y.n19 VGND 0.03243f
C5160 XThC.XTB3.Y.n20 VGND 0.02691f
C5161 XThC.XTB3.Y.n21 VGND 1.39635f
C5162 XThC.XTB3.Y.n22 VGND 0.14933f
C5163 XThR.Tn[8].t6 VGND 0.02288f
C5164 XThR.Tn[8].t4 VGND 0.02288f
C5165 XThR.Tn[8].n0 VGND 0.06947f
C5166 XThR.Tn[8].t7 VGND 0.02288f
C5167 XThR.Tn[8].t5 VGND 0.02288f
C5168 XThR.Tn[8].n1 VGND 0.05086f
C5169 XThR.Tn[8].n2 VGND 0.23126f
C5170 XThR.Tn[8].t11 VGND 0.01487f
C5171 XThR.Tn[8].t8 VGND 0.01487f
C5172 XThR.Tn[8].n3 VGND 0.03709f
C5173 XThR.Tn[8].t1 VGND 0.01487f
C5174 XThR.Tn[8].t2 VGND 0.01487f
C5175 XThR.Tn[8].n4 VGND 0.02974f
C5176 XThR.Tn[8].n5 VGND 0.06858f
C5177 XThR.Tn[8].t39 VGND 0.01788f
C5178 XThR.Tn[8].t33 VGND 0.01958f
C5179 XThR.Tn[8].n6 VGND 0.04781f
C5180 XThR.Tn[8].n7 VGND 0.07431f
C5181 XThR.Tn[8].t59 VGND 0.01788f
C5182 XThR.Tn[8].t49 VGND 0.01958f
C5183 XThR.Tn[8].n8 VGND 0.04781f
C5184 XThR.Tn[8].t13 VGND 0.01782f
C5185 XThR.Tn[8].t45 VGND 0.01952f
C5186 XThR.Tn[8].n9 VGND 0.04975f
C5187 XThR.Tn[8].n10 VGND 0.03495f
C5188 XThR.Tn[8].n12 VGND 0.11215f
C5189 XThR.Tn[8].t34 VGND 0.01788f
C5190 XThR.Tn[8].t26 VGND 0.01958f
C5191 XThR.Tn[8].n13 VGND 0.04781f
C5192 XThR.Tn[8].t53 VGND 0.01782f
C5193 XThR.Tn[8].t22 VGND 0.01952f
C5194 XThR.Tn[8].n14 VGND 0.04975f
C5195 XThR.Tn[8].n15 VGND 0.03495f
C5196 XThR.Tn[8].n17 VGND 0.11215f
C5197 XThR.Tn[8].t50 VGND 0.01788f
C5198 XThR.Tn[8].t43 VGND 0.01958f
C5199 XThR.Tn[8].n18 VGND 0.04781f
C5200 XThR.Tn[8].t65 VGND 0.01782f
C5201 XThR.Tn[8].t40 VGND 0.01952f
C5202 XThR.Tn[8].n19 VGND 0.04975f
C5203 XThR.Tn[8].n20 VGND 0.03495f
C5204 XThR.Tn[8].n22 VGND 0.11215f
C5205 XThR.Tn[8].t12 VGND 0.01788f
C5206 XThR.Tn[8].t70 VGND 0.01958f
C5207 XThR.Tn[8].n23 VGND 0.04781f
C5208 XThR.Tn[8].t36 VGND 0.01782f
C5209 XThR.Tn[8].t66 VGND 0.01952f
C5210 XThR.Tn[8].n24 VGND 0.04975f
C5211 XThR.Tn[8].n25 VGND 0.03495f
C5212 XThR.Tn[8].n27 VGND 0.11215f
C5213 XThR.Tn[8].t52 VGND 0.01788f
C5214 XThR.Tn[8].t44 VGND 0.01958f
C5215 XThR.Tn[8].n28 VGND 0.04781f
C5216 XThR.Tn[8].t68 VGND 0.01782f
C5217 XThR.Tn[8].t41 VGND 0.01952f
C5218 XThR.Tn[8].n29 VGND 0.04975f
C5219 XThR.Tn[8].n30 VGND 0.03495f
C5220 XThR.Tn[8].n32 VGND 0.11215f
C5221 XThR.Tn[8].t28 VGND 0.01788f
C5222 XThR.Tn[8].t61 VGND 0.01958f
C5223 XThR.Tn[8].n33 VGND 0.04781f
C5224 XThR.Tn[8].t47 VGND 0.01782f
C5225 XThR.Tn[8].t58 VGND 0.01952f
C5226 XThR.Tn[8].n34 VGND 0.04975f
C5227 XThR.Tn[8].n35 VGND 0.03495f
C5228 XThR.Tn[8].n37 VGND 0.11215f
C5229 XThR.Tn[8].t60 VGND 0.01788f
C5230 XThR.Tn[8].t56 VGND 0.01958f
C5231 XThR.Tn[8].n38 VGND 0.04781f
C5232 XThR.Tn[8].t14 VGND 0.01782f
C5233 XThR.Tn[8].t51 VGND 0.01952f
C5234 XThR.Tn[8].n39 VGND 0.04975f
C5235 XThR.Tn[8].n40 VGND 0.03495f
C5236 XThR.Tn[8].n42 VGND 0.11215f
C5237 XThR.Tn[8].t63 VGND 0.01788f
C5238 XThR.Tn[8].t69 VGND 0.01958f
C5239 XThR.Tn[8].n43 VGND 0.04781f
C5240 XThR.Tn[8].t20 VGND 0.01782f
C5241 XThR.Tn[8].t64 VGND 0.01952f
C5242 XThR.Tn[8].n44 VGND 0.04975f
C5243 XThR.Tn[8].n45 VGND 0.03495f
C5244 XThR.Tn[8].n47 VGND 0.11215f
C5245 XThR.Tn[8].t17 VGND 0.01788f
C5246 XThR.Tn[8].t27 VGND 0.01958f
C5247 XThR.Tn[8].n48 VGND 0.04781f
C5248 XThR.Tn[8].t38 VGND 0.01782f
C5249 XThR.Tn[8].t24 VGND 0.01952f
C5250 XThR.Tn[8].n49 VGND 0.04975f
C5251 XThR.Tn[8].n50 VGND 0.03495f
C5252 XThR.Tn[8].n52 VGND 0.11215f
C5253 XThR.Tn[8].t72 VGND 0.01788f
C5254 XThR.Tn[8].t46 VGND 0.01958f
C5255 XThR.Tn[8].n53 VGND 0.04781f
C5256 XThR.Tn[8].t31 VGND 0.01782f
C5257 XThR.Tn[8].t42 VGND 0.01952f
C5258 XThR.Tn[8].n54 VGND 0.04975f
C5259 XThR.Tn[8].n55 VGND 0.03495f
C5260 XThR.Tn[8].n57 VGND 0.11215f
C5261 XThR.Tn[8].t30 VGND 0.01788f
C5262 XThR.Tn[8].t21 VGND 0.01958f
C5263 XThR.Tn[8].n58 VGND 0.04781f
C5264 XThR.Tn[8].t48 VGND 0.01782f
C5265 XThR.Tn[8].t16 VGND 0.01952f
C5266 XThR.Tn[8].n59 VGND 0.04975f
C5267 XThR.Tn[8].n60 VGND 0.03495f
C5268 XThR.Tn[8].n62 VGND 0.11215f
C5269 XThR.Tn[8].t62 VGND 0.01788f
C5270 XThR.Tn[8].t57 VGND 0.01958f
C5271 XThR.Tn[8].n63 VGND 0.04781f
C5272 XThR.Tn[8].t18 VGND 0.01782f
C5273 XThR.Tn[8].t54 VGND 0.01952f
C5274 XThR.Tn[8].n64 VGND 0.04975f
C5275 XThR.Tn[8].n65 VGND 0.03495f
C5276 XThR.Tn[8].n67 VGND 0.11215f
C5277 XThR.Tn[8].t15 VGND 0.01788f
C5278 XThR.Tn[8].t71 VGND 0.01958f
C5279 XThR.Tn[8].n68 VGND 0.04781f
C5280 XThR.Tn[8].t37 VGND 0.01782f
C5281 XThR.Tn[8].t67 VGND 0.01952f
C5282 XThR.Tn[8].n69 VGND 0.04975f
C5283 XThR.Tn[8].n70 VGND 0.03495f
C5284 XThR.Tn[8].n72 VGND 0.11215f
C5285 XThR.Tn[8].t35 VGND 0.01788f
C5286 XThR.Tn[8].t29 VGND 0.01958f
C5287 XThR.Tn[8].n73 VGND 0.04781f
C5288 XThR.Tn[8].t55 VGND 0.01782f
C5289 XThR.Tn[8].t25 VGND 0.01952f
C5290 XThR.Tn[8].n74 VGND 0.04975f
C5291 XThR.Tn[8].n75 VGND 0.03495f
C5292 XThR.Tn[8].n77 VGND 0.11215f
C5293 XThR.Tn[8].t73 VGND 0.01788f
C5294 XThR.Tn[8].t23 VGND 0.01958f
C5295 XThR.Tn[8].n78 VGND 0.04781f
C5296 XThR.Tn[8].t32 VGND 0.01782f
C5297 XThR.Tn[8].t19 VGND 0.01952f
C5298 XThR.Tn[8].n79 VGND 0.04975f
C5299 XThR.Tn[8].n80 VGND 0.03495f
C5300 XThR.Tn[8].n82 VGND 0.11215f
C5301 XThR.Tn[8].n83 VGND 0.10193f
C5302 XThR.Tn[8].n84 VGND 0.31231f
C5303 XThR.Tn[8].t3 VGND 0.02288f
C5304 XThR.Tn[8].t10 VGND 0.02288f
C5305 XThR.Tn[8].n85 VGND 0.04943f
C5306 XThR.Tn[8].t9 VGND 0.02288f
C5307 XThR.Tn[8].t0 VGND 0.02288f
C5308 XThR.Tn[8].n86 VGND 0.07524f
C5309 XThR.Tn[8].n87 VGND 0.20891f
C5310 XThR.Tn[8].n88 VGND 0.0103f
C5311 XThR.Tn[0].t5 VGND 0.0212f
C5312 XThR.Tn[0].t6 VGND 0.0212f
C5313 XThR.Tn[0].n0 VGND 0.04279f
C5314 XThR.Tn[0].t4 VGND 0.0212f
C5315 XThR.Tn[0].t3 VGND 0.0212f
C5316 XThR.Tn[0].n1 VGND 0.05007f
C5317 XThR.Tn[0].n2 VGND 0.15019f
C5318 XThR.Tn[0].t8 VGND 0.01378f
C5319 XThR.Tn[0].t9 VGND 0.01378f
C5320 XThR.Tn[0].n3 VGND 0.03138f
C5321 XThR.Tn[0].t7 VGND 0.01378f
C5322 XThR.Tn[0].t10 VGND 0.01378f
C5323 XThR.Tn[0].n4 VGND 0.03138f
C5324 XThR.Tn[0].t11 VGND 0.01378f
C5325 XThR.Tn[0].t2 VGND 0.01378f
C5326 XThR.Tn[0].n5 VGND 0.05229f
C5327 XThR.Tn[0].t0 VGND 0.01378f
C5328 XThR.Tn[0].t1 VGND 0.01378f
C5329 XThR.Tn[0].n6 VGND 0.03138f
C5330 XThR.Tn[0].n7 VGND 0.14945f
C5331 XThR.Tn[0].n8 VGND 0.09239f
C5332 XThR.Tn[0].n9 VGND 0.10426f
C5333 XThR.Tn[0].t48 VGND 0.01657f
C5334 XThR.Tn[0].t40 VGND 0.01814f
C5335 XThR.Tn[0].n10 VGND 0.04431f
C5336 XThR.Tn[0].n11 VGND 0.06885f
C5337 XThR.Tn[0].t67 VGND 0.01657f
C5338 XThR.Tn[0].t58 VGND 0.01814f
C5339 XThR.Tn[0].n12 VGND 0.04431f
C5340 XThR.Tn[0].t24 VGND 0.01652f
C5341 XThR.Tn[0].t50 VGND 0.01809f
C5342 XThR.Tn[0].n13 VGND 0.0461f
C5343 XThR.Tn[0].n14 VGND 0.03239f
C5344 XThR.Tn[0].n16 VGND 0.10393f
C5345 XThR.Tn[0].t41 VGND 0.01657f
C5346 XThR.Tn[0].t33 VGND 0.01814f
C5347 XThR.Tn[0].n17 VGND 0.04431f
C5348 XThR.Tn[0].t61 VGND 0.01652f
C5349 XThR.Tn[0].t26 VGND 0.01809f
C5350 XThR.Tn[0].n18 VGND 0.0461f
C5351 XThR.Tn[0].n19 VGND 0.03239f
C5352 XThR.Tn[0].n21 VGND 0.10393f
C5353 XThR.Tn[0].t59 VGND 0.01657f
C5354 XThR.Tn[0].t51 VGND 0.01814f
C5355 XThR.Tn[0].n22 VGND 0.04431f
C5356 XThR.Tn[0].t12 VGND 0.01652f
C5357 XThR.Tn[0].t44 VGND 0.01809f
C5358 XThR.Tn[0].n23 VGND 0.0461f
C5359 XThR.Tn[0].n24 VGND 0.03239f
C5360 XThR.Tn[0].n26 VGND 0.10393f
C5361 XThR.Tn[0].t21 VGND 0.01657f
C5362 XThR.Tn[0].t15 VGND 0.01814f
C5363 XThR.Tn[0].n27 VGND 0.04431f
C5364 XThR.Tn[0].t43 VGND 0.01652f
C5365 XThR.Tn[0].t72 VGND 0.01809f
C5366 XThR.Tn[0].n28 VGND 0.0461f
C5367 XThR.Tn[0].n29 VGND 0.03239f
C5368 XThR.Tn[0].n31 VGND 0.10393f
C5369 XThR.Tn[0].t60 VGND 0.01657f
C5370 XThR.Tn[0].t52 VGND 0.01814f
C5371 XThR.Tn[0].n32 VGND 0.04431f
C5372 XThR.Tn[0].t13 VGND 0.01652f
C5373 XThR.Tn[0].t46 VGND 0.01809f
C5374 XThR.Tn[0].n33 VGND 0.0461f
C5375 XThR.Tn[0].n34 VGND 0.03239f
C5376 XThR.Tn[0].n36 VGND 0.10393f
C5377 XThR.Tn[0].t35 VGND 0.01657f
C5378 XThR.Tn[0].t68 VGND 0.01814f
C5379 XThR.Tn[0].n37 VGND 0.04431f
C5380 XThR.Tn[0].t54 VGND 0.01652f
C5381 XThR.Tn[0].t64 VGND 0.01809f
C5382 XThR.Tn[0].n38 VGND 0.0461f
C5383 XThR.Tn[0].n39 VGND 0.03239f
C5384 XThR.Tn[0].n41 VGND 0.10393f
C5385 XThR.Tn[0].t66 VGND 0.01657f
C5386 XThR.Tn[0].t63 VGND 0.01814f
C5387 XThR.Tn[0].n42 VGND 0.04431f
C5388 XThR.Tn[0].t23 VGND 0.01652f
C5389 XThR.Tn[0].t55 VGND 0.01809f
C5390 XThR.Tn[0].n43 VGND 0.0461f
C5391 XThR.Tn[0].n44 VGND 0.03239f
C5392 XThR.Tn[0].n46 VGND 0.10393f
C5393 XThR.Tn[0].t70 VGND 0.01657f
C5394 XThR.Tn[0].t14 VGND 0.01814f
C5395 XThR.Tn[0].n47 VGND 0.04431f
C5396 XThR.Tn[0].t28 VGND 0.01652f
C5397 XThR.Tn[0].t71 VGND 0.01809f
C5398 XThR.Tn[0].n48 VGND 0.0461f
C5399 XThR.Tn[0].n49 VGND 0.03239f
C5400 XThR.Tn[0].n51 VGND 0.10393f
C5401 XThR.Tn[0].t25 VGND 0.01657f
C5402 XThR.Tn[0].t34 VGND 0.01814f
C5403 XThR.Tn[0].n52 VGND 0.04431f
C5404 XThR.Tn[0].t47 VGND 0.01652f
C5405 XThR.Tn[0].t29 VGND 0.01809f
C5406 XThR.Tn[0].n53 VGND 0.0461f
C5407 XThR.Tn[0].n54 VGND 0.03239f
C5408 XThR.Tn[0].n56 VGND 0.10393f
C5409 XThR.Tn[0].t17 VGND 0.01657f
C5410 XThR.Tn[0].t53 VGND 0.01814f
C5411 XThR.Tn[0].n57 VGND 0.04431f
C5412 XThR.Tn[0].t38 VGND 0.01652f
C5413 XThR.Tn[0].t49 VGND 0.01809f
C5414 XThR.Tn[0].n58 VGND 0.0461f
C5415 XThR.Tn[0].n59 VGND 0.03239f
C5416 XThR.Tn[0].n61 VGND 0.10393f
C5417 XThR.Tn[0].t37 VGND 0.01657f
C5418 XThR.Tn[0].t31 VGND 0.01814f
C5419 XThR.Tn[0].n62 VGND 0.04431f
C5420 XThR.Tn[0].t56 VGND 0.01652f
C5421 XThR.Tn[0].t19 VGND 0.01809f
C5422 XThR.Tn[0].n63 VGND 0.0461f
C5423 XThR.Tn[0].n64 VGND 0.03239f
C5424 XThR.Tn[0].n66 VGND 0.10393f
C5425 XThR.Tn[0].t69 VGND 0.01657f
C5426 XThR.Tn[0].t65 VGND 0.01814f
C5427 XThR.Tn[0].n67 VGND 0.04431f
C5428 XThR.Tn[0].t27 VGND 0.01652f
C5429 XThR.Tn[0].t57 VGND 0.01809f
C5430 XThR.Tn[0].n68 VGND 0.0461f
C5431 XThR.Tn[0].n69 VGND 0.03239f
C5432 XThR.Tn[0].n71 VGND 0.10393f
C5433 XThR.Tn[0].t22 VGND 0.01657f
C5434 XThR.Tn[0].t16 VGND 0.01814f
C5435 XThR.Tn[0].n72 VGND 0.04431f
C5436 XThR.Tn[0].t45 VGND 0.01652f
C5437 XThR.Tn[0].t73 VGND 0.01809f
C5438 XThR.Tn[0].n73 VGND 0.0461f
C5439 XThR.Tn[0].n74 VGND 0.03239f
C5440 XThR.Tn[0].n76 VGND 0.10393f
C5441 XThR.Tn[0].t42 VGND 0.01657f
C5442 XThR.Tn[0].t36 VGND 0.01814f
C5443 XThR.Tn[0].n77 VGND 0.04431f
C5444 XThR.Tn[0].t62 VGND 0.01652f
C5445 XThR.Tn[0].t30 VGND 0.01809f
C5446 XThR.Tn[0].n78 VGND 0.0461f
C5447 XThR.Tn[0].n79 VGND 0.03239f
C5448 XThR.Tn[0].n81 VGND 0.10393f
C5449 XThR.Tn[0].t18 VGND 0.01657f
C5450 XThR.Tn[0].t32 VGND 0.01814f
C5451 XThR.Tn[0].n82 VGND 0.04431f
C5452 XThR.Tn[0].t39 VGND 0.01652f
C5453 XThR.Tn[0].t20 VGND 0.01809f
C5454 XThR.Tn[0].n83 VGND 0.0461f
C5455 XThR.Tn[0].n84 VGND 0.03239f
C5456 XThR.Tn[0].n86 VGND 0.10393f
C5457 XThR.Tn[0].n87 VGND 0.09445f
C5458 XThR.Tn[0].n88 VGND 0.27043f
C5459 XThR.Tn[7].t2 VGND 0.01406f
C5460 XThR.Tn[7].t1 VGND 0.01406f
C5461 XThR.Tn[7].n0 VGND 0.03105f
C5462 XThR.Tn[7].t3 VGND 0.01406f
C5463 XThR.Tn[7].t0 VGND 0.01406f
C5464 XThR.Tn[7].n1 VGND 0.04338f
C5465 XThR.Tn[7].n2 VGND 0.15921f
C5466 XThR.Tn[7].t6 VGND 0.02163f
C5467 XThR.Tn[7].t7 VGND 0.02163f
C5468 XThR.Tn[7].n3 VGND 0.06585f
C5469 XThR.Tn[7].t5 VGND 0.02163f
C5470 XThR.Tn[7].t4 VGND 0.02163f
C5471 XThR.Tn[7].n4 VGND 0.04791f
C5472 XThR.Tn[7].n5 VGND 0.21081f
C5473 XThR.Tn[7].n6 VGND 0.02627f
C5474 XThR.Tn[7].t53 VGND 0.0169f
C5475 XThR.Tn[7].t45 VGND 0.01851f
C5476 XThR.Tn[7].n7 VGND 0.04519f
C5477 XThR.Tn[7].n8 VGND 0.07023f
C5478 XThR.Tn[7].t8 VGND 0.0169f
C5479 XThR.Tn[7].t60 VGND 0.01851f
C5480 XThR.Tn[7].n9 VGND 0.04519f
C5481 XThR.Tn[7].t26 VGND 0.01685f
C5482 XThR.Tn[7].t38 VGND 0.01845f
C5483 XThR.Tn[7].n10 VGND 0.04702f
C5484 XThR.Tn[7].n11 VGND 0.03304f
C5485 XThR.Tn[7].n13 VGND 0.10601f
C5486 XThR.Tn[7].t47 VGND 0.0169f
C5487 XThR.Tn[7].t37 VGND 0.01851f
C5488 XThR.Tn[7].n14 VGND 0.04519f
C5489 XThR.Tn[7].t66 VGND 0.01685f
C5490 XThR.Tn[7].t15 VGND 0.01845f
C5491 XThR.Tn[7].n15 VGND 0.04702f
C5492 XThR.Tn[7].n16 VGND 0.03304f
C5493 XThR.Tn[7].n18 VGND 0.10601f
C5494 XThR.Tn[7].t62 VGND 0.0169f
C5495 XThR.Tn[7].t55 VGND 0.01851f
C5496 XThR.Tn[7].n19 VGND 0.04519f
C5497 XThR.Tn[7].t18 VGND 0.01685f
C5498 XThR.Tn[7].t32 VGND 0.01845f
C5499 XThR.Tn[7].n20 VGND 0.04702f
C5500 XThR.Tn[7].n21 VGND 0.03304f
C5501 XThR.Tn[7].n23 VGND 0.10601f
C5502 XThR.Tn[7].t25 VGND 0.0169f
C5503 XThR.Tn[7].t21 VGND 0.01851f
C5504 XThR.Tn[7].n24 VGND 0.04519f
C5505 XThR.Tn[7].t50 VGND 0.01685f
C5506 XThR.Tn[7].t63 VGND 0.01845f
C5507 XThR.Tn[7].n25 VGND 0.04702f
C5508 XThR.Tn[7].n26 VGND 0.03304f
C5509 XThR.Tn[7].n28 VGND 0.10601f
C5510 XThR.Tn[7].t65 VGND 0.0169f
C5511 XThR.Tn[7].t56 VGND 0.01851f
C5512 XThR.Tn[7].n29 VGND 0.04519f
C5513 XThR.Tn[7].t19 VGND 0.01685f
C5514 XThR.Tn[7].t34 VGND 0.01845f
C5515 XThR.Tn[7].n30 VGND 0.04702f
C5516 XThR.Tn[7].n31 VGND 0.03304f
C5517 XThR.Tn[7].n33 VGND 0.10601f
C5518 XThR.Tn[7].t40 VGND 0.0169f
C5519 XThR.Tn[7].t11 VGND 0.01851f
C5520 XThR.Tn[7].n34 VGND 0.04519f
C5521 XThR.Tn[7].t58 VGND 0.01685f
C5522 XThR.Tn[7].t54 VGND 0.01845f
C5523 XThR.Tn[7].n35 VGND 0.04702f
C5524 XThR.Tn[7].n36 VGND 0.03304f
C5525 XThR.Tn[7].n38 VGND 0.10601f
C5526 XThR.Tn[7].t9 VGND 0.0169f
C5527 XThR.Tn[7].t68 VGND 0.01851f
C5528 XThR.Tn[7].n39 VGND 0.04519f
C5529 XThR.Tn[7].t27 VGND 0.01685f
C5530 XThR.Tn[7].t46 VGND 0.01845f
C5531 XThR.Tn[7].n40 VGND 0.04702f
C5532 XThR.Tn[7].n41 VGND 0.03304f
C5533 XThR.Tn[7].n43 VGND 0.10601f
C5534 XThR.Tn[7].t14 VGND 0.0169f
C5535 XThR.Tn[7].t20 VGND 0.01851f
C5536 XThR.Tn[7].n44 VGND 0.04519f
C5537 XThR.Tn[7].t31 VGND 0.01685f
C5538 XThR.Tn[7].t61 VGND 0.01845f
C5539 XThR.Tn[7].n45 VGND 0.04702f
C5540 XThR.Tn[7].n46 VGND 0.03304f
C5541 XThR.Tn[7].n48 VGND 0.10601f
C5542 XThR.Tn[7].t29 VGND 0.0169f
C5543 XThR.Tn[7].t39 VGND 0.01851f
C5544 XThR.Tn[7].n49 VGND 0.04519f
C5545 XThR.Tn[7].t52 VGND 0.01685f
C5546 XThR.Tn[7].t16 VGND 0.01845f
C5547 XThR.Tn[7].n50 VGND 0.04702f
C5548 XThR.Tn[7].n51 VGND 0.03304f
C5549 XThR.Tn[7].n53 VGND 0.10601f
C5550 XThR.Tn[7].t23 VGND 0.0169f
C5551 XThR.Tn[7].t57 VGND 0.01851f
C5552 XThR.Tn[7].n54 VGND 0.04519f
C5553 XThR.Tn[7].t43 VGND 0.01685f
C5554 XThR.Tn[7].t36 VGND 0.01845f
C5555 XThR.Tn[7].n55 VGND 0.04702f
C5556 XThR.Tn[7].n56 VGND 0.03304f
C5557 XThR.Tn[7].n58 VGND 0.10601f
C5558 XThR.Tn[7].t42 VGND 0.0169f
C5559 XThR.Tn[7].t33 VGND 0.01851f
C5560 XThR.Tn[7].n59 VGND 0.04519f
C5561 XThR.Tn[7].t59 VGND 0.01685f
C5562 XThR.Tn[7].t10 VGND 0.01845f
C5563 XThR.Tn[7].n60 VGND 0.04702f
C5564 XThR.Tn[7].n61 VGND 0.03304f
C5565 XThR.Tn[7].n63 VGND 0.10601f
C5566 XThR.Tn[7].t12 VGND 0.0169f
C5567 XThR.Tn[7].t69 VGND 0.01851f
C5568 XThR.Tn[7].n64 VGND 0.04519f
C5569 XThR.Tn[7].t30 VGND 0.01685f
C5570 XThR.Tn[7].t48 VGND 0.01845f
C5571 XThR.Tn[7].n65 VGND 0.04702f
C5572 XThR.Tn[7].n66 VGND 0.03304f
C5573 XThR.Tn[7].n68 VGND 0.10601f
C5574 XThR.Tn[7].t28 VGND 0.0169f
C5575 XThR.Tn[7].t22 VGND 0.01851f
C5576 XThR.Tn[7].n69 VGND 0.04519f
C5577 XThR.Tn[7].t51 VGND 0.01685f
C5578 XThR.Tn[7].t64 VGND 0.01845f
C5579 XThR.Tn[7].n70 VGND 0.04702f
C5580 XThR.Tn[7].n71 VGND 0.03304f
C5581 XThR.Tn[7].n73 VGND 0.10601f
C5582 XThR.Tn[7].t49 VGND 0.0169f
C5583 XThR.Tn[7].t41 VGND 0.01851f
C5584 XThR.Tn[7].n74 VGND 0.04519f
C5585 XThR.Tn[7].t67 VGND 0.01685f
C5586 XThR.Tn[7].t17 VGND 0.01845f
C5587 XThR.Tn[7].n75 VGND 0.04702f
C5588 XThR.Tn[7].n76 VGND 0.03304f
C5589 XThR.Tn[7].n78 VGND 0.10601f
C5590 XThR.Tn[7].t24 VGND 0.0169f
C5591 XThR.Tn[7].t35 VGND 0.01851f
C5592 XThR.Tn[7].n79 VGND 0.04519f
C5593 XThR.Tn[7].t44 VGND 0.01685f
C5594 XThR.Tn[7].t13 VGND 0.01845f
C5595 XThR.Tn[7].n80 VGND 0.04702f
C5596 XThR.Tn[7].n81 VGND 0.03304f
C5597 XThR.Tn[7].n83 VGND 0.10601f
C5598 XThR.Tn[7].n84 VGND 0.09634f
C5599 XThR.Tn[7].n85 VGND 0.39109f
C5600 XThR.Tn[11].t8 VGND 0.02263f
C5601 XThR.Tn[11].t10 VGND 0.02263f
C5602 XThR.Tn[11].n0 VGND 0.06871f
C5603 XThR.Tn[11].t9 VGND 0.02263f
C5604 XThR.Tn[11].t11 VGND 0.02263f
C5605 XThR.Tn[11].n1 VGND 0.05031f
C5606 XThR.Tn[11].n2 VGND 0.22874f
C5607 XThR.Tn[11].t7 VGND 0.01471f
C5608 XThR.Tn[11].t5 VGND 0.01471f
C5609 XThR.Tn[11].n3 VGND 0.03669f
C5610 XThR.Tn[11].t6 VGND 0.01471f
C5611 XThR.Tn[11].t4 VGND 0.01471f
C5612 XThR.Tn[11].n4 VGND 0.02942f
C5613 XThR.Tn[11].n5 VGND 0.07401f
C5614 XThR.Tn[11].t56 VGND 0.01769f
C5615 XThR.Tn[11].t48 VGND 0.01937f
C5616 XThR.Tn[11].n6 VGND 0.04729f
C5617 XThR.Tn[11].n7 VGND 0.0735f
C5618 XThR.Tn[11].t12 VGND 0.01769f
C5619 XThR.Tn[11].t67 VGND 0.01937f
C5620 XThR.Tn[11].n8 VGND 0.04729f
C5621 XThR.Tn[11].t27 VGND 0.01763f
C5622 XThR.Tn[11].t58 VGND 0.0193f
C5623 XThR.Tn[11].n9 VGND 0.04921f
C5624 XThR.Tn[11].n10 VGND 0.03457f
C5625 XThR.Tn[11].n12 VGND 0.11093f
C5626 XThR.Tn[11].t49 VGND 0.01769f
C5627 XThR.Tn[11].t41 VGND 0.01937f
C5628 XThR.Tn[11].n13 VGND 0.04729f
C5629 XThR.Tn[11].t65 VGND 0.01763f
C5630 XThR.Tn[11].t36 VGND 0.0193f
C5631 XThR.Tn[11].n14 VGND 0.04921f
C5632 XThR.Tn[11].n15 VGND 0.03457f
C5633 XThR.Tn[11].n17 VGND 0.11093f
C5634 XThR.Tn[11].t68 VGND 0.01769f
C5635 XThR.Tn[11].t60 VGND 0.01937f
C5636 XThR.Tn[11].n18 VGND 0.04729f
C5637 XThR.Tn[11].t18 VGND 0.01763f
C5638 XThR.Tn[11].t54 VGND 0.0193f
C5639 XThR.Tn[11].n19 VGND 0.04921f
C5640 XThR.Tn[11].n20 VGND 0.03457f
C5641 XThR.Tn[11].n22 VGND 0.11093f
C5642 XThR.Tn[11].t33 VGND 0.01769f
C5643 XThR.Tn[11].t23 VGND 0.01937f
C5644 XThR.Tn[11].n23 VGND 0.04729f
C5645 XThR.Tn[11].t50 VGND 0.01763f
C5646 XThR.Tn[11].t19 VGND 0.0193f
C5647 XThR.Tn[11].n24 VGND 0.04921f
C5648 XThR.Tn[11].n25 VGND 0.03457f
C5649 XThR.Tn[11].n27 VGND 0.11093f
C5650 XThR.Tn[11].t70 VGND 0.01769f
C5651 XThR.Tn[11].t62 VGND 0.01937f
C5652 XThR.Tn[11].n28 VGND 0.04729f
C5653 XThR.Tn[11].t21 VGND 0.01763f
C5654 XThR.Tn[11].t55 VGND 0.0193f
C5655 XThR.Tn[11].n29 VGND 0.04921f
C5656 XThR.Tn[11].n30 VGND 0.03457f
C5657 XThR.Tn[11].n32 VGND 0.11093f
C5658 XThR.Tn[11].t44 VGND 0.01769f
C5659 XThR.Tn[11].t14 VGND 0.01937f
C5660 XThR.Tn[11].n33 VGND 0.04729f
C5661 XThR.Tn[11].t59 VGND 0.01763f
C5662 XThR.Tn[11].t72 VGND 0.0193f
C5663 XThR.Tn[11].n34 VGND 0.04921f
C5664 XThR.Tn[11].n35 VGND 0.03457f
C5665 XThR.Tn[11].n37 VGND 0.11093f
C5666 XThR.Tn[11].t13 VGND 0.01769f
C5667 XThR.Tn[11].t71 VGND 0.01937f
C5668 XThR.Tn[11].n38 VGND 0.04729f
C5669 XThR.Tn[11].t28 VGND 0.01763f
C5670 XThR.Tn[11].t64 VGND 0.0193f
C5671 XThR.Tn[11].n39 VGND 0.04921f
C5672 XThR.Tn[11].n40 VGND 0.03457f
C5673 XThR.Tn[11].n42 VGND 0.11093f
C5674 XThR.Tn[11].t16 VGND 0.01769f
C5675 XThR.Tn[11].t22 VGND 0.01937f
C5676 XThR.Tn[11].n43 VGND 0.04729f
C5677 XThR.Tn[11].t32 VGND 0.01763f
C5678 XThR.Tn[11].t17 VGND 0.0193f
C5679 XThR.Tn[11].n44 VGND 0.04921f
C5680 XThR.Tn[11].n45 VGND 0.03457f
C5681 XThR.Tn[11].n47 VGND 0.11093f
C5682 XThR.Tn[11].t35 VGND 0.01769f
C5683 XThR.Tn[11].t43 VGND 0.01937f
C5684 XThR.Tn[11].n48 VGND 0.04729f
C5685 XThR.Tn[11].t52 VGND 0.01763f
C5686 XThR.Tn[11].t37 VGND 0.0193f
C5687 XThR.Tn[11].n49 VGND 0.04921f
C5688 XThR.Tn[11].n50 VGND 0.03457f
C5689 XThR.Tn[11].n52 VGND 0.11093f
C5690 XThR.Tn[11].t25 VGND 0.01769f
C5691 XThR.Tn[11].t63 VGND 0.01937f
C5692 XThR.Tn[11].n53 VGND 0.04729f
C5693 XThR.Tn[11].t42 VGND 0.01763f
C5694 XThR.Tn[11].t57 VGND 0.0193f
C5695 XThR.Tn[11].n54 VGND 0.04921f
C5696 XThR.Tn[11].n55 VGND 0.03457f
C5697 XThR.Tn[11].n57 VGND 0.11093f
C5698 XThR.Tn[11].t47 VGND 0.01769f
C5699 XThR.Tn[11].t39 VGND 0.01937f
C5700 XThR.Tn[11].n58 VGND 0.04729f
C5701 XThR.Tn[11].t61 VGND 0.01763f
C5702 XThR.Tn[11].t29 VGND 0.0193f
C5703 XThR.Tn[11].n59 VGND 0.04921f
C5704 XThR.Tn[11].n60 VGND 0.03457f
C5705 XThR.Tn[11].n62 VGND 0.11093f
C5706 XThR.Tn[11].t15 VGND 0.01769f
C5707 XThR.Tn[11].t73 VGND 0.01937f
C5708 XThR.Tn[11].n63 VGND 0.04729f
C5709 XThR.Tn[11].t30 VGND 0.01763f
C5710 XThR.Tn[11].t66 VGND 0.0193f
C5711 XThR.Tn[11].n64 VGND 0.04921f
C5712 XThR.Tn[11].n65 VGND 0.03457f
C5713 XThR.Tn[11].n67 VGND 0.11093f
C5714 XThR.Tn[11].t34 VGND 0.01769f
C5715 XThR.Tn[11].t24 VGND 0.01937f
C5716 XThR.Tn[11].n68 VGND 0.04729f
C5717 XThR.Tn[11].t51 VGND 0.01763f
C5718 XThR.Tn[11].t20 VGND 0.0193f
C5719 XThR.Tn[11].n69 VGND 0.04921f
C5720 XThR.Tn[11].n70 VGND 0.03457f
C5721 XThR.Tn[11].n72 VGND 0.11093f
C5722 XThR.Tn[11].t53 VGND 0.01769f
C5723 XThR.Tn[11].t46 VGND 0.01937f
C5724 XThR.Tn[11].n73 VGND 0.04729f
C5725 XThR.Tn[11].t69 VGND 0.01763f
C5726 XThR.Tn[11].t38 VGND 0.0193f
C5727 XThR.Tn[11].n74 VGND 0.04921f
C5728 XThR.Tn[11].n75 VGND 0.03457f
C5729 XThR.Tn[11].n77 VGND 0.11093f
C5730 XThR.Tn[11].t26 VGND 0.01769f
C5731 XThR.Tn[11].t40 VGND 0.01937f
C5732 XThR.Tn[11].n78 VGND 0.04729f
C5733 XThR.Tn[11].t45 VGND 0.01763f
C5734 XThR.Tn[11].t31 VGND 0.0193f
C5735 XThR.Tn[11].n79 VGND 0.04921f
C5736 XThR.Tn[11].n80 VGND 0.03457f
C5737 XThR.Tn[11].n82 VGND 0.11093f
C5738 XThR.Tn[11].n83 VGND 0.10081f
C5739 XThR.Tn[11].n84 VGND 0.36131f
C5740 XThR.Tn[11].t0 VGND 0.02263f
C5741 XThR.Tn[11].t2 VGND 0.02263f
C5742 XThR.Tn[11].n85 VGND 0.0489f
C5743 XThR.Tn[11].t1 VGND 0.02263f
C5744 XThR.Tn[11].t3 VGND 0.02263f
C5745 XThR.Tn[11].n86 VGND 0.07442f
C5746 XThR.Tn[11].n87 VGND 0.20663f
C5747 XThR.Tn[11].n88 VGND 0.02767f
C5748 XThR.Tn[4].t1 VGND 0.02192f
C5749 XThR.Tn[4].t2 VGND 0.02192f
C5750 XThR.Tn[4].n0 VGND 0.04424f
C5751 XThR.Tn[4].t0 VGND 0.02192f
C5752 XThR.Tn[4].t3 VGND 0.02192f
C5753 XThR.Tn[4].n1 VGND 0.05176f
C5754 XThR.Tn[4].n2 VGND 0.15526f
C5755 XThR.Tn[4].t8 VGND 0.01425f
C5756 XThR.Tn[4].t9 VGND 0.01425f
C5757 XThR.Tn[4].n3 VGND 0.05405f
C5758 XThR.Tn[4].t11 VGND 0.01425f
C5759 XThR.Tn[4].t10 VGND 0.01425f
C5760 XThR.Tn[4].n4 VGND 0.03244f
C5761 XThR.Tn[4].n5 VGND 0.15449f
C5762 XThR.Tn[4].t6 VGND 0.01425f
C5763 XThR.Tn[4].t5 VGND 0.01425f
C5764 XThR.Tn[4].n6 VGND 0.03244f
C5765 XThR.Tn[4].n7 VGND 0.0955f
C5766 XThR.Tn[4].t7 VGND 0.01425f
C5767 XThR.Tn[4].t4 VGND 0.01425f
C5768 XThR.Tn[4].n8 VGND 0.03244f
C5769 XThR.Tn[4].n9 VGND 0.10778f
C5770 XThR.Tn[4].t44 VGND 0.01713f
C5771 XThR.Tn[4].t38 VGND 0.01876f
C5772 XThR.Tn[4].n10 VGND 0.0458f
C5773 XThR.Tn[4].n11 VGND 0.07118f
C5774 XThR.Tn[4].t65 VGND 0.01713f
C5775 XThR.Tn[4].t54 VGND 0.01876f
C5776 XThR.Tn[4].n12 VGND 0.0458f
C5777 XThR.Tn[4].t19 VGND 0.01707f
C5778 XThR.Tn[4].t50 VGND 0.0187f
C5779 XThR.Tn[4].n13 VGND 0.04765f
C5780 XThR.Tn[4].n14 VGND 0.03348f
C5781 XThR.Tn[4].n16 VGND 0.10743f
C5782 XThR.Tn[4].t39 VGND 0.01713f
C5783 XThR.Tn[4].t31 VGND 0.01876f
C5784 XThR.Tn[4].n17 VGND 0.0458f
C5785 XThR.Tn[4].t58 VGND 0.01707f
C5786 XThR.Tn[4].t27 VGND 0.0187f
C5787 XThR.Tn[4].n18 VGND 0.04765f
C5788 XThR.Tn[4].n19 VGND 0.03348f
C5789 XThR.Tn[4].n21 VGND 0.10743f
C5790 XThR.Tn[4].t55 VGND 0.01713f
C5791 XThR.Tn[4].t48 VGND 0.01876f
C5792 XThR.Tn[4].n22 VGND 0.0458f
C5793 XThR.Tn[4].t70 VGND 0.01707f
C5794 XThR.Tn[4].t45 VGND 0.0187f
C5795 XThR.Tn[4].n23 VGND 0.04765f
C5796 XThR.Tn[4].n24 VGND 0.03348f
C5797 XThR.Tn[4].n26 VGND 0.10743f
C5798 XThR.Tn[4].t17 VGND 0.01713f
C5799 XThR.Tn[4].t13 VGND 0.01876f
C5800 XThR.Tn[4].n27 VGND 0.0458f
C5801 XThR.Tn[4].t41 VGND 0.01707f
C5802 XThR.Tn[4].t71 VGND 0.0187f
C5803 XThR.Tn[4].n28 VGND 0.04765f
C5804 XThR.Tn[4].n29 VGND 0.03348f
C5805 XThR.Tn[4].n31 VGND 0.10743f
C5806 XThR.Tn[4].t57 VGND 0.01713f
C5807 XThR.Tn[4].t49 VGND 0.01876f
C5808 XThR.Tn[4].n32 VGND 0.0458f
C5809 XThR.Tn[4].t73 VGND 0.01707f
C5810 XThR.Tn[4].t46 VGND 0.0187f
C5811 XThR.Tn[4].n33 VGND 0.04765f
C5812 XThR.Tn[4].n34 VGND 0.03348f
C5813 XThR.Tn[4].n36 VGND 0.10743f
C5814 XThR.Tn[4].t33 VGND 0.01713f
C5815 XThR.Tn[4].t66 VGND 0.01876f
C5816 XThR.Tn[4].n37 VGND 0.0458f
C5817 XThR.Tn[4].t52 VGND 0.01707f
C5818 XThR.Tn[4].t63 VGND 0.0187f
C5819 XThR.Tn[4].n38 VGND 0.04765f
C5820 XThR.Tn[4].n39 VGND 0.03348f
C5821 XThR.Tn[4].n41 VGND 0.10743f
C5822 XThR.Tn[4].t64 VGND 0.01713f
C5823 XThR.Tn[4].t61 VGND 0.01876f
C5824 XThR.Tn[4].n42 VGND 0.0458f
C5825 XThR.Tn[4].t18 VGND 0.01707f
C5826 XThR.Tn[4].t56 VGND 0.0187f
C5827 XThR.Tn[4].n43 VGND 0.04765f
C5828 XThR.Tn[4].n44 VGND 0.03348f
C5829 XThR.Tn[4].n46 VGND 0.10743f
C5830 XThR.Tn[4].t68 VGND 0.01713f
C5831 XThR.Tn[4].t12 VGND 0.01876f
C5832 XThR.Tn[4].n47 VGND 0.0458f
C5833 XThR.Tn[4].t25 VGND 0.01707f
C5834 XThR.Tn[4].t69 VGND 0.0187f
C5835 XThR.Tn[4].n48 VGND 0.04765f
C5836 XThR.Tn[4].n49 VGND 0.03348f
C5837 XThR.Tn[4].n51 VGND 0.10743f
C5838 XThR.Tn[4].t22 VGND 0.01713f
C5839 XThR.Tn[4].t32 VGND 0.01876f
C5840 XThR.Tn[4].n52 VGND 0.0458f
C5841 XThR.Tn[4].t43 VGND 0.01707f
C5842 XThR.Tn[4].t29 VGND 0.0187f
C5843 XThR.Tn[4].n53 VGND 0.04765f
C5844 XThR.Tn[4].n54 VGND 0.03348f
C5845 XThR.Tn[4].n56 VGND 0.10743f
C5846 XThR.Tn[4].t15 VGND 0.01713f
C5847 XThR.Tn[4].t51 VGND 0.01876f
C5848 XThR.Tn[4].n57 VGND 0.0458f
C5849 XThR.Tn[4].t36 VGND 0.01707f
C5850 XThR.Tn[4].t47 VGND 0.0187f
C5851 XThR.Tn[4].n58 VGND 0.04765f
C5852 XThR.Tn[4].n59 VGND 0.03348f
C5853 XThR.Tn[4].n61 VGND 0.10743f
C5854 XThR.Tn[4].t35 VGND 0.01713f
C5855 XThR.Tn[4].t26 VGND 0.01876f
C5856 XThR.Tn[4].n62 VGND 0.0458f
C5857 XThR.Tn[4].t53 VGND 0.01707f
C5858 XThR.Tn[4].t21 VGND 0.0187f
C5859 XThR.Tn[4].n63 VGND 0.04765f
C5860 XThR.Tn[4].n64 VGND 0.03348f
C5861 XThR.Tn[4].n66 VGND 0.10743f
C5862 XThR.Tn[4].t67 VGND 0.01713f
C5863 XThR.Tn[4].t62 VGND 0.01876f
C5864 XThR.Tn[4].n67 VGND 0.0458f
C5865 XThR.Tn[4].t23 VGND 0.01707f
C5866 XThR.Tn[4].t59 VGND 0.0187f
C5867 XThR.Tn[4].n68 VGND 0.04765f
C5868 XThR.Tn[4].n69 VGND 0.03348f
C5869 XThR.Tn[4].n71 VGND 0.10743f
C5870 XThR.Tn[4].t20 VGND 0.01713f
C5871 XThR.Tn[4].t14 VGND 0.01876f
C5872 XThR.Tn[4].n72 VGND 0.0458f
C5873 XThR.Tn[4].t42 VGND 0.01707f
C5874 XThR.Tn[4].t72 VGND 0.0187f
C5875 XThR.Tn[4].n73 VGND 0.04765f
C5876 XThR.Tn[4].n74 VGND 0.03348f
C5877 XThR.Tn[4].n76 VGND 0.10743f
C5878 XThR.Tn[4].t40 VGND 0.01713f
C5879 XThR.Tn[4].t34 VGND 0.01876f
C5880 XThR.Tn[4].n77 VGND 0.0458f
C5881 XThR.Tn[4].t60 VGND 0.01707f
C5882 XThR.Tn[4].t30 VGND 0.0187f
C5883 XThR.Tn[4].n78 VGND 0.04765f
C5884 XThR.Tn[4].n79 VGND 0.03348f
C5885 XThR.Tn[4].n81 VGND 0.10743f
C5886 XThR.Tn[4].t16 VGND 0.01713f
C5887 XThR.Tn[4].t28 VGND 0.01876f
C5888 XThR.Tn[4].n82 VGND 0.0458f
C5889 XThR.Tn[4].t37 VGND 0.01707f
C5890 XThR.Tn[4].t24 VGND 0.0187f
C5891 XThR.Tn[4].n83 VGND 0.04765f
C5892 XThR.Tn[4].n84 VGND 0.03348f
C5893 XThR.Tn[4].n86 VGND 0.10743f
C5894 XThR.Tn[4].n87 VGND 0.09763f
C5895 XThR.Tn[4].n88 VGND 0.18445f
C5896 XThC.Tn[7].t4 VGND 0.02413f
C5897 XThC.Tn[7].t7 VGND 0.02413f
C5898 XThC.Tn[7].n0 VGND 0.05198f
C5899 XThC.Tn[7].t6 VGND 0.02413f
C5900 XThC.Tn[7].t5 VGND 0.02413f
C5901 XThC.Tn[7].n1 VGND 0.07891f
C5902 XThC.Tn[7].n2 VGND 0.23202f
C5903 XThC.Tn[7].t8 VGND 0.01913f
C5904 XThC.Tn[7].t11 VGND 0.02089f
C5905 XThC.Tn[7].n3 VGND 0.04666f
C5906 XThC.Tn[7].n4 VGND 0.02666f
C5907 XThC.Tn[7].n5 VGND 0.03243f
C5908 XThC.Tn[7].t25 VGND 0.01913f
C5909 XThC.Tn[7].t30 VGND 0.02089f
C5910 XThC.Tn[7].n6 VGND 0.04666f
C5911 XThC.Tn[7].n7 VGND 0.02666f
C5912 XThC.Tn[7].n8 VGND 0.15407f
C5913 XThC.Tn[7].t27 VGND 0.01913f
C5914 XThC.Tn[7].t34 VGND 0.02089f
C5915 XThC.Tn[7].n9 VGND 0.04666f
C5916 XThC.Tn[7].n10 VGND 0.02666f
C5917 XThC.Tn[7].n11 VGND 0.15407f
C5918 XThC.Tn[7].t29 VGND 0.01913f
C5919 XThC.Tn[7].t35 VGND 0.02089f
C5920 XThC.Tn[7].n12 VGND 0.04666f
C5921 XThC.Tn[7].n13 VGND 0.02666f
C5922 XThC.Tn[7].n14 VGND 0.15407f
C5923 XThC.Tn[7].t18 VGND 0.01913f
C5924 XThC.Tn[7].t22 VGND 0.02089f
C5925 XThC.Tn[7].n15 VGND 0.04666f
C5926 XThC.Tn[7].n16 VGND 0.02666f
C5927 XThC.Tn[7].n17 VGND 0.15407f
C5928 XThC.Tn[7].t20 VGND 0.01913f
C5929 XThC.Tn[7].t23 VGND 0.02089f
C5930 XThC.Tn[7].n18 VGND 0.04666f
C5931 XThC.Tn[7].n19 VGND 0.02666f
C5932 XThC.Tn[7].n20 VGND 0.15407f
C5933 XThC.Tn[7].t33 VGND 0.01913f
C5934 XThC.Tn[7].t39 VGND 0.02089f
C5935 XThC.Tn[7].n21 VGND 0.04666f
C5936 XThC.Tn[7].n22 VGND 0.02666f
C5937 XThC.Tn[7].n23 VGND 0.15407f
C5938 XThC.Tn[7].t10 VGND 0.01913f
C5939 XThC.Tn[7].t14 VGND 0.02089f
C5940 XThC.Tn[7].n24 VGND 0.04666f
C5941 XThC.Tn[7].n25 VGND 0.02666f
C5942 XThC.Tn[7].n26 VGND 0.15407f
C5943 XThC.Tn[7].t12 VGND 0.01913f
C5944 XThC.Tn[7].t16 VGND 0.02089f
C5945 XThC.Tn[7].n27 VGND 0.04666f
C5946 XThC.Tn[7].n28 VGND 0.02666f
C5947 XThC.Tn[7].n29 VGND 0.15407f
C5948 XThC.Tn[7].t31 VGND 0.01913f
C5949 XThC.Tn[7].t36 VGND 0.02089f
C5950 XThC.Tn[7].n30 VGND 0.04666f
C5951 XThC.Tn[7].n31 VGND 0.02666f
C5952 XThC.Tn[7].n32 VGND 0.15407f
C5953 XThC.Tn[7].t32 VGND 0.01913f
C5954 XThC.Tn[7].t38 VGND 0.02089f
C5955 XThC.Tn[7].n33 VGND 0.04666f
C5956 XThC.Tn[7].n34 VGND 0.02666f
C5957 XThC.Tn[7].n35 VGND 0.15407f
C5958 XThC.Tn[7].t13 VGND 0.01913f
C5959 XThC.Tn[7].t17 VGND 0.02089f
C5960 XThC.Tn[7].n36 VGND 0.04666f
C5961 XThC.Tn[7].n37 VGND 0.02666f
C5962 XThC.Tn[7].n38 VGND 0.15407f
C5963 XThC.Tn[7].t21 VGND 0.01913f
C5964 XThC.Tn[7].t26 VGND 0.02089f
C5965 XThC.Tn[7].n39 VGND 0.04666f
C5966 XThC.Tn[7].n40 VGND 0.02666f
C5967 XThC.Tn[7].n41 VGND 0.15407f
C5968 XThC.Tn[7].t24 VGND 0.01913f
C5969 XThC.Tn[7].t28 VGND 0.02089f
C5970 XThC.Tn[7].n42 VGND 0.04666f
C5971 XThC.Tn[7].n43 VGND 0.02666f
C5972 XThC.Tn[7].n44 VGND 0.15407f
C5973 XThC.Tn[7].t37 VGND 0.01913f
C5974 XThC.Tn[7].t9 VGND 0.02089f
C5975 XThC.Tn[7].n45 VGND 0.04666f
C5976 XThC.Tn[7].n46 VGND 0.02666f
C5977 XThC.Tn[7].n47 VGND 0.15407f
C5978 XThC.Tn[7].t15 VGND 0.01913f
C5979 XThC.Tn[7].t19 VGND 0.02089f
C5980 XThC.Tn[7].n48 VGND 0.04666f
C5981 XThC.Tn[7].n49 VGND 0.02666f
C5982 XThC.Tn[7].n50 VGND 0.15407f
C5983 XThC.Tn[7].n51 VGND 0.97494f
C5984 XThC.Tn[7].n52 VGND 0.06268f
C5985 XThC.Tn[7].t2 VGND 0.01569f
C5986 XThC.Tn[7].t1 VGND 0.01569f
C5987 XThC.Tn[7].n53 VGND 0.04842f
C5988 XThC.Tn[7].t0 VGND 0.01569f
C5989 XThC.Tn[7].t3 VGND 0.01569f
C5990 XThC.Tn[7].n54 VGND 0.03465f
C5991 XThC.Tn[7].n55 VGND 0.17137f
C5992 XThC.Tn[7].n56 VGND 0.02887f
C5993 XThR.Tn[1].t8 VGND 0.02151f
C5994 XThR.Tn[1].t9 VGND 0.02151f
C5995 XThR.Tn[1].n0 VGND 0.04341f
C5996 XThR.Tn[1].t11 VGND 0.02151f
C5997 XThR.Tn[1].t10 VGND 0.02151f
C5998 XThR.Tn[1].n1 VGND 0.05079f
C5999 XThR.Tn[1].n2 VGND 0.14218f
C6000 XThR.Tn[1].t7 VGND 0.01398f
C6001 XThR.Tn[1].t4 VGND 0.01398f
C6002 XThR.Tn[1].n3 VGND 0.03183f
C6003 XThR.Tn[1].t6 VGND 0.01398f
C6004 XThR.Tn[1].t5 VGND 0.01398f
C6005 XThR.Tn[1].n4 VGND 0.03183f
C6006 XThR.Tn[1].t2 VGND 0.01398f
C6007 XThR.Tn[1].t1 VGND 0.01398f
C6008 XThR.Tn[1].n5 VGND 0.03183f
C6009 XThR.Tn[1].t3 VGND 0.01398f
C6010 XThR.Tn[1].t0 VGND 0.01398f
C6011 XThR.Tn[1].n6 VGND 0.05304f
C6012 XThR.Tn[1].n7 VGND 0.15159f
C6013 XThR.Tn[1].n8 VGND 0.09371f
C6014 XThR.Tn[1].n9 VGND 0.10576f
C6015 XThR.Tn[1].t24 VGND 0.01681f
C6016 XThR.Tn[1].t18 VGND 0.0184f
C6017 XThR.Tn[1].n10 VGND 0.04494f
C6018 XThR.Tn[1].n11 VGND 0.06984f
C6019 XThR.Tn[1].t44 VGND 0.01681f
C6020 XThR.Tn[1].t34 VGND 0.0184f
C6021 XThR.Tn[1].n12 VGND 0.04494f
C6022 XThR.Tn[1].t61 VGND 0.01675f
C6023 XThR.Tn[1].t30 VGND 0.01834f
C6024 XThR.Tn[1].n13 VGND 0.04676f
C6025 XThR.Tn[1].n14 VGND 0.03285f
C6026 XThR.Tn[1].n16 VGND 0.10542f
C6027 XThR.Tn[1].t19 VGND 0.01681f
C6028 XThR.Tn[1].t73 VGND 0.0184f
C6029 XThR.Tn[1].n17 VGND 0.04494f
C6030 XThR.Tn[1].t38 VGND 0.01675f
C6031 XThR.Tn[1].t69 VGND 0.01834f
C6032 XThR.Tn[1].n18 VGND 0.04676f
C6033 XThR.Tn[1].n19 VGND 0.03285f
C6034 XThR.Tn[1].n21 VGND 0.10542f
C6035 XThR.Tn[1].t35 VGND 0.01681f
C6036 XThR.Tn[1].t28 VGND 0.0184f
C6037 XThR.Tn[1].n22 VGND 0.04494f
C6038 XThR.Tn[1].t50 VGND 0.01675f
C6039 XThR.Tn[1].t25 VGND 0.01834f
C6040 XThR.Tn[1].n23 VGND 0.04676f
C6041 XThR.Tn[1].n24 VGND 0.03285f
C6042 XThR.Tn[1].n26 VGND 0.10542f
C6043 XThR.Tn[1].t59 VGND 0.01681f
C6044 XThR.Tn[1].t55 VGND 0.0184f
C6045 XThR.Tn[1].n27 VGND 0.04494f
C6046 XThR.Tn[1].t21 VGND 0.01675f
C6047 XThR.Tn[1].t51 VGND 0.01834f
C6048 XThR.Tn[1].n28 VGND 0.04676f
C6049 XThR.Tn[1].n29 VGND 0.03285f
C6050 XThR.Tn[1].n31 VGND 0.10542f
C6051 XThR.Tn[1].t37 VGND 0.01681f
C6052 XThR.Tn[1].t29 VGND 0.0184f
C6053 XThR.Tn[1].n32 VGND 0.04494f
C6054 XThR.Tn[1].t53 VGND 0.01675f
C6055 XThR.Tn[1].t26 VGND 0.01834f
C6056 XThR.Tn[1].n33 VGND 0.04676f
C6057 XThR.Tn[1].n34 VGND 0.03285f
C6058 XThR.Tn[1].n36 VGND 0.10542f
C6059 XThR.Tn[1].t13 VGND 0.01681f
C6060 XThR.Tn[1].t46 VGND 0.0184f
C6061 XThR.Tn[1].n37 VGND 0.04494f
C6062 XThR.Tn[1].t32 VGND 0.01675f
C6063 XThR.Tn[1].t43 VGND 0.01834f
C6064 XThR.Tn[1].n38 VGND 0.04676f
C6065 XThR.Tn[1].n39 VGND 0.03285f
C6066 XThR.Tn[1].n41 VGND 0.10542f
C6067 XThR.Tn[1].t45 VGND 0.01681f
C6068 XThR.Tn[1].t41 VGND 0.0184f
C6069 XThR.Tn[1].n42 VGND 0.04494f
C6070 XThR.Tn[1].t60 VGND 0.01675f
C6071 XThR.Tn[1].t36 VGND 0.01834f
C6072 XThR.Tn[1].n43 VGND 0.04676f
C6073 XThR.Tn[1].n44 VGND 0.03285f
C6074 XThR.Tn[1].n46 VGND 0.10542f
C6075 XThR.Tn[1].t48 VGND 0.01681f
C6076 XThR.Tn[1].t54 VGND 0.0184f
C6077 XThR.Tn[1].n47 VGND 0.04494f
C6078 XThR.Tn[1].t67 VGND 0.01675f
C6079 XThR.Tn[1].t49 VGND 0.01834f
C6080 XThR.Tn[1].n48 VGND 0.04676f
C6081 XThR.Tn[1].n49 VGND 0.03285f
C6082 XThR.Tn[1].n51 VGND 0.10542f
C6083 XThR.Tn[1].t64 VGND 0.01681f
C6084 XThR.Tn[1].t12 VGND 0.0184f
C6085 XThR.Tn[1].n52 VGND 0.04494f
C6086 XThR.Tn[1].t23 VGND 0.01675f
C6087 XThR.Tn[1].t71 VGND 0.01834f
C6088 XThR.Tn[1].n53 VGND 0.04676f
C6089 XThR.Tn[1].n54 VGND 0.03285f
C6090 XThR.Tn[1].n56 VGND 0.10542f
C6091 XThR.Tn[1].t57 VGND 0.01681f
C6092 XThR.Tn[1].t31 VGND 0.0184f
C6093 XThR.Tn[1].n57 VGND 0.04494f
C6094 XThR.Tn[1].t16 VGND 0.01675f
C6095 XThR.Tn[1].t27 VGND 0.01834f
C6096 XThR.Tn[1].n58 VGND 0.04676f
C6097 XThR.Tn[1].n59 VGND 0.03285f
C6098 XThR.Tn[1].n61 VGND 0.10542f
C6099 XThR.Tn[1].t15 VGND 0.01681f
C6100 XThR.Tn[1].t68 VGND 0.0184f
C6101 XThR.Tn[1].n62 VGND 0.04494f
C6102 XThR.Tn[1].t33 VGND 0.01675f
C6103 XThR.Tn[1].t63 VGND 0.01834f
C6104 XThR.Tn[1].n63 VGND 0.04676f
C6105 XThR.Tn[1].n64 VGND 0.03285f
C6106 XThR.Tn[1].n66 VGND 0.10542f
C6107 XThR.Tn[1].t47 VGND 0.01681f
C6108 XThR.Tn[1].t42 VGND 0.0184f
C6109 XThR.Tn[1].n67 VGND 0.04494f
C6110 XThR.Tn[1].t65 VGND 0.01675f
C6111 XThR.Tn[1].t39 VGND 0.01834f
C6112 XThR.Tn[1].n68 VGND 0.04676f
C6113 XThR.Tn[1].n69 VGND 0.03285f
C6114 XThR.Tn[1].n71 VGND 0.10542f
C6115 XThR.Tn[1].t62 VGND 0.01681f
C6116 XThR.Tn[1].t56 VGND 0.0184f
C6117 XThR.Tn[1].n72 VGND 0.04494f
C6118 XThR.Tn[1].t22 VGND 0.01675f
C6119 XThR.Tn[1].t52 VGND 0.01834f
C6120 XThR.Tn[1].n73 VGND 0.04676f
C6121 XThR.Tn[1].n74 VGND 0.03285f
C6122 XThR.Tn[1].n76 VGND 0.10542f
C6123 XThR.Tn[1].t20 VGND 0.01681f
C6124 XThR.Tn[1].t14 VGND 0.0184f
C6125 XThR.Tn[1].n77 VGND 0.04494f
C6126 XThR.Tn[1].t40 VGND 0.01675f
C6127 XThR.Tn[1].t72 VGND 0.01834f
C6128 XThR.Tn[1].n78 VGND 0.04676f
C6129 XThR.Tn[1].n79 VGND 0.03285f
C6130 XThR.Tn[1].n81 VGND 0.10542f
C6131 XThR.Tn[1].t58 VGND 0.01681f
C6132 XThR.Tn[1].t70 VGND 0.0184f
C6133 XThR.Tn[1].n82 VGND 0.04494f
C6134 XThR.Tn[1].t17 VGND 0.01675f
C6135 XThR.Tn[1].t66 VGND 0.01834f
C6136 XThR.Tn[1].n83 VGND 0.04676f
C6137 XThR.Tn[1].n84 VGND 0.03285f
C6138 XThR.Tn[1].n86 VGND 0.10542f
C6139 XThR.Tn[1].n87 VGND 0.0958f
C6140 XThR.Tn[1].n88 VGND 0.27576f
C6141 XThR.Tn[1].n89 VGND 0.045f
C6142 XThC.Tn[8].t5 VGND 0.01696f
C6143 XThC.Tn[8].t4 VGND 0.01696f
C6144 XThC.Tn[8].n0 VGND 0.04229f
C6145 XThC.Tn[8].t7 VGND 0.01696f
C6146 XThC.Tn[8].t6 VGND 0.01696f
C6147 XThC.Tn[8].n1 VGND 0.03391f
C6148 XThC.Tn[8].n2 VGND 0.08531f
C6149 XThC.Tn[8].t43 VGND 0.02068f
C6150 XThC.Tn[8].t41 VGND 0.02258f
C6151 XThC.Tn[8].n3 VGND 0.05043f
C6152 XThC.Tn[8].n4 VGND 0.02882f
C6153 XThC.Tn[8].n5 VGND 0.03505f
C6154 XThC.Tn[8].t29 VGND 0.02068f
C6155 XThC.Tn[8].t26 VGND 0.02258f
C6156 XThC.Tn[8].n6 VGND 0.05043f
C6157 XThC.Tn[8].n7 VGND 0.02882f
C6158 XThC.Tn[8].n8 VGND 0.16652f
C6159 XThC.Tn[8].t34 VGND 0.02068f
C6160 XThC.Tn[8].t28 VGND 0.02258f
C6161 XThC.Tn[8].n9 VGND 0.05043f
C6162 XThC.Tn[8].n10 VGND 0.02882f
C6163 XThC.Tn[8].n11 VGND 0.16652f
C6164 XThC.Tn[8].t35 VGND 0.02068f
C6165 XThC.Tn[8].t30 VGND 0.02258f
C6166 XThC.Tn[8].n12 VGND 0.05043f
C6167 XThC.Tn[8].n13 VGND 0.02882f
C6168 XThC.Tn[8].n14 VGND 0.16652f
C6169 XThC.Tn[8].t22 VGND 0.02068f
C6170 XThC.Tn[8].t19 VGND 0.02258f
C6171 XThC.Tn[8].n15 VGND 0.05043f
C6172 XThC.Tn[8].n16 VGND 0.02882f
C6173 XThC.Tn[8].n17 VGND 0.16652f
C6174 XThC.Tn[8].t23 VGND 0.02068f
C6175 XThC.Tn[8].t20 VGND 0.02258f
C6176 XThC.Tn[8].n18 VGND 0.05043f
C6177 XThC.Tn[8].n19 VGND 0.02882f
C6178 XThC.Tn[8].n20 VGND 0.16652f
C6179 XThC.Tn[8].t39 VGND 0.02068f
C6180 XThC.Tn[8].t33 VGND 0.02258f
C6181 XThC.Tn[8].n21 VGND 0.05043f
C6182 XThC.Tn[8].n22 VGND 0.02882f
C6183 XThC.Tn[8].n23 VGND 0.16652f
C6184 XThC.Tn[8].t14 VGND 0.02068f
C6185 XThC.Tn[8].t42 VGND 0.02258f
C6186 XThC.Tn[8].n24 VGND 0.05043f
C6187 XThC.Tn[8].n25 VGND 0.02882f
C6188 XThC.Tn[8].n26 VGND 0.16652f
C6189 XThC.Tn[8].t16 VGND 0.02068f
C6190 XThC.Tn[8].t12 VGND 0.02258f
C6191 XThC.Tn[8].n27 VGND 0.05043f
C6192 XThC.Tn[8].n28 VGND 0.02882f
C6193 XThC.Tn[8].n29 VGND 0.16652f
C6194 XThC.Tn[8].t36 VGND 0.02068f
C6195 XThC.Tn[8].t31 VGND 0.02258f
C6196 XThC.Tn[8].n30 VGND 0.05043f
C6197 XThC.Tn[8].n31 VGND 0.02882f
C6198 XThC.Tn[8].n32 VGND 0.16652f
C6199 XThC.Tn[8].t38 VGND 0.02068f
C6200 XThC.Tn[8].t32 VGND 0.02258f
C6201 XThC.Tn[8].n33 VGND 0.05043f
C6202 XThC.Tn[8].n34 VGND 0.02882f
C6203 XThC.Tn[8].n35 VGND 0.16652f
C6204 XThC.Tn[8].t17 VGND 0.02068f
C6205 XThC.Tn[8].t13 VGND 0.02258f
C6206 XThC.Tn[8].n36 VGND 0.05043f
C6207 XThC.Tn[8].n37 VGND 0.02882f
C6208 XThC.Tn[8].n38 VGND 0.16652f
C6209 XThC.Tn[8].t25 VGND 0.02068f
C6210 XThC.Tn[8].t21 VGND 0.02258f
C6211 XThC.Tn[8].n39 VGND 0.05043f
C6212 XThC.Tn[8].n40 VGND 0.02882f
C6213 XThC.Tn[8].n41 VGND 0.16652f
C6214 XThC.Tn[8].t27 VGND 0.02068f
C6215 XThC.Tn[8].t24 VGND 0.02258f
C6216 XThC.Tn[8].n42 VGND 0.05043f
C6217 XThC.Tn[8].n43 VGND 0.02882f
C6218 XThC.Tn[8].n44 VGND 0.16652f
C6219 XThC.Tn[8].t40 VGND 0.02068f
C6220 XThC.Tn[8].t37 VGND 0.02258f
C6221 XThC.Tn[8].n45 VGND 0.05043f
C6222 XThC.Tn[8].n46 VGND 0.02882f
C6223 XThC.Tn[8].n47 VGND 0.16652f
C6224 XThC.Tn[8].t18 VGND 0.02068f
C6225 XThC.Tn[8].t15 VGND 0.02258f
C6226 XThC.Tn[8].n48 VGND 0.05043f
C6227 XThC.Tn[8].n49 VGND 0.02882f
C6228 XThC.Tn[8].n50 VGND 0.16652f
C6229 XThC.Tn[8].n51 VGND 0.07701f
C6230 XThC.Tn[8].n52 VGND 0.72901f
C6231 XThC.Tn[8].n53 VGND 0.05851f
C6232 XThC.Tn[8].t9 VGND 0.02609f
C6233 XThC.Tn[8].t10 VGND 0.02609f
C6234 XThC.Tn[8].n54 VGND 0.05636f
C6235 XThC.Tn[8].t8 VGND 0.02609f
C6236 XThC.Tn[8].t11 VGND 0.02609f
C6237 XThC.Tn[8].n55 VGND 0.08578f
C6238 XThC.Tn[8].n56 VGND 0.23835f
C6239 XThC.Tn[8].n57 VGND 0.03748f
C6240 XThC.Tn[8].t2 VGND 0.02609f
C6241 XThC.Tn[8].t1 VGND 0.02609f
C6242 XThC.Tn[8].n58 VGND 0.05799f
C6243 XThC.Tn[8].t0 VGND 0.02609f
C6244 XThC.Tn[8].t3 VGND 0.02609f
C6245 XThC.Tn[8].n59 VGND 0.0792f
C6246 XThC.Tn[8].n60 VGND 0.25808f
C6247 XThC.XTB1.Y.t1 VGND 0.03224f
C6248 XThC.XTB1.Y.n0 VGND 0.02084f
C6249 XThC.XTB1.Y.n1 VGND 0.02659f
C6250 XThC.XTB1.Y.t2 VGND 0.01618f
C6251 XThC.XTB1.Y.t0 VGND 0.01618f
C6252 XThC.XTB1.Y.n2 VGND 0.03473f
C6253 XThC.XTB1.Y.t17 VGND 0.02517f
C6254 XThC.XTB1.Y.t5 VGND 0.01483f
C6255 XThC.XTB1.Y.n3 VGND 0.02997f
C6256 XThC.XTB1.Y.t6 VGND 0.02517f
C6257 XThC.XTB1.Y.t12 VGND 0.01483f
C6258 XThC.XTB1.Y.n4 VGND 0.01542f
C6259 XThC.XTB1.Y.t8 VGND 0.02517f
C6260 XThC.XTB1.Y.t13 VGND 0.01483f
C6261 XThC.XTB1.Y.n5 VGND 0.03313f
C6262 XThC.XTB1.Y.t11 VGND 0.02517f
C6263 XThC.XTB1.Y.t16 VGND 0.01483f
C6264 XThC.XTB1.Y.n6 VGND 0.03076f
C6265 XThC.XTB1.Y.n7 VGND 0.01871f
C6266 XThC.XTB1.Y.n8 VGND 0.03098f
C6267 XThC.XTB1.Y.n9 VGND 0.01198f
C6268 XThC.XTB1.Y.n10 VGND 0.01463f
C6269 XThC.XTB1.Y.n11 VGND 0.03313f
C6270 XThC.XTB1.Y.n12 VGND 0.01661f
C6271 XThC.XTB1.Y.n13 VGND 0.02824f
C6272 XThC.XTB1.Y.t18 VGND 0.02517f
C6273 XThC.XTB1.Y.t9 VGND 0.01483f
C6274 XThC.XTB1.Y.n14 VGND 0.03392f
C6275 XThC.XTB1.Y.t7 VGND 0.02517f
C6276 XThC.XTB1.Y.t15 VGND 0.01483f
C6277 XThC.XTB1.Y.t14 VGND 0.02517f
C6278 XThC.XTB1.Y.t3 VGND 0.01483f
C6279 XThC.XTB1.Y.t10 VGND 0.02517f
C6280 XThC.XTB1.Y.t4 VGND 0.01483f
C6281 XThC.XTB1.Y.n15 VGND 0.04223f
C6282 XThC.XTB1.Y.n16 VGND 0.0446f
C6283 XThC.XTB1.Y.n17 VGND 0.01719f
C6284 XThC.XTB1.Y.n18 VGND 0.0363f
C6285 XThC.XTB1.Y.n19 VGND 0.01661f
C6286 XThC.XTB1.Y.n20 VGND 0.01378f
C6287 XThC.XTB1.Y.n21 VGND 0.77148f
C6288 XThC.XTB1.Y.n22 VGND 0.07634f
C6289 XThC.Tn[14].t4 VGND 0.01604f
C6290 XThC.Tn[14].t6 VGND 0.01604f
C6291 XThC.Tn[14].n0 VGND 0.04002f
C6292 XThC.Tn[14].t5 VGND 0.01604f
C6293 XThC.Tn[14].t7 VGND 0.01604f
C6294 XThC.Tn[14].n1 VGND 0.03209f
C6295 XThC.Tn[14].n2 VGND 0.08072f
C6296 XThC.Tn[14].t43 VGND 0.01956f
C6297 XThC.Tn[14].t38 VGND 0.02137f
C6298 XThC.Tn[14].n3 VGND 0.04772f
C6299 XThC.Tn[14].n4 VGND 0.02727f
C6300 XThC.Tn[14].n5 VGND 0.03317f
C6301 XThC.Tn[14].t29 VGND 0.01956f
C6302 XThC.Tn[14].t22 VGND 0.02137f
C6303 XThC.Tn[14].n6 VGND 0.04772f
C6304 XThC.Tn[14].n7 VGND 0.02727f
C6305 XThC.Tn[14].n8 VGND 0.15757f
C6306 XThC.Tn[14].t32 VGND 0.01956f
C6307 XThC.Tn[14].t25 VGND 0.02137f
C6308 XThC.Tn[14].n9 VGND 0.04772f
C6309 XThC.Tn[14].n10 VGND 0.02727f
C6310 XThC.Tn[14].n11 VGND 0.15757f
C6311 XThC.Tn[14].t34 VGND 0.01956f
C6312 XThC.Tn[14].t26 VGND 0.02137f
C6313 XThC.Tn[14].n12 VGND 0.04772f
C6314 XThC.Tn[14].n13 VGND 0.02727f
C6315 XThC.Tn[14].n14 VGND 0.15757f
C6316 XThC.Tn[14].t20 VGND 0.01956f
C6317 XThC.Tn[14].t14 VGND 0.02137f
C6318 XThC.Tn[14].n15 VGND 0.04772f
C6319 XThC.Tn[14].n16 VGND 0.02727f
C6320 XThC.Tn[14].n17 VGND 0.15757f
C6321 XThC.Tn[14].t23 VGND 0.01956f
C6322 XThC.Tn[14].t17 VGND 0.02137f
C6323 XThC.Tn[14].n18 VGND 0.04772f
C6324 XThC.Tn[14].n19 VGND 0.02727f
C6325 XThC.Tn[14].n20 VGND 0.15757f
C6326 XThC.Tn[14].t37 VGND 0.01956f
C6327 XThC.Tn[14].t31 VGND 0.02137f
C6328 XThC.Tn[14].n21 VGND 0.04772f
C6329 XThC.Tn[14].n22 VGND 0.02727f
C6330 XThC.Tn[14].n23 VGND 0.15757f
C6331 XThC.Tn[14].t13 VGND 0.01956f
C6332 XThC.Tn[14].t39 VGND 0.02137f
C6333 XThC.Tn[14].n24 VGND 0.04772f
C6334 XThC.Tn[14].n25 VGND 0.02727f
C6335 XThC.Tn[14].n26 VGND 0.15757f
C6336 XThC.Tn[14].t15 VGND 0.01956f
C6337 XThC.Tn[14].t41 VGND 0.02137f
C6338 XThC.Tn[14].n27 VGND 0.04772f
C6339 XThC.Tn[14].n28 VGND 0.02727f
C6340 XThC.Tn[14].n29 VGND 0.15757f
C6341 XThC.Tn[14].t35 VGND 0.01956f
C6342 XThC.Tn[14].t27 VGND 0.02137f
C6343 XThC.Tn[14].n30 VGND 0.04772f
C6344 XThC.Tn[14].n31 VGND 0.02727f
C6345 XThC.Tn[14].n32 VGND 0.15757f
C6346 XThC.Tn[14].t36 VGND 0.01956f
C6347 XThC.Tn[14].t30 VGND 0.02137f
C6348 XThC.Tn[14].n33 VGND 0.04772f
C6349 XThC.Tn[14].n34 VGND 0.02727f
C6350 XThC.Tn[14].n35 VGND 0.15757f
C6351 XThC.Tn[14].t16 VGND 0.01956f
C6352 XThC.Tn[14].t42 VGND 0.02137f
C6353 XThC.Tn[14].n36 VGND 0.04772f
C6354 XThC.Tn[14].n37 VGND 0.02727f
C6355 XThC.Tn[14].n38 VGND 0.15757f
C6356 XThC.Tn[14].t24 VGND 0.01956f
C6357 XThC.Tn[14].t19 VGND 0.02137f
C6358 XThC.Tn[14].n39 VGND 0.04772f
C6359 XThC.Tn[14].n40 VGND 0.02727f
C6360 XThC.Tn[14].n41 VGND 0.15757f
C6361 XThC.Tn[14].t28 VGND 0.01956f
C6362 XThC.Tn[14].t21 VGND 0.02137f
C6363 XThC.Tn[14].n42 VGND 0.04772f
C6364 XThC.Tn[14].n43 VGND 0.02727f
C6365 XThC.Tn[14].n44 VGND 0.15757f
C6366 XThC.Tn[14].t40 VGND 0.01956f
C6367 XThC.Tn[14].t33 VGND 0.02137f
C6368 XThC.Tn[14].n45 VGND 0.04772f
C6369 XThC.Tn[14].n46 VGND 0.02727f
C6370 XThC.Tn[14].n47 VGND 0.15757f
C6371 XThC.Tn[14].t18 VGND 0.01956f
C6372 XThC.Tn[14].t12 VGND 0.02137f
C6373 XThC.Tn[14].n48 VGND 0.04772f
C6374 XThC.Tn[14].n49 VGND 0.02727f
C6375 XThC.Tn[14].n50 VGND 0.15757f
C6376 XThC.Tn[14].n51 VGND 0.94072f
C6377 XThC.Tn[14].n52 VGND 0.06007f
C6378 XThC.Tn[14].t8 VGND 0.02468f
C6379 XThC.Tn[14].t9 VGND 0.02468f
C6380 XThC.Tn[14].n53 VGND 0.05333f
C6381 XThC.Tn[14].t11 VGND 0.02468f
C6382 XThC.Tn[14].t10 VGND 0.02468f
C6383 XThC.Tn[14].n54 VGND 0.08117f
C6384 XThC.Tn[14].n55 VGND 0.22554f
C6385 XThC.Tn[14].n56 VGND 0.03546f
C6386 XThC.Tn[14].t1 VGND 0.02468f
C6387 XThC.Tn[14].t0 VGND 0.02468f
C6388 XThC.Tn[14].n57 VGND 0.05487f
C6389 XThC.Tn[14].t3 VGND 0.02468f
C6390 XThC.Tn[14].t2 VGND 0.02468f
C6391 XThC.Tn[14].n58 VGND 0.07495f
C6392 XThC.Tn[14].n59 VGND 0.24421f
C6393 XThR.Tn[10].t10 VGND 0.02288f
C6394 XThR.Tn[10].t8 VGND 0.02288f
C6395 XThR.Tn[10].n0 VGND 0.06946f
C6396 XThR.Tn[10].t11 VGND 0.02288f
C6397 XThR.Tn[10].t9 VGND 0.02288f
C6398 XThR.Tn[10].n1 VGND 0.05085f
C6399 XThR.Tn[10].n2 VGND 0.23122f
C6400 XThR.Tn[10].t6 VGND 0.02288f
C6401 XThR.Tn[10].t4 VGND 0.02288f
C6402 XThR.Tn[10].n3 VGND 0.04942f
C6403 XThR.Tn[10].t7 VGND 0.02288f
C6404 XThR.Tn[10].t5 VGND 0.02288f
C6405 XThR.Tn[10].n4 VGND 0.07522f
C6406 XThR.Tn[10].n5 VGND 0.20887f
C6407 XThR.Tn[10].n6 VGND 0.01029f
C6408 XThR.Tn[10].t54 VGND 0.01788f
C6409 XThR.Tn[10].t47 VGND 0.01958f
C6410 XThR.Tn[10].n7 VGND 0.0478f
C6411 XThR.Tn[10].n8 VGND 0.07429f
C6412 XThR.Tn[10].t13 VGND 0.01788f
C6413 XThR.Tn[10].t63 VGND 0.01958f
C6414 XThR.Tn[10].n9 VGND 0.0478f
C6415 XThR.Tn[10].t50 VGND 0.01782f
C6416 XThR.Tn[10].t60 VGND 0.01951f
C6417 XThR.Tn[10].n10 VGND 0.04974f
C6418 XThR.Tn[10].n11 VGND 0.03494f
C6419 XThR.Tn[10].n13 VGND 0.11213f
C6420 XThR.Tn[10].t48 VGND 0.01788f
C6421 XThR.Tn[10].t41 VGND 0.01958f
C6422 XThR.Tn[10].n14 VGND 0.0478f
C6423 XThR.Tn[10].t23 VGND 0.01782f
C6424 XThR.Tn[10].t36 VGND 0.01951f
C6425 XThR.Tn[10].n15 VGND 0.04974f
C6426 XThR.Tn[10].n16 VGND 0.03494f
C6427 XThR.Tn[10].n18 VGND 0.11213f
C6428 XThR.Tn[10].t65 VGND 0.01788f
C6429 XThR.Tn[10].t58 VGND 0.01958f
C6430 XThR.Tn[10].n19 VGND 0.0478f
C6431 XThR.Tn[10].t40 VGND 0.01782f
C6432 XThR.Tn[10].t55 VGND 0.01951f
C6433 XThR.Tn[10].n20 VGND 0.04974f
C6434 XThR.Tn[10].n21 VGND 0.03494f
C6435 XThR.Tn[10].n23 VGND 0.11213f
C6436 XThR.Tn[10].t30 VGND 0.01788f
C6437 XThR.Tn[10].t26 VGND 0.01958f
C6438 XThR.Tn[10].n24 VGND 0.0478f
C6439 XThR.Tn[10].t70 VGND 0.01782f
C6440 XThR.Tn[10].t21 VGND 0.01951f
C6441 XThR.Tn[10].n25 VGND 0.04974f
C6442 XThR.Tn[10].n26 VGND 0.03494f
C6443 XThR.Tn[10].n28 VGND 0.11213f
C6444 XThR.Tn[10].t67 VGND 0.01788f
C6445 XThR.Tn[10].t59 VGND 0.01958f
C6446 XThR.Tn[10].n29 VGND 0.0478f
C6447 XThR.Tn[10].t42 VGND 0.01782f
C6448 XThR.Tn[10].t56 VGND 0.01951f
C6449 XThR.Tn[10].n30 VGND 0.04974f
C6450 XThR.Tn[10].n31 VGND 0.03494f
C6451 XThR.Tn[10].n33 VGND 0.11213f
C6452 XThR.Tn[10].t44 VGND 0.01788f
C6453 XThR.Tn[10].t15 VGND 0.01958f
C6454 XThR.Tn[10].n34 VGND 0.0478f
C6455 XThR.Tn[10].t18 VGND 0.01782f
C6456 XThR.Tn[10].t12 VGND 0.01951f
C6457 XThR.Tn[10].n35 VGND 0.04974f
C6458 XThR.Tn[10].n36 VGND 0.03494f
C6459 XThR.Tn[10].n38 VGND 0.11213f
C6460 XThR.Tn[10].t14 VGND 0.01788f
C6461 XThR.Tn[10].t69 VGND 0.01958f
C6462 XThR.Tn[10].n39 VGND 0.0478f
C6463 XThR.Tn[10].t51 VGND 0.01782f
C6464 XThR.Tn[10].t66 VGND 0.01951f
C6465 XThR.Tn[10].n40 VGND 0.04974f
C6466 XThR.Tn[10].n41 VGND 0.03494f
C6467 XThR.Tn[10].n43 VGND 0.11213f
C6468 XThR.Tn[10].t17 VGND 0.01788f
C6469 XThR.Tn[10].t24 VGND 0.01958f
C6470 XThR.Tn[10].n44 VGND 0.0478f
C6471 XThR.Tn[10].t53 VGND 0.01782f
C6472 XThR.Tn[10].t20 VGND 0.01951f
C6473 XThR.Tn[10].n45 VGND 0.04974f
C6474 XThR.Tn[10].n46 VGND 0.03494f
C6475 XThR.Tn[10].n48 VGND 0.11213f
C6476 XThR.Tn[10].t33 VGND 0.01788f
C6477 XThR.Tn[10].t43 VGND 0.01958f
C6478 XThR.Tn[10].n49 VGND 0.0478f
C6479 XThR.Tn[10].t73 VGND 0.01782f
C6480 XThR.Tn[10].t38 VGND 0.01951f
C6481 XThR.Tn[10].n50 VGND 0.04974f
C6482 XThR.Tn[10].n51 VGND 0.03494f
C6483 XThR.Tn[10].n53 VGND 0.11213f
C6484 XThR.Tn[10].t28 VGND 0.01788f
C6485 XThR.Tn[10].t61 VGND 0.01958f
C6486 XThR.Tn[10].n54 VGND 0.0478f
C6487 XThR.Tn[10].t62 VGND 0.01782f
C6488 XThR.Tn[10].t57 VGND 0.01951f
C6489 XThR.Tn[10].n55 VGND 0.04974f
C6490 XThR.Tn[10].n56 VGND 0.03494f
C6491 XThR.Tn[10].n58 VGND 0.11213f
C6492 XThR.Tn[10].t46 VGND 0.01788f
C6493 XThR.Tn[10].t35 VGND 0.01958f
C6494 XThR.Tn[10].n59 VGND 0.0478f
C6495 XThR.Tn[10].t19 VGND 0.01782f
C6496 XThR.Tn[10].t32 VGND 0.01951f
C6497 XThR.Tn[10].n60 VGND 0.04974f
C6498 XThR.Tn[10].n61 VGND 0.03494f
C6499 XThR.Tn[10].n63 VGND 0.11213f
C6500 XThR.Tn[10].t16 VGND 0.01788f
C6501 XThR.Tn[10].t72 VGND 0.01958f
C6502 XThR.Tn[10].n64 VGND 0.0478f
C6503 XThR.Tn[10].t52 VGND 0.01782f
C6504 XThR.Tn[10].t68 VGND 0.01951f
C6505 XThR.Tn[10].n65 VGND 0.04974f
C6506 XThR.Tn[10].n66 VGND 0.03494f
C6507 XThR.Tn[10].n68 VGND 0.11213f
C6508 XThR.Tn[10].t31 VGND 0.01788f
C6509 XThR.Tn[10].t27 VGND 0.01958f
C6510 XThR.Tn[10].n69 VGND 0.0478f
C6511 XThR.Tn[10].t71 VGND 0.01782f
C6512 XThR.Tn[10].t22 VGND 0.01951f
C6513 XThR.Tn[10].n70 VGND 0.04974f
C6514 XThR.Tn[10].n71 VGND 0.03494f
C6515 XThR.Tn[10].n73 VGND 0.11213f
C6516 XThR.Tn[10].t49 VGND 0.01788f
C6517 XThR.Tn[10].t45 VGND 0.01958f
C6518 XThR.Tn[10].n74 VGND 0.0478f
C6519 XThR.Tn[10].t25 VGND 0.01782f
C6520 XThR.Tn[10].t39 VGND 0.01951f
C6521 XThR.Tn[10].n75 VGND 0.04974f
C6522 XThR.Tn[10].n76 VGND 0.03494f
C6523 XThR.Tn[10].n78 VGND 0.11213f
C6524 XThR.Tn[10].t29 VGND 0.01788f
C6525 XThR.Tn[10].t37 VGND 0.01958f
C6526 XThR.Tn[10].n79 VGND 0.0478f
C6527 XThR.Tn[10].t64 VGND 0.01782f
C6528 XThR.Tn[10].t34 VGND 0.01951f
C6529 XThR.Tn[10].n80 VGND 0.04974f
C6530 XThR.Tn[10].n81 VGND 0.03494f
C6531 XThR.Tn[10].n83 VGND 0.11213f
C6532 XThR.Tn[10].n84 VGND 0.1019f
C6533 XThR.Tn[10].n85 VGND 0.31372f
C6534 XThR.Tn[10].t0 VGND 0.01487f
C6535 XThR.Tn[10].t2 VGND 0.01487f
C6536 XThR.Tn[10].n86 VGND 0.02974f
C6537 XThR.Tn[10].t1 VGND 0.01487f
C6538 XThR.Tn[10].t3 VGND 0.01487f
C6539 XThR.Tn[10].n87 VGND 0.03708f
C6540 XThR.Tn[10].n88 VGND 0.06857f
C6541 XThC.Tn[3].t5 VGND 0.02303f
C6542 XThC.Tn[3].t4 VGND 0.02303f
C6543 XThC.Tn[3].n0 VGND 0.04649f
C6544 XThC.Tn[3].t7 VGND 0.02303f
C6545 XThC.Tn[3].t6 VGND 0.02303f
C6546 XThC.Tn[3].n1 VGND 0.0544f
C6547 XThC.Tn[3].n2 VGND 0.16316f
C6548 XThC.Tn[3].t1 VGND 0.01497f
C6549 XThC.Tn[3].t0 VGND 0.01497f
C6550 XThC.Tn[3].n3 VGND 0.03409f
C6551 XThC.Tn[3].t11 VGND 0.01497f
C6552 XThC.Tn[3].t10 VGND 0.01497f
C6553 XThC.Tn[3].n4 VGND 0.0568f
C6554 XThC.Tn[3].t9 VGND 0.01497f
C6555 XThC.Tn[3].t8 VGND 0.01497f
C6556 XThC.Tn[3].n5 VGND 0.03409f
C6557 XThC.Tn[3].n6 VGND 0.16235f
C6558 XThC.Tn[3].t3 VGND 0.01497f
C6559 XThC.Tn[3].t2 VGND 0.01497f
C6560 XThC.Tn[3].n7 VGND 0.03409f
C6561 XThC.Tn[3].n8 VGND 0.10036f
C6562 XThC.Tn[3].n9 VGND 0.11327f
C6563 XThC.Tn[3].t12 VGND 0.01826f
C6564 XThC.Tn[3].t42 VGND 0.01994f
C6565 XThC.Tn[3].n10 VGND 0.04453f
C6566 XThC.Tn[3].n11 VGND 0.02545f
C6567 XThC.Tn[3].n12 VGND 0.03095f
C6568 XThC.Tn[3].t30 VGND 0.01826f
C6569 XThC.Tn[3].t27 VGND 0.01994f
C6570 XThC.Tn[3].n13 VGND 0.04453f
C6571 XThC.Tn[3].n14 VGND 0.02545f
C6572 XThC.Tn[3].n15 VGND 0.14703f
C6573 XThC.Tn[3].t35 VGND 0.01826f
C6574 XThC.Tn[3].t29 VGND 0.01994f
C6575 XThC.Tn[3].n16 VGND 0.04453f
C6576 XThC.Tn[3].n17 VGND 0.02545f
C6577 XThC.Tn[3].n18 VGND 0.14703f
C6578 XThC.Tn[3].t36 VGND 0.01826f
C6579 XThC.Tn[3].t31 VGND 0.01994f
C6580 XThC.Tn[3].n19 VGND 0.04453f
C6581 XThC.Tn[3].n20 VGND 0.02545f
C6582 XThC.Tn[3].n21 VGND 0.14703f
C6583 XThC.Tn[3].t23 VGND 0.01826f
C6584 XThC.Tn[3].t20 VGND 0.01994f
C6585 XThC.Tn[3].n22 VGND 0.04453f
C6586 XThC.Tn[3].n23 VGND 0.02545f
C6587 XThC.Tn[3].n24 VGND 0.14703f
C6588 XThC.Tn[3].t24 VGND 0.01826f
C6589 XThC.Tn[3].t21 VGND 0.01994f
C6590 XThC.Tn[3].n25 VGND 0.04453f
C6591 XThC.Tn[3].n26 VGND 0.02545f
C6592 XThC.Tn[3].n27 VGND 0.14703f
C6593 XThC.Tn[3].t40 VGND 0.01826f
C6594 XThC.Tn[3].t34 VGND 0.01994f
C6595 XThC.Tn[3].n28 VGND 0.04453f
C6596 XThC.Tn[3].n29 VGND 0.02545f
C6597 XThC.Tn[3].n30 VGND 0.14703f
C6598 XThC.Tn[3].t15 VGND 0.01826f
C6599 XThC.Tn[3].t43 VGND 0.01994f
C6600 XThC.Tn[3].n31 VGND 0.04453f
C6601 XThC.Tn[3].n32 VGND 0.02545f
C6602 XThC.Tn[3].n33 VGND 0.14703f
C6603 XThC.Tn[3].t17 VGND 0.01826f
C6604 XThC.Tn[3].t13 VGND 0.01994f
C6605 XThC.Tn[3].n34 VGND 0.04453f
C6606 XThC.Tn[3].n35 VGND 0.02545f
C6607 XThC.Tn[3].n36 VGND 0.14703f
C6608 XThC.Tn[3].t37 VGND 0.01826f
C6609 XThC.Tn[3].t32 VGND 0.01994f
C6610 XThC.Tn[3].n37 VGND 0.04453f
C6611 XThC.Tn[3].n38 VGND 0.02545f
C6612 XThC.Tn[3].n39 VGND 0.14703f
C6613 XThC.Tn[3].t39 VGND 0.01826f
C6614 XThC.Tn[3].t33 VGND 0.01994f
C6615 XThC.Tn[3].n40 VGND 0.04453f
C6616 XThC.Tn[3].n41 VGND 0.02545f
C6617 XThC.Tn[3].n42 VGND 0.14703f
C6618 XThC.Tn[3].t18 VGND 0.01826f
C6619 XThC.Tn[3].t14 VGND 0.01994f
C6620 XThC.Tn[3].n43 VGND 0.04453f
C6621 XThC.Tn[3].n44 VGND 0.02545f
C6622 XThC.Tn[3].n45 VGND 0.14703f
C6623 XThC.Tn[3].t26 VGND 0.01826f
C6624 XThC.Tn[3].t22 VGND 0.01994f
C6625 XThC.Tn[3].n46 VGND 0.04453f
C6626 XThC.Tn[3].n47 VGND 0.02545f
C6627 XThC.Tn[3].n48 VGND 0.14703f
C6628 XThC.Tn[3].t28 VGND 0.01826f
C6629 XThC.Tn[3].t25 VGND 0.01994f
C6630 XThC.Tn[3].n49 VGND 0.04453f
C6631 XThC.Tn[3].n50 VGND 0.02545f
C6632 XThC.Tn[3].n51 VGND 0.14703f
C6633 XThC.Tn[3].t41 VGND 0.01826f
C6634 XThC.Tn[3].t38 VGND 0.01994f
C6635 XThC.Tn[3].n52 VGND 0.04453f
C6636 XThC.Tn[3].n53 VGND 0.02545f
C6637 XThC.Tn[3].n54 VGND 0.14703f
C6638 XThC.Tn[3].t19 VGND 0.01826f
C6639 XThC.Tn[3].t16 VGND 0.01994f
C6640 XThC.Tn[3].n55 VGND 0.04453f
C6641 XThC.Tn[3].n56 VGND 0.02545f
C6642 XThC.Tn[3].n57 VGND 0.14703f
C6643 XThC.Tn[3].n58 VGND 0.07767f
C6644 XThC.Tn[1].t11 VGND 0.02257f
C6645 XThC.Tn[1].t10 VGND 0.02257f
C6646 XThC.Tn[1].n0 VGND 0.04555f
C6647 XThC.Tn[1].t9 VGND 0.02257f
C6648 XThC.Tn[1].t8 VGND 0.02257f
C6649 XThC.Tn[1].n1 VGND 0.05329f
C6650 XThC.Tn[1].n2 VGND 0.15986f
C6651 XThC.Tn[1].t5 VGND 0.01467f
C6652 XThC.Tn[1].t4 VGND 0.01467f
C6653 XThC.Tn[1].n3 VGND 0.0334f
C6654 XThC.Tn[1].t7 VGND 0.01467f
C6655 XThC.Tn[1].t6 VGND 0.01467f
C6656 XThC.Tn[1].n4 VGND 0.0334f
C6657 XThC.Tn[1].t1 VGND 0.01467f
C6658 XThC.Tn[1].t0 VGND 0.01467f
C6659 XThC.Tn[1].n5 VGND 0.0334f
C6660 XThC.Tn[1].t3 VGND 0.01467f
C6661 XThC.Tn[1].t2 VGND 0.01467f
C6662 XThC.Tn[1].n6 VGND 0.05565f
C6663 XThC.Tn[1].n7 VGND 0.15906f
C6664 XThC.Tn[1].n8 VGND 0.09833f
C6665 XThC.Tn[1].n9 VGND 0.11097f
C6666 XThC.Tn[1].t31 VGND 0.01789f
C6667 XThC.Tn[1].t29 VGND 0.01954f
C6668 XThC.Tn[1].n10 VGND 0.04363f
C6669 XThC.Tn[1].n11 VGND 0.02493f
C6670 XThC.Tn[1].n12 VGND 0.03032f
C6671 XThC.Tn[1].t17 VGND 0.01789f
C6672 XThC.Tn[1].t14 VGND 0.01954f
C6673 XThC.Tn[1].n13 VGND 0.04363f
C6674 XThC.Tn[1].n14 VGND 0.02493f
C6675 XThC.Tn[1].n15 VGND 0.14405f
C6676 XThC.Tn[1].t22 VGND 0.01789f
C6677 XThC.Tn[1].t16 VGND 0.01954f
C6678 XThC.Tn[1].n16 VGND 0.04363f
C6679 XThC.Tn[1].n17 VGND 0.02493f
C6680 XThC.Tn[1].n18 VGND 0.14405f
C6681 XThC.Tn[1].t23 VGND 0.01789f
C6682 XThC.Tn[1].t18 VGND 0.01954f
C6683 XThC.Tn[1].n19 VGND 0.04363f
C6684 XThC.Tn[1].n20 VGND 0.02493f
C6685 XThC.Tn[1].n21 VGND 0.14405f
C6686 XThC.Tn[1].t42 VGND 0.01789f
C6687 XThC.Tn[1].t39 VGND 0.01954f
C6688 XThC.Tn[1].n22 VGND 0.04363f
C6689 XThC.Tn[1].n23 VGND 0.02493f
C6690 XThC.Tn[1].n24 VGND 0.14405f
C6691 XThC.Tn[1].t43 VGND 0.01789f
C6692 XThC.Tn[1].t40 VGND 0.01954f
C6693 XThC.Tn[1].n25 VGND 0.04363f
C6694 XThC.Tn[1].n26 VGND 0.02493f
C6695 XThC.Tn[1].n27 VGND 0.14405f
C6696 XThC.Tn[1].t27 VGND 0.01789f
C6697 XThC.Tn[1].t21 VGND 0.01954f
C6698 XThC.Tn[1].n28 VGND 0.04363f
C6699 XThC.Tn[1].n29 VGND 0.02493f
C6700 XThC.Tn[1].n30 VGND 0.14405f
C6701 XThC.Tn[1].t34 VGND 0.01789f
C6702 XThC.Tn[1].t30 VGND 0.01954f
C6703 XThC.Tn[1].n31 VGND 0.04363f
C6704 XThC.Tn[1].n32 VGND 0.02493f
C6705 XThC.Tn[1].n33 VGND 0.14405f
C6706 XThC.Tn[1].t36 VGND 0.01789f
C6707 XThC.Tn[1].t32 VGND 0.01954f
C6708 XThC.Tn[1].n34 VGND 0.04363f
C6709 XThC.Tn[1].n35 VGND 0.02493f
C6710 XThC.Tn[1].n36 VGND 0.14405f
C6711 XThC.Tn[1].t24 VGND 0.01789f
C6712 XThC.Tn[1].t19 VGND 0.01954f
C6713 XThC.Tn[1].n37 VGND 0.04363f
C6714 XThC.Tn[1].n38 VGND 0.02493f
C6715 XThC.Tn[1].n39 VGND 0.14405f
C6716 XThC.Tn[1].t26 VGND 0.01789f
C6717 XThC.Tn[1].t20 VGND 0.01954f
C6718 XThC.Tn[1].n40 VGND 0.04363f
C6719 XThC.Tn[1].n41 VGND 0.02493f
C6720 XThC.Tn[1].n42 VGND 0.14405f
C6721 XThC.Tn[1].t37 VGND 0.01789f
C6722 XThC.Tn[1].t33 VGND 0.01954f
C6723 XThC.Tn[1].n43 VGND 0.04363f
C6724 XThC.Tn[1].n44 VGND 0.02493f
C6725 XThC.Tn[1].n45 VGND 0.14405f
C6726 XThC.Tn[1].t13 VGND 0.01789f
C6727 XThC.Tn[1].t41 VGND 0.01954f
C6728 XThC.Tn[1].n46 VGND 0.04363f
C6729 XThC.Tn[1].n47 VGND 0.02493f
C6730 XThC.Tn[1].n48 VGND 0.14405f
C6731 XThC.Tn[1].t15 VGND 0.01789f
C6732 XThC.Tn[1].t12 VGND 0.01954f
C6733 XThC.Tn[1].n49 VGND 0.04363f
C6734 XThC.Tn[1].n50 VGND 0.02493f
C6735 XThC.Tn[1].n51 VGND 0.14405f
C6736 XThC.Tn[1].t28 VGND 0.01789f
C6737 XThC.Tn[1].t25 VGND 0.01954f
C6738 XThC.Tn[1].n52 VGND 0.04363f
C6739 XThC.Tn[1].n53 VGND 0.02493f
C6740 XThC.Tn[1].n54 VGND 0.14405f
C6741 XThC.Tn[1].t38 VGND 0.01789f
C6742 XThC.Tn[1].t35 VGND 0.01954f
C6743 XThC.Tn[1].n55 VGND 0.04363f
C6744 XThC.Tn[1].n56 VGND 0.02493f
C6745 XThC.Tn[1].n57 VGND 0.14405f
C6746 XThC.Tn[1].n58 VGND 0.53187f
C6747 XThC.Tn[1].n59 VGND 0.05367f
C6748 Vbias.t266 VGND 0.19156f
C6749 Vbias.n0 VGND 0.20854f
C6750 Vbias.t85 VGND 0.19156f
C6751 Vbias.n1 VGND 0.20891f
C6752 Vbias.n2 VGND 0.13854f
C6753 Vbias.t180 VGND 0.19156f
C6754 Vbias.n3 VGND 0.20891f
C6755 Vbias.n4 VGND 0.13854f
C6756 Vbias.t188 VGND 0.19156f
C6757 Vbias.n5 VGND 0.20891f
C6758 Vbias.n6 VGND 0.13854f
C6759 Vbias.t21 VGND 0.19156f
C6760 Vbias.n7 VGND 0.20891f
C6761 Vbias.n8 VGND 0.13854f
C6762 Vbias.t107 VGND 0.19156f
C6763 Vbias.n9 VGND 0.20891f
C6764 Vbias.n10 VGND 0.13854f
C6765 Vbias.t190 VGND 0.19156f
C6766 Vbias.n11 VGND 0.20891f
C6767 Vbias.n12 VGND 0.13854f
C6768 Vbias.t25 VGND 0.19156f
C6769 Vbias.n13 VGND 0.20891f
C6770 Vbias.n14 VGND 0.13854f
C6771 Vbias.t45 VGND 0.19156f
C6772 Vbias.n15 VGND 0.20891f
C6773 Vbias.n16 VGND 0.13854f
C6774 Vbias.t117 VGND 0.19156f
C6775 Vbias.n17 VGND 0.20891f
C6776 Vbias.n18 VGND 0.13854f
C6777 Vbias.t208 VGND 0.19156f
C6778 Vbias.n19 VGND 0.20891f
C6779 Vbias.n20 VGND 0.13854f
C6780 Vbias.t229 VGND 0.19156f
C6781 Vbias.n21 VGND 0.20891f
C6782 Vbias.n22 VGND 0.13854f
C6783 Vbias.t120 VGND 0.19156f
C6784 Vbias.n23 VGND 0.20891f
C6785 Vbias.n24 VGND 0.13854f
C6786 Vbias.t148 VGND 0.19156f
C6787 Vbias.n25 VGND 0.20891f
C6788 Vbias.n26 VGND 0.13854f
C6789 Vbias.t157 VGND 0.19156f
C6790 Vbias.n27 VGND 0.20891f
C6791 Vbias.n28 VGND 0.13854f
C6792 Vbias.t67 VGND 0.19156f
C6793 Vbias.n29 VGND 0.20891f
C6794 Vbias.n30 VGND 0.13854f
C6795 Vbias.n31 VGND 0.58136f
C6796 Vbias.t146 VGND 0.19156f
C6797 Vbias.n32 VGND 0.20854f
C6798 Vbias.t222 VGND 0.19156f
C6799 Vbias.n33 VGND 0.20891f
C6800 Vbias.n34 VGND 0.13854f
C6801 Vbias.t65 VGND 0.19156f
C6802 Vbias.n35 VGND 0.20891f
C6803 Vbias.n36 VGND 0.13854f
C6804 Vbias.t73 VGND 0.19156f
C6805 Vbias.n37 VGND 0.20891f
C6806 Vbias.n38 VGND 0.13854f
C6807 Vbias.t158 VGND 0.19156f
C6808 Vbias.n39 VGND 0.20891f
C6809 Vbias.n40 VGND 0.13854f
C6810 Vbias.t251 VGND 0.19156f
C6811 Vbias.n41 VGND 0.20891f
C6812 Vbias.n42 VGND 0.13854f
C6813 Vbias.t78 VGND 0.19156f
C6814 Vbias.n43 VGND 0.20891f
C6815 Vbias.n44 VGND 0.13854f
C6816 Vbias.t164 VGND 0.19156f
C6817 Vbias.n45 VGND 0.20891f
C6818 Vbias.n46 VGND 0.13854f
C6819 Vbias.t184 VGND 0.19156f
C6820 Vbias.n47 VGND 0.20891f
C6821 Vbias.n48 VGND 0.13854f
C6822 Vbias.t260 VGND 0.19156f
C6823 Vbias.n49 VGND 0.20891f
C6824 Vbias.n50 VGND 0.13854f
C6825 Vbias.t90 VGND 0.19156f
C6826 Vbias.n51 VGND 0.20891f
C6827 Vbias.n52 VGND 0.13854f
C6828 Vbias.t112 VGND 0.19156f
C6829 Vbias.n53 VGND 0.20891f
C6830 Vbias.n54 VGND 0.13854f
C6831 Vbias.t265 VGND 0.19156f
C6832 Vbias.n55 VGND 0.20891f
C6833 Vbias.n56 VGND 0.13854f
C6834 Vbias.t32 VGND 0.19156f
C6835 Vbias.n57 VGND 0.20891f
C6836 Vbias.n58 VGND 0.13854f
C6837 Vbias.t41 VGND 0.19156f
C6838 Vbias.n59 VGND 0.20891f
C6839 Vbias.n60 VGND 0.13854f
C6840 Vbias.t200 VGND 0.19156f
C6841 Vbias.n61 VGND 0.20891f
C6842 Vbias.n62 VGND 0.13854f
C6843 Vbias.n63 VGND 0.5981f
C6844 Vbias.t221 VGND 0.19156f
C6845 Vbias.n64 VGND 0.20854f
C6846 Vbias.t37 VGND 0.19156f
C6847 Vbias.n65 VGND 0.20891f
C6848 Vbias.n66 VGND 0.13854f
C6849 Vbias.t138 VGND 0.19156f
C6850 Vbias.n67 VGND 0.20891f
C6851 Vbias.n68 VGND 0.13854f
C6852 Vbias.t145 VGND 0.19156f
C6853 Vbias.n69 VGND 0.20891f
C6854 Vbias.n70 VGND 0.13854f
C6855 Vbias.t230 VGND 0.19156f
C6856 Vbias.n71 VGND 0.20891f
C6857 Vbias.n72 VGND 0.13854f
C6858 Vbias.t64 VGND 0.19156f
C6859 Vbias.n73 VGND 0.20891f
C6860 Vbias.n74 VGND 0.13854f
C6861 Vbias.t151 VGND 0.19156f
C6862 Vbias.n75 VGND 0.20891f
C6863 Vbias.n76 VGND 0.13854f
C6864 Vbias.t236 VGND 0.19156f
C6865 Vbias.n77 VGND 0.20891f
C6866 Vbias.n78 VGND 0.13854f
C6867 Vbias.t259 VGND 0.19156f
C6868 Vbias.n79 VGND 0.20891f
C6869 Vbias.n80 VGND 0.13854f
C6870 Vbias.t77 VGND 0.19156f
C6871 Vbias.n81 VGND 0.20891f
C6872 Vbias.n82 VGND 0.13854f
C6873 Vbias.t163 VGND 0.19156f
C6874 Vbias.n83 VGND 0.20891f
C6875 Vbias.n84 VGND 0.13854f
C6876 Vbias.t183 VGND 0.19156f
C6877 Vbias.n85 VGND 0.20891f
C6878 Vbias.n86 VGND 0.13854f
C6879 Vbias.t83 VGND 0.19156f
C6880 Vbias.n87 VGND 0.20891f
C6881 Vbias.n88 VGND 0.13854f
C6882 Vbias.t103 VGND 0.19156f
C6883 Vbias.n89 VGND 0.20891f
C6884 Vbias.n90 VGND 0.13854f
C6885 Vbias.t110 VGND 0.19156f
C6886 Vbias.n91 VGND 0.20891f
C6887 Vbias.n92 VGND 0.13854f
C6888 Vbias.t19 VGND 0.19156f
C6889 Vbias.n93 VGND 0.20891f
C6890 Vbias.n94 VGND 0.13854f
C6891 Vbias.n95 VGND 0.5981f
C6892 Vbias.t36 VGND 0.19156f
C6893 Vbias.n96 VGND 0.20854f
C6894 Vbias.t106 VGND 0.19156f
C6895 Vbias.n97 VGND 0.20891f
C6896 Vbias.n98 VGND 0.13854f
C6897 Vbias.t209 VGND 0.19156f
C6898 Vbias.n99 VGND 0.20891f
C6899 Vbias.n100 VGND 0.13854f
C6900 Vbias.t220 VGND 0.19156f
C6901 Vbias.n101 VGND 0.20891f
C6902 Vbias.n102 VGND 0.13854f
C6903 Vbias.t44 VGND 0.19156f
C6904 Vbias.n103 VGND 0.20891f
C6905 Vbias.n104 VGND 0.13854f
C6906 Vbias.t137 VGND 0.19156f
C6907 Vbias.n105 VGND 0.20891f
C6908 Vbias.n106 VGND 0.13854f
C6909 Vbias.t224 VGND 0.19156f
C6910 Vbias.n107 VGND 0.20891f
C6911 Vbias.n108 VGND 0.13854f
C6912 Vbias.t48 VGND 0.19156f
C6913 Vbias.n109 VGND 0.20891f
C6914 Vbias.n110 VGND 0.13854f
C6915 Vbias.t76 VGND 0.19156f
C6916 Vbias.n111 VGND 0.20891f
C6917 Vbias.n112 VGND 0.13854f
C6918 Vbias.t149 VGND 0.19156f
C6919 Vbias.n113 VGND 0.20891f
C6920 Vbias.n114 VGND 0.13854f
C6921 Vbias.t234 VGND 0.19156f
C6922 Vbias.n115 VGND 0.20891f
C6923 Vbias.n116 VGND 0.13854f
C6924 Vbias.t258 VGND 0.19156f
C6925 Vbias.n117 VGND 0.20891f
C6926 Vbias.n118 VGND 0.13854f
C6927 Vbias.t154 VGND 0.19156f
C6928 Vbias.n119 VGND 0.20891f
C6929 Vbias.n120 VGND 0.13854f
C6930 Vbias.t176 VGND 0.19156f
C6931 Vbias.n121 VGND 0.20891f
C6932 Vbias.n122 VGND 0.13854f
C6933 Vbias.t181 VGND 0.19156f
C6934 Vbias.n123 VGND 0.20891f
C6935 Vbias.n124 VGND 0.13854f
C6936 Vbias.t92 VGND 0.19156f
C6937 Vbias.n125 VGND 0.20891f
C6938 Vbias.n126 VGND 0.13854f
C6939 Vbias.n127 VGND 0.5981f
C6940 Vbias.t192 VGND 0.19156f
C6941 Vbias.n128 VGND 0.20854f
C6942 Vbias.t12 VGND 0.19156f
C6943 Vbias.n129 VGND 0.20891f
C6944 Vbias.n130 VGND 0.13854f
C6945 Vbias.t109 VGND 0.19156f
C6946 Vbias.n131 VGND 0.20891f
C6947 Vbias.n132 VGND 0.13854f
C6948 Vbias.t121 VGND 0.19156f
C6949 Vbias.n133 VGND 0.20891f
C6950 Vbias.n134 VGND 0.13854f
C6951 Vbias.t212 VGND 0.19156f
C6952 Vbias.n135 VGND 0.20891f
C6953 Vbias.n136 VGND 0.13854f
C6954 Vbias.t40 VGND 0.19156f
C6955 Vbias.n137 VGND 0.20891f
C6956 Vbias.n138 VGND 0.13854f
C6957 Vbias.t122 VGND 0.19156f
C6958 Vbias.n139 VGND 0.20891f
C6959 Vbias.n140 VGND 0.13854f
C6960 Vbias.t215 VGND 0.19156f
C6961 Vbias.n141 VGND 0.20891f
C6962 Vbias.n142 VGND 0.13854f
C6963 Vbias.t237 VGND 0.19156f
C6964 Vbias.n143 VGND 0.20891f
C6965 Vbias.n144 VGND 0.13854f
C6966 Vbias.t49 VGND 0.19156f
C6967 Vbias.n145 VGND 0.20891f
C6968 Vbias.n146 VGND 0.13854f
C6969 Vbias.t140 VGND 0.19156f
C6970 Vbias.n147 VGND 0.20891f
C6971 Vbias.n148 VGND 0.13854f
C6972 Vbias.t165 VGND 0.19156f
C6973 Vbias.n149 VGND 0.20891f
C6974 Vbias.n150 VGND 0.13854f
C6975 Vbias.t53 VGND 0.19156f
C6976 Vbias.n151 VGND 0.20891f
C6977 Vbias.n152 VGND 0.13854f
C6978 Vbias.t84 VGND 0.19156f
C6979 Vbias.n153 VGND 0.20891f
C6980 Vbias.n154 VGND 0.13854f
C6981 Vbias.t91 VGND 0.19156f
C6982 Vbias.n155 VGND 0.20891f
C6983 Vbias.n156 VGND 0.13854f
C6984 Vbias.t255 VGND 0.19156f
C6985 Vbias.n157 VGND 0.20891f
C6986 Vbias.n158 VGND 0.13854f
C6987 Vbias.n159 VGND 0.5981f
C6988 Vbias.t61 VGND 0.19156f
C6989 Vbias.n160 VGND 0.20854f
C6990 Vbias.t134 VGND 0.19156f
C6991 Vbias.n161 VGND 0.20891f
C6992 Vbias.n162 VGND 0.13854f
C6993 Vbias.t232 VGND 0.19156f
C6994 Vbias.n163 VGND 0.20891f
C6995 Vbias.n164 VGND 0.13854f
C6996 Vbias.t247 VGND 0.19156f
C6997 Vbias.n165 VGND 0.20891f
C6998 Vbias.n166 VGND 0.13854f
C6999 Vbias.t72 VGND 0.19156f
C7000 Vbias.n167 VGND 0.20891f
C7001 Vbias.n168 VGND 0.13854f
C7002 Vbias.t161 VGND 0.19156f
C7003 Vbias.n169 VGND 0.20891f
C7004 Vbias.n170 VGND 0.13854f
C7005 Vbias.t250 VGND 0.19156f
C7006 Vbias.n171 VGND 0.20891f
C7007 Vbias.n172 VGND 0.13854f
C7008 Vbias.t80 VGND 0.19156f
C7009 Vbias.n173 VGND 0.20891f
C7010 Vbias.n174 VGND 0.13854f
C7011 Vbias.t100 VGND 0.19156f
C7012 Vbias.n175 VGND 0.20891f
C7013 Vbias.n176 VGND 0.13854f
C7014 Vbias.t173 VGND 0.19156f
C7015 Vbias.n177 VGND 0.20891f
C7016 Vbias.n178 VGND 0.13854f
C7017 Vbias.t262 VGND 0.19156f
C7018 Vbias.n179 VGND 0.20891f
C7019 Vbias.n180 VGND 0.13854f
C7020 Vbias.t28 VGND 0.19156f
C7021 Vbias.n181 VGND 0.20891f
C7022 Vbias.n182 VGND 0.13854f
C7023 Vbias.t178 VGND 0.19156f
C7024 Vbias.n183 VGND 0.20891f
C7025 Vbias.n184 VGND 0.13854f
C7026 Vbias.t197 VGND 0.19156f
C7027 Vbias.n185 VGND 0.20891f
C7028 Vbias.n186 VGND 0.13854f
C7029 Vbias.t213 VGND 0.19156f
C7030 Vbias.n187 VGND 0.20891f
C7031 Vbias.n188 VGND 0.13854f
C7032 Vbias.t115 VGND 0.19156f
C7033 Vbias.n189 VGND 0.20891f
C7034 Vbias.n190 VGND 0.13854f
C7035 Vbias.n191 VGND 0.5981f
C7036 Vbias.t195 VGND 0.19156f
C7037 Vbias.n192 VGND 0.20854f
C7038 Vbias.t16 VGND 0.19156f
C7039 Vbias.n193 VGND 0.20891f
C7040 Vbias.n194 VGND 0.13854f
C7041 Vbias.t114 VGND 0.19156f
C7042 Vbias.n195 VGND 0.20891f
C7043 Vbias.n196 VGND 0.13854f
C7044 Vbias.t123 VGND 0.19156f
C7045 Vbias.n197 VGND 0.20891f
C7046 Vbias.n198 VGND 0.13854f
C7047 Vbias.t214 VGND 0.19156f
C7048 Vbias.n199 VGND 0.20891f
C7049 Vbias.n200 VGND 0.13854f
C7050 Vbias.t42 VGND 0.19156f
C7051 Vbias.n201 VGND 0.20891f
C7052 Vbias.n202 VGND 0.13854f
C7053 Vbias.t126 VGND 0.19156f
C7054 Vbias.n203 VGND 0.20891f
C7055 Vbias.n204 VGND 0.13854f
C7056 Vbias.t218 VGND 0.19156f
C7057 Vbias.n205 VGND 0.20891f
C7058 Vbias.n206 VGND 0.13854f
C7059 Vbias.t240 VGND 0.19156f
C7060 Vbias.n207 VGND 0.20891f
C7061 Vbias.n208 VGND 0.13854f
C7062 Vbias.t52 VGND 0.19156f
C7063 Vbias.n209 VGND 0.20891f
C7064 Vbias.n210 VGND 0.13854f
C7065 Vbias.t142 VGND 0.19156f
C7066 Vbias.n211 VGND 0.20891f
C7067 Vbias.n212 VGND 0.13854f
C7068 Vbias.t168 VGND 0.19156f
C7069 Vbias.n213 VGND 0.20891f
C7070 Vbias.n214 VGND 0.13854f
C7071 Vbias.t57 VGND 0.19156f
C7072 Vbias.n215 VGND 0.20891f
C7073 Vbias.n216 VGND 0.13854f
C7074 Vbias.t86 VGND 0.19156f
C7075 Vbias.n217 VGND 0.20891f
C7076 Vbias.n218 VGND 0.13854f
C7077 Vbias.t95 VGND 0.19156f
C7078 Vbias.n219 VGND 0.20891f
C7079 Vbias.n220 VGND 0.13854f
C7080 Vbias.t256 VGND 0.19156f
C7081 Vbias.n221 VGND 0.20891f
C7082 Vbias.n222 VGND 0.13854f
C7083 Vbias.n223 VGND 0.5981f
C7084 Vbias.t15 VGND 0.19156f
C7085 Vbias.n224 VGND 0.20854f
C7086 Vbias.t89 VGND 0.19156f
C7087 Vbias.n225 VGND 0.20891f
C7088 Vbias.n226 VGND 0.13854f
C7089 Vbias.t186 VGND 0.19156f
C7090 Vbias.n227 VGND 0.20891f
C7091 Vbias.n228 VGND 0.13854f
C7092 Vbias.t194 VGND 0.19156f
C7093 Vbias.n229 VGND 0.20891f
C7094 Vbias.n230 VGND 0.13854f
C7095 Vbias.t29 VGND 0.19156f
C7096 Vbias.n231 VGND 0.20891f
C7097 Vbias.n232 VGND 0.13854f
C7098 Vbias.t113 VGND 0.19156f
C7099 Vbias.n233 VGND 0.20891f
C7100 Vbias.n234 VGND 0.13854f
C7101 Vbias.t198 VGND 0.19156f
C7102 Vbias.n235 VGND 0.20891f
C7103 Vbias.n236 VGND 0.13854f
C7104 Vbias.t34 VGND 0.19156f
C7105 Vbias.n237 VGND 0.20891f
C7106 Vbias.n238 VGND 0.13854f
C7107 Vbias.t51 VGND 0.19156f
C7108 Vbias.n239 VGND 0.20891f
C7109 Vbias.n240 VGND 0.13854f
C7110 Vbias.t125 VGND 0.19156f
C7111 Vbias.n241 VGND 0.20891f
C7112 Vbias.n242 VGND 0.13854f
C7113 Vbias.t217 VGND 0.19156f
C7114 Vbias.n243 VGND 0.20891f
C7115 Vbias.n244 VGND 0.13854f
C7116 Vbias.t239 VGND 0.19156f
C7117 Vbias.n245 VGND 0.20891f
C7118 Vbias.n246 VGND 0.13854f
C7119 Vbias.t129 VGND 0.19156f
C7120 Vbias.n247 VGND 0.20891f
C7121 Vbias.n248 VGND 0.13854f
C7122 Vbias.t155 VGND 0.19156f
C7123 Vbias.n249 VGND 0.20891f
C7124 Vbias.n250 VGND 0.13854f
C7125 Vbias.t167 VGND 0.19156f
C7126 Vbias.n251 VGND 0.20891f
C7127 Vbias.n252 VGND 0.13854f
C7128 Vbias.t70 VGND 0.19156f
C7129 Vbias.n253 VGND 0.20891f
C7130 Vbias.n254 VGND 0.13854f
C7131 Vbias.n255 VGND 0.5981f
C7132 Vbias.t88 VGND 0.19156f
C7133 Vbias.n256 VGND 0.20854f
C7134 Vbias.t160 VGND 0.19156f
C7135 Vbias.n257 VGND 0.20891f
C7136 Vbias.n258 VGND 0.13854f
C7137 Vbias.t263 VGND 0.19156f
C7138 Vbias.n259 VGND 0.20891f
C7139 Vbias.n260 VGND 0.13854f
C7140 Vbias.t14 VGND 0.19156f
C7141 Vbias.n261 VGND 0.20891f
C7142 Vbias.n262 VGND 0.13854f
C7143 Vbias.t99 VGND 0.19156f
C7144 Vbias.n263 VGND 0.20891f
C7145 Vbias.n264 VGND 0.13854f
C7146 Vbias.t185 VGND 0.19156f
C7147 Vbias.n265 VGND 0.20891f
C7148 Vbias.n266 VGND 0.13854f
C7149 Vbias.t17 VGND 0.19156f
C7150 Vbias.n267 VGND 0.20891f
C7151 Vbias.n268 VGND 0.13854f
C7152 Vbias.t104 VGND 0.19156f
C7153 Vbias.n269 VGND 0.20891f
C7154 Vbias.n270 VGND 0.13854f
C7155 Vbias.t124 VGND 0.19156f
C7156 Vbias.n271 VGND 0.20891f
C7157 Vbias.n272 VGND 0.13854f
C7158 Vbias.t196 VGND 0.19156f
C7159 Vbias.n273 VGND 0.20891f
C7160 Vbias.n274 VGND 0.13854f
C7161 Vbias.t33 VGND 0.19156f
C7162 Vbias.n275 VGND 0.20891f
C7163 Vbias.n276 VGND 0.13854f
C7164 Vbias.t50 VGND 0.19156f
C7165 Vbias.n277 VGND 0.20891f
C7166 Vbias.n278 VGND 0.13854f
C7167 Vbias.t203 VGND 0.19156f
C7168 Vbias.n279 VGND 0.20891f
C7169 Vbias.n280 VGND 0.13854f
C7170 Vbias.t226 VGND 0.19156f
C7171 Vbias.n281 VGND 0.20891f
C7172 Vbias.n282 VGND 0.13854f
C7173 Vbias.t238 VGND 0.19156f
C7174 Vbias.n283 VGND 0.20891f
C7175 Vbias.n284 VGND 0.13854f
C7176 Vbias.t143 VGND 0.19156f
C7177 Vbias.n285 VGND 0.20891f
C7178 Vbias.n286 VGND 0.13854f
C7179 Vbias.n287 VGND 0.5981f
C7180 Vbias.t55 VGND 0.19156f
C7181 Vbias.n288 VGND 0.20854f
C7182 Vbias.t128 VGND 0.19156f
C7183 Vbias.n289 VGND 0.20891f
C7184 Vbias.n290 VGND 0.13854f
C7185 Vbias.t228 VGND 0.19156f
C7186 Vbias.n291 VGND 0.20891f
C7187 Vbias.n292 VGND 0.13854f
C7188 Vbias.t241 VGND 0.19156f
C7189 Vbias.n293 VGND 0.20891f
C7190 Vbias.n294 VGND 0.13854f
C7191 Vbias.t69 VGND 0.19156f
C7192 Vbias.n295 VGND 0.20891f
C7193 Vbias.n296 VGND 0.13854f
C7194 Vbias.t156 VGND 0.19156f
C7195 Vbias.n297 VGND 0.20891f
C7196 Vbias.n298 VGND 0.13854f
C7197 Vbias.t243 VGND 0.19156f
C7198 Vbias.n299 VGND 0.20891f
C7199 Vbias.n300 VGND 0.13854f
C7200 Vbias.t74 VGND 0.19156f
C7201 Vbias.n301 VGND 0.20891f
C7202 Vbias.n302 VGND 0.13854f
C7203 Vbias.t97 VGND 0.19156f
C7204 Vbias.n303 VGND 0.20891f
C7205 Vbias.n304 VGND 0.13854f
C7206 Vbias.t170 VGND 0.19156f
C7207 Vbias.n305 VGND 0.20891f
C7208 Vbias.n306 VGND 0.13854f
C7209 Vbias.t257 VGND 0.19156f
C7210 Vbias.n307 VGND 0.20891f
C7211 Vbias.n308 VGND 0.13854f
C7212 Vbias.t27 VGND 0.19156f
C7213 Vbias.n309 VGND 0.20891f
C7214 Vbias.n310 VGND 0.13854f
C7215 Vbias.t174 VGND 0.19156f
C7216 Vbias.n311 VGND 0.20891f
C7217 Vbias.n312 VGND 0.13854f
C7218 Vbias.t193 VGND 0.19156f
C7219 Vbias.n313 VGND 0.20891f
C7220 Vbias.n314 VGND 0.13854f
C7221 Vbias.t210 VGND 0.19156f
C7222 Vbias.n315 VGND 0.20891f
C7223 Vbias.n316 VGND 0.13854f
C7224 Vbias.t111 VGND 0.19156f
C7225 Vbias.n317 VGND 0.20891f
C7226 Vbias.n318 VGND 0.13854f
C7227 Vbias.n319 VGND 0.5981f
C7228 Vbias.t127 VGND 0.19156f
C7229 Vbias.n320 VGND 0.20854f
C7230 Vbias.t201 VGND 0.19156f
C7231 Vbias.n321 VGND 0.20891f
C7232 Vbias.n322 VGND 0.13854f
C7233 Vbias.t43 VGND 0.19156f
C7234 Vbias.n323 VGND 0.20891f
C7235 Vbias.n324 VGND 0.13854f
C7236 Vbias.t54 VGND 0.19156f
C7237 Vbias.n325 VGND 0.20891f
C7238 Vbias.n326 VGND 0.13854f
C7239 Vbias.t141 VGND 0.19156f
C7240 Vbias.n327 VGND 0.20891f
C7241 Vbias.n328 VGND 0.13854f
C7242 Vbias.t227 VGND 0.19156f
C7243 Vbias.n329 VGND 0.20891f
C7244 Vbias.n330 VGND 0.13854f
C7245 Vbias.t56 VGND 0.19156f
C7246 Vbias.n331 VGND 0.20891f
C7247 Vbias.n332 VGND 0.13854f
C7248 Vbias.t144 VGND 0.19156f
C7249 Vbias.n333 VGND 0.20891f
C7250 Vbias.n334 VGND 0.13854f
C7251 Vbias.t169 VGND 0.19156f
C7252 Vbias.n335 VGND 0.20891f
C7253 Vbias.n336 VGND 0.13854f
C7254 Vbias.t242 VGND 0.19156f
C7255 Vbias.n337 VGND 0.20891f
C7256 Vbias.n338 VGND 0.13854f
C7257 Vbias.t71 VGND 0.19156f
C7258 Vbias.n339 VGND 0.20891f
C7259 Vbias.n340 VGND 0.13854f
C7260 Vbias.t96 VGND 0.19156f
C7261 Vbias.n341 VGND 0.20891f
C7262 Vbias.n342 VGND 0.13854f
C7263 Vbias.t249 VGND 0.19156f
C7264 Vbias.n343 VGND 0.20891f
C7265 Vbias.n344 VGND 0.13854f
C7266 Vbias.t13 VGND 0.19156f
C7267 Vbias.n345 VGND 0.20891f
C7268 Vbias.n346 VGND 0.13854f
C7269 Vbias.t26 VGND 0.19156f
C7270 Vbias.n347 VGND 0.20891f
C7271 Vbias.n348 VGND 0.13854f
C7272 Vbias.t182 VGND 0.19156f
C7273 Vbias.n349 VGND 0.20891f
C7274 Vbias.n350 VGND 0.13854f
C7275 Vbias.n351 VGND 0.5981f
C7276 Vbias.t204 VGND 0.19156f
C7277 Vbias.n352 VGND 0.20854f
C7278 Vbias.t23 VGND 0.19156f
C7279 Vbias.n353 VGND 0.20891f
C7280 Vbias.n354 VGND 0.13854f
C7281 Vbias.t119 VGND 0.19156f
C7282 Vbias.n355 VGND 0.20891f
C7283 Vbias.n356 VGND 0.13854f
C7284 Vbias.t130 VGND 0.19156f
C7285 Vbias.n357 VGND 0.20891f
C7286 Vbias.n358 VGND 0.13854f
C7287 Vbias.t219 VGND 0.19156f
C7288 Vbias.n359 VGND 0.20891f
C7289 Vbias.n360 VGND 0.13854f
C7290 Vbias.t46 VGND 0.19156f
C7291 Vbias.n361 VGND 0.20891f
C7292 Vbias.n362 VGND 0.13854f
C7293 Vbias.t133 VGND 0.19156f
C7294 Vbias.n363 VGND 0.20891f
C7295 Vbias.n364 VGND 0.13854f
C7296 Vbias.t225 VGND 0.19156f
C7297 Vbias.n365 VGND 0.20891f
C7298 Vbias.n366 VGND 0.13854f
C7299 Vbias.t246 VGND 0.19156f
C7300 Vbias.n367 VGND 0.20891f
C7301 Vbias.n368 VGND 0.13854f
C7302 Vbias.t60 VGND 0.19156f
C7303 Vbias.n369 VGND 0.20891f
C7304 Vbias.n370 VGND 0.13854f
C7305 Vbias.t150 VGND 0.19156f
C7306 Vbias.n371 VGND 0.20891f
C7307 Vbias.n372 VGND 0.13854f
C7308 Vbias.t172 VGND 0.19156f
C7309 Vbias.n373 VGND 0.20891f
C7310 Vbias.n374 VGND 0.13854f
C7311 Vbias.t68 VGND 0.19156f
C7312 Vbias.n375 VGND 0.20891f
C7313 Vbias.n376 VGND 0.13854f
C7314 Vbias.t87 VGND 0.19156f
C7315 Vbias.n377 VGND 0.20891f
C7316 Vbias.n378 VGND 0.13854f
C7317 Vbias.t98 VGND 0.19156f
C7318 Vbias.n379 VGND 0.20891f
C7319 Vbias.n380 VGND 0.13854f
C7320 Vbias.t261 VGND 0.19156f
C7321 Vbias.n381 VGND 0.20891f
C7322 Vbias.n382 VGND 0.13854f
C7323 Vbias.n383 VGND 0.5981f
C7324 Vbias.t22 VGND 0.19156f
C7325 Vbias.n384 VGND 0.20854f
C7326 Vbias.t94 VGND 0.19156f
C7327 Vbias.n385 VGND 0.20891f
C7328 Vbias.n386 VGND 0.13854f
C7329 Vbias.t191 VGND 0.19156f
C7330 Vbias.n387 VGND 0.20891f
C7331 Vbias.n388 VGND 0.13854f
C7332 Vbias.t202 VGND 0.19156f
C7333 Vbias.n389 VGND 0.20891f
C7334 Vbias.n390 VGND 0.13854f
C7335 Vbias.t35 VGND 0.19156f
C7336 Vbias.n391 VGND 0.20891f
C7337 Vbias.n392 VGND 0.13854f
C7338 Vbias.t118 VGND 0.19156f
C7339 Vbias.n393 VGND 0.20891f
C7340 Vbias.n394 VGND 0.13854f
C7341 Vbias.t206 VGND 0.19156f
C7342 Vbias.n395 VGND 0.20891f
C7343 Vbias.n396 VGND 0.13854f
C7344 Vbias.t39 VGND 0.19156f
C7345 Vbias.n397 VGND 0.20891f
C7346 Vbias.n398 VGND 0.13854f
C7347 Vbias.t59 VGND 0.19156f
C7348 Vbias.n399 VGND 0.20891f
C7349 Vbias.n400 VGND 0.13854f
C7350 Vbias.t132 VGND 0.19156f
C7351 Vbias.n401 VGND 0.20891f
C7352 Vbias.n402 VGND 0.13854f
C7353 Vbias.t223 VGND 0.19156f
C7354 Vbias.n403 VGND 0.20891f
C7355 Vbias.n404 VGND 0.13854f
C7356 Vbias.t245 VGND 0.19156f
C7357 Vbias.n405 VGND 0.20891f
C7358 Vbias.n406 VGND 0.13854f
C7359 Vbias.t139 VGND 0.19156f
C7360 Vbias.n407 VGND 0.20891f
C7361 Vbias.n408 VGND 0.13854f
C7362 Vbias.t159 VGND 0.19156f
C7363 Vbias.n409 VGND 0.20891f
C7364 Vbias.n410 VGND 0.13854f
C7365 Vbias.t171 VGND 0.19156f
C7366 Vbias.n411 VGND 0.20891f
C7367 Vbias.n412 VGND 0.13854f
C7368 Vbias.t79 VGND 0.19156f
C7369 Vbias.n413 VGND 0.20891f
C7370 Vbias.n414 VGND 0.13854f
C7371 Vbias.n415 VGND 0.5981f
C7372 Vbias.t93 VGND 0.19156f
C7373 Vbias.n416 VGND 0.20854f
C7374 Vbias.t166 VGND 0.19156f
C7375 Vbias.n417 VGND 0.20891f
C7376 Vbias.n418 VGND 0.13854f
C7377 Vbias.t267 VGND 0.19156f
C7378 Vbias.n419 VGND 0.20891f
C7379 Vbias.n420 VGND 0.13854f
C7380 Vbias.t20 VGND 0.19156f
C7381 Vbias.n421 VGND 0.20891f
C7382 Vbias.n422 VGND 0.13854f
C7383 Vbias.t105 VGND 0.19156f
C7384 Vbias.n423 VGND 0.20891f
C7385 Vbias.n424 VGND 0.13854f
C7386 Vbias.t189 VGND 0.19156f
C7387 Vbias.n425 VGND 0.20891f
C7388 Vbias.n426 VGND 0.13854f
C7389 Vbias.t24 VGND 0.19156f
C7390 Vbias.n427 VGND 0.20891f
C7391 Vbias.n428 VGND 0.13854f
C7392 Vbias.t108 VGND 0.19156f
C7393 Vbias.n429 VGND 0.20891f
C7394 Vbias.n430 VGND 0.13854f
C7395 Vbias.t131 VGND 0.19156f
C7396 Vbias.n431 VGND 0.20891f
C7397 Vbias.n432 VGND 0.13854f
C7398 Vbias.t205 VGND 0.19156f
C7399 Vbias.n433 VGND 0.20891f
C7400 Vbias.n434 VGND 0.13854f
C7401 Vbias.t38 VGND 0.19156f
C7402 Vbias.n435 VGND 0.20891f
C7403 Vbias.n436 VGND 0.13854f
C7404 Vbias.t58 VGND 0.19156f
C7405 Vbias.n437 VGND 0.20891f
C7406 Vbias.n438 VGND 0.13854f
C7407 Vbias.t211 VGND 0.19156f
C7408 Vbias.n439 VGND 0.20891f
C7409 Vbias.n440 VGND 0.13854f
C7410 Vbias.t231 VGND 0.19156f
C7411 Vbias.n441 VGND 0.20891f
C7412 Vbias.n442 VGND 0.13854f
C7413 Vbias.t244 VGND 0.19156f
C7414 Vbias.n443 VGND 0.20891f
C7415 Vbias.n444 VGND 0.13854f
C7416 Vbias.t152 VGND 0.19156f
C7417 Vbias.n445 VGND 0.20891f
C7418 Vbias.n446 VGND 0.13854f
C7419 Vbias.n447 VGND 0.5981f
C7420 Vbias.t63 VGND 0.19156f
C7421 Vbias.n448 VGND 0.20854f
C7422 Vbias.t136 VGND 0.19156f
C7423 Vbias.n449 VGND 0.20891f
C7424 Vbias.n450 VGND 0.13854f
C7425 Vbias.t235 VGND 0.19156f
C7426 Vbias.n451 VGND 0.20891f
C7427 Vbias.n452 VGND 0.13854f
C7428 Vbias.t248 VGND 0.19156f
C7429 Vbias.n453 VGND 0.20891f
C7430 Vbias.n454 VGND 0.13854f
C7431 Vbias.t75 VGND 0.19156f
C7432 Vbias.n455 VGND 0.20891f
C7433 Vbias.n456 VGND 0.13854f
C7434 Vbias.t162 VGND 0.19156f
C7435 Vbias.n457 VGND 0.20891f
C7436 Vbias.n458 VGND 0.13854f
C7437 Vbias.t253 VGND 0.19156f
C7438 Vbias.n459 VGND 0.20891f
C7439 Vbias.n460 VGND 0.13854f
C7440 Vbias.t82 VGND 0.19156f
C7441 Vbias.n461 VGND 0.20891f
C7442 Vbias.n462 VGND 0.13854f
C7443 Vbias.t102 VGND 0.19156f
C7444 Vbias.n463 VGND 0.20891f
C7445 Vbias.n464 VGND 0.13854f
C7446 Vbias.t177 VGND 0.19156f
C7447 Vbias.n465 VGND 0.20891f
C7448 Vbias.n466 VGND 0.13854f
C7449 Vbias.t264 VGND 0.19156f
C7450 Vbias.n467 VGND 0.20891f
C7451 Vbias.n468 VGND 0.13854f
C7452 Vbias.t31 VGND 0.19156f
C7453 Vbias.n469 VGND 0.20891f
C7454 Vbias.n470 VGND 0.13854f
C7455 Vbias.t179 VGND 0.19156f
C7456 Vbias.n471 VGND 0.20891f
C7457 Vbias.n472 VGND 0.13854f
C7458 Vbias.t199 VGND 0.19156f
C7459 Vbias.n473 VGND 0.20891f
C7460 Vbias.n474 VGND 0.13854f
C7461 Vbias.t216 VGND 0.19156f
C7462 Vbias.n475 VGND 0.20891f
C7463 Vbias.n476 VGND 0.13854f
C7464 Vbias.t116 VGND 0.19156f
C7465 Vbias.n477 VGND 0.20891f
C7466 Vbias.n478 VGND 0.13854f
C7467 Vbias.n479 VGND 0.5981f
C7468 Vbias.t135 VGND 0.19156f
C7469 Vbias.n480 VGND 0.20854f
C7470 Vbias.t207 VGND 0.19156f
C7471 Vbias.n481 VGND 0.20891f
C7472 Vbias.n482 VGND 0.13854f
C7473 Vbias.t47 VGND 0.19156f
C7474 Vbias.n483 VGND 0.20891f
C7475 Vbias.n484 VGND 0.13854f
C7476 Vbias.t62 VGND 0.19156f
C7477 Vbias.n485 VGND 0.20891f
C7478 Vbias.n486 VGND 0.13854f
C7479 Vbias.t147 VGND 0.19156f
C7480 Vbias.n487 VGND 0.20891f
C7481 Vbias.n488 VGND 0.13854f
C7482 Vbias.t233 VGND 0.19156f
C7483 Vbias.n489 VGND 0.20891f
C7484 Vbias.n490 VGND 0.13854f
C7485 Vbias.t66 VGND 0.19156f
C7486 Vbias.n491 VGND 0.20891f
C7487 Vbias.n492 VGND 0.13854f
C7488 Vbias.t153 VGND 0.19156f
C7489 Vbias.n493 VGND 0.20891f
C7490 Vbias.n494 VGND 0.13854f
C7491 Vbias.t175 VGND 0.19156f
C7492 Vbias.n495 VGND 0.20891f
C7493 Vbias.n496 VGND 0.13854f
C7494 Vbias.t252 VGND 0.19156f
C7495 Vbias.n497 VGND 0.20891f
C7496 Vbias.n498 VGND 0.13854f
C7497 Vbias.t81 VGND 0.19156f
C7498 Vbias.n499 VGND 0.20891f
C7499 Vbias.n500 VGND 0.13854f
C7500 Vbias.t101 VGND 0.19156f
C7501 Vbias.n501 VGND 0.20891f
C7502 Vbias.n502 VGND 0.13854f
C7503 Vbias.t254 VGND 0.19156f
C7504 Vbias.n503 VGND 0.20891f
C7505 Vbias.n504 VGND 0.13854f
C7506 Vbias.t18 VGND 0.19156f
C7507 Vbias.n505 VGND 0.20891f
C7508 Vbias.n506 VGND 0.13854f
C7509 Vbias.t30 VGND 0.19156f
C7510 Vbias.n507 VGND 0.20891f
C7511 Vbias.n508 VGND 0.13854f
C7512 Vbias.t187 VGND 0.19156f
C7513 Vbias.n509 VGND 0.20891f
C7514 Vbias.n510 VGND 0.13854f
C7515 Vbias.n511 VGND 0.69561f
C7516 Vbias.t5 VGND 0.19054f
C7517 Vbias.n512 VGND 0.64623f
C7518 Vbias.t8 VGND 0.02796f
C7519 Vbias.t3 VGND 0.02796f
C7520 Vbias.n513 VGND 0.05942f
C7521 Vbias.t2 VGND 0.01763f
C7522 Vbias.t9 VGND 0.01763f
C7523 Vbias.n514 VGND 0.0375f
C7524 Vbias.n515 VGND 2.50332f
C7525 Vbias.t4 VGND 0.36737f
C7526 Vbias.n516 VGND 0.42109f
C7527 Vbias.n517 VGND 0.23222f
C7528 Vbias.t7 VGND 0.19054f
C7529 Vbias.n518 VGND 0.59823f
C7530 Vbias.t10 VGND 0.02796f
C7531 Vbias.t11 VGND 0.02796f
C7532 Vbias.n519 VGND 0.05942f
C7533 Vbias.t1 VGND 0.01763f
C7534 Vbias.t0 VGND 0.01763f
C7535 Vbias.n520 VGND 0.0375f
C7536 Vbias.n521 VGND 2.50332f
C7537 Vbias.t6 VGND 0.36731f
C7538 Vbias.n522 VGND 0.42109f
C7539 Vbias.n523 VGND 0.21429f
C7540 Vbias.n524 VGND 1.99477f
C7541 XThC.Tn[2].t10 VGND 0.02306f
C7542 XThC.Tn[2].t9 VGND 0.02306f
C7543 XThC.Tn[2].n0 VGND 0.04655f
C7544 XThC.Tn[2].t8 VGND 0.02306f
C7545 XThC.Tn[2].t7 VGND 0.02306f
C7546 XThC.Tn[2].n1 VGND 0.05447f
C7547 XThC.Tn[2].n2 VGND 0.15249f
C7548 XThC.Tn[2].t6 VGND 0.01499f
C7549 XThC.Tn[2].t5 VGND 0.01499f
C7550 XThC.Tn[2].n3 VGND 0.03414f
C7551 XThC.Tn[2].t4 VGND 0.01499f
C7552 XThC.Tn[2].t3 VGND 0.01499f
C7553 XThC.Tn[2].n4 VGND 0.03414f
C7554 XThC.Tn[2].t1 VGND 0.01499f
C7555 XThC.Tn[2].t2 VGND 0.01499f
C7556 XThC.Tn[2].n5 VGND 0.03414f
C7557 XThC.Tn[2].t11 VGND 0.01499f
C7558 XThC.Tn[2].t0 VGND 0.01499f
C7559 XThC.Tn[2].n6 VGND 0.05688f
C7560 XThC.Tn[2].n7 VGND 0.16258f
C7561 XThC.Tn[2].n8 VGND 0.1005f
C7562 XThC.Tn[2].n9 VGND 0.11343f
C7563 XThC.Tn[2].t20 VGND 0.01828f
C7564 XThC.Tn[2].t18 VGND 0.01997f
C7565 XThC.Tn[2].n10 VGND 0.04459f
C7566 XThC.Tn[2].n11 VGND 0.02548f
C7567 XThC.Tn[2].n12 VGND 0.03099f
C7568 XThC.Tn[2].t38 VGND 0.01828f
C7569 XThC.Tn[2].t35 VGND 0.01997f
C7570 XThC.Tn[2].n13 VGND 0.04459f
C7571 XThC.Tn[2].n14 VGND 0.02548f
C7572 XThC.Tn[2].n15 VGND 0.14724f
C7573 XThC.Tn[2].t43 VGND 0.01828f
C7574 XThC.Tn[2].t37 VGND 0.01997f
C7575 XThC.Tn[2].n16 VGND 0.04459f
C7576 XThC.Tn[2].n17 VGND 0.02548f
C7577 XThC.Tn[2].n18 VGND 0.14724f
C7578 XThC.Tn[2].t12 VGND 0.01828f
C7579 XThC.Tn[2].t39 VGND 0.01997f
C7580 XThC.Tn[2].n19 VGND 0.04459f
C7581 XThC.Tn[2].n20 VGND 0.02548f
C7582 XThC.Tn[2].n21 VGND 0.14724f
C7583 XThC.Tn[2].t31 VGND 0.01828f
C7584 XThC.Tn[2].t28 VGND 0.01997f
C7585 XThC.Tn[2].n22 VGND 0.04459f
C7586 XThC.Tn[2].n23 VGND 0.02548f
C7587 XThC.Tn[2].n24 VGND 0.14724f
C7588 XThC.Tn[2].t32 VGND 0.01828f
C7589 XThC.Tn[2].t29 VGND 0.01997f
C7590 XThC.Tn[2].n25 VGND 0.04459f
C7591 XThC.Tn[2].n26 VGND 0.02548f
C7592 XThC.Tn[2].n27 VGND 0.14724f
C7593 XThC.Tn[2].t16 VGND 0.01828f
C7594 XThC.Tn[2].t42 VGND 0.01997f
C7595 XThC.Tn[2].n28 VGND 0.04459f
C7596 XThC.Tn[2].n29 VGND 0.02548f
C7597 XThC.Tn[2].n30 VGND 0.14724f
C7598 XThC.Tn[2].t23 VGND 0.01828f
C7599 XThC.Tn[2].t19 VGND 0.01997f
C7600 XThC.Tn[2].n31 VGND 0.04459f
C7601 XThC.Tn[2].n32 VGND 0.02548f
C7602 XThC.Tn[2].n33 VGND 0.14724f
C7603 XThC.Tn[2].t25 VGND 0.01828f
C7604 XThC.Tn[2].t21 VGND 0.01997f
C7605 XThC.Tn[2].n34 VGND 0.04459f
C7606 XThC.Tn[2].n35 VGND 0.02548f
C7607 XThC.Tn[2].n36 VGND 0.14724f
C7608 XThC.Tn[2].t13 VGND 0.01828f
C7609 XThC.Tn[2].t40 VGND 0.01997f
C7610 XThC.Tn[2].n37 VGND 0.04459f
C7611 XThC.Tn[2].n38 VGND 0.02548f
C7612 XThC.Tn[2].n39 VGND 0.14724f
C7613 XThC.Tn[2].t15 VGND 0.01828f
C7614 XThC.Tn[2].t41 VGND 0.01997f
C7615 XThC.Tn[2].n40 VGND 0.04459f
C7616 XThC.Tn[2].n41 VGND 0.02548f
C7617 XThC.Tn[2].n42 VGND 0.14724f
C7618 XThC.Tn[2].t26 VGND 0.01828f
C7619 XThC.Tn[2].t22 VGND 0.01997f
C7620 XThC.Tn[2].n43 VGND 0.04459f
C7621 XThC.Tn[2].n44 VGND 0.02548f
C7622 XThC.Tn[2].n45 VGND 0.14724f
C7623 XThC.Tn[2].t34 VGND 0.01828f
C7624 XThC.Tn[2].t30 VGND 0.01997f
C7625 XThC.Tn[2].n46 VGND 0.04459f
C7626 XThC.Tn[2].n47 VGND 0.02548f
C7627 XThC.Tn[2].n48 VGND 0.14724f
C7628 XThC.Tn[2].t36 VGND 0.01828f
C7629 XThC.Tn[2].t33 VGND 0.01997f
C7630 XThC.Tn[2].n49 VGND 0.04459f
C7631 XThC.Tn[2].n50 VGND 0.02548f
C7632 XThC.Tn[2].n51 VGND 0.14724f
C7633 XThC.Tn[2].t17 VGND 0.01828f
C7634 XThC.Tn[2].t14 VGND 0.01997f
C7635 XThC.Tn[2].n52 VGND 0.04459f
C7636 XThC.Tn[2].n53 VGND 0.02548f
C7637 XThC.Tn[2].n54 VGND 0.14724f
C7638 XThC.Tn[2].t27 VGND 0.01828f
C7639 XThC.Tn[2].t24 VGND 0.01997f
C7640 XThC.Tn[2].n55 VGND 0.04459f
C7641 XThC.Tn[2].n56 VGND 0.02548f
C7642 XThC.Tn[2].n57 VGND 0.14724f
C7643 XThC.Tn[2].n58 VGND 0.53552f
C7644 XThC.Tn[2].n59 VGND 0.08697f
C7645 XThC.Tn[2].n60 VGND 0.04826f
C7646 XThC.Tn[4].t9 VGND 0.02356f
C7647 XThC.Tn[4].t8 VGND 0.02356f
C7648 XThC.Tn[4].n0 VGND 0.04755f
C7649 XThC.Tn[4].t11 VGND 0.02356f
C7650 XThC.Tn[4].t10 VGND 0.02356f
C7651 XThC.Tn[4].n1 VGND 0.05564f
C7652 XThC.Tn[4].n2 VGND 0.15575f
C7653 XThC.Tn[4].t5 VGND 0.01531f
C7654 XThC.Tn[4].t4 VGND 0.01531f
C7655 XThC.Tn[4].n3 VGND 0.03487f
C7656 XThC.Tn[4].t7 VGND 0.01531f
C7657 XThC.Tn[4].t6 VGND 0.01531f
C7658 XThC.Tn[4].n4 VGND 0.03487f
C7659 XThC.Tn[4].t2 VGND 0.01531f
C7660 XThC.Tn[4].t1 VGND 0.01531f
C7661 XThC.Tn[4].n5 VGND 0.03487f
C7662 XThC.Tn[4].t0 VGND 0.01531f
C7663 XThC.Tn[4].t3 VGND 0.01531f
C7664 XThC.Tn[4].n6 VGND 0.0581f
C7665 XThC.Tn[4].n7 VGND 0.16606f
C7666 XThC.Tn[4].n8 VGND 0.10265f
C7667 XThC.Tn[4].n9 VGND 0.11585f
C7668 XThC.Tn[4].t28 VGND 0.01867f
C7669 XThC.Tn[4].t26 VGND 0.0204f
C7670 XThC.Tn[4].n10 VGND 0.04555f
C7671 XThC.Tn[4].n11 VGND 0.02603f
C7672 XThC.Tn[4].n12 VGND 0.03166f
C7673 XThC.Tn[4].t14 VGND 0.01867f
C7674 XThC.Tn[4].t43 VGND 0.0204f
C7675 XThC.Tn[4].n13 VGND 0.04555f
C7676 XThC.Tn[4].n14 VGND 0.02603f
C7677 XThC.Tn[4].n15 VGND 0.15039f
C7678 XThC.Tn[4].t19 VGND 0.01867f
C7679 XThC.Tn[4].t13 VGND 0.0204f
C7680 XThC.Tn[4].n16 VGND 0.04555f
C7681 XThC.Tn[4].n17 VGND 0.02603f
C7682 XThC.Tn[4].n18 VGND 0.15039f
C7683 XThC.Tn[4].t20 VGND 0.01867f
C7684 XThC.Tn[4].t15 VGND 0.0204f
C7685 XThC.Tn[4].n19 VGND 0.04555f
C7686 XThC.Tn[4].n20 VGND 0.02603f
C7687 XThC.Tn[4].n21 VGND 0.15039f
C7688 XThC.Tn[4].t39 VGND 0.01867f
C7689 XThC.Tn[4].t36 VGND 0.0204f
C7690 XThC.Tn[4].n22 VGND 0.04555f
C7691 XThC.Tn[4].n23 VGND 0.02603f
C7692 XThC.Tn[4].n24 VGND 0.15039f
C7693 XThC.Tn[4].t40 VGND 0.01867f
C7694 XThC.Tn[4].t37 VGND 0.0204f
C7695 XThC.Tn[4].n25 VGND 0.04555f
C7696 XThC.Tn[4].n26 VGND 0.02603f
C7697 XThC.Tn[4].n27 VGND 0.15039f
C7698 XThC.Tn[4].t24 VGND 0.01867f
C7699 XThC.Tn[4].t18 VGND 0.0204f
C7700 XThC.Tn[4].n28 VGND 0.04555f
C7701 XThC.Tn[4].n29 VGND 0.02603f
C7702 XThC.Tn[4].n30 VGND 0.15039f
C7703 XThC.Tn[4].t31 VGND 0.01867f
C7704 XThC.Tn[4].t27 VGND 0.0204f
C7705 XThC.Tn[4].n31 VGND 0.04555f
C7706 XThC.Tn[4].n32 VGND 0.02603f
C7707 XThC.Tn[4].n33 VGND 0.15039f
C7708 XThC.Tn[4].t33 VGND 0.01867f
C7709 XThC.Tn[4].t29 VGND 0.0204f
C7710 XThC.Tn[4].n34 VGND 0.04555f
C7711 XThC.Tn[4].n35 VGND 0.02603f
C7712 XThC.Tn[4].n36 VGND 0.15039f
C7713 XThC.Tn[4].t21 VGND 0.01867f
C7714 XThC.Tn[4].t16 VGND 0.0204f
C7715 XThC.Tn[4].n37 VGND 0.04555f
C7716 XThC.Tn[4].n38 VGND 0.02603f
C7717 XThC.Tn[4].n39 VGND 0.15039f
C7718 XThC.Tn[4].t23 VGND 0.01867f
C7719 XThC.Tn[4].t17 VGND 0.0204f
C7720 XThC.Tn[4].n40 VGND 0.04555f
C7721 XThC.Tn[4].n41 VGND 0.02603f
C7722 XThC.Tn[4].n42 VGND 0.15039f
C7723 XThC.Tn[4].t34 VGND 0.01867f
C7724 XThC.Tn[4].t30 VGND 0.0204f
C7725 XThC.Tn[4].n43 VGND 0.04555f
C7726 XThC.Tn[4].n44 VGND 0.02603f
C7727 XThC.Tn[4].n45 VGND 0.15039f
C7728 XThC.Tn[4].t42 VGND 0.01867f
C7729 XThC.Tn[4].t38 VGND 0.0204f
C7730 XThC.Tn[4].n46 VGND 0.04555f
C7731 XThC.Tn[4].n47 VGND 0.02603f
C7732 XThC.Tn[4].n48 VGND 0.15039f
C7733 XThC.Tn[4].t12 VGND 0.01867f
C7734 XThC.Tn[4].t41 VGND 0.0204f
C7735 XThC.Tn[4].n49 VGND 0.04555f
C7736 XThC.Tn[4].n50 VGND 0.02603f
C7737 XThC.Tn[4].n51 VGND 0.15039f
C7738 XThC.Tn[4].t25 VGND 0.01867f
C7739 XThC.Tn[4].t22 VGND 0.0204f
C7740 XThC.Tn[4].n52 VGND 0.04555f
C7741 XThC.Tn[4].n53 VGND 0.02603f
C7742 XThC.Tn[4].n54 VGND 0.15039f
C7743 XThC.Tn[4].t35 VGND 0.01867f
C7744 XThC.Tn[4].t32 VGND 0.0204f
C7745 XThC.Tn[4].n55 VGND 0.04555f
C7746 XThC.Tn[4].n56 VGND 0.02603f
C7747 XThC.Tn[4].n57 VGND 0.15039f
C7748 XThC.Tn[4].n58 VGND 0.46855f
C7749 XThC.Tn[4].n59 VGND 0.08903f
C7750 XThC.Tn[4].n60 VGND 0.0493f
C7751 XThR.Tn[5].t8 VGND 0.01426f
C7752 XThR.Tn[5].t9 VGND 0.01426f
C7753 XThR.Tn[5].n0 VGND 0.05411f
C7754 XThR.Tn[5].t11 VGND 0.01426f
C7755 XThR.Tn[5].t10 VGND 0.01426f
C7756 XThR.Tn[5].n1 VGND 0.03247f
C7757 XThR.Tn[5].n2 VGND 0.15464f
C7758 XThR.Tn[5].t6 VGND 0.01426f
C7759 XThR.Tn[5].t5 VGND 0.01426f
C7760 XThR.Tn[5].n3 VGND 0.03247f
C7761 XThR.Tn[5].n4 VGND 0.0956f
C7762 XThR.Tn[5].t7 VGND 0.01426f
C7763 XThR.Tn[5].t4 VGND 0.01426f
C7764 XThR.Tn[5].n5 VGND 0.03247f
C7765 XThR.Tn[5].n6 VGND 0.10789f
C7766 XThR.Tn[5].t17 VGND 0.01715f
C7767 XThR.Tn[5].t72 VGND 0.01877f
C7768 XThR.Tn[5].n7 VGND 0.04585f
C7769 XThR.Tn[5].n8 VGND 0.07125f
C7770 XThR.Tn[5].t39 VGND 0.01715f
C7771 XThR.Tn[5].t26 VGND 0.01877f
C7772 XThR.Tn[5].n9 VGND 0.04585f
C7773 XThR.Tn[5].t13 VGND 0.01709f
C7774 XThR.Tn[5].t23 VGND 0.01871f
C7775 XThR.Tn[5].n10 VGND 0.0477f
C7776 XThR.Tn[5].n11 VGND 0.03351f
C7777 XThR.Tn[5].n13 VGND 0.10754f
C7778 XThR.Tn[5].t73 VGND 0.01715f
C7779 XThR.Tn[5].t66 VGND 0.01877f
C7780 XThR.Tn[5].n14 VGND 0.04585f
C7781 XThR.Tn[5].t48 VGND 0.01709f
C7782 XThR.Tn[5].t61 VGND 0.01871f
C7783 XThR.Tn[5].n15 VGND 0.0477f
C7784 XThR.Tn[5].n16 VGND 0.03351f
C7785 XThR.Tn[5].n18 VGND 0.10754f
C7786 XThR.Tn[5].t28 VGND 0.01715f
C7787 XThR.Tn[5].t21 VGND 0.01877f
C7788 XThR.Tn[5].n19 VGND 0.04585f
C7789 XThR.Tn[5].t65 VGND 0.01709f
C7790 XThR.Tn[5].t18 VGND 0.01871f
C7791 XThR.Tn[5].n20 VGND 0.0477f
C7792 XThR.Tn[5].n21 VGND 0.03351f
C7793 XThR.Tn[5].n23 VGND 0.10754f
C7794 XThR.Tn[5].t55 VGND 0.01715f
C7795 XThR.Tn[5].t51 VGND 0.01877f
C7796 XThR.Tn[5].n24 VGND 0.04585f
C7797 XThR.Tn[5].t33 VGND 0.01709f
C7798 XThR.Tn[5].t46 VGND 0.01871f
C7799 XThR.Tn[5].n25 VGND 0.0477f
C7800 XThR.Tn[5].n26 VGND 0.03351f
C7801 XThR.Tn[5].n28 VGND 0.10754f
C7802 XThR.Tn[5].t30 VGND 0.01715f
C7803 XThR.Tn[5].t22 VGND 0.01877f
C7804 XThR.Tn[5].n29 VGND 0.04585f
C7805 XThR.Tn[5].t67 VGND 0.01709f
C7806 XThR.Tn[5].t19 VGND 0.01871f
C7807 XThR.Tn[5].n30 VGND 0.0477f
C7808 XThR.Tn[5].n31 VGND 0.03351f
C7809 XThR.Tn[5].n33 VGND 0.10754f
C7810 XThR.Tn[5].t69 VGND 0.01715f
C7811 XThR.Tn[5].t40 VGND 0.01877f
C7812 XThR.Tn[5].n34 VGND 0.04585f
C7813 XThR.Tn[5].t43 VGND 0.01709f
C7814 XThR.Tn[5].t37 VGND 0.01871f
C7815 XThR.Tn[5].n35 VGND 0.0477f
C7816 XThR.Tn[5].n36 VGND 0.03351f
C7817 XThR.Tn[5].n38 VGND 0.10754f
C7818 XThR.Tn[5].t38 VGND 0.01715f
C7819 XThR.Tn[5].t32 VGND 0.01877f
C7820 XThR.Tn[5].n39 VGND 0.04585f
C7821 XThR.Tn[5].t14 VGND 0.01709f
C7822 XThR.Tn[5].t29 VGND 0.01871f
C7823 XThR.Tn[5].n40 VGND 0.0477f
C7824 XThR.Tn[5].n41 VGND 0.03351f
C7825 XThR.Tn[5].n43 VGND 0.10754f
C7826 XThR.Tn[5].t42 VGND 0.01715f
C7827 XThR.Tn[5].t49 VGND 0.01877f
C7828 XThR.Tn[5].n44 VGND 0.04585f
C7829 XThR.Tn[5].t16 VGND 0.01709f
C7830 XThR.Tn[5].t45 VGND 0.01871f
C7831 XThR.Tn[5].n45 VGND 0.0477f
C7832 XThR.Tn[5].n46 VGND 0.03351f
C7833 XThR.Tn[5].n48 VGND 0.10754f
C7834 XThR.Tn[5].t58 VGND 0.01715f
C7835 XThR.Tn[5].t68 VGND 0.01877f
C7836 XThR.Tn[5].n49 VGND 0.04585f
C7837 XThR.Tn[5].t36 VGND 0.01709f
C7838 XThR.Tn[5].t63 VGND 0.01871f
C7839 XThR.Tn[5].n50 VGND 0.0477f
C7840 XThR.Tn[5].n51 VGND 0.03351f
C7841 XThR.Tn[5].n53 VGND 0.10754f
C7842 XThR.Tn[5].t53 VGND 0.01715f
C7843 XThR.Tn[5].t24 VGND 0.01877f
C7844 XThR.Tn[5].n54 VGND 0.04585f
C7845 XThR.Tn[5].t25 VGND 0.01709f
C7846 XThR.Tn[5].t20 VGND 0.01871f
C7847 XThR.Tn[5].n55 VGND 0.0477f
C7848 XThR.Tn[5].n56 VGND 0.03351f
C7849 XThR.Tn[5].n58 VGND 0.10754f
C7850 XThR.Tn[5].t71 VGND 0.01715f
C7851 XThR.Tn[5].t60 VGND 0.01877f
C7852 XThR.Tn[5].n59 VGND 0.04585f
C7853 XThR.Tn[5].t44 VGND 0.01709f
C7854 XThR.Tn[5].t57 VGND 0.01871f
C7855 XThR.Tn[5].n60 VGND 0.0477f
C7856 XThR.Tn[5].n61 VGND 0.03351f
C7857 XThR.Tn[5].n63 VGND 0.10754f
C7858 XThR.Tn[5].t41 VGND 0.01715f
C7859 XThR.Tn[5].t35 VGND 0.01877f
C7860 XThR.Tn[5].n64 VGND 0.04585f
C7861 XThR.Tn[5].t15 VGND 0.01709f
C7862 XThR.Tn[5].t31 VGND 0.01871f
C7863 XThR.Tn[5].n65 VGND 0.0477f
C7864 XThR.Tn[5].n66 VGND 0.03351f
C7865 XThR.Tn[5].n68 VGND 0.10754f
C7866 XThR.Tn[5].t56 VGND 0.01715f
C7867 XThR.Tn[5].t52 VGND 0.01877f
C7868 XThR.Tn[5].n69 VGND 0.04585f
C7869 XThR.Tn[5].t34 VGND 0.01709f
C7870 XThR.Tn[5].t47 VGND 0.01871f
C7871 XThR.Tn[5].n70 VGND 0.0477f
C7872 XThR.Tn[5].n71 VGND 0.03351f
C7873 XThR.Tn[5].n73 VGND 0.10754f
C7874 XThR.Tn[5].t12 VGND 0.01715f
C7875 XThR.Tn[5].t70 VGND 0.01877f
C7876 XThR.Tn[5].n74 VGND 0.04585f
C7877 XThR.Tn[5].t50 VGND 0.01709f
C7878 XThR.Tn[5].t64 VGND 0.01871f
C7879 XThR.Tn[5].n75 VGND 0.0477f
C7880 XThR.Tn[5].n76 VGND 0.03351f
C7881 XThR.Tn[5].n78 VGND 0.10754f
C7882 XThR.Tn[5].t54 VGND 0.01715f
C7883 XThR.Tn[5].t62 VGND 0.01877f
C7884 XThR.Tn[5].n79 VGND 0.04585f
C7885 XThR.Tn[5].t27 VGND 0.01709f
C7886 XThR.Tn[5].t59 VGND 0.01871f
C7887 XThR.Tn[5].n80 VGND 0.0477f
C7888 XThR.Tn[5].n81 VGND 0.03351f
C7889 XThR.Tn[5].n83 VGND 0.10754f
C7890 XThR.Tn[5].n84 VGND 0.09773f
C7891 XThR.Tn[5].n85 VGND 0.18927f
C7892 XThR.Tn[5].t2 VGND 0.02194f
C7893 XThR.Tn[5].t3 VGND 0.02194f
C7894 XThR.Tn[5].n86 VGND 0.04428f
C7895 XThR.Tn[5].t1 VGND 0.02194f
C7896 XThR.Tn[5].t0 VGND 0.02194f
C7897 XThR.Tn[5].n87 VGND 0.05181f
C7898 XThR.Tn[5].n88 VGND 0.14505f
C7899 XThR.Tn[5].n89 VGND 0.04591f
C7900 XThR.Tn[3].t9 VGND 0.02182f
C7901 XThR.Tn[3].t10 VGND 0.02182f
C7902 XThR.Tn[3].n0 VGND 0.04405f
C7903 XThR.Tn[3].t8 VGND 0.02182f
C7904 XThR.Tn[3].t11 VGND 0.02182f
C7905 XThR.Tn[3].n1 VGND 0.05154f
C7906 XThR.Tn[3].n2 VGND 0.14427f
C7907 XThR.Tn[3].t7 VGND 0.01418f
C7908 XThR.Tn[3].t4 VGND 0.01418f
C7909 XThR.Tn[3].n3 VGND 0.0323f
C7910 XThR.Tn[3].t6 VGND 0.01418f
C7911 XThR.Tn[3].t5 VGND 0.01418f
C7912 XThR.Tn[3].n4 VGND 0.0323f
C7913 XThR.Tn[3].t0 VGND 0.01418f
C7914 XThR.Tn[3].t1 VGND 0.01418f
C7915 XThR.Tn[3].n5 VGND 0.05382f
C7916 XThR.Tn[3].t3 VGND 0.01418f
C7917 XThR.Tn[3].t2 VGND 0.01418f
C7918 XThR.Tn[3].n6 VGND 0.0323f
C7919 XThR.Tn[3].n7 VGND 0.15382f
C7920 XThR.Tn[3].n8 VGND 0.09509f
C7921 XThR.Tn[3].n9 VGND 0.10731f
C7922 XThR.Tn[3].t64 VGND 0.01705f
C7923 XThR.Tn[3].t57 VGND 0.01867f
C7924 XThR.Tn[3].n10 VGND 0.0456f
C7925 XThR.Tn[3].n11 VGND 0.07087f
C7926 XThR.Tn[3].t18 VGND 0.01705f
C7927 XThR.Tn[3].t70 VGND 0.01867f
C7928 XThR.Tn[3].n12 VGND 0.0456f
C7929 XThR.Tn[3].t24 VGND 0.017f
C7930 XThR.Tn[3].t55 VGND 0.01861f
C7931 XThR.Tn[3].n13 VGND 0.04745f
C7932 XThR.Tn[3].n14 VGND 0.03333f
C7933 XThR.Tn[3].n16 VGND 0.10697f
C7934 XThR.Tn[3].t59 VGND 0.01705f
C7935 XThR.Tn[3].t49 VGND 0.01867f
C7936 XThR.Tn[3].n17 VGND 0.0456f
C7937 XThR.Tn[3].t62 VGND 0.017f
C7938 XThR.Tn[3].t29 VGND 0.01861f
C7939 XThR.Tn[3].n18 VGND 0.04745f
C7940 XThR.Tn[3].n19 VGND 0.03333f
C7941 XThR.Tn[3].n21 VGND 0.10697f
C7942 XThR.Tn[3].t71 VGND 0.01705f
C7943 XThR.Tn[3].t67 VGND 0.01867f
C7944 XThR.Tn[3].n22 VGND 0.0456f
C7945 XThR.Tn[3].t12 VGND 0.017f
C7946 XThR.Tn[3].t47 VGND 0.01861f
C7947 XThR.Tn[3].n23 VGND 0.04745f
C7948 XThR.Tn[3].n24 VGND 0.03333f
C7949 XThR.Tn[3].n26 VGND 0.10697f
C7950 XThR.Tn[3].t39 VGND 0.01705f
C7951 XThR.Tn[3].t33 VGND 0.01867f
C7952 XThR.Tn[3].n27 VGND 0.0456f
C7953 XThR.Tn[3].t42 VGND 0.017f
C7954 XThR.Tn[3].t13 VGND 0.01861f
C7955 XThR.Tn[3].n28 VGND 0.04745f
C7956 XThR.Tn[3].n29 VGND 0.03333f
C7957 XThR.Tn[3].n31 VGND 0.10697f
C7958 XThR.Tn[3].t72 VGND 0.01705f
C7959 XThR.Tn[3].t68 VGND 0.01867f
C7960 XThR.Tn[3].n32 VGND 0.0456f
C7961 XThR.Tn[3].t16 VGND 0.017f
C7962 XThR.Tn[3].t48 VGND 0.01861f
C7963 XThR.Tn[3].n33 VGND 0.04745f
C7964 XThR.Tn[3].n34 VGND 0.03333f
C7965 XThR.Tn[3].n36 VGND 0.10697f
C7966 XThR.Tn[3].t52 VGND 0.01705f
C7967 XThR.Tn[3].t20 VGND 0.01867f
C7968 XThR.Tn[3].n37 VGND 0.0456f
C7969 XThR.Tn[3].t56 VGND 0.017f
C7970 XThR.Tn[3].t66 VGND 0.01861f
C7971 XThR.Tn[3].n38 VGND 0.04745f
C7972 XThR.Tn[3].n39 VGND 0.03333f
C7973 XThR.Tn[3].n41 VGND 0.10697f
C7974 XThR.Tn[3].t19 VGND 0.01705f
C7975 XThR.Tn[3].t14 VGND 0.01867f
C7976 XThR.Tn[3].n42 VGND 0.0456f
C7977 XThR.Tn[3].t23 VGND 0.017f
C7978 XThR.Tn[3].t61 VGND 0.01861f
C7979 XThR.Tn[3].n43 VGND 0.04745f
C7980 XThR.Tn[3].n44 VGND 0.03333f
C7981 XThR.Tn[3].n46 VGND 0.10697f
C7982 XThR.Tn[3].t22 VGND 0.01705f
C7983 XThR.Tn[3].t31 VGND 0.01867f
C7984 XThR.Tn[3].n47 VGND 0.0456f
C7985 XThR.Tn[3].t28 VGND 0.017f
C7986 XThR.Tn[3].t73 VGND 0.01861f
C7987 XThR.Tn[3].n48 VGND 0.04745f
C7988 XThR.Tn[3].n49 VGND 0.03333f
C7989 XThR.Tn[3].n51 VGND 0.10697f
C7990 XThR.Tn[3].t41 VGND 0.01705f
C7991 XThR.Tn[3].t51 VGND 0.01867f
C7992 XThR.Tn[3].n52 VGND 0.0456f
C7993 XThR.Tn[3].t45 VGND 0.017f
C7994 XThR.Tn[3].t30 VGND 0.01861f
C7995 XThR.Tn[3].n53 VGND 0.04745f
C7996 XThR.Tn[3].n54 VGND 0.03333f
C7997 XThR.Tn[3].n56 VGND 0.10697f
C7998 XThR.Tn[3].t35 VGND 0.01705f
C7999 XThR.Tn[3].t69 VGND 0.01867f
C8000 XThR.Tn[3].n57 VGND 0.0456f
C8001 XThR.Tn[3].t37 VGND 0.017f
C8002 XThR.Tn[3].t50 VGND 0.01861f
C8003 XThR.Tn[3].n58 VGND 0.04745f
C8004 XThR.Tn[3].n59 VGND 0.03333f
C8005 XThR.Tn[3].n61 VGND 0.10697f
C8006 XThR.Tn[3].t54 VGND 0.01705f
C8007 XThR.Tn[3].t44 VGND 0.01867f
C8008 XThR.Tn[3].n62 VGND 0.0456f
C8009 XThR.Tn[3].t58 VGND 0.017f
C8010 XThR.Tn[3].t25 VGND 0.01861f
C8011 XThR.Tn[3].n63 VGND 0.04745f
C8012 XThR.Tn[3].n64 VGND 0.03333f
C8013 XThR.Tn[3].n66 VGND 0.10697f
C8014 XThR.Tn[3].t21 VGND 0.01705f
C8015 XThR.Tn[3].t17 VGND 0.01867f
C8016 XThR.Tn[3].n67 VGND 0.0456f
C8017 XThR.Tn[3].t26 VGND 0.017f
C8018 XThR.Tn[3].t63 VGND 0.01861f
C8019 XThR.Tn[3].n68 VGND 0.04745f
C8020 XThR.Tn[3].n69 VGND 0.03333f
C8021 XThR.Tn[3].n71 VGND 0.10697f
C8022 XThR.Tn[3].t40 VGND 0.01705f
C8023 XThR.Tn[3].t34 VGND 0.01867f
C8024 XThR.Tn[3].n72 VGND 0.0456f
C8025 XThR.Tn[3].t43 VGND 0.017f
C8026 XThR.Tn[3].t15 VGND 0.01861f
C8027 XThR.Tn[3].n73 VGND 0.04745f
C8028 XThR.Tn[3].n74 VGND 0.03333f
C8029 XThR.Tn[3].n76 VGND 0.10697f
C8030 XThR.Tn[3].t60 VGND 0.01705f
C8031 XThR.Tn[3].t53 VGND 0.01867f
C8032 XThR.Tn[3].n77 VGND 0.0456f
C8033 XThR.Tn[3].t65 VGND 0.017f
C8034 XThR.Tn[3].t32 VGND 0.01861f
C8035 XThR.Tn[3].n78 VGND 0.04745f
C8036 XThR.Tn[3].n79 VGND 0.03333f
C8037 XThR.Tn[3].n81 VGND 0.10697f
C8038 XThR.Tn[3].t36 VGND 0.01705f
C8039 XThR.Tn[3].t46 VGND 0.01867f
C8040 XThR.Tn[3].n82 VGND 0.0456f
C8041 XThR.Tn[3].t38 VGND 0.017f
C8042 XThR.Tn[3].t27 VGND 0.01861f
C8043 XThR.Tn[3].n83 VGND 0.04745f
C8044 XThR.Tn[3].n84 VGND 0.03333f
C8045 XThR.Tn[3].n86 VGND 0.10697f
C8046 XThR.Tn[3].n87 VGND 0.09721f
C8047 XThR.Tn[3].n88 VGND 0.2153f
C8048 XThR.Tn[3].n89 VGND 0.04566f
C8049 XThC.XTB4.Y.t1 VGND 0.12238f
C8050 XThC.XTB4.Y.n0 VGND 0.16166f
C8051 XThC.XTB4.Y.t4 VGND 0.02956f
C8052 XThC.XTB4.Y.t13 VGND 0.05016f
C8053 XThC.XTB4.Y.n1 VGND 0.05972f
C8054 XThC.XTB4.Y.t7 VGND 0.02956f
C8055 XThC.XTB4.Y.t17 VGND 0.05016f
C8056 XThC.XTB4.Y.n2 VGND 0.03074f
C8057 XThC.XTB4.Y.t10 VGND 0.02956f
C8058 XThC.XTB4.Y.t2 VGND 0.05016f
C8059 XThC.XTB4.Y.n3 VGND 0.06603f
C8060 XThC.XTB4.Y.t14 VGND 0.02956f
C8061 XThC.XTB4.Y.t3 VGND 0.05016f
C8062 XThC.XTB4.Y.n4 VGND 0.0613f
C8063 XThC.XTB4.Y.n5 VGND 0.03729f
C8064 XThC.XTB4.Y.n6 VGND 0.06174f
C8065 XThC.XTB4.Y.n7 VGND 0.02389f
C8066 XThC.XTB4.Y.n8 VGND 0.02916f
C8067 XThC.XTB4.Y.n9 VGND 0.06603f
C8068 XThC.XTB4.Y.n10 VGND 0.0331f
C8069 XThC.XTB4.Y.n11 VGND 0.06459f
C8070 XThC.XTB4.Y.t5 VGND 0.02956f
C8071 XThC.XTB4.Y.t16 VGND 0.05016f
C8072 XThC.XTB4.Y.n12 VGND 0.06761f
C8073 XThC.XTB4.Y.t9 VGND 0.02956f
C8074 XThC.XTB4.Y.t6 VGND 0.05016f
C8075 XThC.XTB4.Y.t15 VGND 0.02956f
C8076 XThC.XTB4.Y.t12 VGND 0.05016f
C8077 XThC.XTB4.Y.t11 VGND 0.02956f
C8078 XThC.XTB4.Y.t8 VGND 0.05016f
C8079 XThC.XTB4.Y.n13 VGND 0.08416f
C8080 XThC.XTB4.Y.n14 VGND 0.08889f
C8081 XThC.XTB4.Y.n15 VGND 0.03426f
C8082 XThC.XTB4.Y.n16 VGND 0.07234f
C8083 XThC.XTB4.Y.n17 VGND 0.0331f
C8084 XThC.XTB4.Y.n18 VGND 0.02701f
C8085 XThC.XTB4.Y.n19 VGND 0.63971f
C8086 XThC.XTB4.Y.n20 VGND 1.29767f
C8087 XThC.XTB4.Y.n21 VGND 0.08408f
C8088 XThC.XTB4.Y.t0 VGND 0.06491f
C8089 XThC.XTB4.Y.n22 VGND 0.04329f
C8090 XThC.Tn[0].t11 VGND 0.01472f
C8091 XThC.Tn[0].t8 VGND 0.01472f
C8092 XThC.Tn[0].n0 VGND 0.05586f
C8093 XThC.Tn[0].t9 VGND 0.01472f
C8094 XThC.Tn[0].t10 VGND 0.01472f
C8095 XThC.Tn[0].n1 VGND 0.03353f
C8096 XThC.Tn[0].n2 VGND 0.15966f
C8097 XThC.Tn[0].t7 VGND 0.01472f
C8098 XThC.Tn[0].t6 VGND 0.01472f
C8099 XThC.Tn[0].n3 VGND 0.03353f
C8100 XThC.Tn[0].n4 VGND 0.0987f
C8101 XThC.Tn[0].t5 VGND 0.01472f
C8102 XThC.Tn[0].t4 VGND 0.01472f
C8103 XThC.Tn[0].n5 VGND 0.03353f
C8104 XThC.Tn[0].n6 VGND 0.11139f
C8105 XThC.Tn[0].t18 VGND 0.01795f
C8106 XThC.Tn[0].t22 VGND 0.01961f
C8107 XThC.Tn[0].n7 VGND 0.04379f
C8108 XThC.Tn[0].n8 VGND 0.02502f
C8109 XThC.Tn[0].n9 VGND 0.03044f
C8110 XThC.Tn[0].t35 VGND 0.01795f
C8111 XThC.Tn[0].t41 VGND 0.01961f
C8112 XThC.Tn[0].n10 VGND 0.04379f
C8113 XThC.Tn[0].n11 VGND 0.02502f
C8114 XThC.Tn[0].n12 VGND 0.14459f
C8115 XThC.Tn[0].t37 VGND 0.01795f
C8116 XThC.Tn[0].t12 VGND 0.01961f
C8117 XThC.Tn[0].n13 VGND 0.04379f
C8118 XThC.Tn[0].n14 VGND 0.02502f
C8119 XThC.Tn[0].n15 VGND 0.14459f
C8120 XThC.Tn[0].t39 VGND 0.01795f
C8121 XThC.Tn[0].t13 VGND 0.01961f
C8122 XThC.Tn[0].n16 VGND 0.04379f
C8123 XThC.Tn[0].n17 VGND 0.02502f
C8124 XThC.Tn[0].n18 VGND 0.14459f
C8125 XThC.Tn[0].t28 VGND 0.01795f
C8126 XThC.Tn[0].t32 VGND 0.01961f
C8127 XThC.Tn[0].n19 VGND 0.04379f
C8128 XThC.Tn[0].n20 VGND 0.02502f
C8129 XThC.Tn[0].n21 VGND 0.14459f
C8130 XThC.Tn[0].t30 VGND 0.01795f
C8131 XThC.Tn[0].t34 VGND 0.01961f
C8132 XThC.Tn[0].n22 VGND 0.04379f
C8133 XThC.Tn[0].n23 VGND 0.02502f
C8134 XThC.Tn[0].n24 VGND 0.14459f
C8135 XThC.Tn[0].t43 VGND 0.01795f
C8136 XThC.Tn[0].t17 VGND 0.01961f
C8137 XThC.Tn[0].n25 VGND 0.04379f
C8138 XThC.Tn[0].n26 VGND 0.02502f
C8139 XThC.Tn[0].n27 VGND 0.14459f
C8140 XThC.Tn[0].t20 VGND 0.01795f
C8141 XThC.Tn[0].t25 VGND 0.01961f
C8142 XThC.Tn[0].n28 VGND 0.04379f
C8143 XThC.Tn[0].n29 VGND 0.02502f
C8144 XThC.Tn[0].n30 VGND 0.14459f
C8145 XThC.Tn[0].t21 VGND 0.01795f
C8146 XThC.Tn[0].t26 VGND 0.01961f
C8147 XThC.Tn[0].n31 VGND 0.04379f
C8148 XThC.Tn[0].n32 VGND 0.02502f
C8149 XThC.Tn[0].n33 VGND 0.14459f
C8150 XThC.Tn[0].t40 VGND 0.01795f
C8151 XThC.Tn[0].t15 VGND 0.01961f
C8152 XThC.Tn[0].n34 VGND 0.04379f
C8153 XThC.Tn[0].n35 VGND 0.02502f
C8154 XThC.Tn[0].n36 VGND 0.14459f
C8155 XThC.Tn[0].t42 VGND 0.01795f
C8156 XThC.Tn[0].t16 VGND 0.01961f
C8157 XThC.Tn[0].n37 VGND 0.04379f
C8158 XThC.Tn[0].n38 VGND 0.02502f
C8159 XThC.Tn[0].n39 VGND 0.14459f
C8160 XThC.Tn[0].t23 VGND 0.01795f
C8161 XThC.Tn[0].t27 VGND 0.01961f
C8162 XThC.Tn[0].n40 VGND 0.04379f
C8163 XThC.Tn[0].n41 VGND 0.02502f
C8164 XThC.Tn[0].n42 VGND 0.14459f
C8165 XThC.Tn[0].t31 VGND 0.01795f
C8166 XThC.Tn[0].t36 VGND 0.01961f
C8167 XThC.Tn[0].n43 VGND 0.04379f
C8168 XThC.Tn[0].n44 VGND 0.02502f
C8169 XThC.Tn[0].n45 VGND 0.14459f
C8170 XThC.Tn[0].t33 VGND 0.01795f
C8171 XThC.Tn[0].t38 VGND 0.01961f
C8172 XThC.Tn[0].n46 VGND 0.04379f
C8173 XThC.Tn[0].n47 VGND 0.02502f
C8174 XThC.Tn[0].n48 VGND 0.14459f
C8175 XThC.Tn[0].t14 VGND 0.01795f
C8176 XThC.Tn[0].t19 VGND 0.01961f
C8177 XThC.Tn[0].n49 VGND 0.04379f
C8178 XThC.Tn[0].n50 VGND 0.02502f
C8179 XThC.Tn[0].n51 VGND 0.14459f
C8180 XThC.Tn[0].t24 VGND 0.01795f
C8181 XThC.Tn[0].t29 VGND 0.01961f
C8182 XThC.Tn[0].n52 VGND 0.04379f
C8183 XThC.Tn[0].n53 VGND 0.02502f
C8184 XThC.Tn[0].n54 VGND 0.14459f
C8185 XThC.Tn[0].n55 VGND 0.25855f
C8186 XThC.Tn[0].n56 VGND 0.06554f
C8187 XThC.Tn[0].t1 VGND 0.02265f
C8188 XThC.Tn[0].t0 VGND 0.02265f
C8189 XThC.Tn[0].n57 VGND 0.04572f
C8190 XThC.Tn[0].t3 VGND 0.02265f
C8191 XThC.Tn[0].t2 VGND 0.02265f
C8192 XThC.Tn[0].n58 VGND 0.05349f
C8193 XThC.Tn[0].n59 VGND 0.14975f
C8194 XThC.Tn[0].n60 VGND 0.0474f
C8195 XThC.Tn[13].t7 VGND 0.01633f
C8196 XThC.Tn[13].t5 VGND 0.01633f
C8197 XThC.Tn[13].n0 VGND 0.04073f
C8198 XThC.Tn[13].t4 VGND 0.01633f
C8199 XThC.Tn[13].t6 VGND 0.01633f
C8200 XThC.Tn[13].n1 VGND 0.03266f
C8201 XThC.Tn[13].n2 VGND 0.07532f
C8202 XThC.Tn[13].t29 VGND 0.01991f
C8203 XThC.Tn[13].t27 VGND 0.02175f
C8204 XThC.Tn[13].n3 VGND 0.04858f
C8205 XThC.Tn[13].n4 VGND 0.02776f
C8206 XThC.Tn[13].n5 VGND 0.03376f
C8207 XThC.Tn[13].t15 VGND 0.01991f
C8208 XThC.Tn[13].t12 VGND 0.02175f
C8209 XThC.Tn[13].n6 VGND 0.04858f
C8210 XThC.Tn[13].n7 VGND 0.02776f
C8211 XThC.Tn[13].n8 VGND 0.1604f
C8212 XThC.Tn[13].t20 VGND 0.01991f
C8213 XThC.Tn[13].t14 VGND 0.02175f
C8214 XThC.Tn[13].n9 VGND 0.04858f
C8215 XThC.Tn[13].n10 VGND 0.02776f
C8216 XThC.Tn[13].n11 VGND 0.1604f
C8217 XThC.Tn[13].t21 VGND 0.01991f
C8218 XThC.Tn[13].t16 VGND 0.02175f
C8219 XThC.Tn[13].n12 VGND 0.04858f
C8220 XThC.Tn[13].n13 VGND 0.02776f
C8221 XThC.Tn[13].n14 VGND 0.1604f
C8222 XThC.Tn[13].t40 VGND 0.01991f
C8223 XThC.Tn[13].t37 VGND 0.02175f
C8224 XThC.Tn[13].n15 VGND 0.04858f
C8225 XThC.Tn[13].n16 VGND 0.02776f
C8226 XThC.Tn[13].n17 VGND 0.1604f
C8227 XThC.Tn[13].t41 VGND 0.01991f
C8228 XThC.Tn[13].t38 VGND 0.02175f
C8229 XThC.Tn[13].n18 VGND 0.04858f
C8230 XThC.Tn[13].n19 VGND 0.02776f
C8231 XThC.Tn[13].n20 VGND 0.1604f
C8232 XThC.Tn[13].t25 VGND 0.01991f
C8233 XThC.Tn[13].t19 VGND 0.02175f
C8234 XThC.Tn[13].n21 VGND 0.04858f
C8235 XThC.Tn[13].n22 VGND 0.02776f
C8236 XThC.Tn[13].n23 VGND 0.1604f
C8237 XThC.Tn[13].t32 VGND 0.01991f
C8238 XThC.Tn[13].t28 VGND 0.02175f
C8239 XThC.Tn[13].n24 VGND 0.04858f
C8240 XThC.Tn[13].n25 VGND 0.02776f
C8241 XThC.Tn[13].n26 VGND 0.1604f
C8242 XThC.Tn[13].t34 VGND 0.01991f
C8243 XThC.Tn[13].t30 VGND 0.02175f
C8244 XThC.Tn[13].n27 VGND 0.04858f
C8245 XThC.Tn[13].n28 VGND 0.02776f
C8246 XThC.Tn[13].n29 VGND 0.1604f
C8247 XThC.Tn[13].t22 VGND 0.01991f
C8248 XThC.Tn[13].t17 VGND 0.02175f
C8249 XThC.Tn[13].n30 VGND 0.04858f
C8250 XThC.Tn[13].n31 VGND 0.02776f
C8251 XThC.Tn[13].n32 VGND 0.1604f
C8252 XThC.Tn[13].t24 VGND 0.01991f
C8253 XThC.Tn[13].t18 VGND 0.02175f
C8254 XThC.Tn[13].n33 VGND 0.04858f
C8255 XThC.Tn[13].n34 VGND 0.02776f
C8256 XThC.Tn[13].n35 VGND 0.1604f
C8257 XThC.Tn[13].t35 VGND 0.01991f
C8258 XThC.Tn[13].t31 VGND 0.02175f
C8259 XThC.Tn[13].n36 VGND 0.04858f
C8260 XThC.Tn[13].n37 VGND 0.02776f
C8261 XThC.Tn[13].n38 VGND 0.1604f
C8262 XThC.Tn[13].t43 VGND 0.01991f
C8263 XThC.Tn[13].t39 VGND 0.02175f
C8264 XThC.Tn[13].n39 VGND 0.04858f
C8265 XThC.Tn[13].n40 VGND 0.02776f
C8266 XThC.Tn[13].n41 VGND 0.1604f
C8267 XThC.Tn[13].t13 VGND 0.01991f
C8268 XThC.Tn[13].t42 VGND 0.02175f
C8269 XThC.Tn[13].n42 VGND 0.04858f
C8270 XThC.Tn[13].n43 VGND 0.02776f
C8271 XThC.Tn[13].n44 VGND 0.1604f
C8272 XThC.Tn[13].t26 VGND 0.01991f
C8273 XThC.Tn[13].t23 VGND 0.02175f
C8274 XThC.Tn[13].n45 VGND 0.04858f
C8275 XThC.Tn[13].n46 VGND 0.02776f
C8276 XThC.Tn[13].n47 VGND 0.1604f
C8277 XThC.Tn[13].t36 VGND 0.01991f
C8278 XThC.Tn[13].t33 VGND 0.02175f
C8279 XThC.Tn[13].n48 VGND 0.04858f
C8280 XThC.Tn[13].n49 VGND 0.02776f
C8281 XThC.Tn[13].n50 VGND 0.1604f
C8282 XThC.Tn[13].n51 VGND 0.88865f
C8283 XThC.Tn[13].n52 VGND 0.07271f
C8284 XThC.Tn[13].t10 VGND 0.02513f
C8285 XThC.Tn[13].t9 VGND 0.02513f
C8286 XThC.Tn[13].n53 VGND 0.05429f
C8287 XThC.Tn[13].t8 VGND 0.02513f
C8288 XThC.Tn[13].t11 VGND 0.02513f
C8289 XThC.Tn[13].n54 VGND 0.08557f
C8290 XThC.Tn[13].n55 VGND 0.22664f
C8291 XThC.Tn[13].n56 VGND 0.01669f
C8292 XThC.Tn[13].t1 VGND 0.02513f
C8293 XThC.Tn[13].t0 VGND 0.02513f
C8294 XThC.Tn[13].n57 VGND 0.07629f
C8295 XThC.Tn[13].t3 VGND 0.02513f
C8296 XThC.Tn[13].t2 VGND 0.02513f
C8297 XThC.Tn[13].n58 VGND 0.05585f
C8298 XThC.Tn[13].n59 VGND 0.24859f
C8299 XThC.Tn[12].t1 VGND 0.01637f
C8300 XThC.Tn[12].t0 VGND 0.01637f
C8301 XThC.Tn[12].n0 VGND 0.03274f
C8302 XThC.Tn[12].t3 VGND 0.01637f
C8303 XThC.Tn[12].t2 VGND 0.01637f
C8304 XThC.Tn[12].n1 VGND 0.04083f
C8305 XThC.Tn[12].n2 VGND 0.08236f
C8306 XThC.Tn[12].t5 VGND 0.02519f
C8307 XThC.Tn[12].t6 VGND 0.02519f
C8308 XThC.Tn[12].n3 VGND 0.05442f
C8309 XThC.Tn[12].t4 VGND 0.02519f
C8310 XThC.Tn[12].t7 VGND 0.02519f
C8311 XThC.Tn[12].n4 VGND 0.08282f
C8312 XThC.Tn[12].n5 VGND 0.23013f
C8313 XThC.Tn[12].t9 VGND 0.02519f
C8314 XThC.Tn[12].t8 VGND 0.02519f
C8315 XThC.Tn[12].n6 VGND 0.07647f
C8316 XThC.Tn[12].t11 VGND 0.02519f
C8317 XThC.Tn[12].t10 VGND 0.02519f
C8318 XThC.Tn[12].n7 VGND 0.05599f
C8319 XThC.Tn[12].n8 VGND 0.24918f
C8320 XThC.Tn[12].n9 VGND 0.03618f
C8321 XThC.Tn[12].t37 VGND 0.01996f
C8322 XThC.Tn[12].t35 VGND 0.0218f
C8323 XThC.Tn[12].n10 VGND 0.04869f
C8324 XThC.Tn[12].n11 VGND 0.02783f
C8325 XThC.Tn[12].n12 VGND 0.03384f
C8326 XThC.Tn[12].t23 VGND 0.01996f
C8327 XThC.Tn[12].t20 VGND 0.0218f
C8328 XThC.Tn[12].n13 VGND 0.04869f
C8329 XThC.Tn[12].n14 VGND 0.02783f
C8330 XThC.Tn[12].n15 VGND 0.16078f
C8331 XThC.Tn[12].t28 VGND 0.01996f
C8332 XThC.Tn[12].t22 VGND 0.0218f
C8333 XThC.Tn[12].n16 VGND 0.04869f
C8334 XThC.Tn[12].n17 VGND 0.02783f
C8335 XThC.Tn[12].n18 VGND 0.16078f
C8336 XThC.Tn[12].t29 VGND 0.01996f
C8337 XThC.Tn[12].t24 VGND 0.0218f
C8338 XThC.Tn[12].n19 VGND 0.04869f
C8339 XThC.Tn[12].n20 VGND 0.02783f
C8340 XThC.Tn[12].n21 VGND 0.16078f
C8341 XThC.Tn[12].t16 VGND 0.01996f
C8342 XThC.Tn[12].t13 VGND 0.0218f
C8343 XThC.Tn[12].n22 VGND 0.04869f
C8344 XThC.Tn[12].n23 VGND 0.02783f
C8345 XThC.Tn[12].n24 VGND 0.16078f
C8346 XThC.Tn[12].t17 VGND 0.01996f
C8347 XThC.Tn[12].t14 VGND 0.0218f
C8348 XThC.Tn[12].n25 VGND 0.04869f
C8349 XThC.Tn[12].n26 VGND 0.02783f
C8350 XThC.Tn[12].n27 VGND 0.16078f
C8351 XThC.Tn[12].t33 VGND 0.01996f
C8352 XThC.Tn[12].t27 VGND 0.0218f
C8353 XThC.Tn[12].n28 VGND 0.04869f
C8354 XThC.Tn[12].n29 VGND 0.02783f
C8355 XThC.Tn[12].n30 VGND 0.16078f
C8356 XThC.Tn[12].t40 VGND 0.01996f
C8357 XThC.Tn[12].t36 VGND 0.0218f
C8358 XThC.Tn[12].n31 VGND 0.04869f
C8359 XThC.Tn[12].n32 VGND 0.02783f
C8360 XThC.Tn[12].n33 VGND 0.16078f
C8361 XThC.Tn[12].t42 VGND 0.01996f
C8362 XThC.Tn[12].t38 VGND 0.0218f
C8363 XThC.Tn[12].n34 VGND 0.04869f
C8364 XThC.Tn[12].n35 VGND 0.02783f
C8365 XThC.Tn[12].n36 VGND 0.16078f
C8366 XThC.Tn[12].t30 VGND 0.01996f
C8367 XThC.Tn[12].t25 VGND 0.0218f
C8368 XThC.Tn[12].n37 VGND 0.04869f
C8369 XThC.Tn[12].n38 VGND 0.02783f
C8370 XThC.Tn[12].n39 VGND 0.16078f
C8371 XThC.Tn[12].t32 VGND 0.01996f
C8372 XThC.Tn[12].t26 VGND 0.0218f
C8373 XThC.Tn[12].n40 VGND 0.04869f
C8374 XThC.Tn[12].n41 VGND 0.02783f
C8375 XThC.Tn[12].n42 VGND 0.16078f
C8376 XThC.Tn[12].t43 VGND 0.01996f
C8377 XThC.Tn[12].t39 VGND 0.0218f
C8378 XThC.Tn[12].n43 VGND 0.04869f
C8379 XThC.Tn[12].n44 VGND 0.02783f
C8380 XThC.Tn[12].n45 VGND 0.16078f
C8381 XThC.Tn[12].t19 VGND 0.01996f
C8382 XThC.Tn[12].t15 VGND 0.0218f
C8383 XThC.Tn[12].n46 VGND 0.04869f
C8384 XThC.Tn[12].n47 VGND 0.02783f
C8385 XThC.Tn[12].n48 VGND 0.16078f
C8386 XThC.Tn[12].t21 VGND 0.01996f
C8387 XThC.Tn[12].t18 VGND 0.0218f
C8388 XThC.Tn[12].n49 VGND 0.04869f
C8389 XThC.Tn[12].n50 VGND 0.02783f
C8390 XThC.Tn[12].n51 VGND 0.16078f
C8391 XThC.Tn[12].t34 VGND 0.01996f
C8392 XThC.Tn[12].t31 VGND 0.0218f
C8393 XThC.Tn[12].n52 VGND 0.04869f
C8394 XThC.Tn[12].n53 VGND 0.02783f
C8395 XThC.Tn[12].n54 VGND 0.16078f
C8396 XThC.Tn[12].t12 VGND 0.01996f
C8397 XThC.Tn[12].t41 VGND 0.0218f
C8398 XThC.Tn[12].n55 VGND 0.04869f
C8399 XThC.Tn[12].n56 VGND 0.02783f
C8400 XThC.Tn[12].n57 VGND 0.16078f
C8401 XThC.Tn[12].n58 VGND 0.88122f
C8402 XThC.Tn[12].n59 VGND 0.0612f
C8403 XThC.Tn[11].t6 VGND 0.01667f
C8404 XThC.Tn[11].t9 VGND 0.01667f
C8405 XThC.Tn[11].n0 VGND 0.04157f
C8406 XThC.Tn[11].t4 VGND 0.01667f
C8407 XThC.Tn[11].t10 VGND 0.01667f
C8408 XThC.Tn[11].n1 VGND 0.03334f
C8409 XThC.Tn[11].n2 VGND 0.07687f
C8410 XThC.Tn[11].t20 VGND 0.02032f
C8411 XThC.Tn[11].t18 VGND 0.0222f
C8412 XThC.Tn[11].n3 VGND 0.04958f
C8413 XThC.Tn[11].n4 VGND 0.02833f
C8414 XThC.Tn[11].n5 VGND 0.03446f
C8415 XThC.Tn[11].t38 VGND 0.02032f
C8416 XThC.Tn[11].t35 VGND 0.0222f
C8417 XThC.Tn[11].n6 VGND 0.04958f
C8418 XThC.Tn[11].n7 VGND 0.02833f
C8419 XThC.Tn[11].n8 VGND 0.1637f
C8420 XThC.Tn[11].t43 VGND 0.02032f
C8421 XThC.Tn[11].t37 VGND 0.0222f
C8422 XThC.Tn[11].n9 VGND 0.04958f
C8423 XThC.Tn[11].n10 VGND 0.02833f
C8424 XThC.Tn[11].n11 VGND 0.1637f
C8425 XThC.Tn[11].t12 VGND 0.02032f
C8426 XThC.Tn[11].t39 VGND 0.0222f
C8427 XThC.Tn[11].n12 VGND 0.04958f
C8428 XThC.Tn[11].n13 VGND 0.02833f
C8429 XThC.Tn[11].n14 VGND 0.1637f
C8430 XThC.Tn[11].t31 VGND 0.02032f
C8431 XThC.Tn[11].t28 VGND 0.0222f
C8432 XThC.Tn[11].n15 VGND 0.04958f
C8433 XThC.Tn[11].n16 VGND 0.02833f
C8434 XThC.Tn[11].n17 VGND 0.1637f
C8435 XThC.Tn[11].t32 VGND 0.02032f
C8436 XThC.Tn[11].t29 VGND 0.0222f
C8437 XThC.Tn[11].n18 VGND 0.04958f
C8438 XThC.Tn[11].n19 VGND 0.02833f
C8439 XThC.Tn[11].n20 VGND 0.1637f
C8440 XThC.Tn[11].t16 VGND 0.02032f
C8441 XThC.Tn[11].t42 VGND 0.0222f
C8442 XThC.Tn[11].n21 VGND 0.04958f
C8443 XThC.Tn[11].n22 VGND 0.02833f
C8444 XThC.Tn[11].n23 VGND 0.1637f
C8445 XThC.Tn[11].t23 VGND 0.02032f
C8446 XThC.Tn[11].t19 VGND 0.0222f
C8447 XThC.Tn[11].n24 VGND 0.04958f
C8448 XThC.Tn[11].n25 VGND 0.02833f
C8449 XThC.Tn[11].n26 VGND 0.1637f
C8450 XThC.Tn[11].t25 VGND 0.02032f
C8451 XThC.Tn[11].t21 VGND 0.0222f
C8452 XThC.Tn[11].n27 VGND 0.04958f
C8453 XThC.Tn[11].n28 VGND 0.02833f
C8454 XThC.Tn[11].n29 VGND 0.1637f
C8455 XThC.Tn[11].t13 VGND 0.02032f
C8456 XThC.Tn[11].t40 VGND 0.0222f
C8457 XThC.Tn[11].n30 VGND 0.04958f
C8458 XThC.Tn[11].n31 VGND 0.02833f
C8459 XThC.Tn[11].n32 VGND 0.1637f
C8460 XThC.Tn[11].t15 VGND 0.02032f
C8461 XThC.Tn[11].t41 VGND 0.0222f
C8462 XThC.Tn[11].n33 VGND 0.04958f
C8463 XThC.Tn[11].n34 VGND 0.02833f
C8464 XThC.Tn[11].n35 VGND 0.1637f
C8465 XThC.Tn[11].t26 VGND 0.02032f
C8466 XThC.Tn[11].t22 VGND 0.0222f
C8467 XThC.Tn[11].n36 VGND 0.04958f
C8468 XThC.Tn[11].n37 VGND 0.02833f
C8469 XThC.Tn[11].n38 VGND 0.1637f
C8470 XThC.Tn[11].t34 VGND 0.02032f
C8471 XThC.Tn[11].t30 VGND 0.0222f
C8472 XThC.Tn[11].n39 VGND 0.04958f
C8473 XThC.Tn[11].n40 VGND 0.02833f
C8474 XThC.Tn[11].n41 VGND 0.1637f
C8475 XThC.Tn[11].t36 VGND 0.02032f
C8476 XThC.Tn[11].t33 VGND 0.0222f
C8477 XThC.Tn[11].n42 VGND 0.04958f
C8478 XThC.Tn[11].n43 VGND 0.02833f
C8479 XThC.Tn[11].n44 VGND 0.1637f
C8480 XThC.Tn[11].t17 VGND 0.02032f
C8481 XThC.Tn[11].t14 VGND 0.0222f
C8482 XThC.Tn[11].n45 VGND 0.04958f
C8483 XThC.Tn[11].n46 VGND 0.02833f
C8484 XThC.Tn[11].n47 VGND 0.1637f
C8485 XThC.Tn[11].t27 VGND 0.02032f
C8486 XThC.Tn[11].t24 VGND 0.0222f
C8487 XThC.Tn[11].n48 VGND 0.04958f
C8488 XThC.Tn[11].n49 VGND 0.02833f
C8489 XThC.Tn[11].n50 VGND 0.1637f
C8490 XThC.Tn[11].n51 VGND 0.07482f
C8491 XThC.Tn[11].t11 VGND 0.02564f
C8492 XThC.Tn[11].t8 VGND 0.02564f
C8493 XThC.Tn[11].n52 VGND 0.0554f
C8494 XThC.Tn[11].t5 VGND 0.02564f
C8495 XThC.Tn[11].t7 VGND 0.02564f
C8496 XThC.Tn[11].n53 VGND 0.08733f
C8497 XThC.Tn[11].n54 VGND 0.23129f
C8498 XThC.Tn[11].n55 VGND 0.01703f
C8499 XThC.Tn[11].t2 VGND 0.02564f
C8500 XThC.Tn[11].t1 VGND 0.02564f
C8501 XThC.Tn[11].n56 VGND 0.057f
C8502 XThC.Tn[11].t0 VGND 0.02564f
C8503 XThC.Tn[11].t3 VGND 0.02564f
C8504 XThC.Tn[11].n57 VGND 0.07786f
C8505 XThC.Tn[11].n58 VGND 0.2537f
C8506 XThC.Tn[9].t4 VGND 0.02612f
C8507 XThC.Tn[9].t7 VGND 0.02612f
C8508 XThC.Tn[9].n0 VGND 0.05643f
C8509 XThC.Tn[9].t6 VGND 0.02612f
C8510 XThC.Tn[9].t5 VGND 0.02612f
C8511 XThC.Tn[9].n1 VGND 0.08894f
C8512 XThC.Tn[9].n2 VGND 0.23556f
C8513 XThC.Tn[9].t9 VGND 0.02612f
C8514 XThC.Tn[9].t8 VGND 0.02612f
C8515 XThC.Tn[9].n3 VGND 0.0793f
C8516 XThC.Tn[9].t11 VGND 0.02612f
C8517 XThC.Tn[9].t10 VGND 0.02612f
C8518 XThC.Tn[9].n4 VGND 0.05805f
C8519 XThC.Tn[9].n5 VGND 0.25838f
C8520 XThC.Tn[9].n6 VGND 0.01734f
C8521 XThC.Tn[9].t26 VGND 0.0207f
C8522 XThC.Tn[9].t12 VGND 0.02261f
C8523 XThC.Tn[9].n7 VGND 0.05049f
C8524 XThC.Tn[9].n8 VGND 0.02885f
C8525 XThC.Tn[9].n9 VGND 0.03509f
C8526 XThC.Tn[9].t13 VGND 0.0207f
C8527 XThC.Tn[9].t30 VGND 0.02261f
C8528 XThC.Tn[9].n10 VGND 0.05049f
C8529 XThC.Tn[9].n11 VGND 0.02885f
C8530 XThC.Tn[9].n12 VGND 0.16672f
C8531 XThC.Tn[9].t15 VGND 0.0207f
C8532 XThC.Tn[9].t34 VGND 0.02261f
C8533 XThC.Tn[9].n13 VGND 0.05049f
C8534 XThC.Tn[9].n14 VGND 0.02885f
C8535 XThC.Tn[9].n15 VGND 0.16672f
C8536 XThC.Tn[9].t17 VGND 0.0207f
C8537 XThC.Tn[9].t35 VGND 0.02261f
C8538 XThC.Tn[9].n16 VGND 0.05049f
C8539 XThC.Tn[9].n17 VGND 0.02885f
C8540 XThC.Tn[9].n18 VGND 0.16672f
C8541 XThC.Tn[9].t39 VGND 0.0207f
C8542 XThC.Tn[9].t24 VGND 0.02261f
C8543 XThC.Tn[9].n19 VGND 0.05049f
C8544 XThC.Tn[9].n20 VGND 0.02885f
C8545 XThC.Tn[9].n21 VGND 0.16672f
C8546 XThC.Tn[9].t40 VGND 0.0207f
C8547 XThC.Tn[9].t25 VGND 0.02261f
C8548 XThC.Tn[9].n22 VGND 0.05049f
C8549 XThC.Tn[9].n23 VGND 0.02885f
C8550 XThC.Tn[9].n24 VGND 0.16672f
C8551 XThC.Tn[9].t22 VGND 0.0207f
C8552 XThC.Tn[9].t38 VGND 0.02261f
C8553 XThC.Tn[9].n25 VGND 0.05049f
C8554 XThC.Tn[9].n26 VGND 0.02885f
C8555 XThC.Tn[9].n27 VGND 0.16672f
C8556 XThC.Tn[9].t28 VGND 0.0207f
C8557 XThC.Tn[9].t14 VGND 0.02261f
C8558 XThC.Tn[9].n28 VGND 0.05049f
C8559 XThC.Tn[9].n29 VGND 0.02885f
C8560 XThC.Tn[9].n30 VGND 0.16672f
C8561 XThC.Tn[9].t31 VGND 0.0207f
C8562 XThC.Tn[9].t16 VGND 0.02261f
C8563 XThC.Tn[9].n31 VGND 0.05049f
C8564 XThC.Tn[9].n32 VGND 0.02885f
C8565 XThC.Tn[9].n33 VGND 0.16672f
C8566 XThC.Tn[9].t19 VGND 0.0207f
C8567 XThC.Tn[9].t36 VGND 0.02261f
C8568 XThC.Tn[9].n34 VGND 0.05049f
C8569 XThC.Tn[9].n35 VGND 0.02885f
C8570 XThC.Tn[9].n36 VGND 0.16672f
C8571 XThC.Tn[9].t21 VGND 0.0207f
C8572 XThC.Tn[9].t37 VGND 0.02261f
C8573 XThC.Tn[9].n37 VGND 0.05049f
C8574 XThC.Tn[9].n38 VGND 0.02885f
C8575 XThC.Tn[9].n39 VGND 0.16672f
C8576 XThC.Tn[9].t32 VGND 0.0207f
C8577 XThC.Tn[9].t18 VGND 0.02261f
C8578 XThC.Tn[9].n40 VGND 0.05049f
C8579 XThC.Tn[9].n41 VGND 0.02885f
C8580 XThC.Tn[9].n42 VGND 0.16672f
C8581 XThC.Tn[9].t42 VGND 0.0207f
C8582 XThC.Tn[9].t27 VGND 0.02261f
C8583 XThC.Tn[9].n43 VGND 0.05049f
C8584 XThC.Tn[9].n44 VGND 0.02885f
C8585 XThC.Tn[9].n45 VGND 0.16672f
C8586 XThC.Tn[9].t43 VGND 0.0207f
C8587 XThC.Tn[9].t29 VGND 0.02261f
C8588 XThC.Tn[9].n46 VGND 0.05049f
C8589 XThC.Tn[9].n47 VGND 0.02885f
C8590 XThC.Tn[9].n48 VGND 0.16672f
C8591 XThC.Tn[9].t23 VGND 0.0207f
C8592 XThC.Tn[9].t41 VGND 0.02261f
C8593 XThC.Tn[9].n49 VGND 0.05049f
C8594 XThC.Tn[9].n50 VGND 0.02885f
C8595 XThC.Tn[9].n51 VGND 0.16672f
C8596 XThC.Tn[9].t33 VGND 0.0207f
C8597 XThC.Tn[9].t20 VGND 0.02261f
C8598 XThC.Tn[9].n52 VGND 0.05049f
C8599 XThC.Tn[9].n53 VGND 0.02885f
C8600 XThC.Tn[9].n54 VGND 0.16672f
C8601 XThC.Tn[9].n55 VGND 0.0762f
C8602 XThC.Tn[9].t1 VGND 0.01698f
C8603 XThC.Tn[9].t0 VGND 0.01698f
C8604 XThC.Tn[9].n56 VGND 0.04234f
C8605 XThC.Tn[9].t2 VGND 0.01698f
C8606 XThC.Tn[9].t3 VGND 0.01698f
C8607 XThC.Tn[9].n57 VGND 0.03395f
C8608 XThC.Tn[9].n58 VGND 0.07828f
C8609 XThC.Tn[5].t7 VGND 0.02353f
C8610 XThC.Tn[5].t6 VGND 0.02353f
C8611 XThC.Tn[5].n0 VGND 0.04749f
C8612 XThC.Tn[5].t5 VGND 0.02353f
C8613 XThC.Tn[5].t4 VGND 0.02353f
C8614 XThC.Tn[5].n1 VGND 0.05557f
C8615 XThC.Tn[5].n2 VGND 0.16669f
C8616 XThC.Tn[5].t1 VGND 0.01529f
C8617 XThC.Tn[5].t0 VGND 0.01529f
C8618 XThC.Tn[5].n3 VGND 0.03483f
C8619 XThC.Tn[5].t8 VGND 0.01529f
C8620 XThC.Tn[5].t11 VGND 0.01529f
C8621 XThC.Tn[5].n4 VGND 0.05803f
C8622 XThC.Tn[5].t10 VGND 0.01529f
C8623 XThC.Tn[5].t9 VGND 0.01529f
C8624 XThC.Tn[5].n5 VGND 0.03483f
C8625 XThC.Tn[5].n6 VGND 0.16586f
C8626 XThC.Tn[5].t3 VGND 0.01529f
C8627 XThC.Tn[5].t2 VGND 0.01529f
C8628 XThC.Tn[5].n7 VGND 0.03483f
C8629 XThC.Tn[5].n8 VGND 0.10253f
C8630 XThC.Tn[5].n9 VGND 0.11572f
C8631 XThC.Tn[5].t15 VGND 0.01865f
C8632 XThC.Tn[5].t33 VGND 0.02037f
C8633 XThC.Tn[5].n10 VGND 0.04549f
C8634 XThC.Tn[5].n11 VGND 0.026f
C8635 XThC.Tn[5].n12 VGND 0.03162f
C8636 XThC.Tn[5].t34 VGND 0.01865f
C8637 XThC.Tn[5].t19 VGND 0.02037f
C8638 XThC.Tn[5].n13 VGND 0.04549f
C8639 XThC.Tn[5].n14 VGND 0.026f
C8640 XThC.Tn[5].n15 VGND 0.15021f
C8641 XThC.Tn[5].t36 VGND 0.01865f
C8642 XThC.Tn[5].t23 VGND 0.02037f
C8643 XThC.Tn[5].n16 VGND 0.04549f
C8644 XThC.Tn[5].n17 VGND 0.026f
C8645 XThC.Tn[5].n18 VGND 0.15021f
C8646 XThC.Tn[5].t38 VGND 0.01865f
C8647 XThC.Tn[5].t24 VGND 0.02037f
C8648 XThC.Tn[5].n19 VGND 0.04549f
C8649 XThC.Tn[5].n20 VGND 0.026f
C8650 XThC.Tn[5].n21 VGND 0.15021f
C8651 XThC.Tn[5].t28 VGND 0.01865f
C8652 XThC.Tn[5].t13 VGND 0.02037f
C8653 XThC.Tn[5].n22 VGND 0.04549f
C8654 XThC.Tn[5].n23 VGND 0.026f
C8655 XThC.Tn[5].n24 VGND 0.15021f
C8656 XThC.Tn[5].t29 VGND 0.01865f
C8657 XThC.Tn[5].t14 VGND 0.02037f
C8658 XThC.Tn[5].n25 VGND 0.04549f
C8659 XThC.Tn[5].n26 VGND 0.026f
C8660 XThC.Tn[5].n27 VGND 0.15021f
C8661 XThC.Tn[5].t43 VGND 0.01865f
C8662 XThC.Tn[5].t27 VGND 0.02037f
C8663 XThC.Tn[5].n28 VGND 0.04549f
C8664 XThC.Tn[5].n29 VGND 0.026f
C8665 XThC.Tn[5].n30 VGND 0.15021f
C8666 XThC.Tn[5].t17 VGND 0.01865f
C8667 XThC.Tn[5].t35 VGND 0.02037f
C8668 XThC.Tn[5].n31 VGND 0.04549f
C8669 XThC.Tn[5].n32 VGND 0.026f
C8670 XThC.Tn[5].n33 VGND 0.15021f
C8671 XThC.Tn[5].t20 VGND 0.01865f
C8672 XThC.Tn[5].t37 VGND 0.02037f
C8673 XThC.Tn[5].n34 VGND 0.04549f
C8674 XThC.Tn[5].n35 VGND 0.026f
C8675 XThC.Tn[5].n36 VGND 0.15021f
C8676 XThC.Tn[5].t40 VGND 0.01865f
C8677 XThC.Tn[5].t25 VGND 0.02037f
C8678 XThC.Tn[5].n37 VGND 0.04549f
C8679 XThC.Tn[5].n38 VGND 0.026f
C8680 XThC.Tn[5].n39 VGND 0.15021f
C8681 XThC.Tn[5].t42 VGND 0.01865f
C8682 XThC.Tn[5].t26 VGND 0.02037f
C8683 XThC.Tn[5].n40 VGND 0.04549f
C8684 XThC.Tn[5].n41 VGND 0.026f
C8685 XThC.Tn[5].n42 VGND 0.15021f
C8686 XThC.Tn[5].t21 VGND 0.01865f
C8687 XThC.Tn[5].t39 VGND 0.02037f
C8688 XThC.Tn[5].n43 VGND 0.04549f
C8689 XThC.Tn[5].n44 VGND 0.026f
C8690 XThC.Tn[5].n45 VGND 0.15021f
C8691 XThC.Tn[5].t31 VGND 0.01865f
C8692 XThC.Tn[5].t16 VGND 0.02037f
C8693 XThC.Tn[5].n46 VGND 0.04549f
C8694 XThC.Tn[5].n47 VGND 0.026f
C8695 XThC.Tn[5].n48 VGND 0.15021f
C8696 XThC.Tn[5].t32 VGND 0.01865f
C8697 XThC.Tn[5].t18 VGND 0.02037f
C8698 XThC.Tn[5].n49 VGND 0.04549f
C8699 XThC.Tn[5].n50 VGND 0.026f
C8700 XThC.Tn[5].n51 VGND 0.15021f
C8701 XThC.Tn[5].t12 VGND 0.01865f
C8702 XThC.Tn[5].t30 VGND 0.02037f
C8703 XThC.Tn[5].n52 VGND 0.04549f
C8704 XThC.Tn[5].n53 VGND 0.026f
C8705 XThC.Tn[5].n54 VGND 0.15021f
C8706 XThC.Tn[5].t22 VGND 0.01865f
C8707 XThC.Tn[5].t41 VGND 0.02037f
C8708 XThC.Tn[5].n55 VGND 0.04549f
C8709 XThC.Tn[5].n56 VGND 0.026f
C8710 XThC.Tn[5].n57 VGND 0.15021f
C8711 XThC.Tn[5].n58 VGND 0.42506f
C8712 XThC.Tn[5].n59 VGND 0.07847f
C8713 XThR.Tn[9].t0 VGND 0.0148f
C8714 XThR.Tn[9].t2 VGND 0.0148f
C8715 XThR.Tn[9].n0 VGND 0.02959f
C8716 XThR.Tn[9].t1 VGND 0.0148f
C8717 XThR.Tn[9].t3 VGND 0.0148f
C8718 XThR.Tn[9].n1 VGND 0.0369f
C8719 XThR.Tn[9].n2 VGND 0.07444f
C8720 XThR.Tn[9].t10 VGND 0.02276f
C8721 XThR.Tn[9].t8 VGND 0.02276f
C8722 XThR.Tn[9].n3 VGND 0.06911f
C8723 XThR.Tn[9].t11 VGND 0.02276f
C8724 XThR.Tn[9].t9 VGND 0.02276f
C8725 XThR.Tn[9].n4 VGND 0.0506f
C8726 XThR.Tn[9].n5 VGND 0.23008f
C8727 XThR.Tn[9].t6 VGND 0.02276f
C8728 XThR.Tn[9].t4 VGND 0.02276f
C8729 XThR.Tn[9].n6 VGND 0.04918f
C8730 XThR.Tn[9].t7 VGND 0.02276f
C8731 XThR.Tn[9].t5 VGND 0.02276f
C8732 XThR.Tn[9].n7 VGND 0.07485f
C8733 XThR.Tn[9].n8 VGND 0.20785f
C8734 XThR.Tn[9].n9 VGND 0.02783f
C8735 XThR.Tn[9].t17 VGND 0.01779f
C8736 XThR.Tn[9].t71 VGND 0.01948f
C8737 XThR.Tn[9].n10 VGND 0.04757f
C8738 XThR.Tn[9].n11 VGND 0.07393f
C8739 XThR.Tn[9].t35 VGND 0.01779f
C8740 XThR.Tn[9].t28 VGND 0.01948f
C8741 XThR.Tn[9].n12 VGND 0.04757f
C8742 XThR.Tn[9].t50 VGND 0.01773f
C8743 XThR.Tn[9].t19 VGND 0.01942f
C8744 XThR.Tn[9].n13 VGND 0.04949f
C8745 XThR.Tn[9].n14 VGND 0.03477f
C8746 XThR.Tn[9].n16 VGND 0.11158f
C8747 XThR.Tn[9].t72 VGND 0.01779f
C8748 XThR.Tn[9].t64 VGND 0.01948f
C8749 XThR.Tn[9].n17 VGND 0.04757f
C8750 XThR.Tn[9].t26 VGND 0.01773f
C8751 XThR.Tn[9].t59 VGND 0.01942f
C8752 XThR.Tn[9].n18 VGND 0.04949f
C8753 XThR.Tn[9].n19 VGND 0.03477f
C8754 XThR.Tn[9].n21 VGND 0.11158f
C8755 XThR.Tn[9].t29 VGND 0.01779f
C8756 XThR.Tn[9].t21 VGND 0.01948f
C8757 XThR.Tn[9].n22 VGND 0.04757f
C8758 XThR.Tn[9].t41 VGND 0.01773f
C8759 XThR.Tn[9].t15 VGND 0.01942f
C8760 XThR.Tn[9].n23 VGND 0.04949f
C8761 XThR.Tn[9].n24 VGND 0.03477f
C8762 XThR.Tn[9].n26 VGND 0.11158f
C8763 XThR.Tn[9].t56 VGND 0.01779f
C8764 XThR.Tn[9].t46 VGND 0.01948f
C8765 XThR.Tn[9].n27 VGND 0.04757f
C8766 XThR.Tn[9].t73 VGND 0.01773f
C8767 XThR.Tn[9].t42 VGND 0.01942f
C8768 XThR.Tn[9].n28 VGND 0.04949f
C8769 XThR.Tn[9].n29 VGND 0.03477f
C8770 XThR.Tn[9].n31 VGND 0.11158f
C8771 XThR.Tn[9].t31 VGND 0.01779f
C8772 XThR.Tn[9].t23 VGND 0.01948f
C8773 XThR.Tn[9].n32 VGND 0.04757f
C8774 XThR.Tn[9].t44 VGND 0.01773f
C8775 XThR.Tn[9].t16 VGND 0.01942f
C8776 XThR.Tn[9].n33 VGND 0.04949f
C8777 XThR.Tn[9].n34 VGND 0.03477f
C8778 XThR.Tn[9].n36 VGND 0.11158f
C8779 XThR.Tn[9].t67 VGND 0.01779f
C8780 XThR.Tn[9].t37 VGND 0.01948f
C8781 XThR.Tn[9].n37 VGND 0.04757f
C8782 XThR.Tn[9].t20 VGND 0.01773f
C8783 XThR.Tn[9].t33 VGND 0.01942f
C8784 XThR.Tn[9].n38 VGND 0.04949f
C8785 XThR.Tn[9].n39 VGND 0.03477f
C8786 XThR.Tn[9].n41 VGND 0.11158f
C8787 XThR.Tn[9].t36 VGND 0.01779f
C8788 XThR.Tn[9].t32 VGND 0.01948f
C8789 XThR.Tn[9].n42 VGND 0.04757f
C8790 XThR.Tn[9].t51 VGND 0.01773f
C8791 XThR.Tn[9].t25 VGND 0.01942f
C8792 XThR.Tn[9].n43 VGND 0.04949f
C8793 XThR.Tn[9].n44 VGND 0.03477f
C8794 XThR.Tn[9].n46 VGND 0.11158f
C8795 XThR.Tn[9].t39 VGND 0.01779f
C8796 XThR.Tn[9].t45 VGND 0.01948f
C8797 XThR.Tn[9].n47 VGND 0.04757f
C8798 XThR.Tn[9].t55 VGND 0.01773f
C8799 XThR.Tn[9].t40 VGND 0.01942f
C8800 XThR.Tn[9].n48 VGND 0.04949f
C8801 XThR.Tn[9].n49 VGND 0.03477f
C8802 XThR.Tn[9].n51 VGND 0.11158f
C8803 XThR.Tn[9].t58 VGND 0.01779f
C8804 XThR.Tn[9].t66 VGND 0.01948f
C8805 XThR.Tn[9].n52 VGND 0.04757f
C8806 XThR.Tn[9].t13 VGND 0.01773f
C8807 XThR.Tn[9].t60 VGND 0.01942f
C8808 XThR.Tn[9].n53 VGND 0.04949f
C8809 XThR.Tn[9].n54 VGND 0.03477f
C8810 XThR.Tn[9].n56 VGND 0.11158f
C8811 XThR.Tn[9].t48 VGND 0.01779f
C8812 XThR.Tn[9].t24 VGND 0.01948f
C8813 XThR.Tn[9].n57 VGND 0.04757f
C8814 XThR.Tn[9].t65 VGND 0.01773f
C8815 XThR.Tn[9].t18 VGND 0.01942f
C8816 XThR.Tn[9].n58 VGND 0.04949f
C8817 XThR.Tn[9].n59 VGND 0.03477f
C8818 XThR.Tn[9].n61 VGND 0.11158f
C8819 XThR.Tn[9].t70 VGND 0.01779f
C8820 XThR.Tn[9].t62 VGND 0.01948f
C8821 XThR.Tn[9].n62 VGND 0.04757f
C8822 XThR.Tn[9].t22 VGND 0.01773f
C8823 XThR.Tn[9].t52 VGND 0.01942f
C8824 XThR.Tn[9].n63 VGND 0.04949f
C8825 XThR.Tn[9].n64 VGND 0.03477f
C8826 XThR.Tn[9].n66 VGND 0.11158f
C8827 XThR.Tn[9].t38 VGND 0.01779f
C8828 XThR.Tn[9].t34 VGND 0.01948f
C8829 XThR.Tn[9].n67 VGND 0.04757f
C8830 XThR.Tn[9].t53 VGND 0.01773f
C8831 XThR.Tn[9].t27 VGND 0.01942f
C8832 XThR.Tn[9].n68 VGND 0.04949f
C8833 XThR.Tn[9].n69 VGND 0.03477f
C8834 XThR.Tn[9].n71 VGND 0.11158f
C8835 XThR.Tn[9].t57 VGND 0.01779f
C8836 XThR.Tn[9].t47 VGND 0.01948f
C8837 XThR.Tn[9].n72 VGND 0.04757f
C8838 XThR.Tn[9].t12 VGND 0.01773f
C8839 XThR.Tn[9].t43 VGND 0.01942f
C8840 XThR.Tn[9].n73 VGND 0.04949f
C8841 XThR.Tn[9].n74 VGND 0.03477f
C8842 XThR.Tn[9].n76 VGND 0.11158f
C8843 XThR.Tn[9].t14 VGND 0.01779f
C8844 XThR.Tn[9].t69 VGND 0.01948f
C8845 XThR.Tn[9].n77 VGND 0.04757f
C8846 XThR.Tn[9].t30 VGND 0.01773f
C8847 XThR.Tn[9].t61 VGND 0.01942f
C8848 XThR.Tn[9].n78 VGND 0.04949f
C8849 XThR.Tn[9].n79 VGND 0.03477f
C8850 XThR.Tn[9].n81 VGND 0.11158f
C8851 XThR.Tn[9].t49 VGND 0.01779f
C8852 XThR.Tn[9].t63 VGND 0.01948f
C8853 XThR.Tn[9].n82 VGND 0.04757f
C8854 XThR.Tn[9].t68 VGND 0.01773f
C8855 XThR.Tn[9].t54 VGND 0.01942f
C8856 XThR.Tn[9].n83 VGND 0.04949f
C8857 XThR.Tn[9].n84 VGND 0.03477f
C8858 XThR.Tn[9].n86 VGND 0.11158f
C8859 XThR.Tn[9].n87 VGND 0.1014f
C8860 XThR.Tn[9].n88 VGND 0.32895f
C8861 XThC.Tn[6].t7 VGND 0.02407f
C8862 XThC.Tn[6].t6 VGND 0.02407f
C8863 XThC.Tn[6].n0 VGND 0.04859f
C8864 XThC.Tn[6].t5 VGND 0.02407f
C8865 XThC.Tn[6].t4 VGND 0.02407f
C8866 XThC.Tn[6].n1 VGND 0.05685f
C8867 XThC.Tn[6].n2 VGND 0.15916f
C8868 XThC.Tn[6].t11 VGND 0.01565f
C8869 XThC.Tn[6].t10 VGND 0.01565f
C8870 XThC.Tn[6].n3 VGND 0.05937f
C8871 XThC.Tn[6].t9 VGND 0.01565f
C8872 XThC.Tn[6].t8 VGND 0.01565f
C8873 XThC.Tn[6].n4 VGND 0.03563f
C8874 XThC.Tn[6].n5 VGND 0.16969f
C8875 XThC.Tn[6].t2 VGND 0.01565f
C8876 XThC.Tn[6].t1 VGND 0.01565f
C8877 XThC.Tn[6].n6 VGND 0.03563f
C8878 XThC.Tn[6].n7 VGND 0.1049f
C8879 XThC.Tn[6].t0 VGND 0.01565f
C8880 XThC.Tn[6].t3 VGND 0.01565f
C8881 XThC.Tn[6].n8 VGND 0.03563f
C8882 XThC.Tn[6].n9 VGND 0.11839f
C8883 XThC.Tn[6].t23 VGND 0.01908f
C8884 XThC.Tn[6].t26 VGND 0.02084f
C8885 XThC.Tn[6].n10 VGND 0.04654f
C8886 XThC.Tn[6].n11 VGND 0.0266f
C8887 XThC.Tn[6].n12 VGND 0.03235f
C8888 XThC.Tn[6].t40 VGND 0.01908f
C8889 XThC.Tn[6].t13 VGND 0.02084f
C8890 XThC.Tn[6].n13 VGND 0.04654f
C8891 XThC.Tn[6].n14 VGND 0.0266f
C8892 XThC.Tn[6].n15 VGND 0.15368f
C8893 XThC.Tn[6].t42 VGND 0.01908f
C8894 XThC.Tn[6].t17 VGND 0.02084f
C8895 XThC.Tn[6].n16 VGND 0.04654f
C8896 XThC.Tn[6].n17 VGND 0.0266f
C8897 XThC.Tn[6].n18 VGND 0.15368f
C8898 XThC.Tn[6].t12 VGND 0.01908f
C8899 XThC.Tn[6].t18 VGND 0.02084f
C8900 XThC.Tn[6].n19 VGND 0.04654f
C8901 XThC.Tn[6].n20 VGND 0.0266f
C8902 XThC.Tn[6].n21 VGND 0.15368f
C8903 XThC.Tn[6].t33 VGND 0.01908f
C8904 XThC.Tn[6].t37 VGND 0.02084f
C8905 XThC.Tn[6].n22 VGND 0.04654f
C8906 XThC.Tn[6].n23 VGND 0.0266f
C8907 XThC.Tn[6].n24 VGND 0.15368f
C8908 XThC.Tn[6].t35 VGND 0.01908f
C8909 XThC.Tn[6].t38 VGND 0.02084f
C8910 XThC.Tn[6].n25 VGND 0.04654f
C8911 XThC.Tn[6].n26 VGND 0.0266f
C8912 XThC.Tn[6].n27 VGND 0.15368f
C8913 XThC.Tn[6].t16 VGND 0.01908f
C8914 XThC.Tn[6].t22 VGND 0.02084f
C8915 XThC.Tn[6].n28 VGND 0.04654f
C8916 XThC.Tn[6].n29 VGND 0.0266f
C8917 XThC.Tn[6].n30 VGND 0.15368f
C8918 XThC.Tn[6].t25 VGND 0.01908f
C8919 XThC.Tn[6].t29 VGND 0.02084f
C8920 XThC.Tn[6].n31 VGND 0.04654f
C8921 XThC.Tn[6].n32 VGND 0.0266f
C8922 XThC.Tn[6].n33 VGND 0.15368f
C8923 XThC.Tn[6].t27 VGND 0.01908f
C8924 XThC.Tn[6].t31 VGND 0.02084f
C8925 XThC.Tn[6].n34 VGND 0.04654f
C8926 XThC.Tn[6].n35 VGND 0.0266f
C8927 XThC.Tn[6].n36 VGND 0.15368f
C8928 XThC.Tn[6].t14 VGND 0.01908f
C8929 XThC.Tn[6].t19 VGND 0.02084f
C8930 XThC.Tn[6].n37 VGND 0.04654f
C8931 XThC.Tn[6].n38 VGND 0.0266f
C8932 XThC.Tn[6].n39 VGND 0.15368f
C8933 XThC.Tn[6].t15 VGND 0.01908f
C8934 XThC.Tn[6].t21 VGND 0.02084f
C8935 XThC.Tn[6].n40 VGND 0.04654f
C8936 XThC.Tn[6].n41 VGND 0.0266f
C8937 XThC.Tn[6].n42 VGND 0.15368f
C8938 XThC.Tn[6].t28 VGND 0.01908f
C8939 XThC.Tn[6].t32 VGND 0.02084f
C8940 XThC.Tn[6].n43 VGND 0.04654f
C8941 XThC.Tn[6].n44 VGND 0.0266f
C8942 XThC.Tn[6].n45 VGND 0.15368f
C8943 XThC.Tn[6].t36 VGND 0.01908f
C8944 XThC.Tn[6].t41 VGND 0.02084f
C8945 XThC.Tn[6].n46 VGND 0.04654f
C8946 XThC.Tn[6].n47 VGND 0.0266f
C8947 XThC.Tn[6].n48 VGND 0.15368f
C8948 XThC.Tn[6].t39 VGND 0.01908f
C8949 XThC.Tn[6].t43 VGND 0.02084f
C8950 XThC.Tn[6].n49 VGND 0.04654f
C8951 XThC.Tn[6].n50 VGND 0.0266f
C8952 XThC.Tn[6].n51 VGND 0.15368f
C8953 XThC.Tn[6].t20 VGND 0.01908f
C8954 XThC.Tn[6].t24 VGND 0.02084f
C8955 XThC.Tn[6].n52 VGND 0.04654f
C8956 XThC.Tn[6].n53 VGND 0.0266f
C8957 XThC.Tn[6].n54 VGND 0.15368f
C8958 XThC.Tn[6].t30 VGND 0.01908f
C8959 XThC.Tn[6].t34 VGND 0.02084f
C8960 XThC.Tn[6].n55 VGND 0.04654f
C8961 XThC.Tn[6].n56 VGND 0.0266f
C8962 XThC.Tn[6].n57 VGND 0.15368f
C8963 XThC.Tn[6].n58 VGND 0.40004f
C8964 XThC.Tn[6].n59 VGND 0.09091f
C8965 XThC.Tn[6].n60 VGND 0.05038f
C8966 XThC.XTBN.Y.n0 VGND 0.01531f
C8967 XThC.XTBN.Y.t50 VGND 0.01024f
C8968 XThC.XTBN.Y.t18 VGND 0.01024f
C8969 XThC.XTBN.Y.n1 VGND 0.01477f
C8970 XThC.XTBN.Y.t120 VGND 0.01024f
C8971 XThC.XTBN.Y.t114 VGND 0.01024f
C8972 XThC.XTBN.Y.n3 VGND 0.0138f
C8973 XThC.XTBN.Y.n5 VGND 0.01477f
C8974 XThC.XTBN.Y.n10 VGND 0.02164f
C8975 XThC.XTBN.Y.t79 VGND 0.01024f
C8976 XThC.XTBN.Y.t36 VGND 0.01024f
C8977 XThC.XTBN.Y.n13 VGND 0.01477f
C8978 XThC.XTBN.Y.t26 VGND 0.01024f
C8979 XThC.XTBN.Y.t21 VGND 0.01024f
C8980 XThC.XTBN.Y.n15 VGND 0.0138f
C8981 XThC.XTBN.Y.n17 VGND 0.01477f
C8982 XThC.XTBN.Y.n22 VGND 0.02164f
C8983 XThC.XTBN.Y.n25 VGND 0.11789f
C8984 XThC.XTBN.Y.t106 VGND 0.01024f
C8985 XThC.XTBN.Y.t70 VGND 0.01024f
C8986 XThC.XTBN.Y.n26 VGND 0.01477f
C8987 XThC.XTBN.Y.t56 VGND 0.01024f
C8988 XThC.XTBN.Y.t48 VGND 0.01024f
C8989 XThC.XTBN.Y.n28 VGND 0.0138f
C8990 XThC.XTBN.Y.n30 VGND 0.01477f
C8991 XThC.XTBN.Y.n35 VGND 0.02164f
C8992 XThC.XTBN.Y.n38 VGND 0.07443f
C8993 XThC.XTBN.Y.t39 VGND 0.01024f
C8994 XThC.XTBN.Y.t122 VGND 0.01024f
C8995 XThC.XTBN.Y.n39 VGND 0.01477f
C8996 XThC.XTBN.Y.t109 VGND 0.01024f
C8997 XThC.XTBN.Y.t102 VGND 0.01024f
C8998 XThC.XTBN.Y.n41 VGND 0.0138f
C8999 XThC.XTBN.Y.n43 VGND 0.01477f
C9000 XThC.XTBN.Y.n48 VGND 0.02164f
C9001 XThC.XTBN.Y.n51 VGND 0.07443f
C9002 XThC.XTBN.Y.t47 VGND 0.01024f
C9003 XThC.XTBN.Y.t17 VGND 0.01024f
C9004 XThC.XTBN.Y.n52 VGND 0.01477f
C9005 XThC.XTBN.Y.t116 VGND 0.01024f
C9006 XThC.XTBN.Y.t111 VGND 0.01024f
C9007 XThC.XTBN.Y.n54 VGND 0.0138f
C9008 XThC.XTBN.Y.n56 VGND 0.01477f
C9009 XThC.XTBN.Y.n61 VGND 0.02164f
C9010 XThC.XTBN.Y.n64 VGND 0.07443f
C9011 XThC.XTBN.Y.t101 VGND 0.01024f
C9012 XThC.XTBN.Y.t63 VGND 0.01024f
C9013 XThC.XTBN.Y.n65 VGND 0.01477f
C9014 XThC.XTBN.Y.t52 VGND 0.01024f
C9015 XThC.XTBN.Y.t44 VGND 0.01024f
C9016 XThC.XTBN.Y.n67 VGND 0.0138f
C9017 XThC.XTBN.Y.n69 VGND 0.01477f
C9018 XThC.XTBN.Y.n74 VGND 0.02164f
C9019 XThC.XTBN.Y.n77 VGND 0.07443f
C9020 XThC.XTBN.Y.t25 VGND 0.01024f
C9021 XThC.XTBN.Y.t100 VGND 0.01024f
C9022 XThC.XTBN.Y.n78 VGND 0.01477f
C9023 XThC.XTBN.Y.t93 VGND 0.01024f
C9024 XThC.XTBN.Y.t90 VGND 0.01024f
C9025 XThC.XTBN.Y.n80 VGND 0.0138f
C9026 XThC.XTBN.Y.n82 VGND 0.01477f
C9027 XThC.XTBN.Y.n87 VGND 0.02164f
C9028 XThC.XTBN.Y.n90 VGND 0.06646f
C9029 XThC.XTBN.Y.t46 VGND 0.01024f
C9030 XThC.XTBN.Y.t6 VGND 0.01024f
C9031 XThC.XTBN.Y.n92 VGND 0.01243f
C9032 XThC.XTBN.Y.t12 VGND 0.01024f
C9033 XThC.XTBN.Y.n93 VGND 0.01348f
C9034 XThC.XTBN.Y.n95 VGND 0.01252f
C9035 XThC.XTBN.Y.n98 VGND 0.01348f
C9036 XThC.XTBN.Y.t54 VGND 0.01024f
C9037 XThC.XTBN.Y.n99 VGND 0.01227f
C9038 XThC.XTBN.Y.n101 VGND 0.01009f
C9039 XThC.XTBN.Y.t38 VGND 0.01024f
C9040 XThC.XTBN.Y.t113 VGND 0.01024f
C9041 XThC.XTBN.Y.n103 VGND 0.01243f
C9042 XThC.XTBN.Y.t119 VGND 0.01024f
C9043 XThC.XTBN.Y.n104 VGND 0.01348f
C9044 XThC.XTBN.Y.n106 VGND 0.01252f
C9045 XThC.XTBN.Y.n109 VGND 0.01348f
C9046 XThC.XTBN.Y.t42 VGND 0.01024f
C9047 XThC.XTBN.Y.n110 VGND 0.01227f
C9048 XThC.XTBN.Y.n113 VGND 0.11256f
C9049 XThC.XTBN.Y.t30 VGND 0.01024f
C9050 XThC.XTBN.Y.t98 VGND 0.01024f
C9051 XThC.XTBN.Y.n115 VGND 0.01243f
C9052 XThC.XTBN.Y.t103 VGND 0.01024f
C9053 XThC.XTBN.Y.n116 VGND 0.01348f
C9054 XThC.XTBN.Y.n118 VGND 0.01252f
C9055 XThC.XTBN.Y.n121 VGND 0.01348f
C9056 XThC.XTBN.Y.t34 VGND 0.01024f
C9057 XThC.XTBN.Y.n122 VGND 0.01227f
C9058 XThC.XTBN.Y.n125 VGND 0.07521f
C9059 XThC.XTBN.Y.t96 VGND 0.01024f
C9060 XThC.XTBN.Y.t51 VGND 0.01024f
C9061 XThC.XTBN.Y.n127 VGND 0.01243f
C9062 XThC.XTBN.Y.t58 VGND 0.01024f
C9063 XThC.XTBN.Y.n128 VGND 0.01348f
C9064 XThC.XTBN.Y.n130 VGND 0.01252f
C9065 XThC.XTBN.Y.n133 VGND 0.01348f
C9066 XThC.XTBN.Y.t99 VGND 0.01024f
C9067 XThC.XTBN.Y.n134 VGND 0.01227f
C9068 XThC.XTBN.Y.n137 VGND 0.07521f
C9069 XThC.XTBN.Y.t88 VGND 0.01024f
C9070 XThC.XTBN.Y.t37 VGND 0.01024f
C9071 XThC.XTBN.Y.n139 VGND 0.01243f
C9072 XThC.XTBN.Y.t40 VGND 0.01024f
C9073 XThC.XTBN.Y.n140 VGND 0.01348f
C9074 XThC.XTBN.Y.n142 VGND 0.01252f
C9075 XThC.XTBN.Y.n145 VGND 0.01348f
C9076 XThC.XTBN.Y.t91 VGND 0.01024f
C9077 XThC.XTBN.Y.n146 VGND 0.01227f
C9078 XThC.XTBN.Y.n149 VGND 0.07534f
C9079 XThC.XTBN.Y.t7 VGND 0.01024f
C9080 XThC.XTBN.Y.t81 VGND 0.01024f
C9081 XThC.XTBN.Y.n151 VGND 0.01243f
C9082 XThC.XTBN.Y.t86 VGND 0.01024f
C9083 XThC.XTBN.Y.n152 VGND 0.01348f
C9084 XThC.XTBN.Y.n154 VGND 0.01252f
C9085 XThC.XTBN.Y.n157 VGND 0.01348f
C9086 XThC.XTBN.Y.t13 VGND 0.01024f
C9087 XThC.XTBN.Y.n158 VGND 0.01227f
C9088 XThC.XTBN.Y.n161 VGND 0.07521f
C9089 XThC.XTBN.Y.t23 VGND 0.01024f
C9090 XThC.XTBN.Y.t95 VGND 0.01024f
C9091 XThC.XTBN.Y.n163 VGND 0.01243f
C9092 XThC.XTBN.Y.t97 VGND 0.01024f
C9093 XThC.XTBN.Y.n164 VGND 0.01348f
C9094 XThC.XTBN.Y.n166 VGND 0.01252f
C9095 XThC.XTBN.Y.n169 VGND 0.01348f
C9096 XThC.XTBN.Y.t28 VGND 0.01024f
C9097 XThC.XTBN.Y.n170 VGND 0.01227f
C9098 XThC.XTBN.Y.n173 VGND 0.08751f
C9099 XThC.XTBN.Y.n174 VGND 0.11019f
C9100 XThC.XTBN.Y.t75 VGND 0.01024f
C9101 XThC.XTBN.Y.t33 VGND 0.01024f
C9102 XThC.XTBN.Y.n175 VGND 0.01477f
C9103 XThC.XTBN.Y.t27 VGND 0.01024f
C9104 XThC.XTBN.Y.n176 VGND 0.02293f
C9105 XThC.XTBN.Y.n181 VGND 0.01477f
C9106 XThC.XTBN.Y.t9 VGND 0.01024f
C9107 XThC.XTBN.Y.n182 VGND 0.0138f
C9108 XThC.XTBN.Y.n186 VGND 0.11129f
C9109 XThC.XTBN.Y.n187 VGND 0.02169f
C9110 XThC.XTBN.Y.n188 VGND 0.01513f
C9111 XThC.XTBN.Y.n189 VGND 0.0307f
C9112 XThR.Tn[12].t0 VGND 0.02276f
C9113 XThR.Tn[12].t2 VGND 0.02276f
C9114 XThR.Tn[12].n0 VGND 0.0506f
C9115 XThR.Tn[12].t3 VGND 0.02276f
C9116 XThR.Tn[12].t1 VGND 0.02276f
C9117 XThR.Tn[12].n1 VGND 0.06912f
C9118 XThR.Tn[12].n2 VGND 0.23009f
C9119 XThR.Tn[12].t7 VGND 0.0148f
C9120 XThR.Tn[12].t5 VGND 0.0148f
C9121 XThR.Tn[12].n3 VGND 0.0369f
C9122 XThR.Tn[12].t6 VGND 0.0148f
C9123 XThR.Tn[12].t4 VGND 0.0148f
C9124 XThR.Tn[12].n4 VGND 0.02959f
C9125 XThR.Tn[12].n5 VGND 0.06824f
C9126 XThR.Tn[12].t36 VGND 0.01779f
C9127 XThR.Tn[12].t28 VGND 0.01948f
C9128 XThR.Tn[12].n6 VGND 0.04757f
C9129 XThR.Tn[12].n7 VGND 0.07393f
C9130 XThR.Tn[12].t53 VGND 0.01779f
C9131 XThR.Tn[12].t43 VGND 0.01948f
C9132 XThR.Tn[12].n8 VGND 0.04757f
C9133 XThR.Tn[12].t71 VGND 0.01773f
C9134 XThR.Tn[12].t21 VGND 0.01942f
C9135 XThR.Tn[12].n9 VGND 0.0495f
C9136 XThR.Tn[12].n10 VGND 0.03477f
C9137 XThR.Tn[12].n12 VGND 0.11159f
C9138 XThR.Tn[12].t30 VGND 0.01779f
C9139 XThR.Tn[12].t20 VGND 0.01948f
C9140 XThR.Tn[12].n13 VGND 0.04757f
C9141 XThR.Tn[12].t49 VGND 0.01773f
C9142 XThR.Tn[12].t60 VGND 0.01942f
C9143 XThR.Tn[12].n14 VGND 0.0495f
C9144 XThR.Tn[12].n15 VGND 0.03477f
C9145 XThR.Tn[12].n17 VGND 0.11159f
C9146 XThR.Tn[12].t45 VGND 0.01779f
C9147 XThR.Tn[12].t38 VGND 0.01948f
C9148 XThR.Tn[12].n18 VGND 0.04757f
C9149 XThR.Tn[12].t63 VGND 0.01773f
C9150 XThR.Tn[12].t15 VGND 0.01942f
C9151 XThR.Tn[12].n19 VGND 0.0495f
C9152 XThR.Tn[12].n20 VGND 0.03477f
C9153 XThR.Tn[12].n22 VGND 0.11159f
C9154 XThR.Tn[12].t70 VGND 0.01779f
C9155 XThR.Tn[12].t66 VGND 0.01948f
C9156 XThR.Tn[12].n23 VGND 0.04757f
C9157 XThR.Tn[12].t33 VGND 0.01773f
C9158 XThR.Tn[12].t46 VGND 0.01942f
C9159 XThR.Tn[12].n24 VGND 0.0495f
C9160 XThR.Tn[12].n25 VGND 0.03477f
C9161 XThR.Tn[12].n27 VGND 0.11159f
C9162 XThR.Tn[12].t48 VGND 0.01779f
C9163 XThR.Tn[12].t39 VGND 0.01948f
C9164 XThR.Tn[12].n28 VGND 0.04757f
C9165 XThR.Tn[12].t64 VGND 0.01773f
C9166 XThR.Tn[12].t17 VGND 0.01942f
C9167 XThR.Tn[12].n29 VGND 0.0495f
C9168 XThR.Tn[12].n30 VGND 0.03477f
C9169 XThR.Tn[12].n32 VGND 0.11159f
C9170 XThR.Tn[12].t23 VGND 0.01779f
C9171 XThR.Tn[12].t56 VGND 0.01948f
C9172 XThR.Tn[12].n33 VGND 0.04757f
C9173 XThR.Tn[12].t41 VGND 0.01773f
C9174 XThR.Tn[12].t37 VGND 0.01942f
C9175 XThR.Tn[12].n34 VGND 0.0495f
C9176 XThR.Tn[12].n35 VGND 0.03477f
C9177 XThR.Tn[12].n37 VGND 0.11159f
C9178 XThR.Tn[12].t54 VGND 0.01779f
C9179 XThR.Tn[12].t51 VGND 0.01948f
C9180 XThR.Tn[12].n38 VGND 0.04757f
C9181 XThR.Tn[12].t72 VGND 0.01773f
C9182 XThR.Tn[12].t29 VGND 0.01942f
C9183 XThR.Tn[12].n39 VGND 0.0495f
C9184 XThR.Tn[12].n40 VGND 0.03477f
C9185 XThR.Tn[12].n42 VGND 0.11159f
C9186 XThR.Tn[12].t59 VGND 0.01779f
C9187 XThR.Tn[12].t65 VGND 0.01948f
C9188 XThR.Tn[12].n43 VGND 0.04757f
C9189 XThR.Tn[12].t14 VGND 0.01773f
C9190 XThR.Tn[12].t44 VGND 0.01942f
C9191 XThR.Tn[12].n44 VGND 0.0495f
C9192 XThR.Tn[12].n45 VGND 0.03477f
C9193 XThR.Tn[12].n47 VGND 0.11159f
C9194 XThR.Tn[12].t12 VGND 0.01779f
C9195 XThR.Tn[12].t22 VGND 0.01948f
C9196 XThR.Tn[12].n48 VGND 0.04757f
C9197 XThR.Tn[12].t35 VGND 0.01773f
C9198 XThR.Tn[12].t61 VGND 0.01942f
C9199 XThR.Tn[12].n49 VGND 0.0495f
C9200 XThR.Tn[12].n50 VGND 0.03477f
C9201 XThR.Tn[12].n52 VGND 0.11159f
C9202 XThR.Tn[12].t68 VGND 0.01779f
C9203 XThR.Tn[12].t40 VGND 0.01948f
C9204 XThR.Tn[12].n53 VGND 0.04757f
C9205 XThR.Tn[12].t26 VGND 0.01773f
C9206 XThR.Tn[12].t19 VGND 0.01942f
C9207 XThR.Tn[12].n54 VGND 0.0495f
C9208 XThR.Tn[12].n55 VGND 0.03477f
C9209 XThR.Tn[12].n57 VGND 0.11159f
C9210 XThR.Tn[12].t25 VGND 0.01779f
C9211 XThR.Tn[12].t16 VGND 0.01948f
C9212 XThR.Tn[12].n58 VGND 0.04757f
C9213 XThR.Tn[12].t42 VGND 0.01773f
C9214 XThR.Tn[12].t55 VGND 0.01942f
C9215 XThR.Tn[12].n59 VGND 0.0495f
C9216 XThR.Tn[12].n60 VGND 0.03477f
C9217 XThR.Tn[12].n62 VGND 0.11159f
C9218 XThR.Tn[12].t57 VGND 0.01779f
C9219 XThR.Tn[12].t52 VGND 0.01948f
C9220 XThR.Tn[12].n63 VGND 0.04757f
C9221 XThR.Tn[12].t13 VGND 0.01773f
C9222 XThR.Tn[12].t31 VGND 0.01942f
C9223 XThR.Tn[12].n64 VGND 0.0495f
C9224 XThR.Tn[12].n65 VGND 0.03477f
C9225 XThR.Tn[12].n67 VGND 0.11159f
C9226 XThR.Tn[12].t73 VGND 0.01779f
C9227 XThR.Tn[12].t67 VGND 0.01948f
C9228 XThR.Tn[12].n68 VGND 0.04757f
C9229 XThR.Tn[12].t34 VGND 0.01773f
C9230 XThR.Tn[12].t47 VGND 0.01942f
C9231 XThR.Tn[12].n69 VGND 0.0495f
C9232 XThR.Tn[12].n70 VGND 0.03477f
C9233 XThR.Tn[12].n72 VGND 0.11159f
C9234 XThR.Tn[12].t32 VGND 0.01779f
C9235 XThR.Tn[12].t24 VGND 0.01948f
C9236 XThR.Tn[12].n73 VGND 0.04757f
C9237 XThR.Tn[12].t50 VGND 0.01773f
C9238 XThR.Tn[12].t62 VGND 0.01942f
C9239 XThR.Tn[12].n74 VGND 0.0495f
C9240 XThR.Tn[12].n75 VGND 0.03477f
C9241 XThR.Tn[12].n77 VGND 0.11159f
C9242 XThR.Tn[12].t69 VGND 0.01779f
C9243 XThR.Tn[12].t18 VGND 0.01948f
C9244 XThR.Tn[12].n78 VGND 0.04757f
C9245 XThR.Tn[12].t27 VGND 0.01773f
C9246 XThR.Tn[12].t58 VGND 0.01942f
C9247 XThR.Tn[12].n79 VGND 0.0495f
C9248 XThR.Tn[12].n80 VGND 0.03477f
C9249 XThR.Tn[12].n82 VGND 0.11159f
C9250 XThR.Tn[12].n83 VGND 0.10141f
C9251 XThR.Tn[12].n84 VGND 0.34586f
C9252 XThR.Tn[12].t10 VGND 0.02276f
C9253 XThR.Tn[12].t8 VGND 0.02276f
C9254 XThR.Tn[12].n85 VGND 0.04918f
C9255 XThR.Tn[12].t11 VGND 0.02276f
C9256 XThR.Tn[12].t9 VGND 0.02276f
C9257 XThR.Tn[12].n86 VGND 0.07486f
C9258 XThR.Tn[12].n87 VGND 0.20785f
C9259 XThR.Tn[12].n88 VGND 0.01024f
C9260 XThR.Tn[14].t8 VGND 0.0231f
C9261 XThR.Tn[14].t9 VGND 0.0231f
C9262 XThR.Tn[14].n0 VGND 0.07015f
C9263 XThR.Tn[14].t10 VGND 0.0231f
C9264 XThR.Tn[14].t11 VGND 0.0231f
C9265 XThR.Tn[14].n1 VGND 0.05136f
C9266 XThR.Tn[14].n2 VGND 0.23353f
C9267 XThR.Tn[14].t6 VGND 0.0231f
C9268 XThR.Tn[14].t7 VGND 0.0231f
C9269 XThR.Tn[14].n3 VGND 0.04992f
C9270 XThR.Tn[14].t4 VGND 0.0231f
C9271 XThR.Tn[14].t5 VGND 0.0231f
C9272 XThR.Tn[14].n4 VGND 0.07598f
C9273 XThR.Tn[14].n5 VGND 0.21096f
C9274 XThR.Tn[14].n6 VGND 0.0104f
C9275 XThR.Tn[14].t69 VGND 0.01806f
C9276 XThR.Tn[14].t62 VGND 0.01977f
C9277 XThR.Tn[14].n7 VGND 0.04828f
C9278 XThR.Tn[14].n8 VGND 0.07503f
C9279 XThR.Tn[14].t24 VGND 0.01806f
C9280 XThR.Tn[14].t13 VGND 0.01977f
C9281 XThR.Tn[14].n9 VGND 0.04828f
C9282 XThR.Tn[14].t28 VGND 0.018f
C9283 XThR.Tn[14].t60 VGND 0.01971f
C9284 XThR.Tn[14].n10 VGND 0.05024f
C9285 XThR.Tn[14].n11 VGND 0.03529f
C9286 XThR.Tn[14].n13 VGND 0.11325f
C9287 XThR.Tn[14].t64 VGND 0.01806f
C9288 XThR.Tn[14].t54 VGND 0.01977f
C9289 XThR.Tn[14].n14 VGND 0.04828f
C9290 XThR.Tn[14].t67 VGND 0.018f
C9291 XThR.Tn[14].t34 VGND 0.01971f
C9292 XThR.Tn[14].n15 VGND 0.05024f
C9293 XThR.Tn[14].n16 VGND 0.03529f
C9294 XThR.Tn[14].n18 VGND 0.11325f
C9295 XThR.Tn[14].t14 VGND 0.01806f
C9296 XThR.Tn[14].t72 VGND 0.01977f
C9297 XThR.Tn[14].n19 VGND 0.04828f
C9298 XThR.Tn[14].t17 VGND 0.018f
C9299 XThR.Tn[14].t52 VGND 0.01971f
C9300 XThR.Tn[14].n20 VGND 0.05024f
C9301 XThR.Tn[14].n21 VGND 0.03529f
C9302 XThR.Tn[14].n23 VGND 0.11325f
C9303 XThR.Tn[14].t44 VGND 0.01806f
C9304 XThR.Tn[14].t38 VGND 0.01977f
C9305 XThR.Tn[14].n24 VGND 0.04828f
C9306 XThR.Tn[14].t47 VGND 0.018f
C9307 XThR.Tn[14].t18 VGND 0.01971f
C9308 XThR.Tn[14].n25 VGND 0.05024f
C9309 XThR.Tn[14].n26 VGND 0.03529f
C9310 XThR.Tn[14].n28 VGND 0.11325f
C9311 XThR.Tn[14].t15 VGND 0.01806f
C9312 XThR.Tn[14].t73 VGND 0.01977f
C9313 XThR.Tn[14].n29 VGND 0.04828f
C9314 XThR.Tn[14].t21 VGND 0.018f
C9315 XThR.Tn[14].t53 VGND 0.01971f
C9316 XThR.Tn[14].n30 VGND 0.05024f
C9317 XThR.Tn[14].n31 VGND 0.03529f
C9318 XThR.Tn[14].n33 VGND 0.11325f
C9319 XThR.Tn[14].t57 VGND 0.01806f
C9320 XThR.Tn[14].t25 VGND 0.01977f
C9321 XThR.Tn[14].n34 VGND 0.04828f
C9322 XThR.Tn[14].t61 VGND 0.018f
C9323 XThR.Tn[14].t71 VGND 0.01971f
C9324 XThR.Tn[14].n35 VGND 0.05024f
C9325 XThR.Tn[14].n36 VGND 0.03529f
C9326 XThR.Tn[14].n38 VGND 0.11325f
C9327 XThR.Tn[14].t23 VGND 0.01806f
C9328 XThR.Tn[14].t19 VGND 0.01977f
C9329 XThR.Tn[14].n39 VGND 0.04828f
C9330 XThR.Tn[14].t29 VGND 0.018f
C9331 XThR.Tn[14].t66 VGND 0.01971f
C9332 XThR.Tn[14].n40 VGND 0.05024f
C9333 XThR.Tn[14].n41 VGND 0.03529f
C9334 XThR.Tn[14].n43 VGND 0.11325f
C9335 XThR.Tn[14].t27 VGND 0.01806f
C9336 XThR.Tn[14].t36 VGND 0.01977f
C9337 XThR.Tn[14].n44 VGND 0.04828f
C9338 XThR.Tn[14].t33 VGND 0.018f
C9339 XThR.Tn[14].t16 VGND 0.01971f
C9340 XThR.Tn[14].n45 VGND 0.05024f
C9341 XThR.Tn[14].n46 VGND 0.03529f
C9342 XThR.Tn[14].n48 VGND 0.11325f
C9343 XThR.Tn[14].t46 VGND 0.01806f
C9344 XThR.Tn[14].t56 VGND 0.01977f
C9345 XThR.Tn[14].n49 VGND 0.04828f
C9346 XThR.Tn[14].t50 VGND 0.018f
C9347 XThR.Tn[14].t35 VGND 0.01971f
C9348 XThR.Tn[14].n50 VGND 0.05024f
C9349 XThR.Tn[14].n51 VGND 0.03529f
C9350 XThR.Tn[14].n53 VGND 0.11325f
C9351 XThR.Tn[14].t40 VGND 0.01806f
C9352 XThR.Tn[14].t12 VGND 0.01977f
C9353 XThR.Tn[14].n54 VGND 0.04828f
C9354 XThR.Tn[14].t42 VGND 0.018f
C9355 XThR.Tn[14].t55 VGND 0.01971f
C9356 XThR.Tn[14].n55 VGND 0.05024f
C9357 XThR.Tn[14].n56 VGND 0.03529f
C9358 XThR.Tn[14].n58 VGND 0.11325f
C9359 XThR.Tn[14].t59 VGND 0.01806f
C9360 XThR.Tn[14].t49 VGND 0.01977f
C9361 XThR.Tn[14].n59 VGND 0.04828f
C9362 XThR.Tn[14].t63 VGND 0.018f
C9363 XThR.Tn[14].t30 VGND 0.01971f
C9364 XThR.Tn[14].n60 VGND 0.05024f
C9365 XThR.Tn[14].n61 VGND 0.03529f
C9366 XThR.Tn[14].n63 VGND 0.11325f
C9367 XThR.Tn[14].t26 VGND 0.01806f
C9368 XThR.Tn[14].t22 VGND 0.01977f
C9369 XThR.Tn[14].n64 VGND 0.04828f
C9370 XThR.Tn[14].t31 VGND 0.018f
C9371 XThR.Tn[14].t68 VGND 0.01971f
C9372 XThR.Tn[14].n65 VGND 0.05024f
C9373 XThR.Tn[14].n66 VGND 0.03529f
C9374 XThR.Tn[14].n68 VGND 0.11325f
C9375 XThR.Tn[14].t45 VGND 0.01806f
C9376 XThR.Tn[14].t39 VGND 0.01977f
C9377 XThR.Tn[14].n69 VGND 0.04828f
C9378 XThR.Tn[14].t48 VGND 0.018f
C9379 XThR.Tn[14].t20 VGND 0.01971f
C9380 XThR.Tn[14].n70 VGND 0.05024f
C9381 XThR.Tn[14].n71 VGND 0.03529f
C9382 XThR.Tn[14].n73 VGND 0.11325f
C9383 XThR.Tn[14].t65 VGND 0.01806f
C9384 XThR.Tn[14].t58 VGND 0.01977f
C9385 XThR.Tn[14].n74 VGND 0.04828f
C9386 XThR.Tn[14].t70 VGND 0.018f
C9387 XThR.Tn[14].t37 VGND 0.01971f
C9388 XThR.Tn[14].n75 VGND 0.05024f
C9389 XThR.Tn[14].n76 VGND 0.03529f
C9390 XThR.Tn[14].n78 VGND 0.11325f
C9391 XThR.Tn[14].t41 VGND 0.01806f
C9392 XThR.Tn[14].t51 VGND 0.01977f
C9393 XThR.Tn[14].n79 VGND 0.04828f
C9394 XThR.Tn[14].t43 VGND 0.018f
C9395 XThR.Tn[14].t32 VGND 0.01971f
C9396 XThR.Tn[14].n80 VGND 0.05024f
C9397 XThR.Tn[14].n81 VGND 0.03529f
C9398 XThR.Tn[14].n83 VGND 0.11325f
C9399 XThR.Tn[14].n84 VGND 0.10292f
C9400 XThR.Tn[14].n85 VGND 0.41345f
C9401 XThR.Tn[14].t0 VGND 0.01502f
C9402 XThR.Tn[14].t1 VGND 0.01502f
C9403 XThR.Tn[14].n86 VGND 0.03003f
C9404 XThR.Tn[14].t2 VGND 0.01502f
C9405 XThR.Tn[14].t3 VGND 0.01502f
C9406 XThR.Tn[14].n87 VGND 0.03745f
C9407 XThR.Tn[14].n88 VGND 0.06926f
C9408 XThR.Tn[6].t7 VGND 0.02178f
C9409 XThR.Tn[6].t4 VGND 0.02178f
C9410 XThR.Tn[6].n0 VGND 0.04396f
C9411 XThR.Tn[6].t6 VGND 0.02178f
C9412 XThR.Tn[6].t5 VGND 0.02178f
C9413 XThR.Tn[6].n1 VGND 0.05143f
C9414 XThR.Tn[6].n2 VGND 0.15428f
C9415 XThR.Tn[6].t8 VGND 0.01416f
C9416 XThR.Tn[6].t9 VGND 0.01416f
C9417 XThR.Tn[6].n3 VGND 0.03223f
C9418 XThR.Tn[6].t11 VGND 0.01416f
C9419 XThR.Tn[6].t10 VGND 0.01416f
C9420 XThR.Tn[6].n4 VGND 0.03223f
C9421 XThR.Tn[6].t0 VGND 0.01416f
C9422 XThR.Tn[6].t1 VGND 0.01416f
C9423 XThR.Tn[6].n5 VGND 0.05371f
C9424 XThR.Tn[6].t3 VGND 0.01416f
C9425 XThR.Tn[6].t2 VGND 0.01416f
C9426 XThR.Tn[6].n6 VGND 0.03223f
C9427 XThR.Tn[6].n7 VGND 0.15351f
C9428 XThR.Tn[6].n8 VGND 0.0949f
C9429 XThR.Tn[6].n9 VGND 0.1071f
C9430 XThR.Tn[6].t62 VGND 0.01702f
C9431 XThR.Tn[6].t56 VGND 0.01864f
C9432 XThR.Tn[6].n10 VGND 0.04551f
C9433 XThR.Tn[6].n11 VGND 0.07073f
C9434 XThR.Tn[6].t20 VGND 0.01702f
C9435 XThR.Tn[6].t72 VGND 0.01864f
C9436 XThR.Tn[6].n12 VGND 0.04551f
C9437 XThR.Tn[6].t36 VGND 0.01696f
C9438 XThR.Tn[6].t68 VGND 0.01858f
C9439 XThR.Tn[6].n13 VGND 0.04735f
C9440 XThR.Tn[6].n14 VGND 0.03327f
C9441 XThR.Tn[6].n16 VGND 0.10675f
C9442 XThR.Tn[6].t57 VGND 0.01702f
C9443 XThR.Tn[6].t49 VGND 0.01864f
C9444 XThR.Tn[6].n17 VGND 0.04551f
C9445 XThR.Tn[6].t14 VGND 0.01696f
C9446 XThR.Tn[6].t45 VGND 0.01858f
C9447 XThR.Tn[6].n18 VGND 0.04735f
C9448 XThR.Tn[6].n19 VGND 0.03327f
C9449 XThR.Tn[6].n21 VGND 0.10675f
C9450 XThR.Tn[6].t73 VGND 0.01702f
C9451 XThR.Tn[6].t66 VGND 0.01864f
C9452 XThR.Tn[6].n22 VGND 0.04551f
C9453 XThR.Tn[6].t26 VGND 0.01696f
C9454 XThR.Tn[6].t63 VGND 0.01858f
C9455 XThR.Tn[6].n23 VGND 0.04735f
C9456 XThR.Tn[6].n24 VGND 0.03327f
C9457 XThR.Tn[6].n26 VGND 0.10675f
C9458 XThR.Tn[6].t35 VGND 0.01702f
C9459 XThR.Tn[6].t31 VGND 0.01864f
C9460 XThR.Tn[6].n27 VGND 0.04551f
C9461 XThR.Tn[6].t59 VGND 0.01696f
C9462 XThR.Tn[6].t27 VGND 0.01858f
C9463 XThR.Tn[6].n28 VGND 0.04735f
C9464 XThR.Tn[6].n29 VGND 0.03327f
C9465 XThR.Tn[6].n31 VGND 0.10675f
C9466 XThR.Tn[6].t13 VGND 0.01702f
C9467 XThR.Tn[6].t67 VGND 0.01864f
C9468 XThR.Tn[6].n32 VGND 0.04551f
C9469 XThR.Tn[6].t29 VGND 0.01696f
C9470 XThR.Tn[6].t64 VGND 0.01858f
C9471 XThR.Tn[6].n33 VGND 0.04735f
C9472 XThR.Tn[6].n34 VGND 0.03327f
C9473 XThR.Tn[6].n36 VGND 0.10675f
C9474 XThR.Tn[6].t51 VGND 0.01702f
C9475 XThR.Tn[6].t22 VGND 0.01864f
C9476 XThR.Tn[6].n37 VGND 0.04551f
C9477 XThR.Tn[6].t70 VGND 0.01696f
C9478 XThR.Tn[6].t19 VGND 0.01858f
C9479 XThR.Tn[6].n38 VGND 0.04735f
C9480 XThR.Tn[6].n39 VGND 0.03327f
C9481 XThR.Tn[6].n41 VGND 0.10675f
C9482 XThR.Tn[6].t21 VGND 0.01702f
C9483 XThR.Tn[6].t17 VGND 0.01864f
C9484 XThR.Tn[6].n42 VGND 0.04551f
C9485 XThR.Tn[6].t37 VGND 0.01696f
C9486 XThR.Tn[6].t12 VGND 0.01858f
C9487 XThR.Tn[6].n43 VGND 0.04735f
C9488 XThR.Tn[6].n44 VGND 0.03327f
C9489 XThR.Tn[6].n46 VGND 0.10675f
C9490 XThR.Tn[6].t24 VGND 0.01702f
C9491 XThR.Tn[6].t30 VGND 0.01864f
C9492 XThR.Tn[6].n47 VGND 0.04551f
C9493 XThR.Tn[6].t43 VGND 0.01696f
C9494 XThR.Tn[6].t25 VGND 0.01858f
C9495 XThR.Tn[6].n48 VGND 0.04735f
C9496 XThR.Tn[6].n49 VGND 0.03327f
C9497 XThR.Tn[6].n51 VGND 0.10675f
C9498 XThR.Tn[6].t40 VGND 0.01702f
C9499 XThR.Tn[6].t50 VGND 0.01864f
C9500 XThR.Tn[6].n52 VGND 0.04551f
C9501 XThR.Tn[6].t61 VGND 0.01696f
C9502 XThR.Tn[6].t47 VGND 0.01858f
C9503 XThR.Tn[6].n53 VGND 0.04735f
C9504 XThR.Tn[6].n54 VGND 0.03327f
C9505 XThR.Tn[6].n56 VGND 0.10675f
C9506 XThR.Tn[6].t33 VGND 0.01702f
C9507 XThR.Tn[6].t69 VGND 0.01864f
C9508 XThR.Tn[6].n57 VGND 0.04551f
C9509 XThR.Tn[6].t54 VGND 0.01696f
C9510 XThR.Tn[6].t65 VGND 0.01858f
C9511 XThR.Tn[6].n58 VGND 0.04735f
C9512 XThR.Tn[6].n59 VGND 0.03327f
C9513 XThR.Tn[6].n61 VGND 0.10675f
C9514 XThR.Tn[6].t53 VGND 0.01702f
C9515 XThR.Tn[6].t44 VGND 0.01864f
C9516 XThR.Tn[6].n62 VGND 0.04551f
C9517 XThR.Tn[6].t71 VGND 0.01696f
C9518 XThR.Tn[6].t39 VGND 0.01858f
C9519 XThR.Tn[6].n63 VGND 0.04735f
C9520 XThR.Tn[6].n64 VGND 0.03327f
C9521 XThR.Tn[6].n66 VGND 0.10675f
C9522 XThR.Tn[6].t23 VGND 0.01702f
C9523 XThR.Tn[6].t18 VGND 0.01864f
C9524 XThR.Tn[6].n67 VGND 0.04551f
C9525 XThR.Tn[6].t41 VGND 0.01696f
C9526 XThR.Tn[6].t15 VGND 0.01858f
C9527 XThR.Tn[6].n68 VGND 0.04735f
C9528 XThR.Tn[6].n69 VGND 0.03327f
C9529 XThR.Tn[6].n71 VGND 0.10675f
C9530 XThR.Tn[6].t38 VGND 0.01702f
C9531 XThR.Tn[6].t32 VGND 0.01864f
C9532 XThR.Tn[6].n72 VGND 0.04551f
C9533 XThR.Tn[6].t60 VGND 0.01696f
C9534 XThR.Tn[6].t28 VGND 0.01858f
C9535 XThR.Tn[6].n73 VGND 0.04735f
C9536 XThR.Tn[6].n74 VGND 0.03327f
C9537 XThR.Tn[6].n76 VGND 0.10675f
C9538 XThR.Tn[6].t58 VGND 0.01702f
C9539 XThR.Tn[6].t52 VGND 0.01864f
C9540 XThR.Tn[6].n77 VGND 0.04551f
C9541 XThR.Tn[6].t16 VGND 0.01696f
C9542 XThR.Tn[6].t48 VGND 0.01858f
C9543 XThR.Tn[6].n78 VGND 0.04735f
C9544 XThR.Tn[6].n79 VGND 0.03327f
C9545 XThR.Tn[6].n81 VGND 0.10675f
C9546 XThR.Tn[6].t34 VGND 0.01702f
C9547 XThR.Tn[6].t46 VGND 0.01864f
C9548 XThR.Tn[6].n82 VGND 0.04551f
C9549 XThR.Tn[6].t55 VGND 0.01696f
C9550 XThR.Tn[6].t42 VGND 0.01858f
C9551 XThR.Tn[6].n83 VGND 0.04735f
C9552 XThR.Tn[6].n84 VGND 0.03327f
C9553 XThR.Tn[6].n86 VGND 0.10675f
C9554 XThR.Tn[6].n87 VGND 0.09701f
C9555 XThR.Tn[6].n88 VGND 0.16149f
C9556 XThR.XTBN.Y.t60 VGND 0.01149f
C9557 XThR.XTBN.Y.n1 VGND 0.01377f
C9558 XThR.XTBN.Y.t12 VGND 0.01149f
C9559 XThR.XTBN.Y.t81 VGND 0.01149f
C9560 XThR.XTBN.Y.n2 VGND 0.01512f
C9561 XThR.XTBN.Y.t121 VGND 0.01149f
C9562 XThR.XTBN.Y.n3 VGND 0.01395f
C9563 XThR.XTBN.Y.n5 VGND 0.01333f
C9564 XThR.XTBN.Y.n8 VGND 0.01512f
C9565 XThR.XTBN.Y.n10 VGND 0.01247f
C9566 XThR.XTBN.Y.t115 VGND 0.01149f
C9567 XThR.XTBN.Y.n12 VGND 0.01377f
C9568 XThR.XTBN.Y.t65 VGND 0.01149f
C9569 XThR.XTBN.Y.t21 VGND 0.01149f
C9570 XThR.XTBN.Y.n13 VGND 0.01512f
C9571 XThR.XTBN.Y.t57 VGND 0.01149f
C9572 XThR.XTBN.Y.n14 VGND 0.01395f
C9573 XThR.XTBN.Y.n16 VGND 0.01333f
C9574 XThR.XTBN.Y.n19 VGND 0.01512f
C9575 XThR.XTBN.Y.n22 VGND 0.12629f
C9576 XThR.XTBN.Y.t27 VGND 0.01149f
C9577 XThR.XTBN.Y.n24 VGND 0.01377f
C9578 XThR.XTBN.Y.t96 VGND 0.01149f
C9579 XThR.XTBN.Y.t46 VGND 0.01149f
C9580 XThR.XTBN.Y.n25 VGND 0.01512f
C9581 XThR.XTBN.Y.t89 VGND 0.01149f
C9582 XThR.XTBN.Y.n26 VGND 0.01395f
C9583 XThR.XTBN.Y.n28 VGND 0.01333f
C9584 XThR.XTBN.Y.n31 VGND 0.01512f
C9585 XThR.XTBN.Y.n34 VGND 0.08438f
C9586 XThR.XTBN.Y.t80 VGND 0.01149f
C9587 XThR.XTBN.Y.n36 VGND 0.01377f
C9588 XThR.XTBN.Y.t31 VGND 0.01149f
C9589 XThR.XTBN.Y.t102 VGND 0.01149f
C9590 XThR.XTBN.Y.n37 VGND 0.01512f
C9591 XThR.XTBN.Y.t25 VGND 0.01149f
C9592 XThR.XTBN.Y.n38 VGND 0.01395f
C9593 XThR.XTBN.Y.n40 VGND 0.01333f
C9594 XThR.XTBN.Y.n43 VGND 0.01512f
C9595 XThR.XTBN.Y.n46 VGND 0.08438f
C9596 XThR.XTBN.Y.t85 VGND 0.01149f
C9597 XThR.XTBN.Y.n48 VGND 0.01377f
C9598 XThR.XTBN.Y.t33 VGND 0.01149f
C9599 XThR.XTBN.Y.t105 VGND 0.01149f
C9600 XThR.XTBN.Y.n49 VGND 0.01512f
C9601 XThR.XTBN.Y.t26 VGND 0.01149f
C9602 XThR.XTBN.Y.n50 VGND 0.01395f
C9603 XThR.XTBN.Y.n52 VGND 0.01333f
C9604 XThR.XTBN.Y.n55 VGND 0.01512f
C9605 XThR.XTBN.Y.n58 VGND 0.08453f
C9606 XThR.XTBN.Y.t54 VGND 0.01149f
C9607 XThR.XTBN.Y.n60 VGND 0.01377f
C9608 XThR.XTBN.Y.t5 VGND 0.01149f
C9609 XThR.XTBN.Y.t73 VGND 0.01149f
C9610 XThR.XTBN.Y.n61 VGND 0.01512f
C9611 XThR.XTBN.Y.t114 VGND 0.01149f
C9612 XThR.XTBN.Y.n62 VGND 0.01395f
C9613 XThR.XTBN.Y.n64 VGND 0.01333f
C9614 XThR.XTBN.Y.n67 VGND 0.01512f
C9615 XThR.XTBN.Y.n70 VGND 0.08438f
C9616 XThR.XTBN.Y.t49 VGND 0.01149f
C9617 XThR.XTBN.Y.n72 VGND 0.01377f
C9618 XThR.XTBN.Y.t119 VGND 0.01149f
C9619 XThR.XTBN.Y.t69 VGND 0.01149f
C9620 XThR.XTBN.Y.n73 VGND 0.01512f
C9621 XThR.XTBN.Y.t108 VGND 0.01149f
C9622 XThR.XTBN.Y.n74 VGND 0.01395f
C9623 XThR.XTBN.Y.n76 VGND 0.01333f
C9624 XThR.XTBN.Y.n79 VGND 0.01512f
C9625 XThR.XTBN.Y.n82 VGND 0.09633f
C9626 XThR.XTBN.Y.t99 VGND 0.01149f
C9627 XThR.XTBN.Y.t87 VGND 0.01149f
C9628 XThR.XTBN.Y.n83 VGND 0.01657f
C9629 XThR.XTBN.Y.t77 VGND 0.01149f
C9630 XThR.XTBN.Y.t68 VGND 0.01149f
C9631 XThR.XTBN.Y.n84 VGND 0.01548f
C9632 XThR.XTBN.Y.n87 VGND 0.01657f
C9633 XThR.XTBN.Y.n92 VGND 0.02428f
C9634 XThR.XTBN.Y.n93 VGND 0.01348f
C9635 XThR.XTBN.Y.t66 VGND 0.01149f
C9636 XThR.XTBN.Y.t23 VGND 0.01149f
C9637 XThR.XTBN.Y.n94 VGND 0.01657f
C9638 XThR.XTBN.Y.t59 VGND 0.01149f
C9639 XThR.XTBN.Y.t97 VGND 0.01149f
C9640 XThR.XTBN.Y.n95 VGND 0.01548f
C9641 XThR.XTBN.Y.n98 VGND 0.01657f
C9642 XThR.XTBN.Y.n103 VGND 0.02428f
C9643 XThR.XTBN.Y.n105 VGND 0.13434f
C9644 XThR.XTBN.Y.t15 VGND 0.01149f
C9645 XThR.XTBN.Y.t83 VGND 0.01149f
C9646 XThR.XTBN.Y.n106 VGND 0.01657f
C9647 XThR.XTBN.Y.t123 VGND 0.01149f
C9648 XThR.XTBN.Y.t39 VGND 0.01149f
C9649 XThR.XTBN.Y.n107 VGND 0.01548f
C9650 XThR.XTBN.Y.n110 VGND 0.01657f
C9651 XThR.XTBN.Y.n115 VGND 0.02428f
C9652 XThR.XTBN.Y.n117 VGND 0.08431f
C9653 XThR.XTBN.Y.t100 VGND 0.01149f
C9654 XThR.XTBN.Y.t50 VGND 0.01149f
C9655 XThR.XTBN.Y.n118 VGND 0.01657f
C9656 XThR.XTBN.Y.t92 VGND 0.01149f
C9657 XThR.XTBN.Y.t13 VGND 0.01149f
C9658 XThR.XTBN.Y.n119 VGND 0.01548f
C9659 XThR.XTBN.Y.n122 VGND 0.01657f
C9660 XThR.XTBN.Y.n127 VGND 0.02428f
C9661 XThR.XTBN.Y.n129 VGND 0.08431f
C9662 XThR.XTBN.Y.t45 VGND 0.01149f
C9663 XThR.XTBN.Y.t117 VGND 0.01149f
C9664 XThR.XTBN.Y.n130 VGND 0.01657f
C9665 XThR.XTBN.Y.t36 VGND 0.01149f
C9666 XThR.XTBN.Y.t75 VGND 0.01149f
C9667 XThR.XTBN.Y.n131 VGND 0.01548f
C9668 XThR.XTBN.Y.n134 VGND 0.01657f
C9669 XThR.XTBN.Y.n139 VGND 0.02428f
C9670 XThR.XTBN.Y.n141 VGND 0.08431f
C9671 XThR.XTBN.Y.t19 VGND 0.01149f
C9672 XThR.XTBN.Y.t86 VGND 0.01149f
C9673 XThR.XTBN.Y.n142 VGND 0.01657f
C9674 XThR.XTBN.Y.t6 VGND 0.01149f
C9675 XThR.XTBN.Y.t43 VGND 0.01149f
C9676 XThR.XTBN.Y.n143 VGND 0.01548f
C9677 XThR.XTBN.Y.n146 VGND 0.01657f
C9678 XThR.XTBN.Y.n151 VGND 0.02428f
C9679 XThR.XTBN.Y.n153 VGND 0.08431f
C9680 XThR.XTBN.Y.t41 VGND 0.01149f
C9681 XThR.XTBN.Y.t113 VGND 0.01149f
C9682 XThR.XTBN.Y.n154 VGND 0.01657f
C9683 XThR.XTBN.Y.t34 VGND 0.01149f
C9684 XThR.XTBN.Y.t72 VGND 0.01149f
C9685 XThR.XTBN.Y.n155 VGND 0.01548f
C9686 XThR.XTBN.Y.n158 VGND 0.01657f
C9687 XThR.XTBN.Y.n163 VGND 0.02428f
C9688 XThR.XTBN.Y.n165 VGND 0.07758f
C9689 XThR.XTBN.Y.n166 VGND 0.12286f
C9690 XThR.XTBN.Y.t106 VGND 0.01149f
C9691 XThR.XTBN.Y.t63 VGND 0.01149f
C9692 XThR.XTBN.Y.n167 VGND 0.01548f
C9693 XThR.XTBN.Y.n169 VGND 0.01657f
C9694 XThR.XTBN.Y.t56 VGND 0.01149f
C9695 XThR.XTBN.Y.t7 VGND 0.01149f
C9696 XThR.XTBN.Y.n170 VGND 0.02573f
C9697 XThR.XTBN.Y.n174 VGND 0.01657f
C9698 XThR.XTBN.Y.n178 VGND 0.12527f
C9699 XThR.XTBN.Y.n179 VGND 0.02292f
C9700 XThR.XTBN.Y.n180 VGND 0.01622f
C9701 XThR.XTBN.Y.n183 VGND 0.01145f
C9702 XThR.XTBN.Y.n184 VGND 0.02249f
C9703 XThC.Tn[10].t2 VGND 0.01671f
C9704 XThC.Tn[10].t6 VGND 0.01671f
C9705 XThC.Tn[10].n0 VGND 0.04168f
C9706 XThC.Tn[10].t10 VGND 0.01671f
C9707 XThC.Tn[10].t3 VGND 0.01671f
C9708 XThC.Tn[10].n1 VGND 0.03342f
C9709 XThC.Tn[10].n2 VGND 0.08408f
C9710 XThC.Tn[10].t38 VGND 0.02038f
C9711 XThC.Tn[10].t36 VGND 0.02226f
C9712 XThC.Tn[10].n3 VGND 0.04971f
C9713 XThC.Tn[10].n4 VGND 0.02841f
C9714 XThC.Tn[10].n5 VGND 0.03455f
C9715 XThC.Tn[10].t24 VGND 0.02038f
C9716 XThC.Tn[10].t21 VGND 0.02226f
C9717 XThC.Tn[10].n6 VGND 0.04971f
C9718 XThC.Tn[10].n7 VGND 0.02841f
C9719 XThC.Tn[10].n8 VGND 0.16413f
C9720 XThC.Tn[10].t29 VGND 0.02038f
C9721 XThC.Tn[10].t23 VGND 0.02226f
C9722 XThC.Tn[10].n9 VGND 0.04971f
C9723 XThC.Tn[10].n10 VGND 0.02841f
C9724 XThC.Tn[10].n11 VGND 0.16413f
C9725 XThC.Tn[10].t30 VGND 0.02038f
C9726 XThC.Tn[10].t25 VGND 0.02226f
C9727 XThC.Tn[10].n12 VGND 0.04971f
C9728 XThC.Tn[10].n13 VGND 0.02841f
C9729 XThC.Tn[10].n14 VGND 0.16413f
C9730 XThC.Tn[10].t17 VGND 0.02038f
C9731 XThC.Tn[10].t14 VGND 0.02226f
C9732 XThC.Tn[10].n15 VGND 0.04971f
C9733 XThC.Tn[10].n16 VGND 0.02841f
C9734 XThC.Tn[10].n17 VGND 0.16413f
C9735 XThC.Tn[10].t18 VGND 0.02038f
C9736 XThC.Tn[10].t15 VGND 0.02226f
C9737 XThC.Tn[10].n18 VGND 0.04971f
C9738 XThC.Tn[10].n19 VGND 0.02841f
C9739 XThC.Tn[10].n20 VGND 0.16413f
C9740 XThC.Tn[10].t34 VGND 0.02038f
C9741 XThC.Tn[10].t28 VGND 0.02226f
C9742 XThC.Tn[10].n21 VGND 0.04971f
C9743 XThC.Tn[10].n22 VGND 0.02841f
C9744 XThC.Tn[10].n23 VGND 0.16413f
C9745 XThC.Tn[10].t41 VGND 0.02038f
C9746 XThC.Tn[10].t37 VGND 0.02226f
C9747 XThC.Tn[10].n24 VGND 0.04971f
C9748 XThC.Tn[10].n25 VGND 0.02841f
C9749 XThC.Tn[10].n26 VGND 0.16413f
C9750 XThC.Tn[10].t43 VGND 0.02038f
C9751 XThC.Tn[10].t39 VGND 0.02226f
C9752 XThC.Tn[10].n27 VGND 0.04971f
C9753 XThC.Tn[10].n28 VGND 0.02841f
C9754 XThC.Tn[10].n29 VGND 0.16413f
C9755 XThC.Tn[10].t31 VGND 0.02038f
C9756 XThC.Tn[10].t26 VGND 0.02226f
C9757 XThC.Tn[10].n30 VGND 0.04971f
C9758 XThC.Tn[10].n31 VGND 0.02841f
C9759 XThC.Tn[10].n32 VGND 0.16413f
C9760 XThC.Tn[10].t33 VGND 0.02038f
C9761 XThC.Tn[10].t27 VGND 0.02226f
C9762 XThC.Tn[10].n33 VGND 0.04971f
C9763 XThC.Tn[10].n34 VGND 0.02841f
C9764 XThC.Tn[10].n35 VGND 0.16413f
C9765 XThC.Tn[10].t12 VGND 0.02038f
C9766 XThC.Tn[10].t40 VGND 0.02226f
C9767 XThC.Tn[10].n36 VGND 0.04971f
C9768 XThC.Tn[10].n37 VGND 0.02841f
C9769 XThC.Tn[10].n38 VGND 0.16413f
C9770 XThC.Tn[10].t20 VGND 0.02038f
C9771 XThC.Tn[10].t16 VGND 0.02226f
C9772 XThC.Tn[10].n39 VGND 0.04971f
C9773 XThC.Tn[10].n40 VGND 0.02841f
C9774 XThC.Tn[10].n41 VGND 0.16413f
C9775 XThC.Tn[10].t22 VGND 0.02038f
C9776 XThC.Tn[10].t19 VGND 0.02226f
C9777 XThC.Tn[10].n42 VGND 0.04971f
C9778 XThC.Tn[10].n43 VGND 0.02841f
C9779 XThC.Tn[10].n44 VGND 0.16413f
C9780 XThC.Tn[10].t35 VGND 0.02038f
C9781 XThC.Tn[10].t32 VGND 0.02226f
C9782 XThC.Tn[10].n45 VGND 0.04971f
C9783 XThC.Tn[10].n46 VGND 0.02841f
C9784 XThC.Tn[10].n47 VGND 0.16413f
C9785 XThC.Tn[10].t13 VGND 0.02038f
C9786 XThC.Tn[10].t42 VGND 0.02226f
C9787 XThC.Tn[10].n48 VGND 0.04971f
C9788 XThC.Tn[10].n49 VGND 0.02841f
C9789 XThC.Tn[10].n50 VGND 0.16413f
C9790 XThC.Tn[10].n51 VGND 0.81978f
C9791 XThC.Tn[10].n52 VGND 0.06249f
C9792 XThC.Tn[10].t5 VGND 0.02571f
C9793 XThC.Tn[10].t4 VGND 0.02571f
C9794 XThC.Tn[10].n53 VGND 0.05555f
C9795 XThC.Tn[10].t7 VGND 0.02571f
C9796 XThC.Tn[10].t0 VGND 0.02571f
C9797 XThC.Tn[10].n54 VGND 0.08455f
C9798 XThC.Tn[10].n55 VGND 0.23493f
C9799 XThC.Tn[10].n56 VGND 0.03694f
C9800 XThC.Tn[10].t1 VGND 0.02571f
C9801 XThC.Tn[10].t8 VGND 0.02571f
C9802 XThC.Tn[10].n57 VGND 0.07807f
C9803 XThC.Tn[10].t11 VGND 0.02571f
C9804 XThC.Tn[10].t9 VGND 0.02571f
C9805 XThC.Tn[10].n58 VGND 0.05715f
C9806 XThC.Tn[10].n59 VGND 0.25438f
C9807 Iout.n0 VGND 0.24452f
C9808 Iout.n1 VGND 1.27854f
C9809 Iout.n2 VGND 0.24452f
C9810 Iout.n3 VGND 0.24452f
C9811 Iout.t170 VGND 0.02354f
C9812 Iout.n4 VGND 0.05236f
C9813 Iout.n5 VGND 0.20684f
C9814 Iout.n6 VGND 0.24452f
C9815 Iout.n7 VGND 1.27854f
C9816 Iout.n8 VGND 0.24452f
C9817 Iout.t92 VGND 0.02354f
C9818 Iout.n9 VGND 0.05236f
C9819 Iout.n10 VGND 0.20684f
C9820 Iout.n11 VGND 0.24452f
C9821 Iout.n12 VGND 1.27854f
C9822 Iout.n13 VGND 0.24452f
C9823 Iout.t14 VGND 0.02354f
C9824 Iout.n14 VGND 0.05236f
C9825 Iout.n15 VGND 0.20684f
C9826 Iout.n16 VGND 0.24452f
C9827 Iout.n17 VGND 1.27854f
C9828 Iout.n18 VGND 0.24452f
C9829 Iout.t6 VGND 0.02354f
C9830 Iout.n19 VGND 0.05236f
C9831 Iout.n20 VGND 0.20684f
C9832 Iout.n21 VGND 0.50694f
C9833 Iout.t116 VGND 0.02354f
C9834 Iout.n22 VGND 0.05236f
C9835 Iout.n23 VGND 0.30503f
C9836 Iout.n24 VGND 0.24452f
C9837 Iout.n25 VGND 0.24452f
C9838 Iout.n26 VGND 0.24452f
C9839 Iout.n27 VGND 0.24452f
C9840 Iout.n28 VGND 0.24452f
C9841 Iout.n29 VGND 0.24452f
C9842 Iout.n30 VGND 0.24452f
C9843 Iout.n31 VGND 0.24452f
C9844 Iout.n32 VGND 0.24452f
C9845 Iout.n33 VGND 0.24452f
C9846 Iout.n34 VGND 0.24452f
C9847 Iout.n35 VGND 0.24452f
C9848 Iout.n36 VGND 0.24452f
C9849 Iout.n37 VGND 0.24452f
C9850 Iout.t112 VGND 0.02354f
C9851 Iout.n38 VGND 0.05236f
C9852 Iout.n39 VGND 0.02663f
C9853 Iout.n40 VGND 0.24452f
C9854 Iout.n41 VGND 0.04879f
C9855 Iout.t196 VGND 0.02354f
C9856 Iout.n42 VGND 0.05236f
C9857 Iout.n43 VGND 0.02663f
C9858 Iout.t120 VGND 0.02354f
C9859 Iout.n44 VGND 0.05236f
C9860 Iout.n45 VGND 0.02663f
C9861 Iout.n46 VGND 0.24452f
C9862 Iout.t36 VGND 0.02354f
C9863 Iout.n47 VGND 0.05236f
C9864 Iout.n48 VGND 0.02663f
C9865 Iout.n49 VGND 0.24452f
C9866 Iout.t202 VGND 0.02354f
C9867 Iout.n50 VGND 0.05236f
C9868 Iout.n51 VGND 0.02663f
C9869 Iout.n52 VGND 0.24452f
C9870 Iout.t227 VGND 0.02354f
C9871 Iout.n53 VGND 0.05236f
C9872 Iout.n54 VGND 0.02663f
C9873 Iout.n55 VGND 0.24452f
C9874 Iout.t100 VGND 0.02354f
C9875 Iout.n56 VGND 0.05236f
C9876 Iout.n57 VGND 0.02663f
C9877 Iout.n58 VGND 0.24452f
C9878 Iout.t57 VGND 0.02354f
C9879 Iout.n59 VGND 0.05236f
C9880 Iout.n60 VGND 0.02663f
C9881 Iout.n61 VGND 0.24452f
C9882 Iout.t119 VGND 0.02354f
C9883 Iout.n62 VGND 0.05236f
C9884 Iout.n63 VGND 0.02663f
C9885 Iout.n64 VGND 0.24452f
C9886 Iout.t109 VGND 0.02354f
C9887 Iout.n65 VGND 0.05236f
C9888 Iout.n66 VGND 0.02663f
C9889 Iout.n67 VGND 0.24452f
C9890 Iout.t61 VGND 0.02354f
C9891 Iout.n68 VGND 0.05236f
C9892 Iout.n69 VGND 0.02663f
C9893 Iout.n70 VGND 0.24452f
C9894 Iout.t38 VGND 0.02354f
C9895 Iout.n71 VGND 0.05236f
C9896 Iout.n72 VGND 0.02663f
C9897 Iout.n73 VGND 0.24452f
C9898 Iout.t138 VGND 0.02354f
C9899 Iout.n74 VGND 0.05236f
C9900 Iout.n75 VGND 0.02663f
C9901 Iout.n76 VGND 0.24452f
C9902 Iout.t187 VGND 0.02354f
C9903 Iout.n77 VGND 0.05236f
C9904 Iout.n78 VGND 0.02663f
C9905 Iout.n79 VGND 0.24452f
C9906 Iout.n80 VGND 0.24452f
C9907 Iout.t186 VGND 0.02354f
C9908 Iout.n81 VGND 0.05236f
C9909 Iout.n82 VGND 0.02663f
C9910 Iout.n83 VGND 0.24452f
C9911 Iout.n84 VGND 0.04879f
C9912 Iout.t90 VGND 0.02354f
C9913 Iout.n85 VGND 0.05236f
C9914 Iout.n86 VGND 0.02663f
C9915 Iout.t247 VGND 0.02354f
C9916 Iout.n87 VGND 0.05236f
C9917 Iout.n88 VGND 0.02663f
C9918 Iout.n89 VGND 0.24452f
C9919 Iout.t52 VGND 0.02354f
C9920 Iout.n90 VGND 0.05236f
C9921 Iout.n91 VGND 0.02663f
C9922 Iout.n92 VGND 0.24452f
C9923 Iout.t115 VGND 0.02354f
C9924 Iout.n93 VGND 0.05236f
C9925 Iout.n94 VGND 0.02663f
C9926 Iout.n95 VGND 0.24452f
C9927 Iout.t126 VGND 0.02354f
C9928 Iout.n96 VGND 0.05236f
C9929 Iout.n97 VGND 0.02663f
C9930 Iout.n98 VGND 0.24452f
C9931 Iout.t148 VGND 0.02354f
C9932 Iout.n99 VGND 0.05236f
C9933 Iout.n100 VGND 0.02663f
C9934 Iout.n101 VGND 0.24452f
C9935 Iout.t35 VGND 0.02354f
C9936 Iout.n102 VGND 0.05236f
C9937 Iout.n103 VGND 0.02663f
C9938 Iout.n104 VGND 0.24452f
C9939 Iout.t180 VGND 0.02354f
C9940 Iout.n105 VGND 0.05236f
C9941 Iout.n106 VGND 0.02663f
C9942 Iout.n107 VGND 0.24452f
C9943 Iout.t153 VGND 0.02354f
C9944 Iout.n108 VGND 0.05236f
C9945 Iout.n109 VGND 0.02663f
C9946 Iout.n110 VGND 0.24452f
C9947 Iout.t193 VGND 0.02354f
C9948 Iout.n111 VGND 0.05236f
C9949 Iout.n112 VGND 0.02663f
C9950 Iout.n113 VGND 0.24452f
C9951 Iout.t10 VGND 0.02354f
C9952 Iout.n114 VGND 0.05236f
C9953 Iout.n115 VGND 0.02663f
C9954 Iout.n116 VGND 0.24452f
C9955 Iout.t191 VGND 0.02354f
C9956 Iout.n117 VGND 0.05236f
C9957 Iout.n118 VGND 0.02663f
C9958 Iout.n119 VGND 0.24452f
C9959 Iout.t81 VGND 0.02354f
C9960 Iout.n120 VGND 0.05236f
C9961 Iout.n121 VGND 0.02663f
C9962 Iout.n122 VGND 0.04879f
C9963 Iout.t239 VGND 0.02354f
C9964 Iout.n123 VGND 0.05236f
C9965 Iout.n124 VGND 0.02663f
C9966 Iout.n125 VGND 0.24452f
C9967 Iout.n126 VGND 0.24452f
C9968 Iout.t88 VGND 0.02354f
C9969 Iout.n127 VGND 0.05236f
C9970 Iout.n128 VGND 0.02663f
C9971 Iout.n129 VGND 0.04879f
C9972 Iout.t234 VGND 0.02354f
C9973 Iout.n130 VGND 0.05236f
C9974 Iout.n131 VGND 0.02663f
C9975 Iout.n132 VGND 0.24452f
C9976 Iout.t26 VGND 0.02354f
C9977 Iout.n133 VGND 0.05236f
C9978 Iout.n134 VGND 0.02663f
C9979 Iout.n135 VGND 0.04879f
C9980 Iout.t78 VGND 0.02354f
C9981 Iout.n136 VGND 0.05236f
C9982 Iout.n137 VGND 0.02663f
C9983 Iout.n138 VGND 0.24452f
C9984 Iout.n139 VGND 0.24452f
C9985 Iout.t68 VGND 0.02354f
C9986 Iout.n140 VGND 0.05236f
C9987 Iout.n141 VGND 0.02663f
C9988 Iout.n142 VGND 0.04879f
C9989 Iout.t39 VGND 0.02354f
C9990 Iout.n143 VGND 0.05236f
C9991 Iout.n144 VGND 0.02663f
C9992 Iout.n145 VGND 0.14435f
C9993 Iout.t33 VGND 0.02354f
C9994 Iout.n146 VGND 0.05236f
C9995 Iout.n147 VGND 0.02663f
C9996 Iout.n148 VGND 0.04879f
C9997 Iout.t21 VGND 0.02354f
C9998 Iout.n149 VGND 0.05236f
C9999 Iout.n150 VGND 0.02663f
C10000 Iout.n151 VGND 0.24452f
C10001 Iout.n152 VGND 0.14435f
C10002 Iout.n153 VGND 0.24452f
C10003 Iout.n154 VGND 0.24452f
C10004 Iout.n155 VGND 0.24452f
C10005 Iout.t178 VGND 0.02354f
C10006 Iout.n156 VGND 0.05236f
C10007 Iout.n157 VGND 0.02663f
C10008 Iout.n158 VGND 0.24452f
C10009 Iout.n159 VGND 0.24452f
C10010 Iout.n160 VGND 0.24452f
C10011 Iout.n161 VGND 0.24452f
C10012 Iout.n162 VGND 0.24452f
C10013 Iout.n163 VGND 0.24452f
C10014 Iout.n164 VGND 0.24452f
C10015 Iout.n165 VGND 0.24452f
C10016 Iout.n166 VGND 0.24452f
C10017 Iout.n167 VGND 0.24452f
C10018 Iout.t22 VGND 0.02354f
C10019 Iout.n168 VGND 0.05236f
C10020 Iout.n169 VGND 0.02663f
C10021 Iout.n170 VGND 0.24452f
C10022 Iout.n171 VGND 0.04879f
C10023 Iout.t124 VGND 0.02354f
C10024 Iout.n172 VGND 0.05236f
C10025 Iout.n173 VGND 0.02663f
C10026 Iout.t135 VGND 0.02354f
C10027 Iout.n174 VGND 0.05236f
C10028 Iout.n175 VGND 0.02663f
C10029 Iout.n176 VGND 0.24452f
C10030 Iout.t84 VGND 0.02354f
C10031 Iout.n177 VGND 0.05236f
C10032 Iout.n178 VGND 0.02663f
C10033 Iout.n179 VGND 0.24452f
C10034 Iout.t60 VGND 0.02354f
C10035 Iout.n180 VGND 0.05236f
C10036 Iout.n181 VGND 0.02663f
C10037 Iout.n182 VGND 0.24452f
C10038 Iout.t0 VGND 0.02354f
C10039 Iout.n183 VGND 0.05236f
C10040 Iout.n184 VGND 0.02663f
C10041 Iout.n185 VGND 0.24452f
C10042 Iout.t204 VGND 0.02354f
C10043 Iout.n186 VGND 0.05236f
C10044 Iout.n187 VGND 0.02663f
C10045 Iout.n188 VGND 0.24452f
C10046 Iout.t64 VGND 0.02354f
C10047 Iout.n189 VGND 0.05236f
C10048 Iout.n190 VGND 0.02663f
C10049 Iout.n191 VGND 0.14435f
C10050 Iout.t43 VGND 0.02354f
C10051 Iout.n192 VGND 0.05236f
C10052 Iout.n193 VGND 0.02663f
C10053 Iout.n194 VGND 0.04879f
C10054 Iout.t232 VGND 0.02354f
C10055 Iout.n195 VGND 0.05236f
C10056 Iout.n196 VGND 0.02663f
C10057 Iout.n197 VGND 0.14435f
C10058 Iout.n198 VGND 0.04879f
C10059 Iout.t169 VGND 0.02354f
C10060 Iout.n199 VGND 0.05236f
C10061 Iout.n200 VGND 0.02663f
C10062 Iout.n201 VGND 0.04879f
C10063 Iout.t225 VGND 0.02354f
C10064 Iout.n202 VGND 0.05236f
C10065 Iout.n203 VGND 0.02663f
C10066 Iout.n204 VGND 0.14435f
C10067 Iout.n205 VGND 0.04879f
C10068 Iout.t56 VGND 0.02354f
C10069 Iout.n206 VGND 0.05236f
C10070 Iout.n207 VGND 0.02663f
C10071 Iout.n208 VGND 0.14435f
C10072 Iout.n209 VGND 0.04879f
C10073 Iout.t69 VGND 0.02354f
C10074 Iout.n210 VGND 0.05236f
C10075 Iout.n211 VGND 0.02663f
C10076 Iout.n212 VGND 0.14435f
C10077 Iout.n213 VGND 0.04879f
C10078 Iout.t128 VGND 0.02354f
C10079 Iout.n214 VGND 0.05236f
C10080 Iout.n215 VGND 0.02663f
C10081 Iout.n216 VGND 0.14435f
C10082 Iout.n217 VGND 0.04879f
C10083 Iout.t46 VGND 0.02354f
C10084 Iout.n218 VGND 0.05236f
C10085 Iout.n219 VGND 0.02663f
C10086 Iout.n220 VGND 0.14435f
C10087 Iout.n221 VGND 0.04879f
C10088 Iout.t233 VGND 0.02354f
C10089 Iout.n222 VGND 0.05236f
C10090 Iout.n223 VGND 0.02663f
C10091 Iout.n224 VGND 0.14435f
C10092 Iout.n225 VGND 0.04879f
C10093 Iout.t252 VGND 0.02354f
C10094 Iout.n226 VGND 0.05236f
C10095 Iout.n227 VGND 0.02663f
C10096 Iout.n228 VGND 0.04879f
C10097 Iout.n229 VGND 0.14435f
C10098 Iout.n230 VGND 0.24452f
C10099 Iout.n231 VGND 0.04879f
C10100 Iout.t136 VGND 0.02354f
C10101 Iout.n232 VGND 0.05236f
C10102 Iout.n233 VGND 0.02663f
C10103 Iout.n234 VGND 0.04879f
C10104 Iout.t157 VGND 0.02354f
C10105 Iout.n235 VGND 0.05236f
C10106 Iout.n236 VGND 0.02663f
C10107 Iout.n237 VGND 0.04879f
C10108 Iout.t15 VGND 0.02354f
C10109 Iout.n238 VGND 0.05236f
C10110 Iout.n239 VGND 0.02663f
C10111 Iout.n240 VGND 0.04879f
C10112 Iout.t1 VGND 0.02354f
C10113 Iout.n241 VGND 0.05236f
C10114 Iout.n242 VGND 0.02663f
C10115 Iout.n243 VGND 0.04879f
C10116 Iout.t221 VGND 0.02354f
C10117 Iout.n244 VGND 0.05236f
C10118 Iout.n245 VGND 0.02663f
C10119 Iout.n246 VGND 0.04879f
C10120 Iout.t18 VGND 0.02354f
C10121 Iout.n247 VGND 0.05236f
C10122 Iout.n248 VGND 0.02663f
C10123 Iout.n249 VGND 0.04879f
C10124 Iout.t238 VGND 0.02354f
C10125 Iout.n250 VGND 0.05236f
C10126 Iout.n251 VGND 0.02663f
C10127 Iout.t212 VGND 0.02354f
C10128 Iout.n252 VGND 0.05236f
C10129 Iout.n253 VGND 0.02663f
C10130 Iout.n254 VGND 0.04879f
C10131 Iout.t237 VGND 0.02354f
C10132 Iout.n255 VGND 0.05236f
C10133 Iout.n256 VGND 0.02663f
C10134 Iout.n257 VGND 0.04879f
C10135 Iout.n258 VGND 0.24452f
C10136 Iout.t198 VGND 0.02354f
C10137 Iout.n259 VGND 0.05236f
C10138 Iout.n260 VGND 0.02663f
C10139 Iout.n261 VGND 0.04879f
C10140 Iout.n262 VGND 0.24452f
C10141 Iout.n263 VGND 0.24452f
C10142 Iout.n264 VGND 0.04879f
C10143 Iout.t144 VGND 0.02354f
C10144 Iout.n265 VGND 0.05236f
C10145 Iout.n266 VGND 0.02663f
C10146 Iout.n267 VGND 0.04879f
C10147 Iout.n268 VGND 0.24452f
C10148 Iout.n269 VGND 0.24452f
C10149 Iout.n270 VGND 0.04879f
C10150 Iout.t65 VGND 0.02354f
C10151 Iout.n271 VGND 0.05236f
C10152 Iout.n272 VGND 0.02663f
C10153 Iout.n273 VGND 0.04879f
C10154 Iout.n274 VGND 0.24452f
C10155 Iout.n275 VGND 0.24452f
C10156 Iout.n276 VGND 0.04879f
C10157 Iout.t154 VGND 0.02354f
C10158 Iout.n277 VGND 0.05236f
C10159 Iout.n278 VGND 0.02663f
C10160 Iout.n279 VGND 0.04879f
C10161 Iout.n280 VGND 0.24452f
C10162 Iout.n281 VGND 0.24452f
C10163 Iout.n282 VGND 0.04879f
C10164 Iout.t140 VGND 0.02354f
C10165 Iout.n283 VGND 0.05236f
C10166 Iout.n284 VGND 0.02663f
C10167 Iout.n285 VGND 0.04879f
C10168 Iout.n286 VGND 0.24452f
C10169 Iout.n287 VGND 0.24452f
C10170 Iout.n288 VGND 0.04879f
C10171 Iout.t215 VGND 0.02354f
C10172 Iout.n289 VGND 0.05236f
C10173 Iout.n290 VGND 0.02663f
C10174 Iout.n291 VGND 0.04879f
C10175 Iout.n292 VGND 0.24452f
C10176 Iout.n293 VGND 0.24452f
C10177 Iout.n294 VGND 0.04879f
C10178 Iout.t149 VGND 0.02354f
C10179 Iout.n295 VGND 0.05236f
C10180 Iout.n296 VGND 0.02663f
C10181 Iout.n297 VGND 0.04879f
C10182 Iout.n298 VGND 0.24452f
C10183 Iout.n299 VGND 0.24452f
C10184 Iout.n300 VGND 0.04879f
C10185 Iout.t7 VGND 0.02354f
C10186 Iout.n301 VGND 0.05236f
C10187 Iout.n302 VGND 0.02663f
C10188 Iout.n303 VGND 0.04879f
C10189 Iout.n304 VGND 0.24452f
C10190 Iout.t118 VGND 0.02354f
C10191 Iout.n305 VGND 0.05236f
C10192 Iout.n306 VGND 0.02663f
C10193 Iout.n307 VGND 0.04879f
C10194 Iout.t91 VGND 0.02354f
C10195 Iout.n308 VGND 0.05236f
C10196 Iout.n309 VGND 0.02663f
C10197 Iout.n310 VGND 0.04879f
C10198 Iout.t222 VGND 0.02354f
C10199 Iout.n311 VGND 0.05236f
C10200 Iout.n312 VGND 0.02663f
C10201 Iout.n313 VGND 0.04879f
C10202 Iout.t67 VGND 0.02354f
C10203 Iout.n314 VGND 0.05236f
C10204 Iout.n315 VGND 0.02663f
C10205 Iout.n316 VGND 0.04879f
C10206 Iout.t8 VGND 0.02354f
C10207 Iout.n317 VGND 0.05236f
C10208 Iout.n318 VGND 0.02663f
C10209 Iout.n319 VGND 0.04879f
C10210 Iout.t182 VGND 0.02354f
C10211 Iout.n320 VGND 0.05236f
C10212 Iout.n321 VGND 0.02663f
C10213 Iout.n322 VGND 0.04879f
C10214 Iout.t130 VGND 0.02354f
C10215 Iout.n323 VGND 0.05236f
C10216 Iout.n324 VGND 0.02663f
C10217 Iout.n325 VGND 0.04879f
C10218 Iout.t145 VGND 0.02354f
C10219 Iout.n326 VGND 0.05236f
C10220 Iout.n327 VGND 0.02663f
C10221 Iout.n328 VGND 0.04879f
C10222 Iout.t2 VGND 0.02354f
C10223 Iout.n329 VGND 0.05236f
C10224 Iout.n330 VGND 0.02663f
C10225 Iout.n331 VGND 0.04879f
C10226 Iout.n332 VGND 0.24452f
C10227 Iout.t41 VGND 0.02354f
C10228 Iout.n333 VGND 0.05236f
C10229 Iout.n334 VGND 0.02663f
C10230 Iout.n335 VGND 0.04879f
C10231 Iout.t230 VGND 0.02354f
C10232 Iout.n336 VGND 0.05236f
C10233 Iout.n337 VGND 0.02663f
C10234 Iout.n338 VGND 0.04879f
C10235 Iout.t141 VGND 0.02354f
C10236 Iout.n339 VGND 0.05236f
C10237 Iout.n340 VGND 0.02663f
C10238 Iout.n341 VGND 0.04879f
C10239 Iout.t190 VGND 0.02354f
C10240 Iout.n342 VGND 0.05236f
C10241 Iout.n343 VGND 0.02663f
C10242 Iout.n344 VGND 0.04879f
C10243 Iout.t229 VGND 0.02354f
C10244 Iout.n345 VGND 0.05236f
C10245 Iout.n346 VGND 0.02663f
C10246 Iout.n347 VGND 0.04879f
C10247 Iout.t32 VGND 0.02354f
C10248 Iout.n348 VGND 0.05236f
C10249 Iout.n349 VGND 0.02663f
C10250 Iout.n350 VGND 0.04879f
C10251 Iout.t224 VGND 0.02354f
C10252 Iout.n351 VGND 0.05236f
C10253 Iout.n352 VGND 0.02663f
C10254 Iout.n353 VGND 0.04879f
C10255 Iout.t93 VGND 0.02354f
C10256 Iout.n354 VGND 0.05236f
C10257 Iout.n355 VGND 0.02663f
C10258 Iout.n356 VGND 0.04879f
C10259 Iout.t86 VGND 0.02354f
C10260 Iout.n357 VGND 0.05236f
C10261 Iout.n358 VGND 0.02663f
C10262 Iout.n359 VGND 0.04879f
C10263 Iout.t37 VGND 0.02354f
C10264 Iout.n360 VGND 0.05236f
C10265 Iout.n361 VGND 0.02663f
C10266 Iout.n362 VGND 0.04879f
C10267 Iout.t146 VGND 0.02354f
C10268 Iout.n363 VGND 0.05236f
C10269 Iout.n364 VGND 0.02663f
C10270 Iout.n365 VGND 0.04879f
C10271 Iout.t30 VGND 0.02354f
C10272 Iout.n366 VGND 0.05236f
C10273 Iout.n367 VGND 0.02663f
C10274 Iout.n368 VGND 0.04879f
C10275 Iout.n369 VGND 0.24452f
C10276 Iout.t77 VGND 0.02354f
C10277 Iout.n370 VGND 0.05236f
C10278 Iout.n371 VGND 0.02663f
C10279 Iout.n372 VGND 0.04879f
C10280 Iout.n373 VGND 0.24452f
C10281 Iout.n374 VGND 0.24452f
C10282 Iout.n375 VGND 0.04879f
C10283 Iout.t223 VGND 0.02354f
C10284 Iout.n376 VGND 0.05236f
C10285 Iout.n377 VGND 0.02663f
C10286 Iout.t29 VGND 0.02354f
C10287 Iout.n378 VGND 0.05236f
C10288 Iout.n379 VGND 0.02663f
C10289 Iout.n380 VGND 0.04879f
C10290 Iout.n381 VGND 0.24452f
C10291 Iout.n382 VGND 0.24452f
C10292 Iout.n383 VGND 0.04879f
C10293 Iout.t183 VGND 0.02354f
C10294 Iout.n384 VGND 0.05236f
C10295 Iout.n385 VGND 0.02663f
C10296 Iout.t99 VGND 0.02354f
C10297 Iout.n386 VGND 0.05236f
C10298 Iout.n387 VGND 0.02663f
C10299 Iout.n388 VGND 0.04879f
C10300 Iout.n389 VGND 0.24452f
C10301 Iout.n390 VGND 0.24452f
C10302 Iout.n391 VGND 0.04879f
C10303 Iout.t104 VGND 0.02354f
C10304 Iout.n392 VGND 0.05236f
C10305 Iout.n393 VGND 0.02663f
C10306 Iout.t244 VGND 0.02354f
C10307 Iout.n394 VGND 0.05236f
C10308 Iout.n395 VGND 0.02663f
C10309 Iout.n396 VGND 0.04879f
C10310 Iout.n397 VGND 0.24452f
C10311 Iout.n398 VGND 0.24452f
C10312 Iout.n399 VGND 0.04879f
C10313 Iout.t254 VGND 0.02354f
C10314 Iout.n400 VGND 0.05236f
C10315 Iout.n401 VGND 0.02663f
C10316 Iout.t55 VGND 0.02354f
C10317 Iout.n402 VGND 0.05236f
C10318 Iout.n403 VGND 0.02663f
C10319 Iout.n404 VGND 0.04879f
C10320 Iout.n405 VGND 0.24452f
C10321 Iout.n406 VGND 0.24452f
C10322 Iout.n407 VGND 0.04879f
C10323 Iout.t16 VGND 0.02354f
C10324 Iout.n408 VGND 0.05236f
C10325 Iout.n409 VGND 0.02663f
C10326 Iout.t240 VGND 0.02354f
C10327 Iout.n410 VGND 0.05236f
C10328 Iout.n411 VGND 0.02663f
C10329 Iout.n412 VGND 0.04879f
C10330 Iout.n413 VGND 0.24452f
C10331 Iout.n414 VGND 0.24452f
C10332 Iout.n415 VGND 0.04879f
C10333 Iout.t70 VGND 0.02354f
C10334 Iout.n416 VGND 0.05236f
C10335 Iout.n417 VGND 0.02663f
C10336 Iout.t132 VGND 0.02354f
C10337 Iout.n418 VGND 0.05236f
C10338 Iout.n419 VGND 0.02663f
C10339 Iout.n420 VGND 0.04879f
C10340 Iout.n421 VGND 0.24452f
C10341 Iout.n422 VGND 0.24452f
C10342 Iout.n423 VGND 0.04879f
C10343 Iout.t152 VGND 0.02354f
C10344 Iout.n424 VGND 0.05236f
C10345 Iout.n425 VGND 0.02663f
C10346 Iout.t206 VGND 0.02354f
C10347 Iout.n426 VGND 0.05236f
C10348 Iout.n427 VGND 0.02663f
C10349 Iout.n428 VGND 0.04879f
C10350 Iout.n429 VGND 0.24452f
C10351 Iout.n430 VGND 0.24452f
C10352 Iout.n431 VGND 0.04879f
C10353 Iout.t142 VGND 0.02354f
C10354 Iout.n432 VGND 0.05236f
C10355 Iout.n433 VGND 0.02663f
C10356 Iout.t194 VGND 0.02354f
C10357 Iout.n434 VGND 0.05236f
C10358 Iout.n435 VGND 0.02663f
C10359 Iout.n436 VGND 0.24452f
C10360 Iout.n437 VGND 0.04879f
C10361 Iout.t156 VGND 0.02354f
C10362 Iout.n438 VGND 0.05236f
C10363 Iout.n439 VGND 0.02663f
C10364 Iout.n440 VGND 0.04879f
C10365 Iout.t76 VGND 0.02354f
C10366 Iout.n441 VGND 0.05236f
C10367 Iout.n442 VGND 0.02663f
C10368 Iout.n443 VGND 0.04879f
C10369 Iout.n444 VGND 0.24452f
C10370 Iout.n445 VGND 0.24452f
C10371 Iout.n446 VGND 0.04879f
C10372 Iout.t226 VGND 0.02354f
C10373 Iout.n447 VGND 0.05236f
C10374 Iout.n448 VGND 0.02663f
C10375 Iout.t184 VGND 0.02354f
C10376 Iout.n449 VGND 0.05236f
C10377 Iout.n450 VGND 0.02663f
C10378 Iout.n451 VGND 0.04879f
C10379 Iout.t173 VGND 0.02354f
C10380 Iout.n452 VGND 0.05236f
C10381 Iout.n453 VGND 0.02663f
C10382 Iout.n454 VGND 0.04879f
C10383 Iout.n455 VGND 0.24452f
C10384 Iout.n456 VGND 0.24452f
C10385 Iout.n457 VGND 0.04879f
C10386 Iout.t25 VGND 0.02354f
C10387 Iout.n458 VGND 0.05236f
C10388 Iout.n459 VGND 0.02663f
C10389 Iout.t158 VGND 0.02354f
C10390 Iout.n460 VGND 0.05236f
C10391 Iout.n461 VGND 0.02663f
C10392 Iout.n462 VGND 0.04879f
C10393 Iout.t63 VGND 0.02354f
C10394 Iout.n463 VGND 0.05236f
C10395 Iout.n464 VGND 0.02663f
C10396 Iout.n465 VGND 0.04879f
C10397 Iout.n466 VGND 0.24452f
C10398 Iout.n467 VGND 0.24452f
C10399 Iout.n468 VGND 0.04879f
C10400 Iout.t249 VGND 0.02354f
C10401 Iout.n469 VGND 0.05236f
C10402 Iout.n470 VGND 0.02663f
C10403 Iout.n471 VGND 0.04879f
C10404 Iout.t53 VGND 0.02354f
C10405 Iout.n472 VGND 0.05236f
C10406 Iout.n473 VGND 0.02663f
C10407 Iout.n474 VGND 0.04879f
C10408 Iout.n475 VGND 0.24452f
C10409 Iout.n476 VGND 0.24452f
C10410 Iout.n477 VGND 0.04879f
C10411 Iout.t200 VGND 0.02354f
C10412 Iout.n478 VGND 0.05236f
C10413 Iout.n479 VGND 0.02663f
C10414 Iout.t147 VGND 0.02354f
C10415 Iout.n480 VGND 0.05236f
C10416 Iout.n481 VGND 0.02663f
C10417 Iout.n482 VGND 0.04879f
C10418 Iout.t192 VGND 0.02354f
C10419 Iout.n483 VGND 0.05236f
C10420 Iout.n484 VGND 0.02663f
C10421 Iout.n485 VGND 0.04879f
C10422 Iout.n486 VGND 0.24452f
C10423 Iout.n487 VGND 0.24452f
C10424 Iout.n488 VGND 0.04879f
C10425 Iout.t228 VGND 0.02354f
C10426 Iout.n489 VGND 0.05236f
C10427 Iout.n490 VGND 0.02663f
C10428 Iout.t28 VGND 0.02354f
C10429 Iout.n491 VGND 0.05236f
C10430 Iout.n492 VGND 0.02663f
C10431 Iout.n493 VGND 0.04879f
C10432 Iout.t197 VGND 0.02354f
C10433 Iout.n494 VGND 0.05236f
C10434 Iout.n495 VGND 0.02663f
C10435 Iout.n496 VGND 0.04879f
C10436 Iout.n497 VGND 0.24452f
C10437 Iout.n498 VGND 0.14435f
C10438 Iout.n499 VGND 0.04879f
C10439 Iout.t80 VGND 0.02354f
C10440 Iout.n500 VGND 0.05236f
C10441 Iout.n501 VGND 0.02663f
C10442 Iout.n502 VGND 0.14435f
C10443 Iout.n503 VGND 0.04879f
C10444 Iout.t114 VGND 0.02354f
C10445 Iout.n504 VGND 0.05236f
C10446 Iout.n505 VGND 0.02663f
C10447 Iout.n506 VGND 0.04879f
C10448 Iout.t108 VGND 0.02354f
C10449 Iout.n507 VGND 0.05236f
C10450 Iout.n508 VGND 0.02663f
C10451 Iout.t210 VGND 0.02354f
C10452 Iout.n509 VGND 0.05236f
C10453 Iout.n510 VGND 0.02663f
C10454 Iout.n511 VGND 0.14435f
C10455 Iout.n512 VGND 0.04879f
C10456 Iout.t175 VGND 0.02354f
C10457 Iout.n513 VGND 0.05236f
C10458 Iout.n514 VGND 0.02663f
C10459 Iout.n515 VGND 0.04879f
C10460 Iout.n516 VGND 0.14435f
C10461 Iout.n517 VGND 0.24452f
C10462 Iout.n518 VGND 0.04879f
C10463 Iout.t250 VGND 0.02354f
C10464 Iout.n519 VGND 0.05236f
C10465 Iout.n520 VGND 0.02663f
C10466 Iout.n521 VGND 0.04879f
C10467 Iout.n522 VGND 0.24452f
C10468 Iout.n523 VGND 0.24452f
C10469 Iout.n524 VGND 0.04879f
C10470 Iout.t27 VGND 0.02354f
C10471 Iout.n525 VGND 0.05236f
C10472 Iout.n526 VGND 0.02663f
C10473 Iout.n527 VGND 0.04879f
C10474 Iout.n528 VGND 0.24452f
C10475 Iout.n529 VGND 0.24452f
C10476 Iout.n530 VGND 0.04879f
C10477 Iout.t236 VGND 0.02354f
C10478 Iout.n531 VGND 0.05236f
C10479 Iout.n532 VGND 0.02663f
C10480 Iout.n533 VGND 0.04879f
C10481 Iout.t105 VGND 0.02354f
C10482 Iout.n534 VGND 0.05236f
C10483 Iout.n535 VGND 0.02663f
C10484 Iout.t44 VGND 0.02354f
C10485 Iout.n536 VGND 0.05236f
C10486 Iout.n537 VGND 0.02663f
C10487 Iout.n538 VGND 0.04879f
C10488 Iout.n539 VGND 0.24452f
C10489 Iout.n540 VGND 0.24452f
C10490 Iout.n541 VGND 0.04879f
C10491 Iout.t161 VGND 0.02354f
C10492 Iout.n542 VGND 0.05236f
C10493 Iout.n543 VGND 0.02663f
C10494 Iout.n544 VGND 0.04879f
C10495 Iout.n545 VGND 0.24452f
C10496 Iout.n546 VGND 0.24452f
C10497 Iout.n547 VGND 0.04879f
C10498 Iout.t75 VGND 0.02354f
C10499 Iout.n548 VGND 0.05236f
C10500 Iout.n549 VGND 0.02663f
C10501 Iout.n550 VGND 0.04879f
C10502 Iout.n551 VGND 0.24452f
C10503 Iout.n552 VGND 0.24452f
C10504 Iout.n553 VGND 0.04879f
C10505 Iout.t151 VGND 0.02354f
C10506 Iout.n554 VGND 0.05236f
C10507 Iout.n555 VGND 0.02663f
C10508 Iout.n556 VGND 0.04879f
C10509 Iout.t231 VGND 0.02354f
C10510 Iout.n557 VGND 0.05236f
C10511 Iout.n558 VGND 0.02663f
C10512 Iout.t131 VGND 0.02354f
C10513 Iout.n559 VGND 0.05236f
C10514 Iout.n560 VGND 0.02663f
C10515 Iout.n561 VGND 0.04879f
C10516 Iout.n562 VGND 0.24452f
C10517 Iout.t85 VGND 0.02354f
C10518 Iout.n563 VGND 0.05236f
C10519 Iout.n564 VGND 0.02663f
C10520 Iout.n565 VGND 0.04879f
C10521 Iout.n566 VGND 0.24452f
C10522 Iout.n567 VGND 0.24452f
C10523 Iout.n568 VGND 0.04879f
C10524 Iout.t242 VGND 0.02354f
C10525 Iout.n569 VGND 0.05236f
C10526 Iout.n570 VGND 0.02663f
C10527 Iout.n571 VGND 0.04879f
C10528 Iout.n572 VGND 0.24452f
C10529 Iout.t19 VGND 0.02354f
C10530 Iout.n573 VGND 0.05236f
C10531 Iout.n574 VGND 0.02663f
C10532 Iout.n575 VGND 0.04879f
C10533 Iout.t172 VGND 0.02354f
C10534 Iout.n576 VGND 0.05236f
C10535 Iout.n577 VGND 0.02663f
C10536 Iout.n578 VGND 0.04879f
C10537 Iout.n579 VGND 0.24452f
C10538 Iout.n580 VGND 0.24452f
C10539 Iout.n581 VGND 0.04879f
C10540 Iout.t235 VGND 0.02354f
C10541 Iout.n582 VGND 0.05236f
C10542 Iout.n583 VGND 0.02663f
C10543 Iout.n584 VGND 0.04879f
C10544 Iout.n585 VGND 0.24452f
C10545 Iout.n586 VGND 0.24452f
C10546 Iout.n587 VGND 0.04879f
C10547 Iout.t48 VGND 0.02354f
C10548 Iout.n588 VGND 0.05236f
C10549 Iout.n589 VGND 0.02663f
C10550 Iout.n590 VGND 0.04879f
C10551 Iout.n591 VGND 0.24452f
C10552 Iout.n592 VGND 0.24452f
C10553 Iout.n593 VGND 0.04879f
C10554 Iout.t34 VGND 0.02354f
C10555 Iout.n594 VGND 0.05236f
C10556 Iout.n595 VGND 0.02663f
C10557 Iout.n596 VGND 0.04879f
C10558 Iout.n597 VGND 0.24452f
C10559 Iout.n598 VGND 0.24452f
C10560 Iout.n599 VGND 0.04879f
C10561 Iout.t143 VGND 0.02354f
C10562 Iout.n600 VGND 0.05236f
C10563 Iout.n601 VGND 0.02663f
C10564 Iout.n602 VGND 0.04879f
C10565 Iout.n603 VGND 0.24452f
C10566 Iout.n604 VGND 0.24452f
C10567 Iout.n605 VGND 0.04879f
C10568 Iout.t203 VGND 0.02354f
C10569 Iout.n606 VGND 0.05236f
C10570 Iout.n607 VGND 0.02663f
C10571 Iout.n608 VGND 0.04879f
C10572 Iout.n609 VGND 0.24452f
C10573 Iout.n610 VGND 0.24452f
C10574 Iout.n611 VGND 0.04879f
C10575 Iout.t31 VGND 0.02354f
C10576 Iout.n612 VGND 0.05236f
C10577 Iout.n613 VGND 0.02663f
C10578 Iout.n614 VGND 0.04879f
C10579 Iout.n615 VGND 0.24452f
C10580 Iout.n616 VGND 0.24452f
C10581 Iout.n617 VGND 0.04879f
C10582 Iout.t255 VGND 0.02354f
C10583 Iout.n618 VGND 0.05236f
C10584 Iout.n619 VGND 0.02663f
C10585 Iout.n620 VGND 0.04879f
C10586 Iout.n621 VGND 0.24452f
C10587 Iout.n622 VGND 0.24452f
C10588 Iout.n623 VGND 0.04879f
C10589 Iout.t155 VGND 0.02354f
C10590 Iout.n624 VGND 0.05236f
C10591 Iout.n625 VGND 0.02663f
C10592 Iout.n626 VGND 0.04879f
C10593 Iout.n627 VGND 0.24452f
C10594 Iout.n628 VGND 0.24452f
C10595 Iout.n629 VGND 0.04879f
C10596 Iout.t82 VGND 0.02354f
C10597 Iout.n630 VGND 0.05236f
C10598 Iout.n631 VGND 0.02663f
C10599 Iout.n632 VGND 0.04879f
C10600 Iout.n633 VGND 0.24452f
C10601 Iout.n634 VGND 0.24452f
C10602 Iout.n635 VGND 0.04879f
C10603 Iout.t107 VGND 0.02354f
C10604 Iout.n636 VGND 0.05236f
C10605 Iout.n637 VGND 0.02663f
C10606 Iout.n638 VGND 0.04879f
C10607 Iout.n639 VGND 0.24452f
C10608 Iout.n640 VGND 0.24452f
C10609 Iout.n641 VGND 0.04879f
C10610 Iout.t23 VGND 0.02354f
C10611 Iout.n642 VGND 0.05236f
C10612 Iout.n643 VGND 0.02663f
C10613 Iout.n644 VGND 0.04879f
C10614 Iout.n645 VGND 0.24452f
C10615 Iout.n646 VGND 0.24452f
C10616 Iout.n647 VGND 0.04879f
C10617 Iout.t209 VGND 0.02354f
C10618 Iout.n648 VGND 0.05236f
C10619 Iout.n649 VGND 0.02663f
C10620 Iout.n650 VGND 0.04879f
C10621 Iout.n651 VGND 0.24452f
C10622 Iout.n652 VGND 0.24452f
C10623 Iout.n653 VGND 0.04879f
C10624 Iout.t164 VGND 0.02354f
C10625 Iout.n654 VGND 0.05236f
C10626 Iout.n655 VGND 0.02663f
C10627 Iout.n656 VGND 0.04879f
C10628 Iout.t113 VGND 0.02354f
C10629 Iout.n657 VGND 0.05236f
C10630 Iout.n658 VGND 0.02663f
C10631 Iout.n659 VGND 0.04879f
C10632 Iout.t179 VGND 0.02354f
C10633 Iout.n660 VGND 0.05236f
C10634 Iout.n661 VGND 0.02663f
C10635 Iout.n662 VGND 0.04879f
C10636 Iout.t62 VGND 0.02354f
C10637 Iout.n663 VGND 0.05236f
C10638 Iout.n664 VGND 0.02663f
C10639 Iout.n665 VGND 0.04879f
C10640 Iout.t122 VGND 0.02354f
C10641 Iout.n666 VGND 0.05236f
C10642 Iout.n667 VGND 0.02663f
C10643 Iout.n668 VGND 0.04879f
C10644 Iout.t98 VGND 0.02354f
C10645 Iout.n669 VGND 0.05236f
C10646 Iout.n670 VGND 0.02663f
C10647 Iout.n671 VGND 0.04879f
C10648 Iout.t168 VGND 0.02354f
C10649 Iout.n672 VGND 0.05236f
C10650 Iout.n673 VGND 0.02663f
C10651 Iout.n674 VGND 0.04879f
C10652 Iout.t199 VGND 0.02354f
C10653 Iout.n675 VGND 0.05236f
C10654 Iout.n676 VGND 0.02663f
C10655 Iout.n677 VGND 0.04879f
C10656 Iout.t71 VGND 0.02354f
C10657 Iout.n678 VGND 0.05236f
C10658 Iout.n679 VGND 0.02663f
C10659 Iout.n680 VGND 0.04879f
C10660 Iout.t167 VGND 0.02354f
C10661 Iout.n681 VGND 0.05236f
C10662 Iout.n682 VGND 0.02663f
C10663 Iout.n683 VGND 0.04879f
C10664 Iout.t13 VGND 0.02354f
C10665 Iout.n684 VGND 0.05236f
C10666 Iout.n685 VGND 0.02663f
C10667 Iout.n686 VGND 0.04879f
C10668 Iout.t89 VGND 0.02354f
C10669 Iout.n687 VGND 0.05236f
C10670 Iout.n688 VGND 0.02663f
C10671 Iout.n689 VGND 0.04879f
C10672 Iout.t188 VGND 0.02354f
C10673 Iout.n690 VGND 0.05236f
C10674 Iout.n691 VGND 0.02663f
C10675 Iout.t163 VGND 0.02354f
C10676 Iout.n692 VGND 0.05236f
C10677 Iout.n693 VGND 0.02663f
C10678 Iout.n694 VGND 0.04879f
C10679 Iout.t47 VGND 0.02354f
C10680 Iout.n695 VGND 0.05236f
C10681 Iout.n696 VGND 0.02663f
C10682 Iout.n697 VGND 0.04879f
C10683 Iout.n698 VGND 0.24452f
C10684 Iout.t166 VGND 0.02354f
C10685 Iout.n699 VGND 0.05236f
C10686 Iout.n700 VGND 0.02663f
C10687 Iout.n701 VGND 0.04879f
C10688 Iout.n702 VGND 0.24452f
C10689 Iout.n703 VGND 0.24452f
C10690 Iout.n704 VGND 0.04879f
C10691 Iout.t123 VGND 0.02354f
C10692 Iout.n705 VGND 0.05236f
C10693 Iout.n706 VGND 0.02663f
C10694 Iout.n707 VGND 0.04879f
C10695 Iout.n708 VGND 0.24452f
C10696 Iout.n709 VGND 0.24452f
C10697 Iout.n710 VGND 0.04879f
C10698 Iout.t49 VGND 0.02354f
C10699 Iout.n711 VGND 0.05236f
C10700 Iout.n712 VGND 0.02663f
C10701 Iout.n713 VGND 0.04879f
C10702 Iout.n714 VGND 0.24452f
C10703 Iout.n715 VGND 0.24452f
C10704 Iout.n716 VGND 0.04879f
C10705 Iout.t134 VGND 0.02354f
C10706 Iout.n717 VGND 0.05236f
C10707 Iout.n718 VGND 0.02663f
C10708 Iout.n719 VGND 0.04879f
C10709 Iout.n720 VGND 0.24452f
C10710 Iout.n721 VGND 0.24452f
C10711 Iout.n722 VGND 0.04879f
C10712 Iout.t12 VGND 0.02354f
C10713 Iout.n723 VGND 0.05236f
C10714 Iout.n724 VGND 0.02663f
C10715 Iout.n725 VGND 0.04879f
C10716 Iout.n726 VGND 0.24452f
C10717 Iout.n727 VGND 0.24452f
C10718 Iout.n728 VGND 0.04879f
C10719 Iout.t217 VGND 0.02354f
C10720 Iout.n729 VGND 0.05236f
C10721 Iout.n730 VGND 0.02663f
C10722 Iout.n731 VGND 0.04879f
C10723 Iout.n732 VGND 0.24452f
C10724 Iout.n733 VGND 0.24452f
C10725 Iout.n734 VGND 0.04879f
C10726 Iout.t213 VGND 0.02354f
C10727 Iout.n735 VGND 0.05236f
C10728 Iout.n736 VGND 0.02663f
C10729 Iout.n737 VGND 0.04879f
C10730 Iout.n738 VGND 0.24452f
C10731 Iout.n739 VGND 0.24452f
C10732 Iout.n740 VGND 0.04879f
C10733 Iout.t4 VGND 0.02354f
C10734 Iout.n741 VGND 0.05236f
C10735 Iout.n742 VGND 0.02663f
C10736 Iout.n743 VGND 0.04879f
C10737 Iout.n744 VGND 0.24452f
C10738 Iout.n745 VGND 0.24452f
C10739 Iout.n746 VGND 0.04879f
C10740 Iout.t51 VGND 0.02354f
C10741 Iout.n747 VGND 0.05236f
C10742 Iout.n748 VGND 0.02663f
C10743 Iout.n749 VGND 0.04879f
C10744 Iout.n750 VGND 0.24452f
C10745 Iout.n751 VGND 0.24452f
C10746 Iout.n752 VGND 0.04879f
C10747 Iout.t110 VGND 0.02354f
C10748 Iout.n753 VGND 0.05236f
C10749 Iout.n754 VGND 0.02663f
C10750 Iout.n755 VGND 0.04879f
C10751 Iout.n756 VGND 0.24452f
C10752 Iout.n757 VGND 0.24452f
C10753 Iout.n758 VGND 0.04879f
C10754 Iout.t139 VGND 0.02354f
C10755 Iout.n759 VGND 0.05236f
C10756 Iout.n760 VGND 0.02663f
C10757 Iout.n761 VGND 0.04879f
C10758 Iout.n762 VGND 0.24452f
C10759 Iout.n763 VGND 0.24452f
C10760 Iout.n764 VGND 0.04879f
C10761 Iout.t150 VGND 0.02354f
C10762 Iout.n765 VGND 0.05236f
C10763 Iout.n766 VGND 0.02663f
C10764 Iout.n767 VGND 0.04879f
C10765 Iout.n768 VGND 0.24452f
C10766 Iout.n769 VGND 0.24452f
C10767 Iout.n770 VGND 0.04879f
C10768 Iout.t165 VGND 0.02354f
C10769 Iout.n771 VGND 0.05236f
C10770 Iout.n772 VGND 0.02663f
C10771 Iout.n773 VGND 0.04879f
C10772 Iout.n774 VGND 0.24452f
C10773 Iout.n775 VGND 0.24452f
C10774 Iout.n776 VGND 0.04879f
C10775 Iout.t58 VGND 0.02354f
C10776 Iout.n777 VGND 0.05236f
C10777 Iout.n778 VGND 0.02663f
C10778 Iout.n779 VGND 0.04879f
C10779 Iout.n780 VGND 0.24452f
C10780 Iout.t218 VGND 0.02354f
C10781 Iout.n781 VGND 0.05236f
C10782 Iout.n782 VGND 0.02663f
C10783 Iout.n783 VGND 0.04879f
C10784 Iout.t174 VGND 0.02354f
C10785 Iout.n784 VGND 0.05236f
C10786 Iout.n785 VGND 0.02663f
C10787 Iout.n786 VGND 0.04879f
C10788 Iout.t20 VGND 0.02354f
C10789 Iout.n787 VGND 0.05236f
C10790 Iout.n788 VGND 0.02663f
C10791 Iout.n789 VGND 0.04879f
C10792 Iout.t73 VGND 0.02354f
C10793 Iout.n790 VGND 0.05236f
C10794 Iout.n791 VGND 0.02663f
C10795 Iout.n792 VGND 0.04879f
C10796 Iout.t94 VGND 0.02354f
C10797 Iout.n793 VGND 0.05236f
C10798 Iout.n794 VGND 0.02663f
C10799 Iout.n795 VGND 0.04879f
C10800 Iout.t95 VGND 0.02354f
C10801 Iout.n796 VGND 0.05236f
C10802 Iout.n797 VGND 0.02663f
C10803 Iout.n798 VGND 0.04879f
C10804 Iout.t50 VGND 0.02354f
C10805 Iout.n799 VGND 0.05236f
C10806 Iout.n800 VGND 0.02663f
C10807 Iout.n801 VGND 0.04879f
C10808 Iout.t189 VGND 0.02354f
C10809 Iout.n802 VGND 0.05236f
C10810 Iout.n803 VGND 0.02663f
C10811 Iout.n804 VGND 0.04879f
C10812 Iout.t205 VGND 0.02354f
C10813 Iout.n805 VGND 0.05236f
C10814 Iout.n806 VGND 0.02663f
C10815 Iout.n807 VGND 0.04879f
C10816 Iout.t54 VGND 0.02354f
C10817 Iout.n808 VGND 0.05236f
C10818 Iout.n809 VGND 0.02663f
C10819 Iout.n810 VGND 0.04879f
C10820 Iout.t211 VGND 0.02354f
C10821 Iout.n811 VGND 0.05236f
C10822 Iout.n812 VGND 0.02663f
C10823 Iout.n813 VGND 0.04879f
C10824 Iout.t171 VGND 0.02354f
C10825 Iout.n814 VGND 0.05236f
C10826 Iout.n815 VGND 0.02663f
C10827 Iout.n816 VGND 0.04879f
C10828 Iout.t40 VGND 0.02354f
C10829 Iout.n817 VGND 0.05236f
C10830 Iout.n818 VGND 0.02663f
C10831 Iout.n819 VGND 0.04879f
C10832 Iout.t160 VGND 0.02354f
C10833 Iout.n820 VGND 0.05236f
C10834 Iout.n821 VGND 0.02663f
C10835 Iout.n822 VGND 0.04879f
C10836 Iout.t42 VGND 0.02354f
C10837 Iout.n823 VGND 0.05236f
C10838 Iout.n824 VGND 0.02663f
C10839 Iout.n825 VGND 0.04879f
C10840 Iout.n826 VGND 0.24452f
C10841 Iout.t208 VGND 0.02354f
C10842 Iout.n827 VGND 0.05236f
C10843 Iout.n828 VGND 0.02663f
C10844 Iout.n829 VGND 0.08346f
C10845 Iout.n830 VGND 0.50694f
C10846 Iout.n831 VGND 0.04879f
C10847 Iout.t246 VGND 0.02354f
C10848 Iout.n832 VGND 0.05236f
C10849 Iout.n833 VGND 0.02663f
C10850 Iout.t195 VGND 0.02354f
C10851 Iout.n834 VGND 0.05236f
C10852 Iout.n835 VGND 0.02663f
C10853 Iout.n836 VGND 0.04879f
C10854 Iout.n837 VGND 0.50694f
C10855 Iout.n838 VGND 0.08346f
C10856 Iout.t83 VGND 0.02354f
C10857 Iout.n839 VGND 0.05236f
C10858 Iout.n840 VGND 0.02663f
C10859 Iout.t251 VGND 0.02354f
C10860 Iout.n841 VGND 0.05236f
C10861 Iout.n842 VGND 0.02663f
C10862 Iout.n843 VGND 0.08346f
C10863 Iout.n844 VGND 0.50694f
C10864 Iout.n845 VGND 0.04879f
C10865 Iout.t45 VGND 0.02354f
C10866 Iout.n846 VGND 0.05236f
C10867 Iout.n847 VGND 0.02663f
C10868 Iout.t181 VGND 0.02354f
C10869 Iout.n848 VGND 0.05236f
C10870 Iout.n849 VGND 0.02663f
C10871 Iout.n850 VGND 0.04879f
C10872 Iout.n851 VGND 0.50694f
C10873 Iout.n852 VGND 0.08346f
C10874 Iout.t79 VGND 0.02354f
C10875 Iout.n853 VGND 0.05236f
C10876 Iout.n854 VGND 0.02663f
C10877 Iout.t185 VGND 0.02354f
C10878 Iout.n855 VGND 0.05236f
C10879 Iout.n856 VGND 0.02663f
C10880 Iout.n857 VGND 0.08346f
C10881 Iout.n858 VGND 0.50694f
C10882 Iout.n859 VGND 0.04879f
C10883 Iout.t17 VGND 0.02354f
C10884 Iout.n860 VGND 0.05236f
C10885 Iout.n861 VGND 0.02663f
C10886 Iout.t101 VGND 0.02354f
C10887 Iout.n862 VGND 0.05236f
C10888 Iout.n863 VGND 0.02663f
C10889 Iout.n864 VGND 0.04879f
C10890 Iout.n865 VGND 0.50694f
C10891 Iout.n866 VGND 0.08346f
C10892 Iout.t103 VGND 0.02354f
C10893 Iout.n867 VGND 0.05236f
C10894 Iout.n868 VGND 0.02663f
C10895 Iout.t117 VGND 0.02354f
C10896 Iout.n869 VGND 0.05236f
C10897 Iout.n870 VGND 0.02663f
C10898 Iout.n871 VGND 0.08346f
C10899 Iout.n872 VGND 0.50694f
C10900 Iout.n873 VGND 0.04879f
C10901 Iout.t106 VGND 0.02354f
C10902 Iout.n874 VGND 0.05236f
C10903 Iout.n875 VGND 0.02663f
C10904 Iout.t121 VGND 0.02354f
C10905 Iout.n876 VGND 0.05236f
C10906 Iout.n877 VGND 0.02663f
C10907 Iout.n878 VGND 0.04879f
C10908 Iout.n879 VGND 0.50694f
C10909 Iout.n880 VGND 0.08346f
C10910 Iout.t129 VGND 0.02354f
C10911 Iout.n881 VGND 0.05236f
C10912 Iout.n882 VGND 0.02663f
C10913 Iout.t3 VGND 0.02354f
C10914 Iout.n883 VGND 0.05236f
C10915 Iout.n884 VGND 0.02663f
C10916 Iout.n885 VGND 0.08346f
C10917 Iout.n886 VGND 0.50694f
C10918 Iout.n887 VGND 0.04879f
C10919 Iout.t137 VGND 0.02354f
C10920 Iout.n888 VGND 0.05236f
C10921 Iout.n889 VGND 0.02663f
C10922 Iout.t59 VGND 0.02354f
C10923 Iout.n890 VGND 0.05236f
C10924 Iout.n891 VGND 0.02663f
C10925 Iout.n892 VGND 0.04879f
C10926 Iout.n893 VGND 0.50694f
C10927 Iout.n894 VGND 0.08346f
C10928 Iout.t162 VGND 0.02354f
C10929 Iout.n895 VGND 0.05236f
C10930 Iout.n896 VGND 0.02663f
C10931 Iout.t248 VGND 0.02354f
C10932 Iout.n897 VGND 0.05236f
C10933 Iout.n898 VGND 0.02663f
C10934 Iout.n899 VGND 0.08346f
C10935 Iout.n900 VGND 0.50694f
C10936 Iout.n901 VGND 0.04879f
C10937 Iout.t241 VGND 0.02354f
C10938 Iout.n902 VGND 0.05236f
C10939 Iout.n903 VGND 0.02663f
C10940 Iout.t87 VGND 0.02354f
C10941 Iout.n904 VGND 0.05236f
C10942 Iout.n905 VGND 0.02663f
C10943 Iout.n906 VGND 0.04879f
C10944 Iout.n907 VGND 0.50694f
C10945 Iout.n908 VGND 0.08346f
C10946 Iout.t216 VGND 0.02354f
C10947 Iout.n909 VGND 0.05236f
C10948 Iout.n910 VGND 0.02663f
C10949 Iout.t159 VGND 0.02354f
C10950 Iout.n911 VGND 0.05236f
C10951 Iout.n912 VGND 0.02663f
C10952 Iout.n913 VGND 0.08346f
C10953 Iout.n914 VGND 0.50694f
C10954 Iout.n915 VGND 0.04879f
C10955 Iout.t219 VGND 0.02354f
C10956 Iout.n916 VGND 0.05236f
C10957 Iout.n917 VGND 0.02663f
C10958 Iout.t11 VGND 0.02354f
C10959 Iout.n918 VGND 0.05236f
C10960 Iout.n919 VGND 0.02663f
C10961 Iout.n920 VGND 0.04879f
C10962 Iout.n921 VGND 0.50694f
C10963 Iout.n922 VGND 0.08346f
C10964 Iout.t125 VGND 0.02354f
C10965 Iout.n923 VGND 0.05236f
C10966 Iout.n924 VGND 0.02663f
C10967 Iout.n925 VGND 0.08346f
C10968 Iout.t214 VGND 0.02354f
C10969 Iout.n926 VGND 0.05236f
C10970 Iout.n927 VGND 0.02663f
C10971 Iout.n928 VGND 0.08346f
C10972 Iout.n929 VGND 0.50694f
C10973 Iout.n930 VGND 0.04879f
C10974 Iout.t201 VGND 0.02354f
C10975 Iout.n931 VGND 0.05236f
C10976 Iout.n932 VGND 0.02663f
C10977 Iout.n933 VGND 0.04879f
C10978 Iout.t207 VGND 0.02354f
C10979 Iout.n934 VGND 0.05236f
C10980 Iout.n935 VGND 0.20684f
C10981 Iout.n936 VGND 2.70928f
C10982 Iout.n937 VGND 1.27854f
C10983 Iout.t97 VGND 0.02354f
C10984 Iout.n938 VGND 0.05236f
C10985 Iout.n939 VGND 0.20684f
C10986 Iout.n940 VGND 0.04879f
C10987 Iout.n941 VGND 0.24452f
C10988 Iout.n942 VGND 0.24452f
C10989 Iout.n943 VGND 0.04879f
C10990 Iout.t5 VGND 0.02354f
C10991 Iout.n944 VGND 0.05236f
C10992 Iout.n945 VGND 0.02663f
C10993 Iout.n946 VGND 0.04879f
C10994 Iout.n947 VGND 0.24452f
C10995 Iout.n948 VGND 0.24452f
C10996 Iout.n949 VGND 0.04879f
C10997 Iout.t243 VGND 0.02354f
C10998 Iout.n950 VGND 0.05236f
C10999 Iout.n951 VGND 0.02663f
C11000 Iout.n952 VGND 0.04879f
C11001 Iout.t74 VGND 0.02354f
C11002 Iout.n953 VGND 0.05236f
C11003 Iout.n954 VGND 0.20684f
C11004 Iout.n955 VGND 1.27854f
C11005 Iout.n956 VGND 1.27854f
C11006 Iout.t102 VGND 0.02354f
C11007 Iout.n957 VGND 0.05236f
C11008 Iout.n958 VGND 0.20684f
C11009 Iout.n959 VGND 0.04879f
C11010 Iout.n960 VGND 0.24452f
C11011 Iout.n961 VGND 0.24452f
C11012 Iout.n962 VGND 0.04879f
C11013 Iout.t111 VGND 0.02354f
C11014 Iout.n963 VGND 0.05236f
C11015 Iout.n964 VGND 0.02663f
C11016 Iout.n965 VGND 0.04879f
C11017 Iout.n966 VGND 0.24452f
C11018 Iout.n967 VGND 0.24452f
C11019 Iout.n968 VGND 0.04879f
C11020 Iout.t96 VGND 0.02354f
C11021 Iout.n969 VGND 0.05236f
C11022 Iout.n970 VGND 0.02663f
C11023 Iout.n971 VGND 0.04879f
C11024 Iout.t24 VGND 0.02354f
C11025 Iout.n972 VGND 0.05236f
C11026 Iout.n973 VGND 0.20684f
C11027 Iout.n974 VGND 1.27854f
C11028 Iout.n975 VGND 1.27854f
C11029 Iout.t177 VGND 0.02354f
C11030 Iout.n976 VGND 0.05236f
C11031 Iout.n977 VGND 0.20684f
C11032 Iout.n978 VGND 0.04879f
C11033 Iout.n979 VGND 0.24452f
C11034 Iout.n980 VGND 0.24452f
C11035 Iout.n981 VGND 0.04879f
C11036 Iout.t245 VGND 0.02354f
C11037 Iout.n982 VGND 0.05236f
C11038 Iout.n983 VGND 0.02663f
C11039 Iout.n984 VGND 0.04879f
C11040 Iout.n985 VGND 0.24452f
C11041 Iout.n986 VGND 0.24452f
C11042 Iout.n987 VGND 0.04879f
C11043 Iout.t253 VGND 0.02354f
C11044 Iout.n988 VGND 0.05236f
C11045 Iout.n989 VGND 0.02663f
C11046 Iout.n990 VGND 0.04879f
C11047 Iout.t133 VGND 0.02354f
C11048 Iout.n991 VGND 0.05236f
C11049 Iout.n992 VGND 0.20684f
C11050 Iout.n993 VGND 1.27854f
C11051 Iout.n994 VGND 1.27854f
C11052 Iout.t127 VGND 0.02354f
C11053 Iout.n995 VGND 0.05236f
C11054 Iout.n996 VGND 0.20684f
C11055 Iout.n997 VGND 0.04879f
C11056 Iout.n998 VGND 0.24452f
C11057 Iout.n999 VGND 0.24452f
C11058 Iout.n1000 VGND 0.04879f
C11059 Iout.t9 VGND 0.02354f
C11060 Iout.n1001 VGND 0.05236f
C11061 Iout.n1002 VGND 0.02663f
C11062 Iout.n1003 VGND 0.04879f
C11063 Iout.n1004 VGND 0.24452f
C11064 Iout.n1005 VGND 0.24452f
C11065 Iout.n1006 VGND 0.04879f
C11066 Iout.t66 VGND 0.02354f
C11067 Iout.n1007 VGND 0.05236f
C11068 Iout.n1008 VGND 0.02663f
C11069 Iout.n1009 VGND 0.04879f
C11070 Iout.t176 VGND 0.02354f
C11071 Iout.n1010 VGND 0.05236f
C11072 Iout.n1011 VGND 0.20684f
C11073 Iout.n1012 VGND 1.27854f
C11074 Iout.n1013 VGND 1.14803f
C11075 Iout.t220 VGND 0.02354f
C11076 Iout.n1014 VGND 0.05236f
C11077 Iout.n1015 VGND 0.20684f
C11078 Iout.n1016 VGND 0.04879f
C11079 Iout.n1017 VGND 0.24452f
C11080 Iout.n1018 VGND 0.14435f
C11081 Iout.n1019 VGND 0.04879f
C11082 Iout.t72 VGND 0.02354f
C11083 Iout.n1020 VGND 0.05236f
C11084 Iout.n1021 VGND 0.20684f
C11085 Iout.n1022 VGND 0.23752f
C11086 VPWR.n0 VGND 0.03811f
C11087 VPWR.t831 VGND 0.24101f
C11088 VPWR.t555 VGND 0.10665f
C11089 VPWR.t229 VGND 0.30749f
C11090 VPWR.t1752 VGND 0.11635f
C11091 VPWR.t341 VGND 0.11635f
C11092 VPWR.t338 VGND 0.11635f
C11093 VPWR.t694 VGND 0.11635f
C11094 VPWR.t1734 VGND 0.11635f
C11095 VPWR.t1730 VGND 0.11635f
C11096 VPWR.t784 VGND 0.08172f
C11097 VPWR.n1 VGND 0.14848f
C11098 VPWR.n2 VGND 0.07856f
C11099 VPWR.t556 VGND 0.04648f
C11100 VPWR.t785 VGND 0.01165f
C11101 VPWR.t1731 VGND 0.01165f
C11102 VPWR.n4 VGND 0.02558f
C11103 VPWR.t1735 VGND 0.01165f
C11104 VPWR.t695 VGND 0.01165f
C11105 VPWR.n5 VGND 0.02554f
C11106 VPWR.n6 VGND 0.05245f
C11107 VPWR.n7 VGND 0.14784f
C11108 VPWR.n8 VGND 0.04681f
C11109 VPWR.n9 VGND 0.03438f
C11110 VPWR.n10 VGND 0.06162f
C11111 VPWR.n12 VGND 0.01326f
C11112 VPWR.n13 VGND 0.01553f
C11113 VPWR.n14 VGND 0.02278f
C11114 VPWR.n15 VGND 0.06897f
C11115 VPWR.t832 VGND 0.04646f
C11116 VPWR.n17 VGND 0.05976f
C11117 VPWR.n18 VGND 0.27291f
C11118 VPWR.n19 VGND 0.79581f
C11119 VPWR.n20 VGND 0.87881f
C11120 VPWR.n21 VGND 0.09629f
C11121 VPWR.n22 VGND 0.07371f
C11122 VPWR.n23 VGND 0.13453f
C11123 VPWR.n24 VGND 0.08754f
C11124 VPWR.n25 VGND 0.08514f
C11125 VPWR.n26 VGND 0.0998f
C11126 VPWR.t799 VGND 0.03926f
C11127 VPWR.n27 VGND 0.14793f
C11128 VPWR.n28 VGND 0.14793f
C11129 VPWR.t798 VGND 1.04272f
C11130 VPWR.n29 VGND 0.14793f
C11131 VPWR.n30 VGND 0.14793f
C11132 VPWR.n31 VGND 0.08792f
C11133 VPWR.t1711 VGND 0.03926f
C11134 VPWR.t223 VGND 0.011f
C11135 VPWR.t1032 VGND 0.011f
C11136 VPWR.n32 VGND 0.02201f
C11137 VPWR.n33 VGND 0.01833f
C11138 VPWR.n34 VGND 0.01817f
C11139 VPWR.n35 VGND 0.08754f
C11140 VPWR.n36 VGND 0.19403f
C11141 VPWR.n37 VGND 0.78459f
C11142 VPWR.n38 VGND 1.17383f
C11143 VPWR.n39 VGND 0.25904f
C11144 VPWR.n40 VGND 0.82597f
C11145 VPWR.n41 VGND 0.30027f
C11146 VPWR.n42 VGND 0.05635f
C11147 VPWR.t1223 VGND 0.02709f
C11148 VPWR.t1331 VGND 0.02407f
C11149 VPWR.n43 VGND 0.07442f
C11150 VPWR.t1091 VGND 0.07496f
C11151 VPWR.t1098 VGND 0.02709f
C11152 VPWR.t1092 VGND 0.02407f
C11153 VPWR.n44 VGND 0.07442f
C11154 VPWR.n45 VGND 0.05649f
C11155 VPWR.n46 VGND 0.30049f
C11156 VPWR.n47 VGND 0.30049f
C11157 VPWR.n48 VGND 0.05649f
C11158 VPWR.t1079 VGND 0.02709f
C11159 VPWR.t1452 VGND 0.02407f
C11160 VPWR.n49 VGND 0.07442f
C11161 VPWR.t1318 VGND 0.07496f
C11162 VPWR.t1229 VGND 0.02709f
C11163 VPWR.t1319 VGND 0.02407f
C11164 VPWR.n50 VGND 0.07442f
C11165 VPWR.n51 VGND 0.05649f
C11166 VPWR.n52 VGND 0.30049f
C11167 VPWR.n53 VGND 0.30049f
C11168 VPWR.n54 VGND 0.05649f
C11169 VPWR.t1199 VGND 0.02709f
C11170 VPWR.t1191 VGND 0.02407f
C11171 VPWR.n55 VGND 0.07442f
C11172 VPWR.t1172 VGND 0.07496f
C11173 VPWR.t1455 VGND 0.02709f
C11174 VPWR.t1173 VGND 0.02407f
C11175 VPWR.n56 VGND 0.07442f
C11176 VPWR.n57 VGND 0.05649f
C11177 VPWR.n58 VGND 0.30049f
C11178 VPWR.n59 VGND 0.30049f
C11179 VPWR.n60 VGND 0.05649f
C11180 VPWR.t1328 VGND 0.02709f
C11181 VPWR.t1367 VGND 0.02407f
C11182 VPWR.n61 VGND 0.07442f
C11183 VPWR.t1295 VGND 0.07496f
C11184 VPWR.t1309 VGND 0.02709f
C11185 VPWR.t1296 VGND 0.02407f
C11186 VPWR.n62 VGND 0.07442f
C11187 VPWR.n63 VGND 0.05649f
C11188 VPWR.n64 VGND 0.30049f
C11189 VPWR.n65 VGND 0.30049f
C11190 VPWR.n66 VGND 0.05649f
C11191 VPWR.t1149 VGND 0.02709f
C11192 VPWR.t1168 VGND 0.02407f
C11193 VPWR.n67 VGND 0.07442f
C11194 VPWR.t1132 VGND 0.07496f
C11195 VPWR.t1428 VGND 0.02709f
C11196 VPWR.t1133 VGND 0.02407f
C11197 VPWR.n68 VGND 0.07442f
C11198 VPWR.n69 VGND 0.05649f
C11199 VPWR.n70 VGND 0.30049f
C11200 VPWR.n71 VGND 0.30049f
C11201 VPWR.n72 VGND 0.05649f
C11202 VPWR.t1272 VGND 0.02709f
C11203 VPWR.t1415 VGND 0.02407f
C11204 VPWR.n73 VGND 0.07442f
C11205 VPWR.t1253 VGND 0.07496f
C11206 VPWR.t1260 VGND 0.02709f
C11207 VPWR.t1254 VGND 0.02407f
C11208 VPWR.n74 VGND 0.07442f
C11209 VPWR.n75 VGND 0.05649f
C11210 VPWR.n76 VGND 0.30049f
C11211 VPWR.n77 VGND 0.30049f
C11212 VPWR.n78 VGND 0.05649f
C11213 VPWR.t1152 VGND 0.02709f
C11214 VPWR.t1146 VGND 0.02407f
C11215 VPWR.n79 VGND 0.07442f
C11216 VPWR.t1380 VGND 0.07496f
C11217 VPWR.t1396 VGND 0.02709f
C11218 VPWR.t1381 VGND 0.02407f
C11219 VPWR.n80 VGND 0.07442f
C11220 VPWR.n81 VGND 0.05649f
C11221 VPWR.n82 VGND 0.30049f
C11222 VPWR.n83 VGND 0.30049f
C11223 VPWR.n84 VGND 0.05649f
C11224 VPWR.t1275 VGND 0.02709f
C11225 VPWR.t1375 VGND 0.02407f
C11226 VPWR.n85 VGND 0.07442f
C11227 VPWR.t1129 VGND 0.118f
C11228 VPWR.t1105 VGND 0.06383f
C11229 VPWR.t1236 VGND 0.07496f
C11230 VPWR.t1130 VGND 0.02709f
C11231 VPWR.t1237 VGND 0.02407f
C11232 VPWR.n86 VGND 0.07442f
C11233 VPWR.n87 VGND 0.02434f
C11234 VPWR.n88 VGND 0.0267f
C11235 VPWR.n90 VGND 0.01481f
C11236 VPWR.n91 VGND 0.02434f
C11237 VPWR.n92 VGND 0.0267f
C11238 VPWR.n93 VGND 0.02533f
C11239 VPWR.n94 VGND 0.01601f
C11240 VPWR.t1104 VGND 0.01009f
C11241 VPWR.n95 VGND 0.02251f
C11242 VPWR.n96 VGND 0.02292f
C11243 VPWR.n97 VGND 0.01444f
C11244 VPWR.n99 VGND 0.01481f
C11245 VPWR.n100 VGND 0.02158f
C11246 VPWR.n101 VGND 0.14299f
C11247 VPWR.n102 VGND 0.02434f
C11248 VPWR.n103 VGND 0.0267f
C11249 VPWR.n105 VGND 0.01481f
C11250 VPWR.n106 VGND 0.14299f
C11251 VPWR.n107 VGND 0.02434f
C11252 VPWR.n108 VGND 0.0267f
C11253 VPWR.n110 VGND 0.01481f
C11254 VPWR.n111 VGND 0.14299f
C11255 VPWR.n112 VGND 0.02434f
C11256 VPWR.n113 VGND 0.0267f
C11257 VPWR.n115 VGND 0.01481f
C11258 VPWR.n116 VGND 0.14299f
C11259 VPWR.n117 VGND 0.02434f
C11260 VPWR.n118 VGND 0.0267f
C11261 VPWR.n120 VGND 0.01481f
C11262 VPWR.n121 VGND 0.02066f
C11263 VPWR.n122 VGND 0.02434f
C11264 VPWR.n123 VGND 0.0267f
C11265 VPWR.n124 VGND 0.01481f
C11266 VPWR.n126 VGND 0.01444f
C11267 VPWR.t1205 VGND 0.01009f
C11268 VPWR.n127 VGND 0.02251f
C11269 VPWR.n128 VGND 0.02292f
C11270 VPWR.n130 VGND 0.02533f
C11271 VPWR.n131 VGND 0.03003f
C11272 VPWR.n132 VGND 0.02774f
C11273 VPWR.n133 VGND 0.02434f
C11274 VPWR.n134 VGND 0.0267f
C11275 VPWR.n135 VGND 0.02774f
C11276 VPWR.n136 VGND 0.02533f
C11277 VPWR.n137 VGND 0.03003f
C11278 VPWR.t1354 VGND 0.01009f
C11279 VPWR.n139 VGND 0.02251f
C11280 VPWR.n140 VGND 0.02292f
C11281 VPWR.n141 VGND 0.01444f
C11282 VPWR.n143 VGND 0.01481f
C11283 VPWR.n144 VGND 0.01938f
C11284 VPWR.n145 VGND 0.17208f
C11285 VPWR.n146 VGND 0.14299f
C11286 VPWR.n147 VGND 0.01938f
C11287 VPWR.n148 VGND 0.01444f
C11288 VPWR.t1332 VGND 0.01009f
C11289 VPWR.n149 VGND 0.02251f
C11290 VPWR.n150 VGND 0.02292f
C11291 VPWR.n152 VGND 0.02533f
C11292 VPWR.n153 VGND 0.03003f
C11293 VPWR.n154 VGND 0.02774f
C11294 VPWR.n155 VGND 0.02434f
C11295 VPWR.n156 VGND 0.0267f
C11296 VPWR.n158 VGND 0.01481f
C11297 VPWR.n159 VGND 0.01938f
C11298 VPWR.n160 VGND 0.01444f
C11299 VPWR.t1310 VGND 0.01009f
C11300 VPWR.n161 VGND 0.02251f
C11301 VPWR.n162 VGND 0.02292f
C11302 VPWR.n164 VGND 0.02533f
C11303 VPWR.n165 VGND 0.03003f
C11304 VPWR.n166 VGND 0.02774f
C11305 VPWR.n167 VGND 0.02434f
C11306 VPWR.n168 VGND 0.0267f
C11307 VPWR.n169 VGND 0.02774f
C11308 VPWR.n170 VGND 0.02533f
C11309 VPWR.n171 VGND 0.03003f
C11310 VPWR.t1456 VGND 0.01009f
C11311 VPWR.n173 VGND 0.02251f
C11312 VPWR.n174 VGND 0.02292f
C11313 VPWR.n175 VGND 0.01444f
C11314 VPWR.n177 VGND 0.01481f
C11315 VPWR.n178 VGND 0.01938f
C11316 VPWR.n179 VGND 0.14299f
C11317 VPWR.n180 VGND 0.14299f
C11318 VPWR.n181 VGND 0.01938f
C11319 VPWR.n182 VGND 0.01444f
C11320 VPWR.t1437 VGND 0.01009f
C11321 VPWR.n183 VGND 0.02251f
C11322 VPWR.n184 VGND 0.02292f
C11323 VPWR.n186 VGND 0.02533f
C11324 VPWR.n187 VGND 0.03003f
C11325 VPWR.n188 VGND 0.02774f
C11326 VPWR.n189 VGND 0.02434f
C11327 VPWR.n190 VGND 0.0267f
C11328 VPWR.n192 VGND 0.01481f
C11329 VPWR.n193 VGND 0.01938f
C11330 VPWR.n194 VGND 0.01444f
C11331 VPWR.t1276 VGND 0.01009f
C11332 VPWR.n195 VGND 0.02251f
C11333 VPWR.n196 VGND 0.02292f
C11334 VPWR.n198 VGND 0.02533f
C11335 VPWR.n199 VGND 0.03003f
C11336 VPWR.n200 VGND 0.02774f
C11337 VPWR.n201 VGND 0.02434f
C11338 VPWR.n202 VGND 0.0267f
C11339 VPWR.n203 VGND 0.02774f
C11340 VPWR.n204 VGND 0.02533f
C11341 VPWR.n205 VGND 0.03003f
C11342 VPWR.t1174 VGND 0.01009f
C11343 VPWR.n207 VGND 0.02251f
C11344 VPWR.n208 VGND 0.02292f
C11345 VPWR.n209 VGND 0.01444f
C11346 VPWR.n211 VGND 0.01481f
C11347 VPWR.n212 VGND 0.01938f
C11348 VPWR.n213 VGND 0.14299f
C11349 VPWR.n214 VGND 0.14299f
C11350 VPWR.n215 VGND 0.01938f
C11351 VPWR.n216 VGND 0.01444f
C11352 VPWR.t1139 VGND 0.01009f
C11353 VPWR.n217 VGND 0.02251f
C11354 VPWR.n218 VGND 0.02292f
C11355 VPWR.n220 VGND 0.02533f
C11356 VPWR.n221 VGND 0.03003f
C11357 VPWR.n222 VGND 0.02774f
C11358 VPWR.n223 VGND 0.02434f
C11359 VPWR.n224 VGND 0.0267f
C11360 VPWR.n226 VGND 0.01481f
C11361 VPWR.n227 VGND 0.01938f
C11362 VPWR.n228 VGND 0.01444f
C11363 VPWR.t1302 VGND 0.01009f
C11364 VPWR.n229 VGND 0.02251f
C11365 VPWR.n230 VGND 0.02292f
C11366 VPWR.n232 VGND 0.02533f
C11367 VPWR.n233 VGND 0.03003f
C11368 VPWR.n234 VGND 0.02774f
C11369 VPWR.n235 VGND 0.02434f
C11370 VPWR.n236 VGND 0.0267f
C11371 VPWR.n237 VGND 0.02774f
C11372 VPWR.n238 VGND 0.02533f
C11373 VPWR.n239 VGND 0.03003f
C11374 VPWR.t1278 VGND 0.01009f
C11375 VPWR.n241 VGND 0.02251f
C11376 VPWR.n242 VGND 0.02292f
C11377 VPWR.n243 VGND 0.01444f
C11378 VPWR.n245 VGND 0.01481f
C11379 VPWR.n246 VGND 0.01938f
C11380 VPWR.n247 VGND 0.14299f
C11381 VPWR.n248 VGND 0.14299f
C11382 VPWR.n249 VGND 0.01938f
C11383 VPWR.n250 VGND 0.01444f
C11384 VPWR.t1134 VGND 0.01009f
C11385 VPWR.n251 VGND 0.02251f
C11386 VPWR.n252 VGND 0.02292f
C11387 VPWR.n254 VGND 0.02533f
C11388 VPWR.n255 VGND 0.03003f
C11389 VPWR.n256 VGND 0.02774f
C11390 VPWR.n257 VGND 0.02434f
C11391 VPWR.n258 VGND 0.0267f
C11392 VPWR.n260 VGND 0.01481f
C11393 VPWR.n261 VGND 0.01938f
C11394 VPWR.n262 VGND 0.01444f
C11395 VPWR.t1416 VGND 0.01009f
C11396 VPWR.n263 VGND 0.02251f
C11397 VPWR.n264 VGND 0.02292f
C11398 VPWR.n266 VGND 0.02533f
C11399 VPWR.n267 VGND 0.03003f
C11400 VPWR.n268 VGND 0.02774f
C11401 VPWR.n269 VGND 0.02434f
C11402 VPWR.n270 VGND 0.0267f
C11403 VPWR.n271 VGND 0.02774f
C11404 VPWR.n272 VGND 0.02533f
C11405 VPWR.n273 VGND 0.03003f
C11406 VPWR.t1382 VGND 0.01009f
C11407 VPWR.n275 VGND 0.02251f
C11408 VPWR.n276 VGND 0.02292f
C11409 VPWR.n277 VGND 0.01444f
C11410 VPWR.n279 VGND 0.01481f
C11411 VPWR.n280 VGND 0.01938f
C11412 VPWR.n281 VGND 0.14299f
C11413 VPWR.n282 VGND 0.19291f
C11414 VPWR.n283 VGND 0.01938f
C11415 VPWR.n284 VGND 0.01444f
C11416 VPWR.t1240 VGND 0.01009f
C11417 VPWR.n285 VGND 0.02251f
C11418 VPWR.n286 VGND 0.02292f
C11419 VPWR.n288 VGND 0.02533f
C11420 VPWR.n289 VGND 0.03003f
C11421 VPWR.n290 VGND 0.02764f
C11422 VPWR.t608 VGND 0.02709f
C11423 VPWR.t488 VGND 0.02407f
C11424 VPWR.n291 VGND 0.07442f
C11425 VPWR.t1694 VGND 0.02709f
C11426 VPWR.t507 VGND 0.02407f
C11427 VPWR.n294 VGND 0.07442f
C11428 VPWR.t607 VGND 0.118f
C11429 VPWR.t736 VGND 0.06383f
C11430 VPWR.t487 VGND 0.07496f
C11431 VPWR.n295 VGND 0.088f
C11432 VPWR.t1693 VGND 0.09722f
C11433 VPWR.t624 VGND 0.06383f
C11434 VPWR.t506 VGND 0.07496f
C11435 VPWR.t1512 VGND 0.09722f
C11436 VPWR.t257 VGND 0.02709f
C11437 VPWR.t1489 VGND 0.02407f
C11438 VPWR.n296 VGND 0.07442f
C11439 VPWR.t1513 VGND 0.02709f
C11440 VPWR.t813 VGND 0.02407f
C11441 VPWR.n298 VGND 0.07442f
C11442 VPWR.t739 VGND 0.06383f
C11443 VPWR.t812 VGND 0.07496f
C11444 VPWR.t500 VGND 0.09722f
C11445 VPWR.t1065 VGND 0.02709f
C11446 VPWR.t1778 VGND 0.02407f
C11447 VPWR.n299 VGND 0.07442f
C11448 VPWR.t501 VGND 0.02709f
C11449 VPWR.t431 VGND 0.02407f
C11450 VPWR.n301 VGND 0.07442f
C11451 VPWR.t1921 VGND 0.06383f
C11452 VPWR.t430 VGND 0.07496f
C11453 VPWR.t70 VGND 0.09722f
C11454 VPWR.t1884 VGND 0.02709f
C11455 VPWR.t77 VGND 0.02407f
C11456 VPWR.n302 VGND 0.07442f
C11457 VPWR.t71 VGND 0.02709f
C11458 VPWR.t811 VGND 0.02407f
C11459 VPWR.n304 VGND 0.07442f
C11460 VPWR.t627 VGND 0.06383f
C11461 VPWR.t810 VGND 0.07496f
C11462 VPWR.t1038 VGND 0.09722f
C11463 VPWR.t871 VGND 0.02709f
C11464 VPWR.t1045 VGND 0.02407f
C11465 VPWR.n305 VGND 0.07442f
C11466 VPWR.t1039 VGND 0.02709f
C11467 VPWR.t1555 VGND 0.02407f
C11468 VPWR.n307 VGND 0.07442f
C11469 VPWR.t623 VGND 0.06383f
C11470 VPWR.t1554 VGND 0.07496f
C11471 VPWR.t1010 VGND 0.09722f
C11472 VPWR.t304 VGND 0.02709f
C11473 VPWR.t1017 VGND 0.02407f
C11474 VPWR.n308 VGND 0.07442f
C11475 VPWR.t1011 VGND 0.02709f
C11476 VPWR.t1829 VGND 0.02407f
C11477 VPWR.n310 VGND 0.07442f
C11478 VPWR.t737 VGND 0.06383f
C11479 VPWR.t1828 VGND 0.07496f
C11480 VPWR.t206 VGND 0.09722f
C11481 VPWR.t905 VGND 0.02709f
C11482 VPWR.t1471 VGND 0.02407f
C11483 VPWR.n311 VGND 0.07442f
C11484 VPWR.t207 VGND 0.02709f
C11485 VPWR.t1640 VGND 0.02407f
C11486 VPWR.n313 VGND 0.07442f
C11487 VPWR.t1918 VGND 0.06383f
C11488 VPWR.t1639 VGND 0.07496f
C11489 VPWR.t994 VGND 0.09722f
C11490 VPWR.t972 VGND 0.02709f
C11491 VPWR.t1715 VGND 0.02407f
C11492 VPWR.n314 VGND 0.07442f
C11493 VPWR.t995 VGND 0.02709f
C11494 VPWR.t1436 VGND 0.02407f
C11495 VPWR.n316 VGND 0.07442f
C11496 VPWR.t625 VGND 0.06383f
C11497 VPWR.t1435 VGND 0.10842f
C11498 VPWR.n317 VGND 0.06192f
C11499 VPWR.n318 VGND 0.0512f
C11500 VPWR.n320 VGND 0.0512f
C11501 VPWR.n322 VGND 0.088f
C11502 VPWR.t1714 VGND 0.07496f
C11503 VPWR.t1076 VGND 0.06383f
C11504 VPWR.t971 VGND 0.09722f
C11505 VPWR.n323 VGND 0.088f
C11506 VPWR.n325 VGND 0.0512f
C11507 VPWR.n327 VGND 0.0512f
C11508 VPWR.n329 VGND 0.088f
C11509 VPWR.t1470 VGND 0.07496f
C11510 VPWR.t1919 VGND 0.06383f
C11511 VPWR.t904 VGND 0.09722f
C11512 VPWR.n330 VGND 0.088f
C11513 VPWR.n332 VGND 0.0512f
C11514 VPWR.n334 VGND 0.0512f
C11515 VPWR.n336 VGND 0.088f
C11516 VPWR.t1016 VGND 0.07496f
C11517 VPWR.t738 VGND 0.06383f
C11518 VPWR.t303 VGND 0.09722f
C11519 VPWR.n337 VGND 0.088f
C11520 VPWR.n339 VGND 0.0512f
C11521 VPWR.n341 VGND 0.0512f
C11522 VPWR.n343 VGND 0.088f
C11523 VPWR.t1044 VGND 0.07496f
C11524 VPWR.t626 VGND 0.06383f
C11525 VPWR.t870 VGND 0.09722f
C11526 VPWR.n344 VGND 0.088f
C11527 VPWR.n346 VGND 0.0512f
C11528 VPWR.n348 VGND 0.0512f
C11529 VPWR.n350 VGND 0.088f
C11530 VPWR.t76 VGND 0.07496f
C11531 VPWR.t1920 VGND 0.06383f
C11532 VPWR.t1883 VGND 0.09722f
C11533 VPWR.n351 VGND 0.088f
C11534 VPWR.n353 VGND 0.0512f
C11535 VPWR.n355 VGND 0.0512f
C11536 VPWR.n357 VGND 0.088f
C11537 VPWR.t1777 VGND 0.07496f
C11538 VPWR.t628 VGND 0.06383f
C11539 VPWR.t1064 VGND 0.09722f
C11540 VPWR.n358 VGND 0.088f
C11541 VPWR.n360 VGND 0.0512f
C11542 VPWR.n362 VGND 0.0512f
C11543 VPWR.n364 VGND 0.088f
C11544 VPWR.t1488 VGND 0.07496f
C11545 VPWR.t740 VGND 0.06383f
C11546 VPWR.t256 VGND 0.09722f
C11547 VPWR.n365 VGND 0.088f
C11548 VPWR.n367 VGND 0.0512f
C11549 VPWR.n368 VGND -0.05607f
C11550 VPWR.n369 VGND 0.30049f
C11551 VPWR.n370 VGND 0.82079f
C11552 VPWR.n371 VGND 0.2969f
C11553 VPWR.t602 VGND 0.02709f
C11554 VPWR.t494 VGND 0.02407f
C11555 VPWR.n372 VGND 0.07442f
C11556 VPWR.t484 VGND 0.02709f
C11557 VPWR.t452 VGND 0.02407f
C11558 VPWR.n375 VGND 0.07442f
C11559 VPWR.t601 VGND 0.118f
C11560 VPWR.t935 VGND 0.06383f
C11561 VPWR.t493 VGND 0.07496f
C11562 VPWR.n376 VGND 0.088f
C11563 VPWR.t483 VGND 0.09722f
C11564 VPWR.t1762 VGND 0.06383f
C11565 VPWR.t451 VGND 0.07496f
C11566 VPWR.t1504 VGND 0.09722f
C11567 VPWR.t511 VGND 0.02709f
C11568 VPWR.t1481 VGND 0.02407f
C11569 VPWR.n377 VGND 0.07442f
C11570 VPWR.n378 VGND 0.2969f
C11571 VPWR.n379 VGND 0.2969f
C11572 VPWR.n380 VGND 0.0512f
C11573 VPWR.t1073 VGND 0.02709f
C11574 VPWR.t1667 VGND 0.02407f
C11575 VPWR.n382 VGND 0.07442f
C11576 VPWR.t1757 VGND 0.06383f
C11577 VPWR.t824 VGND 0.07496f
C11578 VPWR.t1505 VGND 0.02709f
C11579 VPWR.t825 VGND 0.02407f
C11580 VPWR.n383 VGND 0.07442f
C11581 VPWR.n385 VGND 0.088f
C11582 VPWR.t1072 VGND 0.09722f
C11583 VPWR.t934 VGND 0.06383f
C11584 VPWR.t1666 VGND 0.07496f
C11585 VPWR.t434 VGND 0.09722f
C11586 VPWR.t1782 VGND 0.02709f
C11587 VPWR.t913 VGND 0.02407f
C11588 VPWR.n386 VGND 0.07442f
C11589 VPWR.n387 VGND 0.2969f
C11590 VPWR.n388 VGND 0.2969f
C11591 VPWR.n389 VGND 0.0512f
C11592 VPWR.t81 VGND 0.02709f
C11593 VPWR.t63 VGND 0.02407f
C11594 VPWR.n391 VGND 0.07442f
C11595 VPWR.t1739 VGND 0.06383f
C11596 VPWR.t1833 VGND 0.07496f
C11597 VPWR.t435 VGND 0.02709f
C11598 VPWR.t1834 VGND 0.02407f
C11599 VPWR.n392 VGND 0.07442f
C11600 VPWR.n394 VGND 0.088f
C11601 VPWR.t80 VGND 0.09722f
C11602 VPWR.t933 VGND 0.06383f
C11603 VPWR.t62 VGND 0.07496f
C11604 VPWR.t889 VGND 0.09722f
C11605 VPWR.t722 VGND 0.02709f
C11606 VPWR.t896 VGND 0.02407f
C11607 VPWR.n395 VGND 0.07442f
C11608 VPWR.n396 VGND 0.2969f
C11609 VPWR.n397 VGND 0.2969f
C11610 VPWR.n398 VGND 0.0512f
C11611 VPWR.t310 VGND 0.02709f
C11612 VPWR.t178 VGND 0.02407f
C11613 VPWR.n400 VGND 0.07442f
C11614 VPWR.t1741 VGND 0.06383f
C11615 VPWR.t1560 VGND 0.07496f
C11616 VPWR.t890 VGND 0.02709f
C11617 VPWR.t1561 VGND 0.02407f
C11618 VPWR.n401 VGND 0.07442f
C11619 VPWR.n403 VGND 0.088f
C11620 VPWR.t309 VGND 0.09722f
C11621 VPWR.t1756 VGND 0.06383f
C11622 VPWR.t177 VGND 0.07496f
C11623 VPWR.t1824 VGND 0.09722f
C11624 VPWR.t1021 VGND 0.02709f
C11625 VPWR.t96 VGND 0.02407f
C11626 VPWR.n404 VGND 0.07442f
C11627 VPWR.n405 VGND 0.2969f
C11628 VPWR.n406 VGND 0.2969f
C11629 VPWR.n407 VGND 0.0512f
C11630 VPWR.t213 VGND 0.02709f
C11631 VPWR.t119 VGND 0.02407f
C11632 VPWR.n409 VGND 0.07442f
C11633 VPWR.t1738 VGND 0.06383f
C11634 VPWR.t183 VGND 0.07496f
C11635 VPWR.t1825 VGND 0.02709f
C11636 VPWR.t184 VGND 0.02407f
C11637 VPWR.n410 VGND 0.07442f
C11638 VPWR.n412 VGND 0.088f
C11639 VPWR.t212 VGND 0.09722f
C11640 VPWR.t1737 VGND 0.06383f
C11641 VPWR.t118 VGND 0.07496f
C11642 VPWR.t1002 VGND 0.09722f
C11643 VPWR.t1636 VGND 0.02709f
C11644 VPWR.t1727 VGND 0.02407f
C11645 VPWR.n413 VGND 0.07442f
C11646 VPWR.n414 VGND 0.2969f
C11647 VPWR.n415 VGND 0.82597f
C11648 VPWR.n416 VGND 0.2969f
C11649 VPWR.n418 VGND 0.82597f
C11650 VPWR.n419 VGND 0.2969f
C11651 VPWR.n420 VGND 0.0512f
C11652 VPWR.t583 VGND 0.02709f
C11653 VPWR.t1226 VGND 0.02407f
C11654 VPWR.n422 VGND 0.07442f
C11655 VPWR.t24 VGND 0.07496f
C11656 VPWR.t190 VGND 0.02709f
C11657 VPWR.t25 VGND 0.02407f
C11658 VPWR.n423 VGND 0.07442f
C11659 VPWR.n424 VGND 0.2969f
C11660 VPWR.n425 VGND 0.06791f
C11661 VPWR.n426 VGND 0.2969f
C11662 VPWR.n427 VGND 0.2969f
C11663 VPWR.n428 VGND 0.2969f
C11664 VPWR.t1601 VGND 0.02709f
C11665 VPWR.t1061 VGND 0.02407f
C11666 VPWR.n429 VGND 0.07442f
C11667 VPWR.t1814 VGND 0.07496f
C11668 VPWR.t1578 VGND 0.02709f
C11669 VPWR.t1815 VGND 0.02407f
C11670 VPWR.n430 VGND 0.07442f
C11671 VPWR.n431 VGND 0.2969f
C11672 VPWR.n432 VGND 0.2969f
C11673 VPWR.n435 VGND 0.06791f
C11674 VPWR.n436 VGND 0.2969f
C11675 VPWR.n437 VGND 0.2969f
C11676 VPWR.n438 VGND 0.06791f
C11677 VPWR.n439 VGND 0.2969f
C11678 VPWR.n440 VGND 0.0512f
C11679 VPWR.t1 VGND 0.02709f
C11680 VPWR.t575 VGND 0.02407f
C11681 VPWR.n442 VGND 0.07442f
C11682 VPWR.t475 VGND 0.07496f
C11683 VPWR.t412 VGND 0.02709f
C11684 VPWR.t476 VGND 0.02407f
C11685 VPWR.n443 VGND 0.07442f
C11686 VPWR.t1747 VGND 0.02709f
C11687 VPWR.t1880 VGND 0.02407f
C11688 VPWR.n444 VGND 0.07442f
C11689 VPWR.t1681 VGND 0.07496f
C11690 VPWR.t712 VGND 0.02709f
C11691 VPWR.t1682 VGND 0.02407f
C11692 VPWR.n445 VGND 0.07442f
C11693 VPWR.n446 VGND 0.2969f
C11694 VPWR.n447 VGND 0.06791f
C11695 VPWR.n448 VGND 0.2969f
C11696 VPWR.n449 VGND 0.06791f
C11697 VPWR.n450 VGND 0.2969f
C11698 VPWR.n452 VGND 0.2969f
C11699 VPWR.n453 VGND 0.0512f
C11700 VPWR.t1539 VGND 0.02709f
C11701 VPWR.t714 VGND 0.02407f
C11702 VPWR.n455 VGND 0.07442f
C11703 VPWR.t713 VGND 0.07496f
C11704 VPWR.t161 VGND 0.09722f
C11705 VPWR.t733 VGND 0.02709f
C11706 VPWR.t1698 VGND 0.02407f
C11707 VPWR.n456 VGND 0.07442f
C11708 VPWR.t162 VGND 0.02709f
C11709 VPWR.t1801 VGND 0.02407f
C11710 VPWR.n458 VGND 0.07442f
C11711 VPWR.t102 VGND 0.06383f
C11712 VPWR.t1800 VGND 0.07496f
C11713 VPWR.t481 VGND 0.09722f
C11714 VPWR.t170 VGND 0.02709f
C11715 VPWR.t460 VGND 0.02407f
C11716 VPWR.n459 VGND 0.07442f
C11717 VPWR.n460 VGND 0.2969f
C11718 VPWR.n461 VGND 0.2969f
C11719 VPWR.n462 VGND 0.0512f
C11720 VPWR.n463 VGND 0.2969f
C11721 VPWR.n465 VGND 0.2969f
C11722 VPWR.t993 VGND 0.02709f
C11723 VPWR.t1444 VGND 0.02407f
C11724 VPWR.n466 VGND 0.07442f
C11725 VPWR.t1712 VGND 0.07496f
C11726 VPWR.t970 VGND 0.02709f
C11727 VPWR.t1713 VGND 0.02407f
C11728 VPWR.n467 VGND 0.07442f
C11729 VPWR.t203 VGND 0.02709f
C11730 VPWR.t1638 VGND 0.02407f
C11731 VPWR.n468 VGND 0.07442f
C11732 VPWR.t1466 VGND 0.07496f
C11733 VPWR.t903 VGND 0.02709f
C11734 VPWR.t1467 VGND 0.02407f
C11735 VPWR.n469 VGND 0.07442f
C11736 VPWR.t1009 VGND 0.02709f
C11737 VPWR.t1827 VGND 0.02407f
C11738 VPWR.n470 VGND 0.07442f
C11739 VPWR.t311 VGND 0.07496f
C11740 VPWR.t1574 VGND 0.02709f
C11741 VPWR.t312 VGND 0.02407f
C11742 VPWR.n471 VGND 0.07442f
C11743 VPWR.t867 VGND 0.02709f
C11744 VPWR.t1041 VGND 0.02407f
C11745 VPWR.n472 VGND 0.07442f
C11746 VPWR.t806 VGND 0.07496f
C11747 VPWR.t69 VGND 0.02709f
C11748 VPWR.t807 VGND 0.02407f
C11749 VPWR.n473 VGND 0.07442f
C11750 VPWR.n474 VGND 0.2969f
C11751 VPWR.n475 VGND 0.2969f
C11752 VPWR.n477 VGND 0.2969f
C11753 VPWR.n479 VGND 0.2969f
C11754 VPWR.n480 VGND 0.0512f
C11755 VPWR.t499 VGND 0.02709f
C11756 VPWR.t427 VGND 0.02407f
C11757 VPWR.n481 VGND 0.07442f
C11758 VPWR.t1797 VGND 0.07496f
C11759 VPWR.t1515 VGND 0.02709f
C11760 VPWR.t1798 VGND 0.02407f
C11761 VPWR.n482 VGND 0.07442f
C11762 VPWR.t255 VGND 0.02709f
C11763 VPWR.t1491 VGND 0.02407f
C11764 VPWR.n483 VGND 0.07442f
C11765 VPWR.t502 VGND 0.07496f
C11766 VPWR.t1692 VGND 0.02709f
C11767 VPWR.t503 VGND 0.02407f
C11768 VPWR.n484 VGND 0.07442f
C11769 VPWR.t610 VGND 0.02709f
C11770 VPWR.t486 VGND 0.02407f
C11771 VPWR.n485 VGND 0.07442f
C11772 VPWR.t609 VGND 0.118f
C11773 VPWR.t885 VGND 0.06383f
C11774 VPWR.t485 VGND 0.07496f
C11775 VPWR.t154 VGND 0.06383f
C11776 VPWR.t1691 VGND 0.09722f
C11777 VPWR.n486 VGND 0.088f
C11778 VPWR.n488 VGND 0.2969f
C11779 VPWR.t620 VGND 0.02709f
C11780 VPWR.t245 VGND 0.02407f
C11781 VPWR.n489 VGND 0.07442f
C11782 VPWR.t797 VGND 0.02709f
C11783 VPWR.t773 VGND 0.02407f
C11784 VPWR.n491 VGND 0.07442f
C11785 VPWR.t619 VGND 0.118f
C11786 VPWR.t926 VGND 0.06383f
C11787 VPWR.t244 VGND 0.07496f
C11788 VPWR.n492 VGND 0.088f
C11789 VPWR.t796 VGND 0.09722f
C11790 VPWR.t104 VGND 0.06383f
C11791 VPWR.t772 VGND 0.07496f
C11792 VPWR.t929 VGND 0.06383f
C11793 VPWR.t1538 VGND 0.09722f
C11794 VPWR.t1630 VGND 0.02709f
C11795 VPWR.t1517 VGND 0.02407f
C11796 VPWR.n493 VGND 0.07442f
C11797 VPWR.n495 VGND 0.088f
C11798 VPWR.t1516 VGND 0.07496f
C11799 VPWR.t861 VGND 0.06383f
C11800 VPWR.t1629 VGND 0.09722f
C11801 VPWR.n496 VGND 0.088f
C11802 VPWR.n498 VGND 0.0512f
C11803 VPWR.n499 VGND -0.05607f
C11804 VPWR.n500 VGND 0.2969f
C11805 VPWR.n501 VGND 0.82079f
C11806 VPWR.n502 VGND 0.2969f
C11807 VPWR.n503 VGND 0.0512f
C11808 VPWR.t940 VGND 0.02709f
C11809 VPWR.t1529 VGND 0.02407f
C11810 VPWR.n505 VGND 0.07442f
C11811 VPWR.t595 VGND 0.118f
C11812 VPWR.t1657 VGND 0.06383f
C11813 VPWR.t792 VGND 0.07496f
C11814 VPWR.t596 VGND 0.02709f
C11815 VPWR.t793 VGND 0.02407f
C11816 VPWR.n506 VGND 0.07442f
C11817 VPWR.n507 VGND -0.05607f
C11818 VPWR.n509 VGND 0.088f
C11819 VPWR.t702 VGND 0.09722f
C11820 VPWR.t1652 VGND 0.06383f
C11821 VPWR.t947 VGND 0.07496f
C11822 VPWR.t703 VGND 0.02709f
C11823 VPWR.t948 VGND 0.02407f
C11824 VPWR.n510 VGND 0.07442f
C11825 VPWR.n512 VGND 0.088f
C11826 VPWR.t939 VGND 0.09722f
C11827 VPWR.t328 VGND 0.06383f
C11828 VPWR.t1528 VGND 0.07496f
C11829 VPWR.t820 VGND 0.09722f
C11830 VPWR.t1493 VGND 0.02709f
C11831 VPWR.t1790 VGND 0.02407f
C11832 VPWR.n513 VGND 0.07442f
C11833 VPWR.t821 VGND 0.02709f
C11834 VPWR.t1593 VGND 0.02407f
C11835 VPWR.n515 VGND 0.07442f
C11836 VPWR.t1656 VGND 0.06383f
C11837 VPWR.t1592 VGND 0.07496f
C11838 VPWR.t1851 VGND 0.09722f
C11839 VPWR.t1585 VGND 0.02709f
C11840 VPWR.t164 VGND 0.02407f
C11841 VPWR.n516 VGND 0.07442f
C11842 VPWR.t1852 VGND 0.02709f
C11843 VPWR.t1770 VGND 0.02407f
C11844 VPWR.n518 VGND 0.07442f
C11845 VPWR.t1649 VGND 0.06383f
C11846 VPWR.t1769 VGND 0.07496f
C11847 VPWR.t54 VGND 0.09722f
C11848 VPWR.t1842 VGND 0.02709f
C11849 VPWR.t107 VGND 0.02407f
C11850 VPWR.n519 VGND 0.07442f
C11851 VPWR.t55 VGND 0.02709f
C11852 VPWR.t659 VGND 0.02407f
C11853 VPWR.n521 VGND 0.07442f
C11854 VPWR.t1654 VGND 0.06383f
C11855 VPWR.t658 VGND 0.07496f
C11856 VPWR.t1895 VGND 0.09722f
C11857 VPWR.t671 VGND 0.02709f
C11858 VPWR.t359 VGND 0.02407f
C11859 VPWR.n522 VGND 0.07442f
C11860 VPWR.t1896 VGND 0.02709f
C11861 VPWR.t756 VGND 0.02407f
C11862 VPWR.n524 VGND 0.07442f
C11863 VPWR.t326 VGND 0.06383f
C11864 VPWR.t755 VGND 0.07496f
C11865 VPWR.t1606 VGND 0.09722f
C11866 VPWR.t748 VGND 0.02709f
C11867 VPWR.t1597 VGND 0.02407f
C11868 VPWR.n525 VGND 0.07442f
C11869 VPWR.n526 VGND 0.2969f
C11870 VPWR.n527 VGND 0.2969f
C11871 VPWR.n528 VGND 0.0512f
C11872 VPWR.t1473 VGND 0.02709f
C11873 VPWR.t9 VGND 0.02407f
C11874 VPWR.n530 VGND 0.07442f
C11875 VPWR.t331 VGND 0.06383f
C11876 VPWR.t1048 VGND 0.07496f
C11877 VPWR.t1607 VGND 0.02709f
C11878 VPWR.t1049 VGND 0.02407f
C11879 VPWR.n531 VGND 0.07442f
C11880 VPWR.n533 VGND 0.088f
C11881 VPWR.t1472 VGND 0.09722f
C11882 VPWR.t330 VGND 0.06383f
C11883 VPWR.t8 VGND 0.07496f
C11884 VPWR.t1722 VGND 0.09722f
C11885 VPWR.t1708 VGND 0.02709f
C11886 VPWR.t521 VGND 0.02407f
C11887 VPWR.n534 VGND 0.07442f
C11888 VPWR.t1723 VGND 0.02709f
C11889 VPWR.t1293 VGND 0.02407f
C11890 VPWR.n536 VGND 0.07442f
C11891 VPWR.t1653 VGND 0.06383f
C11892 VPWR.t1292 VGND 0.10842f
C11893 VPWR.n537 VGND 0.06192f
C11894 VPWR.n538 VGND 0.0512f
C11895 VPWR.n539 VGND 0.2969f
C11896 VPWR.n540 VGND 0.82597f
C11897 VPWR.n541 VGND 0.2969f
C11898 VPWR.t999 VGND 0.02709f
C11899 VPWR.t1410 VGND 0.02407f
C11900 VPWR.n542 VGND 0.07442f
C11901 VPWR.t1724 VGND 0.07496f
C11902 VPWR.t1634 VGND 0.02709f
C11903 VPWR.t1725 VGND 0.02407f
C11904 VPWR.n543 VGND 0.07442f
C11905 VPWR.n544 VGND 0.0512f
C11906 VPWR.n545 VGND 0.2969f
C11907 VPWR.n546 VGND 0.06791f
C11908 VPWR.n547 VGND 0.2969f
C11909 VPWR.n548 VGND 0.2969f
C11910 VPWR.n550 VGND 0.2969f
C11911 VPWR.n552 VGND 0.2969f
C11912 VPWR.n553 VGND 0.0512f
C11913 VPWR.t308 VGND 0.02709f
C11914 VPWR.t176 VGND 0.02407f
C11915 VPWR.n554 VGND 0.07442f
C11916 VPWR.t893 VGND 0.07496f
C11917 VPWR.t720 VGND 0.02709f
C11918 VPWR.t894 VGND 0.02407f
C11919 VPWR.n555 VGND 0.07442f
C11920 VPWR.n556 VGND 0.0512f
C11921 VPWR.n557 VGND 0.2969f
C11922 VPWR.n558 VGND 0.2969f
C11923 VPWR.n560 VGND 0.2969f
C11924 VPWR.n562 VGND 0.2969f
C11925 VPWR.n563 VGND 0.0512f
C11926 VPWR.t1069 VGND 0.02709f
C11927 VPWR.t1665 VGND 0.02407f
C11928 VPWR.n565 VGND 0.07442f
C11929 VPWR.t1664 VGND 0.07496f
C11930 VPWR.t432 VGND 0.09722f
C11931 VPWR.t1780 VGND 0.02709f
C11932 VPWR.t439 VGND 0.02407f
C11933 VPWR.n566 VGND 0.07442f
C11934 VPWR.t433 VGND 0.02709f
C11935 VPWR.t85 VGND 0.02407f
C11936 VPWR.n567 VGND 0.07442f
C11937 VPWR.t298 VGND 0.06383f
C11938 VPWR.t84 VGND 0.07496f
C11939 VPWR.t315 VGND 0.06383f
C11940 VPWR.t719 VGND 0.09722f
C11941 VPWR.t79 VGND 0.02709f
C11942 VPWR.t61 VGND 0.02407f
C11943 VPWR.n568 VGND 0.07442f
C11944 VPWR.n570 VGND 0.088f
C11945 VPWR.t60 VGND 0.07496f
C11946 VPWR.t316 VGND 0.06383f
C11947 VPWR.t78 VGND 0.09722f
C11948 VPWR.n571 VGND 0.088f
C11949 VPWR.n573 VGND 0.0512f
C11950 VPWR.n574 VGND 0.2969f
C11951 VPWR.n575 VGND 0.2969f
C11952 VPWR.n577 VGND 0.2969f
C11953 VPWR.n578 VGND 0.0512f
C11954 VPWR.t909 VGND 0.02709f
C11955 VPWR.t215 VGND 0.02407f
C11956 VPWR.n580 VGND 0.07442f
C11957 VPWR.t214 VGND 0.07496f
C11958 VPWR.t1905 VGND 0.09722f
C11959 VPWR.t1053 VGND 0.02709f
C11960 VPWR.t1912 VGND 0.02407f
C11961 VPWR.n581 VGND 0.07442f
C11962 VPWR.n582 VGND 0.2969f
C11963 VPWR.n583 VGND 0.2969f
C11964 VPWR.n585 VGND 0.2969f
C11965 VPWR.n586 VGND 0.0512f
C11966 VPWR.t11 VGND 0.02709f
C11967 VPWR.t529 VGND 0.02407f
C11968 VPWR.n588 VGND 0.07442f
C11969 VPWR.t528 VGND 0.07496f
C11970 VPWR.t581 VGND 0.02709f
C11971 VPWR.t1234 VGND 0.02407f
C11972 VPWR.n589 VGND 0.07442f
C11973 VPWR.n590 VGND 0.2969f
C11974 VPWR.n591 VGND 0.06791f
C11975 VPWR.n592 VGND 0.82597f
C11976 VPWR.n593 VGND 0.2969f
C11977 VPWR.n594 VGND 0.0512f
C11978 VPWR.t585 VGND 0.02709f
C11979 VPWR.t1194 VGND 0.02407f
C11980 VPWR.n596 VGND 0.07442f
C11981 VPWR.t26 VGND 0.07496f
C11982 VPWR.t192 VGND 0.02709f
C11983 VPWR.t27 VGND 0.02407f
C11984 VPWR.n597 VGND 0.07442f
C11985 VPWR.t1813 VGND 0.02709f
C11986 VPWR.t205 VGND 0.02407f
C11987 VPWR.n598 VGND 0.07442f
C11988 VPWR.t906 VGND 0.07496f
C11989 VPWR.t766 VGND 0.02709f
C11990 VPWR.t907 VGND 0.02407f
C11991 VPWR.n599 VGND 0.07442f
C11992 VPWR.n600 VGND 0.2969f
C11993 VPWR.n601 VGND 0.2969f
C11994 VPWR.n604 VGND 0.2969f
C11995 VPWR.n605 VGND 0.0512f
C11996 VPWR.t361 VGND 0.02709f
C11997 VPWR.t1580 VGND 0.02407f
C11998 VPWR.n606 VGND 0.07442f
C11999 VPWR.t122 VGND 0.07496f
C12000 VPWR.t517 VGND 0.02709f
C12001 VPWR.t123 VGND 0.02407f
C12002 VPWR.n607 VGND 0.07442f
C12003 VPWR.n608 VGND 0.2969f
C12004 VPWR.n609 VGND 0.2969f
C12005 VPWR.t480 VGND 0.02709f
C12006 VPWR.t3 VGND 0.02407f
C12007 VPWR.n610 VGND 0.07442f
C12008 VPWR.t457 VGND 0.07496f
C12009 VPWR.t168 VGND 0.02709f
C12010 VPWR.t458 VGND 0.02407f
C12011 VPWR.n611 VGND 0.07442f
C12012 VPWR.n612 VGND 0.2969f
C12013 VPWR.n613 VGND 0.2969f
C12014 VPWR.t160 VGND 0.02709f
C12015 VPWR.t172 VGND 0.02407f
C12016 VPWR.n614 VGND 0.07442f
C12017 VPWR.t1695 VGND 0.07496f
C12018 VPWR.t731 VGND 0.02709f
C12019 VPWR.t1696 VGND 0.02407f
C12020 VPWR.n615 VGND 0.07442f
C12021 VPWR.n616 VGND 0.0512f
C12022 VPWR.n617 VGND 0.2969f
C12023 VPWR.n618 VGND 0.2969f
C12024 VPWR.t1628 VGND 0.02709f
C12025 VPWR.t1519 VGND 0.02407f
C12026 VPWR.n619 VGND 0.07442f
C12027 VPWR.t770 VGND 0.07496f
C12028 VPWR.t795 VGND 0.02709f
C12029 VPWR.t771 VGND 0.02407f
C12030 VPWR.n620 VGND 0.07442f
C12031 VPWR.n621 VGND 0.2969f
C12032 VPWR.n622 VGND 0.2969f
C12033 VPWR.n623 VGND 0.2969f
C12034 VPWR.t622 VGND 0.02709f
C12035 VPWR.t1686 VGND 0.02407f
C12036 VPWR.n624 VGND 0.07442f
C12037 VPWR.t621 VGND 0.118f
C12038 VPWR.t881 VGND 0.06383f
C12039 VPWR.t1685 VGND 0.07496f
C12040 VPWR.t1646 VGND 0.06383f
C12041 VPWR.t794 VGND 0.09722f
C12042 VPWR.n625 VGND 0.088f
C12043 VPWR.n627 VGND -0.05607f
C12044 VPWR.t616 VGND 0.02709f
C12045 VPWR.t801 VGND 0.02407f
C12046 VPWR.n628 VGND 0.07442f
C12047 VPWR.t249 VGND 0.02709f
C12048 VPWR.t1926 VGND 0.02407f
C12049 VPWR.n631 VGND 0.07442f
C12050 VPWR.t615 VGND 0.118f
C12051 VPWR.t850 VGND 0.06383f
C12052 VPWR.t800 VGND 0.07496f
C12053 VPWR.n632 VGND 0.088f
C12054 VPWR.t248 VGND 0.09722f
C12055 VPWR.t105 VGND 0.06383f
C12056 VPWR.t1925 VGND 0.07496f
C12057 VPWR.t1526 VGND 0.09722f
C12058 VPWR.t962 VGND 0.02709f
C12059 VPWR.t1503 VGND 0.02407f
C12060 VPWR.n633 VGND 0.07442f
C12061 VPWR.t1527 VGND 0.02709f
C12062 VPWR.t1071 VGND 0.02407f
C12063 VPWR.n635 VGND 0.07442f
C12064 VPWR.t495 VGND 0.06383f
C12065 VPWR.t1070 VGND 0.07496f
C12066 VPWR.t407 VGND 0.09722f
C12067 VPWR.t1743 VGND 0.02709f
C12068 VPWR.t414 VGND 0.02407f
C12069 VPWR.n636 VGND 0.07442f
C12070 VPWR.t408 VGND 0.02709f
C12071 VPWR.t472 VGND 0.02407f
C12072 VPWR.n638 VGND 0.07442f
C12073 VPWR.t293 VGND 0.06383f
C12074 VPWR.t471 VGND 0.07496f
C12075 VPWR.t110 VGND 0.09722f
C12076 VPWR.t466 VGND 0.02709f
C12077 VPWR.t724 VGND 0.02407f
C12078 VPWR.n639 VGND 0.07442f
C12079 VPWR.t111 VGND 0.02709f
C12080 VPWR.t571 VGND 0.02407f
C12081 VPWR.n641 VGND 0.07442f
C12082 VPWR.t563 VGND 0.06383f
C12083 VPWR.t570 VGND 0.07496f
C12084 VPWR.t265 VGND 0.09722f
C12085 VPWR.t422 VGND 0.02709f
C12086 VPWR.t272 VGND 0.02407f
C12087 VPWR.n642 VGND 0.07442f
C12088 VPWR.t266 VGND 0.02709f
C12089 VPWR.t760 VGND 0.02407f
C12090 VPWR.n644 VGND 0.07442f
C12091 VPWR.t852 VGND 0.06383f
C12092 VPWR.t759 VGND 0.07496f
C12093 VPWR.t292 VGND 0.06383f
C12094 VPWR.t908 VGND 0.09722f
C12095 VPWR.t1023 VGND 0.02709f
C12096 VPWR.t1545 VGND 0.02407f
C12097 VPWR.n645 VGND 0.07442f
C12098 VPWR.n647 VGND 0.088f
C12099 VPWR.t1544 VGND 0.07496f
C12100 VPWR.t851 VGND 0.06383f
C12101 VPWR.t1022 VGND 0.09722f
C12102 VPWR.n648 VGND 0.088f
C12103 VPWR.n650 VGND 0.0512f
C12104 VPWR.n652 VGND 0.0512f
C12105 VPWR.n654 VGND 0.088f
C12106 VPWR.t271 VGND 0.07496f
C12107 VPWR.t1581 VGND 0.06383f
C12108 VPWR.t421 VGND 0.09722f
C12109 VPWR.n655 VGND 0.088f
C12110 VPWR.n657 VGND 0.0512f
C12111 VPWR.n659 VGND 0.0512f
C12112 VPWR.n661 VGND 0.088f
C12113 VPWR.t723 VGND 0.07496f
C12114 VPWR.t564 VGND 0.06383f
C12115 VPWR.t465 VGND 0.09722f
C12116 VPWR.n662 VGND 0.088f
C12117 VPWR.n664 VGND 0.0512f
C12118 VPWR.n666 VGND 0.0512f
C12119 VPWR.n668 VGND 0.088f
C12120 VPWR.t413 VGND 0.07496f
C12121 VPWR.t294 VGND 0.06383f
C12122 VPWR.t1742 VGND 0.09722f
C12123 VPWR.t1794 VGND 0.02709f
C12124 VPWR.t1678 VGND 0.02407f
C12125 VPWR.n669 VGND 0.07442f
C12126 VPWR.n670 VGND 0.0512f
C12127 VPWR.n672 VGND 0.088f
C12128 VPWR.t1677 VGND 0.07496f
C12129 VPWR.t565 VGND 0.06383f
C12130 VPWR.t1793 VGND 0.09722f
C12131 VPWR.n673 VGND 0.088f
C12132 VPWR.n675 VGND 0.0512f
C12133 VPWR.n677 VGND 0.0512f
C12134 VPWR.n679 VGND 0.088f
C12135 VPWR.t1502 VGND 0.07496f
C12136 VPWR.t496 VGND 0.06383f
C12137 VPWR.t961 VGND 0.09722f
C12138 VPWR.n680 VGND 0.088f
C12139 VPWR.n682 VGND 0.0512f
C12140 VPWR.n683 VGND -0.05607f
C12141 VPWR.t604 VGND 0.02709f
C12142 VPWR.t492 VGND 0.02407f
C12143 VPWR.n684 VGND 0.07442f
C12144 VPWR.t253 VGND 0.02709f
C12145 VPWR.t450 VGND 0.02407f
C12146 VPWR.n687 VGND 0.07442f
C12147 VPWR.t603 VGND 0.118f
C12148 VPWR.t318 VGND 0.06383f
C12149 VPWR.t491 VGND 0.07496f
C12150 VPWR.n688 VGND 0.088f
C12151 VPWR.t252 VGND 0.09722f
C12152 VPWR.t313 VGND 0.06383f
C12153 VPWR.t449 VGND 0.07496f
C12154 VPWR.t317 VGND 0.06383f
C12155 VPWR.t1068 VGND 0.09722f
C12156 VPWR.t1507 VGND 0.02709f
C12157 VPWR.t823 VGND 0.02407f
C12158 VPWR.n689 VGND 0.07442f
C12159 VPWR.n691 VGND 0.088f
C12160 VPWR.t822 VGND 0.07496f
C12161 VPWR.t398 VGND 0.06383f
C12162 VPWR.t1506 VGND 0.09722f
C12163 VPWR.t509 VGND 0.02709f
C12164 VPWR.t1483 VGND 0.02407f
C12165 VPWR.n692 VGND 0.07442f
C12166 VPWR.n693 VGND 0.0512f
C12167 VPWR.n695 VGND 0.088f
C12168 VPWR.t1482 VGND 0.07496f
C12169 VPWR.t399 VGND 0.06383f
C12170 VPWR.t508 VGND 0.09722f
C12171 VPWR.n696 VGND 0.088f
C12172 VPWR.n698 VGND 0.0512f
C12173 VPWR.n699 VGND -0.05607f
C12174 VPWR.n700 VGND 0.06791f
C12175 VPWR.n701 VGND 0.06791f
C12176 VPWR.n702 VGND 0.2969f
C12177 VPWR.n703 VGND 0.82079f
C12178 VPWR.n704 VGND 0.06791f
C12179 VPWR.n705 VGND 0.06791f
C12180 VPWR.n706 VGND 0.06791f
C12181 VPWR.n707 VGND 0.06791f
C12182 VPWR.n708 VGND 0.06791f
C12183 VPWR.n709 VGND 0.2969f
C12184 VPWR.n711 VGND 0.2969f
C12185 VPWR.n712 VGND 0.0512f
C12186 VPWR.t1850 VGND 0.02709f
C12187 VPWR.t1846 VGND 0.02407f
C12188 VPWR.n714 VGND 0.07442f
C12189 VPWR.t1845 VGND 0.07496f
C12190 VPWR.t808 VGND 0.09722f
C12191 VPWR.t1840 VGND 0.02709f
C12192 VPWR.t655 VGND 0.02407f
C12193 VPWR.n715 VGND 0.07442f
C12194 VPWR.n716 VGND 0.2969f
C12195 VPWR.n717 VGND 0.2969f
C12196 VPWR.n718 VGND 0.0512f
C12197 VPWR.t669 VGND 0.02709f
C12198 VPWR.t357 VGND 0.02407f
C12199 VPWR.n720 VGND 0.07442f
C12200 VPWR.t1619 VGND 0.06383f
C12201 VPWR.t674 VGND 0.07496f
C12202 VPWR.t809 VGND 0.02709f
C12203 VPWR.t675 VGND 0.02407f
C12204 VPWR.n721 VGND 0.07442f
C12205 VPWR.n723 VGND 0.088f
C12206 VPWR.t668 VGND 0.09722f
C12207 VPWR.t1616 VGND 0.06383f
C12208 VPWR.t356 VGND 0.07496f
C12209 VPWR.t745 VGND 0.09722f
C12210 VPWR.t1894 VGND 0.02709f
C12211 VPWR.t752 VGND 0.02407f
C12212 VPWR.n724 VGND 0.07442f
C12213 VPWR.t746 VGND 0.02709f
C12214 VPWR.t1595 VGND 0.02407f
C12215 VPWR.n726 VGND 0.07442f
C12216 VPWR.t440 VGND 0.06383f
C12217 VPWR.t1594 VGND 0.07496f
C12218 VPWR.t1468 VGND 0.09722f
C12219 VPWR.t1605 VGND 0.02709f
C12220 VPWR.t1047 VGND 0.02407f
C12221 VPWR.n727 VGND 0.07442f
C12222 VPWR.n728 VGND 0.2969f
C12223 VPWR.n729 VGND 0.2969f
C12224 VPWR.n730 VGND 0.0512f
C12225 VPWR.t1706 VGND 0.02709f
C12226 VPWR.t589 VGND 0.02407f
C12227 VPWR.n732 VGND 0.07442f
C12228 VPWR.t445 VGND 0.06383f
C12229 VPWR.t6 VGND 0.07496f
C12230 VPWR.t1469 VGND 0.02709f
C12231 VPWR.t7 VGND 0.02407f
C12232 VPWR.n733 VGND 0.07442f
C12233 VPWR.n735 VGND 0.088f
C12234 VPWR.t1705 VGND 0.09722f
C12235 VPWR.t444 VGND 0.06383f
C12236 VPWR.t588 VGND 0.07496f
C12237 VPWR.t1719 VGND 0.02709f
C12238 VPWR.t1299 VGND 0.02407f
C12239 VPWR.n736 VGND 0.07442f
C12240 VPWR.n737 VGND 0.2969f
C12241 VPWR.n739 VGND 0.82597f
C12242 VPWR.n740 VGND 0.2969f
C12243 VPWR.n743 VGND 0.2969f
C12244 VPWR.n744 VGND 0.0512f
C12245 VPWR.t911 VGND 0.02709f
C12246 VPWR.t217 VGND 0.02407f
C12247 VPWR.n746 VGND 0.07442f
C12248 VPWR.t761 VGND 0.07496f
C12249 VPWR.t268 VGND 0.02709f
C12250 VPWR.t762 VGND 0.02407f
C12251 VPWR.n747 VGND 0.07442f
C12252 VPWR.n748 VGND 0.2969f
C12253 VPWR.n749 VGND 0.2969f
C12254 VPWR.t567 VGND 0.02709f
C12255 VPWR.t274 VGND 0.02407f
C12256 VPWR.n750 VGND 0.07442f
C12257 VPWR.t572 VGND 0.07496f
C12258 VPWR.t113 VGND 0.02709f
C12259 VPWR.t573 VGND 0.02407f
C12260 VPWR.n751 VGND 0.07442f
C12261 VPWR.t468 VGND 0.02709f
C12262 VPWR.t726 VGND 0.02407f
C12263 VPWR.n752 VGND 0.07442f
C12264 VPWR.t473 VGND 0.07496f
C12265 VPWR.t410 VGND 0.02709f
C12266 VPWR.t474 VGND 0.02407f
C12267 VPWR.n753 VGND 0.07442f
C12268 VPWR.n754 VGND 0.2969f
C12269 VPWR.n755 VGND 0.06791f
C12270 VPWR.n756 VGND 0.2969f
C12271 VPWR.n757 VGND 0.2969f
C12272 VPWR.n760 VGND 0.2969f
C12273 VPWR.n761 VGND 0.0512f
C12274 VPWR.t1495 VGND 0.02709f
C12275 VPWR.t1788 VGND 0.02407f
C12276 VPWR.n762 VGND 0.07442f
C12277 VPWR.t943 VGND 0.07496f
C12278 VPWR.t701 VGND 0.02709f
C12279 VPWR.t944 VGND 0.02407f
C12280 VPWR.n763 VGND 0.07442f
C12281 VPWR.n764 VGND 0.2969f
C12282 VPWR.n765 VGND 0.2969f
C12283 VPWR.t614 VGND 0.02709f
C12284 VPWR.t803 VGND 0.02407f
C12285 VPWR.n766 VGND 0.07442f
C12286 VPWR.t1565 VGND 0.02709f
C12287 VPWR.t1928 VGND 0.02407f
C12288 VPWR.n769 VGND 0.07442f
C12289 VPWR.t613 VGND 0.118f
C12290 VPWR.t876 VGND 0.06383f
C12291 VPWR.t802 VGND 0.07496f
C12292 VPWR.n770 VGND 0.088f
C12293 VPWR.t1564 VGND 0.09722f
C12294 VPWR.t1809 VGND 0.06383f
C12295 VPWR.t1927 VGND 0.07496f
C12296 VPWR.t1524 VGND 0.09722f
C12297 VPWR.t964 VGND 0.02709f
C12298 VPWR.t1501 VGND 0.02407f
C12299 VPWR.n771 VGND 0.07442f
C12300 VPWR.t1525 VGND 0.02709f
C12301 VPWR.t1075 VGND 0.02407f
C12302 VPWR.n772 VGND 0.07442f
C12303 VPWR.t684 VGND 0.06383f
C12304 VPWR.t1074 VGND 0.07496f
C12305 VPWR.t1744 VGND 0.09722f
C12306 VPWR.t708 VGND 0.02709f
C12307 VPWR.t1680 VGND 0.02407f
C12308 VPWR.n773 VGND 0.07442f
C12309 VPWR.t1745 VGND 0.02709f
C12310 VPWR.t1878 VGND 0.02407f
C12311 VPWR.n775 VGND 0.07442f
C12312 VPWR.t690 VGND 0.06383f
C12313 VPWR.t1877 VGND 0.07496f
C12314 VPWR.t689 VGND 0.06383f
C12315 VPWR.t409 VGND 0.09722f
C12316 VPWR.n776 VGND 0.088f
C12317 VPWR.n778 VGND 0.0512f
C12318 VPWR.n780 VGND 0.0512f
C12319 VPWR.n782 VGND 0.088f
C12320 VPWR.t1679 VGND 0.07496f
C12321 VPWR.t875 VGND 0.06383f
C12322 VPWR.t707 VGND 0.09722f
C12323 VPWR.n783 VGND 0.088f
C12324 VPWR.n785 VGND 0.0512f
C12325 VPWR.n787 VGND 0.0512f
C12326 VPWR.n789 VGND 0.088f
C12327 VPWR.t1500 VGND 0.07496f
C12328 VPWR.t685 VGND 0.06383f
C12329 VPWR.t963 VGND 0.09722f
C12330 VPWR.n790 VGND 0.088f
C12331 VPWR.n792 VGND 0.0512f
C12332 VPWR.n793 VGND -0.05607f
C12333 VPWR.n794 VGND 0.82079f
C12334 VPWR.n795 VGND 0.2969f
C12335 VPWR.n796 VGND 0.0512f
C12336 VPWR.t1624 VGND 0.02709f
C12337 VPWR.t1533 VGND 0.02407f
C12338 VPWR.n798 VGND 0.07442f
C12339 VPWR.t599 VGND 0.118f
C12340 VPWR.t1808 VGND 0.06383f
C12341 VPWR.t788 VGND 0.07496f
C12342 VPWR.t600 VGND 0.02709f
C12343 VPWR.t789 VGND 0.02407f
C12344 VPWR.n799 VGND 0.07442f
C12345 VPWR.n800 VGND -0.05607f
C12346 VPWR.n802 VGND 0.088f
C12347 VPWR.t698 VGND 0.09722f
C12348 VPWR.t1915 VGND 0.06383f
C12349 VPWR.t941 VGND 0.07496f
C12350 VPWR.t699 VGND 0.02709f
C12351 VPWR.t942 VGND 0.02407f
C12352 VPWR.n803 VGND 0.07442f
C12353 VPWR.n805 VGND 0.088f
C12354 VPWR.t1623 VGND 0.09722f
C12355 VPWR.t197 VGND 0.06383f
C12356 VPWR.t1532 VGND 0.07496f
C12357 VPWR.t814 VGND 0.09722f
C12358 VPWR.t1497 VGND 0.02709f
C12359 VPWR.t1786 VGND 0.02407f
C12360 VPWR.n806 VGND 0.07442f
C12361 VPWR.t815 VGND 0.02709f
C12362 VPWR.t1587 VGND 0.02407f
C12363 VPWR.n808 VGND 0.07442f
C12364 VPWR.t1807 VGND 0.06383f
C12365 VPWR.t1586 VGND 0.07496f
C12366 VPWR.t1847 VGND 0.09722f
C12367 VPWR.t925 VGND 0.02709f
C12368 VPWR.t1854 VGND 0.02407f
C12369 VPWR.n809 VGND 0.07442f
C12370 VPWR.n810 VGND 0.2969f
C12371 VPWR.n811 VGND 0.2969f
C12372 VPWR.n812 VGND 0.0512f
C12373 VPWR.t805 VGND 0.02709f
C12374 VPWR.t673 VGND 0.02407f
C12375 VPWR.n814 VGND 0.07442f
C12376 VPWR.t201 VGND 0.06383f
C12377 VPWR.t1843 VGND 0.07496f
C12378 VPWR.t1848 VGND 0.02709f
C12379 VPWR.t1844 VGND 0.02407f
C12380 VPWR.n815 VGND 0.07442f
C12381 VPWR.n817 VGND 0.0512f
C12382 VPWR.n819 VGND 0.088f
C12383 VPWR.t1837 VGND 0.09722f
C12384 VPWR.t1806 VGND 0.06383f
C12385 VPWR.t652 VGND 0.07496f
C12386 VPWR.t1838 VGND 0.02709f
C12387 VPWR.t653 VGND 0.02407f
C12388 VPWR.n820 VGND 0.07442f
C12389 VPWR.n822 VGND 0.088f
C12390 VPWR.t804 VGND 0.09722f
C12391 VPWR.t1917 VGND 0.06383f
C12392 VPWR.t672 VGND 0.07496f
C12393 VPWR.t1891 VGND 0.09722f
C12394 VPWR.t667 VGND 0.02709f
C12395 VPWR.t355 VGND 0.02407f
C12396 VPWR.n823 VGND 0.07442f
C12397 VPWR.t1892 VGND 0.02709f
C12398 VPWR.t750 VGND 0.02407f
C12399 VPWR.n825 VGND 0.07442f
C12400 VPWR.t195 VGND 0.06383f
C12401 VPWR.t749 VGND 0.07496f
C12402 VPWR.t1614 VGND 0.09722f
C12403 VPWR.t221 VGND 0.02709f
C12404 VPWR.t1611 VGND 0.02407f
C12405 VPWR.n826 VGND 0.07442f
C12406 VPWR.t1615 VGND 0.02709f
C12407 VPWR.t194 VGND 0.02407f
C12408 VPWR.n828 VGND 0.07442f
C12409 VPWR.t200 VGND 0.06383f
C12410 VPWR.t193 VGND 0.07496f
C12411 VPWR.t1703 VGND 0.09722f
C12412 VPWR.t1465 VGND 0.02709f
C12413 VPWR.t23 VGND 0.02407f
C12414 VPWR.n829 VGND 0.07442f
C12415 VPWR.t1704 VGND 0.02709f
C12416 VPWR.t587 VGND 0.02407f
C12417 VPWR.n830 VGND 0.07442f
C12418 VPWR.t198 VGND 0.06383f
C12419 VPWR.t586 VGND 0.07496f
C12420 VPWR.t1717 VGND 0.02709f
C12421 VPWR.t1306 VGND 0.02407f
C12422 VPWR.n831 VGND 0.07442f
C12423 VPWR.n833 VGND 0.0512f
C12424 VPWR.n834 VGND 0.06192f
C12425 VPWR.t1305 VGND 0.10842f
C12426 VPWR.t1916 VGND 0.06383f
C12427 VPWR.t1716 VGND 0.09722f
C12428 VPWR.n835 VGND 0.088f
C12429 VPWR.n837 VGND 0.0512f
C12430 VPWR.n838 VGND 0.2969f
C12431 VPWR.n839 VGND 0.29751f
C12432 VPWR.n841 VGND 0.29751f
C12433 VPWR.t997 VGND 0.02709f
C12434 VPWR.t1420 VGND 0.02407f
C12435 VPWR.n842 VGND 0.07442f
C12436 VPWR.t1720 VGND 0.07496f
C12437 VPWR.t1632 VGND 0.02709f
C12438 VPWR.t1721 VGND 0.02407f
C12439 VPWR.n843 VGND 0.07442f
C12440 VPWR.t209 VGND 0.02709f
C12441 VPWR.t115 VGND 0.02407f
C12442 VPWR.n844 VGND 0.07442f
C12443 VPWR.t1474 VGND 0.07496f
C12444 VPWR.t1821 VGND 0.02709f
C12445 VPWR.t1475 VGND 0.02407f
C12446 VPWR.n845 VGND 0.07442f
C12447 VPWR.n846 VGND 0.0512f
C12448 VPWR.n847 VGND 0.29751f
C12449 VPWR.n848 VGND 0.29751f
C12450 VPWR.t306 VGND 0.02709f
C12451 VPWR.t174 VGND 0.02407f
C12452 VPWR.n849 VGND 0.07442f
C12453 VPWR.t1556 VGND 0.07496f
C12454 VPWR.t1043 VGND 0.02709f
C12455 VPWR.t1557 VGND 0.02407f
C12456 VPWR.n850 VGND 0.07442f
C12457 VPWR.n851 VGND 0.29751f
C12458 VPWR.n852 VGND 0.29751f
C12459 VPWR.n853 VGND 0.06791f
C12460 VPWR.n854 VGND 0.06791f
C12461 VPWR.n855 VGND 0.06791f
C12462 VPWR.n856 VGND 0.06791f
C12463 VPWR.n857 VGND 0.2969f
C12464 VPWR.t718 VGND 0.02709f
C12465 VPWR.t892 VGND 0.02407f
C12466 VPWR.n858 VGND 0.07442f
C12467 VPWR.t56 VGND 0.07496f
C12468 VPWR.t75 VGND 0.02709f
C12469 VPWR.t57 VGND 0.02407f
C12470 VPWR.n859 VGND 0.07442f
C12471 VPWR.n860 VGND 0.0512f
C12472 VPWR.n861 VGND 0.29751f
C12473 VPWR.n862 VGND 0.29751f
C12474 VPWR.n864 VGND 0.29751f
C12475 VPWR.n866 VGND 0.29751f
C12476 VPWR.n867 VGND 0.0512f
C12477 VPWR.t1067 VGND 0.02709f
C12478 VPWR.t1784 VGND 0.02407f
C12479 VPWR.n868 VGND 0.07442f
C12480 VPWR.t1484 VGND 0.07496f
C12481 VPWR.t505 VGND 0.02709f
C12482 VPWR.t1485 VGND 0.02407f
C12483 VPWR.n869 VGND 0.07442f
C12484 VPWR.t251 VGND 0.02709f
C12485 VPWR.t513 VGND 0.02407f
C12486 VPWR.n870 VGND 0.07442f
C12487 VPWR.t605 VGND 0.118f
C12488 VPWR.t101 VGND 0.06383f
C12489 VPWR.t489 VGND 0.07496f
C12490 VPWR.t606 VGND 0.02709f
C12491 VPWR.t490 VGND 0.02407f
C12492 VPWR.n871 VGND 0.07442f
C12493 VPWR.n872 VGND 0.10954f
C12494 VPWR.n873 VGND -0.05607f
C12495 VPWR.n874 VGND 0.10954f
C12496 VPWR.n875 VGND 0.0512f
C12497 VPWR.t946 VGND 0.02709f
C12498 VPWR.t1521 VGND 0.02407f
C12499 VPWR.n877 VGND 0.07442f
C12500 VPWR.t590 VGND 0.118f
C12501 VPWR.t1859 VGND 0.06383f
C12502 VPWR.t1683 VGND 0.07496f
C12503 VPWR.t591 VGND 0.02709f
C12504 VPWR.t1684 VGND 0.02407f
C12505 VPWR.n878 VGND 0.07442f
C12506 VPWR.n880 VGND 0.088f
C12507 VPWR.t704 VGND 0.09722f
C12508 VPWR.t90 VGND 0.06383f
C12509 VPWR.t1625 VGND 0.07496f
C12510 VPWR.t705 VGND 0.02709f
C12511 VPWR.t1626 VGND 0.02407f
C12512 VPWR.n881 VGND 0.07442f
C12513 VPWR.n883 VGND 0.088f
C12514 VPWR.t945 VGND 0.09722f
C12515 VPWR.t1863 VGND 0.06383f
C12516 VPWR.t1520 VGND 0.07496f
C12517 VPWR.t826 VGND 0.09722f
C12518 VPWR.t1487 VGND 0.02709f
C12519 VPWR.t1792 VGND 0.02407f
C12520 VPWR.n884 VGND 0.07442f
C12521 VPWR.t827 VGND 0.02709f
C12522 VPWR.t158 VGND 0.02407f
C12523 VPWR.n886 VGND 0.07442f
C12524 VPWR.t744 VGND 0.06383f
C12525 VPWR.t157 VGND 0.07496f
C12526 VPWR.t1857 VGND 0.09722f
C12527 VPWR.t1591 VGND 0.02709f
C12528 VPWR.t166 VGND 0.02407f
C12529 VPWR.n887 VGND 0.07442f
C12530 VPWR.n888 VGND 0.10954f
C12531 VPWR.n889 VGND 0.06791f
C12532 VPWR.n890 VGND 0.06791f
C12533 VPWR.n891 VGND 0.06791f
C12534 VPWR.n892 VGND 0.10954f
C12535 VPWR.n893 VGND 0.0512f
C12536 VPWR.t59 VGND 0.02709f
C12537 VPWR.t661 VGND 0.02407f
C12538 VPWR.n895 VGND 0.07442f
C12539 VPWR.t87 VGND 0.06383f
C12540 VPWR.t1771 VGND 0.07496f
C12541 VPWR.t1858 VGND 0.02709f
C12542 VPWR.t1772 VGND 0.02407f
C12543 VPWR.n896 VGND 0.07442f
C12544 VPWR.n898 VGND 0.0512f
C12545 VPWR.n900 VGND 0.088f
C12546 VPWR.t1767 VGND 0.09722f
C12547 VPWR.t279 VGND 0.06383f
C12548 VPWR.t108 VGND 0.07496f
C12549 VPWR.t1768 VGND 0.02709f
C12550 VPWR.t109 VGND 0.02407f
C12551 VPWR.n901 VGND 0.07442f
C12552 VPWR.n903 VGND 0.088f
C12553 VPWR.t58 VGND 0.09722f
C12554 VPWR.t278 VGND 0.06383f
C12555 VPWR.t660 VGND 0.07496f
C12556 VPWR.t1897 VGND 0.09722f
C12557 VPWR.t657 VGND 0.02709f
C12558 VPWR.t365 VGND 0.02407f
C12559 VPWR.n904 VGND 0.07442f
C12560 VPWR.t1898 VGND 0.02709f
C12561 VPWR.t758 VGND 0.02407f
C12562 VPWR.n906 VGND 0.07442f
C12563 VPWR.t1861 VGND 0.06383f
C12564 VPWR.t757 VGND 0.07496f
C12565 VPWR.t1608 VGND 0.09722f
C12566 VPWR.t754 VGND 0.02709f
C12567 VPWR.t1603 VGND 0.02407f
C12568 VPWR.n907 VGND 0.07442f
C12569 VPWR.t1609 VGND 0.02709f
C12570 VPWR.t1051 VGND 0.02407f
C12571 VPWR.n909 VGND 0.07442f
C12572 VPWR.t86 VGND 0.06383f
C12573 VPWR.t1050 VGND 0.07496f
C12574 VPWR.t20 VGND 0.09722f
C12575 VPWR.t1477 VGND 0.02709f
C12576 VPWR.t15 VGND 0.02407f
C12577 VPWR.n910 VGND 0.07442f
C12578 VPWR.n911 VGND 0.10954f
C12579 VPWR.n912 VGND 0.06791f
C12580 VPWR.n913 VGND 0.06791f
C12581 VPWR.n914 VGND 0.06791f
C12582 VPWR.n915 VGND 0.06791f
C12583 VPWR.n916 VGND 0.06791f
C12584 VPWR.n917 VGND -0.01517f
C12585 VPWR.n918 VGND 0.04424f
C12586 VPWR.n919 VGND 0.0512f
C12587 VPWR.n921 VGND 0.02474f
C12588 VPWR.t1269 VGND 0.02178f
C12589 VPWR.n923 VGND 0.04654f
C12590 VPWR.t1389 VGND 0.02407f
C12591 VPWR.n924 VGND 0.03816f
C12592 VPWR.t1550 VGND 0.07496f
C12593 VPWR.n925 VGND 0.02474f
C12594 VPWR.t1124 VGND 0.02178f
C12595 VPWR.n927 VGND 0.04654f
C12596 VPWR.t1551 VGND 0.02407f
C12597 VPWR.n928 VGND 0.03816f
C12598 VPWR.n929 VGND 0.0512f
C12599 VPWR.n930 VGND -0.01517f
C12600 VPWR.n931 VGND 0.0534f
C12601 VPWR.n932 VGND 0.0746f
C12602 VPWR.t1392 VGND 0.01009f
C12603 VPWR.n933 VGND 0.02252f
C12604 VPWR.n934 VGND 0.01543f
C12605 VPWR.n935 VGND 0.05077f
C12606 VPWR.n936 VGND 0.07925f
C12607 VPWR.n937 VGND 0.15751f
C12608 VPWR.n938 VGND 0.82597f
C12609 VPWR.n939 VGND 0.82597f
C12610 VPWR.n941 VGND 0.03811f
C12611 VPWR.t150 VGND 0.79335f
C12612 VPWR.n942 VGND 0.4327f
C12613 VPWR.t64 VGND 0.79335f
C12614 VPWR.n943 VGND 0.33651f
C12615 VPWR.n944 VGND 0.23646f
C12616 VPWR.t560 VGND 0.04648f
C12617 VPWR.t664 VGND 0.01165f
C12618 VPWR.t781 VGND 0.01165f
C12619 VPWR.n946 VGND 0.02558f
C12620 VPWR.t782 VGND 0.01165f
C12621 VPWR.t151 VGND 0.01165f
C12622 VPWR.n947 VGND 0.02554f
C12623 VPWR.t384 VGND 0.01165f
C12624 VPWR.t383 VGND 0.01165f
C12625 VPWR.n948 VGND 0.02554f
C12626 VPWR.n949 VGND 0.08473f
C12627 VPWR.n950 VGND 0.14784f
C12628 VPWR.n951 VGND 0.04681f
C12629 VPWR.n952 VGND 0.03438f
C12630 VPWR.t380 VGND 0.01165f
C12631 VPWR.t385 VGND 0.01165f
C12632 VPWR.n953 VGND 0.02558f
C12633 VPWR.n954 VGND 0.10491f
C12634 VPWR.n956 VGND 0.01326f
C12635 VPWR.n957 VGND 0.01553f
C12636 VPWR.n958 VGND 0.02278f
C12637 VPWR.t558 VGND 0.04648f
C12638 VPWR.n959 VGND 0.12245f
C12639 VPWR.t1571 VGND 0.04646f
C12640 VPWR.t65 VGND 0.04646f
C12641 VPWR.n961 VGND 0.10933f
C12642 VPWR.n962 VGND 0.27291f
C12643 VPWR.n963 VGND 1.33431f
C12644 VPWR.n964 VGND 0.03811f
C12645 VPWR.t557 VGND 0.79335f
C12646 VPWR.n965 VGND 0.4327f
C12647 VPWR.t224 VGND 0.79335f
C12648 VPWR.n966 VGND 0.33651f
C12649 VPWR.n967 VGND 0.23859f
C12650 VPWR.t681 VGND 0.01165f
C12651 VPWR.t679 VGND 0.01165f
C12652 VPWR.n969 VGND 0.02558f
C12653 VPWR.t678 VGND 0.01165f
C12654 VPWR.t676 VGND 0.01165f
C12655 VPWR.n970 VGND 0.02554f
C12656 VPWR.t225 VGND 0.01165f
C12657 VPWR.t226 VGND 0.01165f
C12658 VPWR.n971 VGND 0.02554f
C12659 VPWR.n972 VGND 0.08473f
C12660 VPWR.n973 VGND 0.14784f
C12661 VPWR.n974 VGND 0.04681f
C12662 VPWR.n975 VGND 0.03438f
C12663 VPWR.t1461 VGND 0.01165f
C12664 VPWR.t1463 VGND 0.01165f
C12665 VPWR.n976 VGND 0.02558f
C12666 VPWR.n977 VGND 0.10491f
C12667 VPWR.n979 VGND 0.01326f
C12668 VPWR.n980 VGND 0.01553f
C12669 VPWR.n981 VGND 0.02237f
C12670 VPWR.t561 VGND 0.04641f
C12671 VPWR.n983 VGND 0.04961f
C12672 VPWR.t830 VGND 0.04651f
C12673 VPWR.n985 VGND 0.07408f
C12674 VPWR.n986 VGND 0.27291f
C12675 VPWR.n987 VGND 1.33431f
C12676 VPWR.n988 VGND 0.03811f
C12677 VPWR.t559 VGND 0.79335f
C12678 VPWR.n989 VGND 0.4327f
C12679 VPWR.t66 VGND 0.79335f
C12680 VPWR.n990 VGND 0.33651f
C12681 VPWR.n991 VGND 0.23859f
C12682 VPWR.t843 VGND 0.01165f
C12683 VPWR.t841 VGND 0.01165f
C12684 VPWR.n993 VGND 0.02558f
C12685 VPWR.t840 VGND 0.01165f
C12686 VPWR.t839 VGND 0.01165f
C12687 VPWR.n994 VGND 0.02554f
C12688 VPWR.t984 VGND 0.01165f
C12689 VPWR.t991 VGND 0.01165f
C12690 VPWR.n995 VGND 0.02554f
C12691 VPWR.n996 VGND 0.08473f
C12692 VPWR.n997 VGND 0.14784f
C12693 VPWR.n998 VGND 0.04681f
C12694 VPWR.n999 VGND 0.03438f
C12695 VPWR.t988 VGND 0.01165f
C12696 VPWR.t985 VGND 0.01165f
C12697 VPWR.n1000 VGND 0.02558f
C12698 VPWR.n1001 VGND 0.10491f
C12699 VPWR.n1003 VGND 0.01326f
C12700 VPWR.n1004 VGND 0.01553f
C12701 VPWR.n1005 VGND 0.02237f
C12702 VPWR.n1006 VGND 0.01137f
C12703 VPWR.n1007 VGND 0.01064f
C12704 VPWR.t1572 VGND 0.04651f
C12705 VPWR.t67 VGND 0.04651f
C12706 VPWR.n1008 VGND 0.13737f
C12707 VPWR.n1009 VGND 0.27291f
C12708 VPWR.n1010 VGND 1.33431f
C12709 VPWR.t416 VGND 0.04644f
C12710 VPWR.t829 VGND 0.04651f
C12711 VPWR.t418 VGND 0.04612f
C12712 VPWR.n1011 VGND 0.11958f
C12713 VPWR.t954 VGND 0.04559f
C12714 VPWR.n1012 VGND 0.05509f
C12715 VPWR.n1013 VGND 0.03811f
C12716 VPWR.t787 VGND 0.04389f
C12717 VPWR.n1014 VGND 0.04174f
C12718 VPWR.t693 VGND 0.01165f
C12719 VPWR.t919 VGND 0.01165f
C12720 VPWR.n1015 VGND 0.02546f
C12721 VPWR.t340 VGND 0.04078f
C12722 VPWR.n1016 VGND 0.06116f
C12723 VPWR.n1017 VGND 0.03811f
C12724 VPWR.t951 VGND 0.04646f
C12725 VPWR.n1018 VGND 0.05849f
C12726 VPWR.n1019 VGND 0.02237f
C12727 VPWR.n1020 VGND 0.03811f
C12728 VPWR.t921 VGND 0.01165f
C12729 VPWR.t923 VGND 0.01165f
C12730 VPWR.n1022 VGND 0.02546f
C12731 VPWR.n1023 VGND 0.03731f
C12732 VPWR.n1025 VGND 0.02858f
C12733 VPWR.n1026 VGND 0.02858f
C12734 VPWR.n1027 VGND 0.03811f
C12735 VPWR.t1733 VGND 0.01165f
C12736 VPWR.t697 VGND 0.01165f
C12737 VPWR.n1029 VGND 0.02546f
C12738 VPWR.n1030 VGND 0.02931f
C12739 VPWR.t956 VGND 0.01165f
C12740 VPWR.t932 VGND 0.01165f
C12741 VPWR.n1031 VGND 0.02546f
C12742 VPWR.n1032 VGND 0.03239f
C12743 VPWR.n1034 VGND 0.03459f
C12744 VPWR.n1035 VGND 0.01305f
C12745 VPWR.t1799 VGND 0.03908f
C12746 VPWR.t415 VGND 0.08792f
C12747 VPWR.t828 VGND 0.10257f
C12748 VPWR.t417 VGND 0.19049f
C12749 VPWR.t950 VGND 0.1025f
C12750 VPWR.t922 VGND 0.11635f
C12751 VPWR.t920 VGND 0.11311f
C12752 VPWR.t918 VGND 0.1809f
C12753 VPWR.t692 VGND 0.15386f
C12754 VPWR.t339 VGND 0.10257f
C12755 VPWR.t696 VGND 0.10257f
C12756 VPWR.t931 VGND 0.10257f
C12757 VPWR.t1732 VGND 0.10257f
C12758 VPWR.t955 VGND 0.10257f
C12759 VPWR.t786 VGND 0.10257f
C12760 VPWR.t953 VGND 0.10135f
C12761 VPWR.n1037 VGND 0.3486f
C12762 VPWR.n1038 VGND 0.14164f
C12763 VPWR.n1039 VGND 0.01553f
C12764 VPWR.n1040 VGND 0.02858f
C12765 VPWR.n1041 VGND 0.03438f
C12766 VPWR.n1043 VGND 0.05169f
C12767 VPWR.n1044 VGND 0.25738f
C12768 VPWR.n1045 VGND 1.33431f
C12769 VPWR.t727 VGND 0.04569f
C12770 VPWR.t769 VGND 0.04556f
C12771 VPWR.t233 VGND 0.04646f
C12772 VPWR.n1046 VGND 0.06475f
C12773 VPWR.t783 VGND 0.04436f
C12774 VPWR.t386 VGND 0.04436f
C12775 VPWR.n1047 VGND 0.08048f
C12776 VPWR.n1048 VGND 0.03811f
C12777 VPWR.n1050 VGND 0.03811f
C12778 VPWR.t665 VGND 0.01165f
C12779 VPWR.t1872 VGND 0.01165f
C12780 VPWR.n1051 VGND 0.02546f
C12781 VPWR.t387 VGND 0.01165f
C12782 VPWR.t1751 VGND 0.01165f
C12783 VPWR.n1052 VGND 0.02546f
C12784 VPWR.n1053 VGND 0.05187f
C12785 VPWR.t1753 VGND 0.04646f
C12786 VPWR.t1868 VGND 0.04646f
C12787 VPWR.n1054 VGND 0.10708f
C12788 VPWR.n1055 VGND 0.02237f
C12789 VPWR.n1056 VGND 0.03811f
C12790 VPWR.t1759 VGND 0.01165f
C12791 VPWR.t342 VGND 0.01165f
C12792 VPWR.n1058 VGND 0.02546f
C12793 VPWR.t228 VGND 0.01165f
C12794 VPWR.t232 VGND 0.01165f
C12795 VPWR.n1059 VGND 0.02546f
C12796 VPWR.n1060 VGND 0.05862f
C12797 VPWR.n1062 VGND 0.03811f
C12798 VPWR.n1063 VGND 0.03811f
C12799 VPWR.n1064 VGND 0.03811f
C12800 VPWR.t153 VGND 0.01165f
C12801 VPWR.t780 VGND 0.01165f
C12802 VPWR.n1066 VGND 0.02546f
C12803 VPWR.t382 VGND 0.01165f
C12804 VPWR.t381 VGND 0.01165f
C12805 VPWR.n1067 VGND 0.02546f
C12806 VPWR.n1068 VGND 0.05187f
C12807 VPWR.n1071 VGND 0.03811f
C12808 VPWR.n1072 VGND 0.02858f
C12809 VPWR.t152 VGND 0.79335f
C12810 VPWR.n1074 VGND 0.4327f
C12811 VPWR.t227 VGND 0.79335f
C12812 VPWR.n1075 VGND 0.33651f
C12813 VPWR.n1076 VGND 0.23646f
C12814 VPWR.n1077 VGND 0.01553f
C12815 VPWR.n1078 VGND 0.02858f
C12816 VPWR.n1079 VGND 0.03459f
C12817 VPWR.n1081 VGND 0.04738f
C12818 VPWR.n1082 VGND 0.06418f
C12819 VPWR.n1083 VGND 0.25717f
C12820 VPWR.n1084 VGND 1.33431f
C12821 VPWR.t423 VGND 0.04641f
C12822 VPWR.t779 VGND 0.04641f
C12823 VPWR.n1085 VGND 0.01137f
C12824 VPWR.t677 VGND 0.04436f
C12825 VPWR.t1462 VGND 0.04436f
C12826 VPWR.n1086 VGND 0.08048f
C12827 VPWR.n1087 VGND 0.03811f
C12828 VPWR.n1089 VGND 0.03811f
C12829 VPWR.t682 VGND 0.01165f
C12830 VPWR.t1754 VGND 0.01165f
C12831 VPWR.n1090 VGND 0.02546f
C12832 VPWR.t1831 VGND 0.01165f
C12833 VPWR.t1869 VGND 0.01165f
C12834 VPWR.n1091 VGND 0.02546f
C12835 VPWR.n1092 VGND 0.05187f
C12836 VPWR.t1870 VGND 0.04646f
C12837 VPWR.t1750 VGND 0.04646f
C12838 VPWR.n1093 VGND 0.10708f
C12839 VPWR.n1094 VGND 0.02237f
C12840 VPWR.n1095 VGND 0.03811f
C12841 VPWR.t231 VGND 0.01165f
C12842 VPWR.t930 VGND 0.01165f
C12843 VPWR.n1097 VGND 0.02546f
C12844 VPWR.t1871 VGND 0.01165f
C12845 VPWR.t1761 VGND 0.01165f
C12846 VPWR.n1098 VGND 0.02546f
C12847 VPWR.n1099 VGND 0.05862f
C12848 VPWR.n1101 VGND 0.03811f
C12849 VPWR.n1102 VGND 0.03811f
C12850 VPWR.n1103 VGND 0.03811f
C12851 VPWR.t683 VGND 0.01165f
C12852 VPWR.t680 VGND 0.01165f
C12853 VPWR.n1105 VGND 0.02546f
C12854 VPWR.t1830 VGND 0.01165f
C12855 VPWR.t1832 VGND 0.01165f
C12856 VPWR.n1106 VGND 0.02546f
C12857 VPWR.n1107 VGND 0.05187f
C12858 VPWR.n1110 VGND 0.03811f
C12859 VPWR.n1111 VGND 0.02858f
C12860 VPWR.t230 VGND 0.79335f
C12861 VPWR.n1113 VGND 0.4327f
C12862 VPWR.t778 VGND 0.79335f
C12863 VPWR.n1114 VGND 0.33651f
C12864 VPWR.n1115 VGND 0.23859f
C12865 VPWR.n1116 VGND 0.01553f
C12866 VPWR.n1117 VGND 0.02858f
C12867 VPWR.n1118 VGND 0.03459f
C12868 VPWR.n1120 VGND 0.09381f
C12869 VPWR.n1121 VGND 0.26132f
C12870 VPWR.n1122 VGND 1.33431f
C12871 VPWR.t842 VGND 0.04436f
C12872 VPWR.t986 VGND 0.04436f
C12873 VPWR.n1123 VGND 0.08048f
C12874 VPWR.n1124 VGND 0.03811f
C12875 VPWR.n1126 VGND 0.03811f
C12876 VPWR.t837 VGND 0.01165f
C12877 VPWR.t1758 VGND 0.01165f
C12878 VPWR.n1127 VGND 0.02546f
C12879 VPWR.t987 VGND 0.01165f
C12880 VPWR.t949 VGND 0.01165f
C12881 VPWR.n1128 VGND 0.02546f
C12882 VPWR.n1129 VGND 0.05187f
C12883 VPWR.t1755 VGND 0.04646f
C12884 VPWR.t917 VGND 0.04646f
C12885 VPWR.n1130 VGND 0.10708f
C12886 VPWR.n1131 VGND 0.02237f
C12887 VPWR.n1132 VGND 0.03811f
C12888 VPWR.t1760 VGND 0.01165f
C12889 VPWR.t344 VGND 0.01165f
C12890 VPWR.n1134 VGND 0.02546f
C12891 VPWR.t952 VGND 0.01165f
C12892 VPWR.t1749 VGND 0.01165f
C12893 VPWR.n1135 VGND 0.02546f
C12894 VPWR.n1136 VGND 0.05862f
C12895 VPWR.n1138 VGND 0.03811f
C12896 VPWR.n1139 VGND 0.03811f
C12897 VPWR.n1140 VGND 0.03811f
C12898 VPWR.t838 VGND 0.01165f
C12899 VPWR.t836 VGND 0.01165f
C12900 VPWR.n1142 VGND 0.02546f
C12901 VPWR.t990 VGND 0.01165f
C12902 VPWR.t989 VGND 0.01165f
C12903 VPWR.n1143 VGND 0.02546f
C12904 VPWR.n1144 VGND 0.05187f
C12905 VPWR.n1147 VGND 0.03811f
C12906 VPWR.n1148 VGND 0.02858f
C12907 VPWR.t343 VGND 0.60858f
C12908 VPWR.n1150 VGND 0.34819f
C12909 VPWR.t916 VGND 0.60858f
C12910 VPWR.n1151 VGND 0.27284f
C12911 VPWR.n1152 VGND 0.22873f
C12912 VPWR.n1153 VGND 0.34967f
C12913 VPWR.n1154 VGND 5.08436f
C12914 VPWR.n1155 VGND 0.82079f
C12915 VPWR.n1156 VGND 0.82079f
C12916 VPWR.n1157 VGND -0.05416f
C12917 VPWR.n1158 VGND 0.02774f
C12918 VPWR.t1161 VGND 0.02709f
C12919 VPWR.t1244 VGND 0.02407f
C12920 VPWR.n1160 VGND 0.07442f
C12921 VPWR.t1398 VGND 0.118f
C12922 VPWR.t1391 VGND 0.06383f
C12923 VPWR.t1107 VGND 0.07496f
C12924 VPWR.t1399 VGND 0.02709f
C12925 VPWR.t1108 VGND 0.02407f
C12926 VPWR.n1161 VGND 0.07442f
C12927 VPWR.n1163 VGND 0.088f
C12928 VPWR.t1160 VGND 0.09722f
C12929 VPWR.t1121 VGND 0.06383f
C12930 VPWR.t1243 VGND 0.07496f
C12931 VPWR.t1424 VGND 0.09722f
C12932 VPWR.t1263 VGND 0.02709f
C12933 VPWR.t1257 VGND 0.02407f
C12934 VPWR.n1164 VGND 0.07442f
C12935 VPWR.n1165 VGND 0.05649f
C12936 VPWR.n1166 VGND 0.10954f
C12937 VPWR.n1167 VGND -0.01517f
C12938 VPWR.n1168 VGND 0.06791f
C12939 VPWR.n1170 VGND 0.04424f
C12940 VPWR.n1171 VGND 0.0512f
C12941 VPWR.n1173 VGND 0.02474f
C12942 VPWR.t1325 VGND 0.02178f
C12943 VPWR.n1175 VGND 0.04654f
C12944 VPWR.t1669 VGND 0.02407f
C12945 VPWR.n1176 VGND 0.03816f
C12946 VPWR.t1536 VGND 0.07496f
C12947 VPWR.n1177 VGND 0.02474f
C12948 VPWR.t1449 VGND 0.02178f
C12949 VPWR.n1179 VGND 0.04654f
C12950 VPWR.t1537 VGND 0.02407f
C12951 VPWR.n1180 VGND 0.03816f
C12952 VPWR.n1181 VGND 0.02474f
C12953 VPWR.t1322 VGND 0.02178f
C12954 VPWR.n1183 VGND 0.04654f
C12955 VPWR.t454 VGND 0.02407f
C12956 VPWR.n1184 VGND 0.03816f
C12957 VPWR.t1185 VGND 0.118f
C12958 VPWR.t1170 VGND 0.06383f
C12959 VPWR.t844 VGND 0.07496f
C12960 VPWR.n1185 VGND 0.02474f
C12961 VPWR.t1186 VGND 0.02178f
C12962 VPWR.n1187 VGND 0.04654f
C12963 VPWR.t845 VGND 0.02407f
C12964 VPWR.n1188 VGND 0.03816f
C12965 VPWR.n1189 VGND -0.05607f
C12966 VPWR.n1191 VGND 0.088f
C12967 VPWR.t1321 VGND 0.09722f
C12968 VPWR.t1301 VGND 0.06383f
C12969 VPWR.t453 VGND 0.07496f
C12970 VPWR.t1430 VGND 0.06383f
C12971 VPWR.t1448 VGND 0.09722f
C12972 VPWR.n1192 VGND 0.088f
C12973 VPWR.n1194 VGND 0.0512f
C12974 VPWR.n1197 VGND 0.0512f
C12975 VPWR.n1199 VGND 0.088f
C12976 VPWR.t1219 VGND 0.09722f
C12977 VPWR.t1086 VGND 0.06383f
C12978 VPWR.t728 VGND 0.07496f
C12979 VPWR.n1200 VGND 0.02474f
C12980 VPWR.t1220 VGND 0.02178f
C12981 VPWR.n1202 VGND 0.04654f
C12982 VPWR.t729 VGND 0.02407f
C12983 VPWR.n1203 VGND 0.03816f
C12984 VPWR.n1205 VGND 0.088f
C12985 VPWR.t1324 VGND 0.09722f
C12986 VPWR.t1196 VGND 0.06383f
C12987 VPWR.t1668 VGND 0.07496f
C12988 VPWR.t1094 VGND 0.09722f
C12989 VPWR.n1206 VGND 0.02474f
C12990 VPWR.t1347 VGND 0.02178f
C12991 VPWR.n1208 VGND 0.04654f
C12992 VPWR.t915 VGND 0.02407f
C12993 VPWR.n1209 VGND 0.03816f
C12994 VPWR.n1211 VGND 0.02474f
C12995 VPWR.t1095 VGND 0.02178f
C12996 VPWR.n1213 VGND 0.04654f
C12997 VPWR.t1836 VGND 0.02407f
C12998 VPWR.n1214 VGND 0.03816f
C12999 VPWR.t1353 VGND 0.06383f
C13000 VPWR.t1835 VGND 0.07496f
C13001 VPWR.t1357 VGND 0.09722f
C13002 VPWR.n1215 VGND 0.02474f
C13003 VPWR.t1217 VGND 0.02178f
C13004 VPWR.n1217 VGND 0.04654f
C13005 VPWR.t515 VGND 0.02407f
C13006 VPWR.n1218 VGND 0.03816f
C13007 VPWR.n1220 VGND 0.02474f
C13008 VPWR.t1358 VGND 0.02178f
C13009 VPWR.n1222 VGND 0.04654f
C13010 VPWR.t1570 VGND 0.02407f
C13011 VPWR.n1223 VGND 0.03816f
C13012 VPWR.t1231 VGND 0.06383f
C13013 VPWR.t1569 VGND 0.07496f
C13014 VPWR.t1113 VGND 0.09722f
C13015 VPWR.n1224 VGND 0.02474f
C13016 VPWR.t1386 VGND 0.02178f
C13017 VPWR.n1226 VGND 0.04654f
C13018 VPWR.t1563 VGND 0.02407f
C13019 VPWR.n1227 VGND 0.03816f
C13020 VPWR.n1228 VGND -0.01517f
C13021 VPWR.n1229 VGND 0.0534f
C13022 VPWR.n1230 VGND 0.0746f
C13023 VPWR.n1231 VGND -0.01517f
C13024 VPWR.n1232 VGND 0.0512f
C13025 VPWR.n1234 VGND 0.06791f
C13026 VPWR.n1236 VGND 0.02774f
C13027 VPWR.t1378 VGND 0.02709f
C13028 VPWR.t1370 VGND 0.02407f
C13029 VPWR.n1238 VGND 0.07442f
C13030 VPWR.t1369 VGND 0.07496f
C13031 VPWR.t1089 VGND 0.02709f
C13032 VPWR.t1212 VGND 0.02407f
C13033 VPWR.n1239 VGND 0.07442f
C13034 VPWR.n1240 VGND 0.02533f
C13035 VPWR.n1241 VGND 0.03003f
C13036 VPWR.t1083 VGND 0.01009f
C13037 VPWR.n1243 VGND 0.02251f
C13038 VPWR.n1244 VGND 0.02292f
C13039 VPWR.n1245 VGND 0.14299f
C13040 VPWR.n1246 VGND 0.05649f
C13041 VPWR.n1247 VGND 0.05649f
C13042 VPWR.t1187 VGND 0.01009f
C13043 VPWR.n1248 VGND 0.02251f
C13044 VPWR.n1249 VGND 0.02292f
C13045 VPWR.n1250 VGND 0.14299f
C13046 VPWR.t1340 VGND 0.01009f
C13047 VPWR.n1251 VGND 0.02251f
C13048 VPWR.n1252 VGND 0.02292f
C13049 VPWR.t1082 VGND 0.02709f
C13050 VPWR.t1460 VGND 0.02407f
C13051 VPWR.n1253 VGND 0.07442f
C13052 VPWR.t1440 VGND 0.07496f
C13053 VPWR.t1339 VGND 0.02709f
C13054 VPWR.t1441 VGND 0.02407f
C13055 VPWR.n1254 VGND 0.07442f
C13056 VPWR.n1256 VGND 0.02533f
C13057 VPWR.n1257 VGND 0.03003f
C13058 VPWR.n1258 VGND 0.02774f
C13059 VPWR.n1259 VGND 0.05649f
C13060 VPWR.t1209 VGND 0.02709f
C13061 VPWR.t1282 VGND 0.02407f
C13062 VPWR.n1260 VGND 0.07442f
C13063 VPWR.t1177 VGND 0.07496f
C13064 VPWR.t1183 VGND 0.02709f
C13065 VPWR.t1178 VGND 0.02407f
C13066 VPWR.n1261 VGND 0.07442f
C13067 VPWR.n1262 VGND 0.05649f
C13068 VPWR.n1263 VGND 0.10954f
C13069 VPWR.n1264 VGND 0.05649f
C13070 VPWR.t1364 VGND 0.02709f
C13071 VPWR.t1433 VGND 0.02407f
C13072 VPWR.n1265 VGND 0.07442f
C13073 VPWR.t1401 VGND 0.07496f
C13074 VPWR.t1314 VGND 0.02709f
C13075 VPWR.t1402 VGND 0.02407f
C13076 VPWR.n1266 VGND 0.07442f
C13077 VPWR.n1267 VGND 0.05649f
C13078 VPWR.n1268 VGND 0.10954f
C13079 VPWR.n1269 VGND 0.05649f
C13080 VPWR.t1155 VGND 0.02709f
C13081 VPWR.t1285 VGND 0.02407f
C13082 VPWR.n1270 VGND 0.07442f
C13083 VPWR.t1137 VGND 0.07496f
C13084 VPWR.t1143 VGND 0.02709f
C13085 VPWR.t1138 VGND 0.02407f
C13086 VPWR.n1271 VGND 0.07442f
C13087 VPWR.n1272 VGND 0.01938f
C13088 VPWR.n1273 VGND 0.01938f
C13089 VPWR.n1274 VGND 0.01938f
C13090 VPWR.n1275 VGND 0.01938f
C13091 VPWR.n1276 VGND 0.14299f
C13092 VPWR.t1425 VGND 0.02709f
C13093 VPWR.t1361 VGND 0.02407f
C13094 VPWR.n1277 VGND 0.07442f
C13095 VPWR.t1290 VGND 0.06383f
C13096 VPWR.t1360 VGND 0.07496f
C13097 VPWR.t1407 VGND 0.06383f
C13098 VPWR.t1142 VGND 0.09722f
C13099 VPWR.n1278 VGND 0.088f
C13100 VPWR.n1281 VGND 0.05649f
C13101 VPWR.n1282 VGND 0.02533f
C13102 VPWR.n1283 VGND 0.03003f
C13103 VPWR.t1248 VGND 0.01009f
C13104 VPWR.n1285 VGND 0.02251f
C13105 VPWR.n1286 VGND 0.02292f
C13106 VPWR.n1287 VGND 0.02158f
C13107 VPWR.n1288 VGND 0.02533f
C13108 VPWR.n1289 VGND 0.01601f
C13109 VPWR.t1390 VGND 0.01009f
C13110 VPWR.n1290 VGND 0.02251f
C13111 VPWR.n1291 VGND 0.02292f
C13112 VPWR.n1292 VGND 0.01481f
C13113 VPWR.n1294 VGND 0.01444f
C13114 VPWR.n1295 VGND 0.02434f
C13115 VPWR.n1296 VGND 0.0267f
C13116 VPWR.n1297 VGND 0.02764f
C13117 VPWR.n1298 VGND 0.02533f
C13118 VPWR.n1299 VGND 0.03003f
C13119 VPWR.t1120 VGND 0.01009f
C13120 VPWR.n1301 VGND 0.02251f
C13121 VPWR.n1302 VGND 0.02292f
C13122 VPWR.n1303 VGND 0.02434f
C13123 VPWR.n1304 VGND 0.0267f
C13124 VPWR.n1305 VGND 0.01444f
C13125 VPWR.n1307 VGND 0.01481f
C13126 VPWR.n1308 VGND 0.01938f
C13127 VPWR.n1309 VGND 0.19291f
C13128 VPWR.n1310 VGND 0.14299f
C13129 VPWR.n1311 VGND 0.01938f
C13130 VPWR.n1312 VGND 0.01481f
C13131 VPWR.n1314 VGND 0.01444f
C13132 VPWR.n1315 VGND 0.02434f
C13133 VPWR.n1316 VGND 0.0267f
C13134 VPWR.n1317 VGND 0.02774f
C13135 VPWR.n1318 VGND 0.02533f
C13136 VPWR.n1319 VGND 0.03003f
C13137 VPWR.t1289 VGND 0.01009f
C13138 VPWR.n1321 VGND 0.02251f
C13139 VPWR.n1322 VGND 0.02292f
C13140 VPWR.n1323 VGND 0.01938f
C13141 VPWR.n1324 VGND 0.01481f
C13142 VPWR.n1326 VGND 0.01444f
C13143 VPWR.n1327 VGND 0.02434f
C13144 VPWR.n1328 VGND 0.0267f
C13145 VPWR.n1329 VGND 0.02774f
C13146 VPWR.n1330 VGND 0.02533f
C13147 VPWR.n1331 VGND 0.03003f
C13148 VPWR.t1406 VGND 0.01009f
C13149 VPWR.n1333 VGND 0.02251f
C13150 VPWR.n1334 VGND 0.02292f
C13151 VPWR.n1335 VGND 0.02434f
C13152 VPWR.n1336 VGND 0.0267f
C13153 VPWR.n1337 VGND 0.01444f
C13154 VPWR.n1339 VGND 0.01481f
C13155 VPWR.n1340 VGND 0.01938f
C13156 VPWR.n1341 VGND 0.14299f
C13157 VPWR.n1342 VGND 0.14299f
C13158 VPWR.n1343 VGND 0.14299f
C13159 VPWR.n1344 VGND 0.14299f
C13160 VPWR.n1345 VGND 0.14299f
C13161 VPWR.n1346 VGND 0.14299f
C13162 VPWR.n1347 VGND 0.01938f
C13163 VPWR.n1348 VGND 0.01938f
C13164 VPWR.n1349 VGND 0.02434f
C13165 VPWR.n1350 VGND 0.0267f
C13166 VPWR.n1351 VGND 0.01481f
C13167 VPWR.n1353 VGND 0.01444f
C13168 VPWR.t1315 VGND 0.01009f
C13169 VPWR.n1354 VGND 0.02251f
C13170 VPWR.n1355 VGND 0.02292f
C13171 VPWR.n1357 VGND 0.02533f
C13172 VPWR.n1358 VGND 0.03003f
C13173 VPWR.n1359 VGND 0.02774f
C13174 VPWR.n1360 VGND 0.02434f
C13175 VPWR.n1361 VGND 0.0267f
C13176 VPWR.n1362 VGND 0.01481f
C13177 VPWR.n1364 VGND 0.01444f
C13178 VPWR.t1162 VGND 0.01009f
C13179 VPWR.n1365 VGND 0.02251f
C13180 VPWR.n1366 VGND 0.02292f
C13181 VPWR.n1368 VGND 0.02533f
C13182 VPWR.n1369 VGND 0.03003f
C13183 VPWR.n1370 VGND 0.02774f
C13184 VPWR.n1371 VGND 0.02434f
C13185 VPWR.n1372 VGND 0.0267f
C13186 VPWR.n1373 VGND 0.01481f
C13187 VPWR.n1375 VGND 0.01444f
C13188 VPWR.t1445 VGND 0.01009f
C13189 VPWR.n1376 VGND 0.02251f
C13190 VPWR.n1377 VGND 0.02292f
C13191 VPWR.n1379 VGND 0.02533f
C13192 VPWR.n1380 VGND 0.03003f
C13193 VPWR.n1381 VGND 0.02774f
C13194 VPWR.n1382 VGND 0.02434f
C13195 VPWR.n1383 VGND 0.0267f
C13196 VPWR.n1384 VGND 0.01481f
C13197 VPWR.n1386 VGND 0.01444f
C13198 VPWR.t1411 VGND 0.01009f
C13199 VPWR.n1387 VGND 0.02251f
C13200 VPWR.n1388 VGND 0.02292f
C13201 VPWR.n1390 VGND 0.02533f
C13202 VPWR.n1391 VGND 0.03003f
C13203 VPWR.n1392 VGND 0.02774f
C13204 VPWR.n1393 VGND 0.02434f
C13205 VPWR.n1394 VGND 0.0267f
C13206 VPWR.n1395 VGND 0.01481f
C13207 VPWR.n1397 VGND 0.01444f
C13208 VPWR.t1179 VGND 0.01009f
C13209 VPWR.n1398 VGND 0.02251f
C13210 VPWR.n1399 VGND 0.02292f
C13211 VPWR.n1401 VGND 0.02533f
C13212 VPWR.n1402 VGND 0.03003f
C13213 VPWR.n1403 VGND 0.02774f
C13214 VPWR.n1404 VGND 0.02434f
C13215 VPWR.n1405 VGND 0.0267f
C13216 VPWR.n1406 VGND 0.01481f
C13217 VPWR.n1408 VGND 0.01444f
C13218 VPWR.t1164 VGND 0.01009f
C13219 VPWR.n1409 VGND 0.02251f
C13220 VPWR.n1410 VGND 0.02292f
C13221 VPWR.n1412 VGND 0.02533f
C13222 VPWR.n1413 VGND 0.03003f
C13223 VPWR.n1414 VGND 0.02774f
C13224 VPWR.n1415 VGND 0.05649f
C13225 VPWR.n1416 VGND 0.0534f
C13226 VPWR.n1417 VGND 0.0534f
C13227 VPWR.t1300 VGND 0.01009f
C13228 VPWR.n1418 VGND 0.02252f
C13229 VPWR.n1419 VGND 0.01543f
C13230 VPWR.n1420 VGND 0.05077f
C13231 VPWR.n1421 VGND 0.07925f
C13232 VPWR.n1422 VGND 0.04424f
C13233 VPWR.n1423 VGND 0.0746f
C13234 VPWR.t1169 VGND 0.01009f
C13235 VPWR.n1424 VGND 0.02252f
C13236 VPWR.n1425 VGND 0.01543f
C13237 VPWR.n1426 VGND 0.05077f
C13238 VPWR.n1427 VGND 0.06312f
C13239 VPWR.n1428 VGND 0.05271f
C13240 VPWR.n1429 VGND 0.04424f
C13241 VPWR.n1430 VGND 0.0534f
C13242 VPWR.n1431 VGND 0.04424f
C13243 VPWR.n1432 VGND 0.0534f
C13244 VPWR.n1433 VGND 0.0746f
C13245 VPWR.t1429 VGND 0.01009f
C13246 VPWR.n1434 VGND 0.02252f
C13247 VPWR.n1435 VGND 0.01543f
C13248 VPWR.n1436 VGND 0.05077f
C13249 VPWR.n1437 VGND 0.07925f
C13250 VPWR.n1438 VGND 0.0746f
C13251 VPWR.t1085 VGND 0.01009f
C13252 VPWR.n1439 VGND 0.02252f
C13253 VPWR.n1440 VGND 0.01543f
C13254 VPWR.n1441 VGND 0.05077f
C13255 VPWR.n1442 VGND 0.07925f
C13256 VPWR.n1443 VGND 0.0746f
C13257 VPWR.t1195 VGND 0.01009f
C13258 VPWR.n1444 VGND 0.02252f
C13259 VPWR.n1445 VGND 0.01543f
C13260 VPWR.n1446 VGND 0.05077f
C13261 VPWR.n1447 VGND 0.07925f
C13262 VPWR.n1448 VGND 0.0746f
C13263 VPWR.t1350 VGND 0.01009f
C13264 VPWR.n1449 VGND 0.02252f
C13265 VPWR.n1450 VGND 0.01543f
C13266 VPWR.n1451 VGND 0.05077f
C13267 VPWR.n1452 VGND 0.07925f
C13268 VPWR.n1453 VGND 0.0746f
C13269 VPWR.t1352 VGND 0.01009f
C13270 VPWR.n1454 VGND 0.02252f
C13271 VPWR.n1455 VGND 0.01543f
C13272 VPWR.n1456 VGND 0.05077f
C13273 VPWR.n1457 VGND 0.07925f
C13274 VPWR.n1458 VGND 0.0746f
C13275 VPWR.t1200 VGND 0.01009f
C13276 VPWR.n1459 VGND 0.02252f
C13277 VPWR.n1460 VGND 0.01543f
C13278 VPWR.n1461 VGND 0.05077f
C13279 VPWR.n1462 VGND 0.07925f
C13280 VPWR.t1348 VGND 0.01009f
C13281 VPWR.n1463 VGND 0.02252f
C13282 VPWR.n1464 VGND 0.01543f
C13283 VPWR.n1465 VGND 0.05077f
C13284 VPWR.n1466 VGND 0.07925f
C13285 VPWR.n1467 VGND 0.0746f
C13286 VPWR.t1230 VGND 0.01009f
C13287 VPWR.n1468 VGND 0.02252f
C13288 VPWR.n1469 VGND 0.01543f
C13289 VPWR.n1470 VGND 0.05077f
C13290 VPWR.n1471 VGND 0.07925f
C13291 VPWR.n1472 VGND 0.0746f
C13292 VPWR.n1473 VGND 0.04424f
C13293 VPWR.n1474 VGND 0.0534f
C13294 VPWR.n1475 VGND 0.04424f
C13295 VPWR.n1476 VGND 0.0534f
C13296 VPWR.n1477 VGND 0.04424f
C13297 VPWR.n1478 VGND 0.0534f
C13298 VPWR.n1479 VGND 0.04424f
C13299 VPWR.n1480 VGND 0.0534f
C13300 VPWR.n1481 VGND 0.04424f
C13301 VPWR.n1482 VGND 0.10954f
C13302 VPWR.n1483 VGND 0.06791f
C13303 VPWR.n1484 VGND -0.01517f
C13304 VPWR.n1488 VGND 0.088f
C13305 VPWR.t1154 VGND 0.09722f
C13306 VPWR.t1165 VGND 0.06383f
C13307 VPWR.t1284 VGND 0.07496f
C13308 VPWR.t1180 VGND 0.06383f
C13309 VPWR.t1313 VGND 0.09722f
C13310 VPWR.n1489 VGND 0.088f
C13311 VPWR.n1493 VGND -0.01517f
C13312 VPWR.n1494 VGND 0.06791f
C13313 VPWR.n1495 VGND 0.06791f
C13314 VPWR.n1496 VGND -0.01517f
C13315 VPWR.n1500 VGND 0.088f
C13316 VPWR.t1363 VGND 0.09722f
C13317 VPWR.t1412 VGND 0.06383f
C13318 VPWR.t1432 VGND 0.07496f
C13319 VPWR.t1446 VGND 0.06383f
C13320 VPWR.t1182 VGND 0.09722f
C13321 VPWR.n1501 VGND 0.088f
C13322 VPWR.n1505 VGND -0.01517f
C13323 VPWR.n1506 VGND 0.06791f
C13324 VPWR.n1507 VGND 0.06791f
C13325 VPWR.n1508 VGND 0.06791f
C13326 VPWR.n1509 VGND 0.06791f
C13327 VPWR.n1510 VGND -0.01517f
C13328 VPWR.n1514 VGND 0.088f
C13329 VPWR.t1208 VGND 0.09722f
C13330 VPWR.t1163 VGND 0.06383f
C13331 VPWR.t1281 VGND 0.07496f
C13332 VPWR.t1316 VGND 0.06383f
C13333 VPWR.t1338 VGND 0.09722f
C13334 VPWR.n1515 VGND 0.088f
C13335 VPWR.n1519 VGND 0.05649f
C13336 VPWR.n1523 VGND 0.088f
C13337 VPWR.t1081 VGND 0.09722f
C13338 VPWR.t1341 VGND 0.06383f
C13339 VPWR.t1459 VGND 0.07496f
C13340 VPWR.t1239 VGND 0.06383f
C13341 VPWR.t1377 VGND 0.09722f
C13342 VPWR.t1344 VGND 0.02709f
C13343 VPWR.t1336 VGND 0.02407f
C13344 VPWR.n1524 VGND 0.07442f
C13345 VPWR.n1526 VGND 0.088f
C13346 VPWR.t1335 VGND 0.07496f
C13347 VPWR.t1214 VGND 0.06383f
C13348 VPWR.t1343 VGND 0.09722f
C13349 VPWR.t1103 VGND 0.02709f
C13350 VPWR.t1204 VGND 0.02407f
C13351 VPWR.n1527 VGND 0.07442f
C13352 VPWR.n1531 VGND 0.088f
C13353 VPWR.t1203 VGND 0.07496f
C13354 VPWR.t1188 VGND 0.06383f
C13355 VPWR.t1102 VGND 0.09722f
C13356 VPWR.n1532 VGND 0.088f
C13357 VPWR.n1535 VGND 0.05649f
C13358 VPWR.n1537 VGND 0.02533f
C13359 VPWR.n1538 VGND 0.03003f
C13360 VPWR.n1539 VGND 0.02774f
C13361 VPWR.n1540 VGND 0.02434f
C13362 VPWR.n1541 VGND 0.0267f
C13363 VPWR.n1542 VGND 0.01444f
C13364 VPWR.n1544 VGND 0.01481f
C13365 VPWR.n1545 VGND 0.01938f
C13366 VPWR.n1546 VGND 0.14299f
C13367 VPWR.n1547 VGND 0.14299f
C13368 VPWR.n1548 VGND 0.01938f
C13369 VPWR.n1549 VGND 0.01481f
C13370 VPWR.n1551 VGND 0.01444f
C13371 VPWR.n1552 VGND 0.02434f
C13372 VPWR.n1553 VGND 0.0267f
C13373 VPWR.n1554 VGND 0.02774f
C13374 VPWR.n1555 VGND 0.02533f
C13375 VPWR.n1556 VGND 0.03003f
C13376 VPWR.t1213 VGND 0.01009f
C13377 VPWR.n1558 VGND 0.02251f
C13378 VPWR.n1559 VGND 0.02292f
C13379 VPWR.n1560 VGND 0.01938f
C13380 VPWR.n1561 VGND 0.01481f
C13381 VPWR.n1563 VGND 0.01444f
C13382 VPWR.n1564 VGND 0.02434f
C13383 VPWR.n1565 VGND 0.0267f
C13384 VPWR.n1566 VGND 0.02774f
C13385 VPWR.n1567 VGND 0.02533f
C13386 VPWR.n1568 VGND 0.03003f
C13387 VPWR.t1238 VGND 0.01009f
C13388 VPWR.n1570 VGND 0.02251f
C13389 VPWR.n1571 VGND 0.02292f
C13390 VPWR.n1572 VGND 0.02434f
C13391 VPWR.n1573 VGND 0.0267f
C13392 VPWR.n1574 VGND 0.01444f
C13393 VPWR.n1576 VGND 0.01481f
C13394 VPWR.n1577 VGND 0.01938f
C13395 VPWR.n1578 VGND 0.17208f
C13396 VPWR.n1579 VGND 0.02066f
C13397 VPWR.n1580 VGND 0.01481f
C13398 VPWR.n1582 VGND 0.01444f
C13399 VPWR.n1583 VGND 0.02434f
C13400 VPWR.n1584 VGND 0.0267f
C13401 VPWR.n1585 VGND 0.05635f
C13402 VPWR.n1587 VGND 0.06192f
C13403 VPWR.t1211 VGND 0.10842f
C13404 VPWR.t1084 VGND 0.06383f
C13405 VPWR.t1088 VGND 0.09722f
C13406 VPWR.n1588 VGND 0.088f
C13407 VPWR.n1591 VGND 0.05649f
C13408 VPWR.n1593 VGND -0.01517f
C13409 VPWR.n1594 VGND 0.06791f
C13410 VPWR.n1595 VGND 0.06791f
C13411 VPWR.n1596 VGND 0.06791f
C13412 VPWR.n1597 VGND -0.01517f
C13413 VPWR.t1099 VGND 0.01009f
C13414 VPWR.n1598 VGND 0.02252f
C13415 VPWR.n1599 VGND 0.01543f
C13416 VPWR.n1600 VGND 0.05077f
C13417 VPWR.n1601 VGND 0.07925f
C13418 VPWR.t1371 VGND 0.01009f
C13419 VPWR.n1602 VGND 0.02252f
C13420 VPWR.n1603 VGND 0.01543f
C13421 VPWR.n1604 VGND 0.05077f
C13422 VPWR.n1605 VGND 0.07925f
C13423 VPWR.n1606 VGND 0.0746f
C13424 VPWR.t1115 VGND 0.01009f
C13425 VPWR.n1607 VGND 0.02252f
C13426 VPWR.n1608 VGND 0.01543f
C13427 VPWR.n1609 VGND 0.05077f
C13428 VPWR.n1610 VGND 0.07925f
C13429 VPWR.n1611 VGND 0.0746f
C13430 VPWR.n1612 VGND 0.0534f
C13431 VPWR.n1613 VGND 0.04424f
C13432 VPWR.n1614 VGND 0.10954f
C13433 VPWR.n1616 VGND 0.02474f
C13434 VPWR.t1247 VGND 0.02178f
C13435 VPWR.n1618 VGND 0.04654f
C13436 VPWR.t1613 VGND 0.02407f
C13437 VPWR.n1619 VGND 0.03816f
C13438 VPWR.t1100 VGND 0.06383f
C13439 VPWR.t179 VGND 0.07496f
C13440 VPWR.n1620 VGND 0.02474f
C13441 VPWR.t1114 VGND 0.02178f
C13442 VPWR.n1622 VGND 0.04654f
C13443 VPWR.t180 VGND 0.02407f
C13444 VPWR.n1623 VGND 0.03816f
C13445 VPWR.n1625 VGND 0.088f
C13446 VPWR.t1246 VGND 0.09722f
C13447 VPWR.t1116 VGND 0.06383f
C13448 VPWR.t1612 VGND 0.07496f
C13449 VPWR.t1393 VGND 0.06383f
C13450 VPWR.t1123 VGND 0.09722f
C13451 VPWR.n1626 VGND 0.02474f
C13452 VPWR.t1288 VGND 0.02178f
C13453 VPWR.n1628 VGND 0.04654f
C13454 VPWR.t186 VGND 0.02407f
C13455 VPWR.n1629 VGND 0.03816f
C13456 VPWR.n1631 VGND 0.088f
C13457 VPWR.t185 VGND 0.07496f
C13458 VPWR.t1372 VGND 0.06383f
C13459 VPWR.t1287 VGND 0.09722f
C13460 VPWR.n1632 VGND 0.088f
C13461 VPWR.n1634 VGND 0.0512f
C13462 VPWR.n1636 VGND 0.10954f
C13463 VPWR.n1637 VGND 0.04424f
C13464 VPWR.n1638 VGND 0.0534f
C13465 VPWR.n1639 VGND 0.04424f
C13466 VPWR.n1640 VGND 0.10954f
C13467 VPWR.n1642 VGND 0.0512f
C13468 VPWR.n1644 VGND 0.088f
C13469 VPWR.t1562 VGND 0.07496f
C13470 VPWR.t1349 VGND 0.06383f
C13471 VPWR.t1385 VGND 0.09722f
C13472 VPWR.n1645 VGND 0.088f
C13473 VPWR.n1647 VGND 0.0512f
C13474 VPWR.n1649 VGND 0.0512f
C13475 VPWR.n1651 VGND 0.088f
C13476 VPWR.t514 VGND 0.07496f
C13477 VPWR.t1201 VGND 0.06383f
C13478 VPWR.t1216 VGND 0.09722f
C13479 VPWR.n1652 VGND 0.088f
C13480 VPWR.n1654 VGND 0.0512f
C13481 VPWR.n1656 VGND 0.0512f
C13482 VPWR.n1658 VGND 0.088f
C13483 VPWR.t914 VGND 0.07496f
C13484 VPWR.t1351 VGND 0.06383f
C13485 VPWR.t1346 VGND 0.09722f
C13486 VPWR.n1659 VGND 0.088f
C13487 VPWR.n1661 VGND 0.0512f
C13488 VPWR.n1663 VGND 0.10954f
C13489 VPWR.n1664 VGND -0.01517f
C13490 VPWR.n1665 VGND 0.06791f
C13491 VPWR.n1666 VGND 0.06791f
C13492 VPWR.n1667 VGND -0.01517f
C13493 VPWR.n1671 VGND 0.088f
C13494 VPWR.t1256 VGND 0.07496f
C13495 VPWR.t1249 VGND 0.06383f
C13496 VPWR.t1262 VGND 0.09722f
C13497 VPWR.n1672 VGND 0.088f
C13498 VPWR.n1675 VGND 0.05649f
C13499 VPWR.n1677 VGND -0.01517f
C13500 VPWR.n1678 VGND 0.06791f
C13501 VPWR.n1679 VGND 0.89437f
C13502 VPWR.n1680 VGND 7.44332f
C13503 VPWR.n1681 VGND 4.75452f
C13504 VPWR.n1682 VGND 0.15751f
C13505 VPWR.n1683 VGND -0.01517f
C13506 VPWR.n1684 VGND 0.10954f
C13507 VPWR.n1685 VGND 0.13384f
C13508 VPWR.n1686 VGND 0.0534f
C13509 VPWR.t1250 VGND 0.01009f
C13510 VPWR.n1687 VGND 0.02252f
C13511 VPWR.n1688 VGND 0.01543f
C13512 VPWR.n1689 VGND 0.05076f
C13513 VPWR.n1690 VGND 0.04178f
C13514 VPWR.t1421 VGND 0.01009f
C13515 VPWR.n1691 VGND 0.02252f
C13516 VPWR.n1692 VGND 0.01543f
C13517 VPWR.n1693 VGND 0.05077f
C13518 VPWR.n1694 VGND 0.07925f
C13519 VPWR.n1695 VGND 0.0746f
C13520 VPWR.n1696 VGND 0.0534f
C13521 VPWR.n1697 VGND 0.04424f
C13522 VPWR.n1698 VGND 0.0534f
C13523 VPWR.n1699 VGND 0.04424f
C13524 VPWR.n1700 VGND 0.10954f
C13525 VPWR.n1703 VGND 0.0512f
C13526 VPWR.n1705 VGND 0.088f
C13527 VPWR.t1157 VGND 0.09722f
C13528 VPWR.t1422 VGND 0.06383f
C13529 VPWR.t578 VGND 0.07496f
C13530 VPWR.n1706 VGND 0.02474f
C13531 VPWR.t1158 VGND 0.02178f
C13532 VPWR.n1708 VGND 0.04654f
C13533 VPWR.t579 VGND 0.02407f
C13534 VPWR.n1709 VGND 0.03816f
C13535 VPWR.n1711 VGND 0.088f
C13536 VPWR.t1268 VGND 0.09722f
C13537 VPWR.t1251 VGND 0.06383f
C13538 VPWR.t1388 VGND 0.10842f
C13539 VPWR.n1712 VGND 0.06192f
C13540 VPWR.n1713 VGND 0.0512f
C13541 VPWR.n1715 VGND 0.10954f
C13542 VPWR.n1716 VGND 0.0512f
C13543 VPWR.t577 VGND 0.02709f
C13544 VPWR.t1266 VGND 0.02407f
C13545 VPWR.n1718 VGND 0.07442f
C13546 VPWR.t1864 VGND 0.06383f
C13547 VPWR.t522 VGND 0.07496f
C13548 VPWR.t21 VGND 0.02709f
C13549 VPWR.t523 VGND 0.02407f
C13550 VPWR.n1719 VGND 0.07442f
C13551 VPWR.n1721 VGND 0.088f
C13552 VPWR.t576 VGND 0.09722f
C13553 VPWR.t277 VGND 0.06383f
C13554 VPWR.t1265 VGND 0.10842f
C13555 VPWR.n1722 VGND 0.06192f
C13556 VPWR.n1723 VGND 0.0512f
C13557 VPWR.n1725 VGND 0.29751f
C13558 VPWR.n1726 VGND 0.06791f
C13559 VPWR.n1727 VGND 0.06791f
C13560 VPWR.n1728 VGND 0.29751f
C13561 VPWR.n1730 VGND 0.0512f
C13562 VPWR.n1732 VGND 0.088f
C13563 VPWR.t14 VGND 0.07496f
C13564 VPWR.t1865 VGND 0.06383f
C13565 VPWR.t1476 VGND 0.09722f
C13566 VPWR.n1733 VGND 0.088f
C13567 VPWR.n1735 VGND 0.0512f
C13568 VPWR.n1737 VGND 0.0512f
C13569 VPWR.n1739 VGND 0.088f
C13570 VPWR.t1602 VGND 0.07496f
C13571 VPWR.t1860 VGND 0.06383f
C13572 VPWR.t753 VGND 0.09722f
C13573 VPWR.n1740 VGND 0.088f
C13574 VPWR.n1742 VGND 0.0512f
C13575 VPWR.n1744 VGND 0.0512f
C13576 VPWR.n1746 VGND 0.088f
C13577 VPWR.t364 VGND 0.07496f
C13578 VPWR.t89 VGND 0.06383f
C13579 VPWR.t656 VGND 0.09722f
C13580 VPWR.n1747 VGND 0.088f
C13581 VPWR.n1749 VGND 0.0512f
C13582 VPWR.n1751 VGND 0.29751f
C13583 VPWR.n1752 VGND 0.06791f
C13584 VPWR.n1753 VGND 0.06791f
C13585 VPWR.n1754 VGND 0.06791f
C13586 VPWR.n1755 VGND 0.29751f
C13587 VPWR.n1757 VGND 0.0512f
C13588 VPWR.n1759 VGND 0.088f
C13589 VPWR.t165 VGND 0.07496f
C13590 VPWR.t88 VGND 0.06383f
C13591 VPWR.t1590 VGND 0.09722f
C13592 VPWR.n1760 VGND 0.088f
C13593 VPWR.n1762 VGND 0.0512f
C13594 VPWR.n1764 VGND 0.0512f
C13595 VPWR.n1766 VGND 0.088f
C13596 VPWR.t1791 VGND 0.07496f
C13597 VPWR.t1862 VGND 0.06383f
C13598 VPWR.t1486 VGND 0.09722f
C13599 VPWR.n1767 VGND 0.088f
C13600 VPWR.n1769 VGND 0.0512f
C13601 VPWR.n1771 VGND 0.29751f
C13602 VPWR.n1772 VGND 0.06791f
C13603 VPWR.n1773 VGND 0.06791f
C13604 VPWR.n1774 VGND 0.29751f
C13605 VPWR.n1775 VGND 0.06791f
C13606 VPWR.n1776 VGND 0.06791f
C13607 VPWR.n1777 VGND 0.2969f
C13608 VPWR.n1778 VGND -0.05607f
C13609 VPWR.n1780 VGND 0.088f
C13610 VPWR.t250 VGND 0.09722f
C13611 VPWR.t1904 VGND 0.06383f
C13612 VPWR.t512 VGND 0.07496f
C13613 VPWR.t131 VGND 0.06383f
C13614 VPWR.t504 VGND 0.09722f
C13615 VPWR.n1781 VGND 0.088f
C13616 VPWR.n1783 VGND 0.0512f
C13617 VPWR.n1785 VGND 0.0512f
C13618 VPWR.n1787 VGND 0.088f
C13619 VPWR.t1508 VGND 0.09722f
C13620 VPWR.t130 VGND 0.06383f
C13621 VPWR.t818 VGND 0.07496f
C13622 VPWR.t1509 VGND 0.02709f
C13623 VPWR.t819 VGND 0.02407f
C13624 VPWR.n1788 VGND 0.07442f
C13625 VPWR.n1790 VGND 0.088f
C13626 VPWR.t1066 VGND 0.09722f
C13627 VPWR.t100 VGND 0.06383f
C13628 VPWR.t1783 VGND 0.07496f
C13629 VPWR.t99 VGND 0.06383f
C13630 VPWR.t74 VGND 0.09722f
C13631 VPWR.t429 VGND 0.02709f
C13632 VPWR.t83 VGND 0.02407f
C13633 VPWR.n1791 VGND 0.07442f
C13634 VPWR.n1793 VGND 0.088f
C13635 VPWR.t82 VGND 0.07496f
C13636 VPWR.t1901 VGND 0.06383f
C13637 VPWR.t428 VGND 0.09722f
C13638 VPWR.t1776 VGND 0.02709f
C13639 VPWR.t437 VGND 0.02407f
C13640 VPWR.n1794 VGND 0.07442f
C13641 VPWR.n1796 VGND 0.0512f
C13642 VPWR.n1798 VGND 0.088f
C13643 VPWR.t436 VGND 0.07496f
C13644 VPWR.t1902 VGND 0.06383f
C13645 VPWR.t1775 VGND 0.09722f
C13646 VPWR.n1799 VGND 0.088f
C13647 VPWR.n1801 VGND 0.0512f
C13648 VPWR.n1803 VGND 0.2969f
C13649 VPWR.n1804 VGND 0.06791f
C13650 VPWR.n1805 VGND 0.06791f
C13651 VPWR.n1806 VGND 0.2969f
C13652 VPWR.n1807 VGND 0.2969f
C13653 VPWR.n1808 VGND 0.06791f
C13654 VPWR.n1809 VGND 0.06791f
C13655 VPWR.n1810 VGND 0.06791f
C13656 VPWR.n1811 VGND 0.2969f
C13657 VPWR.n1812 VGND 0.2969f
C13658 VPWR.n1813 VGND 0.06791f
C13659 VPWR.n1814 VGND 0.06791f
C13660 VPWR.n1815 VGND 0.06791f
C13661 VPWR.n1816 VGND 0.06791f
C13662 VPWR.n1817 VGND 0.2969f
C13663 VPWR.n1820 VGND 0.0512f
C13664 VPWR.n1822 VGND 0.088f
C13665 VPWR.t717 VGND 0.09722f
C13666 VPWR.t98 VGND 0.06383f
C13667 VPWR.t891 VGND 0.07496f
C13668 VPWR.t1903 VGND 0.06383f
C13669 VPWR.t1042 VGND 0.09722f
C13670 VPWR.n1823 VGND 0.088f
C13671 VPWR.n1825 VGND 0.0512f
C13672 VPWR.n1827 VGND 0.2969f
C13673 VPWR.n1828 VGND 0.06791f
C13674 VPWR.n1829 VGND 0.06791f
C13675 VPWR.n1830 VGND 0.2969f
C13676 VPWR.n1832 VGND 0.0512f
C13677 VPWR.n1834 VGND 0.088f
C13678 VPWR.t305 VGND 0.09722f
C13679 VPWR.t129 VGND 0.06383f
C13680 VPWR.t173 VGND 0.07496f
C13681 VPWR.t1900 VGND 0.06383f
C13682 VPWR.t1820 VGND 0.09722f
C13683 VPWR.t1015 VGND 0.02709f
C13684 VPWR.t92 VGND 0.02407f
C13685 VPWR.n1835 VGND 0.07442f
C13686 VPWR.n1837 VGND 0.088f
C13687 VPWR.t91 VGND 0.07496f
C13688 VPWR.t128 VGND 0.06383f
C13689 VPWR.t1014 VGND 0.09722f
C13690 VPWR.n1838 VGND 0.088f
C13691 VPWR.n1840 VGND 0.0512f
C13692 VPWR.n1842 VGND 0.2969f
C13693 VPWR.n1843 VGND 0.06791f
C13694 VPWR.n1844 VGND 0.06791f
C13695 VPWR.n1845 VGND 0.2969f
C13696 VPWR.n1847 VGND 0.0512f
C13697 VPWR.n1849 VGND 0.088f
C13698 VPWR.t208 VGND 0.09722f
C13699 VPWR.t1899 VGND 0.06383f
C13700 VPWR.t114 VGND 0.07496f
C13701 VPWR.t835 VGND 0.06383f
C13702 VPWR.t1631 VGND 0.09722f
C13703 VPWR.n1850 VGND 0.088f
C13704 VPWR.n1852 VGND 0.0512f
C13705 VPWR.n1855 VGND 0.0512f
C13706 VPWR.n1857 VGND 0.088f
C13707 VPWR.t996 VGND 0.09722f
C13708 VPWR.t97 VGND 0.06383f
C13709 VPWR.t1419 VGND 0.10842f
C13710 VPWR.n1858 VGND 0.06192f
C13711 VPWR.n1859 VGND 0.0512f
C13712 VPWR.n1861 VGND 0.2969f
C13713 VPWR.n1862 VGND 0.15751f
C13714 VPWR.n1863 VGND 0.06791f
C13715 VPWR.n1864 VGND 0.06791f
C13716 VPWR.n1865 VGND 0.06791f
C13717 VPWR.n1866 VGND 0.2969f
C13718 VPWR.n1867 VGND 0.2969f
C13719 VPWR.n1868 VGND 0.06791f
C13720 VPWR.n1869 VGND 0.06791f
C13721 VPWR.n1870 VGND 0.2969f
C13722 VPWR.n1872 VGND 0.0512f
C13723 VPWR.n1874 VGND 0.088f
C13724 VPWR.t22 VGND 0.07496f
C13725 VPWR.t199 VGND 0.06383f
C13726 VPWR.t1464 VGND 0.09722f
C13727 VPWR.n1875 VGND 0.088f
C13728 VPWR.n1877 VGND 0.0512f
C13729 VPWR.n1879 VGND 0.0512f
C13730 VPWR.n1881 VGND 0.088f
C13731 VPWR.t1610 VGND 0.07496f
C13732 VPWR.t1922 VGND 0.06383f
C13733 VPWR.t220 VGND 0.09722f
C13734 VPWR.n1882 VGND 0.088f
C13735 VPWR.n1884 VGND 0.0512f
C13736 VPWR.n1886 VGND 0.0512f
C13737 VPWR.n1888 VGND 0.088f
C13738 VPWR.t354 VGND 0.07496f
C13739 VPWR.t1914 VGND 0.06383f
C13740 VPWR.t666 VGND 0.09722f
C13741 VPWR.n1889 VGND 0.088f
C13742 VPWR.n1891 VGND 0.0512f
C13743 VPWR.n1893 VGND 0.2969f
C13744 VPWR.n1894 VGND 0.06791f
C13745 VPWR.n1895 VGND 0.06791f
C13746 VPWR.n1896 VGND 0.06791f
C13747 VPWR.n1897 VGND 0.2969f
C13748 VPWR.n1899 VGND 0.0512f
C13749 VPWR.n1901 VGND 0.088f
C13750 VPWR.t1853 VGND 0.07496f
C13751 VPWR.t1913 VGND 0.06383f
C13752 VPWR.t924 VGND 0.09722f
C13753 VPWR.n1902 VGND 0.088f
C13754 VPWR.n1904 VGND 0.0512f
C13755 VPWR.n1906 VGND 0.0512f
C13756 VPWR.n1908 VGND 0.088f
C13757 VPWR.t1785 VGND 0.07496f
C13758 VPWR.t196 VGND 0.06383f
C13759 VPWR.t1496 VGND 0.09722f
C13760 VPWR.n1909 VGND 0.088f
C13761 VPWR.n1911 VGND 0.0512f
C13762 VPWR.n1913 VGND 0.2969f
C13763 VPWR.n1914 VGND 0.06791f
C13764 VPWR.n1915 VGND 0.06791f
C13765 VPWR.n1916 VGND 0.82079f
C13766 VPWR.n1917 VGND 0.82079f
C13767 VPWR.n1918 VGND 0.06791f
C13768 VPWR.n1919 VGND 0.06791f
C13769 VPWR.n1920 VGND 0.06791f
C13770 VPWR.n1921 VGND 0.2969f
C13771 VPWR.t598 VGND 0.02709f
C13772 VPWR.t791 VGND 0.02407f
C13773 VPWR.n1922 VGND 0.07442f
C13774 VPWR.t597 VGND 0.118f
C13775 VPWR.t1622 VGND 0.06383f
C13776 VPWR.t790 VGND 0.07496f
C13777 VPWR.t1617 VGND 0.06383f
C13778 VPWR.t700 VGND 0.09722f
C13779 VPWR.n1923 VGND 0.088f
C13780 VPWR.n1925 VGND -0.05607f
C13781 VPWR.n1926 VGND 0.2969f
C13782 VPWR.n1927 VGND 0.06791f
C13783 VPWR.n1928 VGND 0.06791f
C13784 VPWR.n1929 VGND 0.2969f
C13785 VPWR.n1931 VGND 0.0512f
C13786 VPWR.n1933 VGND 0.088f
C13787 VPWR.t937 VGND 0.09722f
C13788 VPWR.t443 VGND 0.06383f
C13789 VPWR.t1530 VGND 0.07496f
C13790 VPWR.t938 VGND 0.02709f
C13791 VPWR.t1531 VGND 0.02407f
C13792 VPWR.n1934 VGND 0.07442f
C13793 VPWR.n1936 VGND 0.088f
C13794 VPWR.t1494 VGND 0.09722f
C13795 VPWR.t442 VGND 0.06383f
C13796 VPWR.t1787 VGND 0.07496f
C13797 VPWR.t447 VGND 0.06383f
C13798 VPWR.t1849 VGND 0.09722f
C13799 VPWR.t1583 VGND 0.02709f
C13800 VPWR.t1856 VGND 0.02407f
C13801 VPWR.n1937 VGND 0.07442f
C13802 VPWR.n1939 VGND 0.088f
C13803 VPWR.t1855 VGND 0.07496f
C13804 VPWR.t448 VGND 0.06383f
C13805 VPWR.t1582 VGND 0.09722f
C13806 VPWR.t817 VGND 0.02709f
C13807 VPWR.t1589 VGND 0.02407f
C13808 VPWR.n1940 VGND 0.07442f
C13809 VPWR.n1941 VGND 0.0512f
C13810 VPWR.n1943 VGND 0.088f
C13811 VPWR.t1588 VGND 0.07496f
C13812 VPWR.t1621 VGND 0.06383f
C13813 VPWR.t816 VGND 0.09722f
C13814 VPWR.n1944 VGND 0.088f
C13815 VPWR.n1946 VGND 0.0512f
C13816 VPWR.n1948 VGND 0.2969f
C13817 VPWR.n1949 VGND 0.06791f
C13818 VPWR.n1950 VGND 0.06791f
C13819 VPWR.n1951 VGND 0.2969f
C13820 VPWR.n1952 VGND 0.2969f
C13821 VPWR.n1953 VGND 0.06791f
C13822 VPWR.n1954 VGND 0.06791f
C13823 VPWR.n1955 VGND 0.06791f
C13824 VPWR.n1956 VGND 0.06791f
C13825 VPWR.n1957 VGND 0.06791f
C13826 VPWR.n1958 VGND 0.06791f
C13827 VPWR.n1959 VGND 0.2969f
C13828 VPWR.n1961 VGND 0.0512f
C13829 VPWR.n1963 VGND 0.088f
C13830 VPWR.t467 VGND 0.09722f
C13831 VPWR.t874 VGND 0.06383f
C13832 VPWR.t725 VGND 0.07496f
C13833 VPWR.t873 VGND 0.06383f
C13834 VPWR.t112 VGND 0.09722f
C13835 VPWR.n1964 VGND 0.088f
C13836 VPWR.n1966 VGND 0.0512f
C13837 VPWR.n1969 VGND 0.0512f
C13838 VPWR.n1971 VGND 0.088f
C13839 VPWR.t566 VGND 0.09722f
C13840 VPWR.t691 VGND 0.06383f
C13841 VPWR.t273 VGND 0.07496f
C13842 VPWR.t878 VGND 0.06383f
C13843 VPWR.t267 VGND 0.09722f
C13844 VPWR.n1972 VGND 0.088f
C13845 VPWR.n1974 VGND 0.0512f
C13846 VPWR.n1976 VGND 0.06791f
C13847 VPWR.n1977 VGND 0.06791f
C13848 VPWR.n1978 VGND 0.06791f
C13849 VPWR.n1979 VGND 0.2969f
C13850 VPWR.n1980 VGND 0.2969f
C13851 VPWR.n1981 VGND 0.06791f
C13852 VPWR.n1982 VGND 0.06791f
C13853 VPWR.n1983 VGND 0.2969f
C13854 VPWR.n1985 VGND 0.0512f
C13855 VPWR.n1987 VGND 0.088f
C13856 VPWR.t1024 VGND 0.09722f
C13857 VPWR.t877 VGND 0.06383f
C13858 VPWR.t1546 VGND 0.07496f
C13859 VPWR.t1025 VGND 0.02709f
C13860 VPWR.t1547 VGND 0.02407f
C13861 VPWR.n1988 VGND 0.07442f
C13862 VPWR.n1990 VGND 0.088f
C13863 VPWR.t910 VGND 0.09722f
C13864 VPWR.t688 VGND 0.06383f
C13865 VPWR.t216 VGND 0.07496f
C13866 VPWR.t1907 VGND 0.09722f
C13867 VPWR.t1055 VGND 0.02709f
C13868 VPWR.t1817 VGND 0.02407f
C13869 VPWR.n1991 VGND 0.07442f
C13870 VPWR.t1908 VGND 0.02709f
C13871 VPWR.t1005 VGND 0.02407f
C13872 VPWR.n1992 VGND 0.07442f
C13873 VPWR.t686 VGND 0.06383f
C13874 VPWR.t1004 VGND 0.07496f
C13875 VPWR.t527 VGND 0.02709f
C13876 VPWR.t1119 VGND 0.02407f
C13877 VPWR.n1993 VGND 0.07442f
C13878 VPWR.n1994 VGND 0.0512f
C13879 VPWR.n1995 VGND 0.06192f
C13880 VPWR.t1118 VGND 0.10842f
C13881 VPWR.t872 VGND 0.06383f
C13882 VPWR.t526 VGND 0.09722f
C13883 VPWR.n1996 VGND 0.088f
C13884 VPWR.n1998 VGND 0.0512f
C13885 VPWR.n2000 VGND 0.0512f
C13886 VPWR.n2002 VGND 0.088f
C13887 VPWR.t1816 VGND 0.07496f
C13888 VPWR.t687 VGND 0.06383f
C13889 VPWR.t1054 VGND 0.09722f
C13890 VPWR.n2003 VGND 0.088f
C13891 VPWR.n2005 VGND 0.0512f
C13892 VPWR.n2007 VGND 0.2969f
C13893 VPWR.n2008 VGND 0.06791f
C13894 VPWR.n2009 VGND 0.06791f
C13895 VPWR.n2010 VGND 0.06791f
C13896 VPWR.n2011 VGND 0.06791f
C13897 VPWR.n2012 VGND 0.2969f
C13898 VPWR.n2013 VGND 0.2969f
C13899 VPWR.n2014 VGND 0.06791f
C13900 VPWR.n2015 VGND 0.15751f
C13901 VPWR.n2016 VGND 0.82597f
C13902 VPWR.n2017 VGND 0.82597f
C13903 VPWR.n2018 VGND 0.15751f
C13904 VPWR.n2019 VGND 0.2969f
C13905 VPWR.n2020 VGND 0.06791f
C13906 VPWR.n2021 VGND 0.15751f
C13907 VPWR.n2022 VGND 0.2969f
C13908 VPWR.n2024 VGND 0.0512f
C13909 VPWR.n2025 VGND 0.06192f
C13910 VPWR.t1298 VGND 0.10842f
C13911 VPWR.t1618 VGND 0.06383f
C13912 VPWR.t1718 VGND 0.09722f
C13913 VPWR.n2026 VGND 0.088f
C13914 VPWR.n2028 VGND 0.0512f
C13915 VPWR.n2030 VGND 0.2969f
C13916 VPWR.n2031 VGND 0.06791f
C13917 VPWR.n2032 VGND 0.06791f
C13918 VPWR.n2033 VGND 0.2969f
C13919 VPWR.n2035 VGND 0.0512f
C13920 VPWR.n2037 VGND 0.088f
C13921 VPWR.t1046 VGND 0.07496f
C13922 VPWR.t446 VGND 0.06383f
C13923 VPWR.t1604 VGND 0.09722f
C13924 VPWR.n2038 VGND 0.088f
C13925 VPWR.n2040 VGND 0.0512f
C13926 VPWR.n2042 VGND 0.0512f
C13927 VPWR.n2044 VGND 0.088f
C13928 VPWR.t751 VGND 0.07496f
C13929 VPWR.t441 VGND 0.06383f
C13930 VPWR.t1893 VGND 0.09722f
C13931 VPWR.n2045 VGND 0.088f
C13932 VPWR.n2047 VGND 0.0512f
C13933 VPWR.n2049 VGND 0.2969f
C13934 VPWR.n2050 VGND 0.06791f
C13935 VPWR.n2051 VGND 0.06791f
C13936 VPWR.n2052 VGND 0.2969f
C13937 VPWR.n2054 VGND 0.0512f
C13938 VPWR.n2056 VGND 0.088f
C13939 VPWR.t654 VGND 0.07496f
C13940 VPWR.t1620 VGND 0.06383f
C13941 VPWR.t1839 VGND 0.09722f
C13942 VPWR.n2057 VGND 0.088f
C13943 VPWR.n2059 VGND 0.0512f
C13944 VPWR.n2061 VGND 0.2969f
C13945 VPWR.n2062 VGND 0.06791f
C13946 VPWR.n2063 VGND 0.06791f
C13947 VPWR.n2064 VGND 0.2969f
C13948 VPWR.n2065 VGND 0.0512f
C13949 VPWR.t1700 VGND 0.02709f
C13950 VPWR.t1805 VGND 0.02407f
C13951 VPWR.n2067 VGND 0.07442f
C13952 VPWR.t715 VGND 0.07496f
C13953 VPWR.t1535 VGND 0.02709f
C13954 VPWR.t716 VGND 0.02407f
C13955 VPWR.n2068 VGND 0.07442f
C13956 VPWR.t775 VGND 0.02709f
C13957 VPWR.t1511 VGND 0.02407f
C13958 VPWR.n2069 VGND 0.07442f
C13959 VPWR.t776 VGND 0.07496f
C13960 VPWR.t1688 VGND 0.02709f
C13961 VPWR.t777 VGND 0.02407f
C13962 VPWR.n2070 VGND 0.07442f
C13963 VPWR.t618 VGND 0.02709f
C13964 VPWR.t247 VGND 0.02407f
C13965 VPWR.n2071 VGND 0.07442f
C13966 VPWR.t617 VGND 0.118f
C13967 VPWR.t901 VGND 0.06383f
C13968 VPWR.t246 VGND 0.07496f
C13969 VPWR.t1037 VGND 0.06383f
C13970 VPWR.t1687 VGND 0.09722f
C13971 VPWR.n2072 VGND 0.088f
C13972 VPWR.n2074 VGND -0.05607f
C13973 VPWR.n2076 VGND 0.0512f
C13974 VPWR.n2078 VGND 0.088f
C13975 VPWR.t774 VGND 0.09722f
C13976 VPWR.t1661 VGND 0.06383f
C13977 VPWR.t1510 VGND 0.07496f
C13978 VPWR.t1660 VGND 0.06383f
C13979 VPWR.t1534 VGND 0.09722f
C13980 VPWR.n2079 VGND 0.088f
C13981 VPWR.n2081 VGND 0.0512f
C13982 VPWR.n2084 VGND 0.0512f
C13983 VPWR.n2086 VGND 0.088f
C13984 VPWR.t734 VGND 0.09722f
C13985 VPWR.t900 VGND 0.06383f
C13986 VPWR.t1701 VGND 0.07496f
C13987 VPWR.t735 VGND 0.02709f
C13988 VPWR.t1702 VGND 0.02407f
C13989 VPWR.n2087 VGND 0.07442f
C13990 VPWR.n2089 VGND 0.088f
C13991 VPWR.t1699 VGND 0.09722f
C13992 VPWR.t1035 VGND 0.06383f
C13993 VPWR.t1804 VGND 0.07496f
C13994 VPWR.t461 VGND 0.09722f
C13995 VPWR.t1803 VGND 0.02709f
C13996 VPWR.t464 VGND 0.02407f
C13997 VPWR.n2090 VGND 0.07442f
C13998 VPWR.t462 VGND 0.02709f
C13999 VPWR.t869 VGND 0.02407f
C14000 VPWR.n2092 VGND 0.07442f
C14001 VPWR.t899 VGND 0.06383f
C14002 VPWR.t868 VGND 0.07496f
C14003 VPWR.t126 VGND 0.09722f
C14004 VPWR.t651 VGND 0.02709f
C14005 VPWR.t420 VGND 0.02407f
C14006 VPWR.n2093 VGND 0.07442f
C14007 VPWR.t127 VGND 0.02709f
C14008 VPWR.t264 VGND 0.02407f
C14009 VPWR.n2095 VGND 0.07442f
C14010 VPWR.t1036 VGND 0.06383f
C14011 VPWR.t263 VGND 0.07496f
C14012 VPWR.t1658 VGND 0.06383f
C14013 VPWR.t765 VGND 0.09722f
C14014 VPWR.t369 VGND 0.02709f
C14015 VPWR.t768 VGND 0.02407f
C14016 VPWR.n2096 VGND 0.07442f
C14017 VPWR.n2097 VGND 0.0512f
C14018 VPWR.n2099 VGND 0.088f
C14019 VPWR.t767 VGND 0.07496f
C14020 VPWR.t1659 VGND 0.06383f
C14021 VPWR.t368 VGND 0.09722f
C14022 VPWR.n2100 VGND 0.088f
C14023 VPWR.n2102 VGND 0.0512f
C14024 VPWR.n2104 VGND 0.0512f
C14025 VPWR.n2106 VGND 0.088f
C14026 VPWR.t419 VGND 0.07496f
C14027 VPWR.t898 VGND 0.06383f
C14028 VPWR.t650 VGND 0.09722f
C14029 VPWR.n2107 VGND 0.088f
C14030 VPWR.n2109 VGND 0.0512f
C14031 VPWR.n2111 VGND 0.0512f
C14032 VPWR.n2113 VGND 0.088f
C14033 VPWR.t463 VGND 0.07496f
C14034 VPWR.t1034 VGND 0.06383f
C14035 VPWR.t1802 VGND 0.09722f
C14036 VPWR.n2114 VGND 0.088f
C14037 VPWR.n2116 VGND 0.0512f
C14038 VPWR.n2118 VGND 0.2969f
C14039 VPWR.n2119 VGND 0.06791f
C14040 VPWR.n2120 VGND 0.06791f
C14041 VPWR.n2121 VGND 0.06791f
C14042 VPWR.n2122 VGND 0.06791f
C14043 VPWR.n2123 VGND 0.06791f
C14044 VPWR.n2124 VGND 0.82079f
C14045 VPWR.n2125 VGND 0.82079f
C14046 VPWR.n2126 VGND 0.82079f
C14047 VPWR.n2127 VGND 0.06791f
C14048 VPWR.n2128 VGND 0.06791f
C14049 VPWR.n2129 VGND 0.06791f
C14050 VPWR.n2130 VGND 0.06791f
C14051 VPWR.n2131 VGND 0.2969f
C14052 VPWR.n2132 VGND 0.2969f
C14053 VPWR.n2133 VGND 0.06791f
C14054 VPWR.n2134 VGND 0.06791f
C14055 VPWR.n2135 VGND 0.2969f
C14056 VPWR.n2137 VGND 0.0512f
C14057 VPWR.n2139 VGND 0.088f
C14058 VPWR.t1627 VGND 0.09722f
C14059 VPWR.t536 VGND 0.06383f
C14060 VPWR.t1518 VGND 0.07496f
C14061 VPWR.t880 VGND 0.06383f
C14062 VPWR.t730 VGND 0.09722f
C14063 VPWR.t1541 VGND 0.02709f
C14064 VPWR.t710 VGND 0.02407f
C14065 VPWR.n2140 VGND 0.07442f
C14066 VPWR.n2142 VGND 0.088f
C14067 VPWR.t709 VGND 0.07496f
C14068 VPWR.t743 VGND 0.06383f
C14069 VPWR.t1540 VGND 0.09722f
C14070 VPWR.n2143 VGND 0.088f
C14071 VPWR.n2145 VGND 0.0512f
C14072 VPWR.n2147 VGND 0.2969f
C14073 VPWR.n2148 VGND 0.06791f
C14074 VPWR.n2149 VGND 0.06791f
C14075 VPWR.n2150 VGND 0.06791f
C14076 VPWR.n2151 VGND 0.2969f
C14077 VPWR.n2154 VGND 0.0512f
C14078 VPWR.n2156 VGND 0.088f
C14079 VPWR.t159 VGND 0.09722f
C14080 VPWR.t32 VGND 0.06383f
C14081 VPWR.t171 VGND 0.07496f
C14082 VPWR.t31 VGND 0.06383f
C14083 VPWR.t167 VGND 0.09722f
C14084 VPWR.n2157 VGND 0.088f
C14085 VPWR.n2159 VGND 0.0512f
C14086 VPWR.n2161 VGND 0.2969f
C14087 VPWR.n2162 VGND 0.06791f
C14088 VPWR.n2163 VGND 0.06791f
C14089 VPWR.n2164 VGND 0.2969f
C14090 VPWR.n2166 VGND 0.0512f
C14091 VPWR.n2168 VGND 0.088f
C14092 VPWR.t479 VGND 0.09722f
C14093 VPWR.t879 VGND 0.06383f
C14094 VPWR.t2 VGND 0.07496f
C14095 VPWR.t1648 VGND 0.06383f
C14096 VPWR.t516 VGND 0.09722f
C14097 VPWR.n2169 VGND 0.088f
C14098 VPWR.n2171 VGND 0.0512f
C14099 VPWR.n2173 VGND 0.2969f
C14100 VPWR.n2174 VGND 0.06791f
C14101 VPWR.n2175 VGND 0.06791f
C14102 VPWR.n2176 VGND 0.2969f
C14103 VPWR.n2178 VGND 0.0512f
C14104 VPWR.n2180 VGND 0.088f
C14105 VPWR.t662 VGND 0.09722f
C14106 VPWR.t33 VGND 0.06383f
C14107 VPWR.t366 VGND 0.07496f
C14108 VPWR.t663 VGND 0.02709f
C14109 VPWR.t367 VGND 0.02407f
C14110 VPWR.n2181 VGND 0.07442f
C14111 VPWR.n2183 VGND 0.088f
C14112 VPWR.t360 VGND 0.09722f
C14113 VPWR.t742 VGND 0.06383f
C14114 VPWR.t1579 VGND 0.07496f
C14115 VPWR.t1598 VGND 0.09722f
C14116 VPWR.t1576 VGND 0.02709f
C14117 VPWR.t1811 VGND 0.02407f
C14118 VPWR.n2184 VGND 0.07442f
C14119 VPWR.t1599 VGND 0.02709f
C14120 VPWR.t1059 VGND 0.02407f
C14121 VPWR.n2185 VGND 0.07442f
C14122 VPWR.t30 VGND 0.06383f
C14123 VPWR.t1058 VGND 0.07496f
C14124 VPWR.t537 VGND 0.06383f
C14125 VPWR.t10 VGND 0.09722f
C14126 VPWR.t188 VGND 0.02709f
C14127 VPWR.t17 VGND 0.02407f
C14128 VPWR.n2186 VGND 0.07442f
C14129 VPWR.n2188 VGND 0.088f
C14130 VPWR.t16 VGND 0.07496f
C14131 VPWR.t538 VGND 0.06383f
C14132 VPWR.t187 VGND 0.09722f
C14133 VPWR.n2189 VGND 0.088f
C14134 VPWR.n2191 VGND 0.0512f
C14135 VPWR.n2193 VGND 0.0512f
C14136 VPWR.n2195 VGND 0.088f
C14137 VPWR.t1810 VGND 0.07496f
C14138 VPWR.t741 VGND 0.06383f
C14139 VPWR.t1575 VGND 0.09722f
C14140 VPWR.n2196 VGND 0.088f
C14141 VPWR.n2198 VGND 0.0512f
C14142 VPWR.n2200 VGND 0.2969f
C14143 VPWR.n2201 VGND 0.06791f
C14144 VPWR.n2202 VGND 0.06791f
C14145 VPWR.n2203 VGND 0.06791f
C14146 VPWR.n2204 VGND 0.2969f
C14147 VPWR.n2205 VGND 0.2969f
C14148 VPWR.n2206 VGND 0.06791f
C14149 VPWR.n2207 VGND 0.06791f
C14150 VPWR.n2208 VGND 0.06791f
C14151 VPWR.n2209 VGND 0.06791f
C14152 VPWR.n2210 VGND 0.2969f
C14153 VPWR.n2212 VGND 0.0512f
C14154 VPWR.n2214 VGND 0.088f
C14155 VPWR.t1812 VGND 0.09722f
C14156 VPWR.t1033 VGND 0.06383f
C14157 VPWR.t204 VGND 0.07496f
C14158 VPWR.t1663 VGND 0.06383f
C14159 VPWR.t191 VGND 0.09722f
C14160 VPWR.n2215 VGND 0.088f
C14161 VPWR.n2217 VGND 0.0512f
C14162 VPWR.n2220 VGND 0.0512f
C14163 VPWR.n2222 VGND 0.088f
C14164 VPWR.t18 VGND 0.09722f
C14165 VPWR.t1662 VGND 0.06383f
C14166 VPWR.t534 VGND 0.07496f
C14167 VPWR.t19 VGND 0.02709f
C14168 VPWR.t535 VGND 0.02407f
C14169 VPWR.n2223 VGND 0.07442f
C14170 VPWR.n2225 VGND 0.088f
C14171 VPWR.t584 VGND 0.09722f
C14172 VPWR.t897 VGND 0.06383f
C14173 VPWR.t1193 VGND 0.10842f
C14174 VPWR.n2226 VGND 0.06192f
C14175 VPWR.n2227 VGND 0.0512f
C14176 VPWR.n2229 VGND 0.2969f
C14177 VPWR.n2230 VGND 0.06791f
C14178 VPWR.n2231 VGND 0.15751f
C14179 VPWR.n2232 VGND 0.82597f
C14180 VPWR.n2233 VGND 0.82597f
C14181 VPWR.n2234 VGND 0.15751f
C14182 VPWR.n2235 VGND 0.2969f
C14183 VPWR.n2237 VGND 0.0512f
C14184 VPWR.n2238 VGND 0.06192f
C14185 VPWR.t1233 VGND 0.10842f
C14186 VPWR.t1647 VGND 0.06383f
C14187 VPWR.t580 VGND 0.09722f
C14188 VPWR.n2239 VGND 0.088f
C14189 VPWR.n2241 VGND 0.0512f
C14190 VPWR.n2243 VGND 0.2969f
C14191 VPWR.n2244 VGND 0.06791f
C14192 VPWR.n2245 VGND 0.06791f
C14193 VPWR.n2246 VGND 0.2969f
C14194 VPWR.n2247 VGND 0.2969f
C14195 VPWR.n2248 VGND 0.06791f
C14196 VPWR.n2249 VGND 0.06791f
C14197 VPWR.n2250 VGND 0.15751f
C14198 VPWR.n2251 VGND 0.06791f
C14199 VPWR.n2252 VGND 0.2969f
C14200 VPWR.t1906 VGND 0.02709f
C14201 VPWR.t1001 VGND 0.02407f
C14202 VPWR.n2254 VGND 0.07442f
C14203 VPWR.t497 VGND 0.06383f
C14204 VPWR.t1000 VGND 0.07496f
C14205 VPWR.t525 VGND 0.02709f
C14206 VPWR.t1127 VGND 0.02407f
C14207 VPWR.n2255 VGND 0.07442f
C14208 VPWR.n2257 VGND 0.0512f
C14209 VPWR.n2258 VGND 0.06192f
C14210 VPWR.t1126 VGND 0.10842f
C14211 VPWR.t562 VGND 0.06383f
C14212 VPWR.t524 VGND 0.09722f
C14213 VPWR.n2259 VGND 0.088f
C14214 VPWR.n2261 VGND 0.0512f
C14215 VPWR.n2263 VGND 0.0512f
C14216 VPWR.n2265 VGND 0.088f
C14217 VPWR.t1911 VGND 0.07496f
C14218 VPWR.t291 VGND 0.06383f
C14219 VPWR.t1052 VGND 0.09722f
C14220 VPWR.n2266 VGND 0.088f
C14221 VPWR.n2268 VGND 0.0512f
C14222 VPWR.n2270 VGND 0.2969f
C14223 VPWR.n2271 VGND 0.06791f
C14224 VPWR.n2272 VGND 0.06791f
C14225 VPWR.n2273 VGND 0.06791f
C14226 VPWR.n2274 VGND 0.06791f
C14227 VPWR.n2275 VGND 0.06791f
C14228 VPWR.n2276 VGND 0.06791f
C14229 VPWR.n2277 VGND 0.06791f
C14230 VPWR.n2278 VGND 0.06791f
C14231 VPWR.n2279 VGND 0.2969f
C14232 VPWR.n2280 VGND 0.2969f
C14233 VPWR.n2281 VGND 0.06791f
C14234 VPWR.n2282 VGND 0.06791f
C14235 VPWR.n2283 VGND 0.2969f
C14236 VPWR.n2285 VGND 0.0512f
C14237 VPWR.n2287 VGND 0.088f
C14238 VPWR.t438 VGND 0.07496f
C14239 VPWR.t299 VGND 0.06383f
C14240 VPWR.t1779 VGND 0.09722f
C14241 VPWR.n2288 VGND 0.088f
C14242 VPWR.n2290 VGND 0.0512f
C14243 VPWR.n2292 VGND 0.2969f
C14244 VPWR.n2293 VGND 0.06791f
C14245 VPWR.n2294 VGND 0.06791f
C14246 VPWR.n2295 VGND 0.2969f
C14247 VPWR.n2296 VGND 0.2969f
C14248 VPWR.n2297 VGND 0.06791f
C14249 VPWR.n2298 VGND 0.06791f
C14250 VPWR.n2299 VGND 0.06791f
C14251 VPWR.n2300 VGND 0.06791f
C14252 VPWR.n2301 VGND 0.06791f
C14253 VPWR.n2302 VGND 0.06791f
C14254 VPWR.n2303 VGND 0.2969f
C14255 VPWR.n2304 VGND 0.2969f
C14256 VPWR.n2305 VGND 0.06791f
C14257 VPWR.n2306 VGND 0.06791f
C14258 VPWR.n2307 VGND 0.2969f
C14259 VPWR.n2309 VGND 0.0512f
C14260 VPWR.n2311 VGND 0.088f
C14261 VPWR.t887 VGND 0.09722f
C14262 VPWR.t300 VGND 0.06383f
C14263 VPWR.t1558 VGND 0.07496f
C14264 VPWR.t888 VGND 0.02709f
C14265 VPWR.t1559 VGND 0.02407f
C14266 VPWR.n2312 VGND 0.07442f
C14267 VPWR.n2314 VGND 0.088f
C14268 VPWR.t307 VGND 0.09722f
C14269 VPWR.t397 VGND 0.06383f
C14270 VPWR.t175 VGND 0.07496f
C14271 VPWR.t1822 VGND 0.09722f
C14272 VPWR.t1019 VGND 0.02709f
C14273 VPWR.t94 VGND 0.02407f
C14274 VPWR.n2315 VGND 0.07442f
C14275 VPWR.t1823 VGND 0.02709f
C14276 VPWR.t1479 VGND 0.02407f
C14277 VPWR.n2317 VGND 0.07442f
C14278 VPWR.t297 VGND 0.06383f
C14279 VPWR.t1478 VGND 0.07496f
C14280 VPWR.t295 VGND 0.06383f
C14281 VPWR.t1633 VGND 0.09722f
C14282 VPWR.t211 VGND 0.02709f
C14283 VPWR.t117 VGND 0.02407f
C14284 VPWR.n2318 VGND 0.07442f
C14285 VPWR.n2320 VGND 0.088f
C14286 VPWR.t116 VGND 0.07496f
C14287 VPWR.t296 VGND 0.06383f
C14288 VPWR.t210 VGND 0.09722f
C14289 VPWR.n2321 VGND 0.088f
C14290 VPWR.n2323 VGND 0.0512f
C14291 VPWR.n2325 VGND 0.0512f
C14292 VPWR.n2327 VGND 0.088f
C14293 VPWR.t93 VGND 0.07496f
C14294 VPWR.t319 VGND 0.06383f
C14295 VPWR.t1018 VGND 0.09722f
C14296 VPWR.n2328 VGND 0.088f
C14297 VPWR.n2330 VGND 0.0512f
C14298 VPWR.n2332 VGND 0.2969f
C14299 VPWR.n2333 VGND 0.06791f
C14300 VPWR.n2334 VGND 0.06791f
C14301 VPWR.n2335 VGND 0.2969f
C14302 VPWR.n2336 VGND 0.2969f
C14303 VPWR.n2337 VGND 0.06791f
C14304 VPWR.n2338 VGND 0.06791f
C14305 VPWR.n2339 VGND 0.06791f
C14306 VPWR.n2340 VGND 0.2969f
C14307 VPWR.n2341 VGND 0.2969f
C14308 VPWR.n2342 VGND 0.06791f
C14309 VPWR.n2343 VGND 0.06791f
C14310 VPWR.n2344 VGND 0.06791f
C14311 VPWR.n2345 VGND 0.06791f
C14312 VPWR.n2346 VGND 0.06791f
C14313 VPWR.n2347 VGND 0.2969f
C14314 VPWR.n2350 VGND 0.0512f
C14315 VPWR.n2352 VGND 0.088f
C14316 VPWR.t998 VGND 0.09722f
C14317 VPWR.t314 VGND 0.06383f
C14318 VPWR.t1409 VGND 0.10842f
C14319 VPWR.n2353 VGND 0.06192f
C14320 VPWR.n2354 VGND 0.0512f
C14321 VPWR.n2356 VGND 0.2969f
C14322 VPWR.n2357 VGND 0.15751f
C14323 VPWR.n2358 VGND 0.82597f
C14324 VPWR.n2359 VGND 0.82597f
C14325 VPWR.n2360 VGND 0.15751f
C14326 VPWR.n2361 VGND 0.06791f
C14327 VPWR.n2362 VGND 0.2969f
C14328 VPWR.n2364 VGND 0.0512f
C14329 VPWR.n2366 VGND 0.088f
C14330 VPWR.t520 VGND 0.07496f
C14331 VPWR.t329 VGND 0.06383f
C14332 VPWR.t1707 VGND 0.09722f
C14333 VPWR.n2367 VGND 0.088f
C14334 VPWR.n2369 VGND 0.0512f
C14335 VPWR.n2371 VGND 0.2969f
C14336 VPWR.n2372 VGND 0.06791f
C14337 VPWR.n2373 VGND 0.06791f
C14338 VPWR.n2374 VGND 0.2969f
C14339 VPWR.n2376 VGND 0.0512f
C14340 VPWR.n2378 VGND 0.088f
C14341 VPWR.t1596 VGND 0.07496f
C14342 VPWR.t325 VGND 0.06383f
C14343 VPWR.t747 VGND 0.09722f
C14344 VPWR.n2379 VGND 0.088f
C14345 VPWR.n2381 VGND 0.0512f
C14346 VPWR.n2383 VGND 0.0512f
C14347 VPWR.n2385 VGND 0.088f
C14348 VPWR.t358 VGND 0.07496f
C14349 VPWR.t1651 VGND 0.06383f
C14350 VPWR.t670 VGND 0.09722f
C14351 VPWR.n2386 VGND 0.088f
C14352 VPWR.n2388 VGND 0.0512f
C14353 VPWR.n2390 VGND 0.0512f
C14354 VPWR.n2392 VGND 0.088f
C14355 VPWR.t106 VGND 0.07496f
C14356 VPWR.t1655 VGND 0.06383f
C14357 VPWR.t1841 VGND 0.09722f
C14358 VPWR.n2393 VGND 0.088f
C14359 VPWR.n2395 VGND 0.0512f
C14360 VPWR.n2397 VGND 0.0512f
C14361 VPWR.n2399 VGND 0.088f
C14362 VPWR.t163 VGND 0.07496f
C14363 VPWR.t1650 VGND 0.06383f
C14364 VPWR.t1584 VGND 0.09722f
C14365 VPWR.n2400 VGND 0.088f
C14366 VPWR.n2402 VGND 0.0512f
C14367 VPWR.n2404 VGND 0.0512f
C14368 VPWR.n2406 VGND 0.088f
C14369 VPWR.t1789 VGND 0.07496f
C14370 VPWR.t327 VGND 0.06383f
C14371 VPWR.t1492 VGND 0.09722f
C14372 VPWR.n2407 VGND 0.088f
C14373 VPWR.n2409 VGND 0.0512f
C14374 VPWR.n2411 VGND 0.2969f
C14375 VPWR.n2412 VGND 0.06791f
C14376 VPWR.n2413 VGND 0.06791f
C14377 VPWR.n2414 VGND 0.82079f
C14378 VPWR.n2415 VGND 0.06791f
C14379 VPWR.n2416 VGND 0.82079f
C14380 VPWR.n2417 VGND 0.82079f
C14381 VPWR.n2418 VGND 0.06791f
C14382 VPWR.n2419 VGND 0.06791f
C14383 VPWR.n2420 VGND 0.06791f
C14384 VPWR.n2421 VGND 0.2969f
C14385 VPWR.n2422 VGND -0.05607f
C14386 VPWR.n2424 VGND 0.0512f
C14387 VPWR.n2426 VGND 0.088f
C14388 VPWR.t254 VGND 0.09722f
C14389 VPWR.t848 VGND 0.06383f
C14390 VPWR.t1490 VGND 0.07496f
C14391 VPWR.t847 VGND 0.06383f
C14392 VPWR.t1514 VGND 0.09722f
C14393 VPWR.n2427 VGND 0.088f
C14394 VPWR.n2429 VGND 0.0512f
C14395 VPWR.n2431 VGND 0.0512f
C14396 VPWR.n2433 VGND 0.088f
C14397 VPWR.t1062 VGND 0.09722f
C14398 VPWR.t884 VGND 0.06383f
C14399 VPWR.t1773 VGND 0.07496f
C14400 VPWR.t1063 VGND 0.02709f
C14401 VPWR.t1774 VGND 0.02407f
C14402 VPWR.n2434 VGND 0.07442f
C14403 VPWR.n2436 VGND 0.088f
C14404 VPWR.t498 VGND 0.09722f
C14405 VPWR.t323 VGND 0.06383f
C14406 VPWR.t426 VGND 0.07496f
C14407 VPWR.t883 VGND 0.06383f
C14408 VPWR.t68 VGND 0.09722f
C14409 VPWR.t1882 VGND 0.02709f
C14410 VPWR.t73 VGND 0.02407f
C14411 VPWR.n2437 VGND 0.07442f
C14412 VPWR.n2439 VGND 0.0512f
C14413 VPWR.n2441 VGND 0.088f
C14414 VPWR.t72 VGND 0.07496f
C14415 VPWR.t322 VGND 0.06383f
C14416 VPWR.t1881 VGND 0.09722f
C14417 VPWR.n2442 VGND 0.088f
C14418 VPWR.n2444 VGND 0.0512f
C14419 VPWR.n2446 VGND 0.2969f
C14420 VPWR.n2447 VGND 0.06791f
C14421 VPWR.n2448 VGND 0.06791f
C14422 VPWR.n2449 VGND 0.2969f
C14423 VPWR.n2450 VGND 0.2969f
C14424 VPWR.n2451 VGND 0.06791f
C14425 VPWR.n2452 VGND 0.06791f
C14426 VPWR.n2453 VGND 0.06791f
C14427 VPWR.n2454 VGND 0.2969f
C14428 VPWR.n2455 VGND 0.2969f
C14429 VPWR.n2456 VGND 0.06791f
C14430 VPWR.n2457 VGND 0.06791f
C14431 VPWR.n2458 VGND 0.06791f
C14432 VPWR.n2459 VGND 0.06791f
C14433 VPWR.n2460 VGND 0.2969f
C14434 VPWR.n2462 VGND 0.0512f
C14435 VPWR.n2464 VGND 0.088f
C14436 VPWR.t866 VGND 0.09722f
C14437 VPWR.t156 VGND 0.06383f
C14438 VPWR.t1040 VGND 0.07496f
C14439 VPWR.t324 VGND 0.06383f
C14440 VPWR.t1573 VGND 0.09722f
C14441 VPWR.n2465 VGND 0.088f
C14442 VPWR.n2467 VGND 0.0512f
C14443 VPWR.n2469 VGND 0.0512f
C14444 VPWR.n2471 VGND 0.088f
C14445 VPWR.t301 VGND 0.09722f
C14446 VPWR.t846 VGND 0.06383f
C14447 VPWR.t1012 VGND 0.07496f
C14448 VPWR.t302 VGND 0.02709f
C14449 VPWR.t1013 VGND 0.02407f
C14450 VPWR.n2472 VGND 0.07442f
C14451 VPWR.n2474 VGND 0.0512f
C14452 VPWR.n2476 VGND 0.088f
C14453 VPWR.t1008 VGND 0.09722f
C14454 VPWR.t886 VGND 0.06383f
C14455 VPWR.t1826 VGND 0.07496f
C14456 VPWR.t321 VGND 0.06383f
C14457 VPWR.t902 VGND 0.09722f
C14458 VPWR.n2477 VGND 0.088f
C14459 VPWR.n2479 VGND 0.0512f
C14460 VPWR.n2482 VGND 0.0512f
C14461 VPWR.n2484 VGND 0.088f
C14462 VPWR.t202 VGND 0.09722f
C14463 VPWR.t320 VGND 0.06383f
C14464 VPWR.t1637 VGND 0.07496f
C14465 VPWR.t849 VGND 0.06383f
C14466 VPWR.t969 VGND 0.09722f
C14467 VPWR.n2485 VGND 0.088f
C14468 VPWR.n2487 VGND 0.0512f
C14469 VPWR.n2490 VGND 0.0512f
C14470 VPWR.n2492 VGND 0.088f
C14471 VPWR.t992 VGND 0.09722f
C14472 VPWR.t155 VGND 0.06383f
C14473 VPWR.t1443 VGND 0.10842f
C14474 VPWR.n2493 VGND 0.06192f
C14475 VPWR.n2494 VGND 0.0512f
C14476 VPWR.n2496 VGND 0.2969f
C14477 VPWR.n2497 VGND 0.15751f
C14478 VPWR.n2498 VGND 0.06791f
C14479 VPWR.n2499 VGND 0.06791f
C14480 VPWR.n2500 VGND 0.06791f
C14481 VPWR.n2501 VGND 0.06791f
C14482 VPWR.n2502 VGND 0.06791f
C14483 VPWR.n2503 VGND 0.06791f
C14484 VPWR.n2504 VGND 0.2969f
C14485 VPWR.n2505 VGND 0.06791f
C14486 VPWR.n2506 VGND 0.2969f
C14487 VPWR.t121 VGND 0.02709f
C14488 VPWR.t371 VGND 0.02407f
C14489 VPWR.n2508 VGND 0.07442f
C14490 VPWR.t1765 VGND 0.06383f
C14491 VPWR.t4 VGND 0.07496f
C14492 VPWR.t482 VGND 0.02709f
C14493 VPWR.t5 VGND 0.02407f
C14494 VPWR.n2509 VGND 0.07442f
C14495 VPWR.n2511 VGND 0.0512f
C14496 VPWR.n2513 VGND 0.088f
C14497 VPWR.t518 VGND 0.09722f
C14498 VPWR.t425 VGND 0.06383f
C14499 VPWR.t124 VGND 0.07496f
C14500 VPWR.t519 VGND 0.02709f
C14501 VPWR.t125 VGND 0.02407f
C14502 VPWR.n2514 VGND 0.07442f
C14503 VPWR.n2516 VGND 0.088f
C14504 VPWR.t120 VGND 0.09722f
C14505 VPWR.t103 VGND 0.06383f
C14506 VPWR.t370 VGND 0.07496f
C14507 VPWR.t927 VGND 0.06383f
C14508 VPWR.t1577 VGND 0.09722f
C14509 VPWR.t363 VGND 0.02709f
C14510 VPWR.t1867 VGND 0.02407f
C14511 VPWR.n2517 VGND 0.07442f
C14512 VPWR.n2518 VGND 0.0512f
C14513 VPWR.n2520 VGND 0.088f
C14514 VPWR.t1866 VGND 0.07496f
C14515 VPWR.t928 VGND 0.06383f
C14516 VPWR.t362 VGND 0.09722f
C14517 VPWR.n2521 VGND 0.088f
C14518 VPWR.n2523 VGND 0.0512f
C14519 VPWR.n2525 VGND 0.2969f
C14520 VPWR.n2526 VGND 0.06791f
C14521 VPWR.n2527 VGND 0.06791f
C14522 VPWR.n2528 VGND 0.06791f
C14523 VPWR.n2529 VGND 0.2969f
C14524 VPWR.n2531 VGND 0.0512f
C14525 VPWR.n2533 VGND 0.088f
C14526 VPWR.t459 VGND 0.07496f
C14527 VPWR.t865 VGND 0.06383f
C14528 VPWR.t169 VGND 0.09722f
C14529 VPWR.n2534 VGND 0.088f
C14530 VPWR.n2536 VGND 0.0512f
C14531 VPWR.n2538 VGND 0.0512f
C14532 VPWR.n2540 VGND 0.088f
C14533 VPWR.t1697 VGND 0.07496f
C14534 VPWR.t1766 VGND 0.06383f
C14535 VPWR.t732 VGND 0.09722f
C14536 VPWR.n2541 VGND 0.088f
C14537 VPWR.n2543 VGND 0.0512f
C14538 VPWR.n2545 VGND 0.2969f
C14539 VPWR.n2546 VGND 0.06791f
C14540 VPWR.n2547 VGND 0.06791f
C14541 VPWR.n2548 VGND 0.2969f
C14542 VPWR.n2549 VGND 0.0512f
C14543 VPWR.t966 VGND 0.02709f
C14544 VPWR.t1499 VGND 0.02407f
C14545 VPWR.n2551 VGND 0.07442f
C14546 VPWR.t611 VGND 0.118f
C14547 VPWR.t1645 VGND 0.06383f
C14548 VPWR.t1689 VGND 0.07496f
C14549 VPWR.t612 VGND 0.02709f
C14550 VPWR.t1690 VGND 0.02407f
C14551 VPWR.n2552 VGND 0.07442f
C14552 VPWR.n2553 VGND -0.05607f
C14553 VPWR.n2555 VGND 0.088f
C14554 VPWR.t1566 VGND 0.09722f
C14555 VPWR.t1670 VGND 0.06383f
C14556 VPWR.t1929 VGND 0.07496f
C14557 VPWR.t1567 VGND 0.02709f
C14558 VPWR.t1930 VGND 0.02407f
C14559 VPWR.n2556 VGND 0.07442f
C14560 VPWR.n2558 VGND 0.088f
C14561 VPWR.t965 VGND 0.09722f
C14562 VPWR.t976 VGND 0.06383f
C14563 VPWR.t1498 VGND 0.07496f
C14564 VPWR.t1644 VGND 0.06383f
C14565 VPWR.t711 VGND 0.09722f
C14566 VPWR.t1523 VGND 0.02709f
C14567 VPWR.t1796 VGND 0.02407f
C14568 VPWR.n2559 VGND 0.07442f
C14569 VPWR.n2561 VGND 0.0512f
C14570 VPWR.n2563 VGND 0.088f
C14571 VPWR.t1795 VGND 0.07496f
C14572 VPWR.t975 VGND 0.06383f
C14573 VPWR.t1522 VGND 0.09722f
C14574 VPWR.n2564 VGND 0.088f
C14575 VPWR.n2566 VGND 0.0512f
C14576 VPWR.n2568 VGND 0.06791f
C14577 VPWR.n2569 VGND 0.2969f
C14578 VPWR.n2570 VGND 0.2969f
C14579 VPWR.n2571 VGND 0.06791f
C14580 VPWR.n2572 VGND 0.06791f
C14581 VPWR.n2573 VGND 0.06791f
C14582 VPWR.n2574 VGND 0.06791f
C14583 VPWR.n2575 VGND 0.06791f
C14584 VPWR.n2576 VGND 0.06791f
C14585 VPWR.n2577 VGND 0.2969f
C14586 VPWR.n2579 VGND 0.0512f
C14587 VPWR.n2581 VGND 0.088f
C14588 VPWR.t1746 VGND 0.09722f
C14589 VPWR.t1675 VGND 0.06383f
C14590 VPWR.t1879 VGND 0.07496f
C14591 VPWR.t1674 VGND 0.06383f
C14592 VPWR.t411 VGND 0.09722f
C14593 VPWR.n2582 VGND 0.088f
C14594 VPWR.n2584 VGND 0.0512f
C14595 VPWR.n2587 VGND 0.0512f
C14596 VPWR.n2589 VGND 0.088f
C14597 VPWR.t469 VGND 0.09722f
C14598 VPWR.t1643 VGND 0.06383f
C14599 VPWR.t1709 VGND 0.07496f
C14600 VPWR.t470 VGND 0.02709f
C14601 VPWR.t1710 VGND 0.02407f
C14602 VPWR.n2590 VGND 0.07442f
C14603 VPWR.n2592 VGND 0.088f
C14604 VPWR.t0 VGND 0.09722f
C14605 VPWR.t1642 VGND 0.06383f
C14606 VPWR.t574 VGND 0.07496f
C14607 VPWR.t269 VGND 0.09722f
C14608 VPWR.t569 VGND 0.02709f
C14609 VPWR.t276 VGND 0.02407f
C14610 VPWR.n2593 VGND 0.07442f
C14611 VPWR.t270 VGND 0.02709f
C14612 VPWR.t764 VGND 0.02407f
C14613 VPWR.n2594 VGND 0.07442f
C14614 VPWR.t974 VGND 0.06383f
C14615 VPWR.t763 VGND 0.07496f
C14616 VPWR.t1542 VGND 0.09722f
C14617 VPWR.t1027 VGND 0.02709f
C14618 VPWR.t1549 VGND 0.02407f
C14619 VPWR.n2595 VGND 0.07442f
C14620 VPWR.t1543 VGND 0.02709f
C14621 VPWR.t219 VGND 0.02407f
C14622 VPWR.n2597 VGND 0.07442f
C14623 VPWR.t1673 VGND 0.06383f
C14624 VPWR.t218 VGND 0.07496f
C14625 VPWR.t1909 VGND 0.09722f
C14626 VPWR.t1057 VGND 0.02709f
C14627 VPWR.t1819 VGND 0.02407f
C14628 VPWR.n2598 VGND 0.07442f
C14629 VPWR.t1910 VGND 0.02709f
C14630 VPWR.t1007 VGND 0.02407f
C14631 VPWR.n2600 VGND 0.07442f
C14632 VPWR.t1671 VGND 0.06383f
C14633 VPWR.t1006 VGND 0.07496f
C14634 VPWR.t531 VGND 0.02709f
C14635 VPWR.t1111 VGND 0.02407f
C14636 VPWR.n2601 VGND 0.07442f
C14637 VPWR.n2602 VGND 0.0512f
C14638 VPWR.n2603 VGND 0.06192f
C14639 VPWR.t1110 VGND 0.10842f
C14640 VPWR.t1641 VGND 0.06383f
C14641 VPWR.t530 VGND 0.09722f
C14642 VPWR.n2604 VGND 0.088f
C14643 VPWR.n2606 VGND 0.0512f
C14644 VPWR.n2608 VGND 0.0512f
C14645 VPWR.n2610 VGND 0.088f
C14646 VPWR.t1818 VGND 0.07496f
C14647 VPWR.t1672 VGND 0.06383f
C14648 VPWR.t1056 VGND 0.09722f
C14649 VPWR.n2611 VGND 0.088f
C14650 VPWR.n2613 VGND 0.0512f
C14651 VPWR.n2615 VGND 0.0512f
C14652 VPWR.n2617 VGND 0.088f
C14653 VPWR.t1548 VGND 0.07496f
C14654 VPWR.t973 VGND 0.06383f
C14655 VPWR.t1026 VGND 0.09722f
C14656 VPWR.n2618 VGND 0.088f
C14657 VPWR.n2620 VGND 0.0512f
C14658 VPWR.n2622 VGND 0.0512f
C14659 VPWR.n2624 VGND 0.088f
C14660 VPWR.t275 VGND 0.07496f
C14661 VPWR.t1676 VGND 0.06383f
C14662 VPWR.t568 VGND 0.09722f
C14663 VPWR.n2625 VGND 0.088f
C14664 VPWR.n2627 VGND 0.0512f
C14665 VPWR.n2629 VGND 0.2969f
C14666 VPWR.n2630 VGND 0.06791f
C14667 VPWR.n2631 VGND 0.06791f
C14668 VPWR.n2632 VGND 0.06791f
C14669 VPWR.n2633 VGND 0.06791f
C14670 VPWR.n2634 VGND 0.06791f
C14671 VPWR.n2635 VGND 0.06791f
C14672 VPWR.n2636 VGND 0.06791f
C14673 VPWR.n2637 VGND 0.06791f
C14674 VPWR.n2638 VGND 0.2969f
C14675 VPWR.n2639 VGND 0.2969f
C14676 VPWR.n2640 VGND 0.06791f
C14677 VPWR.n2641 VGND 0.06791f
C14678 VPWR.n2642 VGND 0.2969f
C14679 VPWR.n2644 VGND 0.0512f
C14680 VPWR.n2646 VGND 0.088f
C14681 VPWR.t1600 VGND 0.09722f
C14682 VPWR.t864 VGND 0.06383f
C14683 VPWR.t1060 VGND 0.07496f
C14684 VPWR.t863 VGND 0.06383f
C14685 VPWR.t189 VGND 0.09722f
C14686 VPWR.n2647 VGND 0.088f
C14687 VPWR.n2649 VGND 0.0512f
C14688 VPWR.n2651 VGND 0.2969f
C14689 VPWR.n2652 VGND 0.06791f
C14690 VPWR.n2653 VGND 0.06791f
C14691 VPWR.n2654 VGND 0.2969f
C14692 VPWR.n2656 VGND 0.0512f
C14693 VPWR.n2658 VGND 0.088f
C14694 VPWR.t12 VGND 0.09722f
C14695 VPWR.t862 VGND 0.06383f
C14696 VPWR.t532 VGND 0.07496f
C14697 VPWR.t13 VGND 0.02709f
C14698 VPWR.t533 VGND 0.02407f
C14699 VPWR.n2659 VGND 0.07442f
C14700 VPWR.n2661 VGND 0.088f
C14701 VPWR.t582 VGND 0.09722f
C14702 VPWR.t424 VGND 0.06383f
C14703 VPWR.t1225 VGND 0.10842f
C14704 VPWR.n2662 VGND 0.06192f
C14705 VPWR.n2663 VGND 0.0512f
C14706 VPWR.n2665 VGND 0.2969f
C14707 VPWR.n2666 VGND 0.06791f
C14708 VPWR.n2667 VGND 0.15751f
C14709 VPWR.n2668 VGND 0.82597f
C14710 VPWR.n2669 VGND 0.82597f
C14711 VPWR.n2670 VGND 0.15751f
C14712 VPWR.n2671 VGND 0.2969f
C14713 VPWR.t1003 VGND 0.02709f
C14714 VPWR.t1405 VGND 0.02407f
C14715 VPWR.n2672 VGND 0.07442f
C14716 VPWR.t1763 VGND 0.06383f
C14717 VPWR.t1404 VGND 0.10842f
C14718 VPWR.n2673 VGND 0.06192f
C14719 VPWR.n2674 VGND 0.0512f
C14720 VPWR.n2676 VGND 0.2969f
C14721 VPWR.n2677 VGND 0.15751f
C14722 VPWR.n2678 VGND 0.06791f
C14723 VPWR.n2679 VGND 0.2969f
C14724 VPWR.n2681 VGND 0.0512f
C14725 VPWR.n2683 VGND 0.088f
C14726 VPWR.t1726 VGND 0.07496f
C14727 VPWR.t1736 VGND 0.06383f
C14728 VPWR.t1635 VGND 0.09722f
C14729 VPWR.n2684 VGND 0.088f
C14730 VPWR.n2686 VGND 0.0512f
C14731 VPWR.n2688 VGND 0.2969f
C14732 VPWR.n2689 VGND 0.06791f
C14733 VPWR.n2690 VGND 0.06791f
C14734 VPWR.n2691 VGND 0.2969f
C14735 VPWR.n2693 VGND 0.0512f
C14736 VPWR.n2695 VGND 0.088f
C14737 VPWR.t95 VGND 0.07496f
C14738 VPWR.t936 VGND 0.06383f
C14739 VPWR.t1020 VGND 0.09722f
C14740 VPWR.n2696 VGND 0.088f
C14741 VPWR.n2698 VGND 0.0512f
C14742 VPWR.n2700 VGND 0.2969f
C14743 VPWR.n2701 VGND 0.06791f
C14744 VPWR.n2702 VGND 0.06791f
C14745 VPWR.n2703 VGND 0.2969f
C14746 VPWR.n2705 VGND 0.0512f
C14747 VPWR.n2707 VGND 0.088f
C14748 VPWR.t895 VGND 0.07496f
C14749 VPWR.t1764 VGND 0.06383f
C14750 VPWR.t721 VGND 0.09722f
C14751 VPWR.n2708 VGND 0.088f
C14752 VPWR.n2710 VGND 0.0512f
C14753 VPWR.n2712 VGND 0.2969f
C14754 VPWR.n2713 VGND 0.06791f
C14755 VPWR.n2714 VGND 0.06791f
C14756 VPWR.n2715 VGND 0.2969f
C14757 VPWR.n2717 VGND 0.0512f
C14758 VPWR.n2719 VGND 0.088f
C14759 VPWR.t912 VGND 0.07496f
C14760 VPWR.t1740 VGND 0.06383f
C14761 VPWR.t1781 VGND 0.09722f
C14762 VPWR.n2720 VGND 0.088f
C14763 VPWR.n2722 VGND 0.0512f
C14764 VPWR.n2724 VGND 0.2969f
C14765 VPWR.n2725 VGND 0.06791f
C14766 VPWR.n2726 VGND 0.06791f
C14767 VPWR.n2727 VGND 0.2969f
C14768 VPWR.n2729 VGND 0.0512f
C14769 VPWR.n2731 VGND 0.088f
C14770 VPWR.t1480 VGND 0.07496f
C14771 VPWR.t1748 VGND 0.06383f
C14772 VPWR.t510 VGND 0.09722f
C14773 VPWR.n2732 VGND 0.088f
C14774 VPWR.n2734 VGND 0.0512f
C14775 VPWR.n2735 VGND -0.05607f
C14776 VPWR.n2736 VGND 0.2969f
C14777 VPWR.n2737 VGND 0.06791f
C14778 VPWR.n2738 VGND 0.82079f
C14779 VPWR.n2739 VGND 0.15751f
C14780 VPWR.n2740 VGND 0.06791f
C14781 VPWR.n2741 VGND 0.06791f
C14782 VPWR.n2742 VGND 0.06791f
C14783 VPWR.n2743 VGND 0.06791f
C14784 VPWR.n2744 VGND 0.06791f
C14785 VPWR.n2745 VGND 0.06791f
C14786 VPWR.n2746 VGND 0.06791f
C14787 VPWR.n2747 VGND 0.06791f
C14788 VPWR.n2748 VGND 0.06791f
C14789 VPWR.n2749 VGND 0.06791f
C14790 VPWR.n2750 VGND 0.06791f
C14791 VPWR.n2751 VGND 0.06791f
C14792 VPWR.n2752 VGND 0.06791f
C14793 VPWR.n2753 VGND 0.06791f
C14794 VPWR.n2754 VGND 0.06791f
C14795 VPWR.n2755 VGND 0.82079f
C14796 VPWR.n2756 VGND 0.46455f
C14797 VPWR.n2757 VGND 0.06791f
C14798 VPWR.n2758 VGND 0.06977f
C14799 VPWR.n2760 VGND -0.05416f
C14800 VPWR.n2762 VGND 0.088f
C14801 VPWR.t1274 VGND 0.09722f
C14802 VPWR.t1241 VGND 0.06383f
C14803 VPWR.t1374 VGND 0.07496f
C14804 VPWR.t1383 VGND 0.06383f
C14805 VPWR.t1395 VGND 0.09722f
C14806 VPWR.n2763 VGND 0.088f
C14807 VPWR.n2767 VGND 0.06977f
C14808 VPWR.n2768 VGND 0.06791f
C14809 VPWR.n2769 VGND 0.06791f
C14810 VPWR.n2770 VGND 0.06977f
C14811 VPWR.n2774 VGND 0.088f
C14812 VPWR.t1151 VGND 0.09722f
C14813 VPWR.t1417 VGND 0.06383f
C14814 VPWR.t1145 VGND 0.07496f
C14815 VPWR.t1135 VGND 0.06383f
C14816 VPWR.t1259 VGND 0.09722f
C14817 VPWR.n2775 VGND 0.088f
C14818 VPWR.n2779 VGND 0.06977f
C14819 VPWR.n2780 VGND 0.06791f
C14820 VPWR.n2781 VGND 0.06791f
C14821 VPWR.n2782 VGND 0.06977f
C14822 VPWR.n2786 VGND 0.088f
C14823 VPWR.t1271 VGND 0.09722f
C14824 VPWR.t1279 VGND 0.06383f
C14825 VPWR.t1414 VGND 0.07496f
C14826 VPWR.t1303 VGND 0.06383f
C14827 VPWR.t1427 VGND 0.09722f
C14828 VPWR.n2787 VGND 0.088f
C14829 VPWR.n2791 VGND 0.06977f
C14830 VPWR.n2792 VGND 0.06791f
C14831 VPWR.n2793 VGND 0.06791f
C14832 VPWR.n2794 VGND 0.06977f
C14833 VPWR.n2798 VGND 0.088f
C14834 VPWR.t1148 VGND 0.09722f
C14835 VPWR.t1140 VGND 0.06383f
C14836 VPWR.t1167 VGND 0.07496f
C14837 VPWR.t1175 VGND 0.06383f
C14838 VPWR.t1308 VGND 0.09722f
C14839 VPWR.n2799 VGND 0.088f
C14840 VPWR.n2803 VGND 0.06977f
C14841 VPWR.n2804 VGND 0.06791f
C14842 VPWR.n2805 VGND 0.06791f
C14843 VPWR.n2806 VGND 0.06977f
C14844 VPWR.n2810 VGND 0.088f
C14845 VPWR.t1327 VGND 0.09722f
C14846 VPWR.t1277 VGND 0.06383f
C14847 VPWR.t1366 VGND 0.07496f
C14848 VPWR.t1438 VGND 0.06383f
C14849 VPWR.t1454 VGND 0.09722f
C14850 VPWR.n2811 VGND 0.088f
C14851 VPWR.n2815 VGND 0.06977f
C14852 VPWR.n2816 VGND 0.06791f
C14853 VPWR.n2817 VGND 0.06791f
C14854 VPWR.n2818 VGND 0.06977f
C14855 VPWR.n2822 VGND 0.088f
C14856 VPWR.t1198 VGND 0.09722f
C14857 VPWR.t1457 VGND 0.06383f
C14858 VPWR.t1190 VGND 0.07496f
C14859 VPWR.t1311 VGND 0.06383f
C14860 VPWR.t1228 VGND 0.09722f
C14861 VPWR.n2823 VGND 0.088f
C14862 VPWR.n2827 VGND 0.06977f
C14863 VPWR.n2828 VGND 0.06791f
C14864 VPWR.n2829 VGND 0.06791f
C14865 VPWR.n2830 VGND 0.06977f
C14866 VPWR.n2834 VGND 0.088f
C14867 VPWR.t1078 VGND 0.09722f
C14868 VPWR.t1333 VGND 0.06383f
C14869 VPWR.t1451 VGND 0.07496f
C14870 VPWR.t1355 VGND 0.06383f
C14871 VPWR.t1097 VGND 0.09722f
C14872 VPWR.n2835 VGND 0.088f
C14873 VPWR.n2839 VGND 0.06977f
C14874 VPWR.n2840 VGND 0.06791f
C14875 VPWR.n2841 VGND 0.06791f
C14876 VPWR.n2842 VGND 0.06977f
C14877 VPWR.n2846 VGND 0.088f
C14878 VPWR.t1222 VGND 0.09722f
C14879 VPWR.t1206 VGND 0.06383f
C14880 VPWR.t1330 VGND 0.10842f
C14881 VPWR.n2847 VGND 0.06192f
C14882 VPWR.n2850 VGND 0.02435f
C14883 VPWR.n2851 VGND 0.05693f
C14884 VPWR.n2852 VGND 0.02435f
C14885 VPWR.n2853 VGND 0.13344f
C14886 VPWR.n2854 VGND 0.02435f
C14887 VPWR.n2855 VGND 0.1037f
C14888 VPWR.n2856 VGND 0.02435f
C14889 VPWR.n2857 VGND 0.1037f
C14890 VPWR.n2858 VGND 0.02435f
C14891 VPWR.n2859 VGND 0.1037f
C14892 VPWR.n2860 VGND 0.02435f
C14893 VPWR.n2861 VGND 0.1037f
C14894 VPWR.n2862 VGND 0.02435f
C14895 VPWR.n2863 VGND 0.1037f
C14896 VPWR.n2864 VGND 0.02435f
C14897 VPWR.n2865 VGND 0.1037f
C14898 VPWR.n2866 VGND 0.02435f
C14899 VPWR.n2867 VGND 0.1037f
C14900 VPWR.n2868 VGND 0.02435f
C14901 VPWR.n2869 VGND 0.1037f
C14902 VPWR.n2870 VGND 0.02435f
C14903 VPWR.n2871 VGND 0.1037f
C14904 VPWR.n2872 VGND 0.02435f
C14905 VPWR.n2873 VGND 0.1037f
C14906 VPWR.n2874 VGND 0.02435f
C14907 VPWR.n2875 VGND 0.1037f
C14908 VPWR.n2876 VGND 0.02435f
C14909 VPWR.n2877 VGND 0.1037f
C14910 VPWR.n2878 VGND 0.02435f
C14911 VPWR.n2879 VGND 0.1037f
C14912 VPWR.n2880 VGND 0.02435f
C14913 VPWR.n2881 VGND 0.11228f
C14914 VPWR.n2882 VGND 0.09374f
C14915 VPWR.n2883 VGND 0.08766f
C14916 VPWR.n2884 VGND 0.15751f
C14917 VPWR.n2885 VGND 2.16512f
C14918 VPWR.n2886 VGND 0.88173f
C14919 VPWR.n2887 VGND 0.36944f
C14920 VPWR.t643 VGND 0.04436f
C14921 VPWR.t137 VGND 0.04436f
C14922 VPWR.n2888 VGND 0.08048f
C14923 VPWR.n2889 VGND 0.03811f
C14924 VPWR.t642 VGND 0.01165f
C14925 VPWR.t646 VGND 0.01165f
C14926 VPWR.n2890 VGND 0.02501f
C14927 VPWR.t147 VGND 0.01165f
C14928 VPWR.t135 VGND 0.01165f
C14929 VPWR.n2891 VGND 0.02501f
C14930 VPWR.n2893 VGND 0.03811f
C14931 VPWR.t1885 VGND 0.01165f
C14932 VPWR.t979 VGND 0.01165f
C14933 VPWR.n2894 VGND 0.02501f
C14934 VPWR.t351 VGND 0.01165f
C14935 VPWR.t406 VGND 0.01165f
C14936 VPWR.n2895 VGND 0.02501f
C14937 VPWR.t983 VGND 0.04646f
C14938 VPWR.t238 VGND 0.04646f
C14939 VPWR.n2896 VGND 0.10714f
C14940 VPWR.n2897 VGND 0.03438f
C14941 VPWR.n2898 VGND 0.01108f
C14942 VPWR.n2899 VGND 0.05028f
C14943 VPWR.t236 VGND 0.01165f
C14944 VPWR.t645 VGND 0.01165f
C14945 VPWR.n2901 VGND 0.02501f
C14946 VPWR.t400 VGND 0.01165f
C14947 VPWR.t143 VGND 0.01165f
C14948 VPWR.n2902 VGND 0.02501f
C14949 VPWR.n2903 VGND 0.05028f
C14950 VPWR.n2904 VGND 0.01159f
C14951 VPWR.n2905 VGND 0.03811f
C14952 VPWR.n2906 VGND 0.03811f
C14953 VPWR.n2907 VGND 0.03811f
C14954 VPWR.n2908 VGND 0.01042f
C14955 VPWR.n2909 VGND 0.05028f
C14956 VPWR.n2912 VGND 0.03811f
C14957 VPWR.n2913 VGND 0.02858f
C14958 VPWR.t237 VGND 0.13921f
C14959 VPWR.t350 VGND 0.20515f
C14960 VPWR.t405 VGND 0.20515f
C14961 VPWR.t235 VGND 0.20515f
C14962 VPWR.t142 VGND 0.20515f
C14963 VPWR.t146 VGND 0.20515f
C14964 VPWR.t134 VGND 0.20515f
C14965 VPWR.t136 VGND 0.45673f
C14966 VPWR.n2915 VGND 0.49851f
C14967 VPWR.n2916 VGND 0.0145f
C14968 VPWR.n2917 VGND 0.87438f
C14969 VPWR.n2918 VGND 0.03811f
C14970 VPWR.t239 VGND 0.13921f
C14971 VPWR.t346 VGND 0.20515f
C14972 VPWR.t261 VGND 0.20515f
C14973 VPWR.t286 VGND 0.20515f
C14974 VPWR.t539 VGND 0.20515f
C14975 VPWR.t549 VGND 0.20515f
C14976 VPWR.t541 VGND 0.20515f
C14977 VPWR.t551 VGND 0.33703f
C14978 VPWR.t258 VGND 0.35779f
C14979 VPWR.n2919 VGND 0.5049f
C14980 VPWR.n2920 VGND 0.14363f
C14981 VPWR.n2921 VGND 0.03811f
C14982 VPWR.t550 VGND 0.01165f
C14983 VPWR.t542 VGND 0.01165f
C14984 VPWR.n2922 VGND 0.02501f
C14985 VPWR.t854 VGND 0.01165f
C14986 VPWR.t860 VGND 0.01165f
C14987 VPWR.n2923 VGND 0.02501f
C14988 VPWR.n2924 VGND 0.05028f
C14989 VPWR.n2925 VGND 0.03811f
C14990 VPWR.t287 VGND 0.01165f
C14991 VPWR.t540 VGND 0.01165f
C14992 VPWR.n2926 VGND 0.02501f
C14993 VPWR.t388 VGND 0.01165f
C14994 VPWR.t858 VGND 0.01165f
C14995 VPWR.n2927 VGND 0.02501f
C14996 VPWR.t240 VGND 0.04646f
C14997 VPWR.t288 VGND 0.04646f
C14998 VPWR.n2929 VGND 0.10714f
C14999 VPWR.t396 VGND 0.01165f
C15000 VPWR.t353 VGND 0.01165f
C15001 VPWR.n2930 VGND 0.02501f
C15002 VPWR.t347 VGND 0.01165f
C15003 VPWR.t262 VGND 0.01165f
C15004 VPWR.n2931 VGND 0.02501f
C15005 VPWR.n2932 VGND 0.05028f
C15006 VPWR.n2933 VGND 0.01108f
C15007 VPWR.n2934 VGND 0.03438f
C15008 VPWR.n2935 VGND 0.03811f
C15009 VPWR.n2936 VGND 0.03811f
C15010 VPWR.n2937 VGND 0.01159f
C15011 VPWR.n2938 VGND 0.05028f
C15012 VPWR.n2940 VGND 0.01042f
C15013 VPWR.n2941 VGND 0.03811f
C15014 VPWR.n2942 VGND 0.03811f
C15015 VPWR.t552 VGND 0.04436f
C15016 VPWR.t856 VGND 0.04436f
C15017 VPWR.n2945 VGND 0.08048f
C15018 VPWR.n2947 VGND 0.02858f
C15019 VPWR.n2948 VGND 0.0145f
C15020 VPWR.n2949 VGND 0.02858f
C15021 VPWR.n2950 VGND 0.01137f
C15022 VPWR.t259 VGND 0.04641f
C15023 VPWR.t1568 VGND 0.04641f
C15024 VPWR.n2952 VGND 0.09381f
C15025 VPWR.n2953 VGND 0.02651f
C15026 VPWR.n2954 VGND 1.33077f
C15027 VPWR.n2955 VGND 0.03811f
C15028 VPWR.t182 VGND 0.04556f
C15029 VPWR.t289 VGND 0.13921f
C15030 VPWR.t336 VGND 0.20515f
C15031 VPWR.t281 VGND 0.20515f
C15032 VPWR.t391 VGND 0.20515f
C15033 VPWR.t48 VGND 0.20515f
C15034 VPWR.t42 VGND 0.20515f
C15035 VPWR.t50 VGND 0.20515f
C15036 VPWR.t44 VGND 0.33703f
C15037 VPWR.t1552 VGND 0.12944f
C15038 VPWR.t181 VGND 0.10257f
C15039 VPWR.t640 VGND 0.22835f
C15040 VPWR.n2956 VGND 0.44751f
C15041 VPWR.n2957 VGND 0.1415f
C15042 VPWR.n2958 VGND 0.03811f
C15043 VPWR.t43 VGND 0.01165f
C15044 VPWR.t51 VGND 0.01165f
C15045 VPWR.n2959 VGND 0.02501f
C15046 VPWR.t374 VGND 0.01165f
C15047 VPWR.t378 VGND 0.01165f
C15048 VPWR.n2960 VGND 0.02501f
C15049 VPWR.n2961 VGND 0.05028f
C15050 VPWR.n2962 VGND 0.03811f
C15051 VPWR.t392 VGND 0.01165f
C15052 VPWR.t49 VGND 0.01165f
C15053 VPWR.n2963 VGND 0.02501f
C15054 VPWR.t404 VGND 0.01165f
C15055 VPWR.t377 VGND 0.01165f
C15056 VPWR.n2964 VGND 0.02501f
C15057 VPWR.t290 VGND 0.04646f
C15058 VPWR.t393 VGND 0.04646f
C15059 VPWR.n2966 VGND 0.10714f
C15060 VPWR.t349 VGND 0.01165f
C15061 VPWR.t282 VGND 0.01165f
C15062 VPWR.n2967 VGND 0.02501f
C15063 VPWR.t337 VGND 0.01165f
C15064 VPWR.t1890 VGND 0.01165f
C15065 VPWR.n2968 VGND 0.02501f
C15066 VPWR.n2969 VGND 0.05028f
C15067 VPWR.n2970 VGND 0.01108f
C15068 VPWR.n2971 VGND 0.03438f
C15069 VPWR.n2972 VGND 0.03811f
C15070 VPWR.n2973 VGND 0.03811f
C15071 VPWR.n2974 VGND 0.01159f
C15072 VPWR.n2975 VGND 0.05028f
C15073 VPWR.n2977 VGND 0.01042f
C15074 VPWR.n2978 VGND 0.03811f
C15075 VPWR.n2979 VGND 0.03811f
C15076 VPWR.t45 VGND 0.04436f
C15077 VPWR.t375 VGND 0.04436f
C15078 VPWR.n2982 VGND 0.08048f
C15079 VPWR.n2984 VGND 0.02858f
C15080 VPWR.n2985 VGND 0.0145f
C15081 VPWR.n2986 VGND 0.02858f
C15082 VPWR.t641 VGND 0.04646f
C15083 VPWR.n2987 VGND 0.06475f
C15084 VPWR.n2989 VGND 0.04738f
C15085 VPWR.t1553 VGND 0.04568f
C15086 VPWR.n2990 VGND 0.0592f
C15087 VPWR.n2991 VGND 0.02258f
C15088 VPWR.n2992 VGND 1.33077f
C15089 VPWR.n2993 VGND 0.03811f
C15090 VPWR.t389 VGND 0.07895f
C15091 VPWR.t333 VGND 0.11635f
C15092 VPWR.t1888 VGND 0.11311f
C15093 VPWR.t402 VGND 0.1809f
C15094 VPWR.t477 VGND 0.15386f
C15095 VPWR.t981 VGND 0.10257f
C15096 VPWR.t1728 VGND 0.10257f
C15097 VPWR.t242 VGND 0.10257f
C15098 VPWR.t1028 VGND 0.10257f
C15099 VPWR.t977 VGND 0.10257f
C15100 VPWR.t28 VGND 0.10257f
C15101 VPWR.t283 VGND 0.14287f
C15102 VPWR.t706 VGND 0.08059f
C15103 VPWR.t1873 VGND 0.08792f
C15104 VPWR.t638 VGND 0.10257f
C15105 VPWR.t1875 VGND 0.19049f
C15106 VPWR.n2994 VGND 0.30708f
C15107 VPWR.n2995 VGND 0.14164f
C15108 VPWR.t1876 VGND 0.04612f
C15109 VPWR.n2996 VGND 0.03811f
C15110 VPWR.t284 VGND 0.04559f
C15111 VPWR.t29 VGND 0.04389f
C15112 VPWR.t243 VGND 0.01165f
C15113 VPWR.t978 VGND 0.01165f
C15114 VPWR.n2997 VGND 0.02501f
C15115 VPWR.t1729 VGND 0.01165f
C15116 VPWR.t1029 VGND 0.01165f
C15117 VPWR.n2998 VGND 0.02501f
C15118 VPWR.n2999 VGND 0.02851f
C15119 VPWR.n3000 VGND 0.03811f
C15120 VPWR.t403 VGND 0.01165f
C15121 VPWR.t478 VGND 0.01165f
C15122 VPWR.n3001 VGND 0.02501f
C15123 VPWR.t390 VGND 0.04646f
C15124 VPWR.n3003 VGND 0.05855f
C15125 VPWR.t334 VGND 0.01165f
C15126 VPWR.t1889 VGND 0.01165f
C15127 VPWR.n3004 VGND 0.02501f
C15128 VPWR.n3005 VGND 0.02851f
C15129 VPWR.n3006 VGND 0.01108f
C15130 VPWR.n3007 VGND 0.03438f
C15131 VPWR.n3008 VGND 0.03811f
C15132 VPWR.n3009 VGND 0.03811f
C15133 VPWR.n3010 VGND 0.01159f
C15134 VPWR.n3011 VGND 0.02785f
C15135 VPWR.t982 VGND 0.04078f
C15136 VPWR.n3012 VGND 0.03251f
C15137 VPWR.n3014 VGND 0.03811f
C15138 VPWR.n3015 VGND 0.03811f
C15139 VPWR.n3016 VGND 0.03159f
C15140 VPWR.n3018 VGND 0.04182f
C15141 VPWR.n3019 VGND 0.05509f
C15142 VPWR.n3021 VGND 0.02258f
C15143 VPWR.n3022 VGND 0.0145f
C15144 VPWR.n3023 VGND 0.02858f
C15145 VPWR.t639 VGND 0.04651f
C15146 VPWR.n3024 VGND 0.11958f
C15147 VPWR.t1874 VGND 0.04644f
C15148 VPWR.n3026 VGND 0.05169f
C15149 VPWR.n3027 VGND 0.02237f
C15150 VPWR.n3028 VGND 1.33077f
C15151 VPWR.n3029 VGND 0.03438f
C15152 VPWR.t395 VGND 0.54218f
C15153 VPWR.t280 VGND 0.20515f
C15154 VPWR.t401 VGND 0.20515f
C15155 VPWR.t332 VGND 0.20515f
C15156 VPWR.t140 VGND 0.20515f
C15157 VPWR.t138 VGND 0.20515f
C15158 VPWR.t144 VGND 0.20515f
C15159 VPWR.t132 VGND 0.18561f
C15160 VPWR.t34 VGND 0.44937f
C15161 VPWR.t631 VGND 0.12455f
C15162 VPWR.n3030 VGND 0.26923f
C15163 VPWR.n3031 VGND 0.14363f
C15164 VPWR.t647 VGND 0.01165f
C15165 VPWR.t644 VGND 0.01165f
C15166 VPWR.n3032 VGND 0.02554f
C15167 VPWR.t141 VGND 0.01165f
C15168 VPWR.t139 VGND 0.01165f
C15169 VPWR.n3033 VGND 0.02554f
C15170 VPWR.n3034 VGND 0.09692f
C15171 VPWR.n3035 VGND 0.07858f
C15172 VPWR.t648 VGND 0.01165f
C15173 VPWR.t649 VGND 0.01165f
C15174 VPWR.n3036 VGND 0.02558f
C15175 VPWR.t145 VGND 0.01165f
C15176 VPWR.t133 VGND 0.01165f
C15177 VPWR.n3037 VGND 0.02558f
C15178 VPWR.n3038 VGND 0.10624f
C15179 VPWR.n3040 VGND 0.30689f
C15180 VPWR.n3041 VGND 0.0145f
C15181 VPWR.n3042 VGND 0.01326f
C15182 VPWR.n3043 VGND 0.01137f
C15183 VPWR.n3044 VGND 0.01064f
C15184 VPWR.t35 VGND 0.04651f
C15185 VPWR.t456 VGND 0.04651f
C15186 VPWR.n3045 VGND 0.13737f
C15187 VPWR.n3046 VGND 0.02858f
C15188 VPWR.n3047 VGND 1.33077f
C15189 VPWR.n3048 VGND 0.03438f
C15190 VPWR.t348 VGND 0.54218f
C15191 VPWR.t1887 VGND 0.20515f
C15192 VPWR.t241 VGND 0.20515f
C15193 VPWR.t1886 VGND 0.20515f
C15194 VPWR.t543 VGND 0.20515f
C15195 VPWR.t553 VGND 0.20515f
C15196 VPWR.t545 VGND 0.20515f
C15197 VPWR.t547 VGND 0.18561f
C15198 VPWR.t959 VGND 0.39931f
C15199 VPWR.t633 VGND 0.08792f
C15200 VPWR.t637 VGND 0.0867f
C15201 VPWR.n3049 VGND 0.268f
C15202 VPWR.n3050 VGND 0.14363f
C15203 VPWR.t544 VGND 0.01165f
C15204 VPWR.t554 VGND 0.01165f
C15205 VPWR.n3051 VGND 0.02554f
C15206 VPWR.t853 VGND 0.01165f
C15207 VPWR.t859 VGND 0.01165f
C15208 VPWR.n3052 VGND 0.02554f
C15209 VPWR.n3053 VGND 0.09692f
C15210 VPWR.n3054 VGND 0.07858f
C15211 VPWR.t546 VGND 0.01165f
C15212 VPWR.t548 VGND 0.01165f
C15213 VPWR.n3055 VGND 0.02558f
C15214 VPWR.t855 VGND 0.01165f
C15215 VPWR.t857 VGND 0.01165f
C15216 VPWR.n3056 VGND 0.02558f
C15217 VPWR.n3057 VGND 0.10624f
C15218 VPWR.n3059 VGND 0.30689f
C15219 VPWR.n3060 VGND 0.0145f
C15220 VPWR.n3061 VGND 0.01305f
C15221 VPWR.t634 VGND 0.04641f
C15222 VPWR.n3063 VGND 0.04961f
C15223 VPWR.t960 VGND 0.04651f
C15224 VPWR.n3065 VGND 0.07408f
C15225 VPWR.n3066 VGND 0.02858f
C15226 VPWR.n3067 VGND 1.33077f
C15227 VPWR.n3068 VGND 0.0348f
C15228 VPWR.t335 VGND 0.54218f
C15229 VPWR.t234 VGND 0.20515f
C15230 VPWR.t394 VGND 0.20515f
C15231 VPWR.t352 VGND 0.20515f
C15232 VPWR.t52 VGND 0.20515f
C15233 VPWR.t46 VGND 0.20515f
C15234 VPWR.t38 VGND 0.20515f
C15235 VPWR.t40 VGND 0.18561f
C15236 VPWR.t36 VGND 0.42495f
C15237 VPWR.t629 VGND 0.14654f
C15238 VPWR.n3069 VGND 0.26678f
C15239 VPWR.n3070 VGND 0.1415f
C15240 VPWR.t632 VGND 0.04648f
C15241 VPWR.t53 VGND 0.01165f
C15242 VPWR.t47 VGND 0.01165f
C15243 VPWR.n3071 VGND 0.02554f
C15244 VPWR.t379 VGND 0.01165f
C15245 VPWR.t376 VGND 0.01165f
C15246 VPWR.n3072 VGND 0.02554f
C15247 VPWR.n3073 VGND 0.09692f
C15248 VPWR.n3074 VGND 0.07858f
C15249 VPWR.t39 VGND 0.01165f
C15250 VPWR.t41 VGND 0.01165f
C15251 VPWR.n3075 VGND 0.02558f
C15252 VPWR.t372 VGND 0.01165f
C15253 VPWR.t373 VGND 0.01165f
C15254 VPWR.n3076 VGND 0.02558f
C15255 VPWR.n3077 VGND 0.10624f
C15256 VPWR.n3079 VGND 0.30689f
C15257 VPWR.n3080 VGND 0.0145f
C15258 VPWR.n3081 VGND 0.01284f
C15259 VPWR.t630 VGND 0.04648f
C15260 VPWR.n3082 VGND 0.12245f
C15261 VPWR.t37 VGND 0.04646f
C15262 VPWR.t455 VGND 0.04646f
C15263 VPWR.n3084 VGND 0.10933f
C15264 VPWR.n3085 VGND 0.02858f
C15265 VPWR.n3086 VGND 1.33077f
C15266 VPWR.n3087 VGND 0.0348f
C15267 VPWR.t958 VGND 0.04646f
C15268 VPWR.n3088 VGND 0.01284f
C15269 VPWR.t636 VGND 0.04648f
C15270 VPWR.n3089 VGND 0.0145f
C15271 VPWR.t980 VGND 0.30749f
C15272 VPWR.t285 VGND 0.11635f
C15273 VPWR.t345 VGND 0.11635f
C15274 VPWR.t260 VGND 0.11635f
C15275 VPWR.t1030 VGND 0.11635f
C15276 VPWR.t148 VGND 0.11635f
C15277 VPWR.t1923 VGND 0.11635f
C15278 VPWR.t967 VGND 0.10527f
C15279 VPWR.t957 VGND 0.24101f
C15280 VPWR.t635 VGND 0.08311f
C15281 VPWR.n3090 VGND 0.14848f
C15282 VPWR.t1924 VGND 0.01165f
C15283 VPWR.t968 VGND 0.01165f
C15284 VPWR.n3091 VGND 0.02558f
C15285 VPWR.n3092 VGND 0.06295f
C15286 VPWR.t1031 VGND 0.01165f
C15287 VPWR.t149 VGND 0.01165f
C15288 VPWR.n3093 VGND 0.02662f
C15289 VPWR.n3094 VGND 0.14214f
C15290 VPWR.n3095 VGND 0.30689f
C15291 VPWR.n3097 VGND 0.07856f
C15292 VPWR.n3098 VGND 0.06897f
C15293 VPWR.n3100 VGND 0.05976f
C15294 VPWR.n3101 VGND 0.02858f
C15295 VPWR.n3102 VGND 1.14955f
C15296 VPWR.n3103 VGND 1.34319f
C15297 VPWR.n3104 VGND 0.08514f
C15298 VPWR.t833 VGND 1.49101f
C15299 VPWR.t222 VGND 0.89906f
C15300 VPWR.n3105 VGND 1.13436f
C15301 VPWR.t592 VGND 1.94178f
C15302 VPWR.n3106 VGND 0.08514f
C15303 VPWR.t593 VGND 0.03926f
C15304 VPWR.n3107 VGND 0.24351f
C15305 VPWR.n3108 VGND 0.15076f
C15306 VPWR.n3109 VGND 1.07739f
C15307 VPWR.n3110 VGND 0.15076f
C15308 VPWR.n3111 VGND 0.08514f
C15309 VPWR.t594 VGND 0.03926f
C15310 VPWR.n3112 VGND 0.24351f
C15311 VPWR.n3113 VGND 0.17097f
C15312 VPWR.n3114 VGND 0.32322f
C15313 VPWR.n3115 VGND 0.09594f
C15314 VPWR.n3116 VGND 0.18244f
C15315 VPWR.n3117 VGND 0.0998f
C15316 VPWR.n3118 VGND 0.10634f
C15317 VPWR.n3119 VGND 0.15076f
C15318 VPWR.n3120 VGND 0.70588f
C15319 VPWR.n3121 VGND 0.15076f
C15320 VPWR.n3122 VGND 0.10634f
C15321 VPWR.n3123 VGND 0.08792f
C15322 VPWR.t882 VGND 0.011f
C15323 VPWR.t834 VGND 0.011f
C15324 VPWR.n3124 VGND 0.02201f
C15325 VPWR.n3125 VGND 0.01833f
C15326 VPWR.n3126 VGND 0.01817f
C15327 VPWR.n3127 VGND 0.09653f
C15328 VPWR.n3128 VGND 0.29252f
C15329 VPWR.n3129 VGND 0.3134f
C15330 VPWR.n3130 VGND 0.33069f
C15331 VPWR.n3131 VGND 2.063f
C15332 XThR.Tn[2].t9 VGND 0.0218f
C15333 XThR.Tn[2].t4 VGND 0.0218f
C15334 XThR.Tn[2].n0 VGND 0.05148f
C15335 XThR.Tn[2].t11 VGND 0.0218f
C15336 XThR.Tn[2].t0 VGND 0.0218f
C15337 XThR.Tn[2].n1 VGND 0.044f
C15338 XThR.Tn[2].n2 VGND 0.15443f
C15339 XThR.Tn[2].t7 VGND 0.01417f
C15340 XThR.Tn[2].t8 VGND 0.01417f
C15341 XThR.Tn[2].n3 VGND 0.05376f
C15342 XThR.Tn[2].t6 VGND 0.01417f
C15343 XThR.Tn[2].t5 VGND 0.01417f
C15344 XThR.Tn[2].n4 VGND 0.03227f
C15345 XThR.Tn[2].n5 VGND 0.15366f
C15346 XThR.Tn[2].t3 VGND 0.01417f
C15347 XThR.Tn[2].t1 VGND 0.01417f
C15348 XThR.Tn[2].n6 VGND 0.03227f
C15349 XThR.Tn[2].n7 VGND 0.09499f
C15350 XThR.Tn[2].t10 VGND 0.01417f
C15351 XThR.Tn[2].t2 VGND 0.01417f
C15352 XThR.Tn[2].n8 VGND 0.03227f
C15353 XThR.Tn[2].n9 VGND 0.10721f
C15354 XThR.Tn[2].t21 VGND 0.01704f
C15355 XThR.Tn[2].t14 VGND 0.01866f
C15356 XThR.Tn[2].n10 VGND 0.04556f
C15357 XThR.Tn[2].n11 VGND 0.0708f
C15358 XThR.Tn[2].t40 VGND 0.01704f
C15359 XThR.Tn[2].t31 VGND 0.01866f
C15360 XThR.Tn[2].n12 VGND 0.04556f
C15361 XThR.Tn[2].t55 VGND 0.01698f
C15362 XThR.Tn[2].t66 VGND 0.0186f
C15363 XThR.Tn[2].n13 VGND 0.0474f
C15364 XThR.Tn[2].n14 VGND 0.0333f
C15365 XThR.Tn[2].n16 VGND 0.10686f
C15366 XThR.Tn[2].t15 VGND 0.01704f
C15367 XThR.Tn[2].t67 VGND 0.01866f
C15368 XThR.Tn[2].n17 VGND 0.04556f
C15369 XThR.Tn[2].t30 VGND 0.01698f
C15370 XThR.Tn[2].t43 VGND 0.0186f
C15371 XThR.Tn[2].n18 VGND 0.0474f
C15372 XThR.Tn[2].n19 VGND 0.0333f
C15373 XThR.Tn[2].n21 VGND 0.10686f
C15374 XThR.Tn[2].t32 VGND 0.01704f
C15375 XThR.Tn[2].t23 VGND 0.01866f
C15376 XThR.Tn[2].n22 VGND 0.04556f
C15377 XThR.Tn[2].t47 VGND 0.01698f
C15378 XThR.Tn[2].t60 VGND 0.0186f
C15379 XThR.Tn[2].n23 VGND 0.0474f
C15380 XThR.Tn[2].n24 VGND 0.0333f
C15381 XThR.Tn[2].n26 VGND 0.10686f
C15382 XThR.Tn[2].t58 VGND 0.01704f
C15383 XThR.Tn[2].t50 VGND 0.01866f
C15384 XThR.Tn[2].n27 VGND 0.04556f
C15385 XThR.Tn[2].t16 VGND 0.01698f
C15386 XThR.Tn[2].t28 VGND 0.0186f
C15387 XThR.Tn[2].n28 VGND 0.0474f
C15388 XThR.Tn[2].n29 VGND 0.0333f
C15389 XThR.Tn[2].n31 VGND 0.10686f
C15390 XThR.Tn[2].t34 VGND 0.01704f
C15391 XThR.Tn[2].t25 VGND 0.01866f
C15392 XThR.Tn[2].n32 VGND 0.04556f
C15393 XThR.Tn[2].t48 VGND 0.01698f
C15394 XThR.Tn[2].t62 VGND 0.0186f
C15395 XThR.Tn[2].n33 VGND 0.0474f
C15396 XThR.Tn[2].n34 VGND 0.0333f
C15397 XThR.Tn[2].n36 VGND 0.10686f
C15398 XThR.Tn[2].t70 VGND 0.01704f
C15399 XThR.Tn[2].t41 VGND 0.01866f
C15400 XThR.Tn[2].n37 VGND 0.04556f
C15401 XThR.Tn[2].t22 VGND 0.01698f
C15402 XThR.Tn[2].t20 VGND 0.0186f
C15403 XThR.Tn[2].n38 VGND 0.0474f
C15404 XThR.Tn[2].n39 VGND 0.0333f
C15405 XThR.Tn[2].n41 VGND 0.10686f
C15406 XThR.Tn[2].t39 VGND 0.01704f
C15407 XThR.Tn[2].t35 VGND 0.01866f
C15408 XThR.Tn[2].n42 VGND 0.04556f
C15409 XThR.Tn[2].t54 VGND 0.01698f
C15410 XThR.Tn[2].t12 VGND 0.0186f
C15411 XThR.Tn[2].n43 VGND 0.0474f
C15412 XThR.Tn[2].n44 VGND 0.0333f
C15413 XThR.Tn[2].n46 VGND 0.10686f
C15414 XThR.Tn[2].t44 VGND 0.01704f
C15415 XThR.Tn[2].t49 VGND 0.01866f
C15416 XThR.Tn[2].n47 VGND 0.04556f
C15417 XThR.Tn[2].t57 VGND 0.01698f
C15418 XThR.Tn[2].t27 VGND 0.0186f
C15419 XThR.Tn[2].n48 VGND 0.0474f
C15420 XThR.Tn[2].n49 VGND 0.0333f
C15421 XThR.Tn[2].n51 VGND 0.10686f
C15422 XThR.Tn[2].t61 VGND 0.01704f
C15423 XThR.Tn[2].t69 VGND 0.01866f
C15424 XThR.Tn[2].n52 VGND 0.04556f
C15425 XThR.Tn[2].t18 VGND 0.01698f
C15426 XThR.Tn[2].t45 VGND 0.0186f
C15427 XThR.Tn[2].n53 VGND 0.0474f
C15428 XThR.Tn[2].n54 VGND 0.0333f
C15429 XThR.Tn[2].n56 VGND 0.10686f
C15430 XThR.Tn[2].t52 VGND 0.01704f
C15431 XThR.Tn[2].t26 VGND 0.01866f
C15432 XThR.Tn[2].n57 VGND 0.04556f
C15433 XThR.Tn[2].t68 VGND 0.01698f
C15434 XThR.Tn[2].t63 VGND 0.0186f
C15435 XThR.Tn[2].n58 VGND 0.0474f
C15436 XThR.Tn[2].n59 VGND 0.0333f
C15437 XThR.Tn[2].n61 VGND 0.10686f
C15438 XThR.Tn[2].t73 VGND 0.01704f
C15439 XThR.Tn[2].t64 VGND 0.01866f
C15440 XThR.Tn[2].n62 VGND 0.04556f
C15441 XThR.Tn[2].t24 VGND 0.01698f
C15442 XThR.Tn[2].t37 VGND 0.0186f
C15443 XThR.Tn[2].n63 VGND 0.0474f
C15444 XThR.Tn[2].n64 VGND 0.0333f
C15445 XThR.Tn[2].n66 VGND 0.10686f
C15446 XThR.Tn[2].t42 VGND 0.01704f
C15447 XThR.Tn[2].t36 VGND 0.01866f
C15448 XThR.Tn[2].n67 VGND 0.04556f
C15449 XThR.Tn[2].t56 VGND 0.01698f
C15450 XThR.Tn[2].t13 VGND 0.0186f
C15451 XThR.Tn[2].n68 VGND 0.0474f
C15452 XThR.Tn[2].n69 VGND 0.0333f
C15453 XThR.Tn[2].n71 VGND 0.10686f
C15454 XThR.Tn[2].t59 VGND 0.01704f
C15455 XThR.Tn[2].t51 VGND 0.01866f
C15456 XThR.Tn[2].n72 VGND 0.04556f
C15457 XThR.Tn[2].t17 VGND 0.01698f
C15458 XThR.Tn[2].t29 VGND 0.0186f
C15459 XThR.Tn[2].n73 VGND 0.0474f
C15460 XThR.Tn[2].n74 VGND 0.0333f
C15461 XThR.Tn[2].n76 VGND 0.10686f
C15462 XThR.Tn[2].t19 VGND 0.01704f
C15463 XThR.Tn[2].t72 VGND 0.01866f
C15464 XThR.Tn[2].n77 VGND 0.04556f
C15465 XThR.Tn[2].t33 VGND 0.01698f
C15466 XThR.Tn[2].t46 VGND 0.0186f
C15467 XThR.Tn[2].n78 VGND 0.0474f
C15468 XThR.Tn[2].n79 VGND 0.0333f
C15469 XThR.Tn[2].n81 VGND 0.10686f
C15470 XThR.Tn[2].t53 VGND 0.01704f
C15471 XThR.Tn[2].t65 VGND 0.01866f
C15472 XThR.Tn[2].n82 VGND 0.04556f
C15473 XThR.Tn[2].t71 VGND 0.01698f
C15474 XThR.Tn[2].t38 VGND 0.0186f
C15475 XThR.Tn[2].n83 VGND 0.0474f
C15476 XThR.Tn[2].n84 VGND 0.0333f
C15477 XThR.Tn[2].n86 VGND 0.10686f
C15478 XThR.Tn[2].n87 VGND 0.09711f
C15479 XThR.Tn[2].n88 VGND 0.21044f
.ends

