magic
tech sky130A
magscale 1 2
timestamp 1760335364
<< locali >>
rect -688 -6230 -640 -6226
rect -688 -6270 -684 -6230
rect -644 -6270 -640 -6230
rect 400 -6234 450 -6216
rect -688 -6274 -640 -6270
rect 400 -6284 412 -6234
rect 1488 -6230 1536 -6226
rect 3056 -6230 3104 -6214
rect 1488 -6270 1492 -6230
rect 1532 -6270 1536 -6230
rect 3056 -6264 3064 -6230
rect 3098 -6264 3104 -6230
rect 772 -6276 820 -6270
rect 1488 -6274 1536 -6270
rect -786 -6312 -738 -6306
rect -786 -6346 -780 -6312
rect -746 -6346 -738 -6312
rect -786 -6354 -738 -6346
rect -316 -6312 -268 -6306
rect -316 -6346 -310 -6312
rect -276 -6346 -268 -6312
rect -316 -6354 -268 -6346
rect 302 -6312 350 -6306
rect 302 -6346 308 -6312
rect 342 -6346 350 -6312
rect 772 -6310 778 -6276
rect 812 -6310 820 -6276
rect 3056 -6282 3104 -6264
rect 3466 -6230 3514 -6226
rect 3466 -6270 3470 -6230
rect 3510 -6270 3514 -6230
rect 3466 -6274 3514 -6270
rect 772 -6318 820 -6310
rect 302 -6354 350 -6346
rect 3056 -6330 3104 -6318
rect 880 -6358 928 -6350
rect 880 -6392 886 -6358
rect 920 -6392 928 -6358
rect 400 -6404 452 -6394
rect 880 -6398 928 -6392
rect 400 -6438 408 -6404
rect 442 -6438 452 -6404
rect 400 -6446 452 -6438
rect 1390 -6402 1438 -6396
rect 1390 -6436 1396 -6402
rect 1430 -6436 1438 -6402
rect 1390 -6444 1438 -6436
rect 1488 -6404 1536 -6396
rect 1488 -6438 1494 -6404
rect 1528 -6438 1536 -6404
rect 1488 -6444 1536 -6438
rect 1968 -6404 2016 -6396
rect 1968 -6438 1974 -6404
rect 2008 -6438 2016 -6404
rect 1968 -6444 2016 -6438
rect 2126 -6402 2174 -6396
rect 2126 -6436 2134 -6402
rect 2168 -6436 2174 -6402
rect 2126 -6444 2174 -6436
rect 2418 -6402 2466 -6396
rect 2418 -6436 2424 -6402
rect 2458 -6436 2466 -6402
rect 2418 -6444 2466 -6436
rect 2576 -6404 2624 -6396
rect 2576 -6438 2582 -6404
rect 2616 -6438 2624 -6404
rect 2576 -6444 2624 -6438
rect 3056 -6442 3060 -6330
rect 3100 -6442 3104 -6330
rect 5110 -6366 5344 -6360
rect 5110 -6414 5122 -6366
rect 5332 -6414 5344 -6366
rect 5110 -6420 5344 -6414
rect 3056 -6454 3104 -6442
rect 874 -6464 922 -6458
rect -684 -6500 -636 -6494
rect -684 -6534 -678 -6500
rect -644 -6534 -636 -6500
rect -684 -6542 -636 -6534
rect -214 -6500 -166 -6494
rect -214 -6534 -208 -6500
rect -174 -6534 -166 -6500
rect -214 -6542 -166 -6534
rect 404 -6500 452 -6494
rect 404 -6534 410 -6500
rect 444 -6534 452 -6500
rect 874 -6498 880 -6464
rect 914 -6498 922 -6464
rect 874 -6506 922 -6498
rect 404 -6542 452 -6534
rect -679 -6632 -639 -6542
rect -209 -6632 -169 -6542
rect 409 -6680 449 -6542
rect 879 -6596 919 -6506
rect 1492 -6518 1540 -6512
rect 1492 -6552 1498 -6518
rect 1532 -6552 1540 -6518
rect 1492 -6560 1540 -6552
rect 1964 -6518 2012 -6512
rect 1964 -6552 1972 -6518
rect 2006 -6552 2012 -6518
rect 1964 -6560 2012 -6552
rect 2580 -6518 2628 -6512
rect 2580 -6552 2586 -6518
rect 2620 -6552 2628 -6518
rect 2580 -6560 2628 -6552
rect 1497 -6650 1537 -6560
rect 1967 -6650 2007 -6560
rect 2585 -6650 2625 -6560
rect 3056 -6630 3100 -6454
rect 3668 -6498 3732 -6492
rect 3668 -6538 3680 -6498
rect 3720 -6538 3732 -6498
rect 3668 -6606 3732 -6538
rect 4132 -6566 4188 -6560
rect 4132 -6606 4140 -6566
rect 4180 -6606 4188 -6566
rect 4132 -6612 4188 -6606
rect 879 -6748 919 -6696
rect 5228 -6702 5280 -6688
rect 5228 -6742 5234 -6702
rect 5274 -6742 5280 -6702
rect 5228 -6756 5280 -6742
rect 1497 -6816 1537 -6764
rect 1969 -6884 2009 -6832
rect 2585 -6952 2625 -6900
rect 2984 -6952 3176 -6946
rect 2984 -7016 2990 -6952
rect 3170 -7016 3176 -6952
rect 2984 -7022 3176 -7016
rect -772 -7302 -570 -7296
rect -772 -7380 -766 -7302
rect -576 -7380 -570 -7302
rect -772 -7386 -570 -7380
rect -278 -7302 -76 -7296
rect -278 -7380 -272 -7302
rect -82 -7380 -76 -7302
rect -278 -7386 -76 -7380
<< viali >>
rect -684 -6270 -644 -6230
rect -202 -6266 -166 -6230
rect 412 -6284 450 -6234
rect 1492 -6270 1532 -6230
rect 1974 -6266 2010 -6230
rect 2583 -6268 2617 -6234
rect 3064 -6264 3098 -6230
rect -780 -6346 -746 -6312
rect -310 -6346 -276 -6312
rect 308 -6346 342 -6312
rect 778 -6310 812 -6276
rect 3470 -6270 3510 -6230
rect 3672 -6266 3706 -6232
rect 4760 -6266 4796 -6230
rect 4146 -6316 4186 -6276
rect 5236 -6312 5272 -6276
rect 5846 -6312 5882 -6276
rect 886 -6392 920 -6358
rect -678 -6438 -644 -6404
rect -204 -6438 -170 -6404
rect 408 -6438 442 -6404
rect 1396 -6436 1430 -6402
rect 1494 -6438 1528 -6404
rect 1974 -6438 2008 -6404
rect 2134 -6436 2168 -6402
rect 2424 -6436 2458 -6402
rect 2582 -6438 2616 -6404
rect 3060 -6442 3100 -6330
rect 4266 -6384 4306 -6344
rect 4849 -6357 4889 -6317
rect 3672 -6436 3706 -6402
rect 4756 -6440 4796 -6400
rect 5122 -6414 5332 -6366
rect 5778 -6402 5886 -6366
rect -678 -6534 -644 -6500
rect -208 -6534 -174 -6500
rect 410 -6534 444 -6500
rect 880 -6498 914 -6464
rect 1498 -6552 1532 -6518
rect 1972 -6552 2006 -6518
rect 2586 -6552 2620 -6518
rect 3680 -6538 3720 -6498
rect 4140 -6606 4180 -6566
rect 4758 -6672 4794 -6636
rect 5234 -6742 5274 -6702
rect 3060 -6898 3100 -6786
rect 5844 -6810 5884 -6770
rect 6324 -6866 6364 -6826
rect 6940 -6866 6980 -6826
rect 2990 -7016 3170 -6952
rect 3600 -6998 3708 -6914
rect 4148 -6998 4256 -6914
rect 4688 -6998 4796 -6914
rect 5236 -6998 5344 -6914
rect 5776 -6998 5884 -6914
rect 6324 -6998 6432 -6914
rect 6864 -6998 6972 -6914
rect -676 -7254 -640 -7214
rect -208 -7254 -172 -7214
rect 412 -7254 448 -7214
rect 880 -7254 916 -7214
rect 1500 -7254 1536 -7214
rect 1970 -7254 2006 -7214
rect 2588 -7254 2624 -7214
rect -766 -7380 -576 -7302
rect -272 -7380 -82 -7302
rect 322 -7368 512 -7302
rect 816 -7368 1006 -7302
rect 1410 -7368 1600 -7302
rect 1904 -7368 2094 -7302
rect 2498 -7368 2688 -7302
rect 3670 -7364 3706 -7324
rect 4150 -7364 4186 -7324
rect 4758 -7364 4794 -7324
rect 5238 -7364 5274 -7324
rect 5846 -7364 5882 -7324
rect 6326 -7364 6362 -7324
rect 6934 -7364 6970 -7324
<< metal1 >>
rect -1016 -5914 -920 -5908
rect -1016 -6142 -1010 -5914
rect -926 -6142 -920 -5914
rect -1016 -6202 -920 -6142
rect -472 -5914 -376 -5908
rect -472 -6142 -466 -5914
rect -382 -6142 -376 -5914
rect -472 -6202 -376 -6142
rect 72 -5914 168 -5908
rect 72 -6142 78 -5914
rect 162 -6142 168 -5914
rect 72 -6202 168 -6142
rect 616 -5914 712 -5908
rect 616 -6142 622 -5914
rect 706 -6142 712 -5914
rect 616 -6202 712 -6142
rect 1160 -5914 1256 -5908
rect 1160 -6142 1166 -5914
rect 1250 -6142 1256 -5914
rect 1160 -6202 1256 -6142
rect 1704 -5914 1800 -5908
rect 1704 -6142 1710 -5914
rect 1794 -6142 1800 -5914
rect 1704 -6202 1800 -6142
rect 2248 -5914 2344 -5908
rect 2248 -6142 2254 -5914
rect 2338 -6142 2344 -5914
rect 2248 -6202 2344 -6142
rect 2792 -5914 2888 -5908
rect 2792 -6142 2798 -5914
rect 2882 -6142 2888 -5914
rect 2792 -6202 2888 -6142
rect 3336 -5914 3432 -5908
rect 3336 -6142 3342 -5914
rect 3426 -6142 3432 -5914
rect 3336 -6202 3432 -6142
rect 1966 -6218 2018 -6212
rect -690 -6224 -638 -6218
rect -690 -6282 -638 -6276
rect -208 -6230 -160 -6218
rect -208 -6266 -202 -6230
rect -166 -6266 -160 -6230
rect -788 -6312 -736 -6298
rect -788 -6346 -780 -6312
rect -746 -6346 -736 -6312
rect -788 -6362 -736 -6346
rect -318 -6312 -266 -6298
rect -318 -6346 -310 -6312
rect -276 -6346 -266 -6312
rect -318 -6362 -266 -6346
rect -208 -6304 -160 -6266
rect 406 -6234 456 -6222
rect 1486 -6224 1538 -6218
rect 406 -6284 412 -6234
rect 450 -6284 551 -6234
rect 406 -6296 456 -6284
rect -208 -6356 -116 -6304
rect -64 -6356 -58 -6304
rect 300 -6312 352 -6298
rect 300 -6346 308 -6312
rect 342 -6346 352 -6312
rect 300 -6362 352 -6346
rect -776 -6504 -748 -6362
rect -688 -6394 -636 -6388
rect -688 -6452 -636 -6446
rect -686 -6492 -634 -6486
rect -692 -6504 -686 -6492
rect -776 -6532 -686 -6504
rect -692 -6544 -686 -6532
rect -634 -6544 -628 -6492
rect -306 -6504 -278 -6362
rect -212 -6394 -160 -6388
rect -212 -6452 -160 -6446
rect -216 -6500 -164 -6486
rect -216 -6504 -208 -6500
rect -306 -6532 -208 -6504
rect -216 -6534 -208 -6532
rect -174 -6534 -164 -6500
rect 312 -6504 340 -6362
rect 400 -6394 452 -6388
rect 400 -6452 452 -6446
rect 402 -6500 454 -6486
rect 402 -6504 410 -6500
rect 312 -6532 410 -6504
rect -686 -6550 -634 -6544
rect -216 -6560 -164 -6534
rect 402 -6534 410 -6532
rect 444 -6534 454 -6500
rect -222 -6612 -216 -6560
rect -164 -6612 -158 -6560
rect -216 -6632 -164 -6612
rect 402 -6628 454 -6534
rect 396 -6680 402 -6628
rect 454 -6680 460 -6628
rect 402 -6700 454 -6680
rect 501 -6982 551 -6284
rect 770 -6276 822 -6262
rect 770 -6310 778 -6276
rect 812 -6310 822 -6276
rect 1486 -6282 1538 -6276
rect 1848 -6230 2018 -6218
rect 1848 -6266 1974 -6230
rect 2010 -6266 2018 -6230
rect 1848 -6282 2018 -6266
rect 2571 -6234 2629 -6228
rect 2571 -6268 2583 -6234
rect 2617 -6236 2629 -6234
rect 3056 -6230 3246 -6214
rect 2617 -6265 2735 -6236
rect 2617 -6268 2629 -6265
rect 2571 -6274 2629 -6268
rect 770 -6326 822 -6310
rect 1848 -6304 1912 -6282
rect 1966 -6284 2018 -6282
rect 782 -6468 810 -6326
rect 878 -6358 930 -6342
rect 1848 -6356 1854 -6304
rect 1906 -6356 1912 -6304
rect 878 -6392 886 -6358
rect 920 -6366 930 -6358
rect 920 -6392 1036 -6366
rect 2706 -6383 2735 -6265
rect 3056 -6264 3064 -6230
rect 3098 -6264 3246 -6230
rect 3056 -6274 3246 -6264
rect 3056 -6276 3104 -6274
rect 3054 -6330 3106 -6304
rect 878 -6394 1036 -6392
rect 878 -6408 978 -6394
rect 972 -6446 978 -6408
rect 1030 -6446 1036 -6394
rect 1388 -6402 1440 -6388
rect 1388 -6436 1396 -6402
rect 1430 -6436 1440 -6402
rect 872 -6464 924 -6450
rect 1388 -6452 1440 -6436
rect 1486 -6394 1538 -6388
rect 1486 -6452 1538 -6446
rect 1966 -6394 2018 -6388
rect 1966 -6452 2018 -6446
rect 2124 -6402 2176 -6388
rect 2124 -6436 2134 -6402
rect 2168 -6436 2176 -6402
rect 2124 -6452 2176 -6436
rect 2416 -6402 2468 -6388
rect 2416 -6436 2424 -6402
rect 2458 -6436 2468 -6402
rect 2416 -6452 2468 -6436
rect 2574 -6394 2626 -6388
rect 2574 -6452 2626 -6446
rect 2694 -6389 2746 -6383
rect 2694 -6447 2746 -6441
rect 3054 -6442 3060 -6330
rect 3100 -6442 3106 -6330
rect 872 -6468 880 -6464
rect 782 -6496 880 -6468
rect 872 -6498 880 -6496
rect 914 -6498 924 -6464
rect 872 -6514 924 -6498
rect 874 -6696 924 -6514
rect 1400 -6522 1428 -6452
rect 1490 -6518 1542 -6504
rect 1490 -6522 1498 -6518
rect 1400 -6550 1498 -6522
rect 1490 -6552 1498 -6550
rect 1532 -6552 1542 -6518
rect 866 -6748 872 -6696
rect 924 -6748 930 -6696
rect 1490 -6764 1542 -6552
rect 1962 -6518 2014 -6504
rect 1962 -6552 1972 -6518
rect 2006 -6522 2014 -6518
rect 2136 -6522 2164 -6452
rect 2006 -6550 2164 -6522
rect 2428 -6522 2456 -6452
rect 2578 -6518 2630 -6504
rect 2578 -6522 2586 -6518
rect 2428 -6550 2586 -6522
rect 2006 -6552 2014 -6550
rect 1484 -6816 1490 -6764
rect 1542 -6816 1548 -6764
rect 1962 -6832 2014 -6552
rect 2578 -6552 2586 -6550
rect 2620 -6552 2630 -6518
rect 1956 -6884 1962 -6832
rect 2014 -6884 2020 -6832
rect 2578 -6900 2630 -6552
rect 2572 -6952 2578 -6900
rect 2630 -6952 2636 -6900
rect 2706 -6977 2735 -6447
rect 3054 -6786 3106 -6442
rect 3186 -6428 3246 -6274
rect 3464 -6224 3516 -6218
rect 3464 -6282 3516 -6276
rect 3590 -6368 3630 -5510
rect 3672 -6212 3712 -5510
rect 3880 -5914 3976 -5908
rect 3880 -6142 3886 -5914
rect 3970 -6142 3976 -5914
rect 3880 -6202 3976 -6142
rect 4424 -5914 4520 -5908
rect 4424 -6142 4430 -5914
rect 4514 -6142 4520 -5914
rect 4424 -6202 4520 -6142
rect 4968 -5914 5064 -5908
rect 4968 -6142 4974 -5914
rect 5058 -6142 5064 -5914
rect 4968 -6202 5064 -6142
rect 3662 -6226 3714 -6212
rect 4752 -6222 4804 -6216
rect 3662 -6284 3714 -6278
rect 4140 -6270 4192 -6264
rect 5238 -6260 5278 -5510
rect 5512 -5914 5608 -5908
rect 5512 -6142 5518 -5914
rect 5602 -6142 5608 -5914
rect 5512 -6202 5608 -6142
rect 5848 -6260 5888 -5510
rect 6056 -5914 6152 -5908
rect 6056 -6142 6062 -5914
rect 6146 -6142 6152 -5914
rect 6056 -6202 6152 -6142
rect 6600 -5914 6696 -5908
rect 6600 -6142 6606 -5914
rect 6690 -6142 6696 -5914
rect 4752 -6280 4804 -6274
rect 5230 -6276 5278 -6260
rect 4140 -6328 4192 -6322
rect 3466 -6420 3472 -6368
rect 3524 -6384 3630 -6368
rect 3524 -6402 3714 -6384
rect 4254 -6390 4260 -6338
rect 4312 -6390 4318 -6338
rect 4837 -6363 4843 -6311
rect 4895 -6363 4901 -6311
rect 5230 -6312 5236 -6276
rect 5272 -6312 5278 -6276
rect 5230 -6326 5278 -6312
rect 5840 -6276 5888 -6260
rect 5840 -6312 5846 -6276
rect 5882 -6312 5888 -6276
rect 5840 -6326 5888 -6312
rect 3524 -6420 3672 -6402
rect 3590 -6436 3672 -6420
rect 3706 -6436 3714 -6402
rect 3590 -6456 3714 -6436
rect 4744 -6446 4750 -6394
rect 4802 -6446 4808 -6394
rect 5110 -6420 5116 -6360
rect 5338 -6420 5344 -6360
rect 5766 -6366 6004 -6360
rect 5766 -6402 5778 -6366
rect 5886 -6402 6004 -6366
rect 5766 -6408 6004 -6402
rect 3186 -6494 3246 -6488
rect 3668 -6544 3674 -6492
rect 3726 -6544 3732 -6492
rect 4128 -6612 4134 -6560
rect 4186 -6612 4192 -6560
rect 4744 -6680 4750 -6628
rect 4802 -6680 4808 -6628
rect 5222 -6696 5286 -6688
rect 5222 -6756 5286 -6748
rect 3054 -6898 3060 -6786
rect 3100 -6860 3106 -6786
rect 5832 -6816 5838 -6764
rect 5890 -6816 5896 -6764
rect 3100 -6898 3296 -6860
rect 3054 -6912 3296 -6898
rect 2984 -6952 3196 -6940
rect 494 -7034 500 -6982
rect 552 -7034 558 -6982
rect 2695 -6983 2747 -6977
rect 501 -7059 551 -7034
rect 2695 -7041 2747 -7035
rect 2984 -7016 2990 -6952
rect 3170 -7016 3196 -6952
rect 3244 -6992 3296 -6912
rect 3498 -6914 3714 -6902
rect -690 -7260 -684 -7208
rect -632 -7260 -626 -7208
rect -222 -7260 -216 -7208
rect -164 -7260 -158 -7208
rect 398 -7260 404 -7208
rect 456 -7260 462 -7208
rect 866 -7260 872 -7208
rect 924 -7260 930 -7208
rect 1486 -7260 1492 -7208
rect 1544 -7260 1550 -7208
rect 1956 -7260 1962 -7208
rect 2014 -7260 2020 -7208
rect 2574 -7260 2580 -7208
rect 2632 -7260 2638 -7208
rect -778 -7302 -564 -7290
rect -778 -7380 -766 -7302
rect -576 -7380 -564 -7302
rect -778 -7430 -564 -7380
rect -284 -7302 -70 -7290
rect -284 -7380 -272 -7302
rect -82 -7380 -70 -7302
rect -284 -7430 -70 -7380
rect 310 -7302 524 -7290
rect 310 -7368 322 -7302
rect 512 -7368 524 -7302
rect 310 -7430 524 -7368
rect 804 -7302 1018 -7290
rect 804 -7368 816 -7302
rect 1006 -7368 1018 -7302
rect 804 -7430 1018 -7368
rect 1398 -7302 1612 -7290
rect 1398 -7368 1410 -7302
rect 1600 -7368 1612 -7302
rect 1398 -7430 1612 -7368
rect 1892 -7302 2106 -7290
rect 1892 -7368 1904 -7302
rect 2094 -7368 2106 -7302
rect 1892 -7430 2106 -7368
rect 2486 -7302 2700 -7290
rect 2486 -7368 2498 -7302
rect 2688 -7368 2700 -7302
rect 2486 -7430 2700 -7368
rect 2984 -7430 3196 -7016
rect 3238 -6998 3302 -6992
rect 3238 -7050 3244 -6998
rect 3296 -7050 3302 -6998
rect 3238 -7056 3302 -7050
rect 3498 -6998 3600 -6914
rect 3708 -6998 3714 -6914
rect 3498 -7012 3714 -6998
rect 4142 -6914 4358 -6902
rect 4142 -6998 4148 -6914
rect 4256 -6998 4358 -6914
rect 4142 -7012 4358 -6998
rect 3498 -7430 3628 -7012
rect 3656 -7370 3662 -7318
rect 3714 -7370 3720 -7318
rect 4136 -7370 4142 -7318
rect 4194 -7370 4200 -7318
rect 4228 -7430 4358 -7012
rect 4586 -6914 4802 -6902
rect 4586 -6998 4688 -6914
rect 4796 -6998 4802 -6914
rect 4586 -7012 4802 -6998
rect 5230 -6914 5446 -6902
rect 5230 -6998 5236 -6914
rect 5344 -6998 5446 -6914
rect 5230 -7012 5446 -6998
rect 4586 -7430 4716 -7012
rect 4744 -7370 4750 -7318
rect 4802 -7370 4808 -7318
rect 5224 -7370 5230 -7318
rect 5282 -7370 5288 -7318
rect 5316 -7430 5446 -7012
rect 5674 -6914 5890 -6902
rect 5674 -6998 5776 -6914
rect 5884 -6998 5890 -6914
rect 5956 -6990 6004 -6408
rect 6600 -6482 6696 -6142
rect 7144 -5914 7240 -5908
rect 7144 -6142 7150 -5914
rect 7234 -6142 7240 -5914
rect 7144 -6482 7240 -6142
rect 6312 -6872 6318 -6820
rect 6370 -6872 6376 -6820
rect 6928 -6872 6934 -6820
rect 6986 -6872 6992 -6820
rect 6318 -6914 6534 -6902
rect 5674 -7012 5890 -6998
rect 5954 -6996 6006 -6990
rect 5674 -7430 5804 -7012
rect 6318 -6998 6324 -6914
rect 6432 -6998 6534 -6914
rect 6318 -7012 6534 -6998
rect 5954 -7054 6006 -7048
rect 5832 -7370 5838 -7318
rect 5890 -7370 5896 -7318
rect 6312 -7370 6318 -7318
rect 6370 -7370 6376 -7318
rect 6404 -7430 6534 -7012
rect 6762 -6914 6978 -6902
rect 6762 -6998 6864 -6914
rect 6972 -6998 6978 -6914
rect 6762 -7012 6978 -6998
rect 6762 -7430 6892 -7012
rect 6920 -7370 6926 -7318
rect 6978 -7370 6984 -7318
<< via1 >>
rect -1010 -6142 -926 -5914
rect -466 -6142 -382 -5914
rect 78 -6142 162 -5914
rect 622 -6142 706 -5914
rect 1166 -6142 1250 -5914
rect 1710 -6142 1794 -5914
rect 2254 -6142 2338 -5914
rect 2798 -6142 2882 -5914
rect 3342 -6142 3426 -5914
rect -690 -6230 -638 -6224
rect -690 -6270 -684 -6230
rect -684 -6270 -644 -6230
rect -644 -6270 -638 -6230
rect -690 -6276 -638 -6270
rect 1486 -6230 1538 -6224
rect -116 -6356 -64 -6304
rect -688 -6404 -636 -6394
rect -688 -6438 -678 -6404
rect -678 -6438 -644 -6404
rect -644 -6438 -636 -6404
rect -688 -6446 -636 -6438
rect -686 -6500 -634 -6492
rect -686 -6534 -678 -6500
rect -678 -6534 -644 -6500
rect -644 -6534 -634 -6500
rect -686 -6544 -634 -6534
rect -212 -6404 -160 -6394
rect -212 -6438 -204 -6404
rect -204 -6438 -170 -6404
rect -170 -6438 -160 -6404
rect -212 -6446 -160 -6438
rect 400 -6404 452 -6394
rect 400 -6438 408 -6404
rect 408 -6438 442 -6404
rect 442 -6438 452 -6404
rect 400 -6446 452 -6438
rect -216 -6612 -164 -6560
rect 402 -6680 454 -6628
rect 1486 -6270 1492 -6230
rect 1492 -6270 1532 -6230
rect 1532 -6270 1538 -6230
rect 1486 -6276 1538 -6270
rect 1854 -6356 1906 -6304
rect 978 -6446 1030 -6394
rect 1486 -6404 1538 -6394
rect 1486 -6438 1494 -6404
rect 1494 -6438 1528 -6404
rect 1528 -6438 1538 -6404
rect 1486 -6446 1538 -6438
rect 1966 -6404 2018 -6394
rect 1966 -6438 1974 -6404
rect 1974 -6438 2008 -6404
rect 2008 -6438 2018 -6404
rect 1966 -6446 2018 -6438
rect 2574 -6404 2626 -6394
rect 2574 -6438 2582 -6404
rect 2582 -6438 2616 -6404
rect 2616 -6438 2626 -6404
rect 2574 -6446 2626 -6438
rect 2694 -6441 2746 -6389
rect 872 -6748 924 -6696
rect 1490 -6816 1542 -6764
rect 1962 -6884 2014 -6832
rect 2578 -6952 2630 -6900
rect 3464 -6230 3516 -6224
rect 3464 -6270 3470 -6230
rect 3470 -6270 3510 -6230
rect 3510 -6270 3516 -6230
rect 3464 -6276 3516 -6270
rect 3886 -6142 3970 -5914
rect 4430 -6142 4514 -5914
rect 4974 -6142 5058 -5914
rect 3662 -6232 3714 -6226
rect 3662 -6266 3672 -6232
rect 3672 -6266 3706 -6232
rect 3706 -6266 3714 -6232
rect 4752 -6230 4804 -6222
rect 3662 -6278 3714 -6266
rect 4140 -6276 4192 -6270
rect 4140 -6316 4146 -6276
rect 4146 -6316 4186 -6276
rect 4186 -6316 4192 -6276
rect 4752 -6266 4760 -6230
rect 4760 -6266 4796 -6230
rect 4796 -6266 4804 -6230
rect 5518 -6142 5602 -5914
rect 6062 -6142 6146 -5914
rect 6606 -6142 6690 -5914
rect 4752 -6274 4804 -6266
rect 4140 -6322 4192 -6316
rect 3472 -6420 3524 -6368
rect 4260 -6344 4312 -6338
rect 4260 -6384 4266 -6344
rect 4266 -6384 4306 -6344
rect 4306 -6384 4312 -6344
rect 4260 -6390 4312 -6384
rect 4843 -6317 4895 -6311
rect 4843 -6357 4849 -6317
rect 4849 -6357 4889 -6317
rect 4889 -6357 4895 -6317
rect 4843 -6363 4895 -6357
rect 3186 -6488 3246 -6428
rect 4750 -6400 4802 -6394
rect 4750 -6440 4756 -6400
rect 4756 -6440 4796 -6400
rect 4796 -6440 4802 -6400
rect 4750 -6446 4802 -6440
rect 5116 -6366 5338 -6360
rect 5116 -6414 5122 -6366
rect 5122 -6414 5332 -6366
rect 5332 -6414 5338 -6366
rect 5116 -6420 5338 -6414
rect 3674 -6498 3726 -6492
rect 3674 -6538 3680 -6498
rect 3680 -6538 3720 -6498
rect 3720 -6538 3726 -6498
rect 3674 -6544 3726 -6538
rect 4134 -6566 4186 -6560
rect 4134 -6606 4140 -6566
rect 4140 -6606 4180 -6566
rect 4180 -6606 4186 -6566
rect 4134 -6612 4186 -6606
rect 4750 -6636 4802 -6628
rect 4750 -6672 4758 -6636
rect 4758 -6672 4794 -6636
rect 4794 -6672 4802 -6636
rect 4750 -6680 4802 -6672
rect 5222 -6702 5286 -6696
rect 5222 -6742 5234 -6702
rect 5234 -6742 5274 -6702
rect 5274 -6742 5286 -6702
rect 5222 -6748 5286 -6742
rect 5838 -6770 5890 -6764
rect 5838 -6810 5844 -6770
rect 5844 -6810 5884 -6770
rect 5884 -6810 5890 -6770
rect 5838 -6816 5890 -6810
rect 500 -7034 552 -6982
rect 2695 -7035 2747 -6983
rect -684 -7214 -632 -7208
rect -684 -7254 -676 -7214
rect -676 -7254 -640 -7214
rect -640 -7254 -632 -7214
rect -684 -7260 -632 -7254
rect -216 -7214 -164 -7208
rect -216 -7254 -208 -7214
rect -208 -7254 -172 -7214
rect -172 -7254 -164 -7214
rect -216 -7260 -164 -7254
rect 404 -7214 456 -7208
rect 404 -7254 412 -7214
rect 412 -7254 448 -7214
rect 448 -7254 456 -7214
rect 404 -7260 456 -7254
rect 872 -7214 924 -7208
rect 872 -7254 880 -7214
rect 880 -7254 916 -7214
rect 916 -7254 924 -7214
rect 872 -7260 924 -7254
rect 1492 -7214 1544 -7208
rect 1492 -7254 1500 -7214
rect 1500 -7254 1536 -7214
rect 1536 -7254 1544 -7214
rect 1492 -7260 1544 -7254
rect 1962 -7214 2014 -7208
rect 1962 -7254 1970 -7214
rect 1970 -7254 2006 -7214
rect 2006 -7254 2014 -7214
rect 1962 -7260 2014 -7254
rect 2580 -7214 2632 -7208
rect 2580 -7254 2588 -7214
rect 2588 -7254 2624 -7214
rect 2624 -7254 2632 -7214
rect 2580 -7260 2632 -7254
rect 3244 -7050 3296 -6998
rect 3662 -7324 3714 -7318
rect 3662 -7364 3670 -7324
rect 3670 -7364 3706 -7324
rect 3706 -7364 3714 -7324
rect 3662 -7370 3714 -7364
rect 4142 -7324 4194 -7318
rect 4142 -7364 4150 -7324
rect 4150 -7364 4186 -7324
rect 4186 -7364 4194 -7324
rect 4142 -7370 4194 -7364
rect 4750 -7324 4802 -7318
rect 4750 -7364 4758 -7324
rect 4758 -7364 4794 -7324
rect 4794 -7364 4802 -7324
rect 4750 -7370 4802 -7364
rect 5230 -7324 5282 -7318
rect 5230 -7364 5238 -7324
rect 5238 -7364 5274 -7324
rect 5274 -7364 5282 -7324
rect 5230 -7370 5282 -7364
rect 7150 -6142 7234 -5914
rect 6318 -6826 6370 -6820
rect 6318 -6866 6324 -6826
rect 6324 -6866 6364 -6826
rect 6364 -6866 6370 -6826
rect 6318 -6872 6370 -6866
rect 6934 -6826 6986 -6820
rect 6934 -6866 6940 -6826
rect 6940 -6866 6980 -6826
rect 6980 -6866 6986 -6826
rect 6934 -6872 6986 -6866
rect 5954 -7048 6006 -6996
rect 5838 -7324 5890 -7318
rect 5838 -7364 5846 -7324
rect 5846 -7364 5882 -7324
rect 5882 -7364 5890 -7324
rect 5838 -7370 5890 -7364
rect 6318 -7324 6370 -7318
rect 6318 -7364 6326 -7324
rect 6326 -7364 6362 -7324
rect 6362 -7364 6370 -7324
rect 6318 -7370 6370 -7364
rect 6926 -7324 6978 -7318
rect 6926 -7364 6934 -7324
rect 6934 -7364 6970 -7324
rect 6970 -7364 6978 -7324
rect 6926 -7370 6978 -7364
<< metal2 >>
rect -1016 -5914 -920 -5908
rect -1016 -6142 -1010 -5914
rect -926 -6142 -920 -5914
rect -1016 -6148 -920 -6142
rect -472 -5914 -376 -5908
rect -472 -6142 -466 -5914
rect -382 -6142 -376 -5914
rect -472 -6148 -376 -6142
rect 72 -5914 168 -5908
rect 72 -6142 78 -5914
rect 162 -6142 168 -5914
rect 72 -6148 168 -6142
rect 616 -5914 712 -5908
rect 616 -6142 622 -5914
rect 706 -6142 712 -5914
rect 616 -6148 712 -6142
rect 1160 -5914 1256 -5908
rect 1160 -6142 1166 -5914
rect 1250 -6142 1256 -5914
rect 1160 -6148 1256 -6142
rect 1704 -5914 1800 -5908
rect 1704 -6142 1710 -5914
rect 1794 -6142 1800 -5914
rect 1704 -6148 1800 -6142
rect 2248 -5914 2344 -5908
rect 2248 -6142 2254 -5914
rect 2338 -6142 2344 -5914
rect 2248 -6148 2344 -6142
rect 2792 -5914 2888 -5908
rect 2792 -6142 2798 -5914
rect 2882 -6142 2888 -5914
rect 2792 -6148 2888 -6142
rect 3336 -5914 3432 -5908
rect 3336 -6142 3342 -5914
rect 3426 -6142 3432 -5914
rect 3336 -6148 3432 -6142
rect 3880 -5914 3976 -5908
rect 3880 -6142 3886 -5914
rect 3970 -6142 3976 -5914
rect 3880 -6148 3976 -6142
rect 4424 -5914 4520 -5908
rect 4424 -6142 4430 -5914
rect 4514 -6142 4520 -5914
rect 4424 -6148 4520 -6142
rect 4968 -5914 5064 -5908
rect 4968 -6142 4974 -5914
rect 5058 -6142 5064 -5914
rect 4968 -6148 5064 -6142
rect 5512 -5914 5608 -5908
rect 5512 -6142 5518 -5914
rect 5602 -6142 5608 -5914
rect 5512 -6148 5608 -6142
rect 6056 -5914 6152 -5908
rect 6056 -6142 6062 -5914
rect 6146 -6142 6152 -5914
rect 6056 -6148 6152 -6142
rect 6600 -5914 6696 -5908
rect 6600 -6142 6606 -5914
rect 6690 -6142 6696 -5914
rect 6600 -6148 6696 -6142
rect 7144 -5914 7240 -5908
rect 7144 -6142 7150 -5914
rect 7234 -6142 7240 -5914
rect 7144 -6148 7240 -6142
rect -690 -6224 -638 -6218
rect 1486 -6224 1538 -6218
rect -638 -6264 1486 -6236
rect -690 -6282 -638 -6276
rect 3464 -6224 3516 -6218
rect 1538 -6264 3464 -6236
rect 1486 -6282 1538 -6276
rect 3464 -6282 3516 -6276
rect 3662 -6226 3714 -6220
rect 4752 -6222 4804 -6216
rect 3714 -6266 4752 -6238
rect 3662 -6284 3714 -6278
rect 4140 -6270 4192 -6266
rect -122 -6356 -116 -6304
rect -64 -6316 -58 -6304
rect 1848 -6316 1854 -6304
rect -64 -6344 1854 -6316
rect -64 -6356 -58 -6344
rect 1848 -6356 1854 -6344
rect 1906 -6312 1912 -6304
rect 1906 -6340 4068 -6312
rect 4752 -6280 4804 -6274
rect 4140 -6328 4192 -6322
rect 4843 -6311 4895 -6305
rect 1906 -6356 1912 -6340
rect 4040 -6356 4068 -6340
rect 4254 -6356 4260 -6338
rect 2480 -6392 2556 -6382
rect 2480 -6394 2490 -6392
rect -694 -6446 -688 -6394
rect -636 -6446 -212 -6394
rect -160 -6446 400 -6394
rect 452 -6446 978 -6394
rect 1030 -6446 1486 -6394
rect 1538 -6446 1966 -6394
rect 2018 -6446 2490 -6394
rect 2480 -6448 2490 -6446
rect 2546 -6394 2556 -6392
rect 2546 -6446 2574 -6394
rect 2626 -6446 2632 -6394
rect 2688 -6441 2694 -6389
rect 2746 -6401 2752 -6389
rect 3118 -6400 3328 -6372
rect 3118 -6401 3146 -6400
rect 2746 -6430 3146 -6401
rect 2746 -6441 2752 -6430
rect 2546 -6448 2556 -6446
rect 2480 -6458 2556 -6448
rect 3174 -6488 3186 -6428
rect 3254 -6488 3266 -6428
rect 3300 -6448 3328 -6400
rect 3466 -6420 3472 -6368
rect 3524 -6380 3530 -6368
rect 3524 -6408 3866 -6380
rect 4040 -6384 4260 -6356
rect 4254 -6390 4260 -6384
rect 4312 -6390 4318 -6338
rect 4843 -6369 4895 -6363
rect 3524 -6420 3530 -6408
rect 3838 -6418 3866 -6408
rect 4744 -6418 4750 -6394
rect 3606 -6448 3790 -6436
rect 3838 -6446 4750 -6418
rect 4802 -6446 4808 -6394
rect 3300 -6464 3790 -6448
rect 3300 -6476 3632 -6464
rect 3761 -6485 3790 -6464
rect 4855 -6485 4884 -6369
rect 5110 -6420 5116 -6360
rect 5338 -6420 5344 -6360
rect -692 -6544 -686 -6492
rect -634 -6504 -628 -6492
rect 3668 -6504 3674 -6492
rect -634 -6516 3146 -6504
rect 3300 -6516 3674 -6504
rect -634 -6532 3674 -6516
rect -634 -6544 -628 -6532
rect 3118 -6544 3328 -6532
rect 3668 -6544 3674 -6532
rect 3726 -6544 3732 -6492
rect 3761 -6514 4884 -6485
rect -222 -6612 -216 -6560
rect -164 -6572 -158 -6560
rect 4128 -6572 4134 -6560
rect -164 -6600 4134 -6572
rect -164 -6612 -158 -6600
rect 4128 -6612 4134 -6600
rect 4186 -6612 4192 -6560
rect 396 -6680 402 -6628
rect 454 -6640 460 -6628
rect 4744 -6640 4750 -6628
rect 454 -6668 4750 -6640
rect 454 -6680 460 -6668
rect 4744 -6680 4750 -6668
rect 4802 -6680 4808 -6628
rect 866 -6748 872 -6696
rect 924 -6708 930 -6696
rect 5216 -6708 5222 -6696
rect 924 -6736 5222 -6708
rect 924 -6748 930 -6736
rect 5216 -6748 5222 -6736
rect 5286 -6748 5292 -6696
rect 1484 -6816 1490 -6764
rect 1542 -6776 1548 -6764
rect 5832 -6776 5838 -6764
rect 1542 -6804 5838 -6776
rect 1542 -6816 1548 -6804
rect 5832 -6816 5838 -6804
rect 5890 -6816 5896 -6764
rect 1956 -6884 1962 -6832
rect 2014 -6844 2020 -6832
rect 6312 -6844 6318 -6820
rect 2014 -6872 6318 -6844
rect 6370 -6872 6376 -6820
rect 6928 -6872 6934 -6820
rect 6986 -6872 6992 -6820
rect 2014 -6884 2020 -6872
rect 2572 -6952 2578 -6900
rect 2630 -6912 2636 -6900
rect 6932 -6912 6988 -6872
rect 2630 -6940 6988 -6912
rect 2630 -6952 2636 -6940
rect 500 -6982 552 -6976
rect 2689 -6994 2695 -6983
rect 552 -7023 2695 -6994
rect 500 -7040 552 -7034
rect 2689 -7035 2695 -7023
rect 2747 -7035 2753 -6983
rect 3520 -6992 3596 -6982
rect 3238 -6998 3302 -6992
rect 3238 -7050 3244 -6998
rect 3296 -7050 3302 -6998
rect 3238 -7056 3302 -7050
rect 3520 -7048 3530 -6992
rect 3586 -6998 3596 -6992
rect 5948 -6998 5954 -6996
rect 3586 -7046 5954 -6998
rect 3586 -7048 3596 -7046
rect 5948 -7048 5954 -7046
rect 6006 -7048 6012 -6996
rect 3244 -7208 3296 -7056
rect 3520 -7058 3596 -7048
rect -690 -7260 -684 -7208
rect -632 -7260 -216 -7208
rect -164 -7260 404 -7208
rect 456 -7260 872 -7208
rect 924 -7260 1492 -7208
rect 1544 -7260 1962 -7208
rect 2014 -7260 2580 -7208
rect 2632 -7260 3296 -7208
rect 3244 -7318 3296 -7260
rect 3244 -7370 3662 -7318
rect 3714 -7370 4142 -7318
rect 4194 -7370 4750 -7318
rect 4802 -7370 5230 -7318
rect 5282 -7370 5838 -7318
rect 5890 -7370 6318 -7318
rect 6370 -7370 6926 -7318
rect 6978 -7370 6984 -7318
<< via2 >>
rect -1006 -6136 -930 -5918
rect 82 -6136 158 -5918
rect 1170 -6136 1246 -5918
rect 1714 -6136 1790 -5918
rect 2258 -6136 2334 -5918
rect 2802 -6136 2878 -5918
rect 3346 -6136 3422 -5918
rect 3890 -6136 3966 -5918
rect 4434 -6136 4510 -5918
rect 4978 -6136 5054 -5918
rect 5522 -6136 5598 -5918
rect 6066 -6136 6142 -5918
rect 6610 -6136 6686 -5918
rect 7154 -6136 7230 -5918
rect 2490 -6448 2546 -6392
rect 3186 -6488 3246 -6428
rect 3246 -6488 3254 -6428
rect 5120 -6418 5176 -6362
rect 3530 -7048 3586 -6992
<< metal3 >>
rect -1016 -5614 -920 -5608
rect -1016 -5842 -1010 -5614
rect -926 -5842 -920 -5614
rect -1016 -5918 -920 -5842
rect 72 -5614 168 -5608
rect 72 -5842 78 -5614
rect 162 -5842 168 -5614
rect -1016 -6136 -1006 -5918
rect -930 -6136 -920 -5918
rect -1016 -6148 -920 -6136
rect -472 -5914 -376 -5908
rect -472 -6142 -466 -5914
rect -382 -6142 -376 -5914
rect -472 -6148 -376 -6142
rect 72 -5918 168 -5842
rect 1160 -5614 1256 -5608
rect 1160 -5842 1166 -5614
rect 1250 -5842 1256 -5614
rect 72 -6136 82 -5918
rect 158 -6136 168 -5918
rect 72 -6148 168 -6136
rect 616 -5914 712 -5908
rect 616 -6142 622 -5914
rect 706 -6142 712 -5914
rect 616 -6148 712 -6142
rect 1160 -5918 1256 -5842
rect 2248 -5614 2344 -5608
rect 2248 -5842 2254 -5614
rect 2338 -5842 2344 -5614
rect 1160 -6136 1170 -5918
rect 1246 -6136 1256 -5918
rect 1160 -6148 1256 -6136
rect 1704 -5914 1800 -5908
rect 1704 -6142 1710 -5914
rect 1794 -6142 1800 -5914
rect 1704 -6148 1800 -6142
rect 2248 -5918 2344 -5842
rect 3336 -5614 3432 -5608
rect 3336 -5842 3342 -5614
rect 3426 -5842 3432 -5614
rect 2248 -6136 2258 -5918
rect 2334 -6136 2344 -5918
rect 2248 -6148 2344 -6136
rect 2792 -5914 2888 -5908
rect 2792 -6142 2798 -5914
rect 2882 -6142 2888 -5914
rect 2792 -6148 2888 -6142
rect 3336 -5918 3432 -5842
rect 4424 -5614 4520 -5608
rect 4424 -5842 4430 -5614
rect 4514 -5842 4520 -5614
rect 3336 -6136 3346 -5918
rect 3422 -6136 3432 -5918
rect 3336 -6148 3432 -6136
rect 3880 -5914 3976 -5908
rect 3880 -6142 3886 -5914
rect 3970 -6142 3976 -5914
rect 3880 -6148 3976 -6142
rect 4424 -5918 4520 -5842
rect 5512 -5614 5608 -5608
rect 5512 -5842 5518 -5614
rect 5602 -5842 5608 -5614
rect 4424 -6136 4434 -5918
rect 4510 -6136 4520 -5918
rect 4424 -6148 4520 -6136
rect 4968 -5914 5064 -5908
rect 4968 -6142 4974 -5914
rect 5058 -6142 5064 -5914
rect 4968 -6148 5064 -6142
rect 5512 -5918 5608 -5842
rect 6600 -5614 6696 -5608
rect 6600 -5842 6606 -5614
rect 6690 -5842 6696 -5614
rect 5512 -6136 5522 -5918
rect 5598 -6136 5608 -5918
rect 5512 -6148 5608 -6136
rect 6056 -5914 6152 -5908
rect 6056 -6142 6062 -5914
rect 6146 -6142 6152 -5914
rect 6056 -6148 6152 -6142
rect 6600 -5918 6696 -5842
rect 6600 -6136 6610 -5918
rect 6686 -6136 6696 -5918
rect 6600 -6148 6696 -6136
rect 7144 -5914 7240 -5908
rect 7144 -6142 7150 -5914
rect 7234 -6142 7240 -5914
rect 7144 -6148 7240 -6142
rect 5115 -6362 5181 -6357
rect 2485 -6392 2551 -6387
rect 2485 -6448 2490 -6392
rect 2546 -6448 2551 -6392
rect 5115 -6418 5120 -6362
rect 5176 -6418 5181 -6362
rect 2485 -6453 2551 -6448
rect 3160 -6428 3282 -6422
rect 5115 -6423 5181 -6418
rect 2488 -7130 2548 -6453
rect 3160 -6488 3186 -6428
rect 3254 -6434 3282 -6428
rect 3254 -6488 3588 -6434
rect 3160 -6494 3588 -6488
rect 3528 -6987 3588 -6494
rect 3525 -6992 3591 -6987
rect 3525 -7048 3530 -6992
rect 3586 -7048 3591 -6992
rect 3525 -7053 3591 -7048
rect 5118 -7130 5178 -6423
rect 2488 -7190 5178 -7130
<< via3 >>
rect -1010 -5842 -926 -5614
rect 78 -5842 162 -5614
rect -466 -6142 -382 -5914
rect 1166 -5842 1250 -5614
rect 622 -6142 706 -5914
rect 2254 -5842 2338 -5614
rect 1710 -5918 1794 -5914
rect 1710 -6136 1714 -5918
rect 1714 -6136 1790 -5918
rect 1790 -6136 1794 -5918
rect 1710 -6142 1794 -6136
rect 3342 -5842 3426 -5614
rect 2798 -5918 2882 -5914
rect 2798 -6136 2802 -5918
rect 2802 -6136 2878 -5918
rect 2878 -6136 2882 -5918
rect 2798 -6142 2882 -6136
rect 4430 -5842 4514 -5614
rect 3886 -5918 3970 -5914
rect 3886 -6136 3890 -5918
rect 3890 -6136 3966 -5918
rect 3966 -6136 3970 -5918
rect 3886 -6142 3970 -6136
rect 5518 -5842 5602 -5614
rect 4974 -5918 5058 -5914
rect 4974 -6136 4978 -5918
rect 4978 -6136 5054 -5918
rect 5054 -6136 5058 -5918
rect 4974 -6142 5058 -6136
rect 6606 -5842 6690 -5614
rect 6062 -5918 6146 -5914
rect 6062 -6136 6066 -5918
rect 6066 -6136 6142 -5918
rect 6142 -6136 6146 -5918
rect 6062 -6142 6146 -6136
rect 7150 -5918 7234 -5914
rect 7150 -6136 7154 -5918
rect 7154 -6136 7230 -5918
rect 7230 -6136 7234 -5918
rect 7150 -6142 7234 -6136
<< metal4 >>
rect -1016 -5614 7240 -5608
rect -1016 -5842 -1010 -5614
rect -926 -5842 78 -5614
rect 162 -5842 1166 -5614
rect 1250 -5842 2254 -5614
rect 2338 -5842 3342 -5614
rect 3426 -5842 4430 -5614
rect 4514 -5842 5518 -5614
rect 5602 -5842 6606 -5614
rect 6690 -5842 7240 -5614
rect -1016 -5848 7240 -5842
rect -1016 -5914 7240 -5908
rect -1016 -6142 -466 -5914
rect -382 -6142 622 -5914
rect 706 -6142 1710 -5914
rect 1794 -6142 2798 -5914
rect 2882 -6142 3886 -5914
rect 3970 -6142 4974 -5914
rect 5058 -6142 6062 -5914
rect 6146 -6142 7150 -5914
rect 7234 -6142 7240 -5914
rect -1016 -6148 7240 -6142
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 1 2840 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_1
timestamp 1757695336
transform 0 -1 3928 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_2
timestamp 1757695336
transform 0 1 3928 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_3
timestamp 1757695336
transform 0 -1 5016 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_4
timestamp 1757695336
transform 0 1 5016 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_5
timestamp 1757695336
transform 0 -1 6104 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_6
timestamp 1757695336
transform 0 1 6104 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_7
timestamp 1757695336
transform 0 -1 7192 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn0
timestamp 1757695336
transform 0 -1 -424 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn1
timestamp 1757695336
transform 0 1 -424 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn2
timestamp 1757695336
transform 0 -1 664 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn3
timestamp 1757695336
transform 0 1 664 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn4
timestamp 1757695336
transform 0 -1 1752 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn5
timestamp 1757695336
transform 0 1 1752 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_oTn6
timestamp 1757695336
transform 0 -1 2840 -1 0 -6472
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  XOTn0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 -1 -424 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn1
timestamp 1757695336
transform 0 1 -424 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn2
timestamp 1757695336
transform 0 -1 664 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn3
timestamp 1757695336
transform 0 1 664 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn4
timestamp 1757695336
transform 0 -1 1752 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn5
timestamp 1757695336
transform 0 1 1752 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  XOTn6
timestamp 1757695336
transform 0 -1 2840 -1 0 -6564
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  XOTn7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 1 2840 -1 0 -6564
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  XOTn8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 -1 3928 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn9
timestamp 1757695336
transform 0 1 3928 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn10
timestamp 1757695336
transform 0 -1 5016 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn11
timestamp 1757695336
transform 0 1 5016 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn12
timestamp 1757695336
transform 0 -1 6104 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn13
timestamp 1757695336
transform 0 1 6104 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  XOTn14
timestamp 1757695336
transform 0 -1 7192 1 0 -7392
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  XTA1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 -1 3928 -1 0 -6196
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTA2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 1 3928 -1 0 -6196
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTA3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 -1 5016 -1 0 -6196
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTAN
timestamp 1757695336
transform 0 1 5016 -1 0 -6196
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTAN2
timestamp 1757695336
transform 0 -1 6104 -1 0 -6196
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB1
timestamp 1757695336
transform 0 -1 -424 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB2
timestamp 1757695336
transform 0 1 -424 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  XTB3
timestamp 1757695336
transform 0 -1 664 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  XTB4
timestamp 1757695336
transform 0 1 664 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB5
timestamp 1757695336
transform 0 -1 1752 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB6
timestamp 1757695336
transform 0 1 1752 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  XTB7
timestamp 1757695336
transform 0 -1 2840 1 0 -6472
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  XTBN $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1757695336
transform 0 1 2840 -1 0 -6196
box -38 -48 314 592
<< labels >>
flabel metal4 -1016 -6148 7240 -5908 0 FreeSans 1600 0 0 0 VGND
port 91 nsew
flabel metal4 -1016 -5848 7240 -5608 0 FreeSans 1600 0 0 0 VPWR
port 90 nsew
flabel metal1 5848 -5550 5888 -5510 0 FreeSans 80 90 0 0 d[3]
port 1104 nsew
flabel metal1 5238 -5550 5278 -5510 0 FreeSans 80 90 0 0 d[2]
port 1103 nsew
flabel metal1 3672 -5550 3712 -5510 0 FreeSans 80 90 0 0 d[1]
port 1102 nsew
flabel metal1 3590 -5550 3630 -5510 0 FreeSans 80 90 0 0 d[0]
port 1101 nsew
flabel metal1 -778 -7430 -564 -7386 0 FreeSans 160 0 0 0 Tn[0]
port 1900 nsew
flabel metal1 -284 -7430 -70 -7386 0 FreeSans 160 0 0 0 Tn[1]
port 1901 nsew
flabel metal1 310 -7430 524 -7386 0 FreeSans 160 0 0 0 Tn[2]
port 1902 nsew
flabel metal1 804 -7430 1018 -7386 0 FreeSans 160 0 0 0 Tn[3]
port 1903 nsew
flabel metal1 1398 -7430 1612 -7386 0 FreeSans 160 0 0 0 Tn[4]
port 1904 nsew
flabel metal1 1892 -7430 2106 -7386 0 FreeSans 160 0 0 0 Tn[5]
port 1905 nsew
flabel metal1 2486 -7430 2700 -7386 0 FreeSans 160 0 0 0 Tn[6]
port 1906 nsew
flabel metal1 2984 -7430 3196 -7386 0 FreeSans 160 0 0 0 Tn[7]
port 1907 nsew
flabel metal1 3498 -7430 3628 -7386 0 FreeSans 160 0 0 0 Tn[8]
port 1908 nsew
flabel metal1 4228 -7430 4358 -7386 0 FreeSans 160 0 0 0 Tn[9]
port 1909 nsew
flabel metal1 4586 -7430 4716 -7386 0 FreeSans 160 0 0 0 Tn[10]
port 1910 nsew
flabel metal1 5316 -7430 5446 -7386 0 FreeSans 160 0 0 0 Tn[11]
port 1911 nsew
flabel metal1 5674 -7430 5804 -7386 0 FreeSans 160 0 0 0 Tn[12]
port 1912 nsew
flabel metal1 6404 -7430 6534 -7386 0 FreeSans 160 0 0 0 Tn[13]
port 1913 nsew
flabel metal1 6762 -7430 6892 -7386 0 FreeSans 160 0 0 0 Tn[14]
port 1914 nsew
<< end >>
