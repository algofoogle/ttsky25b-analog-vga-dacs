* NGSPICE file created from csdac255_parax.ext - technology: sky130A

.subckt csdac255_parax Iout VPWR VGND Vbias data[0] data[1] data[2] data[3] data[4]
+ data[5] data[6] data[7] bias[0] bias[1] bias[2]
X0 XA.XIR[2].XIC_dummy_right.icell.SM XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout VGND.t1876 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1 VPWR.t1096 XThR.Tn[2].t12 XA.XIR[3].XIC[8].icell.PUM VPWR.t1095 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2 XA.XIR[12].XIC[10].icell.SM XA.XIR[12].XIC[10].icell.Ien Iout.t236 VGND.t2534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X3 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1794 VPWR.t1796 VPWR.t1795 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X4 VGND.t510 XThC.Tn[10].t12 XA.XIR[4].XIC[10].icell.PDM VGND.t509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X5 VGND.t669 XThR.XTBN.Y.t4 a_n997_2667# VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VPWR.t453 XThR.Tn[6].t12 XA.XIR[7].XIC[8].icell.PUM VPWR.t452 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X7 XA.XIR[14].XIC[5].icell.Ien XThR.Tn[14].t12 VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X8 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[12].t12 XA.XIR[12].XIC[6].icell.Ien VGND.t1792 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X9 XThC.Tn[6].t11 XThC.XTBN.Y.t4 VGND.t2275 VGND.t2274 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1931 VGND.t682 VGND.t681 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X11 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[9].t12 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X12 VGND.t2276 XThC.XTBN.Y.t5 XThC.Tn[5].t7 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 XA.XIR[15].XIC[9].icell.PUM XThC.Tn[9].t12 XA.XIR[15].XIC[9].icell.Ien VPWR.t804 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X14 XA.XIR[9].XIC[0].icell.SM XA.XIR[9].XIC[0].icell.Ien Iout.t245 VGND.t2607 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X15 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[12].t13 VGND.t1794 VGND.t1793 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X16 VGND.t655 XThC.Tn[11].t12 XA.XIR[12].XIC[11].icell.PDM VGND.t654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X17 XA.XIR[12].XIC[1].icell.SM XA.XIR[12].XIC[1].icell.Ien Iout.t221 VGND.t2206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X18 XA.XIR[8].XIC[12].icell.SM XA.XIR[8].XIC[12].icell.Ien Iout.t106 VGND.t1154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X19 XThC.Tn[12].t7 XThC.XTB5.Y VPWR.t167 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 XA.XIR[8].XIC_15.icell.PDM VPWR.t1932 VGND.t684 VGND.t683 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X21 XA.XIR[7].XIC[13].icell.SM XA.XIR[7].XIC[13].icell.Ien Iout.t223 VGND.t2295 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X22 XA.XIR[14].XIC[13].icell.PUM XThC.Tn[13].t12 XA.XIR[14].XIC[13].icell.Ien VPWR.t170 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X23 a_2979_9615# XThC.XTBN.Y.t6 XThC.Tn[0].t6 VPWR.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1792 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1793 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X25 XA.XIR[10].XIC[14].icell.SM XA.XIR[10].XIC[14].icell.Ien Iout.t51 VGND.t523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X26 a_4861_9615# XThC.XTB4.Y.t2 VPWR.t208 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_5949_9615# XThC.XTBN.Y.t7 XThC.Tn[5].t11 VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[6].t13 XA.XIR[6].XIC[10].icell.Ien VGND.t662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X29 XA.XIR[0].XIC[4].icell.PDM VGND.t1028 VGND.t1030 VGND.t1029 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X30 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[3].t12 VGND.t1193 VGND.t1192 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X31 XThR.Tn[5].t7 XThR.XTBN.Y.t5 a_n1049_5611# VPWR.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X32 XThC.Tn[4].t3 XThC.XTB5.Y VGND.t291 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X33 VGND.t2277 XThC.XTBN.Y.t8 XThC.Tn[2].t11 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X34 XThR.XTB2.Y XThR.XTB6.A VPWR.t964 VPWR.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X35 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[6].t14 VGND.t664 VGND.t663 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X36 XA.XIR[6].XIC[11].icell.SM XA.XIR[6].XIC[11].icell.Ien Iout.t25 VGND.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X37 VGND.t2000 XThC.Tn[2].t12 XA.XIR[12].XIC[2].icell.PDM VGND.t1999 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X38 VPWR.t1791 VPWR.t1789 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1790 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X39 VGND.t686 VPWR.t1933 XA.XIR[7].XIC_dummy_left.icell.PDM VGND.t685 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X40 VPWR.t686 XThR.Tn[3].t13 XA.XIR[4].XIC[11].icell.PUM VPWR.t685 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X41 VGND.t1201 Vbias.t12 XA.XIR[14].XIC[11].icell.SM VGND.t1200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X42 XA.XIR[2].XIC[1].icell.PUM XThC.Tn[1].t12 XA.XIR[2].XIC[1].icell.Ien VPWR.t883 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X43 VGND.t2558 XThC.Tn[3].t12 XA.XIR[15].XIC[3].icell.PDM VGND.t2557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X44 VGND.t688 VPWR.t1934 XA.XIR[10].XIC_15.icell.PDM VGND.t687 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X45 VPWR.t533 XThR.Tn[10].t12 XA.XIR[11].XIC[9].icell.PUM VPWR.t532 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X46 XA.XIR[0].XIC[14].icell.PUM XThC.Tn[14].t12 XA.XIR[0].XIC[14].icell.Ien VPWR.t1292 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X47 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1786 VPWR.t1788 VPWR.t1787 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X48 a_7651_9569# XThC.XTB1.Y.t3 XThC.Tn[8].t3 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X49 VGND.t1878 Vbias.t13 XA.XIR[2].XIC[5].icell.SM VGND.t1877 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X50 XA.XIR[1].XIC[6].icell.Ien XThR.Tn[1].t12 VPWR.t910 VPWR.t909 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X51 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t3 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 VGND.t2250 XThC.Tn[4].t12 XA.XIR[2].XIC[4].icell.PDM VGND.t2249 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X53 XThC.XTB5.Y XThC.XTB7.B VGND.t1336 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X54 XThC.Tn[7].t7 XThC.XTBN.Y.t9 VPWR.t1348 VPWR.t1347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X55 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[9].t13 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X56 VGND.t1752 XThR.XTB7.Y XThR.Tn[6].t11 VGND.t1751 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X57 XA.XIR[4].XIC[7].icell.Ien XThR.Tn[4].t12 VPWR.t1179 VPWR.t1178 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X58 VPWR.t465 XThR.XTBN.Y.t6 XThR.Tn[9].t3 VPWR.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X59 XThR.XTB7.Y XThR.XTB7.A VGND.t2647 VGND.t2646 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X60 XA.XIR[3].XIC[8].icell.Ien XThR.Tn[3].t14 VPWR.t688 VPWR.t687 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X61 VPWR.t690 XThR.Tn[3].t15 XA.XIR[4].XIC[2].icell.PUM VPWR.t689 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X62 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[12].t14 VGND.t1796 VGND.t1795 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X63 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[1].t13 XA.XIR[1].XIC[9].icell.Ien VGND.t1605 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X64 VPWR.t1094 XThR.Tn[2].t13 XA.XIR[3].XIC[3].icell.PUM VPWR.t1093 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X65 XA.XIR[5].XIC_dummy_left.icell.SM XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout VGND.t869 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X66 VPWR.t455 XThR.Tn[6].t15 XA.XIR[7].XIC[3].icell.PUM VPWR.t454 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X67 VPWR.t1785 VPWR.t1783 XA.XIR[2].XIC_15.icell.PUM VPWR.t1784 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X68 a_6243_9615# XThC.XTB7.Y VPWR.t119 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X69 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[11].t12 XA.XIR[11].XIC[14].icell.Ien VGND.t1973 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X70 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[11].t13 XA.XIR[11].XIC[8].icell.Ien VGND.t1974 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X71 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[3].t16 VGND.t1195 VGND.t1194 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X72 XThR.Tn[7].t7 XThR.XTBN.Y.t7 VPWR.t467 VPWR.t466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X73 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[0].t12 VGND.t1122 VGND.t1121 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X74 a_8963_9569# XThC.XTBN.Y.t10 VGND.t2278 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X75 VGND.t1880 Vbias.t14 XA.XIR[12].XIC[7].icell.SM VGND.t1879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X76 VGND.t653 XThC.Tn[6].t12 XA.XIR[12].XIC[6].icell.PDM VGND.t652 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X77 XA.XIR[6].XIC[9].icell.SM XA.XIR[6].XIC[9].icell.Ien Iout.t162 VGND.t1590 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X78 XA.XIR[2].XIC_dummy_left.icell.SM XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout VGND.t1403 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X79 XA.XIR[3].XIC[11].icell.SM XA.XIR[3].XIC[11].icell.Ien Iout.t113 VGND.t1279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X80 VGND.t690 VPWR.t1935 XA.XIR[4].XIC_dummy_left.icell.PDM VGND.t689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X81 VGND.t670 XThR.XTBN.Y.t8 XThR.Tn[5].t11 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X82 VGND.t1882 Vbias.t15 XA.XIR[15].XIC[8].icell.SM VGND.t1881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X83 VGND.t1884 Vbias.t16 XA.XIR[14].XIC[9].icell.SM VGND.t1883 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X84 VGND.t2134 XThC.Tn[7].t8 XA.XIR[15].XIC[7].icell.PDM VGND.t2133 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X85 VGND.t657 XThC.Tn[11].t13 XA.XIR[6].XIC[11].icell.PDM VGND.t656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X86 VGND.t1593 XThC.Tn[1].t13 XA.XIR[3].XIC[1].icell.PDM VGND.t1592 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X87 XA.XIR[4].XIC[11].icell.Ien XThR.Tn[4].t13 VPWR.t1181 VPWR.t1180 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X88 VPWR.t135 XThR.XTB6.Y a_n1049_5611# VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X89 XA.XIR[14].XIC[6].icell.PUM XThC.Tn[6].t13 XA.XIR[14].XIC[6].icell.Ien VPWR.t431 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X90 VGND.t1886 Vbias.t17 XA.XIR[9].XIC[7].icell.SM VGND.t1885 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X91 VGND.t2002 XThC.Tn[2].t13 XA.XIR[6].XIC[2].icell.PDM VGND.t2001 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X92 XA.XIR[11].XIC[9].icell.Ien XThR.Tn[11].t14 VPWR.t1162 VPWR.t1161 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X93 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t1936 XA.XIR[6].XIC_dummy_left.icell.Ien VGND.t691 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X94 a_n1049_7787# XThR.XTB2.Y VPWR.t1177 VPWR.t1176 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X95 VGND.t1467 XThC.Tn[9].t13 XA.XIR[14].XIC[9].icell.PDM VGND.t1466 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X96 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[8].t12 XA.XIR[8].XIC[11].icell.Ien VGND.t1460 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X97 VGND.t1888 Vbias.t18 XA.XIR[2].XIC[0].icell.SM VGND.t1887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X98 XA.XIR[1].XIC[1].icell.Ien XThR.Tn[1].t14 VPWR.t1335 VPWR.t1334 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X99 XA.XIR[13].XIC[4].icell.PUM XThC.Tn[4].t13 XA.XIR[13].XIC[4].icell.Ien VPWR.t1329 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X100 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1781 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1782 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X101 VGND.t1890 Vbias.t19 XA.XIR[0].XIC[13].icell.SM VGND.t1889 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X102 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[0].t13 VGND.t1124 VGND.t1123 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X103 XA.XIR[4].XIC[2].icell.Ien XThR.Tn[4].t14 VPWR.t1183 VPWR.t1182 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X104 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[8].t13 VGND.t1462 VGND.t1461 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X105 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[8].t14 VGND.t1464 VGND.t1463 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X106 XA.XIR[3].XIC[3].icell.Ien XThR.Tn[3].t17 VPWR.t692 VPWR.t691 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X107 VGND.t2670 XThC.Tn[12].t12 XA.XIR[0].XIC[12].icell.PDM VGND.t2669 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X108 VPWR.t29 XThC.XTB3.Y.t3 a_4067_9615# VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X109 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[1].t15 XA.XIR[1].XIC[4].icell.Ien VGND.t2255 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X110 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[5].t12 XA.XIR[5].XIC[1].icell.Ien VGND.t124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X111 VPWR.t99 data[4].t0 a_n1335_4229# VPWR.t98 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X112 XA.XIR[2].XIC_15.icell.Ien XThR.Tn[2].t14 VPWR.t1092 VPWR.t1091 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X113 XA.XIR[3].XIC[9].icell.SM XA.XIR[3].XIC[9].icell.Ien Iout.t181 VGND.t1705 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X114 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[9].t14 XA.XIR[9].XIC[1].icell.Ien VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X115 VGND.t672 XThR.XTBN.Y.t9 XThR.Tn[7].t3 VGND.t671 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X116 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[4].t15 XA.XIR[4].XIC[5].icell.Ien VGND.t1989 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X117 a_n1319_5317# XThR.XTB7.A VPWR.t1890 VPWR.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X118 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[8].t15 XA.XIR[8].XIC[2].icell.Ien VGND.t1155 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X119 VPWR.t635 XThR.Tn[13].t12 XA.XIR[14].XIC[14].icell.PUM VPWR.t634 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X120 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[11].t15 XA.XIR[11].XIC[3].icell.Ien VGND.t1975 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X121 XA.XIR[7].XIC[8].icell.PUM XThC.Tn[8].t12 XA.XIR[7].XIC[8].icell.Ien VPWR.t1149 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X122 XThC.Tn[9].t3 XThC.XTB2.Y VPWR.t109 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X123 XA.XIR[15].XIC[4].icell.Ien VPWR.t1778 VPWR.t1780 VPWR.t1779 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X124 VGND.t1892 Vbias.t20 XA.XIR[12].XIC[2].icell.SM VGND.t1891 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X125 XA.XIR[6].XIC[4].icell.SM XA.XIR[6].XIC[4].icell.Ien Iout.t229 VGND.t2506 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X126 VGND.t1894 Vbias.t21 XA.XIR[11].XIC_15.icell.SM VGND.t1893 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X127 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1775 VPWR.t1777 VPWR.t1776 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X128 XThC.Tn[5].t6 XThC.XTBN.Y.t11 VGND.t2279 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X129 XA.XIR[1].XIC_dummy_right.icell.SM XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout VGND.t1516 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X130 VGND.t1896 Vbias.t22 XA.XIR[15].XIC[3].icell.SM VGND.t1895 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X131 VGND.t1898 Vbias.t23 XA.XIR[14].XIC[4].icell.SM VGND.t1897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X132 VGND.t626 XThC.Tn[6].t14 XA.XIR[6].XIC[6].icell.PDM VGND.t625 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X133 VPWR.t666 XThR.Tn[8].t16 XA.XIR[9].XIC[4].icell.PUM VPWR.t665 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X134 VPWR.t973 XThR.Tn[12].t15 XA.XIR[13].XIC[12].icell.PUM VPWR.t972 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X135 VGND.t1027 VGND.t1025 XA.XIR[13].XIC_dummy_right.icell.SM VGND.t1026 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X136 XThR.Tn[9].t7 XThR.XTB2.Y a_n997_3755# VGND.t1554 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X137 XThC.Tn[0].t5 XThC.XTBN.Y.t12 a_2979_9615# VPWR.t1366 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X138 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t1937 VGND.t693 VGND.t692 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X139 XThC.Tn[5].t10 XThC.XTBN.Y.t13 a_5949_9615# VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X140 VGND.t290 XThC.XTB5.Y XThC.Tn[4].t2 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X141 XA.XIR[14].XIC[1].icell.PUM XThC.Tn[1].t14 XA.XIR[14].XIC[1].icell.Ien VPWR.t884 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X142 VGND.t1900 Vbias.t24 XA.XIR[9].XIC[2].icell.SM VGND.t1899 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X143 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t3 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X144 XA.XIR[13].XIC[0].icell.PUM XThC.Tn[0].t12 XA.XIR[13].XIC[0].icell.Ien VPWR.t741 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X145 XThC.Tn[7].t3 XThC.XTBN.Y.t14 VGND.t2359 VGND.t2358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X146 XThC.Tn[2].t10 XThC.XTBN.Y.t15 VGND.t2360 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X147 VGND.t512 XThC.Tn[10].t13 XA.XIR[0].XIC[10].icell.PDM VGND.t511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X148 a_n997_1579# XThR.XTBN.Y.t10 VGND.t1253 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X149 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[5].t13 VGND.t133 VGND.t132 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X150 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[5].t14 VGND.t135 VGND.t134 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X151 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR.t1773 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X152 XA.XIR[9].XIC[14].icell.SM XA.XIR[9].XIC[14].icell.Ien Iout.t36 VGND.t251 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X153 VGND.t2252 XThC.Tn[4].t14 XA.XIR[14].XIC[4].icell.PDM VGND.t2251 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X154 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[8].t17 XA.XIR[8].XIC[6].icell.Ien VGND.t1156 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X155 XA.XIR[1].XIC[7].icell.PUM XThC.Tn[7].t9 XA.XIR[1].XIC[7].icell.Ien VPWR.t1257 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X156 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[6].t16 VGND.t666 VGND.t665 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X157 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[1].t16 VGND.t2257 VGND.t2256 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X158 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[11].t16 XA.XIR[11].XIC[7].icell.Ien VGND.t1976 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X159 XA.XIR[4].XIC[8].icell.PUM XThC.Tn[8].t13 XA.XIR[4].XIC[8].icell.Ien VPWR.t1150 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X160 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[8].t18 VGND.t1158 VGND.t1157 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X161 XA.XIR[0].XIC_15.icell.SM XA.XIR[0].XIC_15.icell.Ien Iout.t180 VGND.t1704 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X162 XA.XIR[4].XIC[12].icell.SM XA.XIR[4].XIC[12].icell.Ien Iout.t174 VGND.t1636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X163 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[13].t13 VGND.t1110 VGND.t1109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X164 XA.XIR[11].XIC[12].icell.PUM XThC.Tn[12].t13 XA.XIR[11].XIC[12].icell.Ien VPWR.t1913 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X165 XA.XIR[12].XIC[4].icell.Ien XThR.Tn[12].t16 VPWR.t975 VPWR.t974 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X166 XA.XIR[3].XIC[4].icell.SM XA.XIR[3].XIC[4].icell.Ien Iout.t77 VGND.t871 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X167 XA.XIR[15].XIC[0].icell.Ien VPWR.t1770 VPWR.t1772 VPWR.t1771 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X168 VGND.t776 Vbias.t25 XA.XIR[8].XIC_15.icell.SM VGND.t775 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X169 VGND.t2180 XThC.Tn[14].t13 XA.XIR[8].XIC[14].icell.PDM VGND.t2179 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X170 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1767 VPWR.t1769 VPWR.t1768 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X171 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[4].t16 XA.XIR[4].XIC[0].icell.Ien VGND.t1990 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X172 VGND.t2156 XThC.Tn[8].t14 XA.XIR[8].XIC[8].icell.PDM VGND.t2155 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X173 XA.XIR[14].XIC[14].icell.Ien XThR.Tn[14].t13 VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X174 VGND.t2361 XThC.XTBN.Y.t16 XThC.Tn[1].t7 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X175 VGND.t778 Vbias.t26 XA.XIR[1].XIC[5].icell.SM VGND.t777 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X176 VPWR.t977 XThR.Tn[12].t17 XA.XIR[13].XIC[10].icell.PUM VPWR.t976 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X177 XA.XIR[7].XIC[3].icell.PUM XThC.Tn[3].t13 XA.XIR[7].XIC[3].icell.Ien VPWR.t1837 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X178 XA.XIR[2].XIC_15.icell.PUM VPWR.t1765 XA.XIR[2].XIC_15.icell.Ien VPWR.t1766 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X179 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[2].t15 XA.XIR[2].XIC[13].icell.Ien VGND.t811 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X180 VPWR.t1 XThR.Tn[9].t15 XA.XIR[10].XIC[12].icell.PUM VPWR.t0 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X181 VPWR.t668 XThR.Tn[8].t19 XA.XIR[9].XIC[0].icell.PUM VPWR.t667 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X182 VGND.t780 Vbias.t27 XA.XIR[4].XIC[6].icell.SM VGND.t779 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X183 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1938 VGND.t695 VGND.t694 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X184 VPWR.t1764 VPWR.t1762 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1763 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X185 VPWR.t1367 XThC.XTBN.Y.t17 XThC.Tn[10].t11 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VGND.t1254 XThR.XTBN.Y.t11 XThR.Tn[3].t7 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[2].t16 VGND.t99 VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X188 XA.XIR[6].XIC[8].icell.Ien XThR.Tn[6].t17 VPWR.t457 VPWR.t456 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X189 XThR.Tn[0].t4 XThR.XTBN.Y.t12 a_n1049_8581# VPWR.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X190 XA.XIR[13].XIC[12].icell.Ien XThR.Tn[13].t14 VPWR.t637 VPWR.t636 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X191 XA.XIR[13].XIC[7].icell.SM XA.XIR[13].XIC[7].icell.Ien Iout.t48 VGND.t421 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X192 VPWR.t598 VGND.t2689 XA.XIR[0].XIC[8].icell.PUM VPWR.t597 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X193 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[10].t13 XA.XIR[10].XIC[14].icell.Ien VGND.t2526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X194 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[10].t14 XA.XIR[10].XIC[8].icell.Ien VGND.t2527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X195 XThC.Tn[12].t6 XThC.XTB5.Y VPWR.t166 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X196 XA.XIR[1].XIC[11].icell.PUM XThC.Tn[11].t14 XA.XIR[1].XIC[11].icell.Ien VPWR.t451 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X197 XThR.Tn[11].t11 XThR.XTBN.Y.t13 VPWR.t694 VPWR.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 XA.XIR[0].XIC[7].icell.Ien XThR.Tn[0].t14 VPWR.t649 VPWR.t648 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X199 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[2].t17 VGND.t97 VGND.t96 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X200 XA.XIR[8].XIC[9].icell.PUM XThC.Tn[9].t14 XA.XIR[8].XIC[9].icell.Ien VPWR.t805 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X201 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[8].t20 VGND.t1160 VGND.t1159 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X202 XA.XIR[1].XIC_dummy_left.icell.SM XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout VGND.t1957 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X203 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[5].t15 VGND.t137 VGND.t136 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X204 VGND.t659 XThC.Tn[11].t15 XA.XIR[5].XIC[11].icell.PDM VGND.t658 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X205 XA.XIR[11].XIC[10].icell.PUM XThC.Tn[10].t14 XA.XIR[11].XIC[10].icell.Ien VPWR.t321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X206 XThR.Tn[2].t8 XThR.XTBN.Y.t14 VGND.t1255 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X207 VGND.t661 XThC.Tn[11].t16 XA.XIR[9].XIC[11].icell.PDM VGND.t660 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X208 VGND.t1024 VGND.t1022 XA.XIR[13].XIC_dummy_left.icell.SM VGND.t1023 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X209 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12].t18 VPWR.t178 VPWR.t177 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X210 XA.XIR[1].XIC[2].icell.PUM XThC.Tn[2].t14 XA.XIR[1].XIC[2].icell.Ien VPWR.t1190 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X211 VPWR.t695 XThR.XTBN.Y.t15 XThR.Tn[12].t3 VPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X212 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[1].t17 VGND.t2259 VGND.t2258 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X213 XThC.XTB7.A data[0].t0 VPWR.t605 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X214 VPWR.t3 XThR.Tn[9].t16 XA.XIR[10].XIC[10].icell.PUM VPWR.t2 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X215 XA.XIR[4].XIC[3].icell.PUM XThC.Tn[3].t14 XA.XIR[4].XIC[3].icell.Ien VPWR.t1838 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X216 VGND.t782 Vbias.t28 XA.XIR[4].XIC[10].icell.SM VGND.t781 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X217 XA.XIR[0].XIC[13].icell.PDM VGND.t1019 VGND.t1021 VGND.t1020 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X218 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[13].t15 VGND.t1112 VGND.t1111 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X219 VGND.t697 VPWR.t1939 XA.XIR[0].XIC_dummy_left.icell.PDM VGND.t696 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X220 VGND.t2004 XThC.Tn[2].t15 XA.XIR[5].XIC[2].icell.PDM VGND.t2003 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X221 VGND.t784 Vbias.t29 XA.XIR[11].XIC[8].icell.SM VGND.t783 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X222 XThC.Tn[9].t7 XThC.XTB2.Y a_7875_9569# VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 VGND.t1569 XThC.Tn[5].t12 XA.XIR[1].XIC[5].icell.PDM VGND.t1568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X224 XA.XIR[10].XIC[9].icell.Ien XThR.Tn[10].t15 VPWR.t1408 VPWR.t1407 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X225 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1940 VGND.t699 VGND.t698 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X226 VGND.t1624 XThC.Tn[2].t16 XA.XIR[9].XIC[2].icell.PDM VGND.t1623 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X227 VGND.t2560 XThC.Tn[3].t15 XA.XIR[8].XIC[3].icell.PDM VGND.t2559 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X228 VGND.t701 VPWR.t1941 XA.XIR[3].XIC_15.icell.PDM VGND.t700 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X229 a_n1319_5611# XThR.XTB6.A VPWR.t962 VPWR.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X230 XA.XIR[13].XIC[10].icell.Ien XThR.Tn[13].t16 VPWR.t639 VPWR.t638 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X231 VGND.t1257 XThR.XTBN.Y.t16 a_n997_3979# VGND.t1256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X232 XA.XIR[15].XIC_15.icell.SM XA.XIR[15].XIC_15.icell.Ien Iout.t100 VGND.t1140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X233 VPWR.t1368 XThC.XTBN.Y.t18 XThC.Tn[14].t11 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 VGND.t786 Vbias.t30 XA.XIR[1].XIC[0].icell.SM VGND.t785 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X235 VPWR.t180 XThR.Tn[12].t19 XA.XIR[13].XIC[5].icell.PUM VPWR.t179 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X236 XA.XIR[12].XIC[4].icell.PUM XThC.Tn[4].t15 XA.XIR[12].XIC[4].icell.Ien VPWR.t1330 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X237 VGND.t788 Vbias.t31 XA.XIR[4].XIC[1].icell.SM VGND.t787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X238 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[7].t8 XA.XIR[7].XIC[14].icell.Ien VGND.t860 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X239 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[7].t9 XA.XIR[7].XIC[8].icell.Ien VGND.t861 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X240 XA.XIR[0].XIC[11].icell.Ien XThR.Tn[0].t15 VPWR.t836 VPWR.t835 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X241 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[2].t18 VGND.t95 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X242 XA.XIR[6].XIC[3].icell.Ien XThR.Tn[6].t18 VPWR.t459 VPWR.t458 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X243 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[14].t14 XA.XIR[14].XIC[12].icell.Ien VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X244 XA.XIR[11].XIC[6].icell.SM XA.XIR[11].XIC[6].icell.Ien Iout.t168 VGND.t1617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X245 XA.XIR[1].XIC_15.icell.Ien XThR.Tn[1].t18 VPWR.t1337 VPWR.t1336 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X246 VGND.t790 Vbias.t32 XA.XIR[2].XIC[14].icell.SM VGND.t789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X247 VGND.t298 XThC.Tn[13].t13 XA.XIR[2].XIC[13].icell.PDM VGND.t297 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X248 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[5].t16 VGND.t139 VGND.t138 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X249 VPWR.t91 XThR.XTB4.Y a_n1049_6699# VPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X250 VGND.t703 VPWR.t1942 XA.XIR[15].XIC_dummy_right.icell.PDM VGND.t702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X251 XA.XIR[13].XIC[2].icell.SM XA.XIR[13].XIC[2].icell.Ien Iout.t104 VGND.t1152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X252 VPWR.t596 VGND.t2690 XA.XIR[0].XIC[3].icell.PUM VPWR.t595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X253 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[10].t16 XA.XIR[10].XIC[3].icell.Ien VGND.t2528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X254 VPWR.t769 XThC.XTB6.Y a_5949_9615# VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VPWR.t176 XThR.XTB1.Y.t3 a_n1049_8581# VPWR.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X256 XA.XIR[5].XIC_15.icell.PDM XThR.Tn[5].t17 XA.XIR[5].XIC_15.icell.Ien VGND.t140 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X257 VPWR.t1164 XThR.Tn[11].t17 XA.XIR[12].XIC[7].icell.PUM VPWR.t1163 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X258 XA.XIR[0].XIC[2].icell.Ien XThR.Tn[0].t16 VPWR.t838 VPWR.t837 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X259 XA.XIR[9].XIC_15.icell.PDM XThR.Tn[9].t17 XA.XIR[9].XIC_15.icell.Ien VGND.t33 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X260 XA.XIR[0].XIC[8].icell.SM XA.XIR[0].XIC[8].icell.Ien Iout.t70 VGND.t830 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X261 VGND.t792 Vbias.t33 XA.XIR[5].XIC[7].icell.SM VGND.t791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X262 XA.XIR[11].XIC[5].icell.PUM XThC.Tn[5].t13 XA.XIR[11].XIC[5].icell.Ien VPWR.t866 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X263 VGND.t628 XThC.Tn[6].t15 XA.XIR[5].XIC[6].icell.PDM VGND.t627 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X264 VGND.t1589 XThR.XTB7.B a_n1335_8107# VGND.t1583 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X265 VPWR.t542 XThR.Tn[7].t10 XA.XIR[8].XIC[4].icell.PUM VPWR.t541 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X266 XA.XIR[0].XIC[5].icell.PDM XThR.Tn[0].t17 XA.XIR[0].XIC[5].icell.Ien VGND.t1526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X267 VPWR.t1761 VPWR.t1759 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1760 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X268 VGND.t630 XThC.Tn[6].t16 XA.XIR[9].XIC[6].icell.PDM VGND.t629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X269 VGND.t794 Vbias.t34 XA.XIR[8].XIC[8].icell.SM VGND.t793 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X270 XA.XIR[7].XIC[9].icell.Ien XThR.Tn[7].t11 VPWR.t544 VPWR.t543 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X271 XThC.XTB4.Y.t1 XThC.XTB7.B VPWR.t730 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X272 VGND.t1018 VGND.t1016 XA.XIR[12].XIC_dummy_right.icell.SM VGND.t1017 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X273 VGND.t2136 XThC.Tn[7].t10 XA.XIR[8].XIC[7].icell.PDM VGND.t2135 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X274 VPWR.t1753 VPWR.t1751 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1752 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X275 XThR.Tn[2].t9 XThR.XTB3.Y.t3 VGND.t1641 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X276 VGND.t1258 XThR.XTBN.Y.t17 a_n997_2891# VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X277 VPWR.t323 XThR.Tn[9].t18 XA.XIR[10].XIC[5].icell.PUM VPWR.t322 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X278 XA.XIR[5].XIC[5].icell.SM XA.XIR[5].XIC[5].icell.Ien Iout.t37 VGND.t252 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X279 VPWR.t1898 XThR.XTB5.Y XThR.Tn[12].t11 VPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 XA.XIR[12].XIC[0].icell.PUM XThC.Tn[0].t13 XA.XIR[12].XIC[0].icell.Ien VPWR.t742 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X281 VGND.t1377 XThC.Tn[0].t14 XA.XIR[1].XIC[0].icell.PDM VGND.t1376 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X282 VGND.t796 Vbias.t35 XA.XIR[11].XIC[3].icell.SM VGND.t795 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X283 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[14].t15 XA.XIR[14].XIC[10].icell.Ien VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X284 XA.XIR[11].XIC[10].icell.SM XA.XIR[11].XIC[10].icell.Ien Iout.t135 VGND.t1402 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X285 VGND.t1260 XThR.XTBN.Y.t18 XThR.Tn[6].t7 VGND.t1259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X286 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[11].t18 VGND.t2547 VGND.t2546 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X287 VPWR.t696 XThR.XTBN.Y.t19 XThR.Tn[9].t2 VPWR.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 XA.XIR[8].XIC[6].icell.SM XA.XIR[8].XIC[6].icell.Ien Iout.t137 VGND.t1429 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X289 XA.XIR[13].XIC[5].icell.Ien XThR.Tn[13].t17 VPWR.t641 VPWR.t640 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X290 VGND.t1015 VGND.t1013 XA.XIR[9].XIC_dummy_right.icell.SM VGND.t1014 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X291 XA.XIR[14].XIC_15.icell.PUM VPWR.t1757 XA.XIR[14].XIC_15.icell.Ien VPWR.t1758 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X292 a_n997_715# XThR.XTBN.Y.t20 VGND.t1262 VGND.t1261 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X293 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[10].t17 XA.XIR[10].XIC[7].icell.Ien VGND.t2529 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X294 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[7].t12 XA.XIR[7].XIC[3].icell.Ien VGND.t862 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X295 XThC.Tn[1].t6 XThC.XTBN.Y.t19 VGND.t2362 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X296 VPWR.t1806 XThR.Tn[11].t19 XA.XIR[12].XIC[11].icell.PUM VPWR.t1805 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X297 XA.XIR[6].XIC[4].icell.PUM XThC.Tn[4].t16 XA.XIR[6].XIC[4].icell.Ien VPWR.t1331 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X298 XThR.Tn[14].t11 XThR.XTB7.Y VPWR.t947 VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X299 XA.XIR[10].XIC[12].icell.PUM XThC.Tn[12].t14 XA.XIR[10].XIC[12].icell.Ien VPWR.t1914 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X300 XA.XIR[2].XIC[5].icell.SM XA.XIR[2].XIC[5].icell.Ien Iout.t206 VGND.t1955 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X301 XA.XIR[11].XIC[1].icell.SM XA.XIR[11].XIC[1].icell.Ien Iout.t57 VGND.t641 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X302 XA.XIR[7].XIC_15.icell.PDM VPWR.t1943 VGND.t705 VGND.t704 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X303 XA.XIR[6].XIC[13].icell.SM XA.XIR[6].XIC[13].icell.Ien Iout.t91 VGND.t1120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X304 XA.XIR[13].XIC[13].icell.PUM XThC.Tn[13].t14 XA.XIR[13].XIC[13].icell.Ien VPWR.t171 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X305 VGND.t798 Vbias.t36 XA.XIR[15].XIC[12].icell.SM VGND.t797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X306 VGND.t1203 Vbias.t37 XA.XIR[14].XIC[13].icell.SM VGND.t1202 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X307 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[2].t19 XA.XIR[2].XIC[1].icell.Ien VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X308 VPWR.t546 XThR.Tn[7].t13 XA.XIR[8].XIC[0].icell.PUM VPWR.t545 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X309 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[1].t19 XA.XIR[1].XIC[13].icell.Ien VGND.t2260 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X310 VPWR.t1897 XThR.XTB5.Y a_n1049_6405# VPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X311 VPWR.t1808 XThR.Tn[11].t20 XA.XIR[12].XIC[2].icell.PUM VPWR.t1807 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X312 XThR.XTB7.B data[6].t0 VPWR.t169 VPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X313 XA.XIR[0].XIC[8].icell.PUM XThC.Tn[8].t15 XA.XIR[0].XIC[8].icell.Ien VPWR.t1265 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X314 VPWR.t209 XThC.XTB4.Y.t3 a_4861_9615# VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X315 XA.XIR[0].XIC[3].icell.SM XA.XIR[0].XIC[3].icell.Ien Iout.t42 VGND.t279 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X316 VGND.t1205 Vbias.t38 XA.XIR[5].XIC[2].icell.SM VGND.t1204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X317 XA.XIR[8].XIC[4].icell.Ien XThR.Tn[8].t21 VPWR.t670 VPWR.t669 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X318 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1754 VPWR.t1756 VPWR.t1755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X319 VGND.t1980 XThR.XTB2.Y XThR.Tn[1].t11 VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X320 XA.XIR[0].XIC[0].icell.PDM XThR.Tn[0].t18 XA.XIR[0].XIC[0].icell.Ien VGND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X321 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[11].t21 VGND.t2549 VGND.t2548 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X322 XA.XIR[12].XIC[7].icell.SM XA.XIR[12].XIC[7].icell.Ien Iout.t152 VGND.t1522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X323 XThR.XTB7.A data[4].t1 a_n1331_2891# VGND.t202 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X324 XA.XIR[8].XIC[10].icell.SM XA.XIR[8].XIC[10].icell.Ien Iout.t176 VGND.t1638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X325 VGND.t1207 Vbias.t39 XA.XIR[8].XIC[3].icell.SM VGND.t1206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X326 XA.XIR[15].XIC[13].icell.Ien VPWR.t1748 VPWR.t1750 VPWR.t1749 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X327 XA.XIR[15].XIC[8].icell.SM XA.XIR[15].XIC[8].icell.Ien Iout.t204 VGND.t1952 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X328 VPWR.t49 XThR.Tn[5].t18 XA.XIR[6].XIC[12].icell.PUM VPWR.t48 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X329 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t1944 XA.XIR[11].XIC_dummy_right.icell.Ien VGND.t706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X330 VPWR.t1278 XThR.Tn[8].t22 XA.XIR[9].XIC[13].icell.PUM VPWR.t1277 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X331 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[7].t14 XA.XIR[7].XIC[7].icell.Ien VGND.t863 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X332 a_n1049_7787# XThR.XTBN.Y.t21 XThR.Tn[1].t3 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X333 XA.XIR[5].XIC[0].icell.SM XA.XIR[5].XIC[0].icell.Ien Iout.t103 VGND.t1144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X334 XA.XIR[10].XIC[10].icell.PUM XThC.Tn[10].t15 XA.XIR[10].XIC[10].icell.Ien VPWR.t1847 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X335 VGND.t2363 XThC.XTBN.Y.t20 XThC.Tn[4].t7 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X336 XA.XIR[6].XIC[0].icell.PUM XThC.Tn[0].t15 XA.XIR[6].XIC[0].icell.Ien VPWR.t743 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X337 XA.XIR[8].XIC[1].icell.SM XA.XIR[8].XIC[1].icell.Ien Iout.t102 VGND.t1143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X338 XA.XIR[3].XIC[13].icell.SM XA.XIR[3].XIC[13].icell.Ien Iout.t127 VGND.t1338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X339 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1746 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1747 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X340 VGND.t1012 VGND.t1010 XA.XIR[12].XIC_dummy_left.icell.SM VGND.t1011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X341 XThC.XTB5.A data[1].t0 a_7331_10587# VPWR.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X342 VGND.t1299 data[1].t1 a_8739_10571# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 XA.XIR[0].XIC[1].icell.PDM VGND.t1007 VGND.t1009 VGND.t1008 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X344 VPWR.t1175 XThR.XTB2.Y XThR.Tn[9].t11 VPWR.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X345 VGND.t1264 XThR.XTBN.Y.t22 XThR.Tn[7].t2 VGND.t1263 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 VGND.t300 XThC.Tn[13].t15 XA.XIR[14].XIC[13].icell.PDM VGND.t299 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X347 XA.XIR[2].XIC[0].icell.SM XA.XIR[2].XIC[0].icell.Ien Iout.t249 VGND.t2619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X348 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1945 XA.XIR[14].XIC_dummy_left.icell.Ien VGND.t707 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X349 XThR.Tn[13].t11 XThR.XTBN.Y.t23 VPWR.t697 VPWR.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X350 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[10].t18 VGND.t2531 VGND.t2530 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X351 XA.XIR[14].XIC_15.icell.SM XA.XIR[14].XIC_15.icell.Ien Iout.t185 VGND.t1788 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X352 VGND.t1209 Vbias.t40 XA.XIR[10].XIC[11].icell.SM VGND.t1208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X353 VGND.t1006 VGND.t1004 XA.XIR[9].XIC_dummy_left.icell.SM VGND.t1005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X354 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8].t23 VPWR.t1280 VPWR.t1279 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X355 VPWR.t1090 XThR.Tn[2].t20 XA.XIR[3].XIC[9].icell.PUM VPWR.t1089 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X356 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1743 VPWR.t1745 VPWR.t1744 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X357 XA.XIR[12].XIC[13].icell.Ien XThR.Tn[12].t20 VPWR.t182 VPWR.t181 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X358 VPWR.t461 XThR.Tn[6].t19 XA.XIR[7].XIC[9].icell.PUM VPWR.t460 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X359 XA.XIR[0].XIC[3].icell.PUM XThC.Tn[3].t16 XA.XIR[0].XIC[3].icell.Ien VPWR.t138 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X360 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1695 VPWR.t1697 VPWR.t1696 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X361 VPWR.t51 XThR.Tn[5].t19 XA.XIR[6].XIC[10].icell.PUM VPWR.t50 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X362 VGND.t1595 XThC.Tn[1].t15 XA.XIR[2].XIC[1].icell.PDM VGND.t1594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X363 VGND.t265 XThR.XTB6.Y XThR.Tn[5].t3 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X364 XA.XIR[13].XIC[6].icell.PUM XThC.Tn[6].t17 XA.XIR[13].XIC[6].icell.Ien VPWR.t432 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X365 XThR.Tn[9].t6 XThR.XTB2.Y a_n997_3755# VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X366 VGND.t1211 Vbias.t41 XA.XIR[1].XIC[14].icell.SM VGND.t1210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X367 XThR.XTB6.Y XThR.XTB6.A VGND.t1769 VGND.t1634 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X368 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t1946 VGND.t709 VGND.t708 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X369 XA.XIR[12].XIC[2].icell.SM XA.XIR[12].XIC[2].icell.Ien Iout.t147 VGND.t1517 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X370 a_n997_1579# XThR.XTBN.Y.t24 VGND.t1265 VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X371 VGND.t1469 XThC.Tn[9].t15 XA.XIR[13].XIC[9].icell.PDM VGND.t1468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X372 XA.XIR[15].XIC[3].icell.SM XA.XIR[15].XIC[3].icell.Ien Iout.t16 VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X373 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[3].t18 XA.XIR[3].XIC[14].icell.Ien VGND.t1196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X374 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[3].t19 XA.XIR[3].XIC[8].icell.Ien VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X375 VPWR.t17 XThR.Tn[14].t16 XA.XIR[15].XIC[7].icell.PUM VPWR.t16 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X376 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR.t1741 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR.t1742 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X377 XA.XIR[13].XIC_dummy_right.icell.SM XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout VGND.t2606 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X378 VPWR.t1004 XThR.Tn[13].t18 XA.XIR[14].XIC[8].icell.PUM VPWR.t1003 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X379 XA.XIR[10].XIC[5].icell.PUM XThC.Tn[5].t14 XA.XIR[10].XIC[5].icell.Ien VPWR.t867 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X380 XA.XIR[15].XIC[6].icell.Ien VPWR.t1738 VPWR.t1740 VPWR.t1739 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X381 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t1947 VGND.t711 VGND.t710 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X382 VGND.t1213 Vbias.t42 XA.XIR[10].XIC[9].icell.SM VGND.t1212 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X383 VPWR.t184 XThR.Tn[12].t21 XA.XIR[13].XIC[14].icell.PUM VPWR.t183 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X384 VPWR.t1282 XThR.Tn[8].t24 XA.XIR[9].XIC[6].icell.PUM VPWR.t1281 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X385 XA.XIR[15].XIC[9].icell.PDM VPWR.t1948 XA.XIR[15].XIC[9].icell.Ien VGND.t712 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X386 XA.XIR[3].XIC[9].icell.Ien XThR.Tn[3].t20 VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X387 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[10].t19 VGND.t2533 VGND.t2532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X388 XA.XIR[15].XIC[12].icell.PDM XThR.Tn[14].t17 VGND.t2120 VGND.t2119 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X389 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1949 VGND.t714 VGND.t713 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X390 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[13].t19 VGND.t1824 VGND.t1823 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X391 VPWR.t740 XThR.XTBN.A XThR.XTBN.Y.t3 VPWR.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X392 VPWR.t53 XThR.Tn[5].t20 XA.XIR[6].XIC[5].icell.PUM VPWR.t52 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X393 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[4].t17 XA.XIR[4].XIC[11].icell.Ien VGND.t1991 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X394 XA.XIR[5].XIC[4].icell.PUM XThC.Tn[4].t17 XA.XIR[5].XIC[4].icell.Ien VPWR.t1332 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X395 VPWR.t1244 XThR.Tn[14].t18 XA.XIR[15].XIC[11].icell.PUM VPWR.t1243 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X396 XA.XIR[1].XIC[5].icell.SM XA.XIR[1].XIC[5].icell.Ien Iout.t8 VGND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X397 XA.XIR[13].XIC[1].icell.PUM XThC.Tn[1].t16 XA.XIR[13].XIC[1].icell.Ien VPWR.t885 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X398 XA.XIR[9].XIC[4].icell.PUM XThC.Tn[4].t18 XA.XIR[9].XIC[4].icell.Ien VPWR.t1333 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X399 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1736 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1737 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X400 a_3523_10575# XThC.XTB7.B VGND.t1335 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X401 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[4].t18 VGND.t2078 VGND.t2077 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X402 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[4].t19 VGND.t2080 VGND.t2079 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X403 XA.XIR[12].XIC[13].icell.PUM XThC.Tn[13].t16 XA.XIR[12].XIC[13].icell.Ien VPWR.t172 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X404 XA.XIR[4].XIC[6].icell.SM XA.XIR[4].XIC[6].icell.Ien Iout.t239 VGND.t2538 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X405 XA.XIR[11].XIC[14].icell.PUM XThC.Tn[14].t14 XA.XIR[11].XIC[14].icell.Ien VPWR.t1293 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X406 VPWR.t1369 XThC.XTBN.Y.t21 XThC.Tn[13].t11 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X407 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[1].t20 XA.XIR[1].XIC[1].icell.Ien VGND.t2261 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X408 VGND.t1215 Vbias.t43 XA.XIR[13].XIC[5].icell.SM VGND.t1214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X409 VGND.t2254 XThC.Tn[4].t19 XA.XIR[13].XIC[4].icell.PDM VGND.t2253 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X410 XA.XIR[12].XIC[6].icell.Ien XThR.Tn[12].t22 VPWR.t186 VPWR.t185 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X411 XThC.Tn[5].t3 XThC.XTB6.Y VGND.t1398 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X412 XThC.Tn[4].t1 XThC.XTB5.Y VGND.t289 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X413 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[4].t20 XA.XIR[4].XIC[2].icell.Ien VGND.t2081 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X414 VGND.t716 VPWR.t1950 XA.XIR[8].XIC_dummy_right.icell.PDM VGND.t715 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X415 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[3].t21 XA.XIR[3].XIC[3].icell.Ien VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X416 XA.XIR[14].XIC[8].icell.Ien XThR.Tn[14].t19 VPWR.t1246 VPWR.t1245 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X417 VPWR.t1248 XThR.Tn[14].t20 XA.XIR[15].XIC[2].icell.PUM VPWR.t1247 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X418 XA.XIR[2].XIC_15.icell.PDM XThR.Tn[2].t21 XA.XIR[2].XIC_15.icell.Ien VGND.t768 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X419 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t3 VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X420 VPWR.t1006 XThR.Tn[13].t20 XA.XIR[14].XIC[3].icell.PUM VPWR.t1005 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X421 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[12].t23 XA.XIR[12].XIC[9].icell.Ien VGND.t301 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X422 VPWR.t325 XThR.Tn[9].t19 XA.XIR[10].XIC[14].icell.PUM VPWR.t324 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X423 XA.XIR[15].XIC[1].icell.Ien VPWR.t1733 VPWR.t1735 VPWR.t1734 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X424 VGND.t1217 Vbias.t44 XA.XIR[11].XIC[12].icell.SM VGND.t1216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X425 VGND.t1219 Vbias.t45 XA.XIR[7].XIC_15.icell.SM VGND.t1218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X426 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1730 VPWR.t1732 VPWR.t1731 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X427 VGND.t2182 XThC.Tn[14].t15 XA.XIR[7].XIC[14].icell.PDM VGND.t2181 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X428 VGND.t2158 XThC.Tn[8].t16 XA.XIR[7].XIC[8].icell.PDM VGND.t2157 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X429 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t6 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X430 XThC.Tn[4].t6 XThC.XTBN.Y.t22 VGND.t2364 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X431 VPWR.t840 XThR.Tn[0].t19 XA.XIR[1].XIC[4].icell.PUM VPWR.t839 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X432 a_n1049_5317# XThR.XTB7.Y VPWR.t946 VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X433 XA.XIR[13].XIC[14].icell.Ien XThR.Tn[13].t21 VPWR.t1008 VPWR.t1007 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X434 XA.XIR[14].XIC[8].icell.SM XA.XIR[14].XIC[8].icell.Ien Iout.t189 VGND.t1797 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X435 XA.XIR[15].XIC[10].icell.PDM XThR.Tn[14].t21 VGND.t2122 VGND.t2121 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X436 VGND.t1221 Vbias.t46 XA.XIR[10].XIC[4].icell.SM VGND.t1220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X437 VGND.t1003 VGND.t1001 XA.XIR[5].XIC_dummy_right.icell.SM VGND.t1002 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X438 VPWR.t1284 XThR.Tn[8].t25 XA.XIR[9].XIC[1].icell.PUM VPWR.t1283 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X439 VPWR.t1211 XThR.Tn[4].t21 XA.XIR[5].XIC[4].icell.PUM VPWR.t1210 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X440 XThC.XTB6.Y XThC.XTB7.B VGND.t1334 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X441 VPWR.t1729 VPWR.t1727 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1728 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X442 XA.XIR[15].XIC[4].icell.PDM VPWR.t1951 XA.XIR[15].XIC[4].icell.Ien VGND.t717 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X443 VPWR.t235 XThR.Tn[7].t15 XA.XIR[8].XIC[13].icell.PUM VPWR.t234 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X444 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t1952 XA.XIR[10].XIC_dummy_right.icell.Ien VGND.t718 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X445 a_6243_9615# XThC.XTBN.Y.t23 XThC.Tn[6].t7 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 XA.XIR[13].XIC_dummy_left.icell.SM XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout VGND.t1142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X447 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[1].t21 VGND.t1993 VGND.t1992 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X448 XA.XIR[5].XIC[0].icell.PUM XThC.Tn[0].t16 XA.XIR[5].XIC[0].icell.Ien VPWR.t744 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X449 XA.XIR[4].XIC[10].icell.SM XA.XIR[4].XIC[10].icell.Ien Iout.t11 VGND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X450 XA.XIR[9].XIC[0].icell.PUM XThC.Tn[0].t17 XA.XIR[9].XIC[0].icell.Ien VPWR.t745 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X451 XThC.Tn[13].t7 XThC.XTB6.Y VPWR.t768 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X452 XA.XIR[5].XIC[14].icell.SM XA.XIR[5].XIC[14].icell.Ien Iout.t241 VGND.t2540 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X453 VGND.t2365 XThC.XTBN.Y.t24 XThC.Tn[0].t10 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X454 XThR.Tn[3].t11 XThR.XTBN.Y.t25 a_n1049_6699# VPWR.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X455 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[4].t22 XA.XIR[4].XIC[6].icell.Ien VGND.t2082 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X456 VGND.t1597 XThC.Tn[1].t17 XA.XIR[14].XIC[1].icell.PDM VGND.t1596 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X457 VGND.t192 XThR.XTB4.Y XThR.Tn[3].t3 VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X458 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[3].t22 XA.XIR[3].XIC[7].icell.Ien VGND.t61 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X459 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[1].t22 VGND.t1995 VGND.t1994 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X460 XA.XIR[7].XIC[9].icell.PUM XThC.Tn[9].t16 XA.XIR[7].XIC[9].icell.Ien VPWR.t806 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X461 XA.XIR[1].XIC[0].icell.SM XA.XIR[1].XIC[0].icell.Ien Iout.t9 VGND.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X462 XA.XIR[3].XIC[12].icell.PUM XThC.Tn[12].t15 XA.XIR[3].XIC[12].icell.Ien VPWR.t1915 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X463 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[4].t23 VGND.t2084 VGND.t2083 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X464 XA.XIR[0].XIC[12].icell.SM XA.XIR[0].XIC[12].icell.Ien Iout.t4 VGND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X465 XA.XIR[0].XIC_15.icell.PDM VPWR.t1953 VGND.t720 VGND.t719 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X466 XA.XIR[4].XIC[1].icell.SM XA.XIR[4].XIC[1].icell.Ien Iout.t12 VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X467 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[9].t20 VGND.t514 VGND.t513 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X468 VGND.t1223 Vbias.t47 XA.XIR[13].XIC[0].icell.SM VGND.t1222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X469 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12].t24 VPWR.t188 VPWR.t187 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X470 XA.XIR[6].XIC[13].icell.PUM XThC.Tn[13].t17 XA.XIR[6].XIC[13].icell.Ien VPWR.t173 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X471 VGND.t1225 Vbias.t48 XA.XIR[8].XIC[12].icell.SM VGND.t1224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X472 XA.XIR[2].XIC[14].icell.SM XA.XIR[2].XIC[14].icell.Ien Iout.t7 VGND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X473 XThR.Tn[11].t7 XThR.XTB4.Y VPWR.t89 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X474 VGND.t2160 XThC.Tn[8].t17 XA.XIR[4].XIC[8].icell.PDM VGND.t2159 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X475 VGND.t2184 XThC.Tn[14].t16 XA.XIR[4].XIC[14].icell.PDM VGND.t2183 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X476 XThC.Tn[14].t3 XThC.XTB7.Y a_10915_9569# VGND.t223 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X477 VPWR.t842 XThR.Tn[0].t20 XA.XIR[1].XIC[0].icell.PUM VPWR.t841 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X478 XA.XIR[14].XIC[3].icell.Ien XThR.Tn[14].t22 VPWR.t1250 VPWR.t1249 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X479 VGND.t2672 XThC.Tn[12].t16 XA.XIR[11].XIC[12].icell.PDM VGND.t2671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X480 VPWR.t1213 XThR.Tn[4].t24 XA.XIR[5].XIC[0].icell.PUM VPWR.t1212 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X481 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[12].t25 XA.XIR[12].XIC[4].icell.Ien VGND.t302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X482 XA.XIR[12].XIC[6].icell.PUM XThC.Tn[6].t18 XA.XIR[12].XIC[6].icell.Ien VPWR.t433 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X483 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t1954 XA.XIR[7].XIC_dummy_right.icell.Ien VGND.t721 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X484 VPWR.t1726 VPWR.t1724 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1725 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X485 XA.XIR[15].XIC[7].icell.PUM XThC.Tn[7].t11 XA.XIR[15].XIC[7].icell.Ien VPWR.t1258 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X486 VGND.t327 XThC.XTB4.Y.t4 XThC.Tn[3].t11 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X487 VPWR.t108 XThC.XTB2.Y XThC.Tn[9].t2 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X488 XA.XIR[5].XIC[12].icell.Ien XThR.Tn[5].t21 VPWR.t55 VPWR.t54 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X489 VGND.t270 XThC.Tn[3].t17 XA.XIR[7].XIC[3].icell.PDM VGND.t269 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X490 VGND.t1044 Vbias.t49 XA.XIR[6].XIC[11].icell.SM VGND.t1043 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X491 VGND.t723 VPWR.t1955 XA.XIR[2].XIC_15.icell.PDM VGND.t722 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X492 VPWR.t1896 XThR.XTB5.Y XThR.Tn[12].t10 VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VGND.t1471 XThC.Tn[9].t17 XA.XIR[12].XIC[9].icell.PDM VGND.t1470 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X494 XA.XIR[14].XIC[3].icell.SM XA.XIR[14].XIC[3].icell.Ien Iout.t179 VGND.t1642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X495 XA.XIR[9].XIC[12].icell.Ien XThR.Tn[9].t21 VPWR.t327 VPWR.t326 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X496 XA.XIR[8].XIC[13].icell.Ien XThR.Tn[8].t26 VPWR.t1286 VPWR.t1285 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X497 XA.XIR[12].XIC_dummy_right.icell.SM XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout VGND.t1303 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X498 XA.XIR[6].XIC[14].icell.PDM XThR.Tn[6].t20 XA.XIR[6].XIC[14].icell.Ien VGND.t667 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X499 XA.XIR[6].XIC[8].icell.PDM XThR.Tn[6].t21 XA.XIR[6].XIC[8].icell.Ien VGND.t668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X500 VPWR.t945 XThR.XTB7.Y XThR.Tn[14].t10 VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X501 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[1].t23 VGND.t1997 VGND.t1996 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X502 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[13].t22 XA.XIR[13].XIC[12].icell.Ien VGND.t1825 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X503 XA.XIR[4].XIC[9].icell.PUM XThC.Tn[9].t18 XA.XIR[4].XIC[9].icell.Ien VPWR.t807 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X504 XThR.Tn[8].t8 XThR.XTB1.Y.t4 a_n997_3979# VGND.t1554 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X505 XA.XIR[3].XIC[10].icell.PUM XThC.Tn[10].t16 XA.XIR[3].XIC[10].icell.Ien VPWR.t1848 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X506 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[4].t25 VGND.t1604 VGND.t1603 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X507 VGND.t849 XThC.Tn[11].t17 XA.XIR[1].XIC[11].icell.PDM VGND.t848 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X508 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t1956 VGND.t725 VGND.t724 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X509 VPWR.t237 XThR.Tn[7].t16 XA.XIR[8].XIC[6].icell.PUM VPWR.t236 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X510 VPWR.t1268 data[2].t0 XThC.XTB7.B VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X511 VGND.t1000 VGND.t998 XA.XIR[5].XIC_dummy_left.icell.SM VGND.t999 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X512 VPWR.t1410 XThR.Tn[10].t20 XA.XIR[11].XIC[7].icell.PUM VPWR.t1409 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X513 VGND.t2569 XThC.Tn[10].t17 XA.XIR[11].XIC[10].icell.PDM VGND.t2568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X514 XThC.Tn[13].t2 XThC.XTB6.Y a_10051_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X515 XThR.Tn[4].t3 XThR.XTBN.Y.t26 a_n1049_6405# VPWR.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X516 XThR.XTB5.Y XThR.XTB7.B a_n1319_6405# VPWR.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X517 VGND.t1046 Vbias.t50 XA.XIR[4].XIC[7].icell.SM VGND.t1045 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X518 XThC.Tn[8].t11 XThC.XTBN.Y.t25 VPWR.t1371 VPWR.t1370 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X519 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[13].t23 VGND.t1827 VGND.t1826 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X520 XA.XIR[15].XIC[11].icell.PUM XThC.Tn[11].t18 XA.XIR[15].XIC[11].icell.Ien VPWR.t534 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X521 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[9].t22 VGND.t516 VGND.t515 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X522 a_n1335_4229# data[5].t0 XThR.XTB5.A VPWR.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X523 VGND.t1626 XThC.Tn[2].t17 XA.XIR[1].XIC[2].icell.PDM VGND.t1625 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X524 VGND.t1048 Vbias.t51 XA.XIR[7].XIC[8].icell.SM VGND.t1047 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X525 XA.XIR[6].XIC[9].icell.Ien XThR.Tn[6].t22 VPWR.t463 VPWR.t462 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X526 XA.XIR[5].XIC[10].icell.Ien XThR.Tn[5].t22 VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X527 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[12].t26 VGND.t304 VGND.t303 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X528 VGND.t2138 XThC.Tn[7].t12 XA.XIR[7].XIC[7].icell.PDM VGND.t2137 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X529 VGND.t1050 Vbias.t52 XA.XIR[6].XIC[9].icell.SM VGND.t1049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X530 VGND.t1052 Vbias.t53 XA.XIR[3].XIC[11].icell.SM VGND.t1051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X531 XThC.Tn[8].t2 XThC.XTB1.Y.t4 a_7651_9569# VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X532 XThC.Tn[13].t10 XThC.XTBN.Y.t26 VPWR.t1372 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X533 VGND.t272 XThC.Tn[3].t18 XA.XIR[4].XIC[3].icell.PDM VGND.t271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X534 XA.XIR[9].XIC[10].icell.Ien XThR.Tn[9].t23 VPWR.t329 VPWR.t328 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X535 XA.XIR[7].XIC_15.icell.SM XA.XIR[7].XIC_15.icell.Ien Iout.t118 VGND.t1304 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X536 XA.XIR[15].XIC[12].icell.SM XA.XIR[15].XIC[12].icell.Ien Iout.t119 VGND.t1305 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X537 VPWR.t594 VGND.t2691 XA.XIR[0].XIC[9].icell.PUM VPWR.t593 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X538 VGND.t1397 XThC.XTB6.Y XThC.Tn[5].t2 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X539 XA.XIR[12].XIC[1].icell.PUM XThC.Tn[1].t18 XA.XIR[12].XIC[1].icell.Ien VPWR.t886 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X540 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1698 VPWR.t1700 VPWR.t1699 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X541 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[3].t23 VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X542 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[3].t24 VGND.t65 VGND.t64 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X543 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[13].t24 XA.XIR[13].XIC[10].icell.Ien VGND.t1828 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X544 XA.XIR[15].XIC[2].icell.PUM XThC.Tn[2].t18 XA.XIR[15].XIC[2].icell.Ien VPWR.t919 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X545 XA.XIR[6].XIC[6].icell.PUM XThC.Tn[6].t19 XA.XIR[6].XIC[6].icell.Ien VPWR.t434 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X546 XA.XIR[10].XIC[14].icell.PUM XThC.Tn[14].t17 XA.XIR[10].XIC[14].icell.Ien VPWR.t94 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X547 VGND.t1054 Vbias.t54 XA.XIR[12].XIC[5].icell.SM VGND.t1053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X548 VGND.t2098 XThC.Tn[4].t20 XA.XIR[12].XIC[4].icell.PDM VGND.t2097 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X549 a_n1049_5611# XThR.XTB6.Y VPWR.t133 VPWR.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 XA.XIR[13].XIC_15.icell.PUM VPWR.t1722 XA.XIR[13].XIC_15.icell.Ien VPWR.t1723 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X551 XThR.Tn[10].t1 XThR.XTB3.Y.t4 a_n997_2891# VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X552 VGND.t1056 Vbias.t55 XA.XIR[15].XIC[6].icell.SM VGND.t1055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X553 XA.XIR[0].XIC[11].icell.PDM XThR.Tn[0].t21 XA.XIR[0].XIC[11].icell.Ien VGND.t1528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X554 VGND.t1571 XThC.Tn[5].t15 XA.XIR[15].XIC[5].icell.PDM VGND.t1570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X555 VGND.t1473 XThC.Tn[9].t19 XA.XIR[6].XIC[9].icell.PDM VGND.t1472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X556 VPWR.t264 XThC.XTBN.Y.t27 XThC.Tn[7].t6 VPWR.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X557 XA.XIR[6].XIC[3].icell.PDM XThR.Tn[6].t23 XA.XIR[6].XIC[3].icell.Ien VGND.t2655 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X558 XA.XIR[1].XIC_15.icell.PDM XThR.Tn[1].t24 XA.XIR[1].XIC_15.icell.Ien VGND.t1998 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X559 VPWR.t1412 XThR.Tn[10].t21 XA.XIR[11].XIC[11].icell.PUM VPWR.t1411 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X560 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR.t1720 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1721 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X561 VPWR.t1173 XThR.XTB2.Y XThR.Tn[9].t10 VPWR.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X562 XThC.Tn[6].t6 XThC.XTBN.Y.t28 a_6243_9615# VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X563 XA.XIR[3].XIC[5].icell.PUM XThC.Tn[5].t16 XA.XIR[3].XIC[5].icell.Ien VPWR.t868 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X564 VPWR.t748 bias[1].t0 Vbias.t3 VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.1275 pd=1.15 as=0.1955 ps=1.31 w=0.85 l=1
X565 VGND.t1058 Vbias.t56 XA.XIR[9].XIC[5].icell.SM VGND.t1057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X566 XA.XIR[8].XIC[6].icell.Ien XThR.Tn[8].t27 VPWR.t1288 VPWR.t1287 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X567 VGND.t632 XThC.Tn[6].t20 XA.XIR[1].XIC[6].icell.PDM VGND.t631 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X568 VPWR.t7 XThR.Tn[3].t25 XA.XIR[4].XIC[4].icell.PUM VPWR.t6 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X569 VPWR.t239 XThR.Tn[7].t17 XA.XIR[8].XIC[1].icell.PUM VPWR.t238 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X570 XA.XIR[0].XIC[2].icell.PDM XThR.Tn[0].t22 XA.XIR[0].XIC[2].icell.Ien VGND.t1925 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X571 XA.XIR[11].XIC[7].icell.Ien XThR.Tn[11].t22 VPWR.t1810 VPWR.t1809 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X572 VGND.t1060 Vbias.t57 XA.XIR[3].XIC[9].icell.SM VGND.t1059 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X573 VGND.t2140 XThC.Tn[7].t13 XA.XIR[4].XIC[7].icell.PDM VGND.t2139 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X574 XA.XIR[15].XIC_15.icell.Ien VPWR.t1717 VPWR.t1719 VPWR.t1718 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X575 VPWR.t1121 XThR.Tn[10].t22 XA.XIR[11].XIC[2].icell.PUM VPWR.t1120 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X576 XA.XIR[12].XIC_dummy_left.icell.SM XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout VGND.t2141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X577 VPWR.t59 XThR.Tn[5].t23 XA.XIR[6].XIC[14].icell.PUM VPWR.t58 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X578 a_n1049_7493# XThR.XTBN.Y.t27 XThR.Tn[2].t5 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X579 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[8].t28 XA.XIR[8].XIC[9].icell.Ien VGND.t2168 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X580 XThC.Tn[0].t9 XThC.XTBN.Y.t29 VGND.t414 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X581 VGND.t1062 Vbias.t58 XA.XIR[4].XIC[2].icell.SM VGND.t1061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X582 VPWR.t1716 VPWR.t1714 XA.XIR[9].XIC_15.icell.PUM VPWR.t1715 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X583 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[0].t23 VGND.t1927 VGND.t1926 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X584 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[0].t24 VGND.t1929 VGND.t1928 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X585 VGND.t1064 Vbias.t59 XA.XIR[7].XIC[3].icell.SM VGND.t1063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X586 a_4067_9615# XThC.XTBN.Y.t30 XThC.Tn[2].t7 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X587 XThR.Tn[0].t9 XThR.XTB1.Y.t5 VGND.t1556 VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X588 VGND.t544 XThR.XTBN.Y.t28 XThR.Tn[5].t10 VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 XA.XIR[11].XIC[7].icell.SM XA.XIR[11].XIC[7].icell.Ien Iout.t224 VGND.t2310 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X590 XA.XIR[5].XIC[5].icell.Ien XThR.Tn[5].t24 VPWR.t61 VPWR.t60 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X591 VGND.t1066 Vbias.t60 XA.XIR[6].XIC[4].icell.SM VGND.t1065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X592 XThR.Tn[14].t7 XThR.XTB7.Y a_n997_715# VGND.t1750 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X593 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[12].t27 VGND.t306 VGND.t305 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X594 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[7].t18 VGND.t390 VGND.t389 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X595 VGND.t1227 Vbias.t61 XA.XIR[15].XIC[10].icell.SM VGND.t1226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X596 XA.XIR[9].XIC[5].icell.Ien XThR.Tn[9].t24 VPWR.t331 VPWR.t330 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X597 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[10].t23 VGND.t1917 VGND.t1916 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X598 XA.XIR[10].XIC[11].icell.SM XA.XIR[10].XIC[11].icell.Ien Iout.t79 VGND.t873 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X599 VGND.t727 VPWR.t1957 XA.XIR[11].XIC_dummy_left.icell.PDM VGND.t726 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X600 XA.XIR[6].XIC[7].icell.PDM XThR.Tn[6].t24 XA.XIR[6].XIC[7].icell.Ien VGND.t2656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X601 VGND.t546 XThR.XTBN.Y.t29 XThR.Tn[4].t7 VGND.t545 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X602 VPWR.t978 bias[1].t1 Vbias.t9 VPWR.t747 sky130_fd_pr__pfet_01v8 ad=0.1275 pd=1.15 as=0.1955 ps=1.31 w=0.85 l=1
X603 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[3].t26 VGND.t67 VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X604 XA.XIR[6].XIC[1].icell.PUM XThC.Tn[1].t19 XA.XIR[6].XIC[1].icell.Ien VPWR.t887 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X605 VGND.t729 VPWR.t1958 XA.XIR[14].XIC_15.icell.PDM VGND.t728 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X606 a_8963_9569# XThC.XTB4.Y.t5 XThC.Tn[11].t0 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X607 XA.XIR[5].XIC[13].icell.PUM XThC.Tn[13].t18 XA.XIR[5].XIC[13].icell.Ien VPWR.t174 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X608 VGND.t1229 Vbias.t62 XA.XIR[12].XIC[0].icell.SM VGND.t1228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X609 XA.XIR[1].XIC[14].icell.SM XA.XIR[1].XIC[14].icell.Ien Iout.t212 VGND.t2143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X610 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR.t1712 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR.t1713 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X611 XA.XIR[9].XIC[13].icell.PUM XThC.Tn[13].t19 XA.XIR[9].XIC[13].icell.Ien VPWR.t1354 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X612 VGND.t1231 Vbias.t63 XA.XIR[15].XIC[1].icell.SM VGND.t1230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X613 XA.XIR[0].XIC[6].icell.PDM XThR.Tn[0].t25 XA.XIR[0].XIC[6].icell.Ien VGND.t1930 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X614 VGND.t2100 XThC.Tn[4].t21 XA.XIR[6].XIC[4].icell.PDM VGND.t2099 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X615 VGND.t1379 XThC.Tn[0].t18 XA.XIR[15].XIC[0].icell.PDM VGND.t1378 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X616 VGND.t1233 Vbias.t64 XA.XIR[10].XIC[13].icell.SM VGND.t1232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X617 XA.XIR[11].XIC[11].icell.Ien XThR.Tn[11].t23 VPWR.t1812 VPWR.t1811 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X618 VGND.t2674 XThC.Tn[12].t17 XA.XIR[10].XIC[12].icell.PDM VGND.t2673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X619 VPWR.t9 XThR.Tn[3].t27 XA.XIR[4].XIC[0].icell.PUM VPWR.t8 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X620 VGND.t1235 Vbias.t65 XA.XIR[13].XIC[14].icell.SM VGND.t1234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X621 XA.XIR[12].XIC_15.icell.Ien XThR.Tn[12].t28 VPWR.t190 VPWR.t189 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X622 VGND.t415 XThC.XTBN.Y.t31 a_8739_9569# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X623 VGND.t2297 XThC.Tn[13].t20 XA.XIR[13].XIC[13].icell.PDM VGND.t2296 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X624 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t1959 XA.XIR[13].XIC_dummy_left.icell.Ien VGND.t730 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X625 VGND.t1237 Vbias.t66 XA.XIR[9].XIC[0].icell.SM VGND.t1236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X626 XA.XIR[4].XIC[4].icell.Ien XThR.Tn[4].t26 VPWR.t898 VPWR.t897 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X627 XA.XIR[8].XIC[1].icell.Ien XThR.Tn[8].t29 VPWR.t296 VPWR.t295 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X628 VGND.t1239 Vbias.t67 XA.XIR[0].XIC_15.icell.SM VGND.t1238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X629 VGND.t2162 XThC.Tn[8].t18 XA.XIR[0].XIC[8].icell.PDM VGND.t2161 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X630 VGND.t195 XThC.Tn[14].t18 XA.XIR[0].XIC[14].icell.PDM VGND.t194 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X631 XA.XIR[11].XIC[2].icell.Ien XThR.Tn[11].t24 VPWR.t1814 VPWR.t1813 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X632 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[7].t19 VGND.t392 VGND.t391 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X633 XA.XIR[8].XIC[7].icell.SM XA.XIR[8].XIC[7].icell.Ien Iout.t157 VGND.t1532 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X634 a_9827_9569# XThC.XTBN.Y.t32 VGND.t416 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X635 VGND.t1241 Vbias.t68 XA.XIR[3].XIC[4].icell.SM VGND.t1240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X636 XA.XIR[7].XIC[8].icell.SM XA.XIR[7].XIC[8].icell.Ien Iout.t214 VGND.t2145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X637 VPWR.t1185 XThR.Tn[1].t25 XA.XIR[2].XIC[12].icell.PUM VPWR.t1184 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X638 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[8].t30 XA.XIR[8].XIC[4].icell.Ien VGND.t468 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X639 VPWR.t1129 XThR.Tn[0].t26 XA.XIR[1].XIC[13].icell.PUM VPWR.t1128 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X640 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t1960 XA.XIR[3].XIC_dummy_right.icell.Ien VGND.t731 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X641 XA.XIR[10].XIC[9].icell.SM XA.XIR[10].XIC[9].icell.Ien Iout.t18 VGND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X642 VPWR.t900 XThR.Tn[4].t27 XA.XIR[5].XIC[13].icell.PUM VPWR.t899 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X643 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[11].t25 XA.XIR[11].XIC[5].icell.Ien VGND.t166 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X644 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[3].t28 VGND.t69 VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X645 VPWR.t1711 VPWR.t1709 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1710 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X646 XA.XIR[15].XIC[13].icell.PDM VPWR.t1961 XA.XIR[15].XIC[13].icell.Ien VGND.t732 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X647 VGND.t2553 XThC.XTB1.Y.t5 XThC.Tn[0].t11 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X648 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[0].t27 VGND.t1932 VGND.t1931 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X649 XA.XIR[11].XIC[2].icell.SM XA.XIR[11].XIC[2].icell.Ien Iout.t178 VGND.t1640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X650 XThR.XTB7.A data[5].t1 VPWR.t93 VPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X651 VGND.t2571 XThC.Tn[10].t18 XA.XIR[10].XIC[10].icell.PDM VGND.t2570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X652 VPWR.t192 XThR.Tn[12].t29 XA.XIR[13].XIC[8].icell.PUM VPWR.t191 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X653 VGND.t676 XThC.XTBN.A XThC.XTBN.Y.t1 VGND.t675 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X654 XA.XIR[0].XIC[9].icell.PUM XThC.Tn[9].t20 XA.XIR[0].XIC[9].icell.Ien VPWR.t808 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X655 VPWR.t881 XThR.XTB7.B XThR.XTB1.Y.t0 VPWR.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X656 a_n997_1579# XThR.XTB6.Y XThR.Tn[13].t2 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X657 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[2].t22 VGND.t815 VGND.t814 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X658 XA.XIR[4].XIC[0].icell.Ien XThR.Tn[4].t28 VPWR.t902 VPWR.t901 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X659 XA.XIR[14].XIC[12].icell.SM XA.XIR[14].XIC[12].icell.Ien Iout.t123 VGND.t1323 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X660 XA.XIR[14].XIC_15.icell.PDM VPWR.t1962 VGND.t734 VGND.t733 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X661 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1706 VPWR.t1708 VPWR.t1707 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X662 XA.XIR[13].XIC[5].icell.SM XA.XIR[13].XIC[5].icell.Ien Iout.t34 VGND.t224 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X663 VPWR.t1187 XThR.Tn[1].t26 XA.XIR[2].XIC[10].icell.PUM VPWR.t1186 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X664 XA.XIR[5].XIC[6].icell.PUM XThC.Tn[6].t21 XA.XIR[5].XIC[6].icell.Ien VPWR.t435 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X665 XThC.Tn[7].t5 XThC.XTBN.Y.t33 VPWR.t266 VPWR.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X666 VGND.t1588 XThR.XTB7.B a_n1335_7243# VGND.t1587 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X667 XA.XIR[9].XIC[6].icell.PUM XThC.Tn[6].t22 XA.XIR[9].XIC[6].icell.Ien VPWR.t436 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X668 XA.XIR[8].XIC[7].icell.PUM XThC.Tn[7].t14 XA.XIR[8].XIC[7].icell.Ien VPWR.t699 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X669 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[0].t28 VGND.t1934 VGND.t1933 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X670 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t1963 VGND.t736 VGND.t735 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X671 XA.XIR[12].XIC_15.icell.PUM VPWR.t1704 XA.XIR[12].XIC_15.icell.Ien VPWR.t1705 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X672 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[8].t31 VGND.t470 VGND.t469 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X673 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[12].t30 XA.XIR[12].XIC[13].icell.Ien VGND.t307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X674 VGND.t274 XThC.Tn[3].t19 XA.XIR[0].XIC[3].icell.PDM VGND.t273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X675 XA.XIR[11].XIC[8].icell.PUM XThC.Tn[8].t19 XA.XIR[11].XIC[8].icell.Ien VPWR.t1266 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X676 VGND.t1475 XThC.Tn[9].t21 XA.XIR[5].XIC[9].icell.PDM VGND.t1474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X677 XA.XIR[8].XIC[2].icell.SM XA.XIR[8].XIC[2].icell.Ien Iout.t199 VGND.t1914 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X678 XA.XIR[2].XIC[12].icell.Ien XThR.Tn[2].t23 VPWR.t1088 VPWR.t1087 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X679 XA.XIR[7].XIC[3].icell.SM XA.XIR[7].XIC[3].icell.Ien Iout.t27 VGND.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X680 XThC.Tn[11].t1 XThC.XTB4.Y.t6 VPWR.t211 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 VGND.t1774 XThC.Tn[9].t22 XA.XIR[9].XIC[9].icell.PDM VGND.t1773 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X682 XA.XIR[10].XIC[4].icell.SM XA.XIR[10].XIC[4].icell.Ien Iout.t43 VGND.t292 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X683 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1701 VPWR.t1703 VPWR.t1702 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X684 a_n997_1803# XThR.XTBN.Y.t30 VGND.t548 VGND.t547 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X685 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[11].t26 XA.XIR[11].XIC[0].icell.Ien VGND.t167 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X686 XThR.Tn[3].t10 XThR.XTBN.Y.t31 a_n1049_6699# VPWR.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X687 VPWR.t333 XThR.Tn[9].t25 XA.XIR[10].XIC[8].icell.PUM VPWR.t332 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X688 VGND.t549 XThR.XTBN.Y.t32 XThR.Tn[3].t6 VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X689 VGND.t1243 Vbias.t69 XA.XIR[11].XIC[6].icell.SM VGND.t1242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X690 XA.XIR[10].XIC[7].icell.Ien XThR.Tn[10].t24 VPWR.t1123 VPWR.t1122 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X691 VGND.t738 VPWR.t1964 XA.XIR[7].XIC_dummy_right.icell.PDM VGND.t737 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X692 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t1965 VGND.t740 VGND.t739 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X693 XThC.Tn[2].t6 XThC.XTBN.Y.t34 a_4067_9615# VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X694 VPWR.t783 XThR.Tn[0].t29 XA.XIR[1].XIC[6].icell.PUM VPWR.t782 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X695 XA.XIR[13].XIC[8].icell.Ien XThR.Tn[13].t25 VPWR.t1010 VPWR.t1009 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X696 VPWR.t904 XThR.Tn[4].t29 XA.XIR[5].XIC[6].icell.PUM VPWR.t903 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X697 VPWR.t194 XThR.Tn[12].t31 XA.XIR[13].XIC[3].icell.PUM VPWR.t193 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X698 XThR.Tn[11].t6 XThR.XTB4.Y VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X699 VPWR.t1694 VPWR.t1692 XA.XIR[8].XIC_15.icell.PUM VPWR.t1693 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X700 VPWR.t107 XThC.XTB2.Y a_3773_9615# VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X701 a_n1049_8581# XThR.XTB1.Y.t6 VPWR.t855 VPWR.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1690 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1691 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X703 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[2].t24 VGND.t813 VGND.t812 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X704 XA.XIR[8].XIC[11].icell.PUM XThC.Tn[11].t19 XA.XIR[8].XIC[11].icell.Ien VPWR.t535 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X705 VGND.t1245 Vbias.t70 XA.XIR[0].XIC[8].icell.SM VGND.t1244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X706 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[10].t25 VGND.t1919 VGND.t1918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X707 VGND.t1272 XThC.Tn[7].t15 XA.XIR[0].XIC[7].icell.PDM VGND.t1271 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X708 VGND.t997 VGND.t995 XA.XIR[4].XIC_dummy_right.icell.SM VGND.t996 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X709 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[5].t25 VGND.t160 VGND.t159 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X710 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[9].t26 VGND.t518 VGND.t517 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X711 XA.XIR[9].XIC[11].icell.SM XA.XIR[9].XIC[11].icell.Ien Iout.t146 VGND.t1476 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X712 XA.XIR[2].XIC[10].icell.Ien XThR.Tn[2].t25 VPWR.t1086 VPWR.t1085 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X713 XA.XIR[13].XIC[0].icell.SM XA.XIR[13].XIC[0].icell.Ien Iout.t121 VGND.t1321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X714 VGND.t742 VPWR.t1966 XA.XIR[10].XIC_dummy_left.icell.PDM VGND.t741 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X715 VPWR.t1883 XThC.XTB6.A a_5949_10571# VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X716 VPWR.t1189 XThR.Tn[1].t27 XA.XIR[2].XIC[5].icell.PUM VPWR.t1188 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X717 XA.XIR[1].XIC[4].icell.PUM XThC.Tn[4].t22 XA.XIR[1].XIC[4].icell.Ien VPWR.t1220 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X718 XA.XIR[5].XIC[1].icell.PUM XThC.Tn[1].t20 XA.XIR[5].XIC[1].icell.Ien VPWR.t888 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X719 VGND.t1250 XThR.XTB3.Y.t5 XThR.Tn[2].t7 VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X720 VPWR.t1012 XThR.Tn[13].t26 XA.XIR[14].XIC[9].icell.PUM VPWR.t1011 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X721 XA.XIR[9].XIC[1].icell.PUM XThC.Tn[1].t21 XA.XIR[9].XIC[1].icell.Ien VPWR.t1363 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X722 XA.XIR[8].XIC[2].icell.PUM XThC.Tn[2].t19 XA.XIR[8].XIC[2].icell.Ien VPWR.t920 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X723 XA.XIR[3].XIC[14].icell.PUM XThC.Tn[14].t19 XA.XIR[3].XIC[14].icell.Ien VPWR.t95 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X724 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[8].t32 VGND.t472 VGND.t471 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X725 XA.XIR[0].XIC[6].icell.SM XA.XIR[0].XIC[6].icell.Ien Iout.t228 VGND.t2505 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X726 XThC.XTBN.Y.t3 XThC.XTBN.A VPWR.t471 VPWR.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X727 VGND.t1247 Vbias.t71 XA.XIR[5].XIC[5].icell.SM VGND.t1246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X728 XA.XIR[11].XIC[3].icell.PUM XThC.Tn[3].t20 XA.XIR[11].XIC[3].icell.Ien VPWR.t139 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X729 VGND.t2102 XThC.Tn[4].t23 XA.XIR[5].XIC[4].icell.PDM VGND.t2101 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X730 VGND.t1249 Vbias.t72 XA.XIR[11].XIC[10].icell.SM VGND.t1248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X731 XA.XIR[10].XIC[11].icell.Ien XThR.Tn[10].t26 VPWR.t1125 VPWR.t1124 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X732 XThR.Tn[8].t9 XThR.XTB1.Y.t7 a_n997_3979# VGND.t1557 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X733 XA.XIR[6].XIC_15.icell.PUM VPWR.t1688 XA.XIR[6].XIC_15.icell.Ien VPWR.t1689 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X734 VGND.t2323 XThC.Tn[1].t22 XA.XIR[13].XIC[1].icell.PDM VGND.t2322 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X735 VGND.t1073 Vbias.t73 XA.XIR[12].XIC[14].icell.SM VGND.t1072 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X736 VGND.t2104 XThC.Tn[4].t24 XA.XIR[9].XIC[4].icell.PDM VGND.t2103 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X737 VGND.t1075 Vbias.t74 XA.XIR[8].XIC[6].icell.SM VGND.t1074 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X738 XA.XIR[7].XIC[7].icell.Ien XThR.Tn[7].t20 VPWR.t241 VPWR.t240 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X739 VGND.t744 VPWR.t1967 XA.XIR[4].XIC_dummy_right.icell.PDM VGND.t743 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X740 VGND.t1573 XThC.Tn[5].t17 XA.XIR[8].XIC[5].icell.PDM VGND.t1572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X741 VGND.t2299 XThC.Tn[13].t21 XA.XIR[12].XIC[13].icell.PDM VGND.t2298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X742 VGND.t417 XThC.XTBN.Y.t35 a_9827_9569# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X743 XA.XIR[2].XIC[12].icell.PUM XThC.Tn[12].t18 XA.XIR[2].XIC[12].icell.Ien VPWR.t954 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X744 VPWR.t335 XThR.Tn[9].t27 XA.XIR[10].XIC[3].icell.PUM VPWR.t334 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X745 VPWR.t118 XThC.XTB7.Y XThC.Tn[14].t7 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X746 XThR.Tn[4].t2 XThR.XTBN.Y.t33 a_n1049_6405# VPWR.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X747 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[14].t23 XA.XIR[14].XIC[8].icell.Ien VGND.t2123 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X748 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[14].t24 XA.XIR[14].XIC[14].icell.Ien VGND.t2124 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X749 VGND.t1077 Vbias.t75 XA.XIR[11].XIC[1].icell.SM VGND.t1076 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X750 XA.XIR[10].XIC[2].icell.Ien XThR.Tn[10].t27 VPWR.t1127 VPWR.t1126 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X751 VGND.t1079 Vbias.t76 XA.XIR[7].XIC[12].icell.SM VGND.t1078 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X752 VPWR.t85 XThR.XTB4.Y a_n1049_6699# VPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X753 XA.XIR[5].XIC[14].icell.Ien XThR.Tn[5].t26 VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X754 VGND.t1081 Vbias.t77 XA.XIR[6].XIC[13].icell.SM VGND.t1080 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X755 VPWR.t785 XThR.Tn[0].t30 XA.XIR[1].XIC[1].icell.PUM VPWR.t784 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X756 XA.XIR[13].XIC[3].icell.Ien XThR.Tn[13].t27 VPWR.t1014 VPWR.t1013 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X757 XA.XIR[9].XIC[14].icell.Ien XThR.Tn[9].t28 VPWR.t337 VPWR.t336 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X758 VGND.t1083 Vbias.t78 XA.XIR[9].XIC[14].icell.SM VGND.t1082 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X759 VPWR.t906 XThR.Tn[4].t30 XA.XIR[5].XIC[1].icell.PUM VPWR.t905 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X760 XA.XIR[9].XIC[9].icell.SM XA.XIR[9].XIC[9].icell.Ien Iout.t172 VGND.t1631 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X761 XA.XIR[8].XIC_15.icell.Ien XThR.Tn[8].t33 VPWR.t298 VPWR.t297 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X762 XA.XIR[15].XIC[1].icell.PDM VPWR.t1968 XA.XIR[15].XIC[1].icell.Ien VGND.t745 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X763 VPWR.t11 XThR.Tn[3].t29 XA.XIR[4].XIC[13].icell.PUM VPWR.t10 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X764 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[10].t28 XA.XIR[10].XIC[5].icell.Ien VGND.t1920 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X765 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR.t1969 XA.XIR[6].XIC_dummy_right.icell.Ien VGND.t746 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X766 XA.XIR[0].XIC[4].icell.Ien XThR.Tn[0].t31 VPWR.t787 VPWR.t786 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X767 XA.XIR[1].XIC[0].icell.PUM XThC.Tn[0].t19 XA.XIR[1].XIC[0].icell.Ien VPWR.t746 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X768 VGND.t1085 Vbias.t79 XA.XIR[0].XIC[3].icell.SM VGND.t1084 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X769 XA.XIR[4].XIC[7].icell.SM XA.XIR[4].XIC[7].icell.Ien Iout.t29 VGND.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X770 XA.XIR[0].XIC[10].icell.SM XA.XIR[0].XIC[10].icell.Ien Iout.t72 VGND.t845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X771 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[5].t27 VGND.t162 VGND.t161 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X772 XA.XIR[2].XIC[5].icell.Ien XThR.Tn[2].t26 VPWR.t1084 VPWR.t1083 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X773 XA.XIR[11].XIC_dummy_right.icell.SM XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X774 VGND.t1087 Vbias.t80 XA.XIR[8].XIC[10].icell.SM VGND.t1086 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X775 VPWR.t373 XThR.XTBN.Y.t34 XThR.Tn[8].t7 VPWR.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X776 XA.XIR[7].XIC[11].icell.Ien XThR.Tn[7].t21 VPWR.t243 VPWR.t242 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X777 XThR.Tn[10].t8 XThR.XTB3.Y.t6 a_n997_2891# VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X778 XA.XIR[14].XIC[9].icell.Ien XThR.Tn[14].t25 VPWR.t1252 VPWR.t1251 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X779 XA.XIR[2].XIC[10].icell.PUM XThC.Tn[10].t19 XA.XIR[2].XIC[10].icell.Ien VPWR.t1849 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X780 XThC.XTB3.Y.t0 XThC.XTB7.B VPWR.t729 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X781 XA.XIR[0].XIC[1].icell.SM XA.XIR[0].XIC[1].icell.Ien Iout.t196 VGND.t1804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X782 VGND.t1089 Vbias.t81 XA.XIR[5].XIC[0].icell.SM VGND.t1088 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X783 VGND.t994 VGND.t992 XA.XIR[4].XIC_dummy_left.icell.SM VGND.t993 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X784 VGND.t1091 Vbias.t82 XA.XIR[8].XIC[1].icell.SM VGND.t1090 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X785 VPWR.t1882 XThC.XTB6.A XThC.XTB2.Y VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X786 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[11].t27 VGND.t169 VGND.t168 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X787 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[11].t28 VGND.t171 VGND.t170 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X788 XA.XIR[12].XIC[5].icell.SM XA.XIR[12].XIC[5].icell.Ien Iout.t19 VGND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X789 XA.XIR[7].XIC[2].icell.Ien XThR.Tn[7].t22 VPWR.t233 VPWR.t232 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X790 VGND.t1093 Vbias.t83 XA.XIR[3].XIC[13].icell.SM VGND.t1092 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X791 VGND.t1381 XThC.Tn[0].t20 XA.XIR[8].XIC[0].icell.PDM VGND.t1380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X792 VGND.t1760 XThC.Tn[12].t19 XA.XIR[3].XIC[12].icell.PDM VGND.t1759 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X793 XThR.XTB3.Y.t2 XThR.XTB7.A VPWR.t1889 VPWR.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X794 XA.XIR[15].XIC[6].icell.SM XA.XIR[15].XIC[6].icell.Ien Iout.t183 VGND.t1771 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X795 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[12].t32 XA.XIR[12].XIC[1].icell.Ien VGND.t308 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X796 VGND.t2301 XThC.Tn[13].t22 XA.XIR[6].XIC[13].icell.PDM VGND.t2300 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X797 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[7].t23 XA.XIR[7].XIC[5].icell.Ien VGND.t380 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X798 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t1970 VGND.t748 VGND.t747 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X799 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t6 VGND.t1749 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X800 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[14].t26 XA.XIR[14].XIC[3].icell.Ien VGND.t2125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X801 XA.XIR[10].XIC[8].icell.PUM XThC.Tn[8].t20 XA.XIR[10].XIC[8].icell.Ien VPWR.t1267 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X802 XA.XIR[1].XIC[12].icell.Ien XThR.Tn[1].t28 VPWR.t511 VPWR.t510 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X803 VGND.t1095 Vbias.t84 XA.XIR[2].XIC[11].icell.SM VGND.t1094 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X804 XA.XIR[6].XIC_15.icell.SM XA.XIR[6].XIC_15.icell.Ien Iout.t87 VGND.t1099 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X805 XA.XIR[0].XIC[0].icell.Ien XThR.Tn[0].t32 VPWR.t789 VPWR.t788 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X806 XThR.Tn[0].t8 XThR.XTBN.Y.t35 VGND.t550 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X807 VPWR.t1895 XThR.XTB5.Y a_n1049_6405# VPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X808 XA.XIR[4].XIC[13].icell.Ien XThR.Tn[4].t31 VPWR.t908 VPWR.t907 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X809 VGND.t227 Vbias.t85 XA.XIR[14].XIC_15.icell.SM VGND.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X810 XA.XIR[9].XIC[4].icell.SM XA.XIR[9].XIC[4].icell.Ien Iout.t149 VGND.t1519 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X811 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[10].t29 XA.XIR[10].XIC[0].icell.Ien VGND.t1921 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X812 XThC.Tn[10].t0 XThC.XTB3.Y.t4 VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X813 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[5].t28 XA.XIR[5].XIC[12].icell.Ien VGND.t163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X814 VPWR.t375 XThR.XTBN.Y.t36 XThR.Tn[10].t5 VPWR.t374 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X815 XA.XIR[8].XIC_dummy_right.icell.SM XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout VGND.t1534 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X816 VPWR.t67 XThR.Tn[11].t29 XA.XIR[12].XIC[4].icell.PUM VPWR.t66 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X817 VPWR.t268 XThC.XTBN.Y.t36 XThC.Tn[13].t9 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X818 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[9].t29 XA.XIR[9].XIC[12].icell.Ien VGND.t519 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X819 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[8].t34 XA.XIR[8].XIC[13].icell.Ien VGND.t473 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X820 a_3773_9615# XThC.XTB2.Y VPWR.t106 VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X821 XThC.Tn[5].t1 XThC.XTB6.Y VGND.t1396 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X822 XA.XIR[4].XIC[2].icell.SM XA.XIR[4].XIC[2].icell.Ien Iout.t208 VGND.t1958 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X823 XThC.Tn[2].t0 XThC.XTB3.Y.t5 VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X824 VPWR.t750 XThR.Tn[3].t30 XA.XIR[4].XIC[6].icell.PUM VPWR.t749 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X825 VPWR.t1082 XThR.Tn[2].t27 XA.XIR[3].XIC[7].icell.PUM VPWR.t1081 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X826 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[12].t33 VGND.t310 VGND.t309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X827 VGND.t2573 XThC.Tn[10].t20 XA.XIR[3].XIC[10].icell.PDM VGND.t2572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X828 VPWR.t1900 XThR.Tn[6].t25 XA.XIR[7].XIC[7].icell.PUM VPWR.t1899 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X829 XA.XIR[15].XIC[10].icell.SM XA.XIR[15].XIC[10].icell.Ien Iout.t167 VGND.t1616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X830 VPWR.t65 XThR.Tn[5].t29 XA.XIR[6].XIC[8].icell.PUM VPWR.t64 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X831 VGND.t552 XThR.XTBN.Y.t37 a_n997_3755# VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X832 XA.XIR[2].XIC[5].icell.PUM XThC.Tn[5].t18 XA.XIR[2].XIC[5].icell.Ien VPWR.t1338 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X833 VPWR.t1830 XThC.XTB1.Y.t6 a_2979_9615# VPWR.t1829 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[9].t30 VGND.t521 VGND.t520 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X835 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t1971 VGND.t750 VGND.t749 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X836 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[14].t27 XA.XIR[14].XIC[7].icell.Ien VGND.t2126 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X837 XA.XIR[1].XIC[10].icell.Ien XThR.Tn[1].t29 VPWR.t513 VPWR.t512 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X838 VGND.t229 Vbias.t86 XA.XIR[2].XIC[9].icell.SM VGND.t228 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X839 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[12].t34 VGND.t394 VGND.t393 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X840 XA.XIR[12].XIC[0].icell.SM XA.XIR[12].XIC[0].icell.Ien Iout.t64 VGND.t803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X841 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[11].t30 VGND.t173 VGND.t172 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X842 XA.XIR[3].XIC_15.icell.SM XA.XIR[3].XIC_15.icell.Ien Iout.t26 VGND.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X843 XA.XIR[11].XIC_dummy_left.icell.SM XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout VGND.t639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X844 XA.XIR[7].XIC[12].icell.SM XA.XIR[7].XIC[12].icell.Ien Iout.t120 VGND.t1306 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X845 XA.XIR[14].XIC[12].icell.PUM XThC.Tn[12].t20 XA.XIR[14].XIC[12].icell.Ien VPWR.t955 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X846 XA.XIR[15].XIC[1].icell.SM XA.XIR[15].XIC[1].icell.Ien Iout.t0 VGND.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X847 VGND.t851 XThC.Tn[11].t20 XA.XIR[15].XIC[11].icell.PDM VGND.t850 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X848 XA.XIR[11].XIC_15.icell.PDM VPWR.t1972 VGND.t752 VGND.t751 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X849 XA.XIR[10].XIC[13].icell.SM XA.XIR[10].XIC[13].icell.Ien Iout.t138 VGND.t1430 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X850 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[5].t30 XA.XIR[5].XIC[10].icell.Ien VGND.t164 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X851 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[7].t24 XA.XIR[7].XIC[0].icell.Ien VGND.t381 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X852 XA.XIR[13].XIC[14].icell.SM XA.XIR[13].XIC[14].icell.Ien Iout.t17 VGND.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X853 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[9].t31 XA.XIR[9].XIC[10].icell.Ien VGND.t522 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X854 XA.XIR[10].XIC[3].icell.PUM XThC.Tn[3].t21 XA.XIR[10].XIC[3].icell.Ien VPWR.t140 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X855 a_5155_9615# XThC.XTB5.Y VPWR.t165 VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X856 XA.XIR[5].XIC_15.icell.PUM VPWR.t1686 XA.XIR[5].XIC_15.icell.Ien VPWR.t1687 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X857 VPWR.t69 XThR.Tn[11].t31 XA.XIR[12].XIC[0].icell.PUM VPWR.t68 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X858 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[6].t26 VGND.t2658 VGND.t2657 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X859 a_n1049_7493# XThR.XTB3.Y.t7 VPWR.t1888 VPWR.t1176 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X860 VGND.t2325 XThC.Tn[1].t23 XA.XIR[12].XIC[1].icell.PDM VGND.t2324 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X861 XA.XIR[9].XIC_15.icell.PUM VPWR.t1684 XA.XIR[9].XIC_15.icell.Ien VPWR.t1685 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X862 VGND.t1628 XThC.Tn[2].t20 XA.XIR[15].XIC[2].icell.PDM VGND.t1627 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X863 VPWR.t1080 XThR.Tn[2].t28 XA.XIR[3].XIC[11].icell.PUM VPWR.t1079 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X864 VPWR.t1902 XThR.Tn[6].t27 XA.XIR[7].XIC[11].icell.PUM VPWR.t1901 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X865 VGND.t754 VPWR.t1973 XA.XIR[13].XIC_15.icell.PDM VGND.t753 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X866 XThC.Tn[8].t7 XThC.XTB1.Y.t7 VPWR.t1832 VPWR.t1831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X867 XA.XIR[4].XIC[6].icell.Ien XThR.Tn[4].t32 VPWR.t1144 VPWR.t1143 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X868 XA.XIR[3].XIC[7].icell.Ien XThR.Tn[3].t31 VPWR.t752 VPWR.t751 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X869 VGND.t2653 XThR.XTB5.Y XThR.Tn[4].t11 VGND.t264 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X870 a_5155_9615# XThC.XTBN.Y.t37 XThC.Tn[4].t11 VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X871 VGND.t756 VPWR.t1974 XA.XIR[0].XIC_dummy_right.icell.PDM VGND.t755 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X872 VPWR.t754 XThR.Tn[3].t32 XA.XIR[4].XIC[1].icell.PUM VPWR.t753 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X873 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[12].t35 VGND.t396 VGND.t395 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X874 VPWR.t1078 XThR.Tn[2].t29 XA.XIR[3].XIC[2].icell.PUM VPWR.t1077 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X875 XThR.XTB5.Y XThR.XTB5.A VGND.t1635 VGND.t1634 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X876 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[11].t32 VGND.t1105 VGND.t1104 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X877 VPWR.t1904 XThR.Tn[6].t28 XA.XIR[7].XIC[2].icell.PUM VPWR.t1903 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X878 VPWR.t515 XThR.Tn[1].t30 XA.XIR[2].XIC[14].icell.PUM VPWR.t514 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X879 VPWR.t859 XThR.Tn[5].t31 XA.XIR[6].XIC[3].icell.PUM VPWR.t858 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X880 XA.XIR[14].XIC[10].icell.PUM XThC.Tn[10].t21 XA.XIR[14].XIC[10].icell.Ien VPWR.t1850 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X881 XA.XIR[8].XIC_dummy_left.icell.SM XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout VGND.t1327 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X882 VPWR.t1675 VPWR.t1673 XA.XIR[1].XIC_15.icell.PUM VPWR.t1674 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X883 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[4].t33 XA.XIR[4].XIC[9].icell.Ien VGND.t1963 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X884 VPWR.t1683 VPWR.t1681 XA.XIR[5].XIC_15.icell.PUM VPWR.t1682 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X885 XA.XIR[15].XIC_15.icell.PDM VPWR.t1975 XA.XIR[15].XIC_15.icell.Ien VGND.t757 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X886 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[6].t29 VGND.t2660 VGND.t2659 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X887 XA.XIR[1].XIC[5].icell.Ien XThR.Tn[1].t31 VPWR.t517 VPWR.t516 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X888 VGND.t231 Vbias.t87 XA.XIR[2].XIC[4].icell.SM VGND.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X889 XA.XIR[6].XIC[8].icell.SM XA.XIR[6].XIC[8].icell.Ien Iout.t233 VGND.t2520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X890 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[2].t30 VGND.t774 VGND.t773 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X891 VGND.t233 Vbias.t88 XA.XIR[15].XIC[7].icell.SM VGND.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X892 VGND.t759 VPWR.t1976 XA.XIR[3].XIC_dummy_left.icell.PDM VGND.t758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X893 VGND.t235 Vbias.t89 XA.XIR[14].XIC[8].icell.SM VGND.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X894 VGND.t634 XThC.Tn[6].t23 XA.XIR[15].XIC[6].icell.PDM VGND.t633 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X895 VPWR.t1680 VPWR.t1678 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1679 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X896 XThC.Tn[14].t2 XThC.XTB7.Y a_10915_9569# VGND.t222 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X897 XThC.XTB3.Y.t1 XThC.XTB7.A a_4387_10575# VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X898 a_n997_1803# XThR.XTBN.Y.t38 VGND.t554 VGND.t553 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X899 XA.XIR[1].XIC[13].icell.PUM XThC.Tn[13].t23 XA.XIR[1].XIC[13].icell.Ien VPWR.t1355 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X900 XA.XIR[3].XIC[11].icell.Ien XThR.Tn[3].t33 VPWR.t756 VPWR.t755 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X901 XA.XIR[15].XIC[14].icell.PDM XThR.Tn[14].t28 VGND.t2128 VGND.t2127 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X902 a_3773_9615# XThC.XTBN.Y.t38 XThC.Tn[1].t11 VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X903 VGND.t2327 XThC.Tn[1].t24 XA.XIR[6].XIC[1].icell.PDM VGND.t2326 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X904 XA.XIR[14].XIC[6].icell.SM XA.XIR[14].XIC[6].icell.Ien Iout.t39 VGND.t266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X905 XA.XIR[15].XIC[8].icell.PDM XThR.Tn[14].t29 VGND.t2130 VGND.t2129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X906 VGND.t237 Vbias.t90 XA.XIR[5].XIC[14].icell.SM VGND.t236 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X907 VGND.t2303 XThC.Tn[13].t24 XA.XIR[5].XIC[13].icell.PDM VGND.t2302 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X908 VPWR.t761 XThC.XTB5.A XThC.XTB1.Y.t2 VPWR.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X909 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR.t1977 XA.XIR[5].XIC_dummy_left.icell.Ien VGND.t760 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X910 VGND.t2305 XThC.Tn[13].t25 XA.XIR[9].XIC[13].icell.PDM VGND.t2304 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X911 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t1978 XA.XIR[9].XIC_dummy_left.icell.Ien VGND.t761 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X912 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[1].t32 VGND.t836 VGND.t835 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X913 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[11].t33 XA.XIR[11].XIC[11].icell.Ien VGND.t1106 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X914 VGND.t239 Vbias.t91 XA.XIR[1].XIC[11].icell.SM VGND.t238 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X915 XA.XIR[4].XIC[1].icell.Ien XThR.Tn[4].t34 VPWR.t1146 VPWR.t1145 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X916 VGND.t241 Vbias.t92 XA.XIR[0].XIC[12].icell.SM VGND.t240 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X917 XA.XIR[3].XIC[2].icell.Ien XThR.Tn[3].t34 VPWR.t758 VPWR.t757 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X918 XA.XIR[12].XIC_15.icell.PDM XThR.Tn[12].t36 XA.XIR[12].XIC_15.icell.Ien VGND.t397 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X919 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1676 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR.t1677 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X920 XA.XIR[2].XIC[14].icell.Ien XThR.Tn[2].t31 VPWR.t1076 VPWR.t1075 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X921 XA.XIR[3].XIC[8].icell.SM XA.XIR[3].XIC[8].icell.Ien Iout.t251 VGND.t2648 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X922 VGND.t102 XThC.XTB3.Y.t6 XThC.Tn[2].t1 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X923 XA.XIR[14].XIC[5].icell.PUM XThC.Tn[5].t19 XA.XIR[14].XIC[5].icell.Ien VPWR.t1339 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X924 a_8739_9569# XThC.XTB3.Y.t7 XThC.Tn[10].t1 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X925 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[8].t35 XA.XIR[8].XIC[1].icell.Ien VGND.t474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X926 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[4].t35 XA.XIR[4].XIC[4].icell.Ien VGND.t1964 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X927 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[3].t35 XA.XIR[3].XIC[5].icell.Ien VGND.t1384 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X928 a_n1319_6405# XThR.XTB5.A VPWR.t927 VPWR.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X929 VPWR.t1254 XThR.Tn[14].t30 XA.XIR[15].XIC[4].icell.PUM VPWR.t1253 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X930 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[11].t34 XA.XIR[11].XIC[2].icell.Ien VGND.t1107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X931 XA.XIR[7].XIC[7].icell.PUM XThC.Tn[7].t16 XA.XIR[7].XIC[7].icell.Ien VPWR.t700 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X932 VPWR.t1667 VPWR.t1665 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1666 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X933 XA.XIR[6].XIC[3].icell.SM XA.XIR[6].XIC[3].icell.Ien Iout.t101 VGND.t1141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X934 a_2979_9615# XThC.XTB1.Y.t8 VPWR.t1834 VPWR.t1833 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X935 XA.XIR[0].XIC[13].icell.Ien XThR.Tn[0].t33 VPWR.t791 VPWR.t790 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X936 VGND.t243 Vbias.t93 XA.XIR[15].XIC[2].icell.SM VGND.t242 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X937 VGND.t245 Vbias.t94 XA.XIR[14].XIC[3].icell.SM VGND.t244 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X938 XThR.Tn[12].t2 XThR.XTBN.Y.t39 VPWR.t377 VPWR.t376 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X939 XA.XIR[4].XIC_dummy_right.icell.SM XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout VGND.t2536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X940 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1670 VPWR.t1672 VPWR.t1671 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X941 XA.XIR[14].XIC[10].icell.SM XA.XIR[14].XIC[10].icell.Ien Iout.t107 VGND.t1266 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X942 XThC.Tn[11].t7 XThC.XTBN.Y.t39 VPWR.t269 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X943 VGND.t1913 data[4].t2 XThR.XTB5.A VGND.t1912 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X944 XThR.XTBN.Y.t1 XThR.XTBN.A VGND.t1375 VGND.t1374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X945 VGND.t643 data[3].t0 XThC.XTBN.A VGND.t642 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X946 VGND.t247 Vbias.t95 XA.XIR[1].XIC[9].icell.SM VGND.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X947 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t1979 VGND.t763 VGND.t762 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X948 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[8].t36 VGND.t117 VGND.t116 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X949 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t7 VGND.t263 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X950 XA.XIR[15].XIC[3].icell.PDM XThR.Tn[14].t31 VGND.t2132 VGND.t2131 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X951 XA.XIR[14].XIC[1].icell.SM XA.XIR[14].XIC[1].icell.Ien Iout.t2 VGND.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X952 XA.XIR[10].XIC_15.icell.PDM VPWR.t1980 VGND.t765 VGND.t764 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X953 XA.XIR[9].XIC[13].icell.SM XA.XIR[9].XIC[13].icell.Ien Iout.t153 VGND.t1523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X954 a_n997_2667# XThR.XTBN.Y.t40 VGND.t555 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X955 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1668 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR.t1669 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X956 XA.XIR[12].XIC[14].icell.SM XA.XIR[12].XIC[14].icell.Ien Iout.t24 VGND.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X957 XA.XIR[1].XIC[6].icell.PUM XThC.Tn[6].t24 XA.XIR[1].XIC[6].icell.Ien VPWR.t437 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X958 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[1].t33 VGND.t838 VGND.t837 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X959 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[11].t35 XA.XIR[11].XIC[6].icell.Ien VGND.t1108 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X960 XA.XIR[7].XIC[11].icell.PUM XThC.Tn[11].t21 XA.XIR[7].XIC[11].icell.Ien VPWR.t536 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X961 XA.XIR[4].XIC[7].icell.PUM XThC.Tn[7].t17 XA.XIR[4].XIC[7].icell.Ien VPWR.t701 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X962 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[4].t36 VGND.t1966 VGND.t1965 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X963 VPWR.t1256 XThR.Tn[14].t32 XA.XIR[15].XIC[0].icell.PUM VPWR.t1255 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X964 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[8].t37 VGND.t119 VGND.t118 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X965 XA.XIR[3].XIC[8].icell.PUM XThC.Tn[8].t21 XA.XIR[3].XIC[8].icell.Ien VPWR.t1373 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X966 VGND.t1776 XThC.Tn[9].t23 XA.XIR[1].XIC[9].icell.PDM VGND.t1775 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X967 XA.XIR[3].XIC[3].icell.SM XA.XIR[3].XIC[3].icell.Ien Iout.t92 VGND.t1125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X968 XThC.Tn[4].t10 XThC.XTBN.Y.t40 a_5155_9615# VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X969 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[3].t36 XA.XIR[3].XIC[0].icell.Ien VGND.t1385 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X970 VGND.t2411 VPWR.t1981 XA.XIR[12].XIC_15.icell.PDM VGND.t2410 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X971 VPWR.t245 XThR.Tn[12].t37 XA.XIR[13].XIC[9].icell.PUM VPWR.t244 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X972 VPWR.t379 XThR.XTBN.Y.t41 XThR.Tn[8].t6 VPWR.t378 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X973 VGND.t197 XThC.Tn[14].t20 XA.XIR[11].XIC[14].icell.PDM VGND.t196 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X974 VGND.t2391 XThC.Tn[8].t22 XA.XIR[11].XIC[8].icell.PDM VGND.t2390 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X975 XA.XIR[7].XIC[2].icell.PUM XThC.Tn[2].t21 XA.XIR[7].XIC[2].icell.Ien VPWR.t921 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X976 XA.XIR[2].XIC[14].icell.PUM XThC.Tn[14].t21 XA.XIR[2].XIC[14].icell.Ien VPWR.t96 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X977 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1662 VPWR.t1664 VPWR.t1663 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X978 a_7651_9569# XThC.XTB1.Y.t9 XThC.Tn[8].t1 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X979 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[2].t32 XA.XIR[2].XIC[12].icell.Ien VGND.t772 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X980 VGND.t249 Vbias.t96 XA.XIR[4].XIC[5].icell.SM VGND.t248 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X981 VPWR.t164 XThC.XTB5.Y XThC.Tn[12].t5 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t1982 XA.XIR[14].XIC_dummy_right.icell.Ien VGND.t2412 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X983 VPWR.t629 XThR.Tn[11].t36 XA.XIR[12].XIC[13].icell.PUM VPWR.t628 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X984 VPWR.t1661 VPWR.t1659 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1660 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X985 VGND.t1716 Vbias.t97 XA.XIR[7].XIC[6].icell.SM VGND.t1715 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X986 XA.XIR[6].XIC[7].icell.Ien XThR.Tn[6].t30 VPWR.t1906 VPWR.t1905 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X987 XA.XIR[5].XIC[8].icell.Ien XThR.Tn[5].t32 VPWR.t861 VPWR.t860 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X988 VGND.t2263 XThC.Tn[5].t20 XA.XIR[7].XIC[5].icell.PDM VGND.t2262 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X989 VGND.t556 XThR.XTBN.Y.t42 XThR.Tn[1].t7 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X990 XA.XIR[15].XIC[7].icell.PDM XThR.Tn[14].t33 VGND.t1502 VGND.t1501 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X991 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[5].t33 VGND.t1561 VGND.t1560 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X992 XA.XIR[9].XIC[8].icell.Ien XThR.Tn[9].t32 VPWR.t339 VPWR.t338 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X993 VPWR.t592 VGND.t2692 XA.XIR[0].XIC[7].icell.PUM VPWR.t591 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X994 VPWR.t1658 VPWR.t1656 XA.XIR[4].XIC_15.icell.PUM VPWR.t1657 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X995 XA.XIR[0].XIC[6].icell.Ien XThR.Tn[0].t34 VPWR.t793 VPWR.t792 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X996 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[13].t28 XA.XIR[13].XIC[14].icell.Ien VGND.t1829 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X997 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[13].t29 XA.XIR[13].XIC[8].icell.Ien VGND.t1830 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X998 VGND.t1718 Vbias.t98 XA.XIR[1].XIC[4].icell.SM VGND.t1717 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X999 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[2].t33 VGND.t771 VGND.t770 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1000 XThR.Tn[6].t10 XThR.XTB7.Y VGND.t1748 VGND.t1747 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1001 a_9827_9569# XThC.XTBN.Y.t41 VGND.t418 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1002 XA.XIR[4].XIC[11].icell.PUM XThC.Tn[11].t22 XA.XIR[4].XIC[11].icell.Ien VPWR.t537 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1003 XThR.Tn[9].t1 XThR.XTBN.Y.t43 VPWR.t380 VPWR.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1004 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[8].t38 VGND.t121 VGND.t120 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1005 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[5].t34 VGND.t1563 VGND.t1562 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1006 XA.XIR[11].XIC[9].icell.PUM XThC.Tn[9].t24 XA.XIR[11].XIC[9].icell.Ien VPWR.t965 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1007 XA.XIR[4].XIC_dummy_left.icell.SM XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout VGND.t1953 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1008 XA.XIR[5].XIC[11].icell.SM XA.XIR[5].XIC[11].icell.Ien Iout.t154 VGND.t1524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1009 XA.XIR[0].XIC[9].icell.PDM XThR.Tn[0].t35 XA.XIR[0].XIC[9].icell.Ien VGND.t1452 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1010 XThC.Tn[1].t10 XThC.XTBN.Y.t42 a_3773_9615# VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1011 VGND.t853 XThC.Tn[11].t23 XA.XIR[8].XIC[11].icell.PDM VGND.t852 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1012 XThR.Tn[0].t7 XThR.XTBN.Y.t44 VGND.t604 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1013 XThC.Tn[13].t1 XThC.XTB6.Y a_10051_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1014 XA.XIR[1].XIC[1].icell.PUM XThC.Tn[1].t25 XA.XIR[1].XIC[1].icell.Ien VPWR.t1364 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1015 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[2].t34 XA.XIR[2].XIC[10].icell.Ien VGND.t769 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1016 XA.XIR[4].XIC[2].icell.PUM XThC.Tn[2].t22 XA.XIR[4].XIC[2].icell.Ien VPWR.t922 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1017 VPWR.t420 XThR.XTBN.Y.t45 XThR.Tn[10].t4 VPWR.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1018 VPWR.t341 XThR.Tn[9].t33 XA.XIR[10].XIC[9].icell.PUM VPWR.t340 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1019 XA.XIR[3].XIC[3].icell.PUM XThC.Tn[3].t22 XA.XIR[3].XIC[3].icell.Ien VPWR.t141 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1020 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[4].t37 VGND.t1968 VGND.t1967 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1021 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1653 VPWR.t1655 VPWR.t1654 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1022 XA.XIR[0].XIC[12].icell.PDM VGND.t989 VGND.t991 VGND.t990 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1023 VGND.t2106 XThC.Tn[4].t25 XA.XIR[1].XIC[4].icell.PDM VGND.t2105 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1024 VGND.t2329 XThC.Tn[1].t26 XA.XIR[5].XIC[1].icell.PDM VGND.t2328 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1025 VGND.t1720 Vbias.t99 XA.XIR[11].XIC[7].icell.SM VGND.t1719 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1026 VGND.t1722 Vbias.t100 XA.XIR[7].XIC[10].icell.SM VGND.t1721 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1027 XA.XIR[6].XIC[11].icell.Ien XThR.Tn[6].t31 VPWR.t1908 VPWR.t1907 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1028 VPWR.t117 XThC.XTB7.Y a_6243_9615# VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1029 XA.XIR[2].XIC[11].icell.SM XA.XIR[2].XIC[11].icell.Ien Iout.t213 VGND.t2144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1030 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t1983 VGND.t2414 VGND.t2413 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1031 VGND.t2331 XThC.Tn[1].t27 XA.XIR[9].XIC[1].icell.PDM VGND.t2330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1032 VGND.t2265 XThC.Tn[5].t21 XA.XIR[4].XIC[5].icell.PDM VGND.t2264 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1033 XA.XIR[13].XIC[9].icell.Ien XThR.Tn[13].t30 VPWR.t998 VPWR.t997 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1034 VGND.t1630 XThC.Tn[2].t23 XA.XIR[8].XIC[2].icell.PDM VGND.t1629 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1035 VPWR.t590 VGND.t2693 XA.XIR[0].XIC[11].icell.PUM VPWR.t589 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1036 VGND.t276 XThC.Tn[3].t23 XA.XIR[11].XIC[3].icell.PDM VGND.t275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1037 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[10].t30 XA.XIR[10].XIC[11].icell.Ien VGND.t1922 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1038 VGND.t2416 VPWR.t1984 XA.XIR[6].XIC_15.icell.PDM VGND.t2415 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1039 VGND.t1598 XThC.XTBN.Y.t43 a_8963_9569# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1040 VGND.t1724 Vbias.t101 XA.XIR[4].XIC[0].icell.SM VGND.t1723 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1041 XA.XIR[15].XIC[4].icell.PUM XThC.Tn[4].t26 XA.XIR[15].XIC[4].icell.Ien VPWR.t1221 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1042 VPWR.t857 XThR.XTB1.Y.t8 XThR.Tn[8].t10 VPWR.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1043 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR.t1651 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR.t1652 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1044 VGND.t1726 Vbias.t102 XA.XIR[7].XIC[1].icell.SM VGND.t1725 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1045 VGND.t1728 Vbias.t103 XA.XIR[2].XIC[13].icell.SM VGND.t1727 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1046 XA.XIR[6].XIC[2].icell.Ien XThR.Tn[6].t32 VPWR.t1910 VPWR.t1909 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1047 XA.XIR[11].XIC[5].icell.SM XA.XIR[11].XIC[5].icell.Ien Iout.t59 VGND.t645 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1048 VGND.t2086 XThC.Tn[0].t21 XA.XIR[7].XIC[0].icell.PDM VGND.t2085 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1049 XA.XIR[1].XIC[14].icell.Ien XThR.Tn[1].t34 VPWR.t519 VPWR.t518 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1050 XA.XIR[5].XIC[3].icell.Ien XThR.Tn[5].t35 VPWR.t863 VPWR.t862 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1051 VGND.t1762 XThC.Tn[12].t21 XA.XIR[2].XIC[12].icell.PDM VGND.t1761 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1052 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[5].t36 VGND.t1565 VGND.t1564 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1053 XThR.XTBN.A data[7].t0 VPWR.t1798 VPWR.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1054 XA.XIR[9].XIC[3].icell.Ien XThR.Tn[9].t34 VPWR.t343 VPWR.t342 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1055 XA.XIR[4].XIC_15.icell.Ien XThR.Tn[4].t38 VPWR.t1148 VPWR.t1147 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1056 XA.XIR[5].XIC[9].icell.SM XA.XIR[5].XIC[9].icell.Ien Iout.t142 VGND.t1451 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1057 a_6243_10571# XThC.XTB7.B XThC.XTB7.Y VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1058 VPWR.t588 VGND.t2694 XA.XIR[0].XIC[2].icell.PUM VPWR.t587 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1059 VPWR.t1172 XThR.XTB2.Y a_n1049_7787# VPWR.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1060 XA.XIR[10].XIC[2].icell.PDM XThR.Tn[10].t31 XA.XIR[10].XIC[2].icell.Ien VGND.t766 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1061 XA.XIR[6].XIC[5].icell.PDM XThR.Tn[6].t33 XA.XIR[6].XIC[5].icell.Ien VGND.t2661 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1062 XA.XIR[0].XIC[1].icell.Ien XThR.Tn[0].t36 VPWR.t662 VPWR.t661 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1063 XA.XIR[13].XIC[3].icell.PDM XThR.Tn[13].t31 XA.XIR[13].XIC[3].icell.Ien VGND.t1819 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1064 VPWR.t631 XThR.Tn[11].t37 XA.XIR[12].XIC[6].icell.PUM VPWR.t630 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1065 XA.XIR[8].XIC_15.icell.PDM XThR.Tn[8].t39 XA.XIR[8].XIC_15.icell.Ien VGND.t122 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1066 XA.XIR[0].XIC[7].icell.SM XA.XIR[0].XIC[7].icell.Ien Iout.t177 VGND.t1639 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1067 XA.XIR[0].XIC[10].icell.PDM VGND.t986 VGND.t988 VGND.t987 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1068 XA.XIR[0].XIC[4].icell.PDM XThR.Tn[0].t37 XA.XIR[0].XIC[4].icell.Ien VGND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1069 VGND.t1730 Vbias.t104 XA.XIR[8].XIC[7].icell.SM VGND.t1729 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1070 a_n1049_7493# XThR.XTBN.Y.t46 XThR.Tn[2].t6 VPWR.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1071 XA.XIR[2].XIC[9].icell.SM XA.XIR[2].XIC[9].icell.Ien Iout.t61 VGND.t647 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1072 VGND.t636 XThC.Tn[6].t25 XA.XIR[8].XIC[6].icell.PDM VGND.t635 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1073 XThC.Tn[8].t6 XThC.XTB1.Y.t10 VPWR.t1836 VPWR.t1835 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1074 VPWR.t477 XThR.Tn[10].t32 XA.XIR[11].XIC[4].icell.PUM VPWR.t476 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1075 VPWR.t1650 VPWR.t1648 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1649 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1076 VGND.t985 VGND.t983 XA.XIR[15].XIC_dummy_right.icell.SM VGND.t984 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1077 VGND.t1274 XThC.Tn[7].t18 XA.XIR[11].XIC[7].icell.PDM VGND.t1273 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1078 XThR.Tn[0].t10 XThR.XTB1.Y.t9 VGND.t1559 VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1079 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[7].t25 XA.XIR[7].XIC[11].icell.Ien VGND.t382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1080 VGND.t1732 Vbias.t105 XA.XIR[11].XIC[2].icell.SM VGND.t1731 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1081 XA.XIR[15].XIC[0].icell.PUM XThC.Tn[0].t22 XA.XIR[15].XIC[0].icell.Ien VPWR.t1214 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1082 VPWR.t1319 XThR.XTB3.Y.t8 XThR.Tn[10].t7 VPWR.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1083 VGND.t2575 XThC.Tn[10].t22 XA.XIR[2].XIC[10].icell.PDM VGND.t2574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1084 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[7].t26 VGND.t384 VGND.t383 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1085 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[7].t27 VGND.t386 VGND.t385 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1086 XA.XIR[8].XIC[5].icell.SM XA.XIR[8].XIC[5].icell.Ien Iout.t240 VGND.t2539 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1087 VPWR.t105 XThC.XTB2.Y a_3773_9615# VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1088 VGND.t2088 XThC.Tn[0].t23 XA.XIR[4].XIC[0].icell.PDM VGND.t2087 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1089 VGND.t605 XThR.XTBN.Y.t47 XThR.Tn[4].t6 VGND.t543 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1090 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1646 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR.t1647 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1091 XA.XIR[7].XIC[6].icell.SM XA.XIR[7].XIC[6].icell.Ien Iout.t33 VGND.t211 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1092 XA.XIR[14].XIC[14].icell.PUM XThC.Tn[14].t22 XA.XIR[14].XIC[14].icell.Ien VPWR.t97 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1093 XA.XIR[10].XIC[6].icell.PDM XThR.Tn[10].t33 XA.XIR[10].XIC[6].icell.Ien VGND.t767 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1094 VPWR.t889 XThC.XTBN.Y.t44 XThC.Tn[9].t11 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t1985 XA.XIR[2].XIC_dummy_left.icell.Ien VGND.t2417 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1096 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[7].t28 XA.XIR[7].XIC[2].icell.Ien VGND.t387 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1097 VGND.t1599 XThC.XTBN.Y.t45 XThC.Tn[5].t5 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1098 XA.XIR[4].XIC[5].icell.PDM XThR.Tn[3].t37 VGND.t1387 VGND.t1386 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1099 XA.XIR[13].XIC[7].icell.PDM XThR.Tn[13].t32 XA.XIR[13].XIC[7].icell.Ien VGND.t1820 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1100 XA.XIR[11].XIC[0].icell.SM XA.XIR[11].XIC[0].icell.Ien Iout.t99 VGND.t1139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1101 XA.XIR[6].XIC[12].icell.SM XA.XIR[6].XIC[12].icell.Ien Iout.t188 VGND.t1791 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1102 VGND.t606 XThR.XTBN.Y.t48 a_n997_1579# VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1103 XA.XIR[13].XIC[12].icell.PUM XThC.Tn[12].t22 XA.XIR[13].XIC[12].icell.Ien VPWR.t956 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1104 XA.XIR[5].XIC[4].icell.SM XA.XIR[5].XIC[4].icell.Ien Iout.t1 VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1105 VGND.t1734 Vbias.t106 XA.XIR[14].XIC[12].icell.SM VGND.t1733 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1106 VGND.t1736 Vbias.t107 XA.XIR[10].XIC_15.icell.SM VGND.t1735 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1107 a_2979_9615# XThC.XTBN.Y.t46 XThC.Tn[0].t4 VPWR.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1108 VGND.t199 XThC.Tn[14].t23 XA.XIR[10].XIC[14].icell.PDM VGND.t198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1109 XA.XIR[6].XIC[0].icell.PDM XThR.Tn[6].t34 XA.XIR[6].XIC[0].icell.Ien VGND.t2662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1110 VGND.t2393 XThC.Tn[8].t23 XA.XIR[10].XIC[8].icell.PDM VGND.t2392 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1111 XA.XIR[1].XIC[12].icell.PDM XThR.Tn[1].t35 XA.XIR[1].XIC[12].icell.Ien VGND.t2676 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1112 VPWR.t633 XThR.Tn[11].t38 XA.XIR[12].XIC[1].icell.PUM VPWR.t632 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1113 XA.XIR[0].XIC[7].icell.PUM XThC.Tn[7].t19 XA.XIR[0].XIC[7].icell.Ien VPWR.t702 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1114 XThC.Tn[12].t2 XThC.XTB5.Y a_9827_9569# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1115 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[4].t39 XA.XIR[4].XIC[13].icell.Ien VGND.t1706 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1116 VPWR.t479 XThR.Tn[10].t34 XA.XIR[11].XIC[0].icell.PUM VPWR.t478 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1117 XThR.XTB6.A data[5].t2 VPWR.t155 VPWR.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1118 XA.XIR[0].XIC[2].icell.SM XA.XIR[0].XIC[2].icell.Ien Iout.t74 VGND.t865 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1119 VPWR.t1645 VPWR.t1643 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1644 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1120 XThR.Tn[14].t5 XThR.XTB7.Y a_n997_715# VGND.t1746 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1121 VPWR.t822 XThR.Tn[14].t34 XA.XIR[15].XIC[13].icell.PUM VPWR.t821 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1122 a_n1049_5317# XThR.XTBN.Y.t49 XThR.Tn[6].t3 VPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1123 XA.XIR[11].XIC[4].icell.Ien XThR.Tn[11].t39 VPWR.t1024 VPWR.t1023 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1124 VGND.t1738 Vbias.t108 XA.XIR[8].XIC[2].icell.SM VGND.t1737 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1125 XA.XIR[2].XIC[4].icell.SM XA.XIR[2].XIC[4].icell.Ien Iout.t109 VGND.t1268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1126 XA.XIR[15].XIC[12].icell.Ien VPWR.t1640 VPWR.t1642 VPWR.t1641 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1127 XA.XIR[7].XIC[10].icell.SM XA.XIR[7].XIC[10].icell.Ien Iout.t210 VGND.t1988 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1128 XA.XIR[15].XIC[7].icell.SM XA.XIR[15].XIC[7].icell.Ien Iout.t63 VGND.t680 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1129 VPWR.t1917 XThR.Tn[1].t36 XA.XIR[2].XIC[8].icell.PUM VPWR.t1916 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1130 VPWR.t43 XThR.Tn[8].t40 XA.XIR[9].XIC[12].icell.PUM VPWR.t42 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1131 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[7].t29 XA.XIR[7].XIC[6].icell.Ien VGND.t1067 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1132 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t1986 VGND.t2419 VGND.t2418 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1133 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[0].t38 VGND.t1147 VGND.t1146 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1134 XA.XIR[10].XIC[9].icell.PUM XThC.Tn[9].t25 XA.XIR[10].XIC[9].icell.Ien VPWR.t966 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1135 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[7].t30 VGND.t1069 VGND.t1068 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1136 XA.XIR[8].XIC[0].icell.SM XA.XIR[8].XIC[0].icell.Ien Iout.t13 VGND.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1137 XA.XIR[3].XIC[12].icell.SM XA.XIR[3].XIC[12].icell.Ien Iout.t10 VGND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1138 XA.XIR[3].XIC_15.icell.PDM VPWR.t1987 VGND.t2421 VGND.t2420 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1139 XA.XIR[13].XIC[10].icell.PUM XThC.Tn[10].t23 XA.XIR[13].XIC[10].icell.Ien VPWR.t1851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1140 XA.XIR[7].XIC[1].icell.SM XA.XIR[7].XIC[1].icell.Ien Iout.t159 VGND.t1535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1141 a_6243_9615# XThC.XTB7.Y VPWR.t116 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1142 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR.t1638 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1639 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1143 VGND.t982 VGND.t980 XA.XIR[15].XIC_dummy_left.icell.SM VGND.t981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1144 XThC.Tn[10].t10 XThC.XTBN.Y.t47 VPWR.t891 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1145 XA.XIR[1].XIC[10].icell.PDM XThR.Tn[1].t37 XA.XIR[1].XIC[10].icell.Ien VGND.t2677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1146 XA.XIR[0].XIC[11].icell.PUM XThC.Tn[11].t24 XA.XIR[0].XIC[11].icell.Ien VPWR.t538 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1147 XA.XIR[4].XIC[0].icell.PDM XThR.Tn[3].t38 VGND.t1389 VGND.t1388 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1148 VGND.t1764 XThC.Tn[12].t23 XA.XIR[14].XIC[12].icell.PDM VGND.t1763 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1149 XA.XIR[1].XIC_15.icell.PUM VPWR.t1636 XA.XIR[1].XIC_15.icell.Ien VPWR.t1637 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1150 XThC.Tn[10].t2 XThC.XTB3.Y.t8 a_8739_9569# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1151 XA.XIR[2].XIC[13].icell.PDM XThR.Tn[1].t38 VGND.t2679 VGND.t2678 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1152 VGND.t221 XThC.XTB7.Y XThC.Tn[6].t3 VGND.t220 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1153 XA.XIR[1].XIC[11].icell.SM XA.XIR[1].XIC[11].icell.Ien Iout.t230 VGND.t2507 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1154 VGND.t2423 VPWR.t1988 XA.XIR[2].XIC_dummy_left.icell.PDM VGND.t2422 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1155 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t1989 VGND.t2425 VGND.t2424 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1156 XThR.Tn[11].t10 XThR.XTBN.Y.t50 VPWR.t423 VPWR.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1157 VGND.t278 XThC.Tn[3].t24 XA.XIR[10].XIC[3].icell.PDM VGND.t277 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1158 VPWR.t892 XThC.XTBN.Y.t48 XThC.Tn[12].t11 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1159 VGND.t2427 VPWR.t1990 XA.XIR[5].XIC_15.icell.PDM VGND.t2426 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1160 XA.XIR[15].XIC[10].icell.Ien VPWR.t1633 VPWR.t1635 VPWR.t1634 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1161 VGND.t1836 Vbias.t109 XA.XIR[13].XIC[11].icell.SM VGND.t1835 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1162 XA.XIR[12].XIC[12].icell.Ien XThR.Tn[12].t38 VPWR.t247 VPWR.t246 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1163 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11].t40 VPWR.t1026 VPWR.t1025 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1164 VGND.t2429 VPWR.t1991 XA.XIR[9].XIC_15.icell.PDM VGND.t2428 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1165 VPWR.t865 XThR.Tn[5].t37 XA.XIR[6].XIC[9].icell.PUM VPWR.t864 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1166 XA.XIR[0].XIC[2].icell.PUM XThC.Tn[2].t24 XA.XIR[0].XIC[2].icell.Ien VPWR.t923 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1167 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1630 VPWR.t1632 VPWR.t1631 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1168 VPWR.t45 XThR.Tn[8].t41 XA.XIR[9].XIC[10].icell.PUM VPWR.t44 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1169 VGND.t1838 Vbias.t110 XA.XIR[1].XIC[13].icell.SM VGND.t1837 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1170 VGND.t1840 Vbias.t111 XA.XIR[0].XIC[6].icell.SM VGND.t1839 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1171 VGND.t2267 XThC.Tn[5].t22 XA.XIR[0].XIC[5].icell.PDM VGND.t2266 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1172 VGND.t1842 Vbias.t112 XA.XIR[4].XIC[14].icell.SM VGND.t1841 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1173 VGND.t2525 XThC.XTB7.A XThC.XTB7.Y VGND.t2524 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1174 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[7].t31 VGND.t1071 VGND.t1070 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1175 XA.XIR[2].XIC[8].icell.Ien XThR.Tn[2].t35 VPWR.t1074 VPWR.t1073 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1176 VPWR.t1919 XThR.Tn[1].t39 XA.XIR[2].XIC[3].icell.PUM VPWR.t1918 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1177 a_n997_1803# XThR.XTB5.Y XThR.Tn[12].t6 VGND.t262 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1178 XA.XIR[15].XIC[2].icell.SM XA.XIR[15].XIC[2].icell.Ien Iout.t169 VGND.t1618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1179 a_n997_2667# XThR.XTBN.Y.t51 VGND.t607 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1180 VPWR.t824 XThR.Tn[14].t35 XA.XIR[15].XIC[6].icell.PUM VPWR.t823 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1181 VPWR.t1000 XThR.Tn[13].t33 XA.XIR[14].XIC[7].icell.PUM VPWR.t999 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1182 a_7875_9569# XThC.XTBN.Y.t49 VGND.t1600 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1183 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[0].t39 VGND.t1149 VGND.t1148 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1184 VGND.t2577 XThC.Tn[10].t24 XA.XIR[14].XIC[10].icell.PDM VGND.t2576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1185 VGND.t608 XThR.XTBN.Y.t52 a_n997_3979# VGND.t551 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1186 XA.XIR[0].XIC_15.icell.Ien XThR.Tn[0].t40 VPWR.t664 VPWR.t663 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1187 XA.XIR[1].XIC[9].icell.SM XA.XIR[1].XIC[9].icell.Ien Iout.t175 VGND.t1637 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1188 XA.XIR[13].XIC[5].icell.PUM XThC.Tn[5].t23 XA.XIR[13].XIC[5].icell.Ien VPWR.t1340 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1189 XThC.Tn[14].t10 XThC.XTBN.Y.t50 VPWR.t893 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1190 a_n1049_6699# XThR.XTB4.Y VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1191 a_4861_9615# XThC.XTBN.Y.t51 XThC.Tn[3].t7 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1192 VGND.t1844 Vbias.t113 XA.XIR[10].XIC[8].icell.SM VGND.t1843 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1193 VGND.t1276 XThC.Tn[7].t20 XA.XIR[10].XIC[7].icell.PDM VGND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1194 VGND.t1846 Vbias.t114 XA.XIR[13].XIC[9].icell.SM VGND.t1845 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1195 XA.XIR[12].XIC[10].icell.Ien XThR.Tn[12].t39 VPWR.t249 VPWR.t248 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1196 XThC.Tn[2].t2 XThC.XTB3.Y.t9 VGND.t104 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1197 XThC.Tn[9].t10 XThC.XTBN.Y.t52 VPWR.t894 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1198 XThC.Tn[5].t4 XThC.XTBN.Y.t53 VGND.t1601 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1199 a_n1335_8107# XThR.XTB6.A XThR.XTB2.Y VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1200 VGND.t1848 Vbias.t115 XA.XIR[0].XIC[10].icell.SM VGND.t1847 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1201 XA.XIR[14].XIC[12].icell.PDM XThR.Tn[13].t34 VGND.t1822 VGND.t1821 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1202 VGND.t2307 XThC.Tn[13].t26 XA.XIR[1].XIC[13].icell.PDM VGND.t2306 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1203 XA.XIR[15].XIC[5].icell.Ien VPWR.t1627 VPWR.t1629 VPWR.t1628 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1204 VGND.t979 VGND.t977 XA.XIR[11].XIC_dummy_right.icell.SM VGND.t978 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1205 VPWR.t623 XThC.XTB1.Y.t11 a_2979_9615# VPWR.t622 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1206 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR.t1992 XA.XIR[1].XIC_dummy_left.icell.Ien VGND.t2430 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1207 XThC.Tn[0].t3 XThC.XTBN.Y.t54 a_2979_9615# VPWR.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1208 XA.XIR[3].XIC[11].icell.PDM XThR.Tn[3].t39 XA.XIR[3].XIC[11].icell.Ien VGND.t1390 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1209 VPWR.t47 XThR.Tn[8].t42 XA.XIR[9].XIC[5].icell.PUM VPWR.t46 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1210 VPWR.t1002 XThR.Tn[13].t35 XA.XIR[14].XIC[11].icell.PUM VPWR.t1001 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1211 XThR.Tn[12].t9 XThR.XTB5.Y VPWR.t1894 VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1212 XA.XIR[8].XIC[4].icell.PUM XThC.Tn[4].t27 XA.XIR[8].XIC[4].icell.Ien VPWR.t1222 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1213 XA.XIR[12].XIC[12].icell.PUM XThC.Tn[12].t24 XA.XIR[12].XIC[12].icell.Ien VPWR.t957 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1214 VGND.t1850 Vbias.t116 XA.XIR[0].XIC[1].icell.SM VGND.t1849 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1215 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR.t1625 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR.t1626 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1216 XA.XIR[4].XIC[5].icell.SM XA.XIR[4].XIC[5].icell.Ien Iout.t84 VGND.t888 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1217 VGND.t2090 XThC.Tn[0].t24 XA.XIR[0].XIC[0].icell.PDM VGND.t2089 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1218 XThR.Tn[6].t6 XThR.XTBN.Y.t53 VGND.t610 VGND.t609 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1219 a_n1049_5611# XThR.XTBN.Y.t54 XThR.Tn[5].t6 VPWR.t422 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1220 XA.XIR[15].XIC[13].icell.PUM XThC.Tn[13].t27 XA.XIR[15].XIC[13].icell.Ien VPWR.t1356 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1221 VGND.t612 XThR.XTBN.Y.t55 a_n997_2891# VGND.t611 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1222 VGND.t1586 XThR.XTB7.B XThR.XTB7.Y VGND.t1585 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1223 XA.XIR[2].XIC[3].icell.Ien XThR.Tn[2].t36 VPWR.t1072 VPWR.t1071 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1224 XA.XIR[11].XIC[14].icell.SM XA.XIR[11].XIC[14].icell.Ien Iout.t160 VGND.t1536 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1225 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[4].t40 XA.XIR[4].XIC[1].icell.Ien VGND.t1707 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1226 XA.XIR[3].XIC[2].icell.PDM XThR.Tn[3].t40 XA.XIR[3].XIC[2].icell.Ien VGND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1227 XA.XIR[14].XIC[7].icell.Ien XThR.Tn[14].t36 VPWR.t826 VPWR.t825 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1228 VPWR.t828 XThR.Tn[14].t37 XA.XIR[15].XIC[1].icell.PUM VPWR.t827 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1229 VGND.t2432 VPWR.t1993 XA.XIR[11].XIC_dummy_right.icell.PDM VGND.t2431 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1230 XA.XIR[2].XIC[8].icell.PUM XThC.Tn[8].t24 XA.XIR[2].XIC[8].icell.Ien VPWR.t1374 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1231 VPWR.t1194 XThR.Tn[13].t36 XA.XIR[14].XIC[2].icell.PUM VPWR.t1193 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1232 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t3 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1233 VPWR.t1624 VPWR.t1622 XA.XIR[12].XIC_15.icell.PUM VPWR.t1623 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1234 XA.XIR[1].XIC[4].icell.SM XA.XIR[1].XIC[4].icell.Ien Iout.t38 VGND.t253 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1235 XA.XIR[10].XIC[4].icell.Ien XThR.Tn[10].t35 VPWR.t481 VPWR.t480 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1236 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1619 VPWR.t1621 VPWR.t1620 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1237 VGND.t1852 Vbias.t117 XA.XIR[6].XIC_15.icell.SM VGND.t1851 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1238 XA.XIR[0].XIC_dummy_right.icell.SM XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout VGND.t1113 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1239 XA.XIR[14].XIC[7].icell.SM XA.XIR[14].XIC[7].icell.Ien Iout.t124 VGND.t1324 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1240 XA.XIR[14].XIC[10].icell.PDM XThR.Tn[13].t37 VGND.t2040 VGND.t2039 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1241 VGND.t1854 Vbias.t118 XA.XIR[10].XIC[3].icell.SM VGND.t1853 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1242 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1616 VPWR.t1618 VPWR.t1617 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1243 VGND.t1602 XThC.XTBN.Y.t55 XThC.Tn[1].t5 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1244 a_n1049_6405# XThR.XTB5.Y VPWR.t1893 VPWR.t82 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1245 VGND.t1856 Vbias.t119 XA.XIR[13].XIC[4].icell.SM VGND.t1855 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1246 XA.XIR[12].XIC[5].icell.Ien XThR.Tn[12].t40 VPWR.t251 VPWR.t250 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1247 VPWR.t607 XThR.Tn[7].t32 XA.XIR[8].XIC[12].icell.PUM VPWR.t606 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1248 XA.XIR[0].XIC[13].icell.PDM XThR.Tn[0].t41 XA.XIR[0].XIC[13].icell.Ien VGND.t1150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1249 VGND.t976 VGND.t974 XA.XIR[8].XIC_dummy_right.icell.SM VGND.t975 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1250 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR.t1994 XA.XIR[13].XIC_dummy_right.icell.Ien VGND.t2433 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1251 VGND.t2435 VPWR.t1995 XA.XIR[14].XIC_dummy_left.icell.PDM VGND.t2434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1252 VPWR.t483 XThR.Tn[10].t36 XA.XIR[11].XIC[13].icell.PUM VPWR.t482 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1253 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[4].t41 VGND.t1709 VGND.t1708 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1254 XA.XIR[12].XIC[10].icell.PUM XThC.Tn[10].t25 XA.XIR[12].XIC[10].icell.Ien VPWR.t1852 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1255 VPWR.t615 XThR.XTB1.Y.t10 XThR.Tn[8].t0 VPWR.t614 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1256 XA.XIR[8].XIC[0].icell.PUM XThC.Tn[0].t25 XA.XIR[8].XIC[0].icell.Ien VPWR.t1215 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1257 XA.XIR[5].XIC[13].icell.SM XA.XIR[5].XIC[13].icell.Ien Iout.t225 VGND.t2321 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1258 VPWR.t425 XThR.XTBN.Y.t56 XThR.Tn[7].t6 VPWR.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1259 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1614 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR.t1615 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1260 VGND.t209 XThC.XTB2.Y XThC.Tn[1].t3 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1261 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR.t1612 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR.t1613 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1262 XA.XIR[8].XIC[14].icell.SM XA.XIR[8].XIC[14].icell.Ien Iout.t114 VGND.t1290 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1263 XA.XIR[3].XIC[6].icell.PDM XThR.Tn[3].t41 XA.XIR[3].XIC[6].icell.Ien VGND.t1161 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1264 XThC.Tn[12].t10 XThC.XTBN.Y.t56 VPWR.t896 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 XA.XIR[2].XIC[1].icell.PDM XThR.Tn[1].t40 VGND.t2681 VGND.t2680 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1266 XA.XIR[14].XIC[11].icell.Ien XThR.Tn[14].t38 VPWR.t830 VPWR.t829 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1267 VGND.t1979 XThR.XTB2.Y XThR.Tn[1].t10 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1268 XThR.Tn[1].t2 XThR.XTBN.Y.t57 a_n1049_7787# VPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1269 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[4].t42 VGND.t1711 VGND.t1710 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1270 XA.XIR[4].XIC[0].icell.SM XA.XIR[4].XIC[0].icell.Ien Iout.t125 VGND.t1326 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1271 XA.XIR[6].XIC[12].icell.PUM XThC.Tn[12].t25 XA.XIR[6].XIC[12].icell.Ien VPWR.t958 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1272 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[12].t41 VGND.t399 VGND.t398 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1273 VGND.t855 XThC.Tn[11].t25 XA.XIR[7].XIC[11].icell.PDM VGND.t854 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1274 XA.XIR[2].XIC[13].icell.SM XA.XIR[2].XIC[13].icell.Ien Iout.t85 VGND.t889 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1275 XA.XIR[7].XIC[4].icell.Ien XThR.Tn[7].t33 VPWR.t609 VPWR.t608 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1276 VGND.t1858 Vbias.t120 XA.XIR[3].XIC_15.icell.SM VGND.t1857 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1277 VGND.t2621 Vbias.t121 XA.XIR[12].XIC[11].icell.SM VGND.t2620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1278 VGND.t973 VGND.t971 XA.XIR[11].XIC_dummy_left.icell.SM VGND.t972 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1279 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10].t37 VPWR.t485 VPWR.t484 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1280 VGND.t2395 XThC.Tn[8].t25 XA.XIR[3].XIC[8].icell.PDM VGND.t2394 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1281 VGND.t201 XThC.Tn[14].t24 XA.XIR[3].XIC[14].icell.PDM VGND.t200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1282 XA.XIR[14].XIC[2].icell.Ien XThR.Tn[14].t39 VPWR.t832 VPWR.t831 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1283 XThR.Tn[9].t9 XThR.XTB2.Y VPWR.t1171 VPWR.t1170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1284 XThR.Tn[7].t1 XThR.XTBN.Y.t58 VGND.t614 VGND.t613 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1285 VPWR.t1318 data[1].t2 XThC.XTB6.A VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1286 XA.XIR[2].XIC[3].icell.PUM XThC.Tn[3].t25 XA.XIR[2].XIC[3].icell.Ien VPWR.t770 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1287 VPWR.t611 XThR.Tn[7].t34 XA.XIR[8].XIC[10].icell.PUM VPWR.t610 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1288 XA.XIR[15].XIC[6].icell.PUM XThC.Tn[6].t26 XA.XIR[15].XIC[6].icell.Ien VPWR.t438 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1289 VPWR.t1611 VPWR.t1609 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1610 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1290 VGND.t435 XThC.XTBN.Y.t57 a_7875_9569# VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1291 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[14].t40 XA.XIR[14].XIC[5].icell.Ien VGND.t1503 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1292 VPWR.t426 XThR.XTBN.Y.t59 XThR.Tn[13].t10 VPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1293 XA.XIR[1].XIC[8].icell.Ien XThR.Tn[1].t41 VPWR.t1921 VPWR.t1920 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1294 VPWR.t1608 VPWR.t1606 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR.t1607 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1295 VGND.t1281 XThC.Tn[2].t25 XA.XIR[7].XIC[2].icell.PDM VGND.t1280 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1296 a_8739_10571# data[0].t1 XThC.XTB7.A VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1297 XA.XIR[14].XIC[2].icell.SM XA.XIR[14].XIC[2].icell.Ien Iout.t83 VGND.t886 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1298 VGND.t2623 Vbias.t122 XA.XIR[9].XIC[11].icell.SM VGND.t2622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1299 VPWR.t658 XThR.XTB3.Y.t9 XThR.Tn[10].t6 VPWR.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1300 XA.XIR[8].XIC[12].icell.Ien XThR.Tn[8].t43 VPWR.t521 VPWR.t520 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1301 VGND.t1778 XThC.Tn[9].t26 XA.XIR[15].XIC[9].icell.PDM VGND.t1777 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1302 XThC.Tn[3].t6 XThC.XTBN.Y.t58 a_4861_9615# VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1303 XA.XIR[5].XIC[8].icell.PDM XThR.Tn[5].t38 XA.XIR[5].XIC[8].icell.Ien VGND.t1566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1304 XA.XIR[5].XIC[14].icell.PDM XThR.Tn[5].t39 XA.XIR[5].XIC[14].icell.Ien VGND.t1567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1305 XA.XIR[11].XIC[13].icell.Ien XThR.Tn[11].t41 VPWR.t1028 VPWR.t1027 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1306 XThR.Tn[5].t2 XThR.XTB6.Y VGND.t261 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1307 XA.XIR[9].XIC[14].icell.PDM XThR.Tn[9].t35 XA.XIR[9].XIC[14].icell.Ien VGND.t526 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1308 XA.XIR[9].XIC[8].icell.PDM XThR.Tn[9].t36 XA.XIR[9].XIC[8].icell.Ien VGND.t527 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1309 VPWR.t879 XThR.XTB7.B XThR.XTB4.Y VPWR.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1310 XA.XIR[15].XIC_dummy_right.icell.SM XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout VGND.t1612 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1311 XA.XIR[3].XIC[9].icell.PUM XThC.Tn[9].t27 XA.XIR[3].XIC[9].icell.Ien VPWR.t967 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1312 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[4].t43 VGND.t1713 VGND.t1712 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1313 XA.XIR[12].XIC[5].icell.PUM XThC.Tn[5].t24 XA.XIR[12].XIC[5].icell.Ien VPWR.t1341 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1314 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR.t1996 VGND.t2437 VGND.t2436 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1315 XA.XIR[6].XIC[10].icell.PUM XThC.Tn[10].t26 XA.XIR[6].XIC[10].icell.Ien VPWR.t1853 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1316 XA.XIR[0].XIC_dummy_left.icell.SM XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout VGND.t1465 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1317 VGND.t2625 Vbias.t123 XA.XIR[12].XIC[9].icell.SM VGND.t2624 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1318 VGND.t857 XThC.Tn[11].t26 XA.XIR[4].XIC[11].icell.PDM VGND.t856 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1319 VPWR.t487 XThR.Tn[10].t38 XA.XIR[11].XIC[6].icell.PUM VPWR.t486 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1320 VGND.t970 VGND.t968 XA.XIR[8].XIC_dummy_left.icell.SM VGND.t969 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1321 XA.XIR[7].XIC[0].icell.Ien XThR.Tn[7].t35 VPWR.t613 VPWR.t612 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1322 a_n997_715# XThR.XTB7.Y XThR.Tn[14].t4 VGND.t1745 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1323 VGND.t2333 XThC.Tn[1].t28 XA.XIR[1].XIC[1].icell.PDM VGND.t2332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1324 VGND.t2627 Vbias.t124 XA.XIR[7].XIC[7].icell.SM VGND.t2626 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1325 XA.XIR[5].XIC[9].icell.Ien XThR.Tn[5].t40 VPWR.t1098 VPWR.t1097 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1326 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[12].t42 VGND.t401 VGND.t400 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1327 VGND.t477 XThC.Tn[6].t27 XA.XIR[7].XIC[6].icell.PDM VGND.t476 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1328 VGND.t2629 Vbias.t125 XA.XIR[6].XIC[8].icell.SM VGND.t2628 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1329 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[11].t42 VGND.t1860 VGND.t1859 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1330 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t1997 VGND.t2439 VGND.t2438 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1331 VGND.t1283 XThC.Tn[2].t26 XA.XIR[4].XIC[2].icell.PDM VGND.t1282 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1332 XA.XIR[9].XIC[9].icell.Ien XThR.Tn[9].t37 VPWR.t345 VPWR.t344 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1333 VGND.t1433 XThC.Tn[3].t26 XA.XIR[3].XIC[3].icell.PDM VGND.t1432 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1334 XA.XIR[14].XIC[8].icell.PUM XThC.Tn[8].t26 XA.XIR[14].XIC[8].icell.Ien VPWR.t1375 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1335 VGND.t2631 Vbias.t126 XA.XIR[9].XIC[9].icell.SM VGND.t2630 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1336 XA.XIR[8].XIC[10].icell.Ien XThR.Tn[8].t44 VPWR.t523 VPWR.t522 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1337 XA.XIR[10].XIC_15.icell.SM XA.XIR[10].XIC_15.icell.Ien Iout.t219 VGND.t2188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1338 VPWR.t931 XThR.Tn[7].t36 XA.XIR[8].XIC[5].icell.PUM VPWR.t930 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1339 XA.XIR[6].XIC[11].icell.PDM XThR.Tn[6].t35 XA.XIR[6].XIC[11].icell.Ien VGND.t2663 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1340 XA.XIR[15].XIC[1].icell.PUM XThC.Tn[1].t29 XA.XIR[15].XIC[1].icell.Ien VPWR.t1365 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1341 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[14].t41 XA.XIR[14].XIC[0].icell.Ien VGND.t1504 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1342 XA.XIR[7].XIC[14].icell.PDM XThR.Tn[6].t36 VGND.t2665 VGND.t2664 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1343 XA.XIR[7].XIC[8].icell.PDM XThR.Tn[6].t37 VGND.t2667 VGND.t2666 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1344 XA.XIR[1].XIC[3].icell.Ien XThR.Tn[1].t42 VPWR.t505 VPWR.t504 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1345 XA.XIR[6].XIC[6].icell.SM XA.XIR[6].XIC[6].icell.Ien Iout.t244 VGND.t2556 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1346 XA.XIR[13].XIC[14].icell.PUM XThC.Tn[14].t25 XA.XIR[13].XIC[14].icell.Ien VPWR.t1295 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1347 VGND.t2633 Vbias.t127 XA.XIR[15].XIC[5].icell.SM VGND.t2632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1348 VGND.t2635 Vbias.t128 XA.XIR[14].XIC[6].icell.SM VGND.t2634 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1349 VGND.t2108 XThC.Tn[4].t28 XA.XIR[15].XIC[4].icell.PDM VGND.t2107 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1350 XA.XIR[6].XIC[2].icell.PDM XThR.Tn[6].t38 XA.XIR[6].XIC[2].icell.Ien VGND.t2668 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1351 VGND.t2441 VPWR.t1998 XA.XIR[10].XIC_dummy_right.icell.PDM VGND.t2440 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1352 XA.XIR[5].XIC[3].icell.PDM XThR.Tn[5].t41 XA.XIR[5].XIC[3].icell.Ien VGND.t1901 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1353 XThC.Tn[1].t4 XThC.XTBN.Y.t59 VGND.t436 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1354 XA.XIR[9].XIC[3].icell.PDM XThR.Tn[9].t38 XA.XIR[9].XIC[3].icell.Ien VGND.t528 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1355 XA.XIR[4].XIC_15.icell.PDM XThR.Tn[4].t44 XA.XIR[4].XIC_15.icell.Ien VGND.t1714 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1356 VPWR.t1605 VPWR.t1603 XA.XIR[15].XIC_15.icell.PUM VPWR.t1604 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1357 XA.XIR[6].XIC[5].icell.PUM XThC.Tn[5].t25 XA.XIR[6].XIC[5].icell.Ien VPWR.t1342 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1358 XA.XIR[0].XIC[1].icell.PDM XThR.Tn[0].t42 XA.XIR[0].XIC[1].icell.Ien VGND.t1151 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1359 XA.XIR[11].XIC[6].icell.Ien XThR.Tn[11].t43 VPWR.t1030 VPWR.t1029 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1360 a_7875_9569# XThC.XTB2.Y XThC.Tn[9].t5 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1361 VPWR.t1070 XThR.Tn[2].t37 XA.XIR[3].XIC[4].icell.PUM VPWR.t1069 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1362 VGND.t2637 Vbias.t129 XA.XIR[3].XIC[8].icell.SM VGND.t2636 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1363 VGND.t479 XThC.Tn[6].t28 XA.XIR[4].XIC[6].icell.PDM VGND.t478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1364 XA.XIR[15].XIC[14].icell.Ien VPWR.t1600 VPWR.t1602 VPWR.t1601 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1365 VGND.t2639 Vbias.t130 XA.XIR[12].XIC[4].icell.SM VGND.t2638 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1366 VPWR.t489 XThR.Tn[10].t39 XA.XIR[11].XIC[1].icell.PUM VPWR.t488 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1367 VGND.t817 XThC.Tn[7].t21 XA.XIR[3].XIC[7].icell.PDM VGND.t816 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1368 VPWR.t1912 XThR.Tn[6].t39 XA.XIR[7].XIC[4].icell.PUM VPWR.t1911 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1369 VPWR.t1599 VPWR.t1597 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1598 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1370 XThR.Tn[13].t1 XThR.XTB6.Y a_n997_1579# VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1371 a_n1049_8581# XThR.XTBN.Y.t60 XThR.Tn[0].t3 VPWR.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1372 XA.XIR[15].XIC_dummy_left.icell.SM XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout VGND.t1924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1373 VPWR.t525 XThR.Tn[8].t45 XA.XIR[9].XIC[14].icell.PUM VPWR.t524 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1374 XA.XIR[11].XIC[9].icell.PDM XThR.Tn[11].t44 XA.XIR[11].XIC[9].icell.Ien VGND.t1861 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1375 XA.XIR[4].XIC[11].icell.PDM XThR.Tn[3].t42 VGND.t1163 VGND.t1162 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1376 VGND.t2641 Vbias.t131 XA.XIR[7].XIC[2].icell.SM VGND.t2640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1377 VGND.t2643 Vbias.t132 XA.XIR[6].XIC[3].icell.SM VGND.t2642 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1378 XA.XIR[6].XIC[10].icell.SM XA.XIR[6].XIC[10].icell.Ien Iout.t88 VGND.t1100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1379 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[11].t45 VGND.t1863 VGND.t1862 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1380 XA.XIR[3].XIC[6].icell.SM XA.XIR[3].XIC[6].icell.Ien Iout.t95 VGND.t1129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1381 XA.XIR[14].XIC[3].icell.PUM XThC.Tn[3].t27 XA.XIR[14].XIC[3].icell.Ien VPWR.t771 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1382 VGND.t343 Vbias.t133 XA.XIR[9].XIC[4].icell.SM VGND.t342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1383 XA.XIR[8].XIC[5].icell.Ien XThR.Tn[8].t46 VPWR.t527 VPWR.t526 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1384 VGND.t345 Vbias.t134 XA.XIR[14].XIC[10].icell.SM VGND.t344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1385 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[10].t40 VGND.t2562 VGND.t2561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1386 XA.XIR[6].XIC[6].icell.PDM XThR.Tn[6].t40 XA.XIR[6].XIC[6].icell.Ien VGND.t2398 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1387 VGND.t1439 data[2].t1 XThC.XTB7.B VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1388 XA.XIR[5].XIC[7].icell.PDM XThR.Tn[5].t42 XA.XIR[5].XIC[7].icell.Ien VGND.t1902 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1389 VGND.t312 XThR.XTBN.Y.t61 XThR.Tn[2].t1 VGND.t311 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1390 XA.XIR[4].XIC[2].icell.PDM XThR.Tn[3].t43 VGND.t1165 VGND.t1164 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1391 XA.XIR[13].XIC[11].icell.SM XA.XIR[13].XIC[11].icell.Ien Iout.t220 VGND.t2195 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1392 a_n1049_5317# XThR.XTB7.Y VPWR.t944 VPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1393 XA.XIR[9].XIC[7].icell.PDM XThR.Tn[9].t39 XA.XIR[9].XIC[7].icell.Ien VGND.t529 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1394 VGND.t437 XThC.XTBN.Y.t60 XThC.Tn[4].t5 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1395 XA.XIR[5].XIC[12].icell.PUM XThC.Tn[12].t26 XA.XIR[5].XIC[12].icell.Ien VPWR.t959 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1396 XA.XIR[7].XIC[3].icell.PDM XThR.Tn[6].t41 VGND.t2400 VGND.t2399 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1397 XA.XIR[2].XIC_15.icell.PDM VPWR.t1999 VGND.t2443 VGND.t2442 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1398 XA.XIR[6].XIC[1].icell.SM XA.XIR[6].XIC[1].icell.Ien Iout.t128 VGND.t1339 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1399 XA.XIR[1].XIC[13].icell.SM XA.XIR[1].XIC[13].icell.Ien Iout.t252 VGND.t2649 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1400 XA.XIR[9].XIC[12].icell.PUM XThC.Tn[12].t27 XA.XIR[9].XIC[12].icell.Ien VPWR.t960 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1401 VGND.t347 Vbias.t135 XA.XIR[15].XIC[0].icell.SM VGND.t346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1402 XA.XIR[8].XIC[13].icell.PUM XThC.Tn[13].t28 XA.XIR[8].XIC[13].icell.Ien VPWR.t1357 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1403 VGND.t349 Vbias.t136 XA.XIR[14].XIC[1].icell.SM VGND.t348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1404 VGND.t351 Vbias.t137 XA.XIR[10].XIC[12].icell.SM VGND.t350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1405 XA.XIR[4].XIC[14].icell.SM XA.XIR[4].XIC[14].icell.Ien Iout.t44 VGND.t293 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1406 XThR.Tn[3].t2 XThR.XTB4.Y VGND.t189 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1407 VGND.t353 Vbias.t138 XA.XIR[13].XIC[13].icell.SM VGND.t352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1408 VPWR.t1068 XThR.Tn[2].t38 XA.XIR[3].XIC[0].icell.PUM VPWR.t1067 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1409 VGND.t1766 XThC.Tn[12].t28 XA.XIR[13].XIC[12].icell.PDM VGND.t1765 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1410 XA.XIR[12].XIC[14].icell.Ien XThR.Tn[12].t43 VPWR.t253 VPWR.t252 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1411 VPWR.t1377 XThR.Tn[6].t42 XA.XIR[7].XIC[0].icell.PUM VPWR.t1376 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1412 VPWR.t115 XThC.XTB7.Y a_6243_9615# VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 VPWR.t767 XThC.XTB6.Y XThC.Tn[13].t6 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1414 VPWR.t1596 VPWR.t1594 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1595 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1415 VGND.t1126 data[1].t3 XThC.XTB5.A VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1416 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[0].t43 VGND.t1342 VGND.t1341 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1417 XA.XIR[3].XIC[4].icell.Ien XThR.Tn[3].t44 VPWR.t672 VPWR.t671 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1418 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[8].t47 VGND.t840 VGND.t839 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1419 Vbias.t11 bias[2].t0 VPWR.t1797 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.1955 pd=1.31 as=0.2465 ps=2.28 w=0.85 l=0.5
X1420 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11].t46 VPWR.t1885 VPWR.t1884 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1421 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1591 VPWR.t1593 VPWR.t1592 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1422 VGND.t355 Vbias.t139 XA.XIR[3].XIC[3].icell.SM VGND.t354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1423 XA.XIR[7].XIC[7].icell.SM XA.XIR[7].XIC[7].icell.Ien Iout.t86 VGND.t1042 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1424 XA.XIR[3].XIC[10].icell.SM XA.XIR[3].XIC[10].icell.Ien Iout.t195 VGND.t1803 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1425 XA.XIR[10].XIC[13].icell.Ien XThR.Tn[10].t41 VPWR.t1840 VPWR.t1839 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1426 VPWR.t732 XThR.Tn[0].t44 XA.XIR[1].XIC[12].icell.PUM VPWR.t731 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1427 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[10].t42 VGND.t2564 VGND.t2563 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1428 XA.XIR[14].XIC_dummy_right.icell.SM XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout VGND.t887 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1429 XA.XIR[10].XIC[8].icell.SM XA.XIR[10].XIC[8].icell.Ien Iout.t215 VGND.t2146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1430 VGND.t439 XThC.XTBN.Y.t61 XThC.Tn[7].t2 VGND.t438 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1431 XA.XIR[4].XIC[6].icell.PDM XThR.Tn[3].t45 VGND.t1167 VGND.t1166 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1432 VPWR.t929 XThR.Tn[4].t45 XA.XIR[5].XIC[12].icell.PUM VPWR.t928 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1433 XA.XIR[11].XIC[4].icell.PDM XThR.Tn[11].t47 XA.XIR[11].XIC[4].icell.Ien VGND.t2608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1434 XA.XIR[13].XIC[9].icell.SM XA.XIR[13].XIC[9].icell.Ien Iout.t108 VGND.t1267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1435 XA.XIR[15].XIC[12].icell.PDM VPWR.t2000 XA.XIR[15].XIC[12].icell.Ien VGND.t2444 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1436 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[0].t45 VGND.t1344 VGND.t1343 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1437 XA.XIR[5].XIC[10].icell.PUM XThC.Tn[10].t27 XA.XIR[5].XIC[10].icell.Ien VPWR.t1854 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1438 XThR.Tn[12].t8 XThR.XTB5.Y VPWR.t1892 VPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1439 XA.XIR[7].XIC[7].icell.PDM XThR.Tn[6].t43 VGND.t2402 VGND.t2401 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1440 a_10915_9569# XThC.XTBN.Y.t62 VGND.t441 VGND.t440 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1441 XA.XIR[3].XIC[1].icell.SM XA.XIR[3].XIC[1].icell.Ien Iout.t165 VGND.t1614 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1442 XA.XIR[9].XIC[10].icell.PUM XThC.Tn[10].t28 XA.XIR[9].XIC[10].icell.Ien VPWR.t1855 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1443 XThR.Tn[6].t5 XThR.XTBN.Y.t62 VGND.t314 VGND.t313 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1444 VPWR.t255 XThR.Tn[12].t44 XA.XIR[13].XIC[7].icell.PUM VPWR.t254 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1445 XThC.Tn[3].t10 XThC.XTB4.Y.t7 VGND.t1909 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1446 XThC.Tn[9].t1 XThC.XTB2.Y VPWR.t104 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1447 VGND.t2579 XThC.Tn[10].t29 XA.XIR[13].XIC[10].icell.PDM VGND.t2578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1448 a_n997_2667# XThR.XTB4.Y XThR.Tn[11].t2 VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1449 VGND.t859 XThC.Tn[11].t27 XA.XIR[0].XIC[11].icell.PDM VGND.t858 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1450 XA.XIR[15].XIC[5].icell.PDM XThR.Tn[14].t42 VGND.t1506 VGND.t1505 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1451 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[5].t43 VGND.t1904 VGND.t1903 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1452 VGND.t357 Vbias.t140 XA.XIR[5].XIC[11].icell.SM VGND.t356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1453 XA.XIR[3].XIC[0].icell.Ien XThR.Tn[3].t46 VPWR.t674 VPWR.t673 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1454 XA.XIR[9].XIC_15.icell.SM XA.XIR[9].XIC_15.icell.Ien Iout.t75 VGND.t866 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1455 VGND.t2446 VPWR.t2001 XA.XIR[1].XIC_15.icell.PDM VGND.t2445 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1456 VPWR.t507 XThR.Tn[1].t43 XA.XIR[2].XIC[9].icell.PUM VPWR.t506 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1457 VPWR.t734 XThR.Tn[0].t46 XA.XIR[1].XIC[10].icell.PUM VPWR.t733 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1458 XA.XIR[7].XIC[13].icell.Ien XThR.Tn[7].t37 VPWR.t933 VPWR.t932 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1459 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1588 VPWR.t1590 VPWR.t1589 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1460 VPWR.t143 XThR.Tn[4].t46 XA.XIR[5].XIC[10].icell.PUM VPWR.t142 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1461 XA.XIR[15].XIC[10].icell.PDM VPWR.t2002 XA.XIR[15].XIC[10].icell.Ien VGND.t2447 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1462 XA.XIR[12].XIC[14].icell.PUM XThC.Tn[14].t26 XA.XIR[12].XIC[14].icell.Ien VPWR.t1296 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1463 XA.XIR[8].XIC[6].icell.PUM XThC.Tn[6].t29 XA.XIR[8].XIC[6].icell.Ien VPWR.t300 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1464 VGND.t1584 XThR.XTB7.B a_n1335_8331# VGND.t1583 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1465 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[0].t47 VGND.t1346 VGND.t1345 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1466 XA.XIR[12].XIC[12].icell.PDM XThR.Tn[12].t45 XA.XIR[12].XIC[12].icell.Ien VGND.t402 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1467 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[8].t48 VGND.t842 VGND.t841 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1468 VGND.t1285 XThC.Tn[2].t27 XA.XIR[0].XIC[2].icell.PDM VGND.t1284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1469 XA.XIR[11].XIC[7].icell.PUM XThC.Tn[7].t22 XA.XIR[11].XIC[7].icell.Ien VPWR.t495 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1470 VPWR.t277 XThC.XTBN.Y.t63 XThC.Tn[9].t9 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1471 XA.XIR[15].XIC_15.icell.PUM VPWR.t1586 XA.XIR[15].XIC_15.icell.Ien VPWR.t1587 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1472 XA.XIR[7].XIC[2].icell.SM XA.XIR[7].XIC[2].icell.Ien Iout.t20 VGND.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1473 a_10051_9569# XThC.XTBN.Y.t64 VGND.t442 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1474 VGND.t1780 XThC.Tn[9].t28 XA.XIR[8].XIC[9].icell.PDM VGND.t1779 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1475 XA.XIR[10].XIC[3].icell.SM XA.XIR[10].XIC[3].icell.Ien Iout.t202 VGND.t1935 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1476 VPWR.t196 XThR.XTBN.Y.t63 XThR.Tn[7].t5 VPWR.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1477 VPWR.t257 XThR.Tn[12].t46 XA.XIR[13].XIC[11].icell.PUM VPWR.t256 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1478 XA.XIR[7].XIC[4].icell.PUM XThC.Tn[4].t29 XA.XIR[7].XIC[4].icell.Ien VPWR.t1877 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1479 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR.t1584 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR.t1585 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1480 XA.XIR[13].XIC[4].icell.SM XA.XIR[13].XIC[4].icell.Ien Iout.t232 VGND.t2509 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1481 VPWR.t347 XThR.Tn[9].t40 XA.XIR[10].XIC[7].icell.PUM VPWR.t346 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1482 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[2].t39 XA.XIR[2].XIC[8].icell.Ien VGND.t801 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1483 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[2].t40 XA.XIR[2].XIC[14].icell.Ien VGND.t800 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1484 XThC.Tn[11].t8 XThC.XTB4.Y.t8 VPWR.t1105 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1485 VGND.t316 XThR.XTBN.Y.t64 XThR.Tn[1].t6 VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1486 XThR.Tn[1].t1 XThR.XTBN.Y.t65 a_n1049_7787# VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1487 a_7651_9569# XThC.XTBN.Y.t65 VGND.t443 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1488 XA.XIR[5].XIC[5].icell.PUM XThC.Tn[5].t26 XA.XIR[5].XIC[5].icell.Ien VPWR.t1343 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1489 VGND.t359 Vbias.t141 XA.XIR[11].XIC[5].icell.SM VGND.t358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1490 XA.XIR[10].XIC[6].icell.Ien XThR.Tn[10].t43 VPWR.t1842 VPWR.t1841 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1491 XA.XIR[9].XIC[5].icell.PUM XThC.Tn[5].t27 XA.XIR[9].XIC[5].icell.Ien VPWR.t1344 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1492 XA.XIR[13].XIC[7].icell.Ien XThR.Tn[13].t38 VPWR.t1196 VPWR.t1195 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1493 VGND.t361 Vbias.t142 XA.XIR[5].XIC[9].icell.SM VGND.t360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1494 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2003 VGND.t2449 VGND.t2448 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1495 VPWR.t259 XThR.Tn[12].t47 XA.XIR[13].XIC[2].icell.PUM VPWR.t258 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1496 XA.XIR[14].XIC_dummy_left.icell.SM XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout VGND.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1497 VPWR.t935 XThR.Tn[7].t38 XA.XIR[8].XIC[14].icell.PUM VPWR.t934 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1498 XA.XIR[0].XIC_15.icell.PDM XThR.Tn[0].t48 XA.XIR[0].XIC_15.icell.Ien VGND.t1347 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1499 XA.XIR[10].XIC[9].icell.PDM XThR.Tn[10].t44 XA.XIR[10].XIC[9].icell.Ien VGND.t2565 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1500 XThR.Tn[6].t9 XThR.XTB7.Y VGND.t1744 VGND.t1743 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1501 a_n1049_5611# XThR.XTB6.Y VPWR.t131 VPWR.t130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 XThR.Tn[9].t8 XThR.XTB2.Y VPWR.t1169 VPWR.t1168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1503 VPWR.t1583 VPWR.t1581 XA.XIR[11].XIC_15.icell.PUM VPWR.t1582 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1504 VGND.t363 Vbias.t143 XA.XIR[0].XIC[7].icell.SM VGND.t362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1505 XA.XIR[12].XIC[10].icell.PDM XThR.Tn[12].t48 XA.XIR[12].XIC[10].icell.Ien VGND.t403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1506 Vbias.t8 bias[0].t0 VPWR.t834 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.12325 pd=1.14 as=0.1275 ps=1.15 w=0.85 l=2
X1507 XThC.Tn[4].t4 XThC.XTBN.Y.t66 VGND.t444 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1508 VGND.t481 XThC.Tn[6].t30 XA.XIR[0].XIC[6].icell.PDM VGND.t480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1509 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[5].t44 VGND.t1906 VGND.t1905 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1510 XA.XIR[15].XIC[0].icell.PDM XThR.Tn[14].t43 VGND.t1508 VGND.t1507 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1511 XA.XIR[11].XIC[11].icell.PUM XThC.Tn[11].t28 XA.XIR[11].XIC[11].icell.Ien VPWR.t539 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1512 VPWR.t199 XThR.XTBN.Y.t66 XThR.Tn[13].t9 VPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1513 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[9].t41 VGND.t531 VGND.t530 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1514 XA.XIR[2].XIC[9].icell.Ien XThR.Tn[2].t41 VPWR.t1066 VPWR.t1065 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1515 VGND.t967 VGND.t965 XA.XIR[7].XIC_dummy_right.icell.SM VGND.t966 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1516 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[12].t49 VGND.t405 VGND.t404 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1517 XA.XIR[12].XIC[11].icell.SM XA.XIR[12].XIC[11].icell.Ien Iout.t226 VGND.t2409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1518 VPWR.t736 XThR.Tn[0].t49 XA.XIR[1].XIC[5].icell.PUM VPWR.t735 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1519 VGND.t2451 VPWR.t2004 XA.XIR[13].XIC_dummy_left.icell.PDM VGND.t2450 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1520 VPWR.t145 XThR.Tn[4].t47 XA.XIR[5].XIC[5].icell.PUM VPWR.t144 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1521 VPWR.t349 XThR.Tn[9].t42 XA.XIR[10].XIC[11].icell.PUM VPWR.t348 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1522 XA.XIR[8].XIC[1].icell.PUM XThC.Tn[1].t30 XA.XIR[8].XIC[1].icell.Ien VPWR.t1359 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1523 XA.XIR[4].XIC[4].icell.PUM XThC.Tn[4].t30 XA.XIR[4].XIC[4].icell.Ien VPWR.t1878 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1524 VGND.t1097 XThR.XTB1.Y.t11 XThR.Tn[0].t0 VGND.t1096 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1525 XA.XIR[0].XIC[5].icell.SM XA.XIR[0].XIC[5].icell.Ien Iout.t134 VGND.t1401 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1526 XThR.Tn[5].t9 XThR.XTBN.Y.t67 VGND.t318 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1527 XA.XIR[7].XIC[0].icell.PUM XThC.Tn[0].t26 XA.XIR[7].XIC[0].icell.Ien VPWR.t1216 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1528 XA.XIR[0].XIC[8].icell.PDM VGND.t962 VGND.t964 VGND.t963 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1529 XA.XIR[0].XIC[14].icell.PDM VGND.t959 VGND.t961 VGND.t960 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1530 VGND.t1582 XThR.XTB7.B XThR.XTB6.Y VGND.t1580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1531 XA.XIR[11].XIC[2].icell.PUM XThC.Tn[2].t28 XA.XIR[11].XIC[2].icell.Ien VPWR.t703 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1532 XA.XIR[6].XIC[14].icell.PUM XThC.Tn[14].t27 XA.XIR[6].XIC[14].icell.Ien VPWR.t1297 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1533 VGND.t445 XThC.XTBN.Y.t67 XThC.Tn[0].t8 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1534 VGND.t365 Vbias.t144 XA.XIR[8].XIC[5].icell.SM VGND.t364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1535 XA.XIR[7].XIC[6].icell.Ien XThR.Tn[7].t39 VPWR.t937 VPWR.t936 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1536 XA.XIR[13].XIC[11].icell.Ien XThR.Tn[13].t39 VPWR.t1198 VPWR.t1197 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1537 VGND.t2006 Vbias.t145 XA.XIR[12].XIC[13].icell.SM VGND.t2005 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1538 VGND.t2598 XThC.Tn[4].t31 XA.XIR[8].XIC[4].icell.PDM VGND.t2597 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1539 VGND.t2453 VPWR.t2005 XA.XIR[3].XIC_dummy_right.icell.PDM VGND.t2452 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1540 VGND.t1768 XThC.Tn[12].t29 XA.XIR[12].XIC[12].icell.PDM VGND.t1767 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1541 VGND.t446 XThC.XTBN.Y.t68 XThC.Tn[3].t3 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1542 VGND.t2008 Vbias.t146 XA.XIR[15].XIC[14].icell.SM VGND.t2007 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1543 VGND.t2269 XThC.Tn[5].t28 XA.XIR[11].XIC[5].icell.PDM VGND.t2268 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1544 VGND.t2309 XThC.Tn[13].t29 XA.XIR[15].XIC[13].icell.PDM VGND.t2308 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1545 VPWR.t351 XThR.Tn[9].t43 XA.XIR[10].XIC[2].icell.PUM VPWR.t350 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1546 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[2].t42 XA.XIR[2].XIC[3].icell.Ien VGND.t799 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1547 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR.t2006 XA.XIR[15].XIC_dummy_left.icell.Ien VGND.t2454 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1548 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[7].t40 XA.XIR[7].XIC[9].icell.Ien VGND.t1739 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1549 XThC.Tn[7].t1 XThC.XTBN.Y.t69 VGND.t448 VGND.t447 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1550 VPWR.t278 XThC.XTBN.Y.t70 XThC.Tn[12].t9 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1551 VGND.t2010 Vbias.t147 XA.XIR[11].XIC[0].icell.SM VGND.t2009 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1552 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10].t45 VPWR.t1844 VPWR.t1843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1553 XA.XIR[6].XIC[4].icell.Ien XThR.Tn[6].t44 VPWR.t1379 VPWR.t1378 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1554 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1578 VPWR.t1580 VPWR.t1579 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1555 VGND.t2012 Vbias.t148 XA.XIR[2].XIC_15.icell.SM VGND.t2011 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1556 VGND.t2014 Vbias.t149 XA.XIR[6].XIC[12].icell.SM VGND.t2013 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1557 VGND.t2397 XThC.Tn[8].t27 XA.XIR[2].XIC[8].icell.PDM VGND.t2396 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1558 VGND.t2190 XThC.Tn[14].t28 XA.XIR[2].XIC[14].icell.PDM VGND.t2189 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1559 VPWR.t1167 XThR.XTB2.Y a_n1049_7787# VPWR.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X1560 XA.XIR[13].XIC[2].icell.Ien XThR.Tn[13].t40 VPWR.t1200 VPWR.t1199 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1561 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[9].t44 VGND.t533 VGND.t532 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1562 VGND.t2016 Vbias.t150 XA.XIR[5].XIC[4].icell.SM VGND.t2015 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1563 VGND.t2018 Vbias.t151 XA.XIR[9].XIC[13].icell.SM VGND.t2017 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1564 XA.XIR[9].XIC[8].icell.SM XA.XIR[9].XIC[8].icell.Ien Iout.t151 VGND.t1521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1565 XA.XIR[8].XIC[14].icell.Ien XThR.Tn[8].t49 VPWR.t529 VPWR.t528 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1566 VGND.t450 XThC.XTBN.Y.t71 a_10915_9569# VGND.t449 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1567 VPWR.t586 VGND.t2695 XA.XIR[0].XIC[4].icell.PUM VPWR.t585 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1568 VPWR.t676 XThR.Tn[3].t47 XA.XIR[4].XIC[12].icell.PUM VPWR.t675 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1569 XA.XIR[10].XIC[4].icell.PDM XThR.Tn[10].t46 XA.XIR[10].XIC[4].icell.Ien VGND.t2566 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1570 VPWR.t1064 XThR.Tn[2].t43 XA.XIR[3].XIC[13].icell.PUM VPWR.t1063 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1571 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR.t2007 XA.XIR[5].XIC_dummy_right.icell.Ien VGND.t2455 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1572 XA.XIR[12].XIC[9].icell.SM XA.XIR[12].XIC[9].icell.Ien Iout.t209 VGND.t1987 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1573 XA.XIR[11].XIC_15.icell.Ien XThR.Tn[11].t48 VPWR.t1887 VPWR.t1886 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1574 XThC.Tn[11].t9 XThC.XTB4.Y.t9 a_8963_9569# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1575 XA.XIR[13].XIC[5].icell.PDM XThR.Tn[13].t41 XA.XIR[13].XIC[5].icell.Ien VGND.t2041 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1576 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR.t2008 XA.XIR[9].XIC_dummy_right.icell.Ien VGND.t2456 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1577 VPWR.t1381 XThR.Tn[6].t45 XA.XIR[7].XIC[13].icell.PUM VPWR.t1380 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1578 VGND.t1910 XThC.XTB4.Y.t10 XThC.Tn[3].t9 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1579 VGND.t2020 Vbias.t152 XA.XIR[0].XIC[2].icell.SM VGND.t2019 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1580 XThR.Tn[14].t3 XThR.XTBN.Y.t68 VPWR.t201 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1581 XA.XIR[4].XIC[0].icell.PUM XThC.Tn[0].t27 XA.XIR[4].XIC[0].icell.Ien VPWR.t1217 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1582 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR.t1576 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR.t1577 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1583 a_7875_9569# XThC.XTBN.Y.t72 VGND.t615 VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1584 VPWR.t129 XThR.XTB6.Y XThR.Tn[13].t7 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1585 VGND.t2581 XThC.Tn[10].t30 XA.XIR[12].XIC[10].icell.PDM VGND.t2580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1586 XA.XIR[2].XIC[9].icell.PUM XThC.Tn[9].t29 XA.XIR[2].XIC[9].icell.Ien VPWR.t968 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1587 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[2].t44 XA.XIR[2].XIC[7].icell.Ien VGND.t802 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1588 XA.XIR[0].XIC[0].icell.SM XA.XIR[0].XIC[0].icell.Ien Iout.t227 VGND.t2504 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1589 XA.XIR[0].XIC[3].icell.PDM VGND.t956 VGND.t958 VGND.t957 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1590 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR.t2009 XA.XIR[12].XIC_dummy_left.icell.Ien VGND.t2457 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1591 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[14].t44 XA.XIR[14].XIC[11].icell.Ien VGND.t1509 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1592 XThC.Tn[11].t10 XThC.XTB4.Y.t11 a_8963_9569# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1593 VGND.t2022 Vbias.t153 XA.XIR[8].XIC[0].icell.SM VGND.t2021 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1594 XA.XIR[7].XIC[1].icell.Ien XThR.Tn[7].t41 VPWR.t939 VPWR.t938 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1595 VGND.t2024 Vbias.t154 XA.XIR[3].XIC[12].icell.SM VGND.t2023 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1596 XA.XIR[6].XIC[0].icell.Ien XThR.Tn[6].t46 VPWR.t1383 VPWR.t1382 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1597 VGND.t955 VGND.t953 XA.XIR[7].XIC_dummy_left.icell.SM VGND.t954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1598 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR.t1574 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR.t1575 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1599 XThC.Tn[0].t0 XThC.XTB1.Y.t12 VGND.t1101 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1600 XA.XIR[15].XIC[5].icell.SM XA.XIR[15].XIC[5].icell.Ien Iout.t93 VGND.t1127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1601 VGND.t616 XThC.XTBN.Y.t73 a_10051_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1602 VGND.t2092 XThC.Tn[0].t28 XA.XIR[11].XIC[0].icell.PDM VGND.t2091 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1603 VPWR.t678 XThR.Tn[3].t48 XA.XIR[4].XIC[10].icell.PUM VPWR.t677 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1604 VGND.t331 XThC.Tn[12].t30 XA.XIR[6].XIC[12].icell.PDM VGND.t330 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1605 XThR.XTB1.Y.t2 XThR.XTB5.A VPWR.t925 VPWR.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 VPWR.t584 VGND.t2696 XA.XIR[0].XIC[0].icell.PUM VPWR.t583 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1607 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[7].t42 XA.XIR[7].XIC[4].icell.Ien VGND.t1740 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1608 XThR.Tn[13].t0 XThR.XTB6.Y a_n997_1579# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1609 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[14].t45 XA.XIR[14].XIC[2].icell.Ien VGND.t1510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1610 XA.XIR[10].XIC[7].icell.PUM XThC.Tn[7].t23 XA.XIR[10].XIC[7].icell.Ien VPWR.t496 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1611 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR.t2010 VGND.t2459 VGND.t2458 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1612 VGND.t1435 XThC.Tn[3].t28 XA.XIR[2].XIC[3].icell.PDM VGND.t1434 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1613 XA.XIR[13].XIC[8].icell.PUM XThC.Tn[8].t28 XA.XIR[13].XIC[8].icell.Ien VPWR.t869 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1614 VGND.t617 XThC.XTBN.Y.t74 a_7651_9569# VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1615 XA.XIR[4].XIC[12].icell.Ien XThR.Tn[4].t48 VPWR.t147 VPWR.t146 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1616 XA.XIR[9].XIC[3].icell.SM XA.XIR[9].XIC[3].icell.Ien Iout.t60 VGND.t646 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1617 XThC.XTBN.Y.t0 XThC.XTBN.A VGND.t674 VGND.t673 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1618 XA.XIR[3].XIC[13].icell.Ien XThR.Tn[3].t49 VPWR.t680 VPWR.t679 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1619 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1571 VPWR.t1573 VPWR.t1572 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1620 XA.XIR[1].XIC[14].icell.PDM XThR.Tn[1].t44 XA.XIR[1].XIC[14].icell.Ien VGND.t831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1621 XA.XIR[12].XIC[4].icell.SM XA.XIR[12].XIC[4].icell.Ien Iout.t76 VGND.t870 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1622 XA.XIR[1].XIC[8].icell.PDM XThR.Tn[1].t45 XA.XIR[1].XIC[8].icell.Ien VGND.t832 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1623 XA.XIR[7].XIC_dummy_right.icell.SM XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout VGND.t1325 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1624 a_n1335_7243# XThR.XTB7.A XThR.XTB3.Y.t1 VGND.t2645 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 XA.XIR[13].XIC[0].icell.PDM XThR.Tn[13].t42 XA.XIR[13].XIC[0].icell.Ien VGND.t1810 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1626 XA.XIR[8].XIC[12].icell.PDM XThR.Tn[8].t50 XA.XIR[8].XIC[12].icell.Ien VGND.t1130 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1627 XA.XIR[0].XIC[7].icell.PDM VGND.t950 VGND.t952 VGND.t951 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1628 a_n1049_5317# XThR.XTBN.Y.t69 XThR.Tn[6].t2 VPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1629 XA.XIR[11].XIC[13].icell.PDM XThR.Tn[11].t49 XA.XIR[11].XIC[13].icell.Ien VGND.t2609 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1630 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2011 VGND.t2461 VGND.t2460 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1631 a_4067_9615# XThC.XTB3.Y.t10 VPWR.t32 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1632 VPWR.t429 XThC.XTBN.Y.t75 XThC.Tn[7].t4 VPWR.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1633 VPWR.t1062 XThR.Tn[2].t45 XA.XIR[3].XIC[6].icell.PUM VPWR.t1061 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1634 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[11].t50 VGND.t2611 VGND.t2610 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1635 XA.XIR[15].XIC[8].icell.Ien VPWR.t1568 VPWR.t1570 VPWR.t1569 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1636 VPWR.t1385 XThR.Tn[6].t47 XA.XIR[7].XIC[6].icell.PUM VPWR.t1384 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1637 VGND.t320 XThR.XTBN.Y.t70 a_n997_1803# VGND.t319 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1638 VPWR.t1100 XThR.Tn[5].t45 XA.XIR[6].XIC[7].icell.PUM VPWR.t1099 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1639 XThR.Tn[3].t5 XThR.XTBN.Y.t71 VGND.t322 VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1640 VGND.t2583 XThC.Tn[10].t31 XA.XIR[6].XIC[10].icell.PDM VGND.t2582 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1641 VPWR.t652 XThR.Tn[8].t51 XA.XIR[9].XIC[8].icell.PUM VPWR.t651 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1642 VPWR.t1106 XThC.XTB4.Y.t12 XThC.Tn[11].t11 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[14].t46 XA.XIR[14].XIC[6].icell.Ien VGND.t1511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1644 XA.XIR[10].XIC[11].icell.PUM XThC.Tn[11].t29 XA.XIR[10].XIC[11].icell.Ien VPWR.t540 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1645 VGND.t2026 Vbias.t155 XA.XIR[2].XIC[8].icell.SM VGND.t2025 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1646 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[12].t50 VGND.t2197 VGND.t2196 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1647 XA.XIR[1].XIC[9].icell.Ien XThR.Tn[1].t46 VPWR.t509 VPWR.t508 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1648 VGND.t819 XThC.Tn[7].t24 XA.XIR[2].XIC[7].icell.PDM VGND.t818 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1649 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[11].t51 VGND.t2613 VGND.t2612 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1650 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[7].t43 VGND.t1754 VGND.t1753 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1651 XA.XIR[4].XIC[10].icell.Ien XThR.Tn[4].t49 VPWR.t149 VPWR.t148 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1652 XA.XIR[15].XIC[0].icell.SM XA.XIR[15].XIC[0].icell.Ien Iout.t139 VGND.t1431 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1653 VGND.t2463 VPWR.t2012 XA.XIR[12].XIC_dummy_left.icell.PDM VGND.t2462 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1654 XThC.Tn[0].t7 XThC.XTBN.Y.t76 VGND.t618 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 XA.XIR[10].XIC[12].icell.SM XA.XIR[10].XIC[12].icell.Ien Iout.t205 VGND.t1954 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1656 VPWR.t682 XThR.Tn[3].t50 XA.XIR[4].XIC[5].icell.PUM VPWR.t681 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1657 XA.XIR[13].XIC[13].icell.SM XA.XIR[13].XIC[13].icell.Ien Iout.t80 VGND.t879 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1658 XThC.Tn[3].t2 XThC.XTBN.Y.t77 VGND.t619 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1659 VGND.t1575 XThC.Tn[8].t29 XA.XIR[14].XIC[8].icell.PDM VGND.t1574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1660 VGND.t2192 XThC.Tn[14].t29 XA.XIR[14].XIC[14].icell.PDM VGND.t2191 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1661 XA.XIR[10].XIC[2].icell.PUM XThC.Tn[2].t29 XA.XIR[10].XIC[2].icell.Ien VPWR.t704 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1662 XA.XIR[8].XIC[10].icell.PDM XThR.Tn[8].t52 XA.XIR[8].XIC[10].icell.Ien VGND.t1131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1663 XA.XIR[5].XIC[14].icell.PUM XThC.Tn[14].t30 XA.XIR[5].XIC[14].icell.Ien VPWR.t1298 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1664 XA.XIR[13].XIC[3].icell.PUM XThC.Tn[3].t29 XA.XIR[13].XIC[3].icell.Ien VPWR.t772 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1665 XA.XIR[9].XIC[14].icell.PUM XThC.Tn[14].t31 XA.XIR[9].XIC[14].icell.Ien VPWR.t1299 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1666 XA.XIR[8].XIC_15.icell.PUM VPWR.t1566 XA.XIR[8].XIC_15.icell.Ien VPWR.t1567 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1667 a_n1049_8581# XThR.XTB1.Y.t12 VPWR.t617 VPWR.t616 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1668 VGND.t2312 XThC.Tn[1].t31 XA.XIR[15].XIC[1].icell.PDM VGND.t2311 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1669 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[8].t53 VGND.t1133 VGND.t1132 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1670 VPWR.t1565 VPWR.t1563 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR.t1564 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1671 VGND.t2028 Vbias.t156 XA.XIR[10].XIC[6].icell.SM VGND.t2027 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1672 VGND.t2271 XThC.Tn[5].t29 XA.XIR[10].XIC[5].icell.PDM VGND.t2270 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1673 XA.XIR[1].XIC[3].icell.PDM XThR.Tn[1].t47 XA.XIR[1].XIC[3].icell.Ien VGND.t833 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1674 XA.XIR[12].XIC[8].icell.Ien XThR.Tn[12].t51 VPWR.t1301 VPWR.t1300 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1675 VPWR.t1102 XThR.Tn[5].t46 XA.XIR[6].XIC[11].icell.PUM VPWR.t1101 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1676 XA.XIR[0].XIC[4].icell.PUM XThC.Tn[4].t32 XA.XIR[0].XIC[4].icell.Ien VPWR.t1879 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1677 VGND.t1169 Vbias.t157 XA.XIR[1].XIC_15.icell.SM VGND.t1168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1678 XA.XIR[7].XIC[13].icell.PUM XThC.Tn[13].t30 XA.XIR[7].XIC[13].icell.Ien VPWR.t1358 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1679 XThC.XTB1.Y.t1 XThC.XTB5.A a_3299_10575# VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1680 XA.XIR[3].XIC[6].icell.Ien XThR.Tn[3].t51 VPWR.t684 VPWR.t683 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1681 VPWR.t1060 XThR.Tn[2].t46 XA.XIR[3].XIC[1].icell.PUM VPWR.t1059 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1682 VGND.t294 XThR.XTB3.Y.t10 XThR.Tn[2].t0 VGND.t191 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 XA.XIR[15].XIC[3].icell.Ien VPWR.t1560 VPWR.t1562 VPWR.t1561 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1684 XA.XIR[12].XIC[6].icell.PDM XThR.Tn[11].t52 VGND.t2615 VGND.t2614 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1685 VGND.t1171 Vbias.t158 XA.XIR[11].XIC[14].icell.SM VGND.t1170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1686 XA.XIR[10].XIC_15.icell.Ien XThR.Tn[10].t47 VPWR.t1846 VPWR.t1845 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1687 XA.XIR[14].XIC[9].icell.PUM XThC.Tn[9].t30 XA.XIR[14].XIC[9].icell.Ien VPWR.t969 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1688 VPWR.t1387 XThR.Tn[6].t48 XA.XIR[7].XIC[1].icell.PUM VPWR.t1386 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1689 VPWR.t1104 XThR.Tn[5].t47 XA.XIR[6].XIC[2].icell.PUM VPWR.t1103 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1690 XA.XIR[7].XIC_dummy_left.icell.SM XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout VGND.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1691 VPWR.t286 XThR.Tn[0].t50 XA.XIR[1].XIC[14].icell.PUM VPWR.t285 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1692 XA.XIR[3].XIC[9].icell.PDM XThR.Tn[3].t52 XA.XIR[3].XIC[9].icell.Ien VGND.t2510 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1693 VPWR.t151 XThR.Tn[4].t50 XA.XIR[5].XIC[14].icell.PUM VPWR.t150 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1694 VPWR.t654 XThR.Tn[8].t54 XA.XIR[9].XIC[3].icell.PUM VPWR.t653 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1695 VGND.t621 XThC.XTBN.Y.t78 XThC.Tn[6].t10 VGND.t620 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1696 VGND.t1173 Vbias.t159 XA.XIR[2].XIC[3].icell.SM VGND.t1172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1697 XA.XIR[6].XIC[7].icell.SM XA.XIR[6].XIC[7].icell.Ien Iout.t55 VGND.t583 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1698 XThC.Tn[10].t3 XThC.XTB3.Y.t11 VPWR.t33 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1699 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[7].t44 VGND.t1756 VGND.t1755 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1700 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[2].t47 VGND.t145 VGND.t144 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1701 XA.XIR[4].XIC[5].icell.Ien XThR.Tn[4].t51 VPWR.t153 VPWR.t152 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1702 VGND.t949 VGND.t947 XA.XIR[0].XIC_dummy_right.icell.SM VGND.t948 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1703 VGND.t1175 Vbias.t160 XA.XIR[14].XIC[7].icell.SM VGND.t1174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1704 VGND.t1177 Vbias.t161 XA.XIR[10].XIC[10].icell.SM VGND.t1176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1705 XThC.Tn[14].t6 XThC.XTB7.Y VPWR.t113 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1706 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[5].t48 VGND.t1908 VGND.t1907 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1707 XA.XIR[1].XIC[7].icell.PDM XThR.Tn[1].t48 XA.XIR[1].XIC[7].icell.Ien VGND.t834 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1708 VGND.t2465 VPWR.t2013 XA.XIR[6].XIC_dummy_left.icell.PDM VGND.t2464 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1709 VGND.t1102 XThC.XTB1.Y.t13 XThC.Tn[0].t1 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1710 VGND.t1437 XThC.Tn[3].t30 XA.XIR[14].XIC[3].icell.PDM VGND.t1436 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1711 XA.XIR[0].XIC[0].icell.PUM XThC.Tn[0].t29 XA.XIR[0].XIC[0].icell.Ien VPWR.t1218 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1712 XA.XIR[1].XIC[12].icell.PUM XThC.Tn[12].t31 XA.XIR[1].XIC[12].icell.Ien VPWR.t212 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1713 XA.XIR[4].XIC[13].icell.PUM XThC.Tn[13].t31 XA.XIR[4].XIC[13].icell.Ien VPWR.t1132 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1714 VGND.t1179 Vbias.t162 XA.XIR[10].XIC[1].icell.SM VGND.t1178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1715 XThR.Tn[8].t5 XThR.XTBN.Y.t72 VPWR.t204 VPWR.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1716 XA.XIR[0].XIC[14].icell.SM XA.XIR[0].XIC[14].icell.Ien Iout.t132 VGND.t1399 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1717 VGND.t1181 Vbias.t163 XA.XIR[5].XIC[13].icell.SM VGND.t1180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1718 XA.XIR[14].XIC[5].icell.SM XA.XIR[14].XIC[5].icell.Ien Iout.t198 VGND.t1875 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1719 XA.XIR[14].XIC[8].icell.PDM XThR.Tn[13].t43 VGND.t1812 VGND.t1811 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1720 XA.XIR[14].XIC[14].icell.PDM XThR.Tn[13].t44 VGND.t1814 VGND.t1813 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1721 VGND.t2094 XThC.Tn[0].t30 XA.XIR[10].XIC[0].icell.PDM VGND.t2093 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1722 VGND.t333 XThC.Tn[12].t32 XA.XIR[5].XIC[12].icell.PDM VGND.t332 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1723 XA.XIR[12].XIC[3].icell.Ien XThR.Tn[12].t52 VPWR.t1303 VPWR.t1302 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1724 VGND.t335 XThC.Tn[12].t33 XA.XIR[9].XIC[12].icell.PDM VGND.t334 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1725 VGND.t1183 Vbias.t164 XA.XIR[8].XIC[14].icell.SM VGND.t1182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1726 XA.XIR[7].XIC_15.icell.Ien XThR.Tn[7].t45 VPWR.t949 VPWR.t948 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1727 VGND.t1940 XThC.Tn[13].t32 XA.XIR[8].XIC[13].icell.PDM VGND.t1939 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1728 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR.t2014 XA.XIR[8].XIC_dummy_left.icell.Ien VGND.t2466 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1729 a_n1049_5611# XThR.XTBN.Y.t73 XThR.Tn[5].t5 VPWR.t202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1730 XA.XIR[3].XIC[1].icell.Ien XThR.Tn[3].t53 VPWR.t1397 VPWR.t1396 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1731 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[4].t52 VGND.t283 VGND.t282 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1732 XA.XIR[12].XIC[8].icell.PUM XThC.Tn[8].t30 XA.XIR[12].XIC[8].icell.Ien VPWR.t870 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1733 VGND.t1185 Vbias.t165 XA.XIR[4].XIC[11].icell.SM VGND.t1184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1734 XA.XIR[3].XIC[7].icell.SM XA.XIR[3].XIC[7].icell.Ien Iout.t6 VGND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1735 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[2].t48 VGND.t143 VGND.t142 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1736 XThR.XTBN.A data[7].t1 VGND.t372 VGND.t371 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1737 XA.XIR[6].XIC[13].icell.Ien XThR.Tn[6].t49 VPWR.t1389 VPWR.t1388 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1738 XA.XIR[3].XIC[4].icell.PDM XThR.Tn[3].t54 XA.XIR[3].XIC[4].icell.Ien VGND.t2511 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1739 XThC.Tn[14].t5 XThC.XTB7.Y VPWR.t112 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1740 VPWR.t984 XThR.Tn[13].t45 XA.XIR[14].XIC[4].icell.PUM VPWR.t983 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1741 XA.XIR[11].XIC[1].icell.PDM XThR.Tn[11].t53 XA.XIR[11].XIC[1].icell.Ien VGND.t2593 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1742 XA.XIR[7].XIC[6].icell.PUM XThC.Tn[6].t31 XA.XIR[7].XIC[6].icell.Ien VPWR.t301 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1743 VPWR.t582 VGND.t2697 XA.XIR[0].XIC[13].icell.PUM VPWR.t581 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1744 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2015 XA.XIR[2].XIC_dummy_right.icell.Ien VGND.t2467 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1745 VGND.t821 XThC.Tn[7].t25 XA.XIR[14].XIC[7].icell.PDM VGND.t820 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1746 XA.XIR[10].XIC[13].icell.PDM XThR.Tn[10].t48 XA.XIR[10].XIC[13].icell.Ien VGND.t2567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1747 XThC.XTB2.Y XThC.XTB7.B VPWR.t728 VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1748 XA.XIR[1].XIC[10].icell.PUM XThC.Tn[10].t32 XA.XIR[1].XIC[10].icell.Ien VPWR.t391 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1749 XA.XIR[6].XIC[2].icell.SM XA.XIR[6].XIC[2].icell.Ien Iout.t31 VGND.t203 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1750 XA.XIR[0].XIC[12].icell.Ien XThR.Tn[0].t51 VPWR.t288 VPWR.t287 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1751 XThR.Tn[5].t8 XThR.XTBN.Y.t74 VGND.t324 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1752 VGND.t1782 XThC.Tn[9].t31 XA.XIR[7].XIC[9].icell.PDM VGND.t1781 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1753 XA.XIR[15].XIC[11].icell.PDM XThR.Tn[14].t47 VGND.t1513 VGND.t1512 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1754 VGND.t1187 Vbias.t166 XA.XIR[14].XIC[2].icell.SM VGND.t1186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1755 VGND.t571 XThC.Tn[10].t33 XA.XIR[5].XIC[10].icell.PDM VGND.t570 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1756 XThR.Tn[10].t3 XThR.XTBN.Y.t75 VPWR.t206 VPWR.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1757 VPWR.t951 XThR.Tn[7].t46 XA.XIR[8].XIC[8].icell.PUM VPWR.t950 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1758 VGND.t573 XThC.Tn[10].t34 XA.XIR[9].XIC[10].icell.PDM VGND.t572 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1759 a_5949_9615# XThC.XTB6.Y VPWR.t766 VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1760 VGND.t1189 Vbias.t167 XA.XIR[1].XIC[8].icell.SM VGND.t1188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1761 VGND.t1191 Vbias.t168 XA.XIR[4].XIC[9].icell.SM VGND.t1190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1762 XA.XIR[14].XIC[0].icell.SM XA.XIR[14].XIC[0].icell.Ien Iout.t50 VGND.t475 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1763 XA.XIR[15].XIC[2].icell.PDM XThR.Tn[14].t48 VGND.t1515 VGND.t1514 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1764 VPWR.t34 XThC.XTB3.Y.t12 XThC.Tn[10].t4 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1765 XA.XIR[14].XIC[3].icell.PDM XThR.Tn[13].t46 VGND.t1816 VGND.t1815 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1766 VGND.t946 VGND.t944 XA.XIR[0].XIC_dummy_left.icell.SM VGND.t945 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1767 XA.XIR[5].XIC_15.icell.SM XA.XIR[5].XIC_15.icell.Ien Iout.t144 VGND.t1454 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1768 XA.XIR[9].XIC[12].icell.SM XA.XIR[9].XIC[12].icell.Ien Iout.t150 VGND.t1520 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1769 XThC.Tn[13].t8 XThC.XTBN.Y.t79 VPWR.t430 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1770 XA.XIR[13].XIC_15.icell.PDM VPWR.t2016 VGND.t2469 VGND.t2468 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1771 a_n997_3755# XThR.XTBN.Y.t76 VGND.t492 VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1772 XA.XIR[12].XIC[13].icell.SM XA.XIR[12].XIC[13].icell.Ien Iout.t14 VGND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1773 VPWR.t307 XThR.XTBN.Y.t77 XThR.Tn[14].t2 VPWR.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 XA.XIR[15].XIC[14].icell.SM XA.XIR[15].XIC[14].icell.Ien Iout.t97 VGND.t1137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1775 XA.XIR[4].XIC[6].icell.PUM XThC.Tn[6].t32 XA.XIR[4].XIC[6].icell.Ien VPWR.t302 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1776 XA.XIR[9].XIC[1].icell.PDM XThR.Tn[8].t55 VGND.t1135 VGND.t1134 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1777 XA.XIR[3].XIC[7].icell.PUM XThC.Tn[7].t26 XA.XIR[3].XIC[7].icell.Ien VPWR.t497 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1778 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[4].t53 VGND.t2148 VGND.t2147 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1779 XA.XIR[12].XIC[3].icell.PUM XThC.Tn[3].t31 XA.XIR[12].XIC[3].icell.Ien VPWR.t773 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1780 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2017 VGND.t2471 VGND.t2470 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1781 VPWR.t986 XThR.Tn[13].t47 XA.XIR[14].XIC[0].icell.PUM VPWR.t985 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1782 XA.XIR[7].XIC[13].icell.PDM XThR.Tn[7].t47 XA.XIR[7].XIC[13].icell.Ien VGND.t1757 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1783 XA.XIR[0].XIC[10].icell.Ien XThR.Tn[0].t52 VPWR.t290 VPWR.t289 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1784 XA.XIR[3].XIC[2].icell.SM XA.XIR[3].XIC[2].icell.Ien Iout.t78 VGND.t872 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1785 XA.XIR[6].XIC[8].icell.PUM XThC.Tn[8].t31 XA.XIR[6].XIC[8].icell.Ien VPWR.t871 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1786 XA.XIR[11].XIC[11].icell.SM XA.XIR[11].XIC[11].icell.Ien Iout.t56 VGND.t640 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1787 XThR.Tn[7].t0 XThR.XTBN.Y.t78 VGND.t494 VGND.t493 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1788 XA.XIR[2].XIC_15.icell.SM XA.XIR[2].XIC_15.icell.Ien Iout.t156 VGND.t1531 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1789 VPWR.t1559 VPWR.t1557 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1558 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1790 VGND.t1784 XThC.Tn[9].t32 XA.XIR[4].XIC[9].icell.PDM VGND.t1783 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1791 XA.XIR[14].XIC[4].icell.Ien XThR.Tn[14].t49 VPWR.t1224 VPWR.t1223 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1792 XA.XIR[7].XIC[1].icell.PUM XThC.Tn[1].t32 XA.XIR[7].XIC[1].icell.Ien VPWR.t1360 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1793 VGND.t2473 VPWR.t2018 XA.XIR[15].XIC_15.icell.PDM VGND.t2472 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1794 XThC.XTB4.Y.t0 XThC.XTB7.B VGND.t1332 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1795 VPWR.t127 XThR.XTB6.Y XThR.Tn[13].t6 VPWR.t126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VPWR.t1111 XThR.XTB3.Y.t11 a_n1049_7493# VPWR.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1797 XA.XIR[1].XIC[5].icell.PUM XThC.Tn[5].t30 XA.XIR[1].XIC[5].icell.Ien VPWR.t1345 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1798 VPWR.t1870 XThR.Tn[11].t54 XA.XIR[12].XIC[12].icell.PUM VPWR.t1869 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1799 VGND.t2367 Vbias.t169 XA.XIR[7].XIC[5].icell.SM VGND.t2366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1800 XA.XIR[6].XIC[6].icell.Ien XThR.Tn[6].t50 VPWR.t1391 VPWR.t1390 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1801 XA.XIR[5].XIC[7].icell.Ien XThR.Tn[5].t49 VPWR.t844 VPWR.t843 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1802 VPWR.t1109 data[4].t3 XThR.XTB7.A VPWR.t1108 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1803 VGND.t2600 XThC.Tn[4].t33 XA.XIR[7].XIC[4].icell.PDM VGND.t2599 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1804 VGND.t2369 Vbias.t170 XA.XIR[6].XIC[6].icell.SM VGND.t2368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1805 VGND.t2475 VPWR.t2019 XA.XIR[2].XIC_dummy_right.icell.PDM VGND.t2474 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1806 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2020 VGND.t2477 VGND.t2476 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1807 XA.XIR[15].XIC[6].icell.PDM XThR.Tn[14].t50 VGND.t2110 VGND.t2109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1808 XThC.Tn[6].t9 XThC.XTBN.Y.t80 VGND.t623 VGND.t622 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1809 XA.XIR[14].XIC[7].icell.PDM XThR.Tn[13].t48 VGND.t1032 VGND.t1031 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1810 XA.XIR[9].XIC[7].icell.Ien XThR.Tn[9].t45 VPWR.t353 VPWR.t352 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1811 XA.XIR[8].XIC[8].icell.Ien XThR.Tn[8].t56 VPWR.t656 VPWR.t655 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1812 VPWR.t580 VGND.t2698 XA.XIR[0].XIC[6].icell.PUM VPWR.t579 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1813 VPWR.t1399 XThR.Tn[3].t55 XA.XIR[4].XIC[14].icell.PUM VPWR.t1398 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1814 XThR.Tn[5].t1 XThR.XTB6.Y VGND.t257 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1815 VPWR.t953 XThR.Tn[7].t48 XA.XIR[8].XIC[3].icell.PUM VPWR.t952 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1816 VPWR.t163 XThC.XTB5.Y a_5155_9615# VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 VPWR.t1556 VPWR.t1554 XA.XIR[3].XIC_15.icell.PUM VPWR.t1555 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1818 XA.XIR[6].XIC[9].icell.PDM XThR.Tn[6].t51 XA.XIR[6].XIC[9].icell.Ien VGND.t2403 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1819 VPWR.t1553 VPWR.t1551 XA.XIR[7].XIC_15.icell.PUM VPWR.t1552 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1820 VGND.t2371 Vbias.t171 XA.XIR[1].XIC[3].icell.SM VGND.t2370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1821 XA.XIR[3].XIC[11].icell.PUM XThC.Tn[11].t30 XA.XIR[3].XIC[11].icell.Ien VPWR.t813 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1822 XThR.Tn[4].t10 XThR.XTB5.Y VGND.t2652 VGND.t260 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1823 a_4861_9615# XThC.XTB4.Y.t13 VPWR.t1107 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X1824 a_5949_9615# XThC.XTBN.Y.t81 XThC.Tn[5].t9 VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1825 VGND.t2373 Vbias.t172 XA.XIR[4].XIC[4].icell.SM VGND.t2372 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1826 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[5].t50 VGND.t1539 VGND.t1538 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1827 VGND.t2479 VPWR.t2021 XA.XIR[5].XIC_dummy_left.icell.PDM VGND.t2478 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1828 XA.XIR[11].XIC[9].icell.SM XA.XIR[11].XIC[9].icell.Ien Iout.t49 VGND.t422 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1829 VGND.t624 XThC.XTBN.Y.t82 XThC.Tn[2].t9 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1830 VGND.t2481 VPWR.t2022 XA.XIR[9].XIC_dummy_left.icell.PDM VGND.t2480 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1831 XA.XIR[8].XIC[11].icell.SM XA.XIR[8].XIC[11].icell.Ien Iout.t216 VGND.t2153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1832 VPWR.t625 XThC.XTB1.Y.t14 XThC.Tn[8].t5 VPWR.t624 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 VGND.t1492 XThC.Tn[11].t31 XA.XIR[11].XIC[11].icell.PDM VGND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1834 a_5155_10571# XThC.XTB7.B XThC.XTB5.Y VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1835 a_10915_9569# XThC.XTBN.Y.t83 VGND.t503 VGND.t502 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1836 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14].t51 VPWR.t1226 VPWR.t1225 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1837 XA.XIR[4].XIC[1].icell.PUM XThC.Tn[1].t33 XA.XIR[4].XIC[1].icell.Ien VPWR.t1361 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1838 XA.XIR[3].XIC[2].icell.PUM XThC.Tn[2].t30 XA.XIR[3].XIC[2].icell.Ien VPWR.t705 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1839 VPWR.t1872 XThR.Tn[11].t55 XA.XIR[12].XIC[10].icell.PUM VPWR.t1871 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1840 XA.XIR[0].XIC[5].icell.Ien XThR.Tn[0].t53 VPWR.t292 VPWR.t291 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1841 XA.XIR[6].XIC[3].icell.PUM XThC.Tn[3].t32 XA.XIR[6].XIC[3].icell.Ien VPWR.t774 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1842 VGND.t2375 Vbias.t173 XA.XIR[6].XIC[10].icell.SM VGND.t2374 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1843 XA.XIR[5].XIC[11].icell.Ien XThR.Tn[5].t51 VPWR.t846 VPWR.t845 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1844 XThC.Tn[3].t8 XThC.XTB4.Y.t14 VGND.t1911 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1845 VGND.t2377 Vbias.t174 XA.XIR[3].XIC[6].icell.SM VGND.t2376 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1846 VGND.t2602 XThC.Tn[4].t34 XA.XIR[4].XIC[4].icell.PDM VGND.t2601 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1847 VGND.t2314 XThC.Tn[1].t34 XA.XIR[8].XIC[1].icell.PDM VGND.t2313 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1848 VGND.t2273 XThC.Tn[5].t31 XA.XIR[3].XIC[5].icell.PDM VGND.t2272 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1849 XA.XIR[9].XIC[11].icell.Ien XThR.Tn[9].t46 VPWR.t382 VPWR.t381 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1850 VGND.t1287 XThC.Tn[2].t31 XA.XIR[11].XIC[2].icell.PDM VGND.t1286 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1851 XA.XIR[4].XIC[9].icell.PDM XThR.Tn[3].t56 VGND.t2513 VGND.t2512 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1852 XA.XIR[13].XIC[11].icell.PDM XThR.Tn[13].t49 XA.XIR[13].XIC[11].icell.Ien VGND.t1033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1853 XThR.Tn[3].t4 XThR.XTBN.Y.t79 VGND.t496 VGND.t495 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1854 XA.XIR[0].XIC[13].icell.PUM XThC.Tn[13].t33 XA.XIR[0].XIC[13].icell.Ien VPWR.t1133 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1855 XA.XIR[6].XIC[1].icell.Ien XThR.Tn[6].t52 VPWR.t1393 VPWR.t1392 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1856 VGND.t2379 Vbias.t175 XA.XIR[7].XIC[0].icell.SM VGND.t2378 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1857 VGND.t2381 Vbias.t176 XA.XIR[2].XIC[12].icell.SM VGND.t2380 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1858 XA.XIR[5].XIC[2].icell.Ien XThR.Tn[5].t52 VPWR.t848 VPWR.t847 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1859 VGND.t2383 Vbias.t177 XA.XIR[6].XIC[1].icell.SM VGND.t2382 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1860 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR.t1549 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR.t1550 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1861 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t1 VGND.t219 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1862 XA.XIR[9].XIC[2].icell.Ien XThR.Tn[9].t47 VPWR.t384 VPWR.t383 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1863 a_4387_10575# XThC.XTB7.B VGND.t1331 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1864 XA.XIR[4].XIC[14].icell.Ien XThR.Tn[4].t54 VPWR.t1260 VPWR.t1259 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1865 XA.XIR[5].XIC[8].icell.SM XA.XIR[5].XIC[8].icell.Ien Iout.t90 VGND.t1119 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1866 XA.XIR[8].XIC[3].icell.Ien XThR.Tn[8].t57 VPWR.t561 VPWR.t560 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1867 VPWR.t578 VGND.t2699 XA.XIR[0].XIC[1].icell.PUM VPWR.t577 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1868 XA.XIR[3].XIC_15.icell.Ien XThR.Tn[3].t57 VPWR.t1401 VPWR.t1400 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1869 XA.XIR[10].XIC[1].icell.PDM XThR.Tn[10].t49 XA.XIR[10].XIC[1].icell.Ien VGND.t1440 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1870 XA.XIR[8].XIC[9].icell.SM XA.XIR[8].XIC[9].icell.Ien Iout.t68 VGND.t807 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1871 XA.XIR[6].XIC[4].icell.PDM XThR.Tn[6].t53 XA.XIR[6].XIC[4].icell.Ien VGND.t2404 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1872 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR.t2023 XA.XIR[1].XIC_dummy_right.icell.Ien VGND.t2482 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1873 XA.XIR[5].XIC[5].icell.PDM XThR.Tn[5].t53 XA.XIR[5].XIC[5].icell.Ien VGND.t1540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1874 XA.XIR[13].XIC[2].icell.PDM XThR.Tn[13].t50 XA.XIR[13].XIC[2].icell.Ien VGND.t1034 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1875 XA.XIR[9].XIC[5].icell.PDM XThR.Tn[9].t48 XA.XIR[9].XIC[5].icell.Ien VGND.t557 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1876 a_10051_9569# XThC.XTBN.Y.t84 VGND.t504 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1877 XA.XIR[11].XIC_15.icell.PDM XThR.Tn[11].t56 XA.XIR[11].XIC_15.icell.Ien VGND.t2594 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1878 XThC.XTB1.Y.t0 XThC.XTB7.B VPWR.t727 VPWR.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1879 a_n1049_6699# XThR.XTBN.Y.t80 XThR.Tn[3].t9 VPWR.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1880 XA.XIR[2].XIC[8].icell.SM XA.XIR[2].XIC[8].icell.Ien Iout.t82 VGND.t881 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1881 XA.XIR[11].XIC[4].icell.SM XA.XIR[11].XIC[4].icell.Ien Iout.t158 VGND.t1533 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1882 VGND.t2385 Vbias.t178 XA.XIR[3].XIC[10].icell.SM VGND.t2384 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1883 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1546 VPWR.t1548 VPWR.t1547 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1884 XA.XIR[6].XIC_dummy_right.icell.SM XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1885 a_n1049_8581# XThR.XTBN.Y.t81 XThR.Tn[0].t2 VPWR.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1886 a_7651_9569# XThC.XTBN.Y.t85 VGND.t505 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1887 VGND.t943 VGND.t941 XA.XIR[14].XIC_dummy_right.icell.SM VGND.t942 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1888 VGND.t483 XThC.Tn[6].t33 XA.XIR[11].XIC[6].icell.PDM VGND.t482 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1889 VPWR.t1406 XThC.XTB7.A a_6243_10571# VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1890 VPWR.t1545 VPWR.t1543 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1544 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1891 XA.XIR[1].XIC[9].icell.PDM XThR.Tn[0].t54 VGND.t465 VGND.t464 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1892 VPWR.t1874 XThR.Tn[11].t57 XA.XIR[12].XIC[5].icell.PUM VPWR.t1873 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1893 XThC.Tn[10].t5 XThC.XTB3.Y.t13 a_8739_9569# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1894 VGND.t2387 Vbias.t179 XA.XIR[3].XIC[1].icell.SM VGND.t2386 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1895 XA.XIR[7].XIC[5].icell.SM XA.XIR[7].XIC[5].icell.Ien Iout.t247 VGND.t2617 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1896 VGND.t2096 XThC.Tn[0].t31 XA.XIR[3].XIC[0].icell.PDM VGND.t2095 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1897 VGND.t498 XThR.XTBN.Y.t82 XThR.Tn[2].t4 VGND.t497 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1898 XA.XIR[11].XIC[14].icell.PDM XThR.Tn[10].t50 VGND.t1442 VGND.t1441 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1899 XA.XIR[11].XIC[8].icell.PDM XThR.Tn[10].t51 VGND.t1444 VGND.t1443 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1900 XA.XIR[10].XIC[6].icell.SM XA.XIR[10].XIC[6].icell.Ien Iout.t81 VGND.t880 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1901 XThR.XTB5.A data[5].t3 VGND.t281 VGND.t280 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 XA.XIR[14].XIC[14].icell.SM XA.XIR[14].XIC[14].icell.Ien Iout.t170 VGND.t1619 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1903 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR.t1541 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR.t1542 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1904 XA.XIR[4].XIC[4].icell.PDM XThR.Tn[3].t58 VGND.t2515 VGND.t2514 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1905 XA.XIR[7].XIC[1].icell.PDM XThR.Tn[7].t49 XA.XIR[7].XIC[1].icell.Ien VGND.t1758 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1906 XA.XIR[13].XIC[6].icell.PDM XThR.Tn[13].t51 XA.XIR[13].XIC[6].icell.Ien VGND.t1035 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1907 XThR.Tn[12].t1 XThR.XTBN.Y.t83 VPWR.t311 VPWR.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1908 VGND.t2484 VPWR.t2024 XA.XIR[14].XIC_dummy_right.icell.PDM VGND.t2483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1909 Vbias.t7 Vbias.t6 VGND.t1199 VGND.t1197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.754 pd=5.78 as=0.754 ps=5.78 w=2.6 l=0.5
X1910 XA.XIR[7].XIC[5].icell.PDM XThR.Tn[6].t54 VGND.t2406 VGND.t2405 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1911 XA.XIR[5].XIC[8].icell.PUM XThC.Tn[8].t32 XA.XIR[5].XIC[8].icell.Ien VPWR.t872 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1912 XThR.Tn[12].t5 XThR.XTB5.Y a_n997_1803# VGND.t259 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1913 XA.XIR[1].XIC_15.icell.SM XA.XIR[1].XIC_15.icell.Ien Iout.t67 VGND.t806 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1914 XA.XIR[9].XIC[8].icell.PUM XThC.Tn[8].t33 XA.XIR[9].XIC[8].icell.Ien VPWR.t873 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1915 XThR.Tn[3].t1 XThR.XTB4.Y VGND.t186 VGND.t185 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X1916 XA.XIR[5].XIC[3].icell.SM XA.XIR[5].XIC[3].icell.Ien Iout.t187 VGND.t1790 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1917 VGND.t500 XThR.XTBN.Y.t84 a_n997_2667# VGND.t499 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1918 XA.XIR[9].XIC_15.icell.PDM VPWR.t2025 VGND.t2486 VGND.t2485 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1919 Vbias.t0 bias[2].t1 VPWR.t494 VPWR.t493 sky130_fd_pr__pfet_01v8 ad=0.1955 pd=1.31 as=0.2465 ps=2.28 w=0.85 l=0.5
X1920 XA.XIR[5].XIC[0].icell.PDM XThR.Tn[5].t54 XA.XIR[5].XIC[0].icell.Ien VGND.t1541 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1921 XA.XIR[8].XIC[4].icell.SM XA.XIR[8].XIC[4].icell.Ien Iout.t211 VGND.t2142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1922 XA.XIR[3].XIC_dummy_right.icell.SM XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout VGND.t1787 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1923 VGND.t2389 Vbias.t180 XA.XIR[13].XIC_15.icell.SM VGND.t2388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1924 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1538 VPWR.t1540 VPWR.t1539 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1925 XA.XIR[0].XIC[6].icell.PUM XThC.Tn[6].t34 XA.XIR[0].XIC[6].icell.Ien VPWR.t303 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1926 VGND.t2194 XThC.Tn[14].t32 XA.XIR[13].XIC[14].icell.PDM VGND.t2193 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1927 VGND.t1577 XThC.Tn[8].t34 XA.XIR[13].XIC[8].icell.PDM VGND.t1576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1928 XA.XIR[9].XIC[0].icell.PDM XThR.Tn[9].t49 XA.XIR[9].XIC[0].icell.Ien VGND.t558 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1929 Vbias.t10 bias[0].t1 VPWR.t1294 VPWR.t833 sky130_fd_pr__pfet_01v8 ad=0.12325 pd=1.14 as=0.1275 ps=1.15 w=0.85 l=2
X1930 a_5155_9615# XThC.XTB5.Y VPWR.t162 VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1931 XA.XIR[4].XIC[12].icell.PDM XThR.Tn[4].t55 XA.XIR[4].XIC[12].icell.Ien VGND.t2149 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1932 VPWR.t161 XThC.XTB5.Y XThC.Tn[12].t4 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1933 XA.XIR[3].XIC[13].icell.PDM XThR.Tn[3].t59 XA.XIR[3].XIC[13].icell.Ien VGND.t2516 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1934 VPWR.t1228 XThR.Tn[14].t52 XA.XIR[15].XIC[12].icell.PUM VPWR.t1227 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1935 XA.XIR[7].XIC_15.icell.PUM VPWR.t1536 XA.XIR[7].XIC_15.icell.Ien VPWR.t1537 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1936 VPWR.t600 XThR.Tn[13].t52 XA.XIR[14].XIC[13].icell.PUM VPWR.t599 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1937 VPWR.t1535 VPWR.t1533 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR.t1534 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1938 VGND.t1786 XThC.Tn[9].t33 XA.XIR[0].XIC[9].icell.PDM VGND.t1785 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1939 XThC.Tn[5].t8 XThC.XTBN.Y.t86 a_5949_9615# VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 XA.XIR[2].XIC[3].icell.SM XA.XIR[2].XIC[3].icell.Ien Iout.t254 VGND.t2675 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1941 XA.XIR[8].XIC[11].icell.PDM XThR.Tn[7].t50 VGND.t374 VGND.t373 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1942 VGND.t288 XThC.XTB5.Y XThC.Tn[4].t0 VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X1943 a_n1049_6405# XThR.XTBN.Y.t85 XThR.Tn[4].t1 VPWR.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X1944 VPWR.t1152 XThR.Tn[1].t49 XA.XIR[2].XIC[7].icell.PUM VPWR.t1151 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1945 VPWR.t294 XThR.Tn[0].t55 XA.XIR[1].XIC[8].icell.PUM VPWR.t293 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1946 XA.XIR[10].XIC[10].icell.SM XA.XIR[10].XIC[10].icell.Ien Iout.t129 VGND.t1340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1947 XThC.Tn[2].t8 XThC.XTBN.Y.t87 VGND.t506 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1948 VPWR.t1262 XThR.Tn[4].t56 XA.XIR[5].XIC[8].icell.PUM VPWR.t1261 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1949 XA.XIR[15].XIC[14].icell.PDM VPWR.t2026 XA.XIR[15].XIC[14].icell.Ien VGND.t2487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1950 XA.XIR[15].XIC[8].icell.PDM VPWR.t2027 XA.XIR[15].XIC[8].icell.Ien VGND.t2488 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1951 a_5155_9615# XThC.XTBN.Y.t88 XThC.Tn[4].t9 VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1952 XA.XIR[1].XIC[4].icell.PDM XThR.Tn[0].t56 VGND.t467 VGND.t466 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1953 XA.XIR[8].XIC[2].icell.PDM XThR.Tn[7].t51 VGND.t376 VGND.t375 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1954 XA.XIR[13].XIC[9].icell.PUM XThC.Tn[9].t34 XA.XIR[13].XIC[9].icell.Ien VPWR.t970 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1955 XA.XIR[7].XIC[0].icell.SM XA.XIR[7].XIC[0].icell.Ien Iout.t28 VGND.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1956 XA.XIR[6].XIC_dummy_left.icell.SM XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout VGND.t1269 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1957 VPWR.t877 XThR.XTB7.B XThR.XTB2.Y VPWR.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1958 XThC.Tn[8].t0 XThC.XTB1.Y.t15 a_7651_9569# VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1959 XA.XIR[11].XIC[3].icell.PDM XThR.Tn[10].t52 VGND.t1446 VGND.t1445 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1960 VGND.t1494 XThC.Tn[11].t32 XA.XIR[10].XIC[11].icell.PDM VGND.t1493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1961 XA.XIR[10].XIC[1].icell.SM XA.XIR[10].XIC[1].icell.Ien Iout.t200 VGND.t1915 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1962 XA.XIR[6].XIC_15.icell.PDM VPWR.t2028 VGND.t2490 VGND.t2489 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1963 VGND.t1393 XThC.XTB5.A XThC.XTB5.Y VGND.t287 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1964 VGND.t940 VGND.t938 XA.XIR[14].XIC_dummy_left.icell.SM VGND.t939 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1965 VGND.t1742 XThR.XTB7.Y XThR.Tn[6].t8 VGND.t1741 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1966 XA.XIR[4].XIC[10].icell.PDM XThR.Tn[4].t57 XA.XIR[4].XIC[10].icell.Ien VGND.t2150 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1967 XA.XIR[1].XIC[14].icell.PUM XThC.Tn[14].t33 XA.XIR[1].XIC[14].icell.Ien VPWR.t1289 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1968 XA.XIR[5].XIC[3].icell.PUM XThC.Tn[3].t33 XA.XIR[5].XIC[3].icell.Ien VPWR.t775 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1969 XA.XIR[7].XIC[0].icell.PDM XThR.Tn[6].t55 VGND.t2408 VGND.t2407 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1970 XA.XIR[2].XIC[12].icell.PDM XThR.Tn[1].t50 VGND.t1970 VGND.t1969 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1971 VPWR.t1230 XThR.Tn[14].t53 XA.XIR[15].XIC[10].icell.PUM VPWR.t1229 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1972 XA.XIR[9].XIC[3].icell.PUM XThC.Tn[3].t34 XA.XIR[9].XIC[3].icell.Ien VPWR.t1320 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1973 XA.XIR[4].XIC_15.icell.PUM VPWR.t1531 XA.XIR[4].XIC_15.icell.Ien VPWR.t1532 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1974 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[4].t58 VGND.t2152 VGND.t2151 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1975 XA.XIR[4].XIC[11].icell.SM XA.XIR[4].XIC[11].icell.Ien Iout.t143 VGND.t1453 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X1976 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR.t2029 VGND.t2492 VGND.t2491 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1977 XA.XIR[15].XIC[9].icell.Ien VPWR.t1528 VPWR.t1530 VPWR.t1529 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1978 VGND.t1289 XThC.Tn[2].t32 XA.XIR[10].XIC[2].icell.PDM VGND.t1288 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1979 XThR.Tn[9].t0 XThR.XTBN.Y.t86 VPWR.t313 VPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1980 VGND.t507 XThC.XTBN.Y.t89 a_9827_9569# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1981 XA.XIR[0].XIC[1].icell.PUM XThC.Tn[1].t35 XA.XIR[0].XIC[1].icell.Ien VPWR.t1362 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1982 VPWR.t1154 XThR.Tn[1].t51 XA.XIR[2].XIC[11].icell.PUM VPWR.t1153 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1983 VGND.t2208 XThC.Tn[3].t35 XA.XIR[13].XIC[3].icell.PDM VGND.t2207 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1984 VGND.t2494 VPWR.t2030 XA.XIR[8].XIC_15.icell.PDM VGND.t2493 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1985 VPWR.t563 XThR.Tn[8].t58 XA.XIR[9].XIC[9].icell.PUM VPWR.t562 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X1986 VGND.t4 Vbias.t181 XA.XIR[1].XIC[12].icell.SM VGND.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1987 XA.XIR[14].XIC[13].icell.Ien XThR.Tn[14].t54 VPWR.t1232 VPWR.t1231 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1988 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR.t1525 VPWR.t1527 VPWR.t1526 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1989 XA.XIR[12].XIC[14].icell.PDM XThR.Tn[12].t53 XA.XIR[12].XIC[14].icell.Ien VGND.t2198 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1990 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1523 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR.t1524 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X1991 XThC.Tn[0].t2 XThC.XTB1.Y.t16 VGND.t1103 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1992 VGND.t6 Vbias.t182 XA.XIR[0].XIC[5].icell.SM VGND.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1993 VGND.t8 Vbias.t183 XA.XIR[4].XIC[13].icell.SM VGND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X1994 XA.XIR[12].XIC[8].icell.PDM XThR.Tn[12].t54 XA.XIR[12].XIC[8].icell.Ien VGND.t2199 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X1995 VGND.t2604 XThC.Tn[4].t35 XA.XIR[0].XIC[4].icell.PDM VGND.t2603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X1996 a_10051_9569# XThC.XTB6.Y XThC.Tn[13].t0 VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1997 XA.XIR[8].XIC[6].icell.PDM XThR.Tn[7].t52 VGND.t378 VGND.t377 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X1998 XA.XIR[2].XIC[7].icell.Ien XThR.Tn[2].t49 VPWR.t1058 VPWR.t1057 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X1999 VGND.t10 Vbias.t184 XA.XIR[7].XIC[14].icell.SM VGND.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2000 XA.XIR[6].XIC_15.icell.Ien XThR.Tn[6].t56 VPWR.t1395 VPWR.t1394 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2001 VPWR.t1156 XThR.Tn[1].t52 XA.XIR[2].XIC[2].icell.PUM VPWR.t1155 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2002 XA.XIR[11].XIC[7].icell.PDM XThR.Tn[10].t53 VGND.t1448 VGND.t1447 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2003 VGND.t1942 XThC.Tn[13].t34 XA.XIR[7].XIC[13].icell.PDM VGND.t1941 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2004 VPWR.t499 XThR.Tn[0].t57 XA.XIR[1].XIC[3].icell.PUM VPWR.t498 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2005 XA.XIR[3].XIC_dummy_left.icell.SM XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout VGND.t420 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2006 XThR.Tn[14].t1 XThR.XTBN.Y.t87 VPWR.t315 VPWR.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2007 VPWR.t1264 XThR.Tn[4].t59 XA.XIR[5].XIC[3].icell.PUM VPWR.t1263 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2008 VPWR.t1522 VPWR.t1520 XA.XIR[0].XIC_15.icell.PUM VPWR.t1521 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2009 VPWR.t602 XThR.Tn[13].t53 XA.XIR[14].XIC[6].icell.PUM VPWR.t601 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2010 XA.XIR[15].XIC[3].icell.PDM VPWR.t2031 XA.XIR[15].XIC[3].icell.Ien VGND.t2495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2011 a_n997_3755# XThR.XTBN.Y.t88 VGND.t501 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2012 XThR.Tn[8].t1 XThR.XTB1.Y.t13 VPWR.t619 VPWR.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2013 XA.XIR[10].XIC_15.icell.PDM XThR.Tn[10].t54 XA.XIR[10].XIC_15.icell.Ien VGND.t1449 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2014 XA.XIR[0].XIC[14].icell.Ien XThR.Tn[0].t58 VPWR.t501 VPWR.t500 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2015 XA.XIR[2].XIC[10].icell.PDM XThR.Tn[1].t53 VGND.t1972 VGND.t1971 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2016 XA.XIR[1].XIC[8].icell.SM XA.XIR[1].XIC[8].icell.Ien Iout.t248 VGND.t2618 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2017 VGND.t12 Vbias.t185 XA.XIR[10].XIC[7].icell.SM VGND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2018 a_n1049_7787# XThR.XTB2.Y VPWR.t1165 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2019 XA.XIR[4].XIC[9].icell.SM XA.XIR[4].XIC[9].icell.Ien Iout.t23 VGND.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2020 VGND.t485 XThC.Tn[6].t35 XA.XIR[10].XIC[6].icell.PDM VGND.t484 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2021 VPWR.t1305 XThR.Tn[12].t55 XA.XIR[13].XIC[4].icell.PUM VPWR.t1304 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2022 a_n1331_2891# data[5].t4 VGND.t1252 VGND.t1251 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2023 VGND.t14 Vbias.t186 XA.XIR[13].XIC[8].icell.SM VGND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2024 XA.XIR[12].XIC[9].icell.Ien XThR.Tn[12].t56 VPWR.t1307 VPWR.t1306 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2025 VPWR.t1519 VPWR.t1517 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR.t1518 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2026 VGND.t823 XThC.Tn[7].t27 XA.XIR[13].XIC[7].icell.PDM VGND.t822 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2027 VPWR.t1234 XThR.Tn[14].t55 XA.XIR[15].XIC[5].icell.PUM VPWR.t1233 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2028 XThR.XTB7.B data[6].t1 VGND.t2186 VGND.t2185 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2029 XThR.Tn[2].t2 XThR.XTBN.Y.t89 a_n1049_7493# VPWR.t270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2030 XA.XIR[10].XIC[14].icell.PDM XThR.Tn[9].t50 VGND.t560 VGND.t559 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2031 XA.XIR[10].XIC[8].icell.PDM XThR.Tn[9].t51 VGND.t562 VGND.t561 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2032 XA.XIR[2].XIC[11].icell.Ien XThR.Tn[2].t50 VPWR.t1056 VPWR.t1055 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2033 XA.XIR[9].XIC[6].icell.SM XA.XIR[9].XIC[6].icell.Ien Iout.t145 VGND.t1455 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2034 VGND.t337 XThC.Tn[12].t34 XA.XIR[1].XIC[12].icell.PDM VGND.t336 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2035 VGND.t1944 XThC.Tn[13].t35 XA.XIR[4].XIC[13].icell.PDM VGND.t1943 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2036 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR.t2032 XA.XIR[4].XIC_dummy_left.icell.Ien VGND.t2496 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2037 XA.XIR[15].XIC[7].icell.PDM VPWR.t2033 XA.XIR[15].XIC[7].icell.Ien VGND.t2497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2038 VGND.t16 Vbias.t187 XA.XIR[0].XIC[0].icell.SM VGND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2039 XA.XIR[12].XIC[3].icell.PDM XThR.Tn[12].t57 XA.XIR[12].XIC[3].icell.Ien VGND.t2200 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2040 VPWR.t318 XThC.XTBN.Y.t90 XThC.Tn[8].t10 VPWR.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2041 XThR.Tn[10].t9 XThR.XTB3.Y.t12 VPWR.t1922 VPWR.t1170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2042 XA.XIR[7].XIC_15.icell.PDM XThR.Tn[7].t53 XA.XIR[7].XIC_15.icell.Ien VGND.t379 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2043 XA.XIR[11].XIC[4].icell.PUM XThC.Tn[4].t36 XA.XIR[11].XIC[4].icell.Ien VPWR.t1880 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2044 XThR.Tn[4].t5 XThR.XTBN.Y.t90 VGND.t423 VGND.t317 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2045 XA.XIR[15].XIC[12].icell.PUM XThC.Tn[12].t35 XA.XIR[15].XIC[12].icell.Ien VPWR.t213 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2046 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR.t1515 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR.t1516 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2047 XA.XIR[2].XIC[2].icell.Ien XThR.Tn[2].t51 VPWR.t1054 VPWR.t1053 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2048 XA.XIR[11].XIC[13].icell.SM XA.XIR[11].XIC[13].icell.Ien Iout.t96 VGND.t1136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2049 VGND.t1581 XThR.XTB7.B XThR.XTB5.Y VGND.t1580 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2050 VGND.t18 Vbias.t188 XA.XIR[12].XIC_15.icell.SM VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2051 VGND.t2170 XThC.Tn[14].t34 XA.XIR[12].XIC[14].icell.PDM VGND.t2169 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2052 XA.XIR[3].XIC[1].icell.PDM XThR.Tn[3].t60 XA.XIR[3].XIC[1].icell.Ien VGND.t2517 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2053 XA.XIR[14].XIC[6].icell.Ien XThR.Tn[14].t56 VPWR.t1236 VPWR.t1235 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2054 VGND.t2030 XThC.Tn[8].t35 XA.XIR[12].XIC[8].icell.PDM VGND.t2029 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2055 VPWR.t988 XThR.Tn[13].t54 XA.XIR[14].XIC[1].icell.PUM VPWR.t987 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2056 XA.XIR[2].XIC[7].icell.PUM XThC.Tn[7].t28 XA.XIR[2].XIC[7].icell.Ien VPWR.t603 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2057 XA.XIR[2].XIC[5].icell.PDM XThR.Tn[2].t52 XA.XIR[2].XIC[5].icell.Ien VGND.t146 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2058 VPWR.t1309 XThR.Tn[12].t58 XA.XIR[13].XIC[0].icell.PUM VPWR.t1308 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2059 VPWR.t386 XThR.Tn[9].t52 XA.XIR[10].XIC[4].icell.PUM VPWR.t385 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2060 XA.XIR[6].XIC[13].icell.PDM XThR.Tn[6].t57 XA.XIR[6].XIC[13].icell.Ien VGND.t1307 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2061 XA.XIR[1].XIC[3].icell.SM XA.XIR[1].XIC[3].icell.Ien Iout.t30 VGND.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2062 XA.XIR[14].XIC[9].icell.PDM XThR.Tn[14].t57 XA.XIR[14].XIC[9].icell.Ien VGND.t2111 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2063 VPWR.t1876 XThR.Tn[11].t58 XA.XIR[12].XIC[14].icell.PUM VPWR.t1875 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2064 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t5 VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2065 XThC.Tn[4].t8 XThC.XTBN.Y.t91 a_5155_9615# VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2066 XA.XIR[13].XIC[4].icell.Ien XThR.Tn[13].t55 VPWR.t990 VPWR.t989 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2067 VGND.t20 Vbias.t189 XA.XIR[10].XIC[2].icell.SM VGND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2068 XA.XIR[4].XIC[4].icell.SM XA.XIR[4].XIC[4].icell.Ien Iout.t186 VGND.t1789 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2069 VGND.t22 Vbias.t190 XA.XIR[9].XIC_15.icell.SM VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2070 XA.XIR[9].XIC[10].icell.SM XA.XIR[9].XIC[10].icell.Ien Iout.t243 VGND.t2555 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2071 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR.t1512 VPWR.t1514 VPWR.t1513 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2072 VGND.t575 XThC.Tn[10].t35 XA.XIR[1].XIC[10].icell.PDM VGND.t574 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2073 VGND.t24 Vbias.t191 XA.XIR[13].XIC[3].icell.SM VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2074 XA.XIR[0].XIC[12].icell.PDM XThR.Tn[0].t59 XA.XIR[0].XIC[12].icell.Ien VGND.t824 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2075 VPWR.t1403 XThR.Tn[3].t61 XA.XIR[4].XIC[8].icell.PUM VPWR.t1402 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2076 VGND.t425 XThR.XTBN.Y.t91 a_n997_1579# VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2077 VPWR.t777 XThR.Tn[10].t55 XA.XIR[11].XIC[12].icell.PUM VPWR.t776 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2078 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR.t2034 VGND.t2499 VGND.t2498 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2079 XA.XIR[12].XIC[9].icell.PUM XThC.Tn[9].t35 XA.XIR[12].XIC[9].icell.Ien VPWR.t971 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2080 XA.XIR[12].XIC[7].icell.PDM XThR.Tn[12].t59 XA.XIR[12].XIC[7].icell.Ien VGND.t2201 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2081 XA.XIR[15].XIC[10].icell.PUM XThC.Tn[10].t36 XA.XIR[15].XIC[10].icell.Ien VPWR.t392 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2082 XA.XIR[10].XIC[3].icell.PDM XThR.Tn[9].t53 VGND.t564 VGND.t563 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2083 XA.XIR[5].XIC[12].icell.SM XA.XIR[5].XIC[12].icell.Ien Iout.t5 VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2084 XA.XIR[9].XIC[1].icell.SM XA.XIR[9].XIC[1].icell.Ien Iout.t163 VGND.t1591 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2085 a_9827_9569# XThC.XTB5.Y XThC.Tn[12].t1 VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2086 XA.XIR[11].XIC[0].icell.PUM XThC.Tn[0].t32 XA.XIR[11].XIC[0].icell.Ien VPWR.t1219 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2087 XA.XIR[8].XIC[13].icell.SM XA.XIR[8].XIC[13].icell.Ien Iout.t117 VGND.t1302 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2088 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR.t1510 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR.t1511 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2089 XA.XIR[7].XIC[14].icell.SM XA.XIR[7].XIC[14].icell.Ien Iout.t250 VGND.t2644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2090 XA.XIR[2].XIC[11].icell.PUM XThC.Tn[11].t33 XA.XIR[2].XIC[11].icell.Ien VPWR.t814 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2091 XA.XIR[5].XIC[1].icell.PDM XThR.Tn[4].t60 VGND.t649 VGND.t648 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2092 XA.XIR[0].XIC[5].icell.PDM VGND.t935 VGND.t937 VGND.t936 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2093 VPWR.t388 XThR.Tn[9].t54 XA.XIR[10].XIC[0].icell.PUM VPWR.t387 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2094 XA.XIR[4].XIC[13].icell.PDM XThR.Tn[3].t62 VGND.t2519 VGND.t2518 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2095 XA.XIR[2].XIC[12].icell.SM XA.XIR[2].XIC[12].icell.Ien Iout.t116 VGND.t1301 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2096 XA.XIR[12].XIC[9].icell.PDM XThR.Tn[11].t59 VGND.t2596 VGND.t2595 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2097 VGND.t2210 XThC.Tn[3].t36 XA.XIR[12].XIC[3].icell.PDM VGND.t2209 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2098 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14].t58 VPWR.t1238 VPWR.t1237 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2099 XThR.XTBN.Y.t2 XThR.XTBN.A VPWR.t738 VPWR.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2100 VGND.t26 Vbias.t192 XA.XIR[15].XIC[11].icell.SM VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2101 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13].t56 VPWR.t992 VPWR.t991 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2102 VPWR.t227 XThR.Tn[7].t54 XA.XIR[8].XIC[9].icell.PUM VPWR.t226 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2103 VGND.t2172 XThC.Tn[14].t35 XA.XIR[6].XIC[14].icell.PDM VGND.t2171 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2104 XA.XIR[0].XIC[10].icell.PDM XThR.Tn[0].t60 XA.XIR[0].XIC[10].icell.Ien VGND.t825 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2105 XA.XIR[2].XIC[2].icell.PUM XThC.Tn[2].t33 XA.XIR[2].XIC[2].icell.Ien VPWR.t706 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2106 XA.XIR[2].XIC[0].icell.PDM XThR.Tn[2].t53 XA.XIR[2].XIC[0].icell.Ien VGND.t157 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2107 VGND.t2032 XThC.Tn[8].t36 XA.XIR[6].XIC[8].icell.PDM VGND.t2031 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2108 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR.t1507 VPWR.t1509 VPWR.t1508 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2109 VPWR.t779 XThR.Tn[10].t56 XA.XIR[11].XIC[10].icell.PUM VPWR.t778 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2110 XA.XIR[0].XIC_15.icell.PUM VPWR.t1505 XA.XIR[0].XIC_15.icell.Ien VPWR.t1506 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2111 XA.XIR[14].XIC[4].icell.PDM XThR.Tn[14].t59 XA.XIR[14].XIC[4].icell.Ien VGND.t2112 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2112 XA.XIR[1].XIC[7].icell.Ien XThR.Tn[1].t54 VPWR.t1158 VPWR.t1157 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2113 VGND.t35 Vbias.t193 XA.XIR[2].XIC[6].icell.SM VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2114 VGND.t2316 XThC.Tn[1].t36 XA.XIR[7].XIC[1].icell.PDM VGND.t2315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2115 VGND.t2281 XThC.Tn[5].t32 XA.XIR[2].XIC[5].icell.PDM VGND.t2280 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2116 VPWR.t272 XThR.XTBN.Y.t92 XThR.Tn[11].t9 VPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2117 XA.XIR[4].XIC[8].icell.Ien XThR.Tn[4].t61 VPWR.t442 VPWR.t441 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2118 XA.XIR[10].XIC[7].icell.PDM XThR.Tn[9].t55 VGND.t566 VGND.t565 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2119 VPWR.t1404 data[1].t4 XThC.XTB7.A VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2120 VPWR.t406 XThR.Tn[3].t63 XA.XIR[4].XIC[3].icell.PUM VPWR.t405 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2121 XA.XIR[11].XIC[12].icell.Ien XThR.Tn[11].t60 VPWR.t1860 VPWR.t1859 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2122 a_8739_9569# XThC.XTBN.Y.t92 VGND.t508 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2123 VGND.t1373 XThR.XTBN.A XThR.XTBN.Y.t0 VGND.t1372 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2124 XThC.Tn[6].t2 XThC.XTB7.Y VGND.t218 VGND.t217 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2125 XA.XIR[8].XIC[14].icell.PDM XThR.Tn[8].t59 XA.XIR[8].XIC[14].icell.Ien VGND.t882 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2126 XA.XIR[8].XIC[8].icell.PDM XThR.Tn[8].t60 XA.XIR[8].XIC[8].icell.Ien VGND.t883 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2127 XA.XIR[15].XIC[5].icell.PUM XThC.Tn[5].t33 XA.XIR[15].XIC[5].icell.Ien VPWR.t1349 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2128 XA.XIR[1].XIC[13].icell.PDM XThR.Tn[0].t61 VGND.t827 VGND.t826 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2129 XA.XIR[6].XIC[9].icell.PUM XThC.Tn[9].t36 XA.XIR[6].XIC[9].icell.Ien VPWR.t1031 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2130 XThR.Tn[12].t4 XThR.XTB5.Y a_n997_1803# VGND.t258 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2131 VGND.t2501 VPWR.t2035 XA.XIR[1].XIC_dummy_left.icell.PDM VGND.t2500 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2132 VGND.t37 Vbias.t194 XA.XIR[12].XIC[8].icell.SM VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2133 VGND.t1496 XThC.Tn[11].t34 XA.XIR[3].XIC[11].icell.PDM VGND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2134 VGND.t1037 XThC.Tn[7].t29 XA.XIR[12].XIC[7].icell.PDM VGND.t1036 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2135 VGND.t39 Vbias.t195 XA.XIR[15].XIC[9].icell.SM VGND.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2136 a_n997_3979# XThR.XTBN.Y.t93 VGND.t427 VGND.t426 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2137 XThC.XTB7.Y XThC.XTB7.B VGND.t1330 VGND.t1329 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2138 XA.XIR[0].XIC[0].icell.PDM VGND.t932 VGND.t934 VGND.t933 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2139 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1502 VPWR.t1504 VPWR.t1503 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2140 VGND.t41 Vbias.t196 XA.XIR[6].XIC[7].icell.SM VGND.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2141 XA.XIR[1].XIC[11].icell.Ien XThR.Tn[1].t55 VPWR.t1160 VPWR.t1159 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2142 VGND.t43 Vbias.t197 XA.XIR[2].XIC[10].icell.SM VGND.t42 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2143 XThC.Tn[8].t9 XThC.XTBN.Y.t93 VPWR.t320 VPWR.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2144 VGND.t2318 XThC.Tn[1].t37 XA.XIR[4].XIC[1].icell.PDM VGND.t2317 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2145 XA.XIR[12].XIC[4].icell.PDM XThR.Tn[11].t61 VGND.t2590 VGND.t2589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2146 VGND.t1607 XThC.Tn[2].t34 XA.XIR[3].XIC[2].icell.PDM VGND.t1606 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2147 VGND.t45 Vbias.t198 XA.XIR[9].XIC[8].icell.SM VGND.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2148 XA.XIR[14].XIC[7].icell.PUM XThC.Tn[7].t30 XA.XIR[14].XIC[7].icell.Ien VPWR.t604 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2149 XA.XIR[8].XIC[9].icell.Ien XThR.Tn[8].t61 VPWR.t565 VPWR.t564 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2150 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR.t2036 VGND.t2503 VGND.t2502 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2151 VGND.t2212 XThC.Tn[3].t37 XA.XIR[6].XIC[3].icell.PDM VGND.t2211 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2152 XA.XIR[5].XIC[11].icell.PDM XThR.Tn[5].t55 XA.XIR[5].XIC[11].icell.Ien VGND.t1542 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2153 XA.XIR[11].XIC[10].icell.Ien XThR.Tn[11].t62 VPWR.t1862 VPWR.t1861 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2154 a_n1049_6699# XThR.XTB4.Y VPWR.t81 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2155 XA.XIR[13].XIC_15.icell.SM XA.XIR[13].XIC_15.icell.Ien Iout.t41 VGND.t268 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2156 VPWR.t569 VGND.t2700 Vbias.t2 VPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.2465 pd=2.28 as=0.12325 ps=1.14 w=0.85 l=2
X2157 VPWR.t781 XThR.Tn[10].t57 XA.XIR[11].XIC[5].icell.PUM VPWR.t780 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2158 XA.XIR[9].XIC[11].icell.PDM XThR.Tn[9].t56 XA.XIR[9].XIC[11].icell.Ien VGND.t567 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2159 XA.XIR[10].XIC[4].icell.PUM XThC.Tn[4].t37 XA.XIR[10].XIC[4].icell.Ien VPWR.t1881 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2160 XA.XIR[1].XIC[2].icell.Ien XThR.Tn[1].t56 VPWR.t709 VPWR.t708 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2161 VGND.t47 Vbias.t199 XA.XIR[2].XIC[1].icell.SM VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2162 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1500 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR.t1501 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2163 XA.XIR[6].XIC[5].icell.SM XA.XIR[6].XIC[5].icell.Ien Iout.t112 VGND.t1278 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2164 VGND.t1478 XThC.Tn[0].t33 XA.XIR[2].XIC[0].icell.PDM VGND.t1477 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2165 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR.t1498 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR.t1499 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2166 XA.XIR[4].XIC[3].icell.Ien XThR.Tn[4].t62 VPWR.t444 VPWR.t443 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2167 VGND.t49 Vbias.t200 XA.XIR[0].XIC[14].icell.SM VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2168 VGND.t51 Vbias.t201 XA.XIR[14].XIC[5].icell.SM VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2169 VGND.t1946 XThC.Tn[13].t36 XA.XIR[0].XIC[13].icell.PDM VGND.t1945 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2170 XA.XIR[6].XIC[1].icell.PDM XThR.Tn[6].t58 XA.XIR[6].XIC[1].icell.Ien VGND.t1308 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2171 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR.t2037 XA.XIR[0].XIC_dummy_left.icell.Ien VGND.t1643 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2172 XA.XIR[1].XIC[5].icell.PDM XThR.Tn[1].t57 XA.XIR[1].XIC[5].icell.Ien VGND.t1291 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2173 XA.XIR[5].XIC[2].icell.PDM XThR.Tn[5].t56 XA.XIR[5].XIC[2].icell.Ien VGND.t1543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2174 VGND.t1645 VPWR.t2038 XA.XIR[13].XIC_dummy_right.icell.PDM VGND.t1644 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2175 XA.XIR[9].XIC[2].icell.PDM XThR.Tn[9].t57 XA.XIR[9].XIC[2].icell.Ien VGND.t568 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2176 XA.XIR[8].XIC[3].icell.PDM XThR.Tn[8].t62 XA.XIR[8].XIC[3].icell.Ien VGND.t884 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2177 XA.XIR[3].XIC_15.icell.PDM XThR.Tn[3].t64 XA.XIR[3].XIC_15.icell.Ien VGND.t599 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2178 VGND.t843 data[1].t5 XThC.XTB6.A VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2179 VPWR.t1240 XThR.Tn[14].t60 XA.XIR[15].XIC[14].icell.PUM VPWR.t1239 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2180 VPWR.t1497 VPWR.t1495 XA.XIR[14].XIC_15.icell.PUM VPWR.t1496 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2181 a_n997_2891# XThR.XTBN.Y.t94 VGND.t429 VGND.t428 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2182 VGND.t53 Vbias.t202 XA.XIR[12].XIC[3].icell.SM VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2183 VGND.t55 Vbias.t203 XA.XIR[3].XIC[7].icell.SM VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2184 VGND.t487 XThC.Tn[6].t36 XA.XIR[3].XIC[6].icell.PDM VGND.t486 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2185 XA.XIR[14].XIC[11].icell.PUM XThC.Tn[11].t35 XA.XIR[14].XIC[11].icell.Ien VPWR.t815 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2186 VPWR.t850 XThR.Tn[5].t57 XA.XIR[6].XIC[4].icell.PUM VPWR.t849 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2187 VPWR.t1494 VPWR.t1492 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1493 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2188 VGND.t57 Vbias.t204 XA.XIR[15].XIC[4].icell.SM VGND.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2189 VGND.t931 VGND.t929 XA.XIR[10].XIC_dummy_right.icell.SM VGND.t930 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2190 VGND.t1039 XThC.Tn[7].t31 XA.XIR[6].XIC[7].icell.PDM VGND.t1038 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2191 VPWR.t1491 VPWR.t1489 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR.t1490 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2192 VPWR.t1311 XThR.Tn[12].t60 XA.XIR[13].XIC[13].icell.PUM VPWR.t1310 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2193 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR.t2039 XA.XIR[15].XIC_dummy_right.icell.Ien VGND.t1646 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2194 XThR.Tn[11].t1 XThR.XTB4.Y a_n997_2667# VGND.t184 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2195 VGND.t1349 Vbias.t205 XA.XIR[6].XIC[2].icell.SM VGND.t1348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2196 XA.XIR[7].XIC[11].icell.PDM XThR.Tn[6].t59 VGND.t1310 VGND.t1309 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2197 VPWR.t159 XThC.XTB5.Y a_5155_9615# VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2198 XA.XIR[10].XIC[0].icell.PUM XThC.Tn[0].t34 XA.XIR[10].XIC[0].icell.Ien VPWR.t809 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2199 XA.XIR[3].XIC[5].icell.SM XA.XIR[3].XIC[5].icell.Ien Iout.t126 VGND.t1337 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2200 XA.XIR[3].XIC[8].icell.PDM XThR.Tn[2].t54 VGND.t156 VGND.t155 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2201 XA.XIR[3].XIC[14].icell.PDM XThR.Tn[2].t55 VGND.t154 VGND.t153 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2202 VGND.t1351 Vbias.t206 XA.XIR[9].XIC[3].icell.SM VGND.t1350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2203 XA.XIR[14].XIC[2].icell.PUM XThC.Tn[2].t35 XA.XIR[14].XIC[2].icell.Ien VPWR.t911 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2204 XA.XIR[5].XIC[6].icell.PDM XThR.Tn[5].t58 XA.XIR[5].XIC[6].icell.Ien VGND.t2550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2205 XA.XIR[11].XIC[5].icell.Ien XThR.Tn[11].t63 VPWR.t1864 VPWR.t1863 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2206 XA.XIR[4].XIC[1].icell.PDM XThR.Tn[3].t65 VGND.t601 VGND.t600 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2207 XA.XIR[9].XIC[6].icell.PDM XThR.Tn[9].t58 XA.XIR[9].XIC[6].icell.Ien VGND.t569 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2208 VGND.t2283 XThC.Tn[5].t34 XA.XIR[14].XIC[5].icell.PDM VGND.t2282 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2209 XA.XIR[8].XIC[7].icell.PDM XThR.Tn[8].t63 XA.XIR[8].XIC[7].icell.Ien VGND.t885 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2210 VGND.t431 XThR.XTBN.Y.t95 XThR.Tn[0].t6 VGND.t430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2211 XA.XIR[7].XIC[2].icell.PDM XThR.Tn[6].t60 VGND.t1312 VGND.t1311 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2212 XA.XIR[1].XIC[8].icell.PUM XThC.Tn[8].t37 XA.XIR[1].XIC[8].icell.Ien VPWR.t1191 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2213 a_n1049_6405# XThR.XTB5.Y VPWR.t1891 VPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2214 XA.XIR[6].XIC[0].icell.SM XA.XIR[6].XIC[0].icell.Ien Iout.t133 VGND.t1400 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2215 XThR.Tn[8].t2 XThR.XTB1.Y.t14 VPWR.t621 VPWR.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2216 XA.XIR[1].XIC[12].icell.SM XA.XIR[1].XIC[12].icell.Ien Iout.t166 VGND.t1615 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2217 XA.XIR[8].XIC[12].icell.PUM XThC.Tn[12].t36 XA.XIR[8].XIC[12].icell.Ien VPWR.t214 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2218 VGND.t1353 Vbias.t207 XA.XIR[14].XIC[0].icell.SM VGND.t1352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2219 XA.XIR[15].XIC[9].icell.PDM XThR.Tn[14].t61 VGND.t2114 VGND.t2113 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2220 XA.XIR[4].XIC[13].icell.SM XA.XIR[4].XIC[13].icell.Ien Iout.t52 VGND.t524 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2221 XA.XIR[5].XIC_15.icell.PDM VPWR.t2040 VGND.t1648 VGND.t1647 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2222 VGND.t1355 Vbias.t208 XA.XIR[5].XIC_15.icell.SM VGND.t1354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2223 XA.XIR[11].XIC[13].icell.PUM XThC.Tn[13].t37 XA.XIR[11].XIC[13].icell.Ien VPWR.t1134 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2224 VGND.t2034 XThC.Tn[8].t38 XA.XIR[5].XIC[8].icell.PDM VGND.t2033 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2225 VGND.t2174 XThC.Tn[14].t36 XA.XIR[5].XIC[14].icell.PDM VGND.t2173 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2226 XA.XIR[1].XIC[0].icell.PDM XThR.Tn[1].t58 XA.XIR[1].XIC[0].icell.Ien VGND.t1292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2227 VGND.t1357 Vbias.t209 XA.XIR[13].XIC[12].icell.SM VGND.t1356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2228 XThR.Tn[1].t9 XThR.XTB2.Y VGND.t1978 VGND.t1555 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2229 VGND.t2176 XThC.Tn[14].t37 XA.XIR[9].XIC[14].icell.PDM VGND.t2175 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2230 VGND.t2036 XThC.Tn[8].t39 XA.XIR[9].XIC[8].icell.PDM VGND.t2035 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2231 VPWR.t1816 XThR.Tn[5].t59 XA.XIR[6].XIC[0].icell.PUM VPWR.t1815 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2232 VGND.t678 XThC.XTBN.Y.t94 a_8739_9569# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2233 XA.XIR[14].XIC_15.icell.Ien XThR.Tn[14].t62 VPWR.t1242 VPWR.t1241 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2234 VGND.t1359 Vbias.t210 XA.XIR[1].XIC[6].icell.SM VGND.t1358 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2235 VPWR.t1488 VPWR.t1486 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR.t1487 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2236 XThC.Tn[1].t2 XThC.XTB2.Y VGND.t208 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2237 VGND.t216 XThC.XTB7.Y XThC.Tn[6].t1 VGND.t215 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2238 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR.t2041 XA.XIR[12].XIC_dummy_right.icell.Ien VGND.t1649 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2239 VPWR.t390 XThR.Tn[9].t59 XA.XIR[10].XIC[13].icell.PUM VPWR.t389 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2240 VPWR.t1485 VPWR.t1483 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1484 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2241 a_6243_9615# XThC.XTBN.Y.t95 XThC.Tn[6].t5 VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2242 VGND.t1361 Vbias.t211 XA.XIR[3].XIC[2].icell.SM VGND.t1360 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2243 VGND.t1363 Vbias.t212 XA.XIR[11].XIC[11].icell.SM VGND.t1362 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2244 XA.XIR[10].XIC[12].icell.Ien XThR.Tn[10].t58 VPWR.t549 VPWR.t548 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2245 XThR.Tn[2].t3 XThR.XTBN.Y.t96 a_n1049_7493# VPWR.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2246 VGND.t1651 VPWR.t2042 XA.XIR[7].XIC_15.icell.PDM VGND.t1650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2247 XA.XIR[10].XIC[7].icell.SM XA.XIR[10].XIC[7].icell.Ien Iout.t155 VGND.t1525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2248 XA.XIR[13].XIC[13].icell.Ien XThR.Tn[13].t57 VPWR.t994 VPWR.t993 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2249 XA.XIR[13].XIC[8].icell.SM XA.XIR[13].XIC[8].icell.Ien Iout.t161 VGND.t1537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2250 XA.XIR[1].XIC[1].icell.PDM XThR.Tn[0].t62 VGND.t829 VGND.t828 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2251 XThR.Tn[13].t8 XThR.XTBN.Y.t97 VPWR.t273 VPWR.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2252 XA.XIR[5].XIC[9].icell.PUM XThC.Tn[9].t37 XA.XIR[5].XIC[9].icell.Ien VPWR.t1032 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2253 XA.XIR[7].XIC[6].icell.PDM XThR.Tn[6].t61 VGND.t1314 VGND.t1313 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2254 XA.XIR[0].XIC[8].icell.Ien XThR.Tn[0].t63 VPWR.t503 VPWR.t502 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2255 XA.XIR[3].XIC[0].icell.SM XA.XIR[3].XIC[0].icell.Ien Iout.t89 VGND.t1118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2256 XA.XIR[9].XIC[9].icell.PUM XThC.Tn[9].t38 XA.XIR[9].XIC[9].icell.Ien VPWR.t1033 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2257 XA.XIR[3].XIC[3].icell.PDM XThR.Tn[2].t56 VGND.t152 VGND.t151 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2258 XThR.Tn[10].t10 XThR.XTB3.Y.t13 VPWR.t1923 VPWR.t1168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2259 XA.XIR[8].XIC[10].icell.PUM XThC.Tn[10].t37 XA.XIR[8].XIC[10].icell.Ien VPWR.t393 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2260 XThR.Tn[4].t4 XThR.XTBN.Y.t98 VGND.t432 VGND.t323 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2261 VPWR.t1313 XThR.Tn[12].t61 XA.XIR[13].XIC[6].icell.PUM VPWR.t1312 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2262 VGND.t928 VGND.t926 XA.XIR[10].XIC_dummy_left.icell.SM VGND.t927 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2263 VGND.t255 XThR.XTB6.Y XThR.Tn[5].t0 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2264 VGND.t1480 XThC.Tn[0].t35 XA.XIR[14].XIC[0].icell.PDM VGND.t1479 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2265 XA.XIR[1].XIC[3].icell.PUM XThC.Tn[3].t38 XA.XIR[1].XIC[3].icell.Ien VPWR.t1321 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2266 VGND.t1365 Vbias.t213 XA.XIR[1].XIC[10].icell.SM VGND.t1364 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2267 a_4861_9615# XThC.XTBN.Y.t96 XThC.Tn[3].t5 VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2268 XA.XIR[15].XIC[4].icell.PDM XThR.Tn[14].t63 VGND.t2116 VGND.t2115 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2269 XA.XIR[0].XIC[11].icell.SM XA.XIR[0].XIC[11].icell.Ien Iout.t47 VGND.t419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2270 XA.XIR[14].XIC[5].icell.PDM XThR.Tn[13].t58 VGND.t1818 VGND.t1817 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2271 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR.t2043 VGND.t1653 VGND.t1652 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2272 a_n997_3755# XThR.XTB2.Y XThR.Tn[9].t4 VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2273 VGND.t2214 XThC.Tn[3].t39 XA.XIR[5].XIC[3].icell.PDM VGND.t2213 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2274 VGND.t1367 Vbias.t214 XA.XIR[11].XIC[9].icell.SM VGND.t1366 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2275 XA.XIR[10].XIC[10].icell.Ien XThR.Tn[10].t59 VPWR.t551 VPWR.t550 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2276 XA.XIR[12].XIC_15.icell.SM XA.XIR[12].XIC_15.icell.Ien Iout.t207 VGND.t1956 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2277 VGND.t2216 XThC.Tn[3].t40 XA.XIR[9].XIC[3].icell.PDM VGND.t2215 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2278 VGND.t1369 Vbias.t215 XA.XIR[8].XIC[11].icell.SM VGND.t1368 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2279 XA.XIR[7].XIC[12].icell.Ien XThR.Tn[7].t55 VPWR.t229 VPWR.t228 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2280 VPWR.t643 XThR.Tn[0].t64 XA.XIR[1].XIC[9].icell.PUM VPWR.t642 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2281 VGND.t1655 VPWR.t2044 XA.XIR[4].XIC_15.icell.PDM VGND.t1654 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2282 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR.t1480 VPWR.t1482 VPWR.t1481 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2283 VGND.t1371 Vbias.t216 XA.XIR[1].XIC[1].icell.SM VGND.t1370 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2284 VPWR.t446 XThR.Tn[4].t63 XA.XIR[5].XIC[9].icell.PUM VPWR.t445 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2285 VGND.t2320 XThC.Tn[1].t38 XA.XIR[0].XIC[1].icell.PDM VGND.t2319 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2286 XA.XIR[11].XIC[6].icell.PUM XThC.Tn[6].t37 XA.XIR[11].XIC[6].icell.Ien VPWR.t304 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2287 XA.XIR[15].XIC[14].icell.PUM XThC.Tn[14].t38 XA.XIR[15].XIC[14].icell.Ien VPWR.t1290 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2288 XA.XIR[3].XIC[7].icell.PDM XThR.Tn[2].t57 VGND.t150 VGND.t149 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2289 XA.XIR[14].XIC[13].icell.PDM XThR.Tn[14].t64 XA.XIR[14].XIC[13].icell.Ien VGND.t2117 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2290 VGND.t1657 VPWR.t2045 XA.XIR[12].XIC_dummy_right.icell.PDM VGND.t1656 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2291 XA.XIR[10].XIC[2].icell.SM XA.XIR[10].XIC[2].icell.Ien Iout.t235 VGND.t2523 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2292 VGND.t1867 XThC.Tn[9].t39 XA.XIR[11].XIC[9].icell.PDM VGND.t1866 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2293 VPWR.t1924 XThR.XTB3.Y.t14 a_n1049_7493# VPWR.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2294 XA.XIR[13].XIC[3].icell.SM XA.XIR[13].XIC[3].icell.Ien Iout.t190 VGND.t1798 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2295 VPWR.t355 XThR.Tn[9].t60 XA.XIR[10].XIC[6].icell.PUM VPWR.t354 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2296 XA.XIR[6].XIC_15.icell.PDM XThR.Tn[6].t62 XA.XIR[6].XIC_15.icell.Ien VGND.t1315 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2297 VPWR.t1866 XThR.Tn[11].t64 XA.XIR[12].XIC[8].icell.PUM VPWR.t1865 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2298 XA.XIR[0].XIC[3].icell.Ien XThR.Tn[0].t65 VPWR.t645 VPWR.t644 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2299 XA.XIR[8].XIC[5].icell.PUM XThC.Tn[5].t35 XA.XIR[8].XIC[5].icell.Ien VPWR.t1350 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2300 XA.XIR[13].XIC[6].icell.Ien XThR.Tn[13].t59 VPWR.t996 VPWR.t995 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2301 XA.XIR[0].XIC[9].icell.SM XA.XIR[0].XIC[9].icell.Ien Iout.t62 VGND.t677 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2302 VGND.t2220 Vbias.t217 XA.XIR[5].XIC[8].icell.SM VGND.t2219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2303 VGND.t1041 XThC.Tn[7].t32 XA.XIR[5].XIC[7].icell.PDM VGND.t1040 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2304 VPWR.t1315 XThR.Tn[12].t62 XA.XIR[13].XIC[1].icell.PUM VPWR.t1314 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2305 XThC.XTB2.Y XThC.XTB6.A a_3523_10575# VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2306 VPWR.t1479 VPWR.t1477 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR.t1478 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2307 VGND.t1960 XThC.Tn[7].t33 XA.XIR[9].XIC[7].icell.PDM VGND.t1959 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2308 VGND.t2222 Vbias.t218 XA.XIR[8].XIC[9].icell.SM VGND.t2221 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2309 XA.XIR[7].XIC[10].icell.Ien XThR.Tn[7].t56 VPWR.t231 VPWR.t230 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2310 XThR.Tn[4].t9 XThR.XTB5.Y VGND.t2651 VGND.t256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2311 VPWR.t274 XThR.XTBN.Y.t99 XThR.Tn[14].t0 VPWR.t198 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2312 VPWR.t553 XThR.Tn[10].t60 XA.XIR[11].XIC[14].icell.PUM VPWR.t552 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2313 XThC.Tn[13].t5 XThC.XTB6.Y VPWR.t765 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2314 XA.XIR[13].XIC[9].icell.PDM XThR.Tn[13].t60 XA.XIR[13].XIC[9].icell.Ien VGND.t1805 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2315 VGND.t1395 XThC.XTB6.Y XThC.Tn[5].t0 VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2316 XA.XIR[14].XIC[0].icell.PDM XThR.Tn[13].t61 VGND.t1807 VGND.t1806 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2317 XA.XIR[5].XIC[6].icell.SM XA.XIR[5].XIC[6].icell.Ien Iout.t94 VGND.t1128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2318 VPWR.t276 XThR.XTBN.Y.t100 XThR.Tn[11].t8 VPWR.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2319 VGND.t2224 Vbias.t219 XA.XIR[11].XIC[4].icell.SM VGND.t2223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2320 XA.XIR[10].XIC[5].icell.Ien XThR.Tn[10].t61 VPWR.t555 VPWR.t554 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2321 XA.XIR[13].XIC[12].icell.PDM XThR.Tn[12].t63 VGND.t2203 VGND.t2202 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2322 VGND.t925 VGND.t923 XA.XIR[6].XIC_dummy_right.icell.SM VGND.t924 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2323 XA.XIR[12].XIC[13].icell.PDM XThR.Tn[11].t65 VGND.t2592 VGND.t2591 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2324 XA.XIR[15].XIC[11].icell.SM XA.XIR[15].XIC[11].icell.Ien Iout.t242 VGND.t2554 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2325 XA.XIR[2].XIC[11].icell.PDM XThR.Tn[2].t58 XA.XIR[2].XIC[11].icell.Ien VGND.t148 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2326 XA.XIR[3].XIC[4].icell.PUM XThC.Tn[4].t38 XA.XIR[3].XIC[4].icell.Ien VPWR.t851 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2327 XThC.Tn[9].t4 XThC.XTB2.Y a_7875_9569# VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2328 XA.XIR[4].XIC_15.icell.PDM VPWR.t2046 VGND.t1659 VGND.t1658 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2329 XA.XIR[11].XIC[1].icell.PUM XThC.Tn[1].t39 XA.XIR[11].XIC[1].icell.Ien VPWR.t1207 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2330 VGND.t2605 XThC.XTB6.A XThC.XTB6.Y VGND.t1333 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2331 VGND.t206 XThC.XTB2.Y XThC.Tn[1].t1 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2332 XA.XIR[10].XIC[13].icell.PUM XThC.Tn[13].t38 XA.XIR[10].XIC[13].icell.Ien VPWR.t1135 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2333 XA.XIR[2].XIC[6].icell.SM XA.XIR[2].XIC[6].icell.Ien Iout.t201 VGND.t1923 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2334 VGND.t2226 Vbias.t220 XA.XIR[12].XIC[12].icell.SM VGND.t2225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2335 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR.t1475 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR.t1476 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2336 XThC.Tn[6].t4 XThC.XTBN.Y.t97 a_6243_9615# VPWR.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2337 XA.XIR[6].XIC[14].icell.SM XA.XIR[6].XIC[14].icell.Ien Iout.t22 VGND.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2338 VGND.t2228 Vbias.t221 XA.XIR[15].XIC[13].icell.SM VGND.t2227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2339 VGND.t2230 Vbias.t222 XA.XIR[14].XIC[14].icell.SM VGND.t2229 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2340 VGND.t339 XThC.Tn[12].t37 XA.XIR[15].XIC[12].icell.PDM VGND.t338 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2341 VGND.t1545 XThC.Tn[4].t39 XA.XIR[11].XIC[4].icell.PDM VGND.t1544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2342 XA.XIR[2].XIC[2].icell.PDM XThR.Tn[2].t59 XA.XIR[2].XIC[2].icell.Ien VGND.t147 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2343 VPWR.t943 XThR.XTB7.Y a_n1049_5317# VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2344 VPWR.t357 XThR.Tn[9].t61 XA.XIR[10].XIC[1].icell.PUM VPWR.t356 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2345 VGND.t1661 VPWR.t2047 XA.XIR[6].XIC_dummy_right.icell.PDM VGND.t1660 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2346 VPWR.t764 XThC.XTB6.Y XThC.Tn[13].t4 VPWR.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2347 VPWR.t1868 XThR.Tn[11].t66 XA.XIR[12].XIC[3].icell.PUM VPWR.t1867 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2348 a_n997_3979# XThR.XTBN.Y.t101 VGND.t434 VGND.t433 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2349 XA.XIR[5].XIC[4].icell.Ien XThR.Tn[5].t60 VPWR.t1818 VPWR.t1817 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2350 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13].t62 VPWR.t980 VPWR.t979 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2351 XA.XIR[9].XIC[4].icell.Ien XThR.Tn[9].t62 VPWR.t359 VPWR.t358 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2352 XA.XIR[0].XIC[4].icell.SM XA.XIR[0].XIC[4].icell.Ien Iout.t71 VGND.t844 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2353 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR.t1472 VPWR.t1474 VPWR.t1473 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2354 VGND.t2232 Vbias.t223 XA.XIR[5].XIC[3].icell.SM VGND.t2231 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2355 VGND.t2234 Vbias.t224 XA.XIR[9].XIC[12].icell.SM VGND.t2233 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2356 XA.XIR[9].XIC[7].icell.SM XA.XIR[9].XIC[7].icell.Ien Iout.t164 VGND.t1613 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2357 VGND.t183 XThR.XTB4.Y XThR.Tn[3].t0 VGND.t182 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2358 XA.XIR[5].XIC[10].icell.SM XA.XIR[5].XIC[10].icell.Ien Iout.t40 VGND.t267 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2359 a_7331_10587# data[0].t2 VPWR.t918 VPWR.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2360 a_4067_9615# XThC.XTBN.Y.t98 XThC.Tn[2].t5 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2361 VPWR.t1052 XThR.Tn[2].t60 XA.XIR[3].XIC[12].icell.PUM VPWR.t1051 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2362 XA.XIR[13].XIC[10].icell.PDM XThR.Tn[12].t64 VGND.t2205 VGND.t2204 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2363 XA.XIR[12].XIC[8].icell.SM XA.XIR[12].XIC[8].icell.Ien Iout.t255 VGND.t2682 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2364 XA.XIR[11].XIC[14].icell.Ien XThR.Tn[11].t67 VPWR.t1016 VPWR.t1015 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2365 VGND.t2236 Vbias.t225 XA.XIR[8].XIC[4].icell.SM VGND.t2235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2366 VGND.t922 VGND.t920 XA.XIR[3].XIC_dummy_right.icell.SM VGND.t921 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2367 XA.XIR[7].XIC[5].icell.Ien XThR.Tn[7].t57 VPWR.t219 VPWR.t218 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2368 VPWR.t711 XThR.Tn[6].t63 XA.XIR[7].XIC[12].icell.PUM VPWR.t710 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2369 XA.XIR[13].XIC[4].icell.PDM XThR.Tn[13].t63 XA.XIR[13].XIC[4].icell.Ien VGND.t1808 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2370 XA.XIR[15].XIC[9].icell.SM XA.XIR[15].XIC[9].icell.Ien Iout.t238 VGND.t2537 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2371 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR.t2048 XA.XIR[8].XIC_dummy_right.icell.Ien VGND.t1662 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2372 VPWR.t1820 XThR.Tn[5].t61 XA.XIR[6].XIC[13].icell.PUM VPWR.t1819 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2373 a_n1049_6699# XThR.XTBN.Y.t102 XThR.Tn[3].t8 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2374 VGND.t1198 Vbias.t4 Vbias.t5 VGND.t1197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.754 pd=5.78 as=0.754 ps=5.78 w=2.6 l=0.5
X2375 XA.XIR[0].XIC[11].icell.PDM VGND.t917 VGND.t919 VGND.t918 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2376 XA.XIR[3].XIC[0].icell.PUM XThC.Tn[0].t36 XA.XIR[3].XIC[0].icell.Ien VPWR.t810 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2377 XA.XIR[1].XIC_15.icell.PDM VPWR.t2049 VGND.t1664 VGND.t1663 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2378 XA.XIR[5].XIC[1].icell.SM XA.XIR[5].XIC[1].icell.Ien Iout.t253 VGND.t2654 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2379 XA.XIR[2].XIC[10].icell.SM XA.XIR[2].XIC[10].icell.Ien Iout.t237 VGND.t2535 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2380 XThC.Tn[3].t4 XThC.XTBN.Y.t99 a_4861_9615# VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2381 XA.XIR[3].XIC[14].icell.SM XA.XIR[3].XIC[14].icell.Ien Iout.t46 VGND.t388 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2382 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR.t1470 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR.t1471 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2383 XThC.XTB5.A data[0].t3 VGND.t1621 VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2384 VGND.t577 XThC.Tn[10].t38 XA.XIR[15].XIC[10].icell.PDM VGND.t576 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2385 VPWR.t79 XThR.XTB4.Y XThR.Tn[11].t5 VPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2386 XA.XIR[2].XIC[6].icell.PDM XThR.Tn[2].t61 XA.XIR[2].XIC[6].icell.Ien VGND.t125 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2387 XA.XIR[0].XIC[2].icell.PDM VGND.t914 VGND.t916 VGND.t915 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2388 XA.XIR[2].XIC[1].icell.SM XA.XIR[2].XIC[1].icell.Ien Iout.t130 VGND.t1392 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2389 VGND.t1498 XThC.Tn[11].t36 XA.XIR[2].XIC[11].icell.PDM VGND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2390 VGND.t452 XThR.XTBN.Y.t103 a_n997_715# VGND.t451 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2391 a_n997_2891# XThR.XTBN.Y.t104 VGND.t454 VGND.t453 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2392 XA.XIR[8].XIC[9].icell.PDM XThR.Tn[7].t58 VGND.t367 VGND.t366 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2393 VGND.t913 VGND.t911 XA.XIR[6].XIC_dummy_left.icell.SM VGND.t912 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2394 XA.XIR[5].XIC[0].icell.Ien XThR.Tn[5].t62 VPWR.t1822 VPWR.t1821 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2395 VPWR.t408 XThR.Tn[3].t66 XA.XIR[4].XIC[9].icell.PUM VPWR.t407 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2396 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9].t63 VPWR.t361 VPWR.t360 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2397 VPWR.t1050 XThR.Tn[2].t62 XA.XIR[3].XIC[10].icell.PUM VPWR.t1049 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2398 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR.t1467 VPWR.t1469 VPWR.t1468 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2399 VPWR.t713 XThR.Tn[6].t64 XA.XIR[7].XIC[10].icell.PUM VPWR.t712 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2400 XA.XIR[14].XIC[1].icell.PDM XThR.Tn[14].t65 XA.XIR[14].XIC[1].icell.Ien VGND.t2118 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2401 XA.XIR[10].XIC[6].icell.PUM XThC.Tn[6].t38 XA.XIR[10].XIC[6].icell.Ien VPWR.t305 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2402 XThR.Tn[11].t0 XThR.XTB4.Y a_n997_2667# VGND.t181 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2403 VPWR.t1466 VPWR.t1464 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1465 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2404 VGND.t1609 XThC.Tn[2].t36 XA.XIR[2].XIC[2].icell.PDM VGND.t1608 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2405 XA.XIR[13].XIC[7].icell.PUM XThC.Tn[7].t34 XA.XIR[13].XIC[7].icell.Ien VPWR.t1138 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2406 XA.XIR[9].XIC[2].icell.SM XA.XIR[9].XIC[2].icell.Ien Iout.t115 VGND.t1300 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2407 VPWR.t103 XThC.XTB2.Y XThC.Tn[9].t0 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2408 XA.XIR[3].XIC[12].icell.Ien XThR.Tn[3].t67 VPWR.t410 VPWR.t409 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2409 a_n997_3979# XThR.XTB1.Y.t15 XThR.Tn[8].t3 VGND.t1098 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2410 VGND.t1666 VPWR.t2050 XA.XIR[0].XIC_15.icell.PDM VGND.t1665 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2411 VGND.t1869 XThC.Tn[9].t40 XA.XIR[10].XIC[9].icell.PDM VGND.t1868 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2412 XA.XIR[12].XIC[3].icell.SM XA.XIR[12].XIC[3].icell.Ien Iout.t234 VGND.t2522 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2413 VPWR.t473 XThC.XTBN.Y.t100 XThC.Tn[8].t8 VPWR.t472 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2414 XA.XIR[15].XIC[4].icell.SM XA.XIR[15].XIC[4].icell.Ien Iout.t32 VGND.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2415 XA.XIR[4].XIC[8].icell.PDM XThR.Tn[4].t64 XA.XIR[4].XIC[8].icell.Ien VGND.t650 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2416 XA.XIR[4].XIC[14].icell.PDM XThR.Tn[4].t65 XA.XIR[4].XIC[14].icell.Ien VGND.t651 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2417 XA.XIR[10].XIC_dummy_right.icell.SM XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout VGND.t846 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2418 a_n1335_8331# XThR.XTB5.A XThR.XTB1.Y.t1 VGND.t1633 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2419 VPWR.t19 XThR.Tn[14].t66 XA.XIR[15].XIC[8].icell.PUM VPWR.t18 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2420 XA.XIR[0].XIC[6].icell.PDM VGND.t908 VGND.t910 VGND.t909 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2421 XA.XIR[11].XIC[12].icell.PDM XThR.Tn[11].t68 XA.XIR[11].XIC[12].icell.Ien VGND.t1831 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2422 a_n1049_6405# XThR.XTBN.Y.t105 XThR.Tn[4].t0 VPWR.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2423 XA.XIR[15].XIC[7].icell.Ien VPWR.t1461 VPWR.t1463 VPWR.t1462 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2424 XThR.Tn[7].t4 XThR.XTBN.Y.t106 VPWR.t281 VPWR.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2425 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR.t2051 VGND.t1668 VGND.t1667 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2426 VPWR.t1824 XThR.Tn[5].t63 XA.XIR[6].XIC[6].icell.PUM VPWR.t1823 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2427 VGND.t907 VGND.t905 XA.XIR[3].XIC_dummy_left.icell.SM VGND.t906 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2428 VPWR.t795 XThR.Tn[8].t64 XA.XIR[9].XIC[7].icell.PUM VPWR.t794 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2429 XThC.Tn[9].t8 XThC.XTBN.Y.t101 VPWR.t474 VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2430 XThR.Tn[1].t5 XThR.XTBN.Y.t107 VGND.t456 VGND.t455 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2431 VPWR.t1460 VPWR.t1458 XA.XIR[13].XIC_15.icell.PUM VPWR.t1459 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2432 VGND.t2238 Vbias.t226 XA.XIR[2].XIC[7].icell.SM VGND.t2237 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2433 VGND.t489 XThC.Tn[6].t39 XA.XIR[2].XIC[6].icell.PDM VGND.t488 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2434 XA.XIR[13].XIC[11].icell.PUM XThC.Tn[11].t37 XA.XIR[13].XIC[11].icell.Ien VPWR.t816 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2435 XA.XIR[12].XIC[1].icell.PDM XThR.Tn[11].t69 VGND.t1833 VGND.t1832 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2436 XA.XIR[8].XIC[4].icell.PDM XThR.Tn[7].t59 VGND.t369 VGND.t368 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2437 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR.t2052 VGND.t1670 VGND.t1669 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2438 XA.XIR[4].XIC[9].icell.Ien XThR.Tn[4].t66 VPWR.t448 VPWR.t447 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2439 XA.XIR[3].XIC[10].icell.Ien XThR.Tn[3].t68 VPWR.t412 VPWR.t411 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2440 XA.XIR[11].XIC[5].icell.PDM XThR.Tn[10].t62 VGND.t875 VGND.t874 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2441 XA.XIR[14].XIC[11].icell.SM XA.XIR[14].XIC[11].icell.Ien Iout.t218 VGND.t2187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2442 XA.XIR[15].XIC[13].icell.PDM XThR.Tn[14].t67 VGND.t89 VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2443 VPWR.t475 XThC.XTBN.Y.t102 XThC.Tn[11].t6 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2444 VPWR.t1048 XThR.Tn[2].t63 XA.XIR[3].XIC[5].icell.PUM VPWR.t1047 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2445 VPWR.t125 XThR.XTB6.Y a_n1049_5611# VPWR.t124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2446 VGND.t1672 VPWR.t2053 XA.XIR[15].XIC_dummy_left.icell.PDM VGND.t1671 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2447 a_n997_2891# XThR.XTB3.Y.t15 XThR.Tn[10].t11 VGND.t190 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2448 XA.XIR[1].XIC[11].icell.PDM XThR.Tn[1].t59 XA.XIR[1].XIC[11].icell.Ien VGND.t1293 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2449 XA.XIR[13].XIC[12].icell.SM XA.XIR[13].XIC[12].icell.Ien Iout.t69 VGND.t808 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2450 VPWR.t715 XThR.Tn[6].t65 XA.XIR[7].XIC[5].icell.PUM VPWR.t714 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2451 XA.XIR[10].XIC[1].icell.PUM XThC.Tn[1].t40 XA.XIR[10].XIC[1].icell.Ien VPWR.t1208 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2452 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR.t1456 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR.t1457 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2453 XA.XIR[1].XIC[6].icell.SM XA.XIR[1].XIC[6].icell.Ien Iout.t131 VGND.t1394 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2454 XA.XIR[2].XIC[8].icell.PDM XThR.Tn[1].t60 VGND.t1295 VGND.t1294 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2455 XA.XIR[2].XIC[14].icell.PDM XThR.Tn[1].t61 VGND.t1297 VGND.t1296 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2456 XA.XIR[13].XIC[2].icell.PUM XThC.Tn[2].t37 XA.XIR[13].XIC[2].icell.Ien VPWR.t912 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2457 XA.XIR[11].XIC[10].icell.PDM XThR.Tn[11].t70 XA.XIR[11].XIC[10].icell.Ien VGND.t1834 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2458 XA.XIR[9].XIC[12].icell.PDM XThR.Tn[8].t65 VGND.t1457 VGND.t1456 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2459 XA.XIR[8].XIC[14].icell.PUM XThC.Tn[14].t39 XA.XIR[8].XIC[14].icell.Ien VPWR.t1291 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2460 VGND.t2240 Vbias.t227 XA.XIR[10].XIC[5].icell.SM VGND.t2239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2461 XA.XIR[15].XIC[11].icell.Ien VPWR.t1453 VPWR.t1455 VPWR.t1454 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2462 VGND.t1547 XThC.Tn[4].t40 XA.XIR[10].XIC[4].icell.PDM VGND.t1546 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2463 VGND.t1674 VPWR.t2054 XA.XIR[5].XIC_dummy_right.icell.PDM VGND.t1673 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2464 XA.XIR[11].XIC_15.icell.PUM VPWR.t1451 XA.XIR[11].XIC_15.icell.Ien VPWR.t1452 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2465 XA.XIR[1].XIC[2].icell.PDM XThR.Tn[1].t62 XA.XIR[1].XIC[2].icell.Ien VGND.t1298 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2466 VGND.t2242 Vbias.t228 XA.XIR[13].XIC[6].icell.SM VGND.t2241 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2467 XA.XIR[12].XIC[7].icell.Ien XThR.Tn[12].t65 VPWR.t1317 VPWR.t1316 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2468 VGND.t2285 XThC.Tn[5].t36 XA.XIR[13].XIC[5].icell.PDM VGND.t2284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2469 VGND.t1676 VPWR.t2055 XA.XIR[9].XIC_dummy_right.icell.PDM VGND.t1675 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2470 XThC.Tn[2].t4 XThC.XTBN.Y.t103 a_4067_9615# VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2471 XA.XIR[4].XIC[3].icell.PDM XThR.Tn[4].t67 XA.XIR[4].XIC[3].icell.Ien VGND.t2243 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2472 VPWR.t797 XThR.Tn[8].t66 XA.XIR[9].XIC[11].icell.PUM VPWR.t796 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2473 VPWR.t21 XThR.Tn[14].t68 XA.XIR[15].XIC[3].icell.PUM VPWR.t20 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2474 XA.XIR[7].XIC[12].icell.PUM XThC.Tn[12].t38 XA.XIR[7].XIC[12].icell.Ien VPWR.t215 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2475 VGND.t1579 XThR.XTB7.B XThR.XTB4.Y VGND.t1578 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2476 VPWR.t1450 VPWR.t1448 XA.XIR[10].XIC_15.icell.PUM VPWR.t1449 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2477 VGND.t1406 Vbias.t229 XA.XIR[4].XIC_15.icell.SM VGND.t1405 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2478 XA.XIR[15].XIC[2].icell.Ien VPWR.t1445 VPWR.t1447 VPWR.t1446 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2479 VGND.t1408 Vbias.t230 XA.XIR[11].XIC[13].icell.SM VGND.t1407 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2480 XA.XIR[10].XIC[14].icell.Ien XThR.Tn[10].t63 VPWR.t557 VPWR.t556 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2481 VGND.t1937 XThR.XTB1.Y.t16 XThR.Tn[0].t11 VGND.t1936 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2482 VPWR.t1270 XThR.Tn[1].t63 XA.XIR[2].XIC[4].icell.PUM VPWR.t1269 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2483 VPWR.t1826 XThR.Tn[5].t64 XA.XIR[6].XIC[1].icell.PUM VPWR.t1825 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2484 XA.XIR[13].XIC_15.icell.Ien XThR.Tn[13].t64 VPWR.t982 VPWR.t981 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2485 XA.XIR[14].XIC[9].icell.SM XA.XIR[14].XIC[9].icell.Ien Iout.t45 VGND.t329 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2486 VPWR.t799 XThR.Tn[8].t67 XA.XIR[9].XIC[2].icell.PUM VPWR.t798 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2487 XA.XIR[15].XIC[5].icell.PDM VPWR.t2056 XA.XIR[15].XIC[5].icell.Ien VGND.t1677 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2488 XA.XIR[10].XIC_dummy_left.icell.SM XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout VGND.t250 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2489 VGND.t1500 XThC.Tn[11].t38 XA.XIR[14].XIC[11].icell.PDM VGND.t1499 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2490 VGND.t1410 Vbias.t231 XA.XIR[2].XIC[2].icell.SM VGND.t1409 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2491 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR.t1442 VPWR.t1444 VPWR.t1443 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2492 XA.XIR[1].XIC[10].icell.SM XA.XIR[1].XIC[10].icell.Ien Iout.t54 VGND.t582 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2493 a_8739_9569# XThC.XTBN.Y.t104 VGND.t679 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2494 XA.XIR[9].XIC[10].icell.PDM XThR.Tn[8].t68 VGND.t1459 VGND.t1458 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2495 XThC.Tn[6].t0 XThC.XTB7.Y VGND.t214 VGND.t213 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2496 XA.XIR[3].XIC[5].icell.Ien XThR.Tn[3].t69 VPWR.t414 VPWR.t413 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2497 XA.XIR[11].XIC[0].icell.PDM XThR.Tn[10].t64 VGND.t877 VGND.t876 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2498 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[5].t65 VGND.t2552 VGND.t2551 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2499 XA.XIR[1].XIC[6].icell.PDM XThR.Tn[1].t64 XA.XIR[1].XIC[6].icell.Ien VGND.t2163 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2500 VGND.t1412 Vbias.t232 XA.XIR[13].XIC[10].icell.SM VGND.t1411 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2501 VGND.t593 XThC.XTBN.Y.t105 XThC.Tn[7].t0 VGND.t592 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2502 XThC.Tn[12].t8 XThC.XTBN.Y.t106 VPWR.t401 VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2503 XA.XIR[12].XIC[11].icell.Ien XThR.Tn[12].t66 VPWR.t398 VPWR.t397 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2504 XA.XIR[4].XIC[7].icell.PDM XThR.Tn[4].t68 XA.XIR[4].XIC[7].icell.Ien VGND.t2244 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2505 VGND.t1611 XThC.Tn[2].t38 XA.XIR[14].XIC[2].icell.PDM VGND.t1610 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2506 XThC.Tn[12].t0 XThC.XTB5.Y a_9827_9569# VGND.t286 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2507 XA.XIR[1].XIC[1].icell.SM XA.XIR[1].XIC[1].icell.Ien Iout.t35 VGND.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2508 XA.XIR[2].XIC[3].icell.PDM XThR.Tn[1].t65 VGND.t2165 VGND.t2164 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2509 XA.XIR[7].XIC[10].icell.PUM XThC.Tn[10].t39 XA.XIR[7].XIC[10].icell.Ien VPWR.t394 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2510 XA.XIR[4].XIC[12].icell.PUM XThC.Tn[12].t39 XA.XIR[4].XIC[12].icell.Ien VPWR.t216 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2511 a_8963_9569# XThC.XTB4.Y.t15 XThC.Tn[11].t2 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2512 XA.XIR[0].XIC[13].icell.SM XA.XIR[0].XIC[13].icell.Ien Iout.t53 VGND.t525 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2513 XA.XIR[3].XIC[13].icell.PUM XThC.Tn[13].t39 XA.XIR[3].XIC[13].icell.Ien VPWR.t1136 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2514 VGND.t1414 Vbias.t233 XA.XIR[10].XIC[0].icell.SM VGND.t1413 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2515 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR.t1440 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR.t1441 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2516 VGND.t1416 Vbias.t234 XA.XIR[5].XIC[12].icell.SM VGND.t1415 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2517 VGND.t2038 XThC.Tn[8].t40 XA.XIR[1].XIC[8].icell.PDM VGND.t2037 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2518 VGND.t2178 XThC.Tn[14].t40 XA.XIR[1].XIC[14].icell.PDM VGND.t2177 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2519 XThR.Tn[13].t5 XThR.XTB6.Y VPWR.t123 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2520 VGND.t1418 Vbias.t235 XA.XIR[13].XIC[1].icell.SM VGND.t1417 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2521 XA.XIR[12].XIC[2].icell.Ien XThR.Tn[12].t67 VPWR.t400 VPWR.t399 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2522 VGND.t1482 XThC.Tn[0].t37 XA.XIR[13].XIC[0].icell.PDM VGND.t1481 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2523 VGND.t1420 Vbias.t236 XA.XIR[8].XIC[13].icell.SM VGND.t1419 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2524 XA.XIR[7].XIC[14].icell.Ien XThR.Tn[7].t60 VPWR.t221 VPWR.t220 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2525 VGND.t341 XThC.Tn[12].t40 XA.XIR[8].XIC[12].icell.PDM VGND.t340 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2526 VPWR.t1272 XThR.Tn[1].t66 XA.XIR[2].XIC[0].icell.PUM VPWR.t1271 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2527 VGND.t1948 XThC.Tn[13].t40 XA.XIR[11].XIC[13].icell.PDM VGND.t1947 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2528 XA.XIR[12].XIC[7].icell.PUM XThC.Tn[7].t35 XA.XIR[12].XIC[7].icell.Ien VPWR.t1139 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2529 VGND.t594 XThC.XTBN.Y.t107 a_7875_9569# VGND.t207 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2530 XA.XIR[12].XIC[5].icell.PDM XThR.Tn[12].t68 XA.XIR[12].XIC[5].icell.Ien VGND.t584 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2531 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR.t2057 XA.XIR[11].XIC_dummy_left.icell.Ien VGND.t1678 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2532 XA.XIR[15].XIC[8].icell.PUM XThC.Tn[8].t41 XA.XIR[15].XIC[8].icell.Ien VPWR.t1192 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2533 XA.XIR[2].XIC[4].icell.Ien XThR.Tn[2].t64 VPWR.t1046 VPWR.t1045 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2534 XA.XIR[14].XIC_15.icell.PDM XThR.Tn[14].t69 XA.XIR[14].XIC_15.icell.Ien VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2535 XA.XIR[11].XIC_15.icell.SM XA.XIR[11].XIC_15.icell.Ien Iout.t246 VGND.t2616 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2536 VGND.t1422 Vbias.t237 XA.XIR[7].XIC[11].icell.SM VGND.t1421 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2537 XA.XIR[6].XIC[12].icell.Ien XThR.Tn[6].t66 VPWR.t717 VPWR.t716 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2538 XA.XIR[5].XIC[13].icell.Ien XThR.Tn[5].t66 VPWR.t1828 VPWR.t1827 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2539 XA.XIR[14].XIC[4].icell.SM XA.XIR[14].XIC[4].icell.Ien Iout.t110 VGND.t1270 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2540 XA.XIR[9].XIC[13].icell.Ien XThR.Tn[9].t64 VPWR.t363 VPWR.t362 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2541 XA.XIR[6].XIC[10].icell.PDM XThR.Tn[5].t67 VGND.t2542 VGND.t2541 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2542 XA.XIR[9].XIC_dummy_right.icell.SM XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout VGND.t2521 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2543 VPWR.t576 VGND.t2701 XA.XIR[0].XIC[12].icell.PUM VPWR.t575 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2544 XA.XIR[15].XIC[0].icell.PDM VPWR.t2058 XA.XIR[15].XIC[0].icell.Ien VGND.t1679 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2545 a_8963_9569# XThC.XTBN.Y.t108 VGND.t595 VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2546 XA.XIR[10].XIC[12].icell.PDM XThR.Tn[10].t65 XA.XIR[10].XIC[12].icell.Ien VGND.t878 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2547 VGND.t491 XThC.Tn[6].t40 XA.XIR[14].XIC[6].icell.PDM VGND.t490 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2548 XA.XIR[1].XIC[9].icell.PUM XThC.Tn[9].t41 XA.XIR[1].XIC[9].icell.Ien VPWR.t1034 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2549 XA.XIR[2].XIC[7].icell.PDM XThR.Tn[1].t67 VGND.t2167 VGND.t2166 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2550 XA.XIR[13].XIC[13].icell.PDM XThR.Tn[13].t65 XA.XIR[13].XIC[13].icell.Ien VGND.t1809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2551 VPWR.t1439 VPWR.t1437 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR.t1438 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2552 XA.XIR[4].XIC[10].icell.PUM XThC.Tn[10].t40 XA.XIR[4].XIC[10].icell.Ien VPWR.t395 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2553 XA.XIR[14].XIC[11].icell.PDM XThR.Tn[13].t66 VGND.t108 VGND.t107 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2554 XA.XIR[0].XIC[8].icell.PDM XThR.Tn[0].t66 XA.XIR[0].XIC[8].icell.Ien VGND.t1114 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2555 XA.XIR[0].XIC[14].icell.PDM XThR.Tn[0].t67 XA.XIR[0].XIC[14].icell.Ien VGND.t1115 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2556 VPWR.t223 XThR.Tn[7].t61 XA.XIR[8].XIC[7].icell.PUM VPWR.t222 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2557 VGND.t579 XThC.Tn[10].t41 XA.XIR[8].XIC[10].icell.PDM VGND.t578 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2558 XThC.Tn[11].t5 XThC.XTBN.Y.t109 VPWR.t402 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2559 VPWR.t559 XThR.Tn[10].t66 XA.XIR[11].XIC[8].icell.PUM VPWR.t558 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2560 VGND.t1424 Vbias.t238 XA.XIR[1].XIC[7].icell.SM VGND.t1423 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2561 XThR.Tn[6].t1 XThR.XTBN.Y.t108 a_n1049_5317# VPWR.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2562 XA.XIR[7].XIC[5].icell.PUM XThC.Tn[5].t37 XA.XIR[7].XIC[5].icell.Ien VPWR.t1351 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2563 VPWR.t659 XThC.XTB4.Y.t16 XThC.Tn[11].t3 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2564 XThR.XTB7.Y XThR.XTB7.B a_n1319_5317# VPWR.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2565 XA.XIR[12].XIC[11].icell.PUM XThC.Tn[11].t39 XA.XIR[12].XIC[11].icell.Ien VPWR.t817 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2566 VGND.t1426 Vbias.t239 XA.XIR[4].XIC[8].icell.SM VGND.t1425 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2567 XA.XIR[15].XIC[1].icell.PDM XThR.Tn[14].t70 VGND.t92 VGND.t91 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2568 XA.XIR[14].XIC[2].icell.PDM XThR.Tn[13].t67 VGND.t110 VGND.t109 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2569 XA.XIR[10].XIC[5].icell.PDM XThR.Tn[9].t65 VGND.t535 VGND.t534 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2570 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR.t2059 VGND.t1681 VGND.t1680 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2571 VGND.t2218 XThC.Tn[3].t41 XA.XIR[1].XIC[3].icell.PDM VGND.t2217 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2572 VGND.t1428 Vbias.t240 XA.XIR[7].XIC[9].icell.SM VGND.t1427 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2573 XA.XIR[6].XIC[10].icell.Ien XThR.Tn[6].t67 VPWR.t719 VPWR.t718 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2574 XA.XIR[2].XIC[0].icell.Ien XThR.Tn[2].t65 VPWR.t1044 VPWR.t1043 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2575 XA.XIR[12].XIC_15.icell.PDM VPWR.t2060 VGND.t1683 VGND.t1682 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2576 XA.XIR[12].XIC[12].icell.SM XA.XIR[12].XIC[12].icell.Ien Iout.t217 VGND.t2154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2577 XA.XIR[8].XIC_15.icell.SM XA.XIR[8].XIC_15.icell.Ien Iout.t194 VGND.t1802 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2578 XA.XIR[15].XIC[13].icell.SM XA.XIR[15].XIC[13].icell.Ien Iout.t203 VGND.t1951 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2579 VPWR.t574 VGND.t2702 XA.XIR[0].XIC[10].icell.PUM VPWR.t573 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2580 VPWR.t35 XThC.XTB3.Y.t14 a_4067_9615# VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2581 XA.XIR[3].XIC[6].icell.PUM XThC.Tn[6].t41 XA.XIR[3].XIC[6].icell.Ien VPWR.t439 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2582 XA.XIR[12].XIC[0].icell.PDM XThR.Tn[12].t69 XA.XIR[12].XIC[0].icell.Ien VGND.t585 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2583 XA.XIR[12].XIC[2].icell.PUM XThC.Tn[2].t39 XA.XIR[12].XIC[2].icell.Ien VPWR.t913 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2584 XA.XIR[10].XIC[10].icell.PDM XThR.Tn[10].t67 XA.XIR[10].XIC[10].icell.Ien VGND.t2042 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2585 VGND.t457 XThR.XTBN.Y.t109 a_n997_1803# VGND.t424 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2586 XA.XIR[7].XIC[12].icell.PDM XThR.Tn[7].t62 XA.XIR[7].XIC[12].icell.Ien VGND.t370 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2587 XA.XIR[0].XIC[9].icell.Ien XThR.Tn[0].t68 VPWR.t647 VPWR.t646 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2588 XA.XIR[15].XIC[3].icell.PUM XThC.Tn[3].t42 XA.XIR[15].XIC[3].icell.Ien VPWR.t1322 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2589 XA.XIR[6].XIC[7].icell.PUM XThC.Tn[7].t36 XA.XIR[6].XIC[7].icell.Ien VPWR.t1140 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2590 XA.XIR[10].XIC_15.icell.PUM VPWR.t1435 XA.XIR[10].XIC_15.icell.Ien VPWR.t1436 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2591 a_3773_9615# XThC.XTB2.Y VPWR.t101 VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2592 VPWR.t1434 VPWR.t1432 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR.t1433 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2593 VGND.t2335 Vbias.t241 XA.XIR[12].XIC[6].icell.SM VGND.t2334 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2594 VGND.t1871 XThC.Tn[9].t42 XA.XIR[3].XIC[9].icell.PDM VGND.t1870 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2595 VGND.t2287 XThC.Tn[5].t38 XA.XIR[12].XIC[5].icell.PDM VGND.t2286 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2596 VPWR.t225 XThR.Tn[7].t63 XA.XIR[8].XIC[11].icell.PUM VPWR.t224 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2597 XA.XIR[2].XIC[4].icell.PUM XThC.Tn[4].t41 XA.XIR[2].XIC[4].icell.Ien VPWR.t852 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2598 VPWR.t77 XThR.XTB4.Y XThR.Tn[11].t4 VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2599 a_n997_715# XThR.XTBN.Y.t110 VGND.t459 VGND.t458 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2600 VGND.t2337 Vbias.t242 XA.XIR[6].XIC[5].icell.SM VGND.t2336 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2601 VPWR.t1131 XThR.XTB1.Y.t17 a_n1049_8581# VPWR.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2602 XA.XIR[4].XIC[5].icell.PUM XThC.Tn[5].t39 XA.XIR[4].XIC[5].icell.Ien VPWR.t1352 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2603 XA.XIR[5].XIC[6].icell.Ien XThR.Tn[5].t68 VPWR.t1800 VPWR.t1799 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2604 XThR.Tn[14].t9 XThR.XTB7.Y VPWR.t942 VPWR.t122 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2605 XA.XIR[14].XIC[6].icell.PDM XThR.Tn[13].t68 VGND.t112 VGND.t111 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2606 XA.XIR[9].XIC[6].icell.Ien XThR.Tn[9].t66 VPWR.t365 VPWR.t364 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2607 VGND.t2339 Vbias.t243 XA.XIR[9].XIC[6].icell.SM VGND.t2338 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2608 VGND.t596 XThC.XTBN.Y.t110 XThC.Tn[3].t1 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2609 XA.XIR[8].XIC[7].icell.Ien XThR.Tn[8].t69 VPWR.t801 VPWR.t800 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2610 VGND.t1962 XThC.Tn[7].t37 XA.XIR[1].XIC[7].icell.PDM VGND.t1961 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2611 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR.t2061 VGND.t1685 VGND.t1684 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2612 XA.XIR[0].XIC[3].icell.PDM XThR.Tn[0].t69 XA.XIR[0].XIC[3].icell.Ien VGND.t1116 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2613 XA.XIR[9].XIC_dummy_left.icell.SM XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout VGND.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2614 VPWR.t1926 XThR.Tn[7].t64 XA.XIR[8].XIC[2].icell.PUM VPWR.t1925 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2615 XThC.Tn[1].t0 XThC.XTB2.Y VGND.t205 VGND.t204 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2616 VPWR.t1042 XThR.Tn[2].t66 XA.XIR[3].XIC[14].icell.PUM VPWR.t1041 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2617 XA.XIR[5].XIC[9].icell.PDM XThR.Tn[5].t69 XA.XIR[5].XIC[9].icell.Ien VGND.t2543 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2618 XA.XIR[11].XIC[8].icell.Ien XThR.Tn[11].t71 VPWR.t1018 VPWR.t1017 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2619 VPWR.t469 XThC.XTBN.A XThC.XTBN.Y.t2 VPWR.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2620 VPWR.t1202 XThR.Tn[10].t68 XA.XIR[11].XIC[3].icell.PUM VPWR.t1201 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2621 XA.XIR[9].XIC[9].icell.PDM XThR.Tn[9].t67 XA.XIR[9].XIC[9].icell.Ien VGND.t536 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2622 VPWR.t721 XThR.Tn[6].t68 XA.XIR[7].XIC[14].icell.PUM VPWR.t720 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2623 VGND.t2341 Vbias.t244 XA.XIR[1].XIC[2].icell.SM VGND.t2340 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2624 VPWR.t1431 VPWR.t1429 XA.XIR[6].XIC_15.icell.PUM VPWR.t1430 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2625 VGND.t2343 Vbias.t245 XA.XIR[4].XIC[3].icell.SM VGND.t2342 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2626 XA.XIR[7].XIC[10].icell.PDM XThR.Tn[7].t65 XA.XIR[7].XIC[10].icell.Ien VGND.t2684 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2627 XThR.Tn[2].t11 XThR.XTB3.Y.t16 VGND.t2683 VGND.t188 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2628 XA.XIR[10].XIC[0].icell.PDM XThR.Tn[9].t68 VGND.t538 VGND.t537 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2629 XA.XIR[6].XIC[11].icell.PUM XThC.Tn[11].t40 XA.XIR[6].XIC[11].icell.Ien VPWR.t818 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2630 XA.XIR[11].XIC[8].icell.SM XA.XIR[11].XIC[8].icell.Ien Iout.t136 VGND.t1404 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2631 VGND.t2345 Vbias.t246 XA.XIR[7].XIC[4].icell.SM VGND.t2344 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2632 XA.XIR[6].XIC[5].icell.Ien XThR.Tn[6].t69 VPWR.t723 VPWR.t722 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2633 VGND.t904 VGND.t902 XA.XIR[2].XIC_dummy_right.icell.SM VGND.t903 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2634 VGND.t2347 Vbias.t247 XA.XIR[12].XIC[10].icell.SM VGND.t2346 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2635 XA.XIR[8].XIC[13].icell.PDM XThR.Tn[7].t66 VGND.t2686 VGND.t2685 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2636 a_n997_3979# XThR.XTB1.Y.t18 XThR.Tn[8].t11 VGND.t1938 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2637 XA.XIR[7].XIC[11].icell.SM XA.XIR[7].XIC[11].icell.Ien Iout.t193 VGND.t1801 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2638 a_3299_10575# XThC.XTB7.B VGND.t1328 VGND.t413 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2639 VGND.t1687 VPWR.t2062 XA.XIR[8].XIC_dummy_left.icell.PDM VGND.t1686 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2640 VGND.t461 XThR.XTBN.Y.t111 XThR.Tn[6].t4 VGND.t460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2641 VPWR.t572 VGND.t2703 XA.XIR[0].XIC[5].icell.PUM VPWR.t571 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2642 XA.XIR[3].XIC[1].icell.PUM XThC.Tn[1].t41 XA.XIR[3].XIC[1].icell.Ien VPWR.t1209 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2643 XA.XIR[2].XIC[0].icell.PUM XThC.Tn[0].t38 XA.XIR[2].XIC[0].icell.Ien VPWR.t811 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2644 VPWR.t1020 XThR.Tn[11].t72 XA.XIR[12].XIC[9].icell.PUM VPWR.t1019 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2645 XA.XIR[6].XIC[2].icell.PUM XThC.Tn[2].t40 XA.XIR[6].XIC[2].icell.Ien VPWR.t914 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2646 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR.t1426 VPWR.t1428 VPWR.t1427 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2647 VGND.t2349 Vbias.t248 XA.XIR[12].XIC[1].icell.SM VGND.t2348 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2648 VGND.t2351 Vbias.t249 XA.XIR[3].XIC[5].icell.SM VGND.t2350 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2649 VGND.t1484 XThC.Tn[0].t39 XA.XIR[12].XIC[0].icell.PDM VGND.t1483 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2650 VPWR.t570 VGND.t2704 Vbias.t1 VPWR.t568 sky130_fd_pr__pfet_01v8 ad=0.2465 pd=2.28 as=0.12325 ps=1.14 w=0.85 l=2
X2651 VGND.t1549 XThC.Tn[4].t42 XA.XIR[3].XIC[4].icell.PDM VGND.t1548 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2652 VGND.t2353 Vbias.t250 XA.XIR[9].XIC[10].icell.SM VGND.t2352 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2653 XA.XIR[8].XIC[11].icell.Ien XThR.Tn[8].t70 VPWR.t803 VPWR.t802 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2654 VGND.t2074 XThC.Tn[1].t42 XA.XIR[11].XIC[1].icell.PDM VGND.t2073 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2655 VGND.t2355 Vbias.t251 XA.XIR[10].XIC[14].icell.SM VGND.t2354 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2656 XA.XIR[0].XIC[7].icell.PDM XThR.Tn[0].t70 XA.XIR[0].XIC[7].icell.Ien VGND.t1117 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2657 VGND.t2289 XThC.Tn[5].t40 XA.XIR[6].XIC[5].icell.PDM VGND.t2288 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2658 VPWR.t403 XThC.XTBN.Y.t111 XThC.Tn[10].t9 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2659 VGND.t1950 XThC.Tn[13].t41 XA.XIR[10].XIC[13].icell.PDM VGND.t1949 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2660 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR.t2063 XA.XIR[10].XIC_dummy_left.icell.Ien VGND.t1688 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2661 XA.XIR[0].XIC[12].icell.PUM XThC.Tn[12].t41 XA.XIR[0].XIC[12].icell.Ien VPWR.t217 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2662 VGND.t597 XThC.XTBN.Y.t112 a_8963_9569# VGND.t328 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2663 XA.XIR[5].XIC[1].icell.Ien XThR.Tn[5].t70 VPWR.t1802 VPWR.t1801 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2664 VGND.t2357 Vbias.t252 XA.XIR[6].XIC[0].icell.SM VGND.t2356 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2665 XA.XIR[7].XIC[9].icell.PDM XThR.Tn[6].t70 VGND.t1317 VGND.t1316 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2666 VPWR.t759 XThC.XTB5.A a_5155_10571# VPWR.t158 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2667 VPWR.t111 XThC.XTB7.Y XThC.Tn[14].t4 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2668 XThR.Tn[1].t4 XThR.XTBN.Y.t112 VGND.t463 VGND.t462 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2669 XA.XIR[1].XIC[4].icell.Ien XThR.Tn[1].t68 VPWR.t1274 VPWR.t1273 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2670 XA.XIR[9].XIC[1].icell.Ien XThR.Tn[9].t69 VPWR.t367 VPWR.t366 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2671 VGND.t2050 Vbias.t253 XA.XIR[9].XIC[1].icell.SM VGND.t2049 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2672 XA.XIR[8].XIC[2].icell.Ien XThR.Tn[8].t71 VPWR.t157 VPWR.t156 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2673 XA.XIR[3].XIC[14].icell.Ien XThR.Tn[3].t70 VPWR.t416 VPWR.t415 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2674 XA.XIR[5].XIC[7].icell.SM XA.XIR[5].XIC[7].icell.Ien Iout.t98 VGND.t1138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2675 VPWR.t1405 XThC.XTB7.A XThC.XTB3.Y.t2 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2676 XA.XIR[11].XIC[3].icell.Ien XThR.Tn[11].t73 VPWR.t1022 VPWR.t1021 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2677 XA.XIR[5].XIC[4].icell.PDM XThR.Tn[5].t71 XA.XIR[5].XIC[4].icell.Ien VGND.t2544 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2678 XA.XIR[8].XIC[8].icell.SM XA.XIR[8].XIC[8].icell.Ien Iout.t184 VGND.t1772 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2679 XA.XIR[7].XIC[9].icell.SM XA.XIR[7].XIC[9].icell.Ien Iout.t58 VGND.t644 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2680 XA.XIR[13].XIC[1].icell.PDM XThR.Tn[13].t69 XA.XIR[13].XIC[1].icell.Ien VGND.t113 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2681 XA.XIR[9].XIC[4].icell.PDM XThR.Tn[9].t70 XA.XIR[9].XIC[4].icell.Ien VGND.t539 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2682 XThR.Tn[8].t4 XThR.XTBN.Y.t113 VPWR.t284 VPWR.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2683 VPWR.t1276 XThR.Tn[1].t69 XA.XIR[2].XIC[13].icell.PUM VPWR.t1275 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2684 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR.t2064 XA.XIR[4].XIC_dummy_right.icell.Ien VGND.t1689 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2685 XThR.Tn[5].t4 XThR.XTBN.Y.t114 a_n1049_5611# VPWR.t282 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2686 a_n997_2891# XThR.XTB3.Y.t17 XThR.Tn[10].t0 VGND.t187 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2687 XA.XIR[8].XIC[5].icell.PDM XThR.Tn[8].t72 XA.XIR[8].XIC[5].icell.Ien VGND.t284 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2688 XThR.XTB6.Y XThR.XTB7.B a_n1319_5611# VPWR.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2689 VPWR.t1425 VPWR.t1423 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1424 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2690 XA.XIR[2].XIC[7].icell.SM XA.XIR[2].XIC[7].icell.Ien Iout.t21 VGND.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2691 XA.XIR[11].XIC[3].icell.SM XA.XIR[11].XIC[3].icell.Ien Iout.t111 VGND.t1277 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2692 a_n1049_7787# XThR.XTBN.Y.t115 XThR.Tn[1].t0 VPWR.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X2693 a_3773_9615# XThC.XTBN.Y.t113 XThC.Tn[1].t9 VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2694 VPWR.t875 XThR.XTB7.B XThR.XTB3.Y.t0 VPWR.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2695 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR.t2065 XA.XIR[7].XIC_dummy_left.icell.Ien VGND.t1690 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2696 XA.XIR[0].XIC[10].icell.PUM XThC.Tn[10].t42 XA.XIR[0].XIC[10].icell.Ien VPWR.t396 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2697 a_4067_9615# XThC.XTB3.Y.t15 VPWR.t36 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2698 VGND.t2052 Vbias.t254 XA.XIR[3].XIC[0].icell.SM VGND.t2051 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2699 VPWR.t37 XThC.XTB3.Y.t16 XThC.Tn[10].t6 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2700 VPWR.t404 XThC.XTBN.Y.t114 XThC.Tn[14].t9 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2701 XA.XIR[1].XIC[0].icell.Ien XThR.Tn[1].t70 VPWR.t1113 VPWR.t1112 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2702 VGND.t901 VGND.t899 XA.XIR[2].XIC_dummy_left.icell.SM VGND.t900 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2703 XA.XIR[14].XIC[4].icell.PUM XThC.Tn[4].t43 XA.XIR[14].XIC[4].icell.Ien VPWR.t853 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2704 XA.XIR[15].XIC_15.icell.PDM VPWR.t2066 VGND.t1692 VGND.t1691 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2705 XA.XIR[10].XIC[5].icell.SM XA.XIR[10].XIC[5].icell.Ien Iout.t182 VGND.t1770 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2706 VGND.t1486 XThC.Tn[0].t40 XA.XIR[6].XIC[0].icell.PDM VGND.t1485 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2707 XA.XIR[14].XIC[13].icell.SM XA.XIR[14].XIC[13].icell.Ien Iout.t222 VGND.t2294 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2708 VGND.t2584 XThR.XTBN.Y.t116 XThR.Tn[0].t5 VGND.t315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2709 XA.XIR[13].XIC[6].icell.SM XA.XIR[13].XIC[6].icell.Ien Iout.t15 VGND.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2710 VGND.t105 XThC.XTB3.Y.t17 XThC.Tn[2].t3 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.08775 ps=0.92 w=0.65 l=0.15
X2711 XA.XIR[5].XIC[7].icell.PUM XThC.Tn[7].t38 XA.XIR[5].XIC[7].icell.Ien VPWR.t1141 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2712 XThR.Tn[10].t2 XThR.XTBN.Y.t117 VPWR.t1856 VPWR.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2713 XA.XIR[7].XIC[4].icell.PDM XThR.Tn[6].t71 VGND.t1319 VGND.t1318 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2714 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR.t2067 VGND.t1694 VGND.t1693 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2715 XA.XIR[9].XIC[7].icell.PUM XThC.Tn[7].t39 XA.XIR[9].XIC[7].icell.Ien VPWR.t1142 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2716 XA.XIR[5].XIC[2].icell.SM XA.XIR[5].XIC[2].icell.Ien Iout.t191 VGND.t1799 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2717 XA.XIR[8].XIC[8].icell.PUM XThC.Tn[8].t42 XA.XIR[8].XIC[8].icell.Ien VPWR.t547 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2718 VGND.t2054 Vbias.t255 XA.XIR[0].XIC[11].icell.SM VGND.t2053 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2719 VPWR.t763 XThC.XTB6.Y a_5949_9615# VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2720 XThR.Tn[1].t8 XThR.XTB2.Y VGND.t1977 VGND.t1558 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X2721 XA.XIR[4].XIC_15.icell.SM XA.XIR[4].XIC_15.icell.Ien Iout.t141 VGND.t1450 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2722 VGND.t2585 XThR.XTBN.Y.t118 a_n997_3755# VGND.t1256 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2723 VPWR.t707 data[3].t1 XThC.XTBN.A VPWR.t160 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2724 XA.XIR[8].XIC[3].icell.SM XA.XIR[8].XIC[3].icell.Ien Iout.t192 VGND.t1800 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2725 a_2979_9615# XThC.XTB1.Y.t17 VPWR.t627 VPWR.t626 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.135 ps=1.27 w=1 l=0.15
X2726 XThC.Tn[3].t0 XThC.XTBN.Y.t115 VGND.t598 VGND.t326 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2727 XA.XIR[2].XIC[13].icell.Ien XThR.Tn[2].t67 VPWR.t1040 VPWR.t1039 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2728 XA.XIR[7].XIC[4].icell.SM XA.XIR[7].XIC[4].icell.Ien Iout.t105 VGND.t1153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2729 XA.XIR[8].XIC[0].icell.PDM XThR.Tn[8].t73 XA.XIR[8].XIC[0].icell.Ien VGND.t285 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2730 XA.XIR[3].XIC[12].icell.PDM XThR.Tn[3].t71 XA.XIR[3].XIC[12].icell.Ien VGND.t602 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2731 XA.XIR[7].XIC[14].icell.PUM XThC.Tn[14].t41 XA.XIR[7].XIC[14].icell.Ien VPWR.t491 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2732 VPWR.t39 XThR.Tn[13].t70 XA.XIR[14].XIC[12].icell.PUM VPWR.t38 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2733 XA.XIR[2].XIC[2].icell.SM XA.XIR[2].XIC[2].icell.Ien Iout.t231 VGND.t2508 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2734 XA.XIR[10].XIC[8].icell.Ien XThR.Tn[10].t69 VPWR.t1204 VPWR.t1203 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2735 a_5949_10571# XThC.XTB7.B XThC.XTB6.Y VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2736 VPWR.t1115 XThR.Tn[1].t71 XA.XIR[2].XIC[6].icell.PUM VPWR.t1114 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2737 VPWR.t71 XThR.Tn[0].t71 XA.XIR[1].XIC[7].icell.PUM VPWR.t70 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2738 XA.XIR[11].XIC[11].icell.PDM XThR.Tn[10].t70 VGND.t2044 VGND.t2043 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2739 XA.XIR[14].XIC[0].icell.PUM XThC.Tn[0].t41 XA.XIR[14].XIC[0].icell.Ien VPWR.t812 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2740 XThR.Tn[13].t4 XThR.XTB6.Y VPWR.t121 VPWR.t120 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2741 VPWR.t1324 XThR.Tn[4].t69 XA.XIR[5].XIC[7].icell.PUM VPWR.t1323 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2742 XA.XIR[13].XIC[10].icell.SM XA.XIR[13].XIC[10].icell.Ien Iout.t173 VGND.t1632 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2743 a_n1049_7493# XThR.XTB3.Y.t18 VPWR.t137 VPWR.t136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2744 XA.XIR[0].XIC[5].icell.PUM XThC.Tn[5].t41 XA.XIR[0].XIC[5].icell.Ien VPWR.t1353 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2745 XA.XIR[5].XIC[11].icell.PUM XThC.Tn[11].t41 XA.XIR[5].XIC[11].icell.Ien VPWR.t819 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2746 XA.XIR[9].XIC[11].icell.PUM XThC.Tn[11].t42 XA.XIR[9].XIC[11].icell.Ien VPWR.t820 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2747 XA.XIR[8].XIC[1].icell.PDM XThR.Tn[7].t67 VGND.t2688 VGND.t2687 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2748 VGND.t898 VGND.t896 XA.XIR[1].XIC_dummy_right.icell.SM VGND.t897 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2749 XA.XIR[3].XIC[5].icell.PDM XThR.Tn[2].t68 VGND.t127 VGND.t126 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2750 VGND.t2056 Vbias.t256 XA.XIR[0].XIC[9].icell.SM VGND.t2055 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2751 XA.XIR[11].XIC[2].icell.PDM XThR.Tn[10].t71 VGND.t2046 VGND.t2045 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2752 XA.XIR[10].XIC[0].icell.SM XA.XIR[10].XIC[0].icell.Ien Iout.t122 VGND.t1322 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2753 VPWR.t450 XThC.XTB1.Y.t18 XThC.Tn[8].t4 VPWR.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2754 VGND.t296 XThC.Tn[11].t43 XA.XIR[13].XIC[11].icell.PDM VGND.t295 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2755 XA.XIR[13].XIC[1].icell.SM XA.XIR[13].XIC[1].icell.Ien Iout.t148 VGND.t1518 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2756 VGND.t2650 XThR.XTB5.Y XThR.Tn[4].t8 VGND.t254 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2757 XThC.Tn[10].t8 XThC.XTBN.Y.t116 VPWR.t260 VPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2758 VGND.t407 XThC.XTBN.Y.t117 XThC.Tn[6].t8 VGND.t406 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2759 XA.XIR[3].XIC[10].icell.PDM XThR.Tn[3].t72 XA.XIR[3].XIC[10].icell.Ien VGND.t603 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2760 XA.XIR[5].XIC[2].icell.PUM XThC.Tn[2].t41 XA.XIR[5].XIC[2].icell.Ien VPWR.t915 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2761 VPWR.t23 XThR.Tn[14].t71 XA.XIR[15].XIC[9].icell.PUM VPWR.t22 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2762 VPWR.t41 XThR.Tn[13].t71 XA.XIR[14].XIC[10].icell.PUM VPWR.t40 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2763 XA.XIR[9].XIC[2].icell.PUM XThC.Tn[2].t42 XA.XIR[9].XIC[2].icell.Ien VPWR.t916 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2764 XA.XIR[4].XIC[14].icell.PUM XThC.Tn[14].t42 XA.XIR[4].XIC[14].icell.Ien VPWR.t492 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2765 XA.XIR[8].XIC[3].icell.PUM XThC.Tn[3].t43 XA.XIR[8].XIC[3].icell.Ien VPWR.t650 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2766 XA.XIR[3].XIC_15.icell.PUM VPWR.t1421 XA.XIR[3].XIC_15.icell.Ien VPWR.t1422 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2767 XA.XIR[5].XIC[12].icell.PDM XThR.Tn[4].t70 VGND.t2246 VGND.t2245 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2768 VGND.t2058 Vbias.t257 XA.XIR[5].XIC[6].icell.SM VGND.t2057 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2769 VGND.t2076 XThC.Tn[1].t43 XA.XIR[10].XIC[1].icell.PDM VGND.t2075 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2770 VGND.t1696 VPWR.t2068 XA.XIR[1].XIC_dummy_right.icell.PDM VGND.t1695 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2771 VGND.t2291 XThC.Tn[5].t42 XA.XIR[5].XIC[5].icell.PDM VGND.t2290 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2772 VGND.t1865 XThC.Tn[2].t43 XA.XIR[13].XIC[2].icell.PDM VGND.t1864 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2773 VGND.t2293 XThC.Tn[5].t43 XA.XIR[9].XIC[5].icell.PDM VGND.t2292 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2774 VPWR.t73 XThR.Tn[0].t72 XA.XIR[1].XIC[11].icell.PUM VPWR.t72 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2775 XA.XIR[7].XIC[8].icell.Ien XThR.Tn[7].t68 VPWR.t1928 VPWR.t1927 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2776 VPWR.t660 XThC.XTB4.Y.t17 a_4861_9615# VPWR.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2777 VPWR.t1326 XThR.Tn[4].t71 XA.XIR[5].XIC[11].icell.PUM VPWR.t1325 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2778 XA.XIR[14].XIC[12].icell.Ien XThR.Tn[14].t72 VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2779 XA.XIR[15].XIC[11].icell.PDM VPWR.t2069 XA.XIR[15].XIC[11].icell.Ien VGND.t1697 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2780 VGND.t1699 VPWR.t2070 XA.XIR[11].XIC_15.icell.PDM VGND.t1698 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2781 XA.XIR[2].XIC[13].icell.PUM XThC.Tn[13].t42 XA.XIR[2].XIC[13].icell.Ien VPWR.t1137 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2782 VGND.t2060 Vbias.t258 XA.XIR[4].XIC[12].icell.SM VGND.t2059 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2783 XThR.Tn[6].t0 XThR.XTBN.Y.t119 a_n1049_5317# VPWR.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2784 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR.t1419 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR.t1420 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2785 a_10915_9569# XThC.XTB7.Y XThC.Tn[14].t0 VGND.t212 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2786 XA.XIR[2].XIC[6].icell.Ien XThR.Tn[2].t69 VPWR.t1038 VPWR.t1037 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2787 XA.XIR[10].XIC[3].icell.Ien XThR.Tn[10].t72 VPWR.t1206 VPWR.t1205 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2788 VGND.t2062 Vbias.t259 XA.XIR[7].XIC[13].icell.SM VGND.t2061 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2789 XA.XIR[6].XIC[14].icell.Ien XThR.Tn[6].t72 VPWR.t725 VPWR.t724 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2790 VGND.t409 XThC.XTBN.Y.t118 a_10915_9569# VGND.t408 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2791 VPWR.t1117 XThR.Tn[1].t72 XA.XIR[2].XIC[1].icell.PUM VPWR.t1116 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2792 XA.XIR[5].XIC_15.icell.Ien XThR.Tn[5].t72 VPWR.t1804 VPWR.t1803 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2793 XA.XIR[11].XIC[6].icell.PDM XThR.Tn[10].t73 VGND.t2048 VGND.t2047 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2794 VGND.t1551 XThC.Tn[12].t42 XA.XIR[7].XIC[12].icell.PDM VGND.t1550 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2795 VGND.t2064 Vbias.t260 XA.XIR[6].XIC[14].icell.SM VGND.t2063 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2796 VPWR.t75 XThR.Tn[0].t73 XA.XIR[1].XIC[2].icell.PUM VPWR.t74 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2797 XA.XIR[9].XIC_15.icell.Ien XThR.Tn[9].t71 VPWR.t369 VPWR.t368 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2798 VPWR.t1328 XThR.Tn[4].t72 XA.XIR[5].XIC[2].icell.PUM VPWR.t1327 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2799 VPWR.t567 VGND.t2705 XA.XIR[0].XIC[14].icell.PUM VPWR.t566 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2800 XA.XIR[15].XIC[2].icell.PDM VPWR.t2071 XA.XIR[15].XIC[2].icell.Ien VGND.t1700 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2801 XA.XIR[2].XIC[9].icell.PDM XThR.Tn[2].t70 XA.XIR[2].XIC[9].icell.Ien VGND.t131 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2802 XThC.Tn[1].t8 XThC.XTBN.Y.t119 a_3773_9615# VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2803 XA.XIR[1].XIC[7].icell.SM XA.XIR[1].XIC[7].icell.Ien Iout.t73 VGND.t864 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2804 XA.XIR[13].XIC_15.icell.PDM XThR.Tn[13].t72 XA.XIR[13].XIC_15.icell.Ien VGND.t847 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2805 XA.XIR[3].XIC[0].icell.PDM XThR.Tn[2].t71 VGND.t130 VGND.t129 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2806 XA.XIR[5].XIC[10].icell.PDM XThR.Tn[4].t73 VGND.t2248 VGND.t2247 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2807 VGND.t2066 Vbias.t261 XA.XIR[0].XIC[4].icell.SM VGND.t2065 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2808 XA.XIR[4].XIC[8].icell.SM XA.XIR[4].XIC[8].icell.Ien Iout.t66 VGND.t805 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2809 XThC.Tn[14].t8 XThC.XTBN.Y.t120 VPWR.t261 VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2810 VGND.t2068 Vbias.t262 XA.XIR[5].XIC[10].icell.SM VGND.t2067 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2811 VGND.t2070 Vbias.t263 XA.XIR[13].XIC[7].icell.SM VGND.t2069 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2812 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR.t2072 XA.XIR[0].XIC_dummy_right.icell.Ien VGND.t1701 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2813 VGND.t638 XThC.Tn[6].t42 XA.XIR[13].XIC[6].icell.PDM VGND.t637 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2814 VGND.t2587 XThR.XTBN.Y.t120 a_n997_715# VGND.t2586 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2815 VPWR.t1418 VPWR.t1416 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR.t1417 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2816 XA.XIR[14].XIC[10].icell.Ien XThR.Tn[14].t73 VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2817 VPWR.t531 XThR.Tn[13].t73 XA.XIR[14].XIC[5].icell.PUM VPWR.t530 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2818 VPWR.t941 XThR.XTB7.Y XThR.Tn[14].t8 VPWR.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2819 XA.XIR[12].XIC[11].icell.PDM XThR.Tn[12].t70 XA.XIR[12].XIC[11].icell.Ien VGND.t586 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2820 VGND.t895 VGND.t893 XA.XIR[1].XIC_dummy_left.icell.SM VGND.t894 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2821 VGND.t2072 Vbias.t264 XA.XIR[5].XIC[1].icell.SM VGND.t2071 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2822 XA.XIR[9].XIC[5].icell.SM XA.XIR[9].XIC[5].icell.Ien Iout.t140 VGND.t1438 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2823 XThR.XTB6.A data[5].t5 VGND.t1530 VGND.t1529 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2824 XThR.Tn[0].t1 XThR.XTBN.Y.t121 a_n1049_8581# VPWR.t1857 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2825 VGND.t1488 XThC.Tn[0].t42 XA.XIR[5].XIC[0].icell.PDM VGND.t1487 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2826 XA.XIR[13].XIC[14].icell.PDM XThR.Tn[12].t71 VGND.t588 VGND.t587 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2827 a_5949_9615# XThC.XTB6.Y VPWR.t762 VPWR.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2828 XA.XIR[13].XIC[8].icell.PDM XThR.Tn[12].t72 VGND.t590 VGND.t589 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2829 XA.XIR[12].XIC[6].icell.SM XA.XIR[12].XIC[6].icell.Ien Iout.t197 VGND.t1874 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2830 VGND.t1490 XThC.Tn[0].t43 XA.XIR[9].XIC[0].icell.PDM VGND.t1489 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2831 VGND.t581 XThC.Tn[10].t43 XA.XIR[7].XIC[10].icell.PDM VGND.t580 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2832 XA.XIR[7].XIC[3].icell.Ien XThR.Tn[7].t69 VPWR.t1930 VPWR.t1929 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2833 VGND.t411 XThC.XTBN.Y.t121 a_10051_9569# VGND.t410 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2834 VGND.t1982 Vbias.t265 XA.XIR[3].XIC[14].icell.SM VGND.t1981 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2835 VGND.t1553 XThC.Tn[12].t43 XA.XIR[4].XIC[12].icell.PDM VGND.t1552 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2836 VGND.t1383 XThC.Tn[13].t43 XA.XIR[3].XIC[13].icell.PDM VGND.t1382 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2837 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR.t2073 XA.XIR[3].XIC_dummy_left.icell.Ien VGND.t1702 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2838 XA.XIR[15].XIC[6].icell.PDM VPWR.t2074 XA.XIR[15].XIC[6].icell.Ien VGND.t1703 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2839 XA.XIR[12].XIC[2].icell.PDM XThR.Tn[12].t73 XA.XIR[12].XIC[2].icell.Ien VGND.t591 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2840 XA.XIR[0].XIC[9].icell.PDM VGND.t890 VGND.t892 VGND.t891 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2841 VPWR.t262 XThC.XTBN.Y.t122 XThC.Tn[11].t4 VPWR.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2842 VGND.t412 XThC.XTBN.Y.t123 a_7651_9569# VGND.t325 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2843 XA.XIR[2].XIC[1].icell.Ien XThR.Tn[2].t72 VPWR.t1036 VPWR.t1035 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2844 XA.XIR[11].XIC[12].icell.SM XA.XIR[11].XIC[12].icell.Ien Iout.t171 VGND.t1620 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2845 XA.XIR[1].XIC[13].icell.Ien XThR.Tn[1].t73 VPWR.t1119 VPWR.t1118 sky130_fd_pr__pfet_01v8 ad=0.0725 pd=0.79 as=0.15 ps=1.6 w=0.5 l=0.15
X2846 XThR.Tn[2].t10 XThR.XTBN.Y.t122 VGND.t2588 VGND.t321 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2847 VPWR.t940 XThR.XTB7.Y a_n1049_5317# VPWR.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X2848 XA.XIR[5].XIC_dummy_right.icell.SM XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout VGND.t1622 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2849 VGND.t1984 Vbias.t266 XA.XIR[15].XIC_15.icell.SM VGND.t1983 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2850 a_8739_9569# XThC.XTB3.Y.t18 XThC.Tn[10].t7 VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2851 XA.XIR[2].XIC[6].icell.PUM XThC.Tn[6].t43 XA.XIR[2].XIC[6].icell.Ien VPWR.t440 sky130_fd_pr__pfet_01v8 ad=0.0675 pd=0.77 as=0.0725 ps=0.79 w=0.5 l=0.15
X2852 VGND.t810 XThC.Tn[14].t43 XA.XIR[15].XIC[14].icell.PDM VGND.t809 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2853 VGND.t868 XThC.Tn[8].t43 XA.XIR[15].XIC[8].icell.PDM VGND.t867 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2854 VPWR.t1858 XThR.XTBN.Y.t123 XThR.Tn[12].t0 VPWR.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2855 XA.XIR[2].XIC[4].icell.PDM XThR.Tn[2].t73 XA.XIR[2].XIC[4].icell.Ien VGND.t128 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2856 XA.XIR[6].XIC[12].icell.PDM XThR.Tn[6].t73 XA.XIR[6].XIC[12].icell.Ien VGND.t1320 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2857 XA.XIR[5].XIC[13].icell.PDM XThR.Tn[5].t73 XA.XIR[5].XIC[13].icell.Ien VGND.t2545 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2858 XA.XIR[1].XIC[2].icell.SM XA.XIR[1].XIC[2].icell.Ien Iout.t65 VGND.t804 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2859 XA.XIR[9].XIC[13].icell.PDM XThR.Tn[9].t72 XA.XIR[9].XIC[13].icell.Ien VGND.t540 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.2304 ps=2.18 w=0.5 l=0.15
X2860 VPWR.t1415 VPWR.t1413 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR.t1414 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
X2861 VGND.t1873 XThC.Tn[9].t43 XA.XIR[2].XIC[9].icell.PDM VGND.t1872 sky130_fd_pr__nfet_01v8 ad=0.0725 pd=0.79 as=0.0725 ps=0.79 w=0.5 l=0.15
X2862 XA.XIR[4].XIC[3].icell.SM XA.XIR[4].XIC[3].icell.Ien Iout.t3 VGND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.0625 pd=0.75 as=0.175 ps=1.7 w=0.5 l=0.5
X2863 XA.XIR[10].XIC[11].icell.PDM XThR.Tn[9].t73 VGND.t542 VGND.t541 sky130_fd_pr__nfet_01v8 ad=0.1312 pd=1.54 as=0.0725 ps=0.79 w=0.5 l=0.15
X2864 VGND.t1986 Vbias.t267 XA.XIR[13].XIC[2].icell.SM VGND.t1985 sky130_fd_pr__nfet_g5v0d10v5 ad=0.175 pd=1.7 as=0.0625 ps=0.75 w=0.5 l=0.5
X2865 VPWR.t418 XThR.Tn[3].t73 XA.XIR[4].XIC[7].icell.PUM VPWR.t417 sky130_fd_pr__pfet_01v8 ad=0.135 pd=1.54 as=0.0675 ps=0.77 w=0.5 l=0.15
R0 VGND.n2839 VGND.n11 1.04433e+06
R1 VGND.n2839 VGND.n2838 74066.7
R2 VGND.n3017 VGND.n3016 21134.4
R3 VGND.n2875 VGND.n2843 13477
R4 VGND.n2843 VGND.n2842 11635.6
R5 VGND.n3010 VGND.n3009 9309.26
R6 VGND.n2908 VGND.n2875 9223.7
R7 VGND.n2909 VGND.n2908 9223.7
R8 VGND.n2962 VGND.n38 9223.7
R9 VGND.n2995 VGND.n2962 9223.7
R10 VGND.n3016 VGND.n11 8212.42
R11 VGND.n2996 VGND.n2995 7447.41
R12 VGND.n1512 VGND.n1511 7387.65
R13 VGND.n1511 VGND.n1510 7387.65
R14 VGND.n2837 VGND.n151 7387.65
R15 VGND.n3015 VGND.n3014 7387.65
R16 VGND.n3014 VGND.n3013 7387.65
R17 VGND.n3013 VGND.n3012 7387.65
R18 VGND.n3012 VGND.n3011 7387.65
R19 VGND.n3011 VGND.n3010 7387.65
R20 VGND.n2838 VGND.n2837 6977.14
R21 VGND.n1514 VGND.t642 6324.96
R22 VGND.n3016 VGND.n3015 5925.11
R23 VGND.n2909 VGND.n38 5231.11
R24 VGND.n1294 VGND.t2470 5168.13
R25 VGND.n3009 VGND.n3008 5074.71
R26 VGND.n1114 VGND.n582 4539.15
R27 VGND.n3009 VGND 4240.58
R28 VGND.n2418 VGND.n277 4077.12
R29 VGND.n1298 VGND.n1296 3417.39
R30 VGND.n1298 VGND.n1297 3417.39
R31 VGND.n1516 VGND.n1515 3417.39
R32 VGND.n964 VGND.n584 3417.39
R33 VGND.n639 VGND.n181 3417.39
R34 VGND.n2836 VGND.n118 3417.39
R35 VGND.n2841 VGND.n2840 3417.39
R36 VGND.n2419 VGND.n2418 3331.79
R37 VGND.n2420 VGND.n2419 3331.79
R38 VGND.n2421 VGND.n2420 3331.79
R39 VGND.n2422 VGND.n2421 3331.79
R40 VGND.n2423 VGND.n2422 3331.79
R41 VGND.n2424 VGND.n2423 3331.79
R42 VGND.n2425 VGND.n2424 3331.79
R43 VGND.n2426 VGND.n2425 3331.79
R44 VGND.n2427 VGND.n2426 3331.79
R45 VGND.n2428 VGND.n2427 3331.79
R46 VGND.n2429 VGND.n2428 3331.79
R47 VGND.n2430 VGND.n2429 3331.79
R48 VGND.n2431 VGND.n2430 3331.79
R49 VGND.n2431 VGND.n36 3331.79
R50 VGND.n2998 VGND.n36 3331.79
R51 VGND.n2998 VGND.n2997 3331.79
R52 VGND.n1297 VGND.n582 3273.91
R53 VGND.n965 VGND.n583 3265.22
R54 VGND.n2842 VGND.n11 3096.3
R55 VGND.n2839 VGND.n118 2756.52
R56 VGND.n2875 VGND.t311 2655.17
R57 VGND.n2908 VGND.t545 2655.17
R58 VGND.n2997 VGND.n2996 2602.7
R59 VGND.n2837 VGND.n2836 2517.39
R60 VGND.n1296 VGND.n1295 2173.91
R61 VGND.n3028 VGND.n3020 2097.71
R62 VGND.n3020 VGND.n3018 2097.71
R63 VGND.n3019 VGND.n3018 2097.71
R64 VGND.n3028 VGND.n3019 2097.71
R65 VGND.n10 VGND.n6 2097.71
R66 VGND.n3029 VGND.n6 2097.71
R67 VGND.n3029 VGND.n5 2097.71
R68 VGND.n10 VGND.n5 2097.71
R69 VGND.n2842 VGND.n2841 2082.61
R70 VGND VGND.n38 1997.7
R71 VGND.n2962 VGND 1997.7
R72 VGND.n2995 VGND 1997.7
R73 VGND.n1509 VGND.n151 1831.57
R74 VGND.t460 VGND.n2909 1807.04
R75 VGND.n2993 VGND.t371 1785.51
R76 VGND.n1510 VGND.n584 1691.3
R77 VGND.n2921 VGND.t1554 1618.39
R78 VGND.t184 VGND.n2961 1618.39
R79 VGND.t259 VGND.n2994 1618.39
R80 VGND.n2843 VGND.t430 1517.24
R81 VGND.n1513 VGND.n1512 1513.49
R82 VGND.n1514 VGND.n1513 1370.36
R83 VGND.n1513 VGND.t891 1270.28
R84 VGND.n1087 VGND.t410 1268.93
R85 VGND.n1087 VGND.t286 1268.93
R86 VGND.n150 VGND.t326 1253.59
R87 VGND.t100 VGND.n150 1253.59
R88 VGND.n618 VGND.t1333 1253.59
R89 VGND.t287 VGND.n618 1253.59
R90 VGND.n1025 VGND.t207 1253.59
R91 VGND.n1025 VGND.t325 1253.59
R92 VGND.n1056 VGND.t328 1253.59
R93 VGND.n1056 VGND.t103 1253.59
R94 VGND.n180 VGND.t204 1253.59
R95 VGND.t413 VGND.n180 1253.59
R96 VGND.n1295 VGND.n1294 1243.48
R97 VGND.n1509 VGND.t936 1237.71
R98 VGND.n2921 VGND.t1912 1213.79
R99 VGND.n1115 VGND.n1114 1198.25
R100 VGND.n3008 VGND.n3007 1198.25
R101 VGND.n2655 VGND.n37 1180.79
R102 VGND.n3000 VGND.n2999 1180.79
R103 VGND.n2494 VGND.n2493 1180.79
R104 VGND.n2433 VGND.n2432 1180.79
R105 VGND.n2316 VGND.n265 1180.79
R106 VGND.n2130 VGND.n266 1180.79
R107 VGND.n2125 VGND.n267 1180.79
R108 VGND.n2341 VGND.n268 1180.79
R109 VGND.n1956 VGND.n269 1180.79
R110 VGND.n1951 VGND.n270 1180.79
R111 VGND.n2366 VGND.n271 1180.79
R112 VGND.n1782 VGND.n272 1180.79
R113 VGND.n1777 VGND.n273 1180.79
R114 VGND.n2391 VGND.n274 1180.79
R115 VGND.n1608 VGND.n275 1180.79
R116 VGND.n2411 VGND.n276 1180.79
R117 VGND.n1236 VGND.n277 1180.79
R118 VGND.n2417 VGND.n2416 1180.79
R119 VGND.n1293 VGND.n1292 1180.46
R120 VGND.n724 VGND.n683 1180.46
R121 VGND.n729 VGND.n728 1180.46
R122 VGND.n734 VGND.n733 1180.46
R123 VGND.n739 VGND.n738 1180.46
R124 VGND.n744 VGND.n743 1180.46
R125 VGND.n749 VGND.n748 1180.46
R126 VGND.n754 VGND.n753 1180.46
R127 VGND.n759 VGND.n758 1180.46
R128 VGND.n764 VGND.n763 1180.46
R129 VGND.n769 VGND.n768 1180.46
R130 VGND.n774 VGND.n773 1180.46
R131 VGND.n779 VGND.n778 1180.46
R132 VGND.n784 VGND.n783 1180.46
R133 VGND.n786 VGND.n785 1180.46
R134 VGND.n1233 VGND.n1232 1180.46
R135 VGND.n1231 VGND.n1230 1180.46
R136 VGND.n1214 VGND.n1213 1180.46
R137 VGND.n1212 VGND.n1211 1180.46
R138 VGND.n1201 VGND.n1200 1180.46
R139 VGND.n1199 VGND.n1198 1180.46
R140 VGND.n1182 VGND.n1181 1180.46
R141 VGND.n1180 VGND.n1179 1180.46
R142 VGND.n1169 VGND.n1168 1180.46
R143 VGND.n1167 VGND.n1166 1180.46
R144 VGND.n1150 VGND.n1149 1180.46
R145 VGND.n1148 VGND.n1147 1180.46
R146 VGND.n1137 VGND.n1136 1180.46
R147 VGND.n1135 VGND.n1134 1180.46
R148 VGND.n1127 VGND.n1126 1180.46
R149 VGND.n2582 VGND.n2581 1180.46
R150 VGND.n2710 VGND.n2709 1180.46
R151 VGND.n2708 VGND.n2707 1180.46
R152 VGND.n2702 VGND.n2701 1180.46
R153 VGND.n2700 VGND.n2699 1180.46
R154 VGND.n2694 VGND.n2693 1180.46
R155 VGND.n2692 VGND.n2691 1180.46
R156 VGND.n2686 VGND.n2685 1180.46
R157 VGND.n2684 VGND.n2683 1180.46
R158 VGND.n2678 VGND.n2677 1180.46
R159 VGND.n2676 VGND.n2675 1180.46
R160 VGND.n2670 VGND.n2669 1180.46
R161 VGND.n2668 VGND.n2667 1180.46
R162 VGND.n2662 VGND.n2661 1180.46
R163 VGND.n2660 VGND.n2659 1180.46
R164 VGND.n238 VGND.n237 1180.46
R165 VGND.n2723 VGND.n2722 1180.46
R166 VGND.n2728 VGND.n2727 1180.46
R167 VGND.n2733 VGND.n2732 1180.46
R168 VGND.n2738 VGND.n2737 1180.46
R169 VGND.n2743 VGND.n2742 1180.46
R170 VGND.n2748 VGND.n2747 1180.46
R171 VGND.n2753 VGND.n2752 1180.46
R172 VGND.n2758 VGND.n2757 1180.46
R173 VGND.n2763 VGND.n2762 1180.46
R174 VGND.n2768 VGND.n2767 1180.46
R175 VGND.n2773 VGND.n2772 1180.46
R176 VGND.n2778 VGND.n2777 1180.46
R177 VGND.n2783 VGND.n2782 1180.46
R178 VGND.n2785 VGND.n2784 1180.46
R179 VGND.n2519 VGND.n2518 1180.46
R180 VGND.n2517 VGND.n2516 1180.46
R181 VGND.n2512 VGND.n2511 1180.46
R182 VGND.n2437 VGND.n248 1180.46
R183 VGND.n2442 VGND.n2441 1180.46
R184 VGND.n2447 VGND.n2446 1180.46
R185 VGND.n2452 VGND.n2451 1180.46
R186 VGND.n2457 VGND.n2456 1180.46
R187 VGND.n2462 VGND.n2461 1180.46
R188 VGND.n2467 VGND.n2466 1180.46
R189 VGND.n2472 VGND.n2471 1180.46
R190 VGND.n2477 VGND.n2476 1180.46
R191 VGND.n2482 VGND.n2481 1180.46
R192 VGND.n2487 VGND.n2486 1180.46
R193 VGND.n2492 VGND.n2491 1180.46
R194 VGND.n2835 VGND.n2834 1180.46
R195 VGND.n375 VGND.n186 1180.46
R196 VGND.n377 VGND.n376 1180.46
R197 VGND.n2175 VGND.n2174 1180.46
R198 VGND.n2177 VGND.n2176 1180.46
R199 VGND.n2201 VGND.n2200 1180.46
R200 VGND.n2203 VGND.n2202 1180.46
R201 VGND.n2227 VGND.n2226 1180.46
R202 VGND.n2229 VGND.n2228 1180.46
R203 VGND.n2253 VGND.n2252 1180.46
R204 VGND.n2255 VGND.n2254 1180.46
R205 VGND.n2284 VGND.n2283 1180.46
R206 VGND.n2289 VGND.n2288 1180.46
R207 VGND.n2294 VGND.n2293 1180.46
R208 VGND.n2296 VGND.n2295 1180.46
R209 VGND.n1432 VGND.n1431 1180.46
R210 VGND.n1434 VGND.n1433 1180.46
R211 VGND.n2162 VGND.n2161 1180.46
R212 VGND.n2164 VGND.n2163 1180.46
R213 VGND.n2188 VGND.n2187 1180.46
R214 VGND.n2190 VGND.n2189 1180.46
R215 VGND.n2214 VGND.n2213 1180.46
R216 VGND.n2216 VGND.n2215 1180.46
R217 VGND.n2240 VGND.n2239 1180.46
R218 VGND.n2242 VGND.n2241 1180.46
R219 VGND.n2266 VGND.n2265 1180.46
R220 VGND.n2273 VGND.n2272 1180.46
R221 VGND.n2271 VGND.n2270 1180.46
R222 VGND.n2311 VGND.n2310 1180.46
R223 VGND.n2313 VGND.n2312 1180.46
R224 VGND.n1446 VGND.n1445 1180.46
R225 VGND.n1498 VGND.n1497 1180.46
R226 VGND.n1496 VGND.n1495 1180.46
R227 VGND.n1491 VGND.n1490 1180.46
R228 VGND.n1486 VGND.n1485 1180.46
R229 VGND.n1481 VGND.n1480 1180.46
R230 VGND.n1476 VGND.n1475 1180.46
R231 VGND.n1471 VGND.n1470 1180.46
R232 VGND.n1466 VGND.n1465 1180.46
R233 VGND.n1461 VGND.n1460 1180.46
R234 VGND.n1456 VGND.n1455 1180.46
R235 VGND.n1451 VGND.n1450 1180.46
R236 VGND.n2141 VGND.n2140 1180.46
R237 VGND.n2139 VGND.n2138 1180.46
R238 VGND.n2134 VGND.n2133 1180.46
R239 VGND.n1508 VGND.n1507 1180.46
R240 VGND.n630 VGND.n623 1180.46
R241 VGND.n632 VGND.n631 1180.46
R242 VGND.n2001 VGND.n2000 1180.46
R243 VGND.n2003 VGND.n2002 1180.46
R244 VGND.n2027 VGND.n2026 1180.46
R245 VGND.n2029 VGND.n2028 1180.46
R246 VGND.n2053 VGND.n2052 1180.46
R247 VGND.n2055 VGND.n2054 1180.46
R248 VGND.n2079 VGND.n2078 1180.46
R249 VGND.n2081 VGND.n2080 1180.46
R250 VGND.n2110 VGND.n2109 1180.46
R251 VGND.n2115 VGND.n2114 1180.46
R252 VGND.n2120 VGND.n2119 1180.46
R253 VGND.n2122 VGND.n2121 1180.46
R254 VGND.n656 VGND.n655 1180.46
R255 VGND.n658 VGND.n657 1180.46
R256 VGND.n1988 VGND.n1987 1180.46
R257 VGND.n1990 VGND.n1989 1180.46
R258 VGND.n2014 VGND.n2013 1180.46
R259 VGND.n2016 VGND.n2015 1180.46
R260 VGND.n2040 VGND.n2039 1180.46
R261 VGND.n2042 VGND.n2041 1180.46
R262 VGND.n2066 VGND.n2065 1180.46
R263 VGND.n2068 VGND.n2067 1180.46
R264 VGND.n2092 VGND.n2091 1180.46
R265 VGND.n2099 VGND.n2098 1180.46
R266 VGND.n2097 VGND.n2096 1180.46
R267 VGND.n2336 VGND.n2335 1180.46
R268 VGND.n2338 VGND.n2337 1180.46
R269 VGND.n963 VGND.n962 1180.46
R270 VGND.n958 VGND.n957 1180.46
R271 VGND.n953 VGND.n952 1180.46
R272 VGND.n948 VGND.n947 1180.46
R273 VGND.n943 VGND.n942 1180.46
R274 VGND.n938 VGND.n937 1180.46
R275 VGND.n933 VGND.n932 1180.46
R276 VGND.n928 VGND.n927 1180.46
R277 VGND.n923 VGND.n922 1180.46
R278 VGND.n918 VGND.n917 1180.46
R279 VGND.n913 VGND.n912 1180.46
R280 VGND.n908 VGND.n907 1180.46
R281 VGND.n1967 VGND.n1966 1180.46
R282 VGND.n1965 VGND.n1964 1180.46
R283 VGND.n1960 VGND.n1959 1180.46
R284 VGND.n1399 VGND.n1398 1180.46
R285 VGND.n1404 VGND.n1403 1180.46
R286 VGND.n1406 VGND.n1405 1180.46
R287 VGND.n1827 VGND.n1826 1180.46
R288 VGND.n1829 VGND.n1828 1180.46
R289 VGND.n1853 VGND.n1852 1180.46
R290 VGND.n1855 VGND.n1854 1180.46
R291 VGND.n1879 VGND.n1878 1180.46
R292 VGND.n1881 VGND.n1880 1180.46
R293 VGND.n1905 VGND.n1904 1180.46
R294 VGND.n1907 VGND.n1906 1180.46
R295 VGND.n1936 VGND.n1935 1180.46
R296 VGND.n1941 VGND.n1940 1180.46
R297 VGND.n1946 VGND.n1945 1180.46
R298 VGND.n1948 VGND.n1947 1180.46
R299 VGND.n1384 VGND.n1383 1180.46
R300 VGND.n1386 VGND.n1385 1180.46
R301 VGND.n1814 VGND.n1813 1180.46
R302 VGND.n1816 VGND.n1815 1180.46
R303 VGND.n1840 VGND.n1839 1180.46
R304 VGND.n1842 VGND.n1841 1180.46
R305 VGND.n1866 VGND.n1865 1180.46
R306 VGND.n1868 VGND.n1867 1180.46
R307 VGND.n1892 VGND.n1891 1180.46
R308 VGND.n1894 VGND.n1893 1180.46
R309 VGND.n1918 VGND.n1917 1180.46
R310 VGND.n1925 VGND.n1924 1180.46
R311 VGND.n1923 VGND.n1922 1180.46
R312 VGND.n2361 VGND.n2360 1180.46
R313 VGND.n2363 VGND.n2362 1180.46
R314 VGND.n1316 VGND.n1315 1180.46
R315 VGND.n1368 VGND.n1367 1180.46
R316 VGND.n1366 VGND.n1365 1180.46
R317 VGND.n1361 VGND.n1360 1180.46
R318 VGND.n1356 VGND.n1355 1180.46
R319 VGND.n1351 VGND.n1350 1180.46
R320 VGND.n1346 VGND.n1345 1180.46
R321 VGND.n1341 VGND.n1340 1180.46
R322 VGND.n1336 VGND.n1335 1180.46
R323 VGND.n1331 VGND.n1330 1180.46
R324 VGND.n1326 VGND.n1325 1180.46
R325 VGND.n1321 VGND.n1320 1180.46
R326 VGND.n1793 VGND.n1792 1180.46
R327 VGND.n1791 VGND.n1790 1180.46
R328 VGND.n1786 VGND.n1785 1180.46
R329 VGND.n1521 VGND.n1520 1180.46
R330 VGND.n1526 VGND.n1525 1180.46
R331 VGND.n1528 VGND.n1527 1180.46
R332 VGND.n1653 VGND.n1652 1180.46
R333 VGND.n1655 VGND.n1654 1180.46
R334 VGND.n1679 VGND.n1678 1180.46
R335 VGND.n1681 VGND.n1680 1180.46
R336 VGND.n1705 VGND.n1704 1180.46
R337 VGND.n1707 VGND.n1706 1180.46
R338 VGND.n1731 VGND.n1730 1180.46
R339 VGND.n1733 VGND.n1732 1180.46
R340 VGND.n1762 VGND.n1761 1180.46
R341 VGND.n1767 VGND.n1766 1180.46
R342 VGND.n1772 VGND.n1771 1180.46
R343 VGND.n1774 VGND.n1773 1180.46
R344 VGND.n1541 VGND.n1540 1180.46
R345 VGND.n1543 VGND.n1542 1180.46
R346 VGND.n1640 VGND.n1639 1180.46
R347 VGND.n1642 VGND.n1641 1180.46
R348 VGND.n1666 VGND.n1665 1180.46
R349 VGND.n1668 VGND.n1667 1180.46
R350 VGND.n1692 VGND.n1691 1180.46
R351 VGND.n1694 VGND.n1693 1180.46
R352 VGND.n1718 VGND.n1717 1180.46
R353 VGND.n1720 VGND.n1719 1180.46
R354 VGND.n1744 VGND.n1743 1180.46
R355 VGND.n1751 VGND.n1750 1180.46
R356 VGND.n1749 VGND.n1748 1180.46
R357 VGND.n2386 VGND.n2385 1180.46
R358 VGND.n2388 VGND.n2387 1180.46
R359 VGND.n1300 VGND.n1299 1180.46
R360 VGND.n1554 VGND.n1553 1180.46
R361 VGND.n1559 VGND.n1558 1180.46
R362 VGND.n1564 VGND.n1563 1180.46
R363 VGND.n1569 VGND.n1568 1180.46
R364 VGND.n1574 VGND.n1573 1180.46
R365 VGND.n1579 VGND.n1578 1180.46
R366 VGND.n1584 VGND.n1583 1180.46
R367 VGND.n1589 VGND.n1588 1180.46
R368 VGND.n1594 VGND.n1593 1180.46
R369 VGND.n1599 VGND.n1598 1180.46
R370 VGND.n1604 VGND.n1603 1180.46
R371 VGND.n1619 VGND.n1618 1180.46
R372 VGND.n1617 VGND.n1616 1180.46
R373 VGND.n1612 VGND.n1611 1180.46
R374 VGND.n839 VGND.n838 1180.46
R375 VGND.n844 VGND.n843 1180.46
R376 VGND.n896 VGND.n895 1180.46
R377 VGND.n894 VGND.n893 1180.46
R378 VGND.n889 VGND.n888 1180.46
R379 VGND.n884 VGND.n883 1180.46
R380 VGND.n879 VGND.n878 1180.46
R381 VGND.n874 VGND.n873 1180.46
R382 VGND.n869 VGND.n868 1180.46
R383 VGND.n864 VGND.n863 1180.46
R384 VGND.n859 VGND.n858 1180.46
R385 VGND.n854 VGND.n853 1180.46
R386 VGND.n849 VGND.n848 1180.46
R387 VGND.n2406 VGND.n2405 1180.46
R388 VGND.n2408 VGND.n2407 1180.46
R389 VGND.n2961 VGND.t202 1180.08
R390 VGND.n1515 VGND.n1514 1169.57
R391 VGND.n3013 VGND.t1634 1146.36
R392 VGND.n3015 VGND.t1633 1112.64
R393 VGND.n3014 VGND.t2645 1112.64
R394 VGND.n2996 VGND 1055.35
R395 VGND.n1510 VGND.n1509 1052.29
R396 VGND.t1197 VGND.n7 1041.38
R397 VGND.t1197 VGND.n3017 1041.38
R398 VGND.t2274 VGND.n965 1032.59
R399 VGND.t694 VGND.n2582 988.926
R400 VGND.n2709 VGND.t2498 988.926
R401 VGND.n2708 VGND.t2476 988.926
R402 VGND.n2701 VGND.t692 988.926
R403 VGND.n2700 VGND.t681 988.926
R404 VGND.n2693 VGND.t1684 988.926
R405 VGND.n2692 VGND.t762 988.926
R406 VGND.n2685 VGND.t739 988.926
R407 VGND.n2684 VGND.t1680 988.926
R408 VGND.n2677 VGND.t2460 988.926
R409 VGND.n2676 VGND.t2448 988.926
R410 VGND.n2669 VGND.t710 988.926
R411 VGND.n2668 VGND.t1667 988.926
R412 VGND.n2661 VGND.t2436 988.926
R413 VGND.n2660 VGND.t724 988.926
R414 VGND.n237 VGND.t1148 988.926
R415 VGND.t2258 VGND.n2723 988.926
R416 VGND.t129 VGND.n2728 988.926
R417 VGND.t1388 VGND.n2733 988.926
R418 VGND.t1967 VGND.n2738 988.926
R419 VGND.t161 VGND.n2743 988.926
R420 VGND.t2407 VGND.n2748 988.926
R421 VGND.t1755 VGND.n2753 988.926
R422 VGND.t471 VGND.n2758 988.926
R423 VGND.t537 VGND.n2763 988.926
R424 VGND.t876 VGND.n2768 988.926
R425 VGND.t1862 VGND.n2773 988.926
R426 VGND.t305 VGND.n2778 988.926
R427 VGND.t1806 VGND.n2783 988.926
R428 VGND.n2784 VGND.t1507 988.926
R429 VGND.n2518 VGND.t828 988.926
R430 VGND.n2517 VGND.t2680 988.926
R431 VGND.n2512 VGND.t770 988.926
R432 VGND.t600 VGND.n2437 988.926
R433 VGND.t648 VGND.n2442 988.926
R434 VGND.t1538 VGND.n2447 988.926
R435 VGND.t665 VGND.n2452 988.926
R436 VGND.t2687 VGND.n2457 988.926
R437 VGND.t1134 VGND.n2462 988.926
R438 VGND.t520 VGND.n2467 988.926
R439 VGND.t1918 VGND.n2472 988.926
R440 VGND.t1832 VGND.n2477 988.926
R441 VGND.t2196 VGND.n2482 988.926
R442 VGND.t1826 VGND.n2487 988.926
R443 VGND.t91 VGND.n2492 988.926
R444 VGND.n2835 VGND.t1343 988.926
R445 VGND.t1994 VGND.n375 988.926
R446 VGND.n376 VGND.t96 988.926
R447 VGND.t1164 VGND.n2175 988.926
R448 VGND.n2176 VGND.t1710 988.926
R449 VGND.t1562 VGND.n2201 988.926
R450 VGND.n2202 VGND.t1311 988.926
R451 VGND.t375 VGND.n2227 988.926
R452 VGND.n2228 VGND.t118 988.926
R453 VGND.t28 VGND.n2253 988.926
R454 VGND.n2254 VGND.t2045 988.926
R455 VGND.t2612 VGND.n2284 988.926
R456 VGND.t393 VGND.n2289 988.926
R457 VGND.t109 VGND.n2294 988.926
R458 VGND.n2295 VGND.t1514 988.926
R459 VGND.t1931 VGND.n1432 988.926
R460 VGND.n1433 VGND.t2164 988.926
R461 VGND.t151 VGND.n2162 988.926
R462 VGND.n2163 VGND.t66 988.926
R463 VGND.t2083 VGND.n2188 988.926
R464 VGND.n2189 VGND.t136 988.926
R465 VGND.t2399 VGND.n2214 988.926
R466 VGND.n2215 VGND.t1068 988.926
R467 VGND.t1157 VGND.n2240 988.926
R468 VGND.n2241 VGND.t563 988.926
R469 VGND.t1445 VGND.n2266 988.926
R470 VGND.n2272 VGND.t172 988.926
R471 VGND.n2271 VGND.t1793 988.926
R472 VGND.t1815 VGND.n2311 988.926
R473 VGND.n2312 VGND.t2131 988.926
R474 VGND.t466 VGND.n1446 988.926
R475 VGND.n1497 VGND.t837 988.926
R476 VGND.n1496 VGND.t812 988.926
R477 VGND.n1491 VGND.t2514 988.926
R478 VGND.n1486 VGND.t2147 988.926
R479 VGND.n1481 VGND.t1905 988.926
R480 VGND.n1476 VGND.t1318 988.926
R481 VGND.n1471 VGND.t368 988.926
R482 VGND.n1466 VGND.t841 988.926
R483 VGND.n1461 VGND.t515 988.926
R484 VGND.n1456 VGND.t2532 988.926
R485 VGND.n1451 VGND.t2589 988.926
R486 VGND.n2140 VGND.t400 988.926
R487 VGND.n2139 VGND.t1111 988.926
R488 VGND.n2134 VGND.t2115 988.926
R489 VGND.n1508 VGND.t1146 988.926
R490 VGND.t2256 VGND.n630 988.926
R491 VGND.n631 VGND.t126 988.926
R492 VGND.t1386 VGND.n2001 988.926
R493 VGND.n2002 VGND.t1965 988.926
R494 VGND.t159 VGND.n2027 988.926
R495 VGND.n2028 VGND.t2405 988.926
R496 VGND.t1753 VGND.n2053 988.926
R497 VGND.n2054 VGND.t469 988.926
R498 VGND.t534 VGND.n2079 988.926
R499 VGND.n2080 VGND.t874 988.926
R500 VGND.t1859 VGND.n2110 988.926
R501 VGND.t303 VGND.n2115 988.926
R502 VGND.t1817 VGND.n2120 988.926
R503 VGND.n2121 VGND.t1505 988.926
R504 VGND.t1345 VGND.n656 988.926
R505 VGND.n657 VGND.t1996 988.926
R506 VGND.t94 VGND.n1988 988.926
R507 VGND.n1989 VGND.t1166 988.926
R508 VGND.t1712 VGND.n2014 988.926
R509 VGND.n2015 VGND.t1564 988.926
R510 VGND.t1313 VGND.n2040 988.926
R511 VGND.n2041 VGND.t377 988.926
R512 VGND.t120 VGND.n2066 988.926
R513 VGND.n2067 VGND.t30 988.926
R514 VGND.t2047 VGND.n2092 988.926
R515 VGND.n2098 VGND.t2614 988.926
R516 VGND.n2097 VGND.t395 988.926
R517 VGND.t111 VGND.n2336 988.926
R518 VGND.n2337 VGND.t2109 988.926
R519 VGND.n963 VGND.t1933 988.926
R520 VGND.n958 VGND.t2166 988.926
R521 VGND.n953 VGND.t149 988.926
R522 VGND.n948 VGND.t68 988.926
R523 VGND.n943 VGND.t1603 988.926
R524 VGND.n938 VGND.t138 988.926
R525 VGND.n933 VGND.t2401 988.926
R526 VGND.n928 VGND.t1070 988.926
R527 VGND.n923 VGND.t1159 988.926
R528 VGND.n918 VGND.t565 988.926
R529 VGND.n913 VGND.t1447 988.926
R530 VGND.n908 VGND.t1104 988.926
R531 VGND.n1966 VGND.t1795 988.926
R532 VGND.n1965 VGND.t1031 988.926
R533 VGND.n1960 VGND.t1501 988.926
R534 VGND.t1926 VGND.n1399 988.926
R535 VGND.t1294 VGND.n1404 988.926
R536 VGND.n1405 VGND.t155 988.926
R537 VGND.t62 VGND.n1827 988.926
R538 VGND.n1828 VGND.t2077 988.926
R539 VGND.t134 VGND.n1853 988.926
R540 VGND.n1854 VGND.t2666 988.926
R541 VGND.t385 VGND.n1879 988.926
R542 VGND.n1880 VGND.t1463 988.926
R543 VGND.t561 VGND.n1905 988.926
R544 VGND.n1906 VGND.t1443 988.926
R545 VGND.t170 VGND.n1936 988.926
R546 VGND.t589 VGND.n1941 988.926
R547 VGND.t1811 VGND.n1946 988.926
R548 VGND.n1947 VGND.t2129 988.926
R549 VGND.t464 VGND.n1384 988.926
R550 VGND.n1385 VGND.t835 988.926
R551 VGND.t814 VGND.n1814 988.926
R552 VGND.n1815 VGND.t2512 988.926
R553 VGND.t282 VGND.n1840 988.926
R554 VGND.n1841 VGND.t1903 988.926
R555 VGND.t1316 VGND.n1866 988.926
R556 VGND.n1867 VGND.t366 988.926
R557 VGND.t839 VGND.n1892 988.926
R558 VGND.n1893 VGND.t513 988.926
R559 VGND.t2530 VGND.n1918 988.926
R560 VGND.n1924 VGND.t2595 988.926
R561 VGND.n1923 VGND.t398 988.926
R562 VGND.t1109 VGND.n2361 988.926
R563 VGND.n2362 VGND.t2113 988.926
R564 VGND.t1123 VGND.n1316 988.926
R565 VGND.n1367 VGND.t1971 988.926
R566 VGND.n1366 VGND.t142 988.926
R567 VGND.n1361 VGND.t1194 988.926
R568 VGND.n1356 VGND.t2247 988.926
R569 VGND.n1351 VGND.t2541 988.926
R570 VGND.n1346 VGND.t2659 988.926
R571 VGND.n1341 VGND.t391 988.926
R572 VGND.n1336 VGND.t1458 988.926
R573 VGND.n1331 VGND.t532 988.926
R574 VGND.n1326 VGND.t2563 988.926
R575 VGND.n1321 VGND.t2548 988.926
R576 VGND.n1792 VGND.t2204 988.926
R577 VGND.n1791 VGND.t2039 988.926
R578 VGND.n1786 VGND.t2121 988.926
R579 VGND.t1341 VGND.n1521 988.926
R580 VGND.t1992 VGND.n1526 988.926
R581 VGND.n1527 VGND.t98 988.926
R582 VGND.t1162 VGND.n1653 988.926
R583 VGND.n1654 VGND.t1708 988.926
R584 VGND.t1560 VGND.n1679 988.926
R585 VGND.n1680 VGND.t1309 988.926
R586 VGND.t373 VGND.n1705 988.926
R587 VGND.n1706 VGND.t116 988.926
R588 VGND.t541 VGND.n1731 988.926
R589 VGND.n1732 VGND.t2043 988.926
R590 VGND.t2610 VGND.n1762 988.926
R591 VGND.t309 VGND.n1767 988.926
R592 VGND.t107 VGND.n1772 988.926
R593 VGND.n1773 VGND.t1512 988.926
R594 VGND.t1121 VGND.n1541 988.926
R595 VGND.n1542 VGND.t1969 988.926
R596 VGND.t144 VGND.n1640 988.926
R597 VGND.n1641 VGND.t1192 988.926
R598 VGND.t2245 VGND.n1666 988.926
R599 VGND.n1667 VGND.t2551 988.926
R600 VGND.t2657 VGND.n1692 988.926
R601 VGND.n1693 VGND.t389 988.926
R602 VGND.t1456 VGND.n1718 988.926
R603 VGND.n1719 VGND.t530 988.926
R604 VGND.t2561 VGND.n1744 988.926
R605 VGND.n1750 VGND.t2546 988.926
R606 VGND.n1749 VGND.t2202 988.926
R607 VGND.t1821 VGND.n2386 988.926
R608 VGND.n2387 VGND.t2119 988.926
R609 VGND.n1299 VGND.t826 988.926
R610 VGND.t2678 VGND.n1554 988.926
R611 VGND.t773 VGND.n1559 988.926
R612 VGND.t2518 VGND.n1564 988.926
R613 VGND.t2151 VGND.n1569 988.926
R614 VGND.t1907 VGND.n1574 988.926
R615 VGND.t663 VGND.n1579 988.926
R616 VGND.t2685 VGND.n1584 988.926
R617 VGND.t1132 VGND.n1589 988.926
R618 VGND.t517 VGND.n1594 988.926
R619 VGND.t1916 VGND.n1599 988.926
R620 VGND.t2591 VGND.n1604 988.926
R621 VGND.n1618 VGND.t404 988.926
R622 VGND.n1617 VGND.t1823 988.926
R623 VGND.n1612 VGND.t88 988.926
R624 VGND.t1928 VGND.n839 988.926
R625 VGND.t1296 VGND.n844 988.926
R626 VGND.n895 VGND.t153 988.926
R627 VGND.n894 VGND.t64 988.926
R628 VGND.n889 VGND.t2079 988.926
R629 VGND.n884 VGND.t132 988.926
R630 VGND.n879 VGND.t2664 988.926
R631 VGND.n874 VGND.t383 988.926
R632 VGND.n869 VGND.t1461 988.926
R633 VGND.n864 VGND.t559 988.926
R634 VGND.n859 VGND.t1441 988.926
R635 VGND.n854 VGND.t168 988.926
R636 VGND.n849 VGND.t587 988.926
R637 VGND.t1813 VGND.n2406 988.926
R638 VGND.n2407 VGND.t2127 988.926
R639 VGND.n1293 VGND.t1663 988.926
R640 VGND.t2442 VGND.n724 988.926
R641 VGND.t2420 VGND.n729 988.926
R642 VGND.t1658 VGND.n734 988.926
R643 VGND.t1647 VGND.n739 988.926
R644 VGND.t2489 VGND.n744 988.926
R645 VGND.t704 VGND.n749 988.926
R646 VGND.t683 VGND.n754 988.926
R647 VGND.t2485 VGND.n759 988.926
R648 VGND.t764 VGND.n764 988.926
R649 VGND.t751 VGND.n769 988.926
R650 VGND.t1682 VGND.n774 988.926
R651 VGND.t2468 VGND.n779 988.926
R652 VGND.t733 VGND.n784 988.926
R653 VGND.n785 VGND.t1691 988.926
R654 VGND.n1512 VGND.n583 934.784
R655 VGND.n2907 VGND 927.203
R656 VGND.n2910 VGND 927.203
R657 VGND.n966 VGND 918.774
R658 VGND.n117 VGND 910.346
R659 VGND.n2874 VGND 910.346
R660 VGND.n3008 VGND.t1750 909.365
R661 VGND.n2837 VGND.n181 900
R662 VGND.n2582 VGND.t1465 852.769
R663 VGND.n2709 VGND.t1957 852.769
R664 VGND.t1403 VGND.n2708 852.769
R665 VGND.n2701 VGND.t420 852.769
R666 VGND.t1953 VGND.n2700 852.769
R667 VGND.n2693 VGND.t869 852.769
R668 VGND.t1269 VGND.n2692 852.769
R669 VGND.n2685 VGND.t158 852.769
R670 VGND.t1327 VGND.n2684 852.769
R671 VGND.n2677 VGND.t75 852.769
R672 VGND.t250 VGND.n2676 852.769
R673 VGND.n2669 VGND.t639 852.769
R674 VGND.t2141 VGND.n2668 852.769
R675 VGND.n2661 VGND.t1142 852.769
R676 VGND.t175 VGND.n2660 852.769
R677 VGND.t1924 VGND.n37 852.769
R678 VGND.n237 VGND.t2504 852.769
R679 VGND.n2723 VGND.t79 852.769
R680 VGND.n2728 VGND.t2619 852.769
R681 VGND.n2733 VGND.t1118 852.769
R682 VGND.n2738 VGND.t1326 852.769
R683 VGND.n2743 VGND.t1144 852.769
R684 VGND.n2748 VGND.t1400 852.769
R685 VGND.n2753 VGND.t179 852.769
R686 VGND.n2758 VGND.t83 852.769
R687 VGND.n2763 VGND.t2607 852.769
R688 VGND.n2768 VGND.t1322 852.769
R689 VGND.n2773 VGND.t1139 852.769
R690 VGND.n2778 VGND.t803 852.769
R691 VGND.n2783 VGND.t1321 852.769
R692 VGND.n2784 VGND.t475 852.769
R693 VGND.n2999 VGND.t1431 852.769
R694 VGND.n2518 VGND.t1804 852.769
R695 VGND.t225 VGND.n2517 852.769
R696 VGND.t1392 VGND.n2512 852.769
R697 VGND.n2437 VGND.t1614 852.769
R698 VGND.n2442 VGND.t82 852.769
R699 VGND.n2447 VGND.t2654 852.769
R700 VGND.n2452 VGND.t1339 852.769
R701 VGND.n2457 VGND.t1535 852.769
R702 VGND.n2462 VGND.t1143 852.769
R703 VGND.n2467 VGND.t1591 852.769
R704 VGND.n2472 VGND.t1915 852.769
R705 VGND.n2477 VGND.t641 852.769
R706 VGND.n2482 VGND.t2206 852.769
R707 VGND.n2487 VGND.t1518 852.769
R708 VGND.n2492 VGND.t58 852.769
R709 VGND.n2493 VGND.t1 852.769
R710 VGND.t865 VGND.n2835 852.769
R711 VGND.n375 VGND.t804 852.769
R712 VGND.n376 VGND.t2508 852.769
R713 VGND.n2175 VGND.t872 852.769
R714 VGND.n2176 VGND.t1958 852.769
R715 VGND.n2201 VGND.t1799 852.769
R716 VGND.n2202 VGND.t203 852.769
R717 VGND.n2227 VGND.t115 852.769
R718 VGND.n2228 VGND.t1914 852.769
R719 VGND.n2253 VGND.t1300 852.769
R720 VGND.n2254 VGND.t2523 852.769
R721 VGND.n2284 VGND.t1640 852.769
R722 VGND.n2289 VGND.t1517 852.769
R723 VGND.n2294 VGND.t1152 852.769
R724 VGND.n2295 VGND.t886 852.769
R725 VGND.n2432 VGND.t1618 852.769
R726 VGND.n1432 VGND.t279 852.769
R727 VGND.n1433 VGND.t193 852.769
R728 VGND.n2162 VGND.t2675 852.769
R729 VGND.n2163 VGND.t1125 852.769
R730 VGND.n2188 VGND.t70 852.769
R731 VGND.n2189 VGND.t1790 852.769
R732 VGND.n2214 VGND.t1141 852.769
R733 VGND.n2215 VGND.t178 852.769
R734 VGND.n2240 VGND.t1800 852.769
R735 VGND.n2241 VGND.t646 852.769
R736 VGND.n2266 VGND.t1935 852.769
R737 VGND.n2272 VGND.t1277 852.769
R738 VGND.t2522 VGND.n2271 852.769
R739 VGND.n2311 VGND.t1798 852.769
R740 VGND.n2312 VGND.t1642 852.769
R741 VGND.t86 VGND.n265 852.769
R742 VGND.n1446 VGND.t844 852.769
R743 VGND.n1497 VGND.t253 852.769
R744 VGND.t1268 VGND.n1496 852.769
R745 VGND.t871 VGND.n1491 852.769
R746 VGND.t1789 VGND.n1486 852.769
R747 VGND.t27 VGND.n1481 852.769
R748 VGND.t2506 VGND.n1476 852.769
R749 VGND.t1153 VGND.n1471 852.769
R750 VGND.t2142 VGND.n1466 852.769
R751 VGND.t1519 VGND.n1461 852.769
R752 VGND.t292 VGND.n1456 852.769
R753 VGND.t1533 VGND.n1451 852.769
R754 VGND.n2140 VGND.t870 852.769
R755 VGND.t2509 VGND.n2139 852.769
R756 VGND.t1270 VGND.n2134 852.769
R757 VGND.t210 VGND.n266 852.769
R758 VGND.t1401 VGND.n1508 852.769
R759 VGND.n630 VGND.t78 852.769
R760 VGND.n631 VGND.t1955 852.769
R761 VGND.n2001 VGND.t1337 852.769
R762 VGND.n2002 VGND.t888 852.769
R763 VGND.n2027 VGND.t252 852.769
R764 VGND.n2028 VGND.t1278 852.769
R765 VGND.n2053 VGND.t2617 852.769
R766 VGND.n2054 VGND.t2539 852.769
R767 VGND.n2079 VGND.t1438 852.769
R768 VGND.n2080 VGND.t1770 852.769
R769 VGND.n2110 VGND.t645 852.769
R770 VGND.n2115 VGND.t114 852.769
R771 VGND.n2120 VGND.t224 852.769
R772 VGND.n2121 VGND.t1875 852.769
R773 VGND.t1127 VGND.n267 852.769
R774 VGND.n656 VGND.t2505 852.769
R775 VGND.n657 VGND.t1394 852.769
R776 VGND.n1988 VGND.t1923 852.769
R777 VGND.n1989 VGND.t1129 852.769
R778 VGND.n2014 VGND.t2538 852.769
R779 VGND.n2015 VGND.t1128 852.769
R780 VGND.n2040 VGND.t2556 852.769
R781 VGND.n2041 VGND.t211 852.769
R782 VGND.n2066 VGND.t1429 852.769
R783 VGND.n2067 VGND.t1455 852.769
R784 VGND.n2092 VGND.t880 852.769
R785 VGND.n2098 VGND.t1617 852.769
R786 VGND.t1874 VGND.n2097 852.769
R787 VGND.n2336 VGND.t85 852.769
R788 VGND.n2337 VGND.t266 852.769
R789 VGND.t1771 VGND.n268 852.769
R790 VGND.t1639 VGND.n963 852.769
R791 VGND.t864 VGND.n958 852.769
R792 VGND.t123 VGND.n953 852.769
R793 VGND.t76 VGND.n948 852.769
R794 VGND.t180 VGND.n943 852.769
R795 VGND.t1138 VGND.n938 852.769
R796 VGND.t583 VGND.n933 852.769
R797 VGND.t1042 VGND.n928 852.769
R798 VGND.t1532 VGND.n923 852.769
R799 VGND.t1613 VGND.n918 852.769
R800 VGND.t1525 VGND.n913 852.769
R801 VGND.t2310 VGND.n908 852.769
R802 VGND.n1966 VGND.t1522 852.769
R803 VGND.t421 VGND.n1965 852.769
R804 VGND.t1324 VGND.n1960 852.769
R805 VGND.t680 VGND.n269 852.769
R806 VGND.n1399 VGND.t830 852.769
R807 VGND.n1404 VGND.t2618 852.769
R808 VGND.n1405 VGND.t881 852.769
R809 VGND.n1827 VGND.t2648 852.769
R810 VGND.n1828 VGND.t805 852.769
R811 VGND.n1853 VGND.t1119 852.769
R812 VGND.n1854 VGND.t2520 852.769
R813 VGND.n1879 VGND.t2145 852.769
R814 VGND.n1880 VGND.t1772 852.769
R815 VGND.n1905 VGND.t1521 852.769
R816 VGND.n1906 VGND.t2146 852.769
R817 VGND.n1936 VGND.t1404 852.769
R818 VGND.n1941 VGND.t2682 852.769
R819 VGND.n1946 VGND.t1537 852.769
R820 VGND.n1947 VGND.t1797 852.769
R821 VGND.t1952 VGND.n270 852.769
R822 VGND.n1384 VGND.t677 852.769
R823 VGND.n1385 VGND.t1637 852.769
R824 VGND.n1814 VGND.t647 852.769
R825 VGND.n1815 VGND.t1705 852.769
R826 VGND.n1840 VGND.t165 852.769
R827 VGND.n1841 VGND.t1451 852.769
R828 VGND.n1866 VGND.t1590 852.769
R829 VGND.n1867 VGND.t644 852.769
R830 VGND.n1892 VGND.t807 852.769
R831 VGND.n1893 VGND.t1631 852.769
R832 VGND.n1918 VGND.t106 852.769
R833 VGND.n1924 VGND.t422 852.769
R834 VGND.t1987 VGND.n1923 852.769
R835 VGND.n2361 VGND.t1267 852.769
R836 VGND.n2362 VGND.t329 852.769
R837 VGND.t2537 VGND.n271 852.769
R838 VGND.n1316 VGND.t845 852.769
R839 VGND.n1367 VGND.t582 852.769
R840 VGND.t2535 VGND.n1366 852.769
R841 VGND.t1803 VGND.n1361 852.769
R842 VGND.t81 VGND.n1356 852.769
R843 VGND.t267 VGND.n1351 852.769
R844 VGND.t1100 VGND.n1346 852.769
R845 VGND.t1988 VGND.n1341 852.769
R846 VGND.t1638 VGND.n1336 852.769
R847 VGND.t2555 VGND.n1331 852.769
R848 VGND.t1340 VGND.n1326 852.769
R849 VGND.t1402 VGND.n1321 852.769
R850 VGND.n1792 VGND.t2534 852.769
R851 VGND.t1632 VGND.n1791 852.769
R852 VGND.t1266 VGND.n1786 852.769
R853 VGND.t1616 VGND.n272 852.769
R854 VGND.n1521 VGND.t419 852.769
R855 VGND.n1526 VGND.t2507 852.769
R856 VGND.n1527 VGND.t2144 852.769
R857 VGND.n1653 VGND.t1279 852.769
R858 VGND.n1654 VGND.t1453 852.769
R859 VGND.n1679 VGND.t1524 852.769
R860 VGND.n1680 VGND.t176 852.769
R861 VGND.n1705 VGND.t1801 852.769
R862 VGND.n1706 VGND.t2153 852.769
R863 VGND.n1731 VGND.t1476 852.769
R864 VGND.n1732 VGND.t873 852.769
R865 VGND.n1762 VGND.t640 852.769
R866 VGND.n1767 VGND.t2409 852.769
R867 VGND.n1772 VGND.t2195 852.769
R868 VGND.n1773 VGND.t2187 852.769
R869 VGND.t2554 VGND.n273 852.769
R870 VGND.n1541 VGND.t71 852.769
R871 VGND.n1542 VGND.t1615 852.769
R872 VGND.n1640 VGND.t1301 852.769
R873 VGND.n1641 VGND.t80 852.769
R874 VGND.n1666 VGND.t1636 852.769
R875 VGND.n1667 VGND.t74 852.769
R876 VGND.n1692 VGND.t1791 852.769
R877 VGND.n1693 VGND.t1306 852.769
R878 VGND.n1718 VGND.t1154 852.769
R879 VGND.n1719 VGND.t1520 852.769
R880 VGND.n1744 VGND.t1954 852.769
R881 VGND.n1750 VGND.t1620 852.769
R882 VGND.t2154 VGND.n1749 852.769
R883 VGND.n2386 VGND.t808 852.769
R884 VGND.n2387 VGND.t1323 852.769
R885 VGND.t1305 VGND.n274 852.769
R886 VGND.n1299 VGND.t525 852.769
R887 VGND.n1554 VGND.t2649 852.769
R888 VGND.n1559 VGND.t889 852.769
R889 VGND.n1564 VGND.t1338 852.769
R890 VGND.n1569 VGND.t524 852.769
R891 VGND.n1574 VGND.t2321 852.769
R892 VGND.n1579 VGND.t1120 852.769
R893 VGND.n1584 VGND.t2295 852.769
R894 VGND.n1589 VGND.t1302 852.769
R895 VGND.n1594 VGND.t1523 852.769
R896 VGND.n1599 VGND.t1430 852.769
R897 VGND.n1604 VGND.t1136 852.769
R898 VGND.n1618 VGND.t84 852.769
R899 VGND.t879 VGND.n1617 852.769
R900 VGND.t2294 VGND.n1612 852.769
R901 VGND.t1951 VGND.n275 852.769
R902 VGND.n839 VGND.t1399 852.769
R903 VGND.n844 VGND.t2143 852.769
R904 VGND.n895 VGND.t77 852.769
R905 VGND.t388 VGND.n894 852.769
R906 VGND.t293 VGND.n889 852.769
R907 VGND.t2540 VGND.n884 852.769
R908 VGND.t141 VGND.n879 852.769
R909 VGND.t2644 VGND.n874 852.769
R910 VGND.t1290 VGND.n869 852.769
R911 VGND.t251 VGND.n864 852.769
R912 VGND.t523 VGND.n859 852.769
R913 VGND.t1536 VGND.n854 852.769
R914 VGND.t174 VGND.n849 852.769
R915 VGND.n2406 VGND.t87 852.769
R916 VGND.n2407 VGND.t1619 852.769
R917 VGND.t1137 VGND.n276 852.769
R918 VGND.t1704 VGND.n1293 852.769
R919 VGND.n724 VGND.t806 852.769
R920 VGND.n729 VGND.t1531 852.769
R921 VGND.n734 VGND.t177 852.769
R922 VGND.n739 VGND.t1450 852.769
R923 VGND.n744 VGND.t1454 852.769
R924 VGND.n749 VGND.t1099 852.769
R925 VGND.n754 VGND.t1304 852.769
R926 VGND.n759 VGND.t1802 852.769
R927 VGND.n764 VGND.t866 852.769
R928 VGND.n769 VGND.t2188 852.769
R929 VGND.n774 VGND.t2616 852.769
R930 VGND.n779 VGND.t1956 852.769
R931 VGND.n784 VGND.t268 852.769
R932 VGND.n785 VGND.t1788 852.769
R933 VGND.n2417 VGND.t1140 852.769
R934 VGND.n1511 VGND 851.341
R935 VGND.n2841 VGND.t2418 809.773
R936 VGND.n2840 VGND.t933 809.773
R937 VGND.t1008 VGND.n118 809.773
R938 VGND.n2836 VGND.t915 809.773
R939 VGND.t957 VGND.n181 809.773
R940 VGND.t1029 VGND.n639 809.773
R941 VGND.t909 VGND.n584 809.773
R942 VGND.n964 VGND.t951 809.773
R943 VGND.t963 VGND.n583 809.773
R944 VGND.n1515 VGND.t987 809.773
R945 VGND.t918 VGND.n1516 809.773
R946 VGND.n1297 VGND.t990 809.773
R947 VGND.t1020 VGND.n1298 809.773
R948 VGND.n1296 VGND.t960 809.773
R949 VGND.n1294 VGND.t719 809.773
R950 VGND.t430 VGND.t462 708.047
R951 VGND.t462 VGND.t315 708.047
R952 VGND.t315 VGND.t455 708.047
R953 VGND.t455 VGND.t1936 708.047
R954 VGND.t1936 VGND.t1555 708.047
R955 VGND.t1555 VGND.t1096 708.047
R956 VGND.t1096 VGND.t1558 708.047
R957 VGND.t1583 VGND.t1633 708.047
R958 VGND.t311 VGND.t495 708.047
R959 VGND.t495 VGND.t497 708.047
R960 VGND.t497 VGND.t321 708.047
R961 VGND.t321 VGND.t191 708.047
R962 VGND.t191 VGND.t188 708.047
R963 VGND.t188 VGND.t182 708.047
R964 VGND.t182 VGND.t185 708.047
R965 VGND.t545 VGND.t323 708.047
R966 VGND.t323 VGND.t543 708.047
R967 VGND.t543 VGND.t317 708.047
R968 VGND.t317 VGND.t264 708.047
R969 VGND.t264 VGND.t260 708.047
R970 VGND.t260 VGND.t254 708.047
R971 VGND.t254 VGND.t256 708.047
R972 VGND.t1580 VGND.t1634 708.047
R973 VGND.t551 VGND.t433 708.047
R974 VGND.t426 VGND.t551 708.047
R975 VGND.t1256 VGND.t426 708.047
R976 VGND.t1938 VGND.t1256 708.047
R977 VGND.t1557 VGND.t1938 708.047
R978 VGND.t1098 VGND.t1557 708.047
R979 VGND.t1554 VGND.t1098 708.047
R980 VGND.t453 VGND.t611 708.047
R981 VGND.t611 VGND.t428 708.047
R982 VGND.t428 VGND.t499 708.047
R983 VGND.t499 VGND.t187 708.047
R984 VGND.t187 VGND.t181 708.047
R985 VGND.t181 VGND.t190 708.047
R986 VGND.t190 VGND.t184 708.047
R987 VGND.t553 VGND.t424 708.047
R988 VGND.t424 VGND.t547 708.047
R989 VGND.t547 VGND.t319 708.047
R990 VGND.t319 VGND.t262 708.047
R991 VGND.t262 VGND.t258 708.047
R992 VGND.t258 VGND.t263 708.047
R993 VGND.t263 VGND.t259 708.047
R994 VGND.n2994 VGND.n2993 708.047
R995 VGND.t673 VGND.t2524 691.188
R996 VGND.t1372 VGND.t2646 691.188
R997 VGND.n2840 VGND.n2839 660.87
R998 VGND.t438 VGND.t217 657.471
R999 VGND.t447 VGND.t215 657.471
R1000 VGND.t592 VGND.t213 657.471
R1001 VGND.t2358 VGND.t620 657.471
R1002 VGND.t1263 VGND.t609 657.471
R1003 VGND.t613 VGND.t1751 657.471
R1004 VGND.t671 VGND.t1747 657.471
R1005 VGND.t493 VGND.t1741 657.471
R1006 VGND.t620 VGND.t622 654.197
R1007 VGND.t609 VGND.t1259 654.197
R1008 VGND.n966 VGND 640.614
R1009 VGND VGND.n117 640.614
R1010 VGND VGND.n2874 640.614
R1011 VGND VGND.n2907 640.614
R1012 VGND.n2910 VGND 632.184
R1013 VGND.t1643 VGND.t696 630.62
R1014 VGND.t2430 VGND.t2500 630.62
R1015 VGND.t2422 VGND.t2417 630.62
R1016 VGND.t1702 VGND.t758 630.62
R1017 VGND.t689 VGND.t2496 630.62
R1018 VGND.t760 VGND.t2478 630.62
R1019 VGND.t2464 VGND.t691 630.62
R1020 VGND.t1690 VGND.t685 630.62
R1021 VGND.t1686 VGND.t2466 630.62
R1022 VGND.t761 VGND.t2480 630.62
R1023 VGND.t741 VGND.t1688 630.62
R1024 VGND.t1678 VGND.t726 630.62
R1025 VGND.t2462 VGND.t2457 630.62
R1026 VGND.t730 VGND.t2450 630.62
R1027 VGND.t2434 VGND.t707 630.62
R1028 VGND.t1671 VGND.t2454 630.62
R1029 VGND.t1527 VGND.t2089 630.62
R1030 VGND.t1376 VGND.t1292 630.62
R1031 VGND.t157 VGND.t1477 630.62
R1032 VGND.t1385 VGND.t2095 630.62
R1033 VGND.t1990 VGND.t2087 630.62
R1034 VGND.t1541 VGND.t1487 630.62
R1035 VGND.t2662 VGND.t1485 630.62
R1036 VGND.t381 VGND.t2085 630.62
R1037 VGND.t285 VGND.t1380 630.62
R1038 VGND.t558 VGND.t1489 630.62
R1039 VGND.t1921 VGND.t2093 630.62
R1040 VGND.t167 VGND.t2091 630.62
R1041 VGND.t585 VGND.t1483 630.62
R1042 VGND.t1810 VGND.t1481 630.62
R1043 VGND.t1504 VGND.t1479 630.62
R1044 VGND.t1378 VGND.t1679 630.62
R1045 VGND.t1151 VGND.t2319 630.62
R1046 VGND.t2332 VGND.t2261 630.62
R1047 VGND.t1594 VGND.t93 630.62
R1048 VGND.t2517 VGND.t1592 630.62
R1049 VGND.t1707 VGND.t2317 630.62
R1050 VGND.t124 VGND.t2328 630.62
R1051 VGND.t1308 VGND.t2326 630.62
R1052 VGND.t1758 VGND.t2315 630.62
R1053 VGND.t474 VGND.t2313 630.62
R1054 VGND.t32 VGND.t2330 630.62
R1055 VGND.t1440 VGND.t2075 630.62
R1056 VGND.t2593 VGND.t2073 630.62
R1057 VGND.t308 VGND.t2324 630.62
R1058 VGND.t113 VGND.t2322 630.62
R1059 VGND.t2118 VGND.t1596 630.62
R1060 VGND.t745 VGND.t2311 630.62
R1061 VGND.t1284 VGND.t1925 630.62
R1062 VGND.t1298 VGND.t1625 630.62
R1063 VGND.t147 VGND.t1608 630.62
R1064 VGND.t1606 VGND.t1391 630.62
R1065 VGND.t2081 VGND.t1282 630.62
R1066 VGND.t2003 VGND.t1543 630.62
R1067 VGND.t2668 VGND.t2001 630.62
R1068 VGND.t1280 VGND.t387 630.62
R1069 VGND.t1155 VGND.t1629 630.62
R1070 VGND.t1623 VGND.t568 630.62
R1071 VGND.t766 VGND.t1288 630.62
R1072 VGND.t1286 VGND.t1107 630.62
R1073 VGND.t591 VGND.t1999 630.62
R1074 VGND.t1034 VGND.t1864 630.62
R1075 VGND.t1510 VGND.t1610 630.62
R1076 VGND.t1627 VGND.t1700 630.62
R1077 VGND.t1116 VGND.t273 630.62
R1078 VGND.t833 VGND.t2217 630.62
R1079 VGND.t1434 VGND.t799 630.62
R1080 VGND.t60 VGND.t1432 630.62
R1081 VGND.t271 VGND.t2243 630.62
R1082 VGND.t1901 VGND.t2213 630.62
R1083 VGND.t2211 VGND.t2655 630.62
R1084 VGND.t862 VGND.t269 630.62
R1085 VGND.t2559 VGND.t884 630.62
R1086 VGND.t528 VGND.t2215 630.62
R1087 VGND.t277 VGND.t2528 630.62
R1088 VGND.t1975 VGND.t275 630.62
R1089 VGND.t2209 VGND.t2200 630.62
R1090 VGND.t2207 VGND.t1819 630.62
R1091 VGND.t2125 VGND.t1436 630.62
R1092 VGND.t2557 VGND.t2495 630.62
R1093 VGND.t1145 VGND.t2603 630.62
R1094 VGND.t2255 VGND.t2105 630.62
R1095 VGND.t2249 VGND.t128 630.62
R1096 VGND.t1548 VGND.t2511 630.62
R1097 VGND.t2601 VGND.t1964 630.62
R1098 VGND.t2101 VGND.t2544 630.62
R1099 VGND.t2099 VGND.t2404 630.62
R1100 VGND.t2599 VGND.t1740 630.62
R1101 VGND.t2597 VGND.t468 630.62
R1102 VGND.t2103 VGND.t539 630.62
R1103 VGND.t1546 VGND.t2566 630.62
R1104 VGND.t1544 VGND.t2608 630.62
R1105 VGND.t2097 VGND.t302 630.62
R1106 VGND.t2253 VGND.t1808 630.62
R1107 VGND.t2251 VGND.t2112 630.62
R1108 VGND.t2107 VGND.t717 630.62
R1109 VGND.t2266 VGND.t1526 630.62
R1110 VGND.t1291 VGND.t1568 630.62
R1111 VGND.t146 VGND.t2280 630.62
R1112 VGND.t2272 VGND.t1384 630.62
R1113 VGND.t1989 VGND.t2264 630.62
R1114 VGND.t2290 VGND.t1540 630.62
R1115 VGND.t2661 VGND.t2288 630.62
R1116 VGND.t2262 VGND.t380 630.62
R1117 VGND.t284 VGND.t1572 630.62
R1118 VGND.t2292 VGND.t557 630.62
R1119 VGND.t1920 VGND.t2270 630.62
R1120 VGND.t2268 VGND.t166 630.62
R1121 VGND.t584 VGND.t2286 630.62
R1122 VGND.t2041 VGND.t2284 630.62
R1123 VGND.t1503 VGND.t2282 630.62
R1124 VGND.t1570 VGND.t1677 630.62
R1125 VGND.t1930 VGND.t480 630.62
R1126 VGND.t2163 VGND.t631 630.62
R1127 VGND.t488 VGND.t125 630.62
R1128 VGND.t1161 VGND.t486 630.62
R1129 VGND.t478 VGND.t2082 630.62
R1130 VGND.t2550 VGND.t627 630.62
R1131 VGND.t625 VGND.t2398 630.62
R1132 VGND.t1067 VGND.t476 630.62
R1133 VGND.t635 VGND.t1156 630.62
R1134 VGND.t569 VGND.t629 630.62
R1135 VGND.t484 VGND.t767 630.62
R1136 VGND.t1108 VGND.t482 630.62
R1137 VGND.t652 VGND.t1792 630.62
R1138 VGND.t637 VGND.t1035 630.62
R1139 VGND.t1511 VGND.t490 630.62
R1140 VGND.t633 VGND.t1703 630.62
R1141 VGND.t1271 VGND.t1117 630.62
R1142 VGND.t1961 VGND.t834 630.62
R1143 VGND.t818 VGND.t802 630.62
R1144 VGND.t816 VGND.t61 630.62
R1145 VGND.t2139 VGND.t2244 630.62
R1146 VGND.t1040 VGND.t1902 630.62
R1147 VGND.t1038 VGND.t2656 630.62
R1148 VGND.t2137 VGND.t863 630.62
R1149 VGND.t2135 VGND.t885 630.62
R1150 VGND.t1959 VGND.t529 630.62
R1151 VGND.t1275 VGND.t2529 630.62
R1152 VGND.t1273 VGND.t1976 630.62
R1153 VGND.t1036 VGND.t2201 630.62
R1154 VGND.t822 VGND.t1820 630.62
R1155 VGND.t820 VGND.t2126 630.62
R1156 VGND.t2133 VGND.t2497 630.62
R1157 VGND.t1114 VGND.t2161 630.62
R1158 VGND.t832 VGND.t2037 630.62
R1159 VGND.t801 VGND.t2396 630.62
R1160 VGND.t2394 VGND.t59 630.62
R1161 VGND.t650 VGND.t2159 630.62
R1162 VGND.t2033 VGND.t1566 630.62
R1163 VGND.t668 VGND.t2031 630.62
R1164 VGND.t2157 VGND.t861 630.62
R1165 VGND.t883 VGND.t2155 630.62
R1166 VGND.t2035 VGND.t527 630.62
R1167 VGND.t2527 VGND.t2392 630.62
R1168 VGND.t2390 VGND.t1974 630.62
R1169 VGND.t2199 VGND.t2029 630.62
R1170 VGND.t1830 VGND.t1576 630.62
R1171 VGND.t2123 VGND.t1574 630.62
R1172 VGND.t867 VGND.t2488 630.62
R1173 VGND.t1452 VGND.t1785 630.62
R1174 VGND.t1605 VGND.t1775 630.62
R1175 VGND.t1872 VGND.t131 630.62
R1176 VGND.t2510 VGND.t1870 630.62
R1177 VGND.t1783 VGND.t1963 630.62
R1178 VGND.t2543 VGND.t1474 630.62
R1179 VGND.t1472 VGND.t2403 630.62
R1180 VGND.t1739 VGND.t1781 630.62
R1181 VGND.t1779 VGND.t2168 630.62
R1182 VGND.t536 VGND.t1773 630.62
R1183 VGND.t1868 VGND.t2565 630.62
R1184 VGND.t1861 VGND.t1866 630.62
R1185 VGND.t1470 VGND.t301 630.62
R1186 VGND.t1468 VGND.t1805 630.62
R1187 VGND.t2111 VGND.t1466 630.62
R1188 VGND.t1777 VGND.t712 630.62
R1189 VGND.t825 VGND.t511 630.62
R1190 VGND.t2677 VGND.t574 630.62
R1191 VGND.t2574 VGND.t769 630.62
R1192 VGND.t2572 VGND.t603 630.62
R1193 VGND.t509 VGND.t2150 630.62
R1194 VGND.t570 VGND.t164 630.62
R1195 VGND.t2582 VGND.t662 630.62
R1196 VGND.t580 VGND.t2684 630.62
R1197 VGND.t578 VGND.t1131 630.62
R1198 VGND.t572 VGND.t522 630.62
R1199 VGND.t2570 VGND.t2042 630.62
R1200 VGND.t2568 VGND.t1834 630.62
R1201 VGND.t2580 VGND.t403 630.62
R1202 VGND.t2578 VGND.t1828 630.62
R1203 VGND.t2576 VGND.t73 630.62
R1204 VGND.t576 VGND.t2447 630.62
R1205 VGND.t1528 VGND.t858 630.62
R1206 VGND.t1293 VGND.t848 630.62
R1207 VGND.t148 VGND.t1497 630.62
R1208 VGND.t1495 VGND.t1390 630.62
R1209 VGND.t1991 VGND.t856 630.62
R1210 VGND.t658 VGND.t1542 630.62
R1211 VGND.t2663 VGND.t656 630.62
R1212 VGND.t854 VGND.t382 630.62
R1213 VGND.t1460 VGND.t852 630.62
R1214 VGND.t660 VGND.t567 630.62
R1215 VGND.t1922 VGND.t1493 630.62
R1216 VGND.t1491 VGND.t1106 630.62
R1217 VGND.t586 VGND.t654 630.62
R1218 VGND.t1033 VGND.t295 630.62
R1219 VGND.t1509 VGND.t1499 630.62
R1220 VGND.t850 VGND.t1697 630.62
R1221 VGND.t2669 VGND.t824 630.62
R1222 VGND.t2676 VGND.t336 630.62
R1223 VGND.t1761 VGND.t772 630.62
R1224 VGND.t602 VGND.t1759 630.62
R1225 VGND.t1552 VGND.t2149 630.62
R1226 VGND.t163 VGND.t332 630.62
R1227 VGND.t330 VGND.t1320 630.62
R1228 VGND.t370 VGND.t1550 630.62
R1229 VGND.t340 VGND.t1130 630.62
R1230 VGND.t519 VGND.t334 630.62
R1231 VGND.t2673 VGND.t878 630.62
R1232 VGND.t1831 VGND.t2671 630.62
R1233 VGND.t1767 VGND.t402 630.62
R1234 VGND.t1765 VGND.t1825 630.62
R1235 VGND.t72 VGND.t1763 630.62
R1236 VGND.t338 VGND.t2444 630.62
R1237 VGND.t1150 VGND.t1945 630.62
R1238 VGND.t2306 VGND.t2260 630.62
R1239 VGND.t811 VGND.t297 630.62
R1240 VGND.t2516 VGND.t1382 630.62
R1241 VGND.t1706 VGND.t1943 630.62
R1242 VGND.t2545 VGND.t2302 630.62
R1243 VGND.t1307 VGND.t2300 630.62
R1244 VGND.t1757 VGND.t1941 630.62
R1245 VGND.t473 VGND.t1939 630.62
R1246 VGND.t540 VGND.t2304 630.62
R1247 VGND.t2567 VGND.t1949 630.62
R1248 VGND.t2609 VGND.t1947 630.62
R1249 VGND.t307 VGND.t2298 630.62
R1250 VGND.t2296 VGND.t1809 630.62
R1251 VGND.t299 VGND.t2117 630.62
R1252 VGND.t2308 VGND.t732 630.62
R1253 VGND.t1115 VGND.t194 630.62
R1254 VGND.t831 VGND.t2177 630.62
R1255 VGND.t800 VGND.t2189 630.62
R1256 VGND.t200 VGND.t1196 630.62
R1257 VGND.t2183 VGND.t651 630.62
R1258 VGND.t2173 VGND.t1567 630.62
R1259 VGND.t2171 VGND.t667 630.62
R1260 VGND.t2181 VGND.t860 630.62
R1261 VGND.t2179 VGND.t882 630.62
R1262 VGND.t2175 VGND.t526 630.62
R1263 VGND.t198 VGND.t2526 630.62
R1264 VGND.t196 VGND.t1973 630.62
R1265 VGND.t2169 VGND.t2198 630.62
R1266 VGND.t2193 VGND.t1829 630.62
R1267 VGND.t2124 VGND.t2191 630.62
R1268 VGND.t809 VGND.t2487 630.62
R1269 VGND.t1665 VGND.t1347 630.62
R1270 VGND.t1998 VGND.t2445 630.62
R1271 VGND.t768 VGND.t722 630.62
R1272 VGND.t599 VGND.t700 630.62
R1273 VGND.t1714 VGND.t1654 630.62
R1274 VGND.t140 VGND.t2426 630.62
R1275 VGND.t1315 VGND.t2415 630.62
R1276 VGND.t379 VGND.t1650 630.62
R1277 VGND.t122 VGND.t2493 630.62
R1278 VGND.t33 VGND.t2428 630.62
R1279 VGND.t1449 VGND.t687 630.62
R1280 VGND.t2594 VGND.t1698 630.62
R1281 VGND.t397 VGND.t2410 630.62
R1282 VGND.t847 VGND.t753 630.62
R1283 VGND.t90 VGND.t728 630.62
R1284 VGND.t2472 VGND.t757 630.62
R1285 VGND.n994 VGND.n966 599.125
R1286 VGND.n117 VGND.n116 599.125
R1287 VGND.n2874 VGND.n2873 599.125
R1288 VGND.n2907 VGND.n2906 599.125
R1289 VGND.n2911 VGND.n2910 599.125
R1290 VGND.n2922 VGND.n2921 599.125
R1291 VGND.n2994 VGND.n2992 599.125
R1292 VGND.n2961 VGND.n2960 599.125
R1293 VGND.t1251 VGND 581.61
R1294 VGND.t1558 VGND 573.181
R1295 VGND.t185 VGND 573.181
R1296 VGND.t256 VGND 573.181
R1297 VGND VGND.t1743 573.181
R1298 VGND.t1374 VGND 564.751
R1299 VGND.n3012 VGND 564.751
R1300 VGND.n3011 VGND 564.751
R1301 VGND.n3010 VGND 556.322
R1302 VGND VGND.t1329 539.465
R1303 VGND.t280 VGND 539.465
R1304 VGND.t410 VGND.n582 494.779
R1305 VGND.n2838 VGND.n7 494.253
R1306 VGND.n1126 VGND.t749 492.058
R1307 VGND.t1693 VGND.n1135 492.058
R1308 VGND.n1136 VGND.t1669 492.058
R1309 VGND.t747 VGND.n1148 492.058
R1310 VGND.n1149 VGND.t735 492.058
R1311 VGND.t713 VGND.n1167 492.058
R1312 VGND.n1168 VGND.t2458 492.058
R1313 VGND.t2438 VGND.n1180 492.058
R1314 VGND.n1181 VGND.t708 492.058
R1315 VGND.t1652 VGND.n1199 492.058
R1316 VGND.n1200 VGND.t2502 492.058
R1317 VGND.t2413 VGND.n1212 492.058
R1318 VGND.n1213 VGND.t698 492.058
R1319 VGND.t2491 VGND.n1231 492.058
R1320 VGND.n1232 VGND.t2424 492.058
R1321 VGND.t622 VGND.t406 481.877
R1322 VGND.t406 VGND.t2274 481.877
R1323 VGND.t313 VGND.t460 481.877
R1324 VGND.t1259 VGND.t313 481.877
R1325 VGND.t642 VGND 452.382
R1326 VGND.n1126 VGND.t1113 424.312
R1327 VGND.n1135 VGND.t1516 424.312
R1328 VGND.n1136 VGND.t1876 424.312
R1329 VGND.n1148 VGND.t1787 424.312
R1330 VGND.n1149 VGND.t2536 424.312
R1331 VGND.n1167 VGND.t1622 424.312
R1332 VGND.n1168 VGND.t2 424.312
R1333 VGND.n1180 VGND.t1325 424.312
R1334 VGND.n1181 VGND.t1534 424.312
R1335 VGND.n1199 VGND.t2521 424.312
R1336 VGND.n1200 VGND.t846 424.312
R1337 VGND.n1212 VGND.t0 424.312
R1338 VGND.n1213 VGND.t1303 424.312
R1339 VGND.n1231 VGND.t2606 424.312
R1340 VGND.n1232 VGND.t887 424.312
R1341 VGND.t1612 VGND.n277 424.312
R1342 VGND.t286 VGND 419.68
R1343 VGND.n639 VGND.n151 413.043
R1344 VGND.t945 VGND.t2418 408.469
R1345 VGND.t894 VGND.t694 408.469
R1346 VGND.t2498 VGND.t900 408.469
R1347 VGND.t906 VGND.t2476 408.469
R1348 VGND.t692 VGND.t993 408.469
R1349 VGND.t999 VGND.t681 408.469
R1350 VGND.t1684 VGND.t912 408.469
R1351 VGND.t954 VGND.t762 408.469
R1352 VGND.t739 VGND.t969 408.469
R1353 VGND.t1005 VGND.t1680 408.469
R1354 VGND.t2460 VGND.t927 408.469
R1355 VGND.t972 VGND.t2448 408.469
R1356 VGND.t710 VGND.t1011 408.469
R1357 VGND.t1023 VGND.t1667 408.469
R1358 VGND.t2436 VGND.t939 408.469
R1359 VGND.t724 VGND.t981 408.469
R1360 VGND.t15 VGND.t933 408.469
R1361 VGND.t1148 VGND.t785 408.469
R1362 VGND.t1887 VGND.t2258 408.469
R1363 VGND.t2051 VGND.t129 408.469
R1364 VGND.t1723 VGND.t1388 408.469
R1365 VGND.t1088 VGND.t1967 408.469
R1366 VGND.t2356 VGND.t161 408.469
R1367 VGND.t2378 VGND.t2407 408.469
R1368 VGND.t2021 VGND.t1755 408.469
R1369 VGND.t1236 VGND.t471 408.469
R1370 VGND.t1413 VGND.t537 408.469
R1371 VGND.t2009 VGND.t876 408.469
R1372 VGND.t1228 VGND.t1862 408.469
R1373 VGND.t1222 VGND.t305 408.469
R1374 VGND.t1352 VGND.t1806 408.469
R1375 VGND.t1507 VGND.t346 408.469
R1376 VGND.t1849 VGND.t1008 408.469
R1377 VGND.t828 VGND.t1370 408.469
R1378 VGND.t2680 VGND.t46 408.469
R1379 VGND.t2386 VGND.t770 408.469
R1380 VGND.t787 VGND.t600 408.469
R1381 VGND.t2071 VGND.t648 408.469
R1382 VGND.t2382 VGND.t1538 408.469
R1383 VGND.t1725 VGND.t665 408.469
R1384 VGND.t1090 VGND.t2687 408.469
R1385 VGND.t2049 VGND.t1134 408.469
R1386 VGND.t1178 VGND.t520 408.469
R1387 VGND.t1076 VGND.t1918 408.469
R1388 VGND.t2348 VGND.t1832 408.469
R1389 VGND.t1417 VGND.t2196 408.469
R1390 VGND.t348 VGND.t1826 408.469
R1391 VGND.t1230 VGND.t91 408.469
R1392 VGND.t915 VGND.t2019 408.469
R1393 VGND.t2340 VGND.t1343 408.469
R1394 VGND.t1409 VGND.t1994 408.469
R1395 VGND.t96 VGND.t1360 408.469
R1396 VGND.t1061 VGND.t1164 408.469
R1397 VGND.t1710 VGND.t1204 408.469
R1398 VGND.t1348 VGND.t1562 408.469
R1399 VGND.t1311 VGND.t2640 408.469
R1400 VGND.t1737 VGND.t375 408.469
R1401 VGND.t118 VGND.t1899 408.469
R1402 VGND.t19 VGND.t28 408.469
R1403 VGND.t2045 VGND.t1731 408.469
R1404 VGND.t1891 VGND.t2612 408.469
R1405 VGND.t1985 VGND.t393 408.469
R1406 VGND.t1186 VGND.t109 408.469
R1407 VGND.t1514 VGND.t242 408.469
R1408 VGND.t1084 VGND.t957 408.469
R1409 VGND.t2370 VGND.t1931 408.469
R1410 VGND.t2164 VGND.t1172 408.469
R1411 VGND.t354 VGND.t151 408.469
R1412 VGND.t66 VGND.t2342 408.469
R1413 VGND.t2231 VGND.t2083 408.469
R1414 VGND.t136 VGND.t2642 408.469
R1415 VGND.t1063 VGND.t2399 408.469
R1416 VGND.t1068 VGND.t1206 408.469
R1417 VGND.t1350 VGND.t1157 408.469
R1418 VGND.t563 VGND.t1853 408.469
R1419 VGND.t795 VGND.t1445 408.469
R1420 VGND.t172 VGND.t52 408.469
R1421 VGND.t1793 VGND.t23 408.469
R1422 VGND.t244 VGND.t1815 408.469
R1423 VGND.t2131 VGND.t1895 408.469
R1424 VGND.t2065 VGND.t1029 408.469
R1425 VGND.t1717 VGND.t466 408.469
R1426 VGND.t837 VGND.t230 408.469
R1427 VGND.t812 VGND.t1240 408.469
R1428 VGND.t2514 VGND.t2372 408.469
R1429 VGND.t2147 VGND.t2015 408.469
R1430 VGND.t1905 VGND.t1065 408.469
R1431 VGND.t1318 VGND.t2344 408.469
R1432 VGND.t368 VGND.t2235 408.469
R1433 VGND.t841 VGND.t342 408.469
R1434 VGND.t515 VGND.t1220 408.469
R1435 VGND.t2532 VGND.t2223 408.469
R1436 VGND.t2589 VGND.t2638 408.469
R1437 VGND.t400 VGND.t1855 408.469
R1438 VGND.t1111 VGND.t1897 408.469
R1439 VGND.t2115 VGND.t56 408.469
R1440 VGND.t936 VGND.t5 408.469
R1441 VGND.t777 VGND.t1146 408.469
R1442 VGND.t1877 VGND.t2256 408.469
R1443 VGND.t126 VGND.t2350 408.469
R1444 VGND.t248 VGND.t1386 408.469
R1445 VGND.t1965 VGND.t1246 408.469
R1446 VGND.t2336 VGND.t159 408.469
R1447 VGND.t2405 VGND.t2366 408.469
R1448 VGND.t364 VGND.t1753 408.469
R1449 VGND.t469 VGND.t1057 408.469
R1450 VGND.t2239 VGND.t534 408.469
R1451 VGND.t874 VGND.t358 408.469
R1452 VGND.t1053 VGND.t1859 408.469
R1453 VGND.t1214 VGND.t303 408.469
R1454 VGND.t50 VGND.t1817 408.469
R1455 VGND.t1505 VGND.t2632 408.469
R1456 VGND.t1839 VGND.t909 408.469
R1457 VGND.t1358 VGND.t1345 408.469
R1458 VGND.t1996 VGND.t34 408.469
R1459 VGND.t2376 VGND.t94 408.469
R1460 VGND.t1166 VGND.t779 408.469
R1461 VGND.t2057 VGND.t1712 408.469
R1462 VGND.t1564 VGND.t2368 408.469
R1463 VGND.t1715 VGND.t1313 408.469
R1464 VGND.t377 VGND.t1074 408.469
R1465 VGND.t2338 VGND.t120 408.469
R1466 VGND.t30 VGND.t2027 408.469
R1467 VGND.t1242 VGND.t2047 408.469
R1468 VGND.t2614 VGND.t2334 408.469
R1469 VGND.t395 VGND.t2241 408.469
R1470 VGND.t2634 VGND.t111 408.469
R1471 VGND.t2109 VGND.t1055 408.469
R1472 VGND.t951 VGND.t362 408.469
R1473 VGND.t1933 VGND.t1423 408.469
R1474 VGND.t2166 VGND.t2237 408.469
R1475 VGND.t149 VGND.t54 408.469
R1476 VGND.t68 VGND.t1045 408.469
R1477 VGND.t1603 VGND.t791 408.469
R1478 VGND.t138 VGND.t40 408.469
R1479 VGND.t2401 VGND.t2626 408.469
R1480 VGND.t1070 VGND.t1729 408.469
R1481 VGND.t1159 VGND.t1885 408.469
R1482 VGND.t565 VGND.t11 408.469
R1483 VGND.t1447 VGND.t1719 408.469
R1484 VGND.t1104 VGND.t1879 408.469
R1485 VGND.t1795 VGND.t2069 408.469
R1486 VGND.t1031 VGND.t1174 408.469
R1487 VGND.t1501 VGND.t232 408.469
R1488 VGND.t1244 VGND.t963 408.469
R1489 VGND.t1188 VGND.t1926 408.469
R1490 VGND.t2025 VGND.t1294 408.469
R1491 VGND.t155 VGND.t2636 408.469
R1492 VGND.t1425 VGND.t62 408.469
R1493 VGND.t2077 VGND.t2219 408.469
R1494 VGND.t2628 VGND.t134 408.469
R1495 VGND.t2666 VGND.t1047 408.469
R1496 VGND.t793 VGND.t385 408.469
R1497 VGND.t1463 VGND.t44 408.469
R1498 VGND.t1843 VGND.t561 408.469
R1499 VGND.t1443 VGND.t783 408.469
R1500 VGND.t36 VGND.t170 408.469
R1501 VGND.t13 VGND.t589 408.469
R1502 VGND.t234 VGND.t1811 408.469
R1503 VGND.t2129 VGND.t1881 408.469
R1504 VGND.t2055 VGND.t891 408.469
R1505 VGND.t246 VGND.t464 408.469
R1506 VGND.t835 VGND.t228 408.469
R1507 VGND.t1059 VGND.t814 408.469
R1508 VGND.t2512 VGND.t1190 408.469
R1509 VGND.t360 VGND.t282 408.469
R1510 VGND.t1903 VGND.t1049 408.469
R1511 VGND.t1427 VGND.t1316 408.469
R1512 VGND.t366 VGND.t2221 408.469
R1513 VGND.t2630 VGND.t839 408.469
R1514 VGND.t513 VGND.t1212 408.469
R1515 VGND.t1366 VGND.t2530 408.469
R1516 VGND.t2595 VGND.t2624 408.469
R1517 VGND.t398 VGND.t1845 408.469
R1518 VGND.t1883 VGND.t1109 408.469
R1519 VGND.t2113 VGND.t38 408.469
R1520 VGND.t1847 VGND.t987 408.469
R1521 VGND.t1364 VGND.t1123 408.469
R1522 VGND.t1971 VGND.t42 408.469
R1523 VGND.t142 VGND.t2384 408.469
R1524 VGND.t1194 VGND.t781 408.469
R1525 VGND.t2247 VGND.t2067 408.469
R1526 VGND.t2541 VGND.t2374 408.469
R1527 VGND.t2659 VGND.t1721 408.469
R1528 VGND.t391 VGND.t1086 408.469
R1529 VGND.t1458 VGND.t2352 408.469
R1530 VGND.t532 VGND.t1176 408.469
R1531 VGND.t2563 VGND.t1248 408.469
R1532 VGND.t2548 VGND.t2346 408.469
R1533 VGND.t2204 VGND.t1411 408.469
R1534 VGND.t2039 VGND.t344 408.469
R1535 VGND.t2121 VGND.t1226 408.469
R1536 VGND.t2053 VGND.t918 408.469
R1537 VGND.t238 VGND.t1341 408.469
R1538 VGND.t1094 VGND.t1992 408.469
R1539 VGND.t98 VGND.t1051 408.469
R1540 VGND.t1184 VGND.t1162 408.469
R1541 VGND.t1708 VGND.t356 408.469
R1542 VGND.t1043 VGND.t1560 408.469
R1543 VGND.t1309 VGND.t1421 408.469
R1544 VGND.t1368 VGND.t373 408.469
R1545 VGND.t116 VGND.t2622 408.469
R1546 VGND.t1208 VGND.t541 408.469
R1547 VGND.t2043 VGND.t1362 408.469
R1548 VGND.t2620 VGND.t2610 408.469
R1549 VGND.t1835 VGND.t309 408.469
R1550 VGND.t1200 VGND.t107 408.469
R1551 VGND.t1512 VGND.t25 408.469
R1552 VGND.t990 VGND.t240 408.469
R1553 VGND.t3 VGND.t1121 408.469
R1554 VGND.t1969 VGND.t2380 408.469
R1555 VGND.t2023 VGND.t144 408.469
R1556 VGND.t1192 VGND.t2059 408.469
R1557 VGND.t1415 VGND.t2245 408.469
R1558 VGND.t2551 VGND.t2013 408.469
R1559 VGND.t1078 VGND.t2657 408.469
R1560 VGND.t389 VGND.t1224 408.469
R1561 VGND.t2233 VGND.t1456 408.469
R1562 VGND.t530 VGND.t350 408.469
R1563 VGND.t1216 VGND.t2561 408.469
R1564 VGND.t2546 VGND.t2225 408.469
R1565 VGND.t2202 VGND.t1356 408.469
R1566 VGND.t1733 VGND.t1821 408.469
R1567 VGND.t2119 VGND.t797 408.469
R1568 VGND.t1889 VGND.t1020 408.469
R1569 VGND.t826 VGND.t1837 408.469
R1570 VGND.t1727 VGND.t2678 408.469
R1571 VGND.t1092 VGND.t773 408.469
R1572 VGND.t7 VGND.t2518 408.469
R1573 VGND.t1180 VGND.t2151 408.469
R1574 VGND.t1080 VGND.t1907 408.469
R1575 VGND.t2061 VGND.t663 408.469
R1576 VGND.t1419 VGND.t2685 408.469
R1577 VGND.t2017 VGND.t1132 408.469
R1578 VGND.t1232 VGND.t517 408.469
R1579 VGND.t1407 VGND.t1916 408.469
R1580 VGND.t2005 VGND.t2591 408.469
R1581 VGND.t404 VGND.t352 408.469
R1582 VGND.t1823 VGND.t1202 408.469
R1583 VGND.t88 VGND.t2227 408.469
R1584 VGND.t48 VGND.t960 408.469
R1585 VGND.t1210 VGND.t1928 408.469
R1586 VGND.t789 VGND.t1296 408.469
R1587 VGND.t153 VGND.t1981 408.469
R1588 VGND.t64 VGND.t1841 408.469
R1589 VGND.t2079 VGND.t236 408.469
R1590 VGND.t132 VGND.t2063 408.469
R1591 VGND.t2664 VGND.t9 408.469
R1592 VGND.t383 VGND.t1182 408.469
R1593 VGND.t1461 VGND.t1082 408.469
R1594 VGND.t559 VGND.t2354 408.469
R1595 VGND.t1441 VGND.t1170 408.469
R1596 VGND.t168 VGND.t1072 408.469
R1597 VGND.t587 VGND.t1234 408.469
R1598 VGND.t2229 VGND.t1813 408.469
R1599 VGND.t2127 VGND.t2007 408.469
R1600 VGND.t719 VGND.t1238 408.469
R1601 VGND.t1168 VGND.t1663 408.469
R1602 VGND.t2011 VGND.t2442 408.469
R1603 VGND.t1857 VGND.t2420 408.469
R1604 VGND.t1405 VGND.t1658 408.469
R1605 VGND.t1354 VGND.t1647 408.469
R1606 VGND.t1851 VGND.t2489 408.469
R1607 VGND.t1218 VGND.t704 408.469
R1608 VGND.t775 VGND.t683 408.469
R1609 VGND.t21 VGND.t2485 408.469
R1610 VGND.t1735 VGND.t764 408.469
R1611 VGND.t1893 VGND.t751 408.469
R1612 VGND.t17 VGND.t1682 408.469
R1613 VGND.t2388 VGND.t2468 408.469
R1614 VGND.t226 VGND.t733 408.469
R1615 VGND.t1691 VGND.t1983 408.469
R1616 VGND.t1261 VGND.t2586 397.848
R1617 VGND.t2586 VGND.t458 397.848
R1618 VGND.t458 VGND.t451 397.848
R1619 VGND.t451 VGND.t1745 397.848
R1620 VGND.t1745 VGND.t1746 397.848
R1621 VGND.t1746 VGND.t1749 397.848
R1622 VGND.t1749 VGND.t1750 397.848
R1623 VGND.t1578 VGND.t2645 396.17
R1624 VGND.t202 VGND.t2185 396.17
R1625 VGND.n2997 VGND.n37 394.137
R1626 VGND.n2999 VGND.n2998 394.137
R1627 VGND.n2493 VGND.n36 394.137
R1628 VGND.n2432 VGND.n2431 394.137
R1629 VGND.n2430 VGND.n265 394.137
R1630 VGND.n2429 VGND.n266 394.137
R1631 VGND.n2428 VGND.n267 394.137
R1632 VGND.n2427 VGND.n268 394.137
R1633 VGND.n2426 VGND.n269 394.137
R1634 VGND.n2425 VGND.n270 394.137
R1635 VGND.n2424 VGND.n271 394.137
R1636 VGND.n2423 VGND.n272 394.137
R1637 VGND.n2422 VGND.n273 394.137
R1638 VGND.n2421 VGND.n274 394.137
R1639 VGND.n2420 VGND.n275 394.137
R1640 VGND.n2419 VGND.n276 394.137
R1641 VGND.n2418 VGND.n2417 394.137
R1642 VGND.n151 VGND.t326 387.421
R1643 VGND.n1510 VGND.t1333 387.421
R1644 VGND.n1512 VGND.t207 387.421
R1645 VGND.n1514 VGND.t328 387.421
R1646 VGND.n2837 VGND.t204 387.421
R1647 VGND.t1912 VGND.t1529 362.452
R1648 VGND.t1529 VGND.t280 345.594
R1649 VGND VGND.t100 328.616
R1650 VGND VGND.t287 328.616
R1651 VGND.t325 VGND 328.616
R1652 VGND.t103 VGND 328.616
R1653 VGND VGND.t413 328.616
R1654 VGND.t1701 VGND.t755 313.776
R1655 VGND.t1695 VGND.t2482 313.776
R1656 VGND.t2467 VGND.t2474 313.776
R1657 VGND.t2452 VGND.t731 313.776
R1658 VGND.t1689 VGND.t743 313.776
R1659 VGND.t1673 VGND.t2455 313.776
R1660 VGND.t746 VGND.t1660 313.776
R1661 VGND.t737 VGND.t721 313.776
R1662 VGND.t1662 VGND.t715 313.776
R1663 VGND.t1675 VGND.t2456 313.776
R1664 VGND.t718 VGND.t2440 313.776
R1665 VGND.t2431 VGND.t706 313.776
R1666 VGND.t1649 VGND.t1656 313.776
R1667 VGND.t1644 VGND.t2433 313.776
R1668 VGND.t2412 VGND.t2483 313.776
R1669 VGND.t702 VGND.t1646 313.776
R1670 VGND.t1587 VGND.t1578 311.877
R1671 VGND.t2185 VGND.t1251 311.877
R1672 VGND VGND.t1583 303.449
R1673 VGND VGND.t1587 295.019
R1674 VGND.n74 VGND.t461 287.832
R1675 VGND VGND.t220 286.591
R1676 VGND.n968 VGND.t439 282.327
R1677 VGND.n66 VGND.t494 282.327
R1678 VGND.n973 VGND.t2359 281.13
R1679 VGND.n77 VGND.t1264 281.13
R1680 VGND.n130 VGND.t2360 280.978
R1681 VGND.n130 VGND.t598 280.978
R1682 VGND.n598 VGND.t444 280.978
R1683 VGND.n598 VGND.t1601 280.978
R1684 VGND.n978 VGND.t2275 280.978
R1685 VGND.n160 VGND.t618 280.978
R1686 VGND.n160 VGND.t436 280.978
R1687 VGND.n100 VGND.t431 280.978
R1688 VGND.n100 VGND.t556 280.978
R1689 VGND.n2855 VGND.t312 280.978
R1690 VGND.n2855 VGND.t1254 280.978
R1691 VGND.n2887 VGND.t546 280.978
R1692 VGND.n2887 VGND.t670 280.978
R1693 VGND.t675 VGND 278.161
R1694 VGND.n2993 VGND 271.014
R1695 VGND VGND.t1580 252.875
R1696 VGND VGND.t1585 252.875
R1697 VGND.t433 VGND 252.875
R1698 VGND VGND.t453 252.875
R1699 VGND VGND.t553 252.875
R1700 VGND.n3027 VGND.n3026 244.329
R1701 VGND.n3024 VGND.n3023 244.329
R1702 VGND.n3030 VGND.n4 244.329
R1703 VGND.n9 VGND.n3 244.329
R1704 VGND.n680 VGND.t1239 241.393
R1705 VGND.n2578 VGND.t946 241.393
R1706 VGND.n233 VGND.t16 241.393
R1707 VGND.n243 VGND.t1850 241.393
R1708 VGND.n183 VGND.t2020 241.393
R1709 VGND.n1423 VGND.t1085 241.393
R1710 VGND.n641 VGND.t2066 241.393
R1711 VGND.n620 VGND.t6 241.393
R1712 VGND.n647 VGND.t1840 241.393
R1713 VGND.n663 VGND.t363 241.393
R1714 VGND.n672 VGND.t1245 241.393
R1715 VGND.n1375 VGND.t2056 241.393
R1716 VGND.n1307 VGND.t1848 241.393
R1717 VGND.n576 VGND.t2054 241.393
R1718 VGND.n572 VGND.t241 241.393
R1719 VGND.n675 VGND.t1890 241.393
R1720 VGND.n829 VGND.t49 241.393
R1721 VGND.n819 VGND.t949 241.393
R1722 VGND.n1291 VGND.t1169 241.284
R1723 VGND.n687 VGND.t2012 241.284
R1724 VGND.n727 VGND.t1858 241.284
R1725 VGND.n732 VGND.t1406 241.284
R1726 VGND.n737 VGND.t1355 241.284
R1727 VGND.n742 VGND.t1852 241.284
R1728 VGND.n747 VGND.t1219 241.284
R1729 VGND.n752 VGND.t776 241.284
R1730 VGND.n757 VGND.t22 241.284
R1731 VGND.n762 VGND.t1736 241.284
R1732 VGND.n767 VGND.t1894 241.284
R1733 VGND.n772 VGND.t18 241.284
R1734 VGND.n777 VGND.t2389 241.284
R1735 VGND.n782 VGND.t227 241.284
R1736 VGND.n1234 VGND.t985 241.284
R1737 VGND.n1229 VGND.t943 241.284
R1738 VGND.n798 VGND.t1027 241.284
R1739 VGND.n1210 VGND.t1018 241.284
R1740 VGND.n1202 VGND.t979 241.284
R1741 VGND.n1197 VGND.t931 241.284
R1742 VGND.n806 VGND.t1015 241.284
R1743 VGND.n1178 VGND.t976 241.284
R1744 VGND.n1170 VGND.t967 241.284
R1745 VGND.n1165 VGND.t925 241.284
R1746 VGND.n814 VGND.t1003 241.284
R1747 VGND.n1146 VGND.t997 241.284
R1748 VGND.n1138 VGND.t922 241.284
R1749 VGND.n1133 VGND.t904 241.284
R1750 VGND.n1128 VGND.t898 241.284
R1751 VGND.n2580 VGND.t895 241.284
R1752 VGND.n2576 VGND.t901 241.284
R1753 VGND.n2706 VGND.t907 241.284
R1754 VGND.n2631 VGND.t994 241.284
R1755 VGND.n2698 VGND.t1000 241.284
R1756 VGND.n2635 VGND.t913 241.284
R1757 VGND.n2690 VGND.t955 241.284
R1758 VGND.n2639 VGND.t970 241.284
R1759 VGND.n2682 VGND.t1006 241.284
R1760 VGND.n2643 VGND.t928 241.284
R1761 VGND.n2674 VGND.t973 241.284
R1762 VGND.n2647 VGND.t1012 241.284
R1763 VGND.n2666 VGND.t1024 241.284
R1764 VGND.n2651 VGND.t940 241.284
R1765 VGND.n2658 VGND.t982 241.284
R1766 VGND.n236 VGND.t786 241.284
R1767 VGND.n2721 VGND.t1888 241.284
R1768 VGND.n2726 VGND.t2052 241.284
R1769 VGND.n2731 VGND.t1724 241.284
R1770 VGND.n2736 VGND.t1089 241.284
R1771 VGND.n2741 VGND.t2357 241.284
R1772 VGND.n2746 VGND.t2379 241.284
R1773 VGND.n2751 VGND.t2022 241.284
R1774 VGND.n2756 VGND.t1237 241.284
R1775 VGND.n2761 VGND.t1414 241.284
R1776 VGND.n2766 VGND.t2010 241.284
R1777 VGND.n2771 VGND.t1229 241.284
R1778 VGND.n2776 VGND.t1223 241.284
R1779 VGND.n2781 VGND.t1353 241.284
R1780 VGND.n231 VGND.t347 241.284
R1781 VGND.n246 VGND.t1371 241.284
R1782 VGND.n2515 VGND.t47 241.284
R1783 VGND.n2510 VGND.t2387 241.284
R1784 VGND.n250 VGND.t788 241.284
R1785 VGND.n2440 VGND.t2072 241.284
R1786 VGND.n2445 VGND.t2383 241.284
R1787 VGND.n2450 VGND.t1726 241.284
R1788 VGND.n2455 VGND.t1091 241.284
R1789 VGND.n2460 VGND.t2050 241.284
R1790 VGND.n2465 VGND.t1179 241.284
R1791 VGND.n2470 VGND.t1077 241.284
R1792 VGND.n2475 VGND.t2349 241.284
R1793 VGND.n2480 VGND.t1418 241.284
R1794 VGND.n2485 VGND.t349 241.284
R1795 VGND.n2490 VGND.t1231 241.284
R1796 VGND.n2833 VGND.t2341 241.284
R1797 VGND.n370 VGND.t1410 241.284
R1798 VGND.n374 VGND.t1361 241.284
R1799 VGND.n2173 VGND.t1062 241.284
R1800 VGND.n368 VGND.t1205 241.284
R1801 VGND.n2199 VGND.t1349 241.284
R1802 VGND.n360 VGND.t2641 241.284
R1803 VGND.n2225 VGND.t1738 241.284
R1804 VGND.n352 VGND.t1900 241.284
R1805 VGND.n2251 VGND.t20 241.284
R1806 VGND.n344 VGND.t1732 241.284
R1807 VGND.n2282 VGND.t1892 241.284
R1808 VGND.n2287 VGND.t1986 241.284
R1809 VGND.n2292 VGND.t1187 241.284
R1810 VGND.n336 VGND.t243 241.284
R1811 VGND.n1430 VGND.t2371 241.284
R1812 VGND.n1427 VGND.t1173 241.284
R1813 VGND.n2160 VGND.t355 241.284
R1814 VGND.n383 VGND.t2343 241.284
R1815 VGND.n2186 VGND.t2232 241.284
R1816 VGND.n364 VGND.t2643 241.284
R1817 VGND.n2212 VGND.t1064 241.284
R1818 VGND.n356 VGND.t1207 241.284
R1819 VGND.n2238 VGND.t1351 241.284
R1820 VGND.n348 VGND.t1854 241.284
R1821 VGND.n2264 VGND.t796 241.284
R1822 VGND.n340 VGND.t53 241.284
R1823 VGND.n2269 VGND.t24 241.284
R1824 VGND.n2309 VGND.t245 241.284
R1825 VGND.n2314 VGND.t1896 241.284
R1826 VGND.n1444 VGND.t1718 241.284
R1827 VGND.n638 VGND.t231 241.284
R1828 VGND.n1494 VGND.t1241 241.284
R1829 VGND.n1489 VGND.t2373 241.284
R1830 VGND.n1484 VGND.t2016 241.284
R1831 VGND.n1479 VGND.t1066 241.284
R1832 VGND.n1474 VGND.t2345 241.284
R1833 VGND.n1469 VGND.t2236 241.284
R1834 VGND.n1464 VGND.t343 241.284
R1835 VGND.n1459 VGND.t1221 241.284
R1836 VGND.n1454 VGND.t2224 241.284
R1837 VGND.n1449 VGND.t2639 241.284
R1838 VGND.n397 VGND.t1856 241.284
R1839 VGND.n2137 VGND.t1898 241.284
R1840 VGND.n2132 VGND.t57 241.284
R1841 VGND.n1506 VGND.t778 241.284
R1842 VGND.n625 VGND.t1878 241.284
R1843 VGND.n629 VGND.t2351 241.284
R1844 VGND.n1999 VGND.t249 241.284
R1845 VGND.n435 VGND.t1247 241.284
R1846 VGND.n2025 VGND.t2337 241.284
R1847 VGND.n427 VGND.t2367 241.284
R1848 VGND.n2051 VGND.t365 241.284
R1849 VGND.n419 VGND.t1058 241.284
R1850 VGND.n2077 VGND.t2240 241.284
R1851 VGND.n411 VGND.t359 241.284
R1852 VGND.n2108 VGND.t1054 241.284
R1853 VGND.n2113 VGND.t1215 241.284
R1854 VGND.n2118 VGND.t51 241.284
R1855 VGND.n2123 VGND.t2633 241.284
R1856 VGND.n654 VGND.t1359 241.284
R1857 VGND.n651 VGND.t35 241.284
R1858 VGND.n1986 VGND.t2377 241.284
R1859 VGND.n439 VGND.t780 241.284
R1860 VGND.n2012 VGND.t2058 241.284
R1861 VGND.n431 VGND.t2369 241.284
R1862 VGND.n2038 VGND.t1716 241.284
R1863 VGND.n423 VGND.t1075 241.284
R1864 VGND.n2064 VGND.t2339 241.284
R1865 VGND.n415 VGND.t2028 241.284
R1866 VGND.n2090 VGND.t1243 241.284
R1867 VGND.n407 VGND.t2335 241.284
R1868 VGND.n2095 VGND.t2242 241.284
R1869 VGND.n2334 VGND.t2635 241.284
R1870 VGND.n2339 VGND.t1056 241.284
R1871 VGND.n961 VGND.t1424 241.284
R1872 VGND.n956 VGND.t2238 241.284
R1873 VGND.n951 VGND.t55 241.284
R1874 VGND.n946 VGND.t1046 241.284
R1875 VGND.n941 VGND.t792 241.284
R1876 VGND.n936 VGND.t41 241.284
R1877 VGND.n931 VGND.t2627 241.284
R1878 VGND.n926 VGND.t1730 241.284
R1879 VGND.n921 VGND.t1886 241.284
R1880 VGND.n916 VGND.t12 241.284
R1881 VGND.n911 VGND.t1720 241.284
R1882 VGND.n906 VGND.t1880 241.284
R1883 VGND.n453 VGND.t2070 241.284
R1884 VGND.n1963 VGND.t1175 241.284
R1885 VGND.n1958 VGND.t233 241.284
R1886 VGND.n1397 VGND.t1189 241.284
R1887 VGND.n1402 VGND.t2026 241.284
R1888 VGND.n670 VGND.t2637 241.284
R1889 VGND.n1825 VGND.t1426 241.284
R1890 VGND.n491 VGND.t2220 241.284
R1891 VGND.n1851 VGND.t2629 241.284
R1892 VGND.n483 VGND.t1048 241.284
R1893 VGND.n1877 VGND.t794 241.284
R1894 VGND.n475 VGND.t45 241.284
R1895 VGND.n1903 VGND.t1844 241.284
R1896 VGND.n467 VGND.t784 241.284
R1897 VGND.n1934 VGND.t37 241.284
R1898 VGND.n1939 VGND.t14 241.284
R1899 VGND.n1944 VGND.t235 241.284
R1900 VGND.n1949 VGND.t1882 241.284
R1901 VGND.n1382 VGND.t247 241.284
R1902 VGND.n1379 VGND.t229 241.284
R1903 VGND.n1812 VGND.t1060 241.284
R1904 VGND.n495 VGND.t1191 241.284
R1905 VGND.n1838 VGND.t361 241.284
R1906 VGND.n487 VGND.t1050 241.284
R1907 VGND.n1864 VGND.t1428 241.284
R1908 VGND.n479 VGND.t2222 241.284
R1909 VGND.n1890 VGND.t2631 241.284
R1910 VGND.n471 VGND.t1213 241.284
R1911 VGND.n1916 VGND.t1367 241.284
R1912 VGND.n463 VGND.t2625 241.284
R1913 VGND.n1921 VGND.t1846 241.284
R1914 VGND.n2359 VGND.t1884 241.284
R1915 VGND.n2364 VGND.t39 241.284
R1916 VGND.n1314 VGND.t1365 241.284
R1917 VGND.n1311 VGND.t43 241.284
R1918 VGND.n1364 VGND.t2385 241.284
R1919 VGND.n1359 VGND.t782 241.284
R1920 VGND.n1354 VGND.t2068 241.284
R1921 VGND.n1349 VGND.t2375 241.284
R1922 VGND.n1344 VGND.t1722 241.284
R1923 VGND.n1339 VGND.t1087 241.284
R1924 VGND.n1334 VGND.t2353 241.284
R1925 VGND.n1329 VGND.t1177 241.284
R1926 VGND.n1324 VGND.t1249 241.284
R1927 VGND.n1319 VGND.t2347 241.284
R1928 VGND.n509 VGND.t1412 241.284
R1929 VGND.n1789 VGND.t345 241.284
R1930 VGND.n1784 VGND.t1227 241.284
R1931 VGND.n1519 VGND.t239 241.284
R1932 VGND.n1524 VGND.t1095 241.284
R1933 VGND.n581 VGND.t1052 241.284
R1934 VGND.n1651 VGND.t1185 241.284
R1935 VGND.n547 VGND.t357 241.284
R1936 VGND.n1677 VGND.t1044 241.284
R1937 VGND.n539 VGND.t1422 241.284
R1938 VGND.n1703 VGND.t1369 241.284
R1939 VGND.n531 VGND.t2623 241.284
R1940 VGND.n1729 VGND.t1209 241.284
R1941 VGND.n523 VGND.t1363 241.284
R1942 VGND.n1760 VGND.t2621 241.284
R1943 VGND.n1765 VGND.t1836 241.284
R1944 VGND.n1770 VGND.t1201 241.284
R1945 VGND.n1775 VGND.t26 241.284
R1946 VGND.n1539 VGND.t4 241.284
R1947 VGND.n570 VGND.t2381 241.284
R1948 VGND.n1638 VGND.t2024 241.284
R1949 VGND.n551 VGND.t2060 241.284
R1950 VGND.n1664 VGND.t1416 241.284
R1951 VGND.n543 VGND.t2014 241.284
R1952 VGND.n1690 VGND.t1079 241.284
R1953 VGND.n535 VGND.t1225 241.284
R1954 VGND.n1716 VGND.t2234 241.284
R1955 VGND.n527 VGND.t351 241.284
R1956 VGND.n1742 VGND.t1217 241.284
R1957 VGND.n519 VGND.t2226 241.284
R1958 VGND.n1747 VGND.t1357 241.284
R1959 VGND.n2384 VGND.t1734 241.284
R1960 VGND.n2389 VGND.t798 241.284
R1961 VGND.n678 VGND.t1838 241.284
R1962 VGND.n1552 VGND.t1728 241.284
R1963 VGND.n1557 VGND.t1093 241.284
R1964 VGND.n1562 VGND.t8 241.284
R1965 VGND.n1567 VGND.t1181 241.284
R1966 VGND.n1572 VGND.t1081 241.284
R1967 VGND.n1577 VGND.t2062 241.284
R1968 VGND.n1582 VGND.t1420 241.284
R1969 VGND.n1587 VGND.t2018 241.284
R1970 VGND.n1592 VGND.t1233 241.284
R1971 VGND.n1597 VGND.t1408 241.284
R1972 VGND.n1602 VGND.t2006 241.284
R1973 VGND.n565 VGND.t353 241.284
R1974 VGND.n1615 VGND.t1203 241.284
R1975 VGND.n1610 VGND.t2228 241.284
R1976 VGND.n837 VGND.t1211 241.284
R1977 VGND.n842 VGND.t790 241.284
R1978 VGND.n834 VGND.t1982 241.284
R1979 VGND.n892 VGND.t1842 241.284
R1980 VGND.n887 VGND.t237 241.284
R1981 VGND.n882 VGND.t2064 241.284
R1982 VGND.n877 VGND.t10 241.284
R1983 VGND.n872 VGND.t1183 241.284
R1984 VGND.n867 VGND.t1083 241.284
R1985 VGND.n862 VGND.t2355 241.284
R1986 VGND.n857 VGND.t1171 241.284
R1987 VGND.n852 VGND.t1073 241.284
R1988 VGND.n847 VGND.t1235 241.284
R1989 VGND.n2404 VGND.t2230 241.284
R1990 VGND.n2409 VGND.t2008 241.284
R1991 VGND.n723 VGND.t1984 241.284
R1992 VGND.t696 VGND.t945 222.15
R1993 VGND.t1465 VGND.t1643 222.15
R1994 VGND.t2500 VGND.t894 222.15
R1995 VGND.t1957 VGND.t2430 222.15
R1996 VGND.t900 VGND.t2422 222.15
R1997 VGND.t2417 VGND.t1403 222.15
R1998 VGND.t758 VGND.t906 222.15
R1999 VGND.t420 VGND.t1702 222.15
R2000 VGND.t993 VGND.t689 222.15
R2001 VGND.t2496 VGND.t1953 222.15
R2002 VGND.t2478 VGND.t999 222.15
R2003 VGND.t869 VGND.t760 222.15
R2004 VGND.t912 VGND.t2464 222.15
R2005 VGND.t691 VGND.t1269 222.15
R2006 VGND.t685 VGND.t954 222.15
R2007 VGND.t158 VGND.t1690 222.15
R2008 VGND.t969 VGND.t1686 222.15
R2009 VGND.t2466 VGND.t1327 222.15
R2010 VGND.t2480 VGND.t1005 222.15
R2011 VGND.t75 VGND.t761 222.15
R2012 VGND.t927 VGND.t741 222.15
R2013 VGND.t1688 VGND.t250 222.15
R2014 VGND.t726 VGND.t972 222.15
R2015 VGND.t639 VGND.t1678 222.15
R2016 VGND.t1011 VGND.t2462 222.15
R2017 VGND.t2457 VGND.t2141 222.15
R2018 VGND.t2450 VGND.t1023 222.15
R2019 VGND.t1142 VGND.t730 222.15
R2020 VGND.t939 VGND.t2434 222.15
R2021 VGND.t707 VGND.t175 222.15
R2022 VGND.t981 VGND.t1671 222.15
R2023 VGND.t2454 VGND.t1924 222.15
R2024 VGND.t2089 VGND.t15 222.15
R2025 VGND.t2504 VGND.t1527 222.15
R2026 VGND.t785 VGND.t1376 222.15
R2027 VGND.t1292 VGND.t79 222.15
R2028 VGND.t1477 VGND.t1887 222.15
R2029 VGND.t2619 VGND.t157 222.15
R2030 VGND.t2095 VGND.t2051 222.15
R2031 VGND.t1118 VGND.t1385 222.15
R2032 VGND.t2087 VGND.t1723 222.15
R2033 VGND.t1326 VGND.t1990 222.15
R2034 VGND.t1487 VGND.t1088 222.15
R2035 VGND.t1144 VGND.t1541 222.15
R2036 VGND.t1485 VGND.t2356 222.15
R2037 VGND.t1400 VGND.t2662 222.15
R2038 VGND.t2085 VGND.t2378 222.15
R2039 VGND.t179 VGND.t381 222.15
R2040 VGND.t1380 VGND.t2021 222.15
R2041 VGND.t83 VGND.t285 222.15
R2042 VGND.t1489 VGND.t1236 222.15
R2043 VGND.t2607 VGND.t558 222.15
R2044 VGND.t2093 VGND.t1413 222.15
R2045 VGND.t1322 VGND.t1921 222.15
R2046 VGND.t2091 VGND.t2009 222.15
R2047 VGND.t1139 VGND.t167 222.15
R2048 VGND.t1483 VGND.t1228 222.15
R2049 VGND.t803 VGND.t585 222.15
R2050 VGND.t1481 VGND.t1222 222.15
R2051 VGND.t1321 VGND.t1810 222.15
R2052 VGND.t1479 VGND.t1352 222.15
R2053 VGND.t475 VGND.t1504 222.15
R2054 VGND.t346 VGND.t1378 222.15
R2055 VGND.t1679 VGND.t1431 222.15
R2056 VGND.t2319 VGND.t1849 222.15
R2057 VGND.t1804 VGND.t1151 222.15
R2058 VGND.t1370 VGND.t2332 222.15
R2059 VGND.t2261 VGND.t225 222.15
R2060 VGND.t46 VGND.t1594 222.15
R2061 VGND.t93 VGND.t1392 222.15
R2062 VGND.t1592 VGND.t2386 222.15
R2063 VGND.t1614 VGND.t2517 222.15
R2064 VGND.t2317 VGND.t787 222.15
R2065 VGND.t82 VGND.t1707 222.15
R2066 VGND.t2328 VGND.t2071 222.15
R2067 VGND.t2654 VGND.t124 222.15
R2068 VGND.t2326 VGND.t2382 222.15
R2069 VGND.t1339 VGND.t1308 222.15
R2070 VGND.t2315 VGND.t1725 222.15
R2071 VGND.t1535 VGND.t1758 222.15
R2072 VGND.t2313 VGND.t1090 222.15
R2073 VGND.t1143 VGND.t474 222.15
R2074 VGND.t2330 VGND.t2049 222.15
R2075 VGND.t1591 VGND.t32 222.15
R2076 VGND.t2075 VGND.t1178 222.15
R2077 VGND.t1915 VGND.t1440 222.15
R2078 VGND.t2073 VGND.t1076 222.15
R2079 VGND.t641 VGND.t2593 222.15
R2080 VGND.t2324 VGND.t2348 222.15
R2081 VGND.t2206 VGND.t308 222.15
R2082 VGND.t2322 VGND.t1417 222.15
R2083 VGND.t1518 VGND.t113 222.15
R2084 VGND.t1596 VGND.t348 222.15
R2085 VGND.t58 VGND.t2118 222.15
R2086 VGND.t2311 VGND.t1230 222.15
R2087 VGND.t1 VGND.t745 222.15
R2088 VGND.t2019 VGND.t1284 222.15
R2089 VGND.t1925 VGND.t865 222.15
R2090 VGND.t1625 VGND.t2340 222.15
R2091 VGND.t804 VGND.t1298 222.15
R2092 VGND.t1608 VGND.t1409 222.15
R2093 VGND.t2508 VGND.t147 222.15
R2094 VGND.t1360 VGND.t1606 222.15
R2095 VGND.t1391 VGND.t872 222.15
R2096 VGND.t1282 VGND.t1061 222.15
R2097 VGND.t1958 VGND.t2081 222.15
R2098 VGND.t1204 VGND.t2003 222.15
R2099 VGND.t1543 VGND.t1799 222.15
R2100 VGND.t2001 VGND.t1348 222.15
R2101 VGND.t203 VGND.t2668 222.15
R2102 VGND.t2640 VGND.t1280 222.15
R2103 VGND.t387 VGND.t115 222.15
R2104 VGND.t1629 VGND.t1737 222.15
R2105 VGND.t1914 VGND.t1155 222.15
R2106 VGND.t1899 VGND.t1623 222.15
R2107 VGND.t568 VGND.t1300 222.15
R2108 VGND.t1288 VGND.t19 222.15
R2109 VGND.t2523 VGND.t766 222.15
R2110 VGND.t1731 VGND.t1286 222.15
R2111 VGND.t1107 VGND.t1640 222.15
R2112 VGND.t1999 VGND.t1891 222.15
R2113 VGND.t1517 VGND.t591 222.15
R2114 VGND.t1864 VGND.t1985 222.15
R2115 VGND.t1152 VGND.t1034 222.15
R2116 VGND.t1610 VGND.t1186 222.15
R2117 VGND.t886 VGND.t1510 222.15
R2118 VGND.t242 VGND.t1627 222.15
R2119 VGND.t1700 VGND.t1618 222.15
R2120 VGND.t273 VGND.t1084 222.15
R2121 VGND.t279 VGND.t1116 222.15
R2122 VGND.t2217 VGND.t2370 222.15
R2123 VGND.t193 VGND.t833 222.15
R2124 VGND.t1172 VGND.t1434 222.15
R2125 VGND.t799 VGND.t2675 222.15
R2126 VGND.t1432 VGND.t354 222.15
R2127 VGND.t1125 VGND.t60 222.15
R2128 VGND.t2342 VGND.t271 222.15
R2129 VGND.t2243 VGND.t70 222.15
R2130 VGND.t2213 VGND.t2231 222.15
R2131 VGND.t1790 VGND.t1901 222.15
R2132 VGND.t2642 VGND.t2211 222.15
R2133 VGND.t2655 VGND.t1141 222.15
R2134 VGND.t269 VGND.t1063 222.15
R2135 VGND.t178 VGND.t862 222.15
R2136 VGND.t1206 VGND.t2559 222.15
R2137 VGND.t884 VGND.t1800 222.15
R2138 VGND.t2215 VGND.t1350 222.15
R2139 VGND.t646 VGND.t528 222.15
R2140 VGND.t1853 VGND.t277 222.15
R2141 VGND.t2528 VGND.t1935 222.15
R2142 VGND.t275 VGND.t795 222.15
R2143 VGND.t1277 VGND.t1975 222.15
R2144 VGND.t52 VGND.t2209 222.15
R2145 VGND.t2200 VGND.t2522 222.15
R2146 VGND.t23 VGND.t2207 222.15
R2147 VGND.t1819 VGND.t1798 222.15
R2148 VGND.t1436 VGND.t244 222.15
R2149 VGND.t1642 VGND.t2125 222.15
R2150 VGND.t1895 VGND.t2557 222.15
R2151 VGND.t2495 VGND.t86 222.15
R2152 VGND.t2603 VGND.t2065 222.15
R2153 VGND.t844 VGND.t1145 222.15
R2154 VGND.t2105 VGND.t1717 222.15
R2155 VGND.t253 VGND.t2255 222.15
R2156 VGND.t230 VGND.t2249 222.15
R2157 VGND.t128 VGND.t1268 222.15
R2158 VGND.t1240 VGND.t1548 222.15
R2159 VGND.t2511 VGND.t871 222.15
R2160 VGND.t2372 VGND.t2601 222.15
R2161 VGND.t1964 VGND.t1789 222.15
R2162 VGND.t2015 VGND.t2101 222.15
R2163 VGND.t2544 VGND.t27 222.15
R2164 VGND.t1065 VGND.t2099 222.15
R2165 VGND.t2404 VGND.t2506 222.15
R2166 VGND.t2344 VGND.t2599 222.15
R2167 VGND.t1740 VGND.t1153 222.15
R2168 VGND.t2235 VGND.t2597 222.15
R2169 VGND.t468 VGND.t2142 222.15
R2170 VGND.t342 VGND.t2103 222.15
R2171 VGND.t539 VGND.t1519 222.15
R2172 VGND.t1220 VGND.t1546 222.15
R2173 VGND.t2566 VGND.t292 222.15
R2174 VGND.t2223 VGND.t1544 222.15
R2175 VGND.t2608 VGND.t1533 222.15
R2176 VGND.t2638 VGND.t2097 222.15
R2177 VGND.t302 VGND.t870 222.15
R2178 VGND.t1855 VGND.t2253 222.15
R2179 VGND.t1808 VGND.t2509 222.15
R2180 VGND.t1897 VGND.t2251 222.15
R2181 VGND.t2112 VGND.t1270 222.15
R2182 VGND.t56 VGND.t2107 222.15
R2183 VGND.t717 VGND.t210 222.15
R2184 VGND.t5 VGND.t2266 222.15
R2185 VGND.t1526 VGND.t1401 222.15
R2186 VGND.t1568 VGND.t777 222.15
R2187 VGND.t78 VGND.t1291 222.15
R2188 VGND.t2280 VGND.t1877 222.15
R2189 VGND.t1955 VGND.t146 222.15
R2190 VGND.t2350 VGND.t2272 222.15
R2191 VGND.t1384 VGND.t1337 222.15
R2192 VGND.t2264 VGND.t248 222.15
R2193 VGND.t888 VGND.t1989 222.15
R2194 VGND.t1246 VGND.t2290 222.15
R2195 VGND.t1540 VGND.t252 222.15
R2196 VGND.t2288 VGND.t2336 222.15
R2197 VGND.t1278 VGND.t2661 222.15
R2198 VGND.t2366 VGND.t2262 222.15
R2199 VGND.t380 VGND.t2617 222.15
R2200 VGND.t1572 VGND.t364 222.15
R2201 VGND.t2539 VGND.t284 222.15
R2202 VGND.t1057 VGND.t2292 222.15
R2203 VGND.t557 VGND.t1438 222.15
R2204 VGND.t2270 VGND.t2239 222.15
R2205 VGND.t1770 VGND.t1920 222.15
R2206 VGND.t358 VGND.t2268 222.15
R2207 VGND.t166 VGND.t645 222.15
R2208 VGND.t2286 VGND.t1053 222.15
R2209 VGND.t114 VGND.t584 222.15
R2210 VGND.t2284 VGND.t1214 222.15
R2211 VGND.t224 VGND.t2041 222.15
R2212 VGND.t2282 VGND.t50 222.15
R2213 VGND.t1875 VGND.t1503 222.15
R2214 VGND.t2632 VGND.t1570 222.15
R2215 VGND.t1677 VGND.t1127 222.15
R2216 VGND.t480 VGND.t1839 222.15
R2217 VGND.t2505 VGND.t1930 222.15
R2218 VGND.t631 VGND.t1358 222.15
R2219 VGND.t1394 VGND.t2163 222.15
R2220 VGND.t34 VGND.t488 222.15
R2221 VGND.t125 VGND.t1923 222.15
R2222 VGND.t486 VGND.t2376 222.15
R2223 VGND.t1129 VGND.t1161 222.15
R2224 VGND.t779 VGND.t478 222.15
R2225 VGND.t2082 VGND.t2538 222.15
R2226 VGND.t627 VGND.t2057 222.15
R2227 VGND.t1128 VGND.t2550 222.15
R2228 VGND.t2368 VGND.t625 222.15
R2229 VGND.t2398 VGND.t2556 222.15
R2230 VGND.t476 VGND.t1715 222.15
R2231 VGND.t211 VGND.t1067 222.15
R2232 VGND.t1074 VGND.t635 222.15
R2233 VGND.t1156 VGND.t1429 222.15
R2234 VGND.t629 VGND.t2338 222.15
R2235 VGND.t1455 VGND.t569 222.15
R2236 VGND.t2027 VGND.t484 222.15
R2237 VGND.t767 VGND.t880 222.15
R2238 VGND.t482 VGND.t1242 222.15
R2239 VGND.t1617 VGND.t1108 222.15
R2240 VGND.t2334 VGND.t652 222.15
R2241 VGND.t1792 VGND.t1874 222.15
R2242 VGND.t2241 VGND.t637 222.15
R2243 VGND.t1035 VGND.t85 222.15
R2244 VGND.t490 VGND.t2634 222.15
R2245 VGND.t266 VGND.t1511 222.15
R2246 VGND.t1055 VGND.t633 222.15
R2247 VGND.t1703 VGND.t1771 222.15
R2248 VGND.t362 VGND.t1271 222.15
R2249 VGND.t1117 VGND.t1639 222.15
R2250 VGND.t1423 VGND.t1961 222.15
R2251 VGND.t834 VGND.t864 222.15
R2252 VGND.t2237 VGND.t818 222.15
R2253 VGND.t802 VGND.t123 222.15
R2254 VGND.t54 VGND.t816 222.15
R2255 VGND.t61 VGND.t76 222.15
R2256 VGND.t1045 VGND.t2139 222.15
R2257 VGND.t2244 VGND.t180 222.15
R2258 VGND.t791 VGND.t1040 222.15
R2259 VGND.t1902 VGND.t1138 222.15
R2260 VGND.t40 VGND.t1038 222.15
R2261 VGND.t2656 VGND.t583 222.15
R2262 VGND.t2626 VGND.t2137 222.15
R2263 VGND.t863 VGND.t1042 222.15
R2264 VGND.t1729 VGND.t2135 222.15
R2265 VGND.t885 VGND.t1532 222.15
R2266 VGND.t1885 VGND.t1959 222.15
R2267 VGND.t529 VGND.t1613 222.15
R2268 VGND.t11 VGND.t1275 222.15
R2269 VGND.t2529 VGND.t1525 222.15
R2270 VGND.t1719 VGND.t1273 222.15
R2271 VGND.t1976 VGND.t2310 222.15
R2272 VGND.t1879 VGND.t1036 222.15
R2273 VGND.t2201 VGND.t1522 222.15
R2274 VGND.t2069 VGND.t822 222.15
R2275 VGND.t1820 VGND.t421 222.15
R2276 VGND.t1174 VGND.t820 222.15
R2277 VGND.t2126 VGND.t1324 222.15
R2278 VGND.t232 VGND.t2133 222.15
R2279 VGND.t2497 VGND.t680 222.15
R2280 VGND.t2161 VGND.t1244 222.15
R2281 VGND.t830 VGND.t1114 222.15
R2282 VGND.t2037 VGND.t1188 222.15
R2283 VGND.t2618 VGND.t832 222.15
R2284 VGND.t2396 VGND.t2025 222.15
R2285 VGND.t881 VGND.t801 222.15
R2286 VGND.t2636 VGND.t2394 222.15
R2287 VGND.t59 VGND.t2648 222.15
R2288 VGND.t2159 VGND.t1425 222.15
R2289 VGND.t805 VGND.t650 222.15
R2290 VGND.t2219 VGND.t2033 222.15
R2291 VGND.t1566 VGND.t1119 222.15
R2292 VGND.t2031 VGND.t2628 222.15
R2293 VGND.t2520 VGND.t668 222.15
R2294 VGND.t1047 VGND.t2157 222.15
R2295 VGND.t861 VGND.t2145 222.15
R2296 VGND.t2155 VGND.t793 222.15
R2297 VGND.t1772 VGND.t883 222.15
R2298 VGND.t44 VGND.t2035 222.15
R2299 VGND.t527 VGND.t1521 222.15
R2300 VGND.t2392 VGND.t1843 222.15
R2301 VGND.t2146 VGND.t2527 222.15
R2302 VGND.t783 VGND.t2390 222.15
R2303 VGND.t1974 VGND.t1404 222.15
R2304 VGND.t2029 VGND.t36 222.15
R2305 VGND.t2682 VGND.t2199 222.15
R2306 VGND.t1576 VGND.t13 222.15
R2307 VGND.t1537 VGND.t1830 222.15
R2308 VGND.t1574 VGND.t234 222.15
R2309 VGND.t1797 VGND.t2123 222.15
R2310 VGND.t1881 VGND.t867 222.15
R2311 VGND.t2488 VGND.t1952 222.15
R2312 VGND.t1785 VGND.t2055 222.15
R2313 VGND.t677 VGND.t1452 222.15
R2314 VGND.t1775 VGND.t246 222.15
R2315 VGND.t1637 VGND.t1605 222.15
R2316 VGND.t228 VGND.t1872 222.15
R2317 VGND.t131 VGND.t647 222.15
R2318 VGND.t1870 VGND.t1059 222.15
R2319 VGND.t1705 VGND.t2510 222.15
R2320 VGND.t1190 VGND.t1783 222.15
R2321 VGND.t1963 VGND.t165 222.15
R2322 VGND.t1474 VGND.t360 222.15
R2323 VGND.t1451 VGND.t2543 222.15
R2324 VGND.t1049 VGND.t1472 222.15
R2325 VGND.t2403 VGND.t1590 222.15
R2326 VGND.t1781 VGND.t1427 222.15
R2327 VGND.t644 VGND.t1739 222.15
R2328 VGND.t2221 VGND.t1779 222.15
R2329 VGND.t2168 VGND.t807 222.15
R2330 VGND.t1773 VGND.t2630 222.15
R2331 VGND.t1631 VGND.t536 222.15
R2332 VGND.t1212 VGND.t1868 222.15
R2333 VGND.t2565 VGND.t106 222.15
R2334 VGND.t1866 VGND.t1366 222.15
R2335 VGND.t422 VGND.t1861 222.15
R2336 VGND.t2624 VGND.t1470 222.15
R2337 VGND.t301 VGND.t1987 222.15
R2338 VGND.t1845 VGND.t1468 222.15
R2339 VGND.t1805 VGND.t1267 222.15
R2340 VGND.t1466 VGND.t1883 222.15
R2341 VGND.t329 VGND.t2111 222.15
R2342 VGND.t38 VGND.t1777 222.15
R2343 VGND.t712 VGND.t2537 222.15
R2344 VGND.t511 VGND.t1847 222.15
R2345 VGND.t845 VGND.t825 222.15
R2346 VGND.t574 VGND.t1364 222.15
R2347 VGND.t582 VGND.t2677 222.15
R2348 VGND.t42 VGND.t2574 222.15
R2349 VGND.t769 VGND.t2535 222.15
R2350 VGND.t2384 VGND.t2572 222.15
R2351 VGND.t603 VGND.t1803 222.15
R2352 VGND.t781 VGND.t509 222.15
R2353 VGND.t2150 VGND.t81 222.15
R2354 VGND.t2067 VGND.t570 222.15
R2355 VGND.t164 VGND.t267 222.15
R2356 VGND.t2374 VGND.t2582 222.15
R2357 VGND.t662 VGND.t1100 222.15
R2358 VGND.t1721 VGND.t580 222.15
R2359 VGND.t2684 VGND.t1988 222.15
R2360 VGND.t1086 VGND.t578 222.15
R2361 VGND.t1131 VGND.t1638 222.15
R2362 VGND.t2352 VGND.t572 222.15
R2363 VGND.t522 VGND.t2555 222.15
R2364 VGND.t1176 VGND.t2570 222.15
R2365 VGND.t2042 VGND.t1340 222.15
R2366 VGND.t1248 VGND.t2568 222.15
R2367 VGND.t1834 VGND.t1402 222.15
R2368 VGND.t2346 VGND.t2580 222.15
R2369 VGND.t403 VGND.t2534 222.15
R2370 VGND.t1411 VGND.t2578 222.15
R2371 VGND.t1828 VGND.t1632 222.15
R2372 VGND.t344 VGND.t2576 222.15
R2373 VGND.t73 VGND.t1266 222.15
R2374 VGND.t1226 VGND.t576 222.15
R2375 VGND.t2447 VGND.t1616 222.15
R2376 VGND.t858 VGND.t2053 222.15
R2377 VGND.t419 VGND.t1528 222.15
R2378 VGND.t848 VGND.t238 222.15
R2379 VGND.t2507 VGND.t1293 222.15
R2380 VGND.t1497 VGND.t1094 222.15
R2381 VGND.t2144 VGND.t148 222.15
R2382 VGND.t1051 VGND.t1495 222.15
R2383 VGND.t1390 VGND.t1279 222.15
R2384 VGND.t856 VGND.t1184 222.15
R2385 VGND.t1453 VGND.t1991 222.15
R2386 VGND.t356 VGND.t658 222.15
R2387 VGND.t1542 VGND.t1524 222.15
R2388 VGND.t656 VGND.t1043 222.15
R2389 VGND.t176 VGND.t2663 222.15
R2390 VGND.t1421 VGND.t854 222.15
R2391 VGND.t382 VGND.t1801 222.15
R2392 VGND.t852 VGND.t1368 222.15
R2393 VGND.t2153 VGND.t1460 222.15
R2394 VGND.t2622 VGND.t660 222.15
R2395 VGND.t567 VGND.t1476 222.15
R2396 VGND.t1493 VGND.t1208 222.15
R2397 VGND.t873 VGND.t1922 222.15
R2398 VGND.t1362 VGND.t1491 222.15
R2399 VGND.t1106 VGND.t640 222.15
R2400 VGND.t654 VGND.t2620 222.15
R2401 VGND.t2409 VGND.t586 222.15
R2402 VGND.t295 VGND.t1835 222.15
R2403 VGND.t2195 VGND.t1033 222.15
R2404 VGND.t1499 VGND.t1200 222.15
R2405 VGND.t2187 VGND.t1509 222.15
R2406 VGND.t25 VGND.t850 222.15
R2407 VGND.t1697 VGND.t2554 222.15
R2408 VGND.t240 VGND.t2669 222.15
R2409 VGND.t824 VGND.t71 222.15
R2410 VGND.t336 VGND.t3 222.15
R2411 VGND.t1615 VGND.t2676 222.15
R2412 VGND.t2380 VGND.t1761 222.15
R2413 VGND.t772 VGND.t1301 222.15
R2414 VGND.t1759 VGND.t2023 222.15
R2415 VGND.t80 VGND.t602 222.15
R2416 VGND.t2059 VGND.t1552 222.15
R2417 VGND.t2149 VGND.t1636 222.15
R2418 VGND.t332 VGND.t1415 222.15
R2419 VGND.t74 VGND.t163 222.15
R2420 VGND.t2013 VGND.t330 222.15
R2421 VGND.t1320 VGND.t1791 222.15
R2422 VGND.t1550 VGND.t1078 222.15
R2423 VGND.t1306 VGND.t370 222.15
R2424 VGND.t1224 VGND.t340 222.15
R2425 VGND.t1130 VGND.t1154 222.15
R2426 VGND.t334 VGND.t2233 222.15
R2427 VGND.t1520 VGND.t519 222.15
R2428 VGND.t350 VGND.t2673 222.15
R2429 VGND.t878 VGND.t1954 222.15
R2430 VGND.t2671 VGND.t1216 222.15
R2431 VGND.t1620 VGND.t1831 222.15
R2432 VGND.t2225 VGND.t1767 222.15
R2433 VGND.t402 VGND.t2154 222.15
R2434 VGND.t1356 VGND.t1765 222.15
R2435 VGND.t1825 VGND.t808 222.15
R2436 VGND.t1763 VGND.t1733 222.15
R2437 VGND.t1323 VGND.t72 222.15
R2438 VGND.t797 VGND.t338 222.15
R2439 VGND.t2444 VGND.t1305 222.15
R2440 VGND.t1945 VGND.t1889 222.15
R2441 VGND.t525 VGND.t1150 222.15
R2442 VGND.t1837 VGND.t2306 222.15
R2443 VGND.t2260 VGND.t2649 222.15
R2444 VGND.t297 VGND.t1727 222.15
R2445 VGND.t889 VGND.t811 222.15
R2446 VGND.t1382 VGND.t1092 222.15
R2447 VGND.t1338 VGND.t2516 222.15
R2448 VGND.t1943 VGND.t7 222.15
R2449 VGND.t524 VGND.t1706 222.15
R2450 VGND.t2302 VGND.t1180 222.15
R2451 VGND.t2321 VGND.t2545 222.15
R2452 VGND.t2300 VGND.t1080 222.15
R2453 VGND.t1120 VGND.t1307 222.15
R2454 VGND.t1941 VGND.t2061 222.15
R2455 VGND.t2295 VGND.t1757 222.15
R2456 VGND.t1939 VGND.t1419 222.15
R2457 VGND.t1302 VGND.t473 222.15
R2458 VGND.t2304 VGND.t2017 222.15
R2459 VGND.t1523 VGND.t540 222.15
R2460 VGND.t1949 VGND.t1232 222.15
R2461 VGND.t1430 VGND.t2567 222.15
R2462 VGND.t1947 VGND.t1407 222.15
R2463 VGND.t1136 VGND.t2609 222.15
R2464 VGND.t2298 VGND.t2005 222.15
R2465 VGND.t84 VGND.t307 222.15
R2466 VGND.t352 VGND.t2296 222.15
R2467 VGND.t1809 VGND.t879 222.15
R2468 VGND.t1202 VGND.t299 222.15
R2469 VGND.t2117 VGND.t2294 222.15
R2470 VGND.t2227 VGND.t2308 222.15
R2471 VGND.t732 VGND.t1951 222.15
R2472 VGND.t194 VGND.t48 222.15
R2473 VGND.t1399 VGND.t1115 222.15
R2474 VGND.t2177 VGND.t1210 222.15
R2475 VGND.t2143 VGND.t831 222.15
R2476 VGND.t2189 VGND.t789 222.15
R2477 VGND.t77 VGND.t800 222.15
R2478 VGND.t1981 VGND.t200 222.15
R2479 VGND.t1196 VGND.t388 222.15
R2480 VGND.t1841 VGND.t2183 222.15
R2481 VGND.t651 VGND.t293 222.15
R2482 VGND.t236 VGND.t2173 222.15
R2483 VGND.t1567 VGND.t2540 222.15
R2484 VGND.t2063 VGND.t2171 222.15
R2485 VGND.t667 VGND.t141 222.15
R2486 VGND.t9 VGND.t2181 222.15
R2487 VGND.t860 VGND.t2644 222.15
R2488 VGND.t1182 VGND.t2179 222.15
R2489 VGND.t882 VGND.t1290 222.15
R2490 VGND.t1082 VGND.t2175 222.15
R2491 VGND.t526 VGND.t251 222.15
R2492 VGND.t2354 VGND.t198 222.15
R2493 VGND.t2526 VGND.t523 222.15
R2494 VGND.t1170 VGND.t196 222.15
R2495 VGND.t1973 VGND.t1536 222.15
R2496 VGND.t1072 VGND.t2169 222.15
R2497 VGND.t2198 VGND.t174 222.15
R2498 VGND.t1234 VGND.t2193 222.15
R2499 VGND.t1829 VGND.t87 222.15
R2500 VGND.t2191 VGND.t2229 222.15
R2501 VGND.t1619 VGND.t2124 222.15
R2502 VGND.t2007 VGND.t809 222.15
R2503 VGND.t2487 VGND.t1137 222.15
R2504 VGND.t1238 VGND.t1665 222.15
R2505 VGND.t1347 VGND.t1704 222.15
R2506 VGND.t2445 VGND.t1168 222.15
R2507 VGND.t806 VGND.t1998 222.15
R2508 VGND.t722 VGND.t2011 222.15
R2509 VGND.t1531 VGND.t768 222.15
R2510 VGND.t700 VGND.t1857 222.15
R2511 VGND.t177 VGND.t599 222.15
R2512 VGND.t1654 VGND.t1405 222.15
R2513 VGND.t1450 VGND.t1714 222.15
R2514 VGND.t2426 VGND.t1354 222.15
R2515 VGND.t1454 VGND.t140 222.15
R2516 VGND.t2415 VGND.t1851 222.15
R2517 VGND.t1099 VGND.t1315 222.15
R2518 VGND.t1650 VGND.t1218 222.15
R2519 VGND.t1304 VGND.t379 222.15
R2520 VGND.t2493 VGND.t775 222.15
R2521 VGND.t1802 VGND.t122 222.15
R2522 VGND.t2428 VGND.t21 222.15
R2523 VGND.t866 VGND.t33 222.15
R2524 VGND.t687 VGND.t1735 222.15
R2525 VGND.t2188 VGND.t1449 222.15
R2526 VGND.t1698 VGND.t1893 222.15
R2527 VGND.t2616 VGND.t2594 222.15
R2528 VGND.t2410 VGND.t17 222.15
R2529 VGND.t1956 VGND.t397 222.15
R2530 VGND.t753 VGND.t2388 222.15
R2531 VGND.t268 VGND.t847 222.15
R2532 VGND.t728 VGND.t226 222.15
R2533 VGND.t1788 VGND.t90 222.15
R2534 VGND.t1983 VGND.t2472 222.15
R2535 VGND.t757 VGND.t1140 222.15
R2536 VGND.n137 VGND.n135 214.365
R2537 VGND.n137 VGND.n136 214.365
R2538 VGND.n127 VGND.n125 214.365
R2539 VGND.n127 VGND.n126 214.365
R2540 VGND.n145 VGND.n143 214.365
R2541 VGND.n145 VGND.n144 214.365
R2542 VGND.n605 VGND.n603 214.365
R2543 VGND.n605 VGND.n604 214.365
R2544 VGND.n595 VGND.n593 214.365
R2545 VGND.n595 VGND.n594 214.365
R2546 VGND.n613 VGND.n611 214.365
R2547 VGND.n613 VGND.n612 214.365
R2548 VGND.n975 VGND.n974 214.365
R2549 VGND.n167 VGND.n165 214.365
R2550 VGND.n167 VGND.n166 214.365
R2551 VGND.n157 VGND.n155 214.365
R2552 VGND.n157 VGND.n156 214.365
R2553 VGND.n175 VGND.n173 214.365
R2554 VGND.n175 VGND.n174 214.365
R2555 VGND.n1100 VGND.n1099 213.613
R2556 VGND.n1102 VGND.n1101 213.613
R2557 VGND.n1072 VGND.n1070 213.613
R2558 VGND.n1072 VGND.n1071 213.613
R2559 VGND.n1075 VGND.n1073 213.613
R2560 VGND.n1075 VGND.n1074 213.613
R2561 VGND.n1010 VGND.n1008 213.613
R2562 VGND.n1010 VGND.n1009 213.613
R2563 VGND.n1013 VGND.n1011 213.613
R2564 VGND.n1013 VGND.n1012 213.613
R2565 VGND.n1041 VGND.n1039 213.613
R2566 VGND.n1041 VGND.n1040 213.613
R2567 VGND.n1044 VGND.n1042 213.613
R2568 VGND.n1044 VGND.n1043 213.613
R2569 VGND.n3023 VGND.n3022 212.329
R2570 VGND.n3031 VGND.n3 212.329
R2571 VGND.n1114 VGND.t212 211.359
R2572 VGND.n972 VGND.n971 207.965
R2573 VGND.n989 VGND.n969 207.965
R2574 VGND.n102 VGND.n98 207.965
R2575 VGND.n102 VGND.n99 207.965
R2576 VGND.n96 VGND.n94 207.965
R2577 VGND.n96 VGND.n95 207.965
R2578 VGND.n109 VGND.n92 207.965
R2579 VGND.n109 VGND.n93 207.965
R2580 VGND.n2857 VGND.n2853 207.965
R2581 VGND.n2857 VGND.n2854 207.965
R2582 VGND.n2851 VGND.n2849 207.965
R2583 VGND.n2851 VGND.n2850 207.965
R2584 VGND.n2864 VGND.n2847 207.965
R2585 VGND.n2864 VGND.n2848 207.965
R2586 VGND.n2889 VGND.n2885 207.965
R2587 VGND.n2889 VGND.n2886 207.965
R2588 VGND.n2883 VGND.n2881 207.965
R2589 VGND.n2883 VGND.n2882 207.965
R2590 VGND.n2896 VGND.n2879 207.965
R2591 VGND.n2896 VGND.n2880 207.965
R2592 VGND.n71 VGND.n70 207.965
R2593 VGND.n83 VGND.n68 207.965
R2594 VGND.n75 VGND.n73 207.965
R2595 VGND.n988 VGND.n970 207.213
R2596 VGND.n18 VGND.n17 207.213
R2597 VGND.n22 VGND.n16 207.213
R2598 VGND.n47 VGND.n45 207.213
R2599 VGND.n47 VGND.n46 207.213
R2600 VGND.n51 VGND.n43 207.213
R2601 VGND.n51 VGND.n44 207.213
R2602 VGND.n82 VGND.n69 207.213
R2603 VGND.n2931 VGND.n2929 207.213
R2604 VGND.n2931 VGND.n2930 207.213
R2605 VGND.n2935 VGND.n2926 207.213
R2606 VGND.n2935 VGND.n2927 207.213
R2607 VGND.n2971 VGND.n2969 207.213
R2608 VGND.n2971 VGND.n2970 207.213
R2609 VGND.n2975 VGND.n2967 207.213
R2610 VGND.n2975 VGND.n2968 207.213
R2611 VGND.t948 VGND.t2470 203.242
R2612 VGND.t749 VGND.t897 203.242
R2613 VGND.t903 VGND.t1693 203.242
R2614 VGND.t1669 VGND.t921 203.242
R2615 VGND.t996 VGND.t747 203.242
R2616 VGND.t735 VGND.t1002 203.242
R2617 VGND.t924 VGND.t713 203.242
R2618 VGND.t2458 VGND.t966 203.242
R2619 VGND.t975 VGND.t2438 203.242
R2620 VGND.t708 VGND.t1014 203.242
R2621 VGND.t930 VGND.t1652 203.242
R2622 VGND.t2502 VGND.t978 203.242
R2623 VGND.t1017 VGND.t2413 203.242
R2624 VGND.t698 VGND.t1026 203.242
R2625 VGND.t942 VGND.t2491 203.242
R2626 VGND.t2424 VGND.t984 203.242
R2627 VGND VGND.n2656 194.419
R2628 VGND VGND.n2652 194.419
R2629 VGND VGND.n2664 194.419
R2630 VGND VGND.n2648 194.419
R2631 VGND VGND.n2672 194.419
R2632 VGND VGND.n2644 194.419
R2633 VGND VGND.n2680 194.419
R2634 VGND VGND.n2640 194.419
R2635 VGND VGND.n2688 194.419
R2636 VGND VGND.n2636 194.419
R2637 VGND VGND.n2696 194.419
R2638 VGND VGND.n2632 194.419
R2639 VGND VGND.n2704 194.419
R2640 VGND VGND.n2583 194.419
R2641 VGND VGND.n2574 194.419
R2642 VGND.n680 VGND.n679 194.391
R2643 VGND.n1290 VGND.n682 194.391
R2644 VGND.n688 VGND.n686 194.391
R2645 VGND.n726 VGND.n725 194.391
R2646 VGND.n731 VGND.n730 194.391
R2647 VGND.n736 VGND.n735 194.391
R2648 VGND.n741 VGND.n740 194.391
R2649 VGND.n746 VGND.n745 194.391
R2650 VGND.n751 VGND.n750 194.391
R2651 VGND.n756 VGND.n755 194.391
R2652 VGND.n761 VGND.n760 194.391
R2653 VGND.n766 VGND.n765 194.391
R2654 VGND.n771 VGND.n770 194.391
R2655 VGND.n776 VGND.n775 194.391
R2656 VGND.n781 VGND.n780 194.391
R2657 VGND.n1235 VGND.n791 194.391
R2658 VGND.n1228 VGND.n1227 194.391
R2659 VGND.n797 VGND.n796 194.391
R2660 VGND.n1209 VGND.n1208 194.391
R2661 VGND.n1203 VGND.n799 194.391
R2662 VGND.n1196 VGND.n1195 194.391
R2663 VGND.n805 VGND.n804 194.391
R2664 VGND.n1177 VGND.n1176 194.391
R2665 VGND.n1171 VGND.n807 194.391
R2666 VGND.n1164 VGND.n1163 194.391
R2667 VGND.n813 VGND.n812 194.391
R2668 VGND.n1145 VGND.n1144 194.391
R2669 VGND.n1139 VGND.n815 194.391
R2670 VGND.n1132 VGND.n1131 194.391
R2671 VGND.n1129 VGND.n817 194.391
R2672 VGND.n2578 VGND.n2577 194.391
R2673 VGND.n233 VGND.n232 194.391
R2674 VGND.n235 VGND.n234 194.391
R2675 VGND.n2720 VGND.n2719 194.391
R2676 VGND.n2725 VGND.n2724 194.391
R2677 VGND.n2730 VGND.n2729 194.391
R2678 VGND.n2735 VGND.n2734 194.391
R2679 VGND.n2740 VGND.n2739 194.391
R2680 VGND.n2745 VGND.n2744 194.391
R2681 VGND.n2750 VGND.n2749 194.391
R2682 VGND.n2755 VGND.n2754 194.391
R2683 VGND.n2760 VGND.n2759 194.391
R2684 VGND.n2765 VGND.n2764 194.391
R2685 VGND.n2770 VGND.n2769 194.391
R2686 VGND.n2775 VGND.n2774 194.391
R2687 VGND.n2780 VGND.n2779 194.391
R2688 VGND.n230 VGND.n229 194.391
R2689 VGND.n243 VGND.n242 194.391
R2690 VGND.n245 VGND.n244 194.391
R2691 VGND.n2514 VGND.n2513 194.391
R2692 VGND.n2509 VGND.n247 194.391
R2693 VGND.n251 VGND.n249 194.391
R2694 VGND.n2439 VGND.n2438 194.391
R2695 VGND.n2444 VGND.n2443 194.391
R2696 VGND.n2449 VGND.n2448 194.391
R2697 VGND.n2454 VGND.n2453 194.391
R2698 VGND.n2459 VGND.n2458 194.391
R2699 VGND.n2464 VGND.n2463 194.391
R2700 VGND.n2469 VGND.n2468 194.391
R2701 VGND.n2474 VGND.n2473 194.391
R2702 VGND.n2479 VGND.n2478 194.391
R2703 VGND.n2484 VGND.n2483 194.391
R2704 VGND.n2489 VGND.n2488 194.391
R2705 VGND.n183 VGND.n182 194.391
R2706 VGND.n2832 VGND.n185 194.391
R2707 VGND.n371 VGND.n369 194.391
R2708 VGND.n373 VGND.n372 194.391
R2709 VGND.n2172 VGND.n2171 194.391
R2710 VGND.n367 VGND.n366 194.391
R2711 VGND.n2198 VGND.n2197 194.391
R2712 VGND.n359 VGND.n358 194.391
R2713 VGND.n2224 VGND.n2223 194.391
R2714 VGND.n351 VGND.n350 194.391
R2715 VGND.n2250 VGND.n2249 194.391
R2716 VGND.n343 VGND.n342 194.391
R2717 VGND.n2281 VGND.n2280 194.391
R2718 VGND.n2286 VGND.n2285 194.391
R2719 VGND.n2291 VGND.n2290 194.391
R2720 VGND.n335 VGND.n334 194.391
R2721 VGND.n1423 VGND.n1422 194.391
R2722 VGND.n1429 VGND.n1428 194.391
R2723 VGND.n1426 VGND.n1425 194.391
R2724 VGND.n2159 VGND.n2158 194.391
R2725 VGND.n382 VGND.n381 194.391
R2726 VGND.n2185 VGND.n2184 194.391
R2727 VGND.n363 VGND.n362 194.391
R2728 VGND.n2211 VGND.n2210 194.391
R2729 VGND.n355 VGND.n354 194.391
R2730 VGND.n2237 VGND.n2236 194.391
R2731 VGND.n347 VGND.n346 194.391
R2732 VGND.n2263 VGND.n2262 194.391
R2733 VGND.n339 VGND.n338 194.391
R2734 VGND.n2268 VGND.n2267 194.391
R2735 VGND.n2308 VGND.n2307 194.391
R2736 VGND.n2315 VGND.n330 194.391
R2737 VGND.n641 VGND.n640 194.391
R2738 VGND.n1443 VGND.n1442 194.391
R2739 VGND.n637 VGND.n636 194.391
R2740 VGND.n1493 VGND.n1492 194.391
R2741 VGND.n1488 VGND.n1487 194.391
R2742 VGND.n1483 VGND.n1482 194.391
R2743 VGND.n1478 VGND.n1477 194.391
R2744 VGND.n1473 VGND.n1472 194.391
R2745 VGND.n1468 VGND.n1467 194.391
R2746 VGND.n1463 VGND.n1462 194.391
R2747 VGND.n1458 VGND.n1457 194.391
R2748 VGND.n1453 VGND.n1452 194.391
R2749 VGND.n1448 VGND.n1447 194.391
R2750 VGND.n396 VGND.n395 194.391
R2751 VGND.n2136 VGND.n2135 194.391
R2752 VGND.n2131 VGND.n398 194.391
R2753 VGND.n620 VGND.n619 194.391
R2754 VGND.n1505 VGND.n622 194.391
R2755 VGND.n626 VGND.n624 194.391
R2756 VGND.n628 VGND.n627 194.391
R2757 VGND.n1998 VGND.n1997 194.391
R2758 VGND.n434 VGND.n433 194.391
R2759 VGND.n2024 VGND.n2023 194.391
R2760 VGND.n426 VGND.n425 194.391
R2761 VGND.n2050 VGND.n2049 194.391
R2762 VGND.n418 VGND.n417 194.391
R2763 VGND.n2076 VGND.n2075 194.391
R2764 VGND.n410 VGND.n409 194.391
R2765 VGND.n2107 VGND.n2106 194.391
R2766 VGND.n2112 VGND.n2111 194.391
R2767 VGND.n2117 VGND.n2116 194.391
R2768 VGND.n2124 VGND.n401 194.391
R2769 VGND.n647 VGND.n646 194.391
R2770 VGND.n653 VGND.n652 194.391
R2771 VGND.n650 VGND.n649 194.391
R2772 VGND.n1985 VGND.n1984 194.391
R2773 VGND.n438 VGND.n437 194.391
R2774 VGND.n2011 VGND.n2010 194.391
R2775 VGND.n430 VGND.n429 194.391
R2776 VGND.n2037 VGND.n2036 194.391
R2777 VGND.n422 VGND.n421 194.391
R2778 VGND.n2063 VGND.n2062 194.391
R2779 VGND.n414 VGND.n413 194.391
R2780 VGND.n2089 VGND.n2088 194.391
R2781 VGND.n406 VGND.n405 194.391
R2782 VGND.n2094 VGND.n2093 194.391
R2783 VGND.n2333 VGND.n2332 194.391
R2784 VGND.n2340 VGND.n319 194.391
R2785 VGND.n663 VGND.n662 194.391
R2786 VGND.n960 VGND.n959 194.391
R2787 VGND.n955 VGND.n954 194.391
R2788 VGND.n950 VGND.n949 194.391
R2789 VGND.n945 VGND.n944 194.391
R2790 VGND.n940 VGND.n939 194.391
R2791 VGND.n935 VGND.n934 194.391
R2792 VGND.n930 VGND.n929 194.391
R2793 VGND.n925 VGND.n924 194.391
R2794 VGND.n920 VGND.n919 194.391
R2795 VGND.n915 VGND.n914 194.391
R2796 VGND.n910 VGND.n909 194.391
R2797 VGND.n905 VGND.n904 194.391
R2798 VGND.n452 VGND.n451 194.391
R2799 VGND.n1962 VGND.n1961 194.391
R2800 VGND.n1957 VGND.n454 194.391
R2801 VGND.n672 VGND.n671 194.391
R2802 VGND.n1396 VGND.n1395 194.391
R2803 VGND.n1401 VGND.n1400 194.391
R2804 VGND.n669 VGND.n668 194.391
R2805 VGND.n1824 VGND.n1823 194.391
R2806 VGND.n490 VGND.n489 194.391
R2807 VGND.n1850 VGND.n1849 194.391
R2808 VGND.n482 VGND.n481 194.391
R2809 VGND.n1876 VGND.n1875 194.391
R2810 VGND.n474 VGND.n473 194.391
R2811 VGND.n1902 VGND.n1901 194.391
R2812 VGND.n466 VGND.n465 194.391
R2813 VGND.n1933 VGND.n1932 194.391
R2814 VGND.n1938 VGND.n1937 194.391
R2815 VGND.n1943 VGND.n1942 194.391
R2816 VGND.n1950 VGND.n457 194.391
R2817 VGND.n1375 VGND.n1374 194.391
R2818 VGND.n1381 VGND.n1380 194.391
R2819 VGND.n1378 VGND.n1377 194.391
R2820 VGND.n1811 VGND.n1810 194.391
R2821 VGND.n494 VGND.n493 194.391
R2822 VGND.n1837 VGND.n1836 194.391
R2823 VGND.n486 VGND.n485 194.391
R2824 VGND.n1863 VGND.n1862 194.391
R2825 VGND.n478 VGND.n477 194.391
R2826 VGND.n1889 VGND.n1888 194.391
R2827 VGND.n470 VGND.n469 194.391
R2828 VGND.n1915 VGND.n1914 194.391
R2829 VGND.n462 VGND.n461 194.391
R2830 VGND.n1920 VGND.n1919 194.391
R2831 VGND.n2358 VGND.n2357 194.391
R2832 VGND.n2365 VGND.n307 194.391
R2833 VGND.n1307 VGND.n1306 194.391
R2834 VGND.n1313 VGND.n1312 194.391
R2835 VGND.n1310 VGND.n1309 194.391
R2836 VGND.n1363 VGND.n1362 194.391
R2837 VGND.n1358 VGND.n1357 194.391
R2838 VGND.n1353 VGND.n1352 194.391
R2839 VGND.n1348 VGND.n1347 194.391
R2840 VGND.n1343 VGND.n1342 194.391
R2841 VGND.n1338 VGND.n1337 194.391
R2842 VGND.n1333 VGND.n1332 194.391
R2843 VGND.n1328 VGND.n1327 194.391
R2844 VGND.n1323 VGND.n1322 194.391
R2845 VGND.n1318 VGND.n1317 194.391
R2846 VGND.n508 VGND.n507 194.391
R2847 VGND.n1788 VGND.n1787 194.391
R2848 VGND.n1783 VGND.n510 194.391
R2849 VGND.n576 VGND.n575 194.391
R2850 VGND.n1518 VGND.n1517 194.391
R2851 VGND.n1523 VGND.n1522 194.391
R2852 VGND.n580 VGND.n579 194.391
R2853 VGND.n1650 VGND.n1649 194.391
R2854 VGND.n546 VGND.n545 194.391
R2855 VGND.n1676 VGND.n1675 194.391
R2856 VGND.n538 VGND.n537 194.391
R2857 VGND.n1702 VGND.n1701 194.391
R2858 VGND.n530 VGND.n529 194.391
R2859 VGND.n1728 VGND.n1727 194.391
R2860 VGND.n522 VGND.n521 194.391
R2861 VGND.n1759 VGND.n1758 194.391
R2862 VGND.n1764 VGND.n1763 194.391
R2863 VGND.n1769 VGND.n1768 194.391
R2864 VGND.n1776 VGND.n513 194.391
R2865 VGND.n572 VGND.n571 194.391
R2866 VGND.n1538 VGND.n1537 194.391
R2867 VGND.n569 VGND.n568 194.391
R2868 VGND.n1637 VGND.n1636 194.391
R2869 VGND.n550 VGND.n549 194.391
R2870 VGND.n1663 VGND.n1662 194.391
R2871 VGND.n542 VGND.n541 194.391
R2872 VGND.n1689 VGND.n1688 194.391
R2873 VGND.n534 VGND.n533 194.391
R2874 VGND.n1715 VGND.n1714 194.391
R2875 VGND.n526 VGND.n525 194.391
R2876 VGND.n1741 VGND.n1740 194.391
R2877 VGND.n518 VGND.n517 194.391
R2878 VGND.n1746 VGND.n1745 194.391
R2879 VGND.n2383 VGND.n2382 194.391
R2880 VGND.n2390 VGND.n294 194.391
R2881 VGND.n675 VGND.n674 194.391
R2882 VGND.n677 VGND.n676 194.391
R2883 VGND.n1551 VGND.n1550 194.391
R2884 VGND.n1556 VGND.n1555 194.391
R2885 VGND.n1561 VGND.n1560 194.391
R2886 VGND.n1566 VGND.n1565 194.391
R2887 VGND.n1571 VGND.n1570 194.391
R2888 VGND.n1576 VGND.n1575 194.391
R2889 VGND.n1581 VGND.n1580 194.391
R2890 VGND.n1586 VGND.n1585 194.391
R2891 VGND.n1591 VGND.n1590 194.391
R2892 VGND.n1596 VGND.n1595 194.391
R2893 VGND.n1601 VGND.n1600 194.391
R2894 VGND.n564 VGND.n563 194.391
R2895 VGND.n1614 VGND.n1613 194.391
R2896 VGND.n1609 VGND.n1605 194.391
R2897 VGND.n829 VGND.n828 194.391
R2898 VGND.n836 VGND.n835 194.391
R2899 VGND.n841 VGND.n840 194.391
R2900 VGND.n833 VGND.n832 194.391
R2901 VGND.n891 VGND.n890 194.391
R2902 VGND.n886 VGND.n885 194.391
R2903 VGND.n881 VGND.n880 194.391
R2904 VGND.n876 VGND.n875 194.391
R2905 VGND.n871 VGND.n870 194.391
R2906 VGND.n866 VGND.n865 194.391
R2907 VGND.n861 VGND.n860 194.391
R2908 VGND.n856 VGND.n855 194.391
R2909 VGND.n851 VGND.n850 194.391
R2910 VGND.n846 VGND.n845 194.391
R2911 VGND.n2403 VGND.n2402 194.391
R2912 VGND.n2410 VGND.n282 194.391
R2913 VGND.n819 VGND.n818 194.391
R2914 VGND.n722 VGND.n721 194.391
R2915 VGND.n3025 VGND.n3024 176.941
R2916 VGND.n9 VGND.n8 176.941
R2917 VGND.n2568 VGND.n2567 161.308
R2918 VGND.n2565 VGND.n2564 161.308
R2919 VGND.n2562 VGND.n2561 161.308
R2920 VGND.n2559 VGND.n2558 161.308
R2921 VGND.n2556 VGND.n2555 161.308
R2922 VGND.n2553 VGND.n2552 161.308
R2923 VGND.n2550 VGND.n2549 161.308
R2924 VGND.n2547 VGND.n2546 161.308
R2925 VGND.n2544 VGND.n2543 161.308
R2926 VGND.n2541 VGND.n2540 161.308
R2927 VGND.n2538 VGND.n2537 161.308
R2928 VGND.n2535 VGND.n2534 161.308
R2929 VGND.n2532 VGND.n2531 161.308
R2930 VGND.n2529 VGND.n2528 161.308
R2931 VGND.n2526 VGND.n2525 161.308
R2932 VGND.n2567 VGND.t2696 159.978
R2933 VGND.n2564 VGND.t2699 159.978
R2934 VGND.n2561 VGND.t2694 159.978
R2935 VGND.n2558 VGND.t2690 159.978
R2936 VGND.n2555 VGND.t2695 159.978
R2937 VGND.n2552 VGND.t2703 159.978
R2938 VGND.n2549 VGND.t2698 159.978
R2939 VGND.n2546 VGND.t2692 159.978
R2940 VGND.n2543 VGND.t2689 159.978
R2941 VGND.n2540 VGND.t2691 159.978
R2942 VGND.n2537 VGND.t2702 159.978
R2943 VGND.n2534 VGND.t2693 159.978
R2944 VGND.n2531 VGND.t2701 159.978
R2945 VGND.n2528 VGND.t2697 159.978
R2946 VGND.n2525 VGND.t2705 159.978
R2947 VGND.n1000 VGND.t676 159.315
R2948 VGND.n2917 VGND.t1375 159.315
R2949 VGND.n1092 VGND.t643 158.361
R2950 VGND.n2987 VGND.t372 158.361
R2951 VGND.n902 VGND.t674 157.291
R2952 VGND.n2915 VGND.t1373 157.291
R2953 VGND.n586 VGND.t1336 156.915
R2954 VGND.n2877 VGND.t1581 156.915
R2955 VGND.n586 VGND.t1334 156.915
R2956 VGND.n2877 VGND.t1582 156.915
R2957 VGND.n588 VGND.t1393 154.131
R2958 VGND.n588 VGND.t2605 154.131
R2959 VGND.n1000 VGND.t2525 154.131
R2960 VGND.n1003 VGND.t1621 154.131
R2961 VGND.n2901 VGND.t1769 154.131
R2962 VGND.n2901 VGND.t1635 154.131
R2963 VGND.n2917 VGND.t2647 154.131
R2964 VGND.n2947 VGND.t1913 154.131
R2965 VGND.n122 VGND.t1332 153.631
R2966 VGND.n1030 VGND.t843 153.631
R2967 VGND.n1061 VGND.t1439 153.631
R2968 VGND.n2869 VGND.t1579 153.631
R2969 VGND.n2949 VGND.t1530 153.631
R2970 VGND.n2954 VGND.t2186 153.631
R2971 VGND.n1031 VGND.t1126 152.757
R2972 VGND.n2950 VGND.t281 152.757
R2973 VGND.n995 VGND.t1330 152.381
R2974 VGND.n65 VGND.t1586 152.381
R2975 VGND.n965 VGND.n964 152.174
R2976 VGND.n153 VGND.t1335 150.922
R2977 VGND.n153 VGND.t1328 150.922
R2978 VGND.n90 VGND.t1589 150.922
R2979 VGND.n90 VGND.t1584 150.922
R2980 VGND.n120 VGND.t327 150.922
R2981 VGND.n585 VGND.t1395 150.922
R2982 VGND.n152 VGND.t209 150.922
R2983 VGND.n89 VGND.t1977 150.922
R2984 VGND.n2844 VGND.t186 150.922
R2985 VGND.n2876 VGND.t257 150.922
R2986 VGND.n120 VGND.t105 150.922
R2987 VGND.n585 VGND.t288 150.922
R2988 VGND.n152 VGND.t2553 150.922
R2989 VGND.n89 VGND.t1559 150.922
R2990 VGND.n2844 VGND.t1641 150.922
R2991 VGND.n2876 VGND.t2651 150.922
R2992 VGND.n121 VGND.t1331 147.411
R2993 VGND.n1062 VGND.t1299 147.411
R2994 VGND.n2868 VGND.t1588 147.411
R2995 VGND.n2955 VGND.t1252 147.411
R2996 VGND.n903 VGND.t221 146.964
R2997 VGND.n88 VGND.t1744 146.964
R2998 VGND.n5 VGND.n3 146.25
R2999 VGND.n7 VGND.n5 146.25
R3000 VGND.n6 VGND.n4 146.25
R3001 VGND.n3017 VGND.n6 146.25
R3002 VGND.n3023 VGND.n3019 146.25
R3003 VGND.n3019 VGND.n7 146.25
R3004 VGND.n3026 VGND.n3020 146.25
R3005 VGND.n3020 VGND.n3017 146.25
R3006 VGND.n2567 VGND.t932 143.911
R3007 VGND.n2564 VGND.t1007 143.911
R3008 VGND.n2561 VGND.t914 143.911
R3009 VGND.n2558 VGND.t956 143.911
R3010 VGND.n2555 VGND.t1028 143.911
R3011 VGND.n2552 VGND.t935 143.911
R3012 VGND.n2549 VGND.t908 143.911
R3013 VGND.n2546 VGND.t950 143.911
R3014 VGND.n2543 VGND.t962 143.911
R3015 VGND.n2540 VGND.t890 143.911
R3016 VGND.n2537 VGND.t986 143.911
R3017 VGND.n2534 VGND.t917 143.911
R3018 VGND.n2531 VGND.t989 143.911
R3019 VGND.n2528 VGND.t1019 143.911
R3020 VGND.n2525 VGND.t959 143.911
R3021 VGND.n1516 VGND.n582 143.478
R3022 VGND VGND.t1261 142.089
R3023 VGND.n826 VGND.t947 119.309
R3024 VGND.n789 VGND.t983 119.309
R3025 VGND.n2589 VGND.t980 119.309
R3026 VGND.n2586 VGND.t944 119.309
R3027 VGND.n2572 VGND.t893 119.309
R3028 VGND.n2585 VGND.t899 119.309
R3029 VGND.n2624 VGND.t905 119.309
R3030 VGND.n2621 VGND.t992 119.309
R3031 VGND.n2618 VGND.t998 119.309
R3032 VGND.n2615 VGND.t911 119.309
R3033 VGND.n2612 VGND.t953 119.309
R3034 VGND.n2609 VGND.t968 119.309
R3035 VGND.n2606 VGND.t1004 119.309
R3036 VGND.n2603 VGND.t926 119.309
R3037 VGND.n2600 VGND.t971 119.309
R3038 VGND.n2597 VGND.t1010 119.309
R3039 VGND.n2594 VGND.t1022 119.309
R3040 VGND.n2591 VGND.t938 119.309
R3041 VGND.n823 VGND.t896 119.309
R3042 VGND.n820 VGND.t902 119.309
R3043 VGND.n1140 VGND.t920 119.309
R3044 VGND.n811 VGND.t995 119.309
R3045 VGND.n809 VGND.t1001 119.309
R3046 VGND.n1155 VGND.t923 119.309
R3047 VGND.n1172 VGND.t965 119.309
R3048 VGND.n803 VGND.t974 119.309
R3049 VGND.n801 VGND.t1013 119.309
R3050 VGND.n1187 VGND.t929 119.309
R3051 VGND.n1204 VGND.t977 119.309
R3052 VGND.n795 VGND.t1016 119.309
R3053 VGND.n793 VGND.t1025 119.309
R3054 VGND.n1219 VGND.t941 119.309
R3055 VGND.t755 VGND.t948 110.535
R3056 VGND.t1113 VGND.t1701 110.535
R3057 VGND.t897 VGND.t1695 110.535
R3058 VGND.t2482 VGND.t1516 110.535
R3059 VGND.t2474 VGND.t903 110.535
R3060 VGND.t1876 VGND.t2467 110.535
R3061 VGND.t921 VGND.t2452 110.535
R3062 VGND.t731 VGND.t1787 110.535
R3063 VGND.t743 VGND.t996 110.535
R3064 VGND.t2536 VGND.t1689 110.535
R3065 VGND.t1002 VGND.t1673 110.535
R3066 VGND.t2455 VGND.t1622 110.535
R3067 VGND.t1660 VGND.t924 110.535
R3068 VGND.t2 VGND.t746 110.535
R3069 VGND.t966 VGND.t737 110.535
R3070 VGND.t721 VGND.t1325 110.535
R3071 VGND.t715 VGND.t975 110.535
R3072 VGND.t1534 VGND.t1662 110.535
R3073 VGND.t1014 VGND.t1675 110.535
R3074 VGND.t2456 VGND.t2521 110.535
R3075 VGND.t2440 VGND.t930 110.535
R3076 VGND.t846 VGND.t718 110.535
R3077 VGND.t978 VGND.t2431 110.535
R3078 VGND.t706 VGND.t0 110.535
R3079 VGND.t1656 VGND.t1017 110.535
R3080 VGND.t1303 VGND.t1649 110.535
R3081 VGND.t1026 VGND.t1644 110.535
R3082 VGND.t2433 VGND.t2606 110.535
R3083 VGND.t2483 VGND.t942 110.535
R3084 VGND.t887 VGND.t2412 110.535
R3085 VGND.t984 VGND.t702 110.535
R3086 VGND.t1646 VGND.t1612 110.535
R3087 VGND.t212 VGND.t222 92.4699
R3088 VGND.t222 VGND.t219 92.4699
R3089 VGND.t219 VGND.t223 92.4699
R3090 VGND.t223 VGND.t440 92.4699
R3091 VGND.t440 VGND.t449 92.4699
R3092 VGND.t449 VGND.t502 92.4699
R3093 VGND.t502 VGND.t408 92.4699
R3094 VGND.n3025 VGND.t2700 88.3562
R3095 VGND.n8 VGND.t2704 88.3562
R3096 VGND VGND.n582 80.9529
R3097 VGND VGND.n582 75.1009
R3098 VGND.n1295 VGND 74.8566
R3099 VGND.t408 VGND 70.4533
R3100 VGND.n3026 VGND.n3025 67.3887
R3101 VGND.n8 VGND.n4 67.3887
R3102 VGND.n151 VGND 58.8055
R3103 VGND.n1510 VGND 58.8055
R3104 VGND.n1512 VGND 58.8055
R3105 VGND.n1514 VGND 58.8055
R3106 VGND.n2837 VGND 58.8055
R3107 VGND.n10 VGND.n9 53.1823
R3108 VGND.t1197 VGND.n10 53.1823
R3109 VGND.n3030 VGND.n3029 53.1823
R3110 VGND.n3029 VGND.t1197 53.1823
R3111 VGND.n3028 VGND.n3027 53.1823
R3112 VGND.t1197 VGND.n3028 53.1823
R3113 VGND.n3024 VGND.n3018 53.1823
R3114 VGND.t1197 VGND.n3018 53.1823
R3115 VGND.t220 VGND.t438 50.5752
R3116 VGND.t217 VGND.t447 50.5752
R3117 VGND.t215 VGND.t592 50.5752
R3118 VGND.t213 VGND.t2358 50.5752
R3119 VGND.t1751 VGND.t1263 50.5752
R3120 VGND.t1747 VGND.t613 50.5752
R3121 VGND.t1741 VGND.t671 50.5752
R3122 VGND.t1743 VGND.t493 50.5752
R3123 VGND VGND.n18 43.2063
R3124 VGND VGND.n47 43.2063
R3125 VGND VGND.n2931 43.2063
R3126 VGND VGND.n2971 43.2063
R3127 VGND.n679 VGND.t720 34.8005
R3128 VGND.n679 VGND.t1666 34.8005
R3129 VGND.n682 VGND.t1664 34.8005
R3130 VGND.n682 VGND.t2446 34.8005
R3131 VGND.n686 VGND.t2443 34.8005
R3132 VGND.n686 VGND.t723 34.8005
R3133 VGND.n725 VGND.t2421 34.8005
R3134 VGND.n725 VGND.t701 34.8005
R3135 VGND.n730 VGND.t1659 34.8005
R3136 VGND.n730 VGND.t1655 34.8005
R3137 VGND.n735 VGND.t1648 34.8005
R3138 VGND.n735 VGND.t2427 34.8005
R3139 VGND.n740 VGND.t2490 34.8005
R3140 VGND.n740 VGND.t2416 34.8005
R3141 VGND.n745 VGND.t705 34.8005
R3142 VGND.n745 VGND.t1651 34.8005
R3143 VGND.n750 VGND.t684 34.8005
R3144 VGND.n750 VGND.t2494 34.8005
R3145 VGND.n755 VGND.t2486 34.8005
R3146 VGND.n755 VGND.t2429 34.8005
R3147 VGND.n760 VGND.t765 34.8005
R3148 VGND.n760 VGND.t688 34.8005
R3149 VGND.n765 VGND.t752 34.8005
R3150 VGND.n765 VGND.t1699 34.8005
R3151 VGND.n770 VGND.t1683 34.8005
R3152 VGND.n770 VGND.t2411 34.8005
R3153 VGND.n775 VGND.t2469 34.8005
R3154 VGND.n775 VGND.t754 34.8005
R3155 VGND.n780 VGND.t734 34.8005
R3156 VGND.n780 VGND.t729 34.8005
R3157 VGND.n791 VGND.t2425 34.8005
R3158 VGND.n791 VGND.t703 34.8005
R3159 VGND.n1227 VGND.t2492 34.8005
R3160 VGND.n1227 VGND.t2484 34.8005
R3161 VGND.n796 VGND.t699 34.8005
R3162 VGND.n796 VGND.t1645 34.8005
R3163 VGND.n1208 VGND.t2414 34.8005
R3164 VGND.n1208 VGND.t1657 34.8005
R3165 VGND.n799 VGND.t2503 34.8005
R3166 VGND.n799 VGND.t2432 34.8005
R3167 VGND.n1195 VGND.t1653 34.8005
R3168 VGND.n1195 VGND.t2441 34.8005
R3169 VGND.n804 VGND.t709 34.8005
R3170 VGND.n804 VGND.t1676 34.8005
R3171 VGND.n1176 VGND.t2439 34.8005
R3172 VGND.n1176 VGND.t716 34.8005
R3173 VGND.n807 VGND.t2459 34.8005
R3174 VGND.n807 VGND.t738 34.8005
R3175 VGND.n1163 VGND.t714 34.8005
R3176 VGND.n1163 VGND.t1661 34.8005
R3177 VGND.n812 VGND.t736 34.8005
R3178 VGND.n812 VGND.t1674 34.8005
R3179 VGND.n1144 VGND.t748 34.8005
R3180 VGND.n1144 VGND.t744 34.8005
R3181 VGND.n815 VGND.t1670 34.8005
R3182 VGND.n815 VGND.t2453 34.8005
R3183 VGND.n1131 VGND.t1694 34.8005
R3184 VGND.n1131 VGND.t2475 34.8005
R3185 VGND.n817 VGND.t750 34.8005
R3186 VGND.n817 VGND.t1696 34.8005
R3187 VGND.n2577 VGND.t2419 34.8005
R3188 VGND.n2577 VGND.t697 34.8005
R3189 VGND.n2656 VGND.t725 34.8005
R3190 VGND.n2656 VGND.t1672 34.8005
R3191 VGND.n2652 VGND.t2437 34.8005
R3192 VGND.n2652 VGND.t2435 34.8005
R3193 VGND.n2664 VGND.t1668 34.8005
R3194 VGND.n2664 VGND.t2451 34.8005
R3195 VGND.n2648 VGND.t711 34.8005
R3196 VGND.n2648 VGND.t2463 34.8005
R3197 VGND.n2672 VGND.t2449 34.8005
R3198 VGND.n2672 VGND.t727 34.8005
R3199 VGND.n2644 VGND.t2461 34.8005
R3200 VGND.n2644 VGND.t742 34.8005
R3201 VGND.n2680 VGND.t1681 34.8005
R3202 VGND.n2680 VGND.t2481 34.8005
R3203 VGND.n2640 VGND.t740 34.8005
R3204 VGND.n2640 VGND.t1687 34.8005
R3205 VGND.n2688 VGND.t763 34.8005
R3206 VGND.n2688 VGND.t686 34.8005
R3207 VGND.n2636 VGND.t1685 34.8005
R3208 VGND.n2636 VGND.t2465 34.8005
R3209 VGND.n2696 VGND.t682 34.8005
R3210 VGND.n2696 VGND.t2479 34.8005
R3211 VGND.n2632 VGND.t693 34.8005
R3212 VGND.n2632 VGND.t690 34.8005
R3213 VGND.n2704 VGND.t2477 34.8005
R3214 VGND.n2704 VGND.t759 34.8005
R3215 VGND.n2583 VGND.t2499 34.8005
R3216 VGND.n2583 VGND.t2423 34.8005
R3217 VGND.n2574 VGND.t695 34.8005
R3218 VGND.n2574 VGND.t2501 34.8005
R3219 VGND.n232 VGND.t934 34.8005
R3220 VGND.n232 VGND.t2090 34.8005
R3221 VGND.n234 VGND.t1149 34.8005
R3222 VGND.n234 VGND.t1377 34.8005
R3223 VGND.n2719 VGND.t2259 34.8005
R3224 VGND.n2719 VGND.t1478 34.8005
R3225 VGND.n2724 VGND.t130 34.8005
R3226 VGND.n2724 VGND.t2096 34.8005
R3227 VGND.n2729 VGND.t1389 34.8005
R3228 VGND.n2729 VGND.t2088 34.8005
R3229 VGND.n2734 VGND.t1968 34.8005
R3230 VGND.n2734 VGND.t1488 34.8005
R3231 VGND.n2739 VGND.t162 34.8005
R3232 VGND.n2739 VGND.t1486 34.8005
R3233 VGND.n2744 VGND.t2408 34.8005
R3234 VGND.n2744 VGND.t2086 34.8005
R3235 VGND.n2749 VGND.t1756 34.8005
R3236 VGND.n2749 VGND.t1381 34.8005
R3237 VGND.n2754 VGND.t472 34.8005
R3238 VGND.n2754 VGND.t1490 34.8005
R3239 VGND.n2759 VGND.t538 34.8005
R3240 VGND.n2759 VGND.t2094 34.8005
R3241 VGND.n2764 VGND.t877 34.8005
R3242 VGND.n2764 VGND.t2092 34.8005
R3243 VGND.n2769 VGND.t1863 34.8005
R3244 VGND.n2769 VGND.t1484 34.8005
R3245 VGND.n2774 VGND.t306 34.8005
R3246 VGND.n2774 VGND.t1482 34.8005
R3247 VGND.n2779 VGND.t1807 34.8005
R3248 VGND.n2779 VGND.t1480 34.8005
R3249 VGND.n229 VGND.t1508 34.8005
R3250 VGND.n229 VGND.t1379 34.8005
R3251 VGND.n242 VGND.t1009 34.8005
R3252 VGND.n242 VGND.t2320 34.8005
R3253 VGND.n244 VGND.t829 34.8005
R3254 VGND.n244 VGND.t2333 34.8005
R3255 VGND.n2513 VGND.t2681 34.8005
R3256 VGND.n2513 VGND.t1595 34.8005
R3257 VGND.n247 VGND.t771 34.8005
R3258 VGND.n247 VGND.t1593 34.8005
R3259 VGND.n249 VGND.t601 34.8005
R3260 VGND.n249 VGND.t2318 34.8005
R3261 VGND.n2438 VGND.t649 34.8005
R3262 VGND.n2438 VGND.t2329 34.8005
R3263 VGND.n2443 VGND.t1539 34.8005
R3264 VGND.n2443 VGND.t2327 34.8005
R3265 VGND.n2448 VGND.t666 34.8005
R3266 VGND.n2448 VGND.t2316 34.8005
R3267 VGND.n2453 VGND.t2688 34.8005
R3268 VGND.n2453 VGND.t2314 34.8005
R3269 VGND.n2458 VGND.t1135 34.8005
R3270 VGND.n2458 VGND.t2331 34.8005
R3271 VGND.n2463 VGND.t521 34.8005
R3272 VGND.n2463 VGND.t2076 34.8005
R3273 VGND.n2468 VGND.t1919 34.8005
R3274 VGND.n2468 VGND.t2074 34.8005
R3275 VGND.n2473 VGND.t1833 34.8005
R3276 VGND.n2473 VGND.t2325 34.8005
R3277 VGND.n2478 VGND.t2197 34.8005
R3278 VGND.n2478 VGND.t2323 34.8005
R3279 VGND.n2483 VGND.t1827 34.8005
R3280 VGND.n2483 VGND.t1597 34.8005
R3281 VGND.n2488 VGND.t92 34.8005
R3282 VGND.n2488 VGND.t2312 34.8005
R3283 VGND.n182 VGND.t916 34.8005
R3284 VGND.n182 VGND.t1285 34.8005
R3285 VGND.n185 VGND.t1344 34.8005
R3286 VGND.n185 VGND.t1626 34.8005
R3287 VGND.n369 VGND.t1995 34.8005
R3288 VGND.n369 VGND.t1609 34.8005
R3289 VGND.n372 VGND.t97 34.8005
R3290 VGND.n372 VGND.t1607 34.8005
R3291 VGND.n2171 VGND.t1165 34.8005
R3292 VGND.n2171 VGND.t1283 34.8005
R3293 VGND.n366 VGND.t1711 34.8005
R3294 VGND.n366 VGND.t2004 34.8005
R3295 VGND.n2197 VGND.t1563 34.8005
R3296 VGND.n2197 VGND.t2002 34.8005
R3297 VGND.n358 VGND.t1312 34.8005
R3298 VGND.n358 VGND.t1281 34.8005
R3299 VGND.n2223 VGND.t376 34.8005
R3300 VGND.n2223 VGND.t1630 34.8005
R3301 VGND.n350 VGND.t119 34.8005
R3302 VGND.n350 VGND.t1624 34.8005
R3303 VGND.n2249 VGND.t29 34.8005
R3304 VGND.n2249 VGND.t1289 34.8005
R3305 VGND.n342 VGND.t2046 34.8005
R3306 VGND.n342 VGND.t1287 34.8005
R3307 VGND.n2280 VGND.t2613 34.8005
R3308 VGND.n2280 VGND.t2000 34.8005
R3309 VGND.n2285 VGND.t394 34.8005
R3310 VGND.n2285 VGND.t1865 34.8005
R3311 VGND.n2290 VGND.t110 34.8005
R3312 VGND.n2290 VGND.t1611 34.8005
R3313 VGND.n334 VGND.t1515 34.8005
R3314 VGND.n334 VGND.t1628 34.8005
R3315 VGND.n1422 VGND.t958 34.8005
R3316 VGND.n1422 VGND.t274 34.8005
R3317 VGND.n1428 VGND.t1932 34.8005
R3318 VGND.n1428 VGND.t2218 34.8005
R3319 VGND.n1425 VGND.t2165 34.8005
R3320 VGND.n1425 VGND.t1435 34.8005
R3321 VGND.n2158 VGND.t152 34.8005
R3322 VGND.n2158 VGND.t1433 34.8005
R3323 VGND.n381 VGND.t67 34.8005
R3324 VGND.n381 VGND.t272 34.8005
R3325 VGND.n2184 VGND.t2084 34.8005
R3326 VGND.n2184 VGND.t2214 34.8005
R3327 VGND.n362 VGND.t137 34.8005
R3328 VGND.n362 VGND.t2212 34.8005
R3329 VGND.n2210 VGND.t2400 34.8005
R3330 VGND.n2210 VGND.t270 34.8005
R3331 VGND.n354 VGND.t1069 34.8005
R3332 VGND.n354 VGND.t2560 34.8005
R3333 VGND.n2236 VGND.t1158 34.8005
R3334 VGND.n2236 VGND.t2216 34.8005
R3335 VGND.n346 VGND.t564 34.8005
R3336 VGND.n346 VGND.t278 34.8005
R3337 VGND.n2262 VGND.t1446 34.8005
R3338 VGND.n2262 VGND.t276 34.8005
R3339 VGND.n338 VGND.t173 34.8005
R3340 VGND.n338 VGND.t2210 34.8005
R3341 VGND.n2267 VGND.t1794 34.8005
R3342 VGND.n2267 VGND.t2208 34.8005
R3343 VGND.n2307 VGND.t1816 34.8005
R3344 VGND.n2307 VGND.t1437 34.8005
R3345 VGND.n330 VGND.t2132 34.8005
R3346 VGND.n330 VGND.t2558 34.8005
R3347 VGND.n640 VGND.t1030 34.8005
R3348 VGND.n640 VGND.t2604 34.8005
R3349 VGND.n1442 VGND.t467 34.8005
R3350 VGND.n1442 VGND.t2106 34.8005
R3351 VGND.n636 VGND.t838 34.8005
R3352 VGND.n636 VGND.t2250 34.8005
R3353 VGND.n1492 VGND.t813 34.8005
R3354 VGND.n1492 VGND.t1549 34.8005
R3355 VGND.n1487 VGND.t2515 34.8005
R3356 VGND.n1487 VGND.t2602 34.8005
R3357 VGND.n1482 VGND.t2148 34.8005
R3358 VGND.n1482 VGND.t2102 34.8005
R3359 VGND.n1477 VGND.t1906 34.8005
R3360 VGND.n1477 VGND.t2100 34.8005
R3361 VGND.n1472 VGND.t1319 34.8005
R3362 VGND.n1472 VGND.t2600 34.8005
R3363 VGND.n1467 VGND.t369 34.8005
R3364 VGND.n1467 VGND.t2598 34.8005
R3365 VGND.n1462 VGND.t842 34.8005
R3366 VGND.n1462 VGND.t2104 34.8005
R3367 VGND.n1457 VGND.t516 34.8005
R3368 VGND.n1457 VGND.t1547 34.8005
R3369 VGND.n1452 VGND.t2533 34.8005
R3370 VGND.n1452 VGND.t1545 34.8005
R3371 VGND.n1447 VGND.t2590 34.8005
R3372 VGND.n1447 VGND.t2098 34.8005
R3373 VGND.n395 VGND.t401 34.8005
R3374 VGND.n395 VGND.t2254 34.8005
R3375 VGND.n2135 VGND.t1112 34.8005
R3376 VGND.n2135 VGND.t2252 34.8005
R3377 VGND.n398 VGND.t2116 34.8005
R3378 VGND.n398 VGND.t2108 34.8005
R3379 VGND.n619 VGND.t937 34.8005
R3380 VGND.n619 VGND.t2267 34.8005
R3381 VGND.n622 VGND.t1147 34.8005
R3382 VGND.n622 VGND.t1569 34.8005
R3383 VGND.n624 VGND.t2257 34.8005
R3384 VGND.n624 VGND.t2281 34.8005
R3385 VGND.n627 VGND.t127 34.8005
R3386 VGND.n627 VGND.t2273 34.8005
R3387 VGND.n1997 VGND.t1387 34.8005
R3388 VGND.n1997 VGND.t2265 34.8005
R3389 VGND.n433 VGND.t1966 34.8005
R3390 VGND.n433 VGND.t2291 34.8005
R3391 VGND.n2023 VGND.t160 34.8005
R3392 VGND.n2023 VGND.t2289 34.8005
R3393 VGND.n425 VGND.t2406 34.8005
R3394 VGND.n425 VGND.t2263 34.8005
R3395 VGND.n2049 VGND.t1754 34.8005
R3396 VGND.n2049 VGND.t1573 34.8005
R3397 VGND.n417 VGND.t470 34.8005
R3398 VGND.n417 VGND.t2293 34.8005
R3399 VGND.n2075 VGND.t535 34.8005
R3400 VGND.n2075 VGND.t2271 34.8005
R3401 VGND.n409 VGND.t875 34.8005
R3402 VGND.n409 VGND.t2269 34.8005
R3403 VGND.n2106 VGND.t1860 34.8005
R3404 VGND.n2106 VGND.t2287 34.8005
R3405 VGND.n2111 VGND.t304 34.8005
R3406 VGND.n2111 VGND.t2285 34.8005
R3407 VGND.n2116 VGND.t1818 34.8005
R3408 VGND.n2116 VGND.t2283 34.8005
R3409 VGND.n401 VGND.t1506 34.8005
R3410 VGND.n401 VGND.t1571 34.8005
R3411 VGND.n646 VGND.t910 34.8005
R3412 VGND.n646 VGND.t481 34.8005
R3413 VGND.n652 VGND.t1346 34.8005
R3414 VGND.n652 VGND.t632 34.8005
R3415 VGND.n649 VGND.t1997 34.8005
R3416 VGND.n649 VGND.t489 34.8005
R3417 VGND.n1984 VGND.t95 34.8005
R3418 VGND.n1984 VGND.t487 34.8005
R3419 VGND.n437 VGND.t1167 34.8005
R3420 VGND.n437 VGND.t479 34.8005
R3421 VGND.n2010 VGND.t1713 34.8005
R3422 VGND.n2010 VGND.t628 34.8005
R3423 VGND.n429 VGND.t1565 34.8005
R3424 VGND.n429 VGND.t626 34.8005
R3425 VGND.n2036 VGND.t1314 34.8005
R3426 VGND.n2036 VGND.t477 34.8005
R3427 VGND.n421 VGND.t378 34.8005
R3428 VGND.n421 VGND.t636 34.8005
R3429 VGND.n2062 VGND.t121 34.8005
R3430 VGND.n2062 VGND.t630 34.8005
R3431 VGND.n413 VGND.t31 34.8005
R3432 VGND.n413 VGND.t485 34.8005
R3433 VGND.n2088 VGND.t2048 34.8005
R3434 VGND.n2088 VGND.t483 34.8005
R3435 VGND.n405 VGND.t2615 34.8005
R3436 VGND.n405 VGND.t653 34.8005
R3437 VGND.n2093 VGND.t396 34.8005
R3438 VGND.n2093 VGND.t638 34.8005
R3439 VGND.n2332 VGND.t112 34.8005
R3440 VGND.n2332 VGND.t491 34.8005
R3441 VGND.n319 VGND.t2110 34.8005
R3442 VGND.n319 VGND.t634 34.8005
R3443 VGND.n662 VGND.t952 34.8005
R3444 VGND.n662 VGND.t1272 34.8005
R3445 VGND.n959 VGND.t1934 34.8005
R3446 VGND.n959 VGND.t1962 34.8005
R3447 VGND.n954 VGND.t2167 34.8005
R3448 VGND.n954 VGND.t819 34.8005
R3449 VGND.n949 VGND.t150 34.8005
R3450 VGND.n949 VGND.t817 34.8005
R3451 VGND.n944 VGND.t69 34.8005
R3452 VGND.n944 VGND.t2140 34.8005
R3453 VGND.n939 VGND.t1604 34.8005
R3454 VGND.n939 VGND.t1041 34.8005
R3455 VGND.n934 VGND.t139 34.8005
R3456 VGND.n934 VGND.t1039 34.8005
R3457 VGND.n929 VGND.t2402 34.8005
R3458 VGND.n929 VGND.t2138 34.8005
R3459 VGND.n924 VGND.t1071 34.8005
R3460 VGND.n924 VGND.t2136 34.8005
R3461 VGND.n919 VGND.t1160 34.8005
R3462 VGND.n919 VGND.t1960 34.8005
R3463 VGND.n914 VGND.t566 34.8005
R3464 VGND.n914 VGND.t1276 34.8005
R3465 VGND.n909 VGND.t1448 34.8005
R3466 VGND.n909 VGND.t1274 34.8005
R3467 VGND.n904 VGND.t1105 34.8005
R3468 VGND.n904 VGND.t1037 34.8005
R3469 VGND.n451 VGND.t1796 34.8005
R3470 VGND.n451 VGND.t823 34.8005
R3471 VGND.n1961 VGND.t1032 34.8005
R3472 VGND.n1961 VGND.t821 34.8005
R3473 VGND.n454 VGND.t1502 34.8005
R3474 VGND.n454 VGND.t2134 34.8005
R3475 VGND.n671 VGND.t964 34.8005
R3476 VGND.n671 VGND.t2162 34.8005
R3477 VGND.n1395 VGND.t1927 34.8005
R3478 VGND.n1395 VGND.t2038 34.8005
R3479 VGND.n1400 VGND.t1295 34.8005
R3480 VGND.n1400 VGND.t2397 34.8005
R3481 VGND.n668 VGND.t156 34.8005
R3482 VGND.n668 VGND.t2395 34.8005
R3483 VGND.n1823 VGND.t63 34.8005
R3484 VGND.n1823 VGND.t2160 34.8005
R3485 VGND.n489 VGND.t2078 34.8005
R3486 VGND.n489 VGND.t2034 34.8005
R3487 VGND.n1849 VGND.t135 34.8005
R3488 VGND.n1849 VGND.t2032 34.8005
R3489 VGND.n481 VGND.t2667 34.8005
R3490 VGND.n481 VGND.t2158 34.8005
R3491 VGND.n1875 VGND.t386 34.8005
R3492 VGND.n1875 VGND.t2156 34.8005
R3493 VGND.n473 VGND.t1464 34.8005
R3494 VGND.n473 VGND.t2036 34.8005
R3495 VGND.n1901 VGND.t562 34.8005
R3496 VGND.n1901 VGND.t2393 34.8005
R3497 VGND.n465 VGND.t1444 34.8005
R3498 VGND.n465 VGND.t2391 34.8005
R3499 VGND.n1932 VGND.t171 34.8005
R3500 VGND.n1932 VGND.t2030 34.8005
R3501 VGND.n1937 VGND.t590 34.8005
R3502 VGND.n1937 VGND.t1577 34.8005
R3503 VGND.n1942 VGND.t1812 34.8005
R3504 VGND.n1942 VGND.t1575 34.8005
R3505 VGND.n457 VGND.t2130 34.8005
R3506 VGND.n457 VGND.t868 34.8005
R3507 VGND.n1374 VGND.t892 34.8005
R3508 VGND.n1374 VGND.t1786 34.8005
R3509 VGND.n1380 VGND.t465 34.8005
R3510 VGND.n1380 VGND.t1776 34.8005
R3511 VGND.n1377 VGND.t836 34.8005
R3512 VGND.n1377 VGND.t1873 34.8005
R3513 VGND.n1810 VGND.t815 34.8005
R3514 VGND.n1810 VGND.t1871 34.8005
R3515 VGND.n493 VGND.t2513 34.8005
R3516 VGND.n493 VGND.t1784 34.8005
R3517 VGND.n1836 VGND.t283 34.8005
R3518 VGND.n1836 VGND.t1475 34.8005
R3519 VGND.n485 VGND.t1904 34.8005
R3520 VGND.n485 VGND.t1473 34.8005
R3521 VGND.n1862 VGND.t1317 34.8005
R3522 VGND.n1862 VGND.t1782 34.8005
R3523 VGND.n477 VGND.t367 34.8005
R3524 VGND.n477 VGND.t1780 34.8005
R3525 VGND.n1888 VGND.t840 34.8005
R3526 VGND.n1888 VGND.t1774 34.8005
R3527 VGND.n469 VGND.t514 34.8005
R3528 VGND.n469 VGND.t1869 34.8005
R3529 VGND.n1914 VGND.t2531 34.8005
R3530 VGND.n1914 VGND.t1867 34.8005
R3531 VGND.n461 VGND.t2596 34.8005
R3532 VGND.n461 VGND.t1471 34.8005
R3533 VGND.n1919 VGND.t399 34.8005
R3534 VGND.n1919 VGND.t1469 34.8005
R3535 VGND.n2357 VGND.t1110 34.8005
R3536 VGND.n2357 VGND.t1467 34.8005
R3537 VGND.n307 VGND.t2114 34.8005
R3538 VGND.n307 VGND.t1778 34.8005
R3539 VGND.n1306 VGND.t988 34.8005
R3540 VGND.n1306 VGND.t512 34.8005
R3541 VGND.n1312 VGND.t1124 34.8005
R3542 VGND.n1312 VGND.t575 34.8005
R3543 VGND.n1309 VGND.t1972 34.8005
R3544 VGND.n1309 VGND.t2575 34.8005
R3545 VGND.n1362 VGND.t143 34.8005
R3546 VGND.n1362 VGND.t2573 34.8005
R3547 VGND.n1357 VGND.t1195 34.8005
R3548 VGND.n1357 VGND.t510 34.8005
R3549 VGND.n1352 VGND.t2248 34.8005
R3550 VGND.n1352 VGND.t571 34.8005
R3551 VGND.n1347 VGND.t2542 34.8005
R3552 VGND.n1347 VGND.t2583 34.8005
R3553 VGND.n1342 VGND.t2660 34.8005
R3554 VGND.n1342 VGND.t581 34.8005
R3555 VGND.n1337 VGND.t392 34.8005
R3556 VGND.n1337 VGND.t579 34.8005
R3557 VGND.n1332 VGND.t1459 34.8005
R3558 VGND.n1332 VGND.t573 34.8005
R3559 VGND.n1327 VGND.t533 34.8005
R3560 VGND.n1327 VGND.t2571 34.8005
R3561 VGND.n1322 VGND.t2564 34.8005
R3562 VGND.n1322 VGND.t2569 34.8005
R3563 VGND.n1317 VGND.t2549 34.8005
R3564 VGND.n1317 VGND.t2581 34.8005
R3565 VGND.n507 VGND.t2205 34.8005
R3566 VGND.n507 VGND.t2579 34.8005
R3567 VGND.n1787 VGND.t2040 34.8005
R3568 VGND.n1787 VGND.t2577 34.8005
R3569 VGND.n510 VGND.t2122 34.8005
R3570 VGND.n510 VGND.t577 34.8005
R3571 VGND.n575 VGND.t919 34.8005
R3572 VGND.n575 VGND.t859 34.8005
R3573 VGND.n1517 VGND.t1342 34.8005
R3574 VGND.n1517 VGND.t849 34.8005
R3575 VGND.n1522 VGND.t1993 34.8005
R3576 VGND.n1522 VGND.t1498 34.8005
R3577 VGND.n579 VGND.t99 34.8005
R3578 VGND.n579 VGND.t1496 34.8005
R3579 VGND.n1649 VGND.t1163 34.8005
R3580 VGND.n1649 VGND.t857 34.8005
R3581 VGND.n545 VGND.t1709 34.8005
R3582 VGND.n545 VGND.t659 34.8005
R3583 VGND.n1675 VGND.t1561 34.8005
R3584 VGND.n1675 VGND.t657 34.8005
R3585 VGND.n537 VGND.t1310 34.8005
R3586 VGND.n537 VGND.t855 34.8005
R3587 VGND.n1701 VGND.t374 34.8005
R3588 VGND.n1701 VGND.t853 34.8005
R3589 VGND.n529 VGND.t117 34.8005
R3590 VGND.n529 VGND.t661 34.8005
R3591 VGND.n1727 VGND.t542 34.8005
R3592 VGND.n1727 VGND.t1494 34.8005
R3593 VGND.n521 VGND.t2044 34.8005
R3594 VGND.n521 VGND.t1492 34.8005
R3595 VGND.n1758 VGND.t2611 34.8005
R3596 VGND.n1758 VGND.t655 34.8005
R3597 VGND.n1763 VGND.t310 34.8005
R3598 VGND.n1763 VGND.t296 34.8005
R3599 VGND.n1768 VGND.t108 34.8005
R3600 VGND.n1768 VGND.t1500 34.8005
R3601 VGND.n513 VGND.t1513 34.8005
R3602 VGND.n513 VGND.t851 34.8005
R3603 VGND.n571 VGND.t991 34.8005
R3604 VGND.n571 VGND.t2670 34.8005
R3605 VGND.n1537 VGND.t1122 34.8005
R3606 VGND.n1537 VGND.t337 34.8005
R3607 VGND.n568 VGND.t1970 34.8005
R3608 VGND.n568 VGND.t1762 34.8005
R3609 VGND.n1636 VGND.t145 34.8005
R3610 VGND.n1636 VGND.t1760 34.8005
R3611 VGND.n549 VGND.t1193 34.8005
R3612 VGND.n549 VGND.t1553 34.8005
R3613 VGND.n1662 VGND.t2246 34.8005
R3614 VGND.n1662 VGND.t333 34.8005
R3615 VGND.n541 VGND.t2552 34.8005
R3616 VGND.n541 VGND.t331 34.8005
R3617 VGND.n1688 VGND.t2658 34.8005
R3618 VGND.n1688 VGND.t1551 34.8005
R3619 VGND.n533 VGND.t390 34.8005
R3620 VGND.n533 VGND.t341 34.8005
R3621 VGND.n1714 VGND.t1457 34.8005
R3622 VGND.n1714 VGND.t335 34.8005
R3623 VGND.n525 VGND.t531 34.8005
R3624 VGND.n525 VGND.t2674 34.8005
R3625 VGND.n1740 VGND.t2562 34.8005
R3626 VGND.n1740 VGND.t2672 34.8005
R3627 VGND.n517 VGND.t2547 34.8005
R3628 VGND.n517 VGND.t1768 34.8005
R3629 VGND.n1745 VGND.t2203 34.8005
R3630 VGND.n1745 VGND.t1766 34.8005
R3631 VGND.n2382 VGND.t1822 34.8005
R3632 VGND.n2382 VGND.t1764 34.8005
R3633 VGND.n294 VGND.t2120 34.8005
R3634 VGND.n294 VGND.t339 34.8005
R3635 VGND.n674 VGND.t1021 34.8005
R3636 VGND.n674 VGND.t1946 34.8005
R3637 VGND.n676 VGND.t827 34.8005
R3638 VGND.n676 VGND.t2307 34.8005
R3639 VGND.n1550 VGND.t2679 34.8005
R3640 VGND.n1550 VGND.t298 34.8005
R3641 VGND.n1555 VGND.t774 34.8005
R3642 VGND.n1555 VGND.t1383 34.8005
R3643 VGND.n1560 VGND.t2519 34.8005
R3644 VGND.n1560 VGND.t1944 34.8005
R3645 VGND.n1565 VGND.t2152 34.8005
R3646 VGND.n1565 VGND.t2303 34.8005
R3647 VGND.n1570 VGND.t1908 34.8005
R3648 VGND.n1570 VGND.t2301 34.8005
R3649 VGND.n1575 VGND.t664 34.8005
R3650 VGND.n1575 VGND.t1942 34.8005
R3651 VGND.n1580 VGND.t2686 34.8005
R3652 VGND.n1580 VGND.t1940 34.8005
R3653 VGND.n1585 VGND.t1133 34.8005
R3654 VGND.n1585 VGND.t2305 34.8005
R3655 VGND.n1590 VGND.t518 34.8005
R3656 VGND.n1590 VGND.t1950 34.8005
R3657 VGND.n1595 VGND.t1917 34.8005
R3658 VGND.n1595 VGND.t1948 34.8005
R3659 VGND.n1600 VGND.t2592 34.8005
R3660 VGND.n1600 VGND.t2299 34.8005
R3661 VGND.n563 VGND.t405 34.8005
R3662 VGND.n563 VGND.t2297 34.8005
R3663 VGND.n1613 VGND.t1824 34.8005
R3664 VGND.n1613 VGND.t300 34.8005
R3665 VGND.n1605 VGND.t89 34.8005
R3666 VGND.n1605 VGND.t2309 34.8005
R3667 VGND.n828 VGND.t961 34.8005
R3668 VGND.n828 VGND.t195 34.8005
R3669 VGND.n835 VGND.t1929 34.8005
R3670 VGND.n835 VGND.t2178 34.8005
R3671 VGND.n840 VGND.t1297 34.8005
R3672 VGND.n840 VGND.t2190 34.8005
R3673 VGND.n832 VGND.t154 34.8005
R3674 VGND.n832 VGND.t201 34.8005
R3675 VGND.n890 VGND.t65 34.8005
R3676 VGND.n890 VGND.t2184 34.8005
R3677 VGND.n885 VGND.t2080 34.8005
R3678 VGND.n885 VGND.t2174 34.8005
R3679 VGND.n880 VGND.t133 34.8005
R3680 VGND.n880 VGND.t2172 34.8005
R3681 VGND.n875 VGND.t2665 34.8005
R3682 VGND.n875 VGND.t2182 34.8005
R3683 VGND.n870 VGND.t384 34.8005
R3684 VGND.n870 VGND.t2180 34.8005
R3685 VGND.n865 VGND.t1462 34.8005
R3686 VGND.n865 VGND.t2176 34.8005
R3687 VGND.n860 VGND.t560 34.8005
R3688 VGND.n860 VGND.t199 34.8005
R3689 VGND.n855 VGND.t1442 34.8005
R3690 VGND.n855 VGND.t197 34.8005
R3691 VGND.n850 VGND.t169 34.8005
R3692 VGND.n850 VGND.t2170 34.8005
R3693 VGND.n845 VGND.t588 34.8005
R3694 VGND.n845 VGND.t2194 34.8005
R3695 VGND.n2402 VGND.t1814 34.8005
R3696 VGND.n2402 VGND.t2192 34.8005
R3697 VGND.n282 VGND.t2128 34.8005
R3698 VGND.n282 VGND.t810 34.8005
R3699 VGND.n818 VGND.t2471 34.8005
R3700 VGND.n818 VGND.t756 34.8005
R3701 VGND.n721 VGND.t1692 34.8005
R3702 VGND.n721 VGND.t2473 34.8005
R3703 VGND.n78 VGND.n76 34.6358
R3704 VGND.n1113 VGND.n1095 34.6358
R3705 VGND.n1109 VGND.n1095 34.6358
R3706 VGND.n1109 VGND.n1108 34.6358
R3707 VGND.n1108 VGND.n1107 34.6358
R3708 VGND.n1107 VGND.n1097 34.6358
R3709 VGND.n1091 VGND.n1065 34.6358
R3710 VGND.n1086 VGND.n1066 34.6358
R3711 VGND.n1082 VGND.n1066 34.6358
R3712 VGND.n1082 VGND.n1081 34.6358
R3713 VGND.n1081 VGND.n1080 34.6358
R3714 VGND.n1080 VGND.n1068 34.6358
R3715 VGND.n134 VGND.n129 34.6358
R3716 VGND.n139 VGND.n138 34.6358
R3717 VGND.n602 VGND.n597 34.6358
R3718 VGND.n607 VGND.n606 34.6358
R3719 VGND.n980 VGND.n979 34.6358
R3720 VGND.n988 VGND.n987 34.6358
R3721 VGND.n984 VGND.n983 34.6358
R3722 VGND.n1024 VGND.n1004 34.6358
R3723 VGND.n1020 VGND.n1004 34.6358
R3724 VGND.n1020 VGND.n1019 34.6358
R3725 VGND.n1019 VGND.n1018 34.6358
R3726 VGND.n1018 VGND.n1006 34.6358
R3727 VGND.n1060 VGND.n1034 34.6358
R3728 VGND.n1055 VGND.n1035 34.6358
R3729 VGND.n1051 VGND.n1035 34.6358
R3730 VGND.n1051 VGND.n1050 34.6358
R3731 VGND.n1050 VGND.n1049 34.6358
R3732 VGND.n1049 VGND.n1037 34.6358
R3733 VGND.n164 VGND.n159 34.6358
R3734 VGND.n169 VGND.n168 34.6358
R3735 VGND.n21 VGND.n20 34.6358
R3736 VGND.n23 VGND.n14 34.6358
R3737 VGND.n27 VGND.n14 34.6358
R3738 VGND.n28 VGND.n27 34.6358
R3739 VGND.n29 VGND.n28 34.6358
R3740 VGND.n29 VGND.n12 34.6358
R3741 VGND.n50 VGND.n49 34.6358
R3742 VGND.n52 VGND.n41 34.6358
R3743 VGND.n56 VGND.n41 34.6358
R3744 VGND.n57 VGND.n56 34.6358
R3745 VGND.n58 VGND.n57 34.6358
R3746 VGND.n58 VGND.n39 34.6358
R3747 VGND.n104 VGND.n103 34.6358
R3748 VGND.n108 VGND.n107 34.6358
R3749 VGND.n2859 VGND.n2858 34.6358
R3750 VGND.n2863 VGND.n2862 34.6358
R3751 VGND.n2891 VGND.n2890 34.6358
R3752 VGND.n2895 VGND.n2894 34.6358
R3753 VGND.n82 VGND.n81 34.6358
R3754 VGND.n2934 VGND.n2928 34.6358
R3755 VGND.n2937 VGND.n2936 34.6358
R3756 VGND.n2937 VGND.n2924 34.6358
R3757 VGND.n2941 VGND.n2924 34.6358
R3758 VGND.n2942 VGND.n2941 34.6358
R3759 VGND.n2943 VGND.n2942 34.6358
R3760 VGND.n2959 VGND.n62 34.6358
R3761 VGND.n2974 VGND.n2973 34.6358
R3762 VGND.n2976 VGND.n2965 34.6358
R3763 VGND.n2980 VGND.n2965 34.6358
R3764 VGND.n2981 VGND.n2980 34.6358
R3765 VGND.n2982 VGND.n2981 34.6358
R3766 VGND.n2982 VGND.n2963 34.6358
R3767 VGND.n2991 VGND.n2986 34.6358
R3768 VGND.n3021 VGND.t1198 34.1632
R3769 VGND.n2 VGND.t1199 34.1153
R3770 VGND.n999 VGND.n902 33.1299
R3771 VGND.n2916 VGND.n2915 33.1299
R3772 VGND.n84 VGND.n66 32.377
R3773 VGND.n990 VGND.n989 32.377
R3774 VGND.n110 VGND.n109 32.377
R3775 VGND.n2865 VGND.n2864 32.377
R3776 VGND.n2897 VGND.n2896 32.377
R3777 VGND.n84 VGND.n83 32.377
R3778 VGND.n3027 VGND.n3022 32.0005
R3779 VGND.n3031 VGND.n3030 32.0005
R3780 VGND.n990 VGND.n968 32.0005
R3781 VGND.n145 VGND.n142 30.4946
R3782 VGND.n613 VGND.n610 30.4946
R3783 VGND.n175 VGND.n172 30.4946
R3784 VGND.n113 VGND.n90 29.8709
R3785 VGND.n1103 VGND.n1102 28.9887
R3786 VGND.n1076 VGND.n1075 28.9887
R3787 VGND.n1014 VGND.n1013 28.9887
R3788 VGND.n1045 VGND.n1044 28.9887
R3789 VGND.n22 VGND.n21 27.8593
R3790 VGND.n51 VGND.n50 27.8593
R3791 VGND.n2935 VGND.n2934 27.8593
R3792 VGND.n2975 VGND.n2974 27.8593
R3793 VGND.n123 VGND.n122 27.0003
R3794 VGND.n2870 VGND.n2869 26.8591
R3795 VGND.n987 VGND.n972 26.3534
R3796 VGND.n107 VGND.n96 26.3534
R3797 VGND.n2862 VGND.n2851 26.3534
R3798 VGND.n2894 VGND.n2883 26.3534
R3799 VGND.n81 VGND.n71 26.3534
R3800 VGND.n146 VGND.n145 25.977
R3801 VGND.n614 VGND.n613 25.977
R3802 VGND.n589 VGND.n586 25.977
R3803 VGND.n176 VGND.n175 25.977
R3804 VGND.n2902 VGND.n2877 25.977
R3805 VGND.n1099 VGND.t441 24.9236
R3806 VGND.n1099 VGND.t450 24.9236
R3807 VGND.n1101 VGND.t503 24.9236
R3808 VGND.n1101 VGND.t409 24.9236
R3809 VGND.n1071 VGND.t416 24.9236
R3810 VGND.n1071 VGND.t417 24.9236
R3811 VGND.n1070 VGND.t442 24.9236
R3812 VGND.n1070 VGND.t616 24.9236
R3813 VGND.n1074 VGND.t418 24.9236
R3814 VGND.n1074 VGND.t507 24.9236
R3815 VGND.n1073 VGND.t504 24.9236
R3816 VGND.n1073 VGND.t411 24.9236
R3817 VGND.n136 VGND.t506 24.9236
R3818 VGND.n136 VGND.t2277 24.9236
R3819 VGND.n135 VGND.t619 24.9236
R3820 VGND.n135 VGND.t596 24.9236
R3821 VGND.n126 VGND.t104 24.9236
R3822 VGND.n126 VGND.t624 24.9236
R3823 VGND.n125 VGND.t1911 24.9236
R3824 VGND.n125 VGND.t446 24.9236
R3825 VGND.n144 VGND.t101 24.9236
R3826 VGND.n144 VGND.t102 24.9236
R3827 VGND.n143 VGND.t1909 24.9236
R3828 VGND.n143 VGND.t1910 24.9236
R3829 VGND.n604 VGND.t2364 24.9236
R3830 VGND.n604 VGND.t437 24.9236
R3831 VGND.n603 VGND.t2279 24.9236
R3832 VGND.n603 VGND.t1599 24.9236
R3833 VGND.n594 VGND.t289 24.9236
R3834 VGND.n594 VGND.t2363 24.9236
R3835 VGND.n593 VGND.t1396 24.9236
R3836 VGND.n593 VGND.t2276 24.9236
R3837 VGND.n612 VGND.t291 24.9236
R3838 VGND.n612 VGND.t290 24.9236
R3839 VGND.n611 VGND.t1398 24.9236
R3840 VGND.n611 VGND.t1397 24.9236
R3841 VGND.n970 VGND.t448 24.9236
R3842 VGND.n970 VGND.t593 24.9236
R3843 VGND.n971 VGND.t214 24.9236
R3844 VGND.n971 VGND.t621 24.9236
R3845 VGND.n969 VGND.t218 24.9236
R3846 VGND.n969 VGND.t216 24.9236
R3847 VGND.n974 VGND.t623 24.9236
R3848 VGND.n974 VGND.t407 24.9236
R3849 VGND.n1009 VGND.t443 24.9236
R3850 VGND.n1009 VGND.t617 24.9236
R3851 VGND.n1008 VGND.t1600 24.9236
R3852 VGND.n1008 VGND.t435 24.9236
R3853 VGND.n1012 VGND.t505 24.9236
R3854 VGND.n1012 VGND.t412 24.9236
R3855 VGND.n1011 VGND.t615 24.9236
R3856 VGND.n1011 VGND.t594 24.9236
R3857 VGND.n1040 VGND.t508 24.9236
R3858 VGND.n1040 VGND.t678 24.9236
R3859 VGND.n1039 VGND.t595 24.9236
R3860 VGND.n1039 VGND.t597 24.9236
R3861 VGND.n1043 VGND.t679 24.9236
R3862 VGND.n1043 VGND.t415 24.9236
R3863 VGND.n1042 VGND.t2278 24.9236
R3864 VGND.n1042 VGND.t1598 24.9236
R3865 VGND.n166 VGND.t414 24.9236
R3866 VGND.n166 VGND.t445 24.9236
R3867 VGND.n165 VGND.t2362 24.9236
R3868 VGND.n165 VGND.t1602 24.9236
R3869 VGND.n156 VGND.t1103 24.9236
R3870 VGND.n156 VGND.t2365 24.9236
R3871 VGND.n155 VGND.t205 24.9236
R3872 VGND.n155 VGND.t2361 24.9236
R3873 VGND.n174 VGND.t1101 24.9236
R3874 VGND.n174 VGND.t1102 24.9236
R3875 VGND.n173 VGND.t208 24.9236
R3876 VGND.n173 VGND.t206 24.9236
R3877 VGND.n17 VGND.t1262 24.9236
R3878 VGND.n17 VGND.t2587 24.9236
R3879 VGND.n16 VGND.t459 24.9236
R3880 VGND.n16 VGND.t452 24.9236
R3881 VGND.n46 VGND.t607 24.9236
R3882 VGND.n46 VGND.t669 24.9236
R3883 VGND.n45 VGND.t454 24.9236
R3884 VGND.n45 VGND.t612 24.9236
R3885 VGND.n44 VGND.t555 24.9236
R3886 VGND.n44 VGND.t500 24.9236
R3887 VGND.n43 VGND.t429 24.9236
R3888 VGND.n43 VGND.t1258 24.9236
R3889 VGND.n99 VGND.t463 24.9236
R3890 VGND.n99 VGND.t316 24.9236
R3891 VGND.n98 VGND.t604 24.9236
R3892 VGND.n98 VGND.t2584 24.9236
R3893 VGND.n95 VGND.t456 24.9236
R3894 VGND.n95 VGND.t1979 24.9236
R3895 VGND.n94 VGND.t550 24.9236
R3896 VGND.n94 VGND.t1937 24.9236
R3897 VGND.n93 VGND.t1978 24.9236
R3898 VGND.n93 VGND.t1980 24.9236
R3899 VGND.n92 VGND.t1556 24.9236
R3900 VGND.n92 VGND.t1097 24.9236
R3901 VGND.n2854 VGND.t496 24.9236
R3902 VGND.n2854 VGND.t549 24.9236
R3903 VGND.n2853 VGND.t1255 24.9236
R3904 VGND.n2853 VGND.t498 24.9236
R3905 VGND.n2850 VGND.t322 24.9236
R3906 VGND.n2850 VGND.t192 24.9236
R3907 VGND.n2849 VGND.t2588 24.9236
R3908 VGND.n2849 VGND.t294 24.9236
R3909 VGND.n2848 VGND.t189 24.9236
R3910 VGND.n2848 VGND.t183 24.9236
R3911 VGND.n2847 VGND.t2683 24.9236
R3912 VGND.n2847 VGND.t1250 24.9236
R3913 VGND.n2886 VGND.t324 24.9236
R3914 VGND.n2886 VGND.t544 24.9236
R3915 VGND.n2885 VGND.t432 24.9236
R3916 VGND.n2885 VGND.t605 24.9236
R3917 VGND.n2882 VGND.t318 24.9236
R3918 VGND.n2882 VGND.t265 24.9236
R3919 VGND.n2881 VGND.t423 24.9236
R3920 VGND.n2881 VGND.t2653 24.9236
R3921 VGND.n2880 VGND.t261 24.9236
R3922 VGND.n2880 VGND.t255 24.9236
R3923 VGND.n2879 VGND.t2652 24.9236
R3924 VGND.n2879 VGND.t2650 24.9236
R3925 VGND.n69 VGND.t614 24.9236
R3926 VGND.n69 VGND.t672 24.9236
R3927 VGND.n70 VGND.t610 24.9236
R3928 VGND.n70 VGND.t1752 24.9236
R3929 VGND.n68 VGND.t1748 24.9236
R3930 VGND.n68 VGND.t1742 24.9236
R3931 VGND.n73 VGND.t314 24.9236
R3932 VGND.n73 VGND.t1260 24.9236
R3933 VGND.n2930 VGND.t501 24.9236
R3934 VGND.n2930 VGND.t552 24.9236
R3935 VGND.n2929 VGND.t434 24.9236
R3936 VGND.n2929 VGND.t608 24.9236
R3937 VGND.n2927 VGND.t492 24.9236
R3938 VGND.n2927 VGND.t2585 24.9236
R3939 VGND.n2926 VGND.t427 24.9236
R3940 VGND.n2926 VGND.t1257 24.9236
R3941 VGND.n2970 VGND.t1265 24.9236
R3942 VGND.n2970 VGND.t425 24.9236
R3943 VGND.n2969 VGND.t554 24.9236
R3944 VGND.n2969 VGND.t457 24.9236
R3945 VGND.n2968 VGND.t1253 24.9236
R3946 VGND.n2968 VGND.t606 24.9236
R3947 VGND.n2967 VGND.t548 24.9236
R3948 VGND.n2967 VGND.t320 24.9236
R3949 VGND.n146 VGND.n120 24.4711
R3950 VGND.n614 VGND.n585 24.4711
R3951 VGND.n589 VGND.n588 24.4711
R3952 VGND.n1000 VGND.n999 24.4711
R3953 VGND.n1029 VGND.n1003 24.4711
R3954 VGND.n176 VGND.n152 24.4711
R3955 VGND.n110 VGND.n89 24.4711
R3956 VGND.n2865 VGND.n2844 24.4711
R3957 VGND.n2897 VGND.n2876 24.4711
R3958 VGND.n2902 VGND.n2901 24.4711
R3959 VGND.n2917 VGND.n2916 24.4711
R3960 VGND.n2948 VGND.n2947 24.4711
R3961 VGND.n2873 VGND.n2845 23.7181
R3962 VGND.n1115 VGND.n1113 23.7181
R3963 VGND.n1087 VGND.n1065 23.7181
R3964 VGND.n1087 VGND.n1086 23.7181
R3965 VGND.n150 VGND.n119 23.7181
R3966 VGND.n994 VGND.n903 23.7181
R3967 VGND.n1025 VGND.n1024 23.7181
R3968 VGND.n1056 VGND.n1034 23.7181
R3969 VGND.n1056 VGND.n1055 23.7181
R3970 VGND.n3007 VGND.n12 23.7181
R3971 VGND.n2960 VGND.n39 23.7181
R3972 VGND.n2943 VGND.n2922 23.7181
R3973 VGND.n2960 VGND.n2959 23.7181
R3974 VGND.n2992 VGND.n2963 23.7181
R3975 VGND.n2992 VGND.n2991 23.7181
R3976 VGND.n995 VGND.n994 23.3417
R3977 VGND.n2911 VGND.n88 23.3417
R3978 VGND.n2911 VGND.n65 23.3417
R3979 VGND.n1103 VGND.n1100 21.4593
R3980 VGND.n1076 VGND.n1072 21.4593
R3981 VGND.n1014 VGND.n1010 21.4593
R3982 VGND.n1045 VGND.n1041 21.4593
R3983 VGND.n102 VGND.n101 21.0905
R3984 VGND.n2857 VGND.n2856 21.0905
R3985 VGND.n2889 VGND.n2888 21.0905
R3986 VGND.n75 VGND.n74 21.0905
R3987 VGND.n103 VGND.n102 20.3299
R3988 VGND.n2858 VGND.n2857 20.3299
R3989 VGND.n2890 VGND.n2889 20.3299
R3990 VGND.n76 VGND.n75 20.3299
R3991 VGND.n142 VGND.n127 19.9534
R3992 VGND.n610 VGND.n595 19.9534
R3993 VGND.n172 VGND.n157 19.9534
R3994 VGND.n1030 VGND.n1029 19.2005
R3995 VGND.n1061 VGND.n1060 19.2005
R3996 VGND.n2949 VGND.n2948 19.2005
R3997 VGND.n2954 VGND.n62 19.2005
R3998 VGND.t2524 VGND.t675 16.8587
R3999 VGND.t1329 VGND.t673 16.8587
R4000 VGND.t1585 VGND.t1372 16.8587
R4001 VGND.t2646 VGND.t1374 16.8587
R4002 VGND.n1093 VGND.n1092 16.077
R4003 VGND.n2988 VGND.n2987 16.077
R4004 VGND.n1031 VGND.n1030 15.4358
R4005 VGND.n2950 VGND.n2949 15.4358
R4006 VGND.n122 VGND.n121 14.6829
R4007 VGND.n1062 VGND.n1061 14.6829
R4008 VGND.n2869 VGND.n2868 14.6829
R4009 VGND.n2955 VGND.n2954 14.6829
R4010 VGND.n131 VGND.n130 14.5711
R4011 VGND.n599 VGND.n598 14.5711
R4012 VGND.n978 VGND.n977 14.5711
R4013 VGND.n161 VGND.n160 14.5711
R4014 VGND.n618 VGND.n586 14.3064
R4015 VGND.n2906 VGND.n2877 14.3064
R4016 VGND.n138 VGND.n137 13.9299
R4017 VGND.n606 VGND.n605 13.9299
R4018 VGND.n983 VGND.n975 13.9299
R4019 VGND.n168 VGND.n167 13.9299
R4020 VGND.n1025 VGND.n1003 13.5534
R4021 VGND.n2947 VGND.n2922 13.5534
R4022 VGND.n150 VGND.n120 13.177
R4023 VGND.n618 VGND.n585 13.177
R4024 VGND.n180 VGND.n152 13.177
R4025 VGND.n116 VGND.n89 13.177
R4026 VGND.n2873 VGND.n2844 13.177
R4027 VGND.n2906 VGND.n2876 13.177
R4028 VGND.n180 VGND.n153 12.8005
R4029 VGND.n116 VGND.n90 12.8005
R4030 VGND.n1092 VGND.n1091 10.5417
R4031 VGND.n2987 VGND.n2986 10.5417
R4032 VGND.n1063 VGND.n1062 10.0534
R4033 VGND.n2956 VGND.n2955 10.0534
R4034 VGND.n1104 VGND.n1103 9.3005
R4035 VGND.n1105 VGND.n1097 9.3005
R4036 VGND.n1107 VGND.n1106 9.3005
R4037 VGND.n1108 VGND.n1096 9.3005
R4038 VGND.n1110 VGND.n1109 9.3005
R4039 VGND.n1111 VGND.n1095 9.3005
R4040 VGND.n1113 VGND.n1112 9.3005
R4041 VGND.n1116 VGND.n1115 9.3005
R4042 VGND.n1077 VGND.n1076 9.3005
R4043 VGND.n1078 VGND.n1068 9.3005
R4044 VGND.n1080 VGND.n1079 9.3005
R4045 VGND.n1081 VGND.n1067 9.3005
R4046 VGND.n1083 VGND.n1082 9.3005
R4047 VGND.n1084 VGND.n1066 9.3005
R4048 VGND.n1086 VGND.n1085 9.3005
R4049 VGND.n1089 VGND.n1065 9.3005
R4050 VGND.n1091 VGND.n1090 9.3005
R4051 VGND.n1088 VGND.n1087 9.3005
R4052 VGND.n148 VGND.n120 9.3005
R4053 VGND.n132 VGND.n129 9.3005
R4054 VGND.n134 VGND.n133 9.3005
R4055 VGND.n138 VGND.n128 9.3005
R4056 VGND.n140 VGND.n139 9.3005
R4057 VGND.n142 VGND.n141 9.3005
R4058 VGND.n145 VGND.n124 9.3005
R4059 VGND.n147 VGND.n146 9.3005
R4060 VGND.n123 VGND.n119 9.3005
R4061 VGND.n150 VGND.n149 9.3005
R4062 VGND.n588 VGND.n587 9.3005
R4063 VGND.n591 VGND.n586 9.3005
R4064 VGND.n616 VGND.n585 9.3005
R4065 VGND.n600 VGND.n597 9.3005
R4066 VGND.n602 VGND.n601 9.3005
R4067 VGND.n606 VGND.n596 9.3005
R4068 VGND.n608 VGND.n607 9.3005
R4069 VGND.n610 VGND.n609 9.3005
R4070 VGND.n613 VGND.n592 9.3005
R4071 VGND.n615 VGND.n614 9.3005
R4072 VGND.n590 VGND.n589 9.3005
R4073 VGND.n618 VGND.n617 9.3005
R4074 VGND.n1001 VGND.n1000 9.3005
R4075 VGND.n992 VGND.n903 9.3005
R4076 VGND.n979 VGND.n976 9.3005
R4077 VGND.n981 VGND.n980 9.3005
R4078 VGND.n983 VGND.n982 9.3005
R4079 VGND.n985 VGND.n984 9.3005
R4080 VGND.n987 VGND.n986 9.3005
R4081 VGND.n988 VGND.n967 9.3005
R4082 VGND.n991 VGND.n990 9.3005
R4083 VGND.n997 VGND.n996 9.3005
R4084 VGND.n999 VGND.n998 9.3005
R4085 VGND.n994 VGND.n993 9.3005
R4086 VGND.n1015 VGND.n1014 9.3005
R4087 VGND.n1016 VGND.n1006 9.3005
R4088 VGND.n1018 VGND.n1017 9.3005
R4089 VGND.n1019 VGND.n1005 9.3005
R4090 VGND.n1021 VGND.n1020 9.3005
R4091 VGND.n1022 VGND.n1004 9.3005
R4092 VGND.n1024 VGND.n1023 9.3005
R4093 VGND.n1027 VGND.n1003 9.3005
R4094 VGND.n1029 VGND.n1028 9.3005
R4095 VGND.n1032 VGND.n1031 9.3005
R4096 VGND.n1026 VGND.n1025 9.3005
R4097 VGND.n1046 VGND.n1045 9.3005
R4098 VGND.n1047 VGND.n1037 9.3005
R4099 VGND.n1049 VGND.n1048 9.3005
R4100 VGND.n1050 VGND.n1036 9.3005
R4101 VGND.n1052 VGND.n1051 9.3005
R4102 VGND.n1053 VGND.n1035 9.3005
R4103 VGND.n1055 VGND.n1054 9.3005
R4104 VGND.n1058 VGND.n1034 9.3005
R4105 VGND.n1060 VGND.n1059 9.3005
R4106 VGND.n1057 VGND.n1056 9.3005
R4107 VGND.n178 VGND.n152 9.3005
R4108 VGND.n162 VGND.n159 9.3005
R4109 VGND.n164 VGND.n163 9.3005
R4110 VGND.n168 VGND.n158 9.3005
R4111 VGND.n170 VGND.n169 9.3005
R4112 VGND.n172 VGND.n171 9.3005
R4113 VGND.n175 VGND.n154 9.3005
R4114 VGND.n177 VGND.n176 9.3005
R4115 VGND.n180 VGND.n179 9.3005
R4116 VGND.n3007 VGND.n3006 9.3005
R4117 VGND.n20 VGND.n19 9.3005
R4118 VGND.n21 VGND.n15 9.3005
R4119 VGND.n24 VGND.n23 9.3005
R4120 VGND.n25 VGND.n14 9.3005
R4121 VGND.n27 VGND.n26 9.3005
R4122 VGND.n28 VGND.n13 9.3005
R4123 VGND.n30 VGND.n29 9.3005
R4124 VGND.n31 VGND.n12 9.3005
R4125 VGND.n114 VGND.n90 9.3005
R4126 VGND.n103 VGND.n97 9.3005
R4127 VGND.n105 VGND.n104 9.3005
R4128 VGND.n107 VGND.n106 9.3005
R4129 VGND.n108 VGND.n91 9.3005
R4130 VGND.n111 VGND.n110 9.3005
R4131 VGND.n112 VGND.n89 9.3005
R4132 VGND.n116 VGND.n115 9.3005
R4133 VGND.n2871 VGND.n2845 9.3005
R4134 VGND.n2858 VGND.n2852 9.3005
R4135 VGND.n2860 VGND.n2859 9.3005
R4136 VGND.n2862 VGND.n2861 9.3005
R4137 VGND.n2863 VGND.n2846 9.3005
R4138 VGND.n2866 VGND.n2865 9.3005
R4139 VGND.n2867 VGND.n2844 9.3005
R4140 VGND.n2873 VGND.n2872 9.3005
R4141 VGND.n2901 VGND.n2900 9.3005
R4142 VGND.n2890 VGND.n2884 9.3005
R4143 VGND.n2892 VGND.n2891 9.3005
R4144 VGND.n2894 VGND.n2893 9.3005
R4145 VGND.n2895 VGND.n2878 9.3005
R4146 VGND.n2898 VGND.n2897 9.3005
R4147 VGND.n2899 VGND.n2876 9.3005
R4148 VGND.n2904 VGND.n2877 9.3005
R4149 VGND.n2903 VGND.n2902 9.3005
R4150 VGND.n2906 VGND.n2905 9.3005
R4151 VGND.n2918 VGND.n2917 9.3005
R4152 VGND.n76 VGND.n72 9.3005
R4153 VGND.n79 VGND.n78 9.3005
R4154 VGND.n81 VGND.n80 9.3005
R4155 VGND.n82 VGND.n67 9.3005
R4156 VGND.n85 VGND.n84 9.3005
R4157 VGND.n87 VGND.n86 9.3005
R4158 VGND.n2914 VGND.n2913 9.3005
R4159 VGND.n2916 VGND.n64 9.3005
R4160 VGND.n2912 VGND.n2911 9.3005
R4161 VGND.n2951 VGND.n2950 9.3005
R4162 VGND.n2932 VGND.n2928 9.3005
R4163 VGND.n2934 VGND.n2933 9.3005
R4164 VGND.n2936 VGND.n2925 9.3005
R4165 VGND.n2938 VGND.n2937 9.3005
R4166 VGND.n2939 VGND.n2924 9.3005
R4167 VGND.n2941 VGND.n2940 9.3005
R4168 VGND.n2942 VGND.n2923 9.3005
R4169 VGND.n2944 VGND.n2943 9.3005
R4170 VGND.n2947 VGND.n2946 9.3005
R4171 VGND.n2948 VGND.n2920 9.3005
R4172 VGND.n2945 VGND.n2922 9.3005
R4173 VGND.n49 VGND.n48 9.3005
R4174 VGND.n50 VGND.n42 9.3005
R4175 VGND.n53 VGND.n52 9.3005
R4176 VGND.n54 VGND.n41 9.3005
R4177 VGND.n56 VGND.n55 9.3005
R4178 VGND.n57 VGND.n40 9.3005
R4179 VGND.n59 VGND.n58 9.3005
R4180 VGND.n60 VGND.n39 9.3005
R4181 VGND.n2960 VGND.n61 9.3005
R4182 VGND.n2959 VGND.n2958 9.3005
R4183 VGND.n2957 VGND.n62 9.3005
R4184 VGND.n2973 VGND.n2972 9.3005
R4185 VGND.n2974 VGND.n2966 9.3005
R4186 VGND.n2977 VGND.n2976 9.3005
R4187 VGND.n2978 VGND.n2965 9.3005
R4188 VGND.n2980 VGND.n2979 9.3005
R4189 VGND.n2981 VGND.n2964 9.3005
R4190 VGND.n2983 VGND.n2982 9.3005
R4191 VGND.n2984 VGND.n2963 9.3005
R4192 VGND.n2992 VGND.n2985 9.3005
R4193 VGND.n2991 VGND.n2990 9.3005
R4194 VGND.n2989 VGND.n2986 9.3005
R4195 VGND.n104 VGND.n96 8.28285
R4196 VGND.n2859 VGND.n2851 8.28285
R4197 VGND.n2891 VGND.n2883 8.28285
R4198 VGND.n2716 VGND.n239 7.9105
R4199 VGND.n2718 VGND.n2717 7.9105
R4200 VGND.n2823 VGND.n193 7.9105
R4201 VGND.n2822 VGND.n194 7.9105
R4202 VGND.n2817 VGND.n199 7.9105
R4203 VGND.n2816 VGND.n200 7.9105
R4204 VGND.n2811 VGND.n205 7.9105
R4205 VGND.n2810 VGND.n206 7.9105
R4206 VGND.n2805 VGND.n211 7.9105
R4207 VGND.n2804 VGND.n212 7.9105
R4208 VGND.n2799 VGND.n217 7.9105
R4209 VGND.n2798 VGND.n218 7.9105
R4210 VGND.n2793 VGND.n223 7.9105
R4211 VGND.n2792 VGND.n224 7.9105
R4212 VGND.n2787 VGND.n2786 7.9105
R4213 VGND.n3001 VGND.n3000 7.9105
R4214 VGND.n2521 VGND.n2520 7.9105
R4215 VGND.n2827 VGND.n189 7.9105
R4216 VGND.n2826 VGND.n190 7.9105
R4217 VGND.n2508 VGND.n2507 7.9105
R4218 VGND.n2506 VGND.n252 7.9105
R4219 VGND.n2505 VGND.n253 7.9105
R4220 VGND.n2504 VGND.n254 7.9105
R4221 VGND.n2503 VGND.n255 7.9105
R4222 VGND.n2502 VGND.n256 7.9105
R4223 VGND.n2501 VGND.n257 7.9105
R4224 VGND.n2500 VGND.n258 7.9105
R4225 VGND.n2499 VGND.n259 7.9105
R4226 VGND.n2498 VGND.n260 7.9105
R4227 VGND.n2497 VGND.n261 7.9105
R4228 VGND.n2496 VGND.n262 7.9105
R4229 VGND.n2495 VGND.n2494 7.9105
R4230 VGND.n643 VGND.n184 7.9105
R4231 VGND.n2831 VGND.n2830 7.9105
R4232 VGND.n379 VGND.n378 7.9105
R4233 VGND.n2170 VGND.n2169 7.9105
R4234 VGND.n2179 VGND.n2178 7.9105
R4235 VGND.n2196 VGND.n2195 7.9105
R4236 VGND.n2205 VGND.n2204 7.9105
R4237 VGND.n2222 VGND.n2221 7.9105
R4238 VGND.n2231 VGND.n2230 7.9105
R4239 VGND.n2248 VGND.n2247 7.9105
R4240 VGND.n2257 VGND.n2256 7.9105
R4241 VGND.n2279 VGND.n2278 7.9105
R4242 VGND.n2301 VGND.n332 7.9105
R4243 VGND.n2300 VGND.n333 7.9105
R4244 VGND.n2298 VGND.n2297 7.9105
R4245 VGND.n2434 VGND.n2433 7.9105
R4246 VGND.n1437 VGND.n1424 7.9105
R4247 VGND.n1436 VGND.n1435 7.9105
R4248 VGND.n2157 VGND.n2156 7.9105
R4249 VGND.n2166 VGND.n2165 7.9105
R4250 VGND.n2183 VGND.n2182 7.9105
R4251 VGND.n2192 VGND.n2191 7.9105
R4252 VGND.n2209 VGND.n2208 7.9105
R4253 VGND.n2218 VGND.n2217 7.9105
R4254 VGND.n2235 VGND.n2234 7.9105
R4255 VGND.n2244 VGND.n2243 7.9105
R4256 VGND.n2261 VGND.n2260 7.9105
R4257 VGND.n2275 VGND.n2274 7.9105
R4258 VGND.n2304 VGND.n331 7.9105
R4259 VGND.n2306 VGND.n2305 7.9105
R4260 VGND.n2318 VGND.n328 7.9105
R4261 VGND.n2317 VGND.n2316 7.9105
R4262 VGND.n1441 VGND.n1440 7.9105
R4263 VGND.n1500 VGND.n1499 7.9105
R4264 VGND.n2153 VGND.n385 7.9105
R4265 VGND.n2152 VGND.n386 7.9105
R4266 VGND.n2151 VGND.n387 7.9105
R4267 VGND.n2150 VGND.n388 7.9105
R4268 VGND.n2149 VGND.n389 7.9105
R4269 VGND.n2148 VGND.n390 7.9105
R4270 VGND.n2147 VGND.n391 7.9105
R4271 VGND.n2146 VGND.n392 7.9105
R4272 VGND.n2145 VGND.n393 7.9105
R4273 VGND.n2144 VGND.n394 7.9105
R4274 VGND.n2143 VGND.n2142 7.9105
R4275 VGND.n2322 VGND.n325 7.9105
R4276 VGND.n2321 VGND.n326 7.9105
R4277 VGND.n2130 VGND.n2129 7.9105
R4278 VGND.n1418 VGND.n621 7.9105
R4279 VGND.n1504 VGND.n1503 7.9105
R4280 VGND.n634 VGND.n633 7.9105
R4281 VGND.n1996 VGND.n1995 7.9105
R4282 VGND.n2005 VGND.n2004 7.9105
R4283 VGND.n2022 VGND.n2021 7.9105
R4284 VGND.n2031 VGND.n2030 7.9105
R4285 VGND.n2048 VGND.n2047 7.9105
R4286 VGND.n2057 VGND.n2056 7.9105
R4287 VGND.n2074 VGND.n2073 7.9105
R4288 VGND.n2083 VGND.n2082 7.9105
R4289 VGND.n2105 VGND.n2104 7.9105
R4290 VGND.n2326 VGND.n322 7.9105
R4291 VGND.n2325 VGND.n323 7.9105
R4292 VGND.n403 VGND.n402 7.9105
R4293 VGND.n2126 VGND.n2125 7.9105
R4294 VGND.n1416 VGND.n648 7.9105
R4295 VGND.n660 VGND.n659 7.9105
R4296 VGND.n1983 VGND.n1982 7.9105
R4297 VGND.n1992 VGND.n1991 7.9105
R4298 VGND.n2009 VGND.n2008 7.9105
R4299 VGND.n2018 VGND.n2017 7.9105
R4300 VGND.n2035 VGND.n2034 7.9105
R4301 VGND.n2044 VGND.n2043 7.9105
R4302 VGND.n2061 VGND.n2060 7.9105
R4303 VGND.n2070 VGND.n2069 7.9105
R4304 VGND.n2087 VGND.n2086 7.9105
R4305 VGND.n2101 VGND.n2100 7.9105
R4306 VGND.n2329 VGND.n320 7.9105
R4307 VGND.n2331 VGND.n2330 7.9105
R4308 VGND.n2343 VGND.n316 7.9105
R4309 VGND.n2342 VGND.n2341 7.9105
R4310 VGND.n1413 VGND.n664 7.9105
R4311 VGND.n1412 VGND.n665 7.9105
R4312 VGND.n1979 VGND.n441 7.9105
R4313 VGND.n1978 VGND.n442 7.9105
R4314 VGND.n1977 VGND.n443 7.9105
R4315 VGND.n1976 VGND.n444 7.9105
R4316 VGND.n1975 VGND.n445 7.9105
R4317 VGND.n1974 VGND.n446 7.9105
R4318 VGND.n1973 VGND.n447 7.9105
R4319 VGND.n1972 VGND.n448 7.9105
R4320 VGND.n1971 VGND.n449 7.9105
R4321 VGND.n1970 VGND.n450 7.9105
R4322 VGND.n1969 VGND.n1968 7.9105
R4323 VGND.n2347 VGND.n313 7.9105
R4324 VGND.n2346 VGND.n314 7.9105
R4325 VGND.n1956 VGND.n1955 7.9105
R4326 VGND.n1394 VGND.n1393 7.9105
R4327 VGND.n1409 VGND.n667 7.9105
R4328 VGND.n1408 VGND.n1407 7.9105
R4329 VGND.n1822 VGND.n1821 7.9105
R4330 VGND.n1831 VGND.n1830 7.9105
R4331 VGND.n1848 VGND.n1847 7.9105
R4332 VGND.n1857 VGND.n1856 7.9105
R4333 VGND.n1874 VGND.n1873 7.9105
R4334 VGND.n1883 VGND.n1882 7.9105
R4335 VGND.n1900 VGND.n1899 7.9105
R4336 VGND.n1909 VGND.n1908 7.9105
R4337 VGND.n1931 VGND.n1930 7.9105
R4338 VGND.n2351 VGND.n310 7.9105
R4339 VGND.n2350 VGND.n311 7.9105
R4340 VGND.n459 VGND.n458 7.9105
R4341 VGND.n1952 VGND.n1951 7.9105
R4342 VGND.n1390 VGND.n1376 7.9105
R4343 VGND.n1388 VGND.n1387 7.9105
R4344 VGND.n1809 VGND.n1808 7.9105
R4345 VGND.n1818 VGND.n1817 7.9105
R4346 VGND.n1835 VGND.n1834 7.9105
R4347 VGND.n1844 VGND.n1843 7.9105
R4348 VGND.n1861 VGND.n1860 7.9105
R4349 VGND.n1870 VGND.n1869 7.9105
R4350 VGND.n1887 VGND.n1886 7.9105
R4351 VGND.n1896 VGND.n1895 7.9105
R4352 VGND.n1913 VGND.n1912 7.9105
R4353 VGND.n1927 VGND.n1926 7.9105
R4354 VGND.n2354 VGND.n308 7.9105
R4355 VGND.n2356 VGND.n2355 7.9105
R4356 VGND.n2368 VGND.n304 7.9105
R4357 VGND.n2367 VGND.n2366 7.9105
R4358 VGND.n1372 VGND.n1308 7.9105
R4359 VGND.n1371 VGND.n1369 7.9105
R4360 VGND.n1805 VGND.n497 7.9105
R4361 VGND.n1804 VGND.n498 7.9105
R4362 VGND.n1803 VGND.n499 7.9105
R4363 VGND.n1802 VGND.n500 7.9105
R4364 VGND.n1801 VGND.n501 7.9105
R4365 VGND.n1800 VGND.n502 7.9105
R4366 VGND.n1799 VGND.n503 7.9105
R4367 VGND.n1798 VGND.n504 7.9105
R4368 VGND.n1797 VGND.n505 7.9105
R4369 VGND.n1796 VGND.n506 7.9105
R4370 VGND.n1795 VGND.n1794 7.9105
R4371 VGND.n2372 VGND.n301 7.9105
R4372 VGND.n2371 VGND.n302 7.9105
R4373 VGND.n1782 VGND.n1781 7.9105
R4374 VGND.n1532 VGND.n577 7.9105
R4375 VGND.n1531 VGND.n578 7.9105
R4376 VGND.n1530 VGND.n1529 7.9105
R4377 VGND.n1648 VGND.n1647 7.9105
R4378 VGND.n1657 VGND.n1656 7.9105
R4379 VGND.n1674 VGND.n1673 7.9105
R4380 VGND.n1683 VGND.n1682 7.9105
R4381 VGND.n1700 VGND.n1699 7.9105
R4382 VGND.n1709 VGND.n1708 7.9105
R4383 VGND.n1726 VGND.n1725 7.9105
R4384 VGND.n1735 VGND.n1734 7.9105
R4385 VGND.n1757 VGND.n1756 7.9105
R4386 VGND.n2376 VGND.n298 7.9105
R4387 VGND.n2375 VGND.n299 7.9105
R4388 VGND.n515 VGND.n514 7.9105
R4389 VGND.n1778 VGND.n1777 7.9105
R4390 VGND.n1536 VGND.n1535 7.9105
R4391 VGND.n1545 VGND.n1544 7.9105
R4392 VGND.n1635 VGND.n1634 7.9105
R4393 VGND.n1644 VGND.n1643 7.9105
R4394 VGND.n1661 VGND.n1660 7.9105
R4395 VGND.n1670 VGND.n1669 7.9105
R4396 VGND.n1687 VGND.n1686 7.9105
R4397 VGND.n1696 VGND.n1695 7.9105
R4398 VGND.n1713 VGND.n1712 7.9105
R4399 VGND.n1722 VGND.n1721 7.9105
R4400 VGND.n1739 VGND.n1738 7.9105
R4401 VGND.n1753 VGND.n1752 7.9105
R4402 VGND.n2379 VGND.n295 7.9105
R4403 VGND.n2381 VGND.n2380 7.9105
R4404 VGND.n2393 VGND.n291 7.9105
R4405 VGND.n2392 VGND.n2391 7.9105
R4406 VGND.n1302 VGND.n1301 7.9105
R4407 VGND.n1549 VGND.n1548 7.9105
R4408 VGND.n1631 VGND.n553 7.9105
R4409 VGND.n1630 VGND.n554 7.9105
R4410 VGND.n1629 VGND.n555 7.9105
R4411 VGND.n1628 VGND.n556 7.9105
R4412 VGND.n1627 VGND.n557 7.9105
R4413 VGND.n1626 VGND.n558 7.9105
R4414 VGND.n1625 VGND.n559 7.9105
R4415 VGND.n1624 VGND.n560 7.9105
R4416 VGND.n1623 VGND.n561 7.9105
R4417 VGND.n1622 VGND.n562 7.9105
R4418 VGND.n1621 VGND.n1620 7.9105
R4419 VGND.n2397 VGND.n286 7.9105
R4420 VGND.n2396 VGND.n287 7.9105
R4421 VGND.n1608 VGND.n1607 7.9105
R4422 VGND.n900 VGND.n830 7.9105
R4423 VGND.n899 VGND.n831 7.9105
R4424 VGND.n898 VGND.n897 7.9105
R4425 VGND.n1279 VGND.n692 7.9105
R4426 VGND.n1278 VGND.n693 7.9105
R4427 VGND.n1271 VGND.n698 7.9105
R4428 VGND.n1270 VGND.n699 7.9105
R4429 VGND.n1263 VGND.n704 7.9105
R4430 VGND.n1262 VGND.n705 7.9105
R4431 VGND.n1255 VGND.n710 7.9105
R4432 VGND.n1254 VGND.n711 7.9105
R4433 VGND.n1247 VGND.n716 7.9105
R4434 VGND.n1246 VGND.n717 7.9105
R4435 VGND.n2401 VGND.n2400 7.9105
R4436 VGND.n288 VGND.n283 7.9105
R4437 VGND.n2412 VGND.n2411 7.9105
R4438 VGND.n1121 VGND.n681 7.9105
R4439 VGND.n1289 VGND.n1288 7.9105
R4440 VGND.n1283 VGND.n689 7.9105
R4441 VGND.n1282 VGND.n690 7.9105
R4442 VGND.n1275 VGND.n695 7.9105
R4443 VGND.n1274 VGND.n696 7.9105
R4444 VGND.n1267 VGND.n701 7.9105
R4445 VGND.n1266 VGND.n702 7.9105
R4446 VGND.n1259 VGND.n707 7.9105
R4447 VGND.n1258 VGND.n708 7.9105
R4448 VGND.n1251 VGND.n713 7.9105
R4449 VGND.n1250 VGND.n714 7.9105
R4450 VGND.n1243 VGND.n719 7.9105
R4451 VGND.n1242 VGND.n720 7.9105
R4452 VGND.n1241 VGND.n787 7.9105
R4453 VGND.n2416 VGND.n2415 7.9105
R4454 VGND.n137 VGND.n134 7.90638
R4455 VGND.n130 VGND.n129 7.90638
R4456 VGND.n605 VGND.n602 7.90638
R4457 VGND.n598 VGND.n597 7.90638
R4458 VGND.n980 VGND.n975 7.90638
R4459 VGND.n979 VGND.n978 7.90638
R4460 VGND.n167 VGND.n164 7.90638
R4461 VGND.n160 VGND.n159 7.90638
R4462 VGND.n1102 VGND.n1098 7.4049
R4463 VGND.n1075 VGND.n1069 7.4049
R4464 VGND.n1013 VGND.n1007 7.4049
R4465 VGND.n1044 VGND.n1038 7.4049
R4466 VGND VGND.n153 7.12482
R4467 VGND.n101 VGND.n100 6.85473
R4468 VGND.n2856 VGND.n2855 6.85473
R4469 VGND.n2888 VGND.n2887 6.85473
R4470 VGND.n23 VGND.n22 6.77697
R4471 VGND.n52 VGND.n51 6.77697
R4472 VGND.n2936 VGND.n2935 6.77697
R4473 VGND.n2976 VGND.n2975 6.77697
R4474 VGND.n973 VGND.n972 5.27109
R4475 VGND.n77 VGND.n71 5.27109
R4476 VGND.n2573 VGND.n2572 4.5005
R4477 VGND.n2628 VGND.n2585 4.5005
R4478 VGND.n2625 VGND.n2624 4.5005
R4479 VGND.n2622 VGND.n2621 4.5005
R4480 VGND.n2619 VGND.n2618 4.5005
R4481 VGND.n2616 VGND.n2615 4.5005
R4482 VGND.n2613 VGND.n2612 4.5005
R4483 VGND.n2610 VGND.n2609 4.5005
R4484 VGND.n2607 VGND.n2606 4.5005
R4485 VGND.n2604 VGND.n2603 4.5005
R4486 VGND.n2601 VGND.n2600 4.5005
R4487 VGND.n2598 VGND.n2597 4.5005
R4488 VGND.n2595 VGND.n2594 4.5005
R4489 VGND.n2592 VGND.n2591 4.5005
R4490 VGND.n2654 VGND.n227 4.5005
R4491 VGND.n2663 VGND.n226 4.5005
R4492 VGND.n2650 VGND.n221 4.5005
R4493 VGND.n2671 VGND.n220 4.5005
R4494 VGND.n2646 VGND.n215 4.5005
R4495 VGND.n2679 VGND.n214 4.5005
R4496 VGND.n2642 VGND.n209 4.5005
R4497 VGND.n2687 VGND.n208 4.5005
R4498 VGND.n2638 VGND.n203 4.5005
R4499 VGND.n2695 VGND.n202 4.5005
R4500 VGND.n2634 VGND.n197 4.5005
R4501 VGND.n2703 VGND.n196 4.5005
R4502 VGND.n2630 VGND.n2629 4.5005
R4503 VGND.n2712 VGND.n2711 4.5005
R4504 VGND.n2527 VGND.n2526 4.5005
R4505 VGND.n2530 VGND.n2529 4.5005
R4506 VGND.n2533 VGND.n2532 4.5005
R4507 VGND.n2536 VGND.n2535 4.5005
R4508 VGND.n2539 VGND.n2538 4.5005
R4509 VGND.n2542 VGND.n2541 4.5005
R4510 VGND.n2545 VGND.n2544 4.5005
R4511 VGND.n2548 VGND.n2547 4.5005
R4512 VGND.n2551 VGND.n2550 4.5005
R4513 VGND.n2554 VGND.n2553 4.5005
R4514 VGND.n2557 VGND.n2556 4.5005
R4515 VGND.n2560 VGND.n2559 4.5005
R4516 VGND.n2563 VGND.n2562 4.5005
R4517 VGND.n2566 VGND.n2565 4.5005
R4518 VGND.n2569 VGND.n2568 4.5005
R4519 VGND.n2579 VGND.n2571 4.5005
R4520 VGND.n2587 VGND.n2586 4.5005
R4521 VGND.n2590 VGND.n2589 4.5005
R4522 VGND.n2655 VGND.n34 4.5005
R4523 VGND.n824 VGND.n823 4.5005
R4524 VGND.n821 VGND.n820 4.5005
R4525 VGND.n1141 VGND.n1140 4.5005
R4526 VGND.n1153 VGND.n811 4.5005
R4527 VGND.n1160 VGND.n809 4.5005
R4528 VGND.n1157 VGND.n1155 4.5005
R4529 VGND.n1173 VGND.n1172 4.5005
R4530 VGND.n1185 VGND.n803 4.5005
R4531 VGND.n1192 VGND.n801 4.5005
R4532 VGND.n1189 VGND.n1187 4.5005
R4533 VGND.n1205 VGND.n1204 4.5005
R4534 VGND.n1217 VGND.n795 4.5005
R4535 VGND.n1223 VGND.n793 4.5005
R4536 VGND.n1220 VGND.n1219 4.5005
R4537 VGND.n790 VGND.n789 4.5005
R4538 VGND.n827 VGND.n826 4.5005
R4539 VGND.n1125 VGND.n1124 4.5005
R4540 VGND.n1130 VGND.n684 4.5005
R4541 VGND.n816 VGND.n685 4.5005
R4542 VGND.n1143 VGND.n1142 4.5005
R4543 VGND.n1152 VGND.n1151 4.5005
R4544 VGND.n1162 VGND.n1161 4.5005
R4545 VGND.n1156 VGND.n808 4.5005
R4546 VGND.n1175 VGND.n1174 4.5005
R4547 VGND.n1184 VGND.n1183 4.5005
R4548 VGND.n1194 VGND.n1193 4.5005
R4549 VGND.n1188 VGND.n800 4.5005
R4550 VGND.n1207 VGND.n1206 4.5005
R4551 VGND.n1216 VGND.n1215 4.5005
R4552 VGND.n1226 VGND.n1225 4.5005
R4553 VGND.n792 VGND.n788 4.5005
R4554 VGND.n1237 VGND.n1236 4.5005
R4555 VGND.n1117 VGND.n1116 4.41365
R4556 VGND VGND.n3005 4.35375
R4557 VGND.n1094 VGND.n1093 4.05427
R4558 VGND.n587 VGND.n0 4.05427
R4559 VGND.n1002 VGND.n1001 4.05427
R4560 VGND.n1033 VGND.n1032 4.05427
R4561 VGND.n1064 VGND.n1063 4.05427
R4562 VGND VGND.n63 3.99438
R4563 VGND.n2919 VGND 3.99438
R4564 VGND.n2952 VGND 3.99438
R4565 VGND VGND.n2953 3.99437
R4566 VGND VGND.n32 3.99437
R4567 VGND.n1238 VGND.n278 3.77268
R4568 VGND.n3003 VGND.n3002 3.77268
R4569 VGND.n1123 VGND.n1122 3.77268
R4570 VGND.n2715 VGND.n2714 3.77268
R4571 VGND.n1285 VGND.n1284 3.77268
R4572 VGND.n2824 VGND.n192 3.77268
R4573 VGND.n1281 VGND.n691 3.77268
R4574 VGND.n2821 VGND.n2820 3.77268
R4575 VGND.n1276 VGND.n694 3.77268
R4576 VGND.n2819 VGND.n2818 3.77268
R4577 VGND.n1273 VGND.n697 3.77268
R4578 VGND.n2815 VGND.n2814 3.77268
R4579 VGND.n1268 VGND.n700 3.77268
R4580 VGND.n2813 VGND.n2812 3.77268
R4581 VGND.n1265 VGND.n703 3.77268
R4582 VGND.n2809 VGND.n2808 3.77268
R4583 VGND.n1260 VGND.n706 3.77268
R4584 VGND.n2807 VGND.n2806 3.77268
R4585 VGND.n1257 VGND.n709 3.77268
R4586 VGND.n2803 VGND.n2802 3.77268
R4587 VGND.n1252 VGND.n712 3.77268
R4588 VGND.n2801 VGND.n2800 3.77268
R4589 VGND.n1249 VGND.n715 3.77268
R4590 VGND.n2797 VGND.n2796 3.77268
R4591 VGND.n1244 VGND.n718 3.77268
R4592 VGND.n2795 VGND.n2794 3.77268
R4593 VGND.n1224 VGND.n284 3.77268
R4594 VGND.n2791 VGND.n2790 3.77268
R4595 VGND.n1240 VGND.n1239 3.77268
R4596 VGND.n2789 VGND.n2788 3.77268
R4597 VGND.n1287 VGND.n1286 3.77268
R4598 VGND.n2713 VGND.n188 3.77268
R4599 VGND.n2588 VGND.n2587 3.75914
R4600 VGND.n2593 VGND.n2590 3.75914
R4601 VGND.n1221 VGND.n790 3.75914
R4602 VGND.n827 VGND.n825 3.75914
R4603 VGND.n2588 VGND.n2573 3.4105
R4604 VGND.n2628 VGND.n2627 3.4105
R4605 VGND.n2626 VGND.n2625 3.4105
R4606 VGND.n2623 VGND.n2622 3.4105
R4607 VGND.n2620 VGND.n2619 3.4105
R4608 VGND.n2617 VGND.n2616 3.4105
R4609 VGND.n2614 VGND.n2613 3.4105
R4610 VGND.n2611 VGND.n2610 3.4105
R4611 VGND.n2608 VGND.n2607 3.4105
R4612 VGND.n2605 VGND.n2604 3.4105
R4613 VGND.n2602 VGND.n2601 3.4105
R4614 VGND.n2599 VGND.n2598 3.4105
R4615 VGND.n2596 VGND.n2595 3.4105
R4616 VGND.n2593 VGND.n2592 3.4105
R4617 VGND.n3003 VGND.n34 3.4105
R4618 VGND.n2789 VGND.n227 3.4105
R4619 VGND.n2790 VGND.n226 3.4105
R4620 VGND.n2795 VGND.n221 3.4105
R4621 VGND.n2796 VGND.n220 3.4105
R4622 VGND.n2801 VGND.n215 3.4105
R4623 VGND.n2802 VGND.n214 3.4105
R4624 VGND.n2807 VGND.n209 3.4105
R4625 VGND.n2808 VGND.n208 3.4105
R4626 VGND.n2813 VGND.n203 3.4105
R4627 VGND.n2814 VGND.n202 3.4105
R4628 VGND.n2819 VGND.n197 3.4105
R4629 VGND.n2820 VGND.n196 3.4105
R4630 VGND.n2629 VGND.n192 3.4105
R4631 VGND.n2713 VGND.n2712 3.4105
R4632 VGND.n2714 VGND.n2571 3.4105
R4633 VGND.n3002 VGND.n3001 3.4105
R4634 VGND.n2716 VGND.n2715 3.4105
R4635 VGND.n2521 VGND.n240 3.4105
R4636 VGND.n2495 VGND.n35 3.4105
R4637 VGND.n2826 VGND.n2825 3.4105
R4638 VGND.n2824 VGND.n2823 3.4105
R4639 VGND.n379 VGND.n191 3.4105
R4640 VGND.n644 VGND.n643 3.4105
R4641 VGND.n2434 VGND.n264 3.4105
R4642 VGND.n2169 VGND.n2168 3.4105
R4643 VGND.n2507 VGND.n195 3.4105
R4644 VGND.n2822 VGND.n2821 3.4105
R4645 VGND.n2167 VGND.n2166 3.4105
R4646 VGND.n2156 VGND.n2155 3.4105
R4647 VGND.n1438 VGND.n1437 3.4105
R4648 VGND.n2317 VGND.n329 3.4105
R4649 VGND.n2182 VGND.n2181 3.4105
R4650 VGND.n2180 VGND.n2179 3.4105
R4651 VGND.n2506 VGND.n198 3.4105
R4652 VGND.n2818 VGND.n2817 3.4105
R4653 VGND.n2151 VGND.n365 3.4105
R4654 VGND.n2152 VGND.n380 3.4105
R4655 VGND.n2154 VGND.n2153 3.4105
R4656 VGND.n1440 VGND.n1439 3.4105
R4657 VGND.n2129 VGND.n399 3.4105
R4658 VGND.n2150 VGND.n361 3.4105
R4659 VGND.n2193 VGND.n2192 3.4105
R4660 VGND.n2195 VGND.n2194 3.4105
R4661 VGND.n2505 VGND.n201 3.4105
R4662 VGND.n2816 VGND.n2815 3.4105
R4663 VGND.n2021 VGND.n2020 3.4105
R4664 VGND.n2006 VGND.n2005 3.4105
R4665 VGND.n1995 VGND.n1994 3.4105
R4666 VGND.n634 VGND.n384 3.4105
R4667 VGND.n1418 VGND.n642 3.4105
R4668 VGND.n2126 VGND.n400 3.4105
R4669 VGND.n2032 VGND.n2031 3.4105
R4670 VGND.n2149 VGND.n357 3.4105
R4671 VGND.n2208 VGND.n2207 3.4105
R4672 VGND.n2206 VGND.n2205 3.4105
R4673 VGND.n2504 VGND.n204 3.4105
R4674 VGND.n2812 VGND.n2811 3.4105
R4675 VGND.n2034 VGND.n2033 3.4105
R4676 VGND.n2019 VGND.n2018 3.4105
R4677 VGND.n2008 VGND.n2007 3.4105
R4678 VGND.n1993 VGND.n1992 3.4105
R4679 VGND.n1982 VGND.n1981 3.4105
R4680 VGND.n1416 VGND.n1415 3.4105
R4681 VGND.n2342 VGND.n317 3.4105
R4682 VGND.n2045 VGND.n2044 3.4105
R4683 VGND.n2047 VGND.n2046 3.4105
R4684 VGND.n2148 VGND.n353 3.4105
R4685 VGND.n2219 VGND.n2218 3.4105
R4686 VGND.n2221 VGND.n2220 3.4105
R4687 VGND.n2503 VGND.n207 3.4105
R4688 VGND.n2810 VGND.n2809 3.4105
R4689 VGND.n1974 VGND.n420 3.4105
R4690 VGND.n1975 VGND.n424 3.4105
R4691 VGND.n1976 VGND.n428 3.4105
R4692 VGND.n1977 VGND.n432 3.4105
R4693 VGND.n1978 VGND.n436 3.4105
R4694 VGND.n1980 VGND.n1979 3.4105
R4695 VGND.n1414 VGND.n1413 3.4105
R4696 VGND.n1955 VGND.n455 3.4105
R4697 VGND.n1973 VGND.n416 3.4105
R4698 VGND.n2060 VGND.n2059 3.4105
R4699 VGND.n2058 VGND.n2057 3.4105
R4700 VGND.n2147 VGND.n349 3.4105
R4701 VGND.n2234 VGND.n2233 3.4105
R4702 VGND.n2232 VGND.n2231 3.4105
R4703 VGND.n2502 VGND.n210 3.4105
R4704 VGND.n2806 VGND.n2805 3.4105
R4705 VGND.n1884 VGND.n1883 3.4105
R4706 VGND.n1873 VGND.n1872 3.4105
R4707 VGND.n1858 VGND.n1857 3.4105
R4708 VGND.n1847 VGND.n1846 3.4105
R4709 VGND.n1832 VGND.n1831 3.4105
R4710 VGND.n1821 VGND.n1820 3.4105
R4711 VGND.n1408 VGND.n440 3.4105
R4712 VGND.n1393 VGND.n661 3.4105
R4713 VGND.n1952 VGND.n456 3.4105
R4714 VGND.n1899 VGND.n1898 3.4105
R4715 VGND.n1972 VGND.n412 3.4105
R4716 VGND.n2071 VGND.n2070 3.4105
R4717 VGND.n2073 VGND.n2072 3.4105
R4718 VGND.n2146 VGND.n345 3.4105
R4719 VGND.n2245 VGND.n2244 3.4105
R4720 VGND.n2247 VGND.n2246 3.4105
R4721 VGND.n2501 VGND.n213 3.4105
R4722 VGND.n2804 VGND.n2803 3.4105
R4723 VGND.n1897 VGND.n1896 3.4105
R4724 VGND.n1886 VGND.n1885 3.4105
R4725 VGND.n1871 VGND.n1870 3.4105
R4726 VGND.n1860 VGND.n1859 3.4105
R4727 VGND.n1845 VGND.n1844 3.4105
R4728 VGND.n1834 VGND.n1833 3.4105
R4729 VGND.n1819 VGND.n1818 3.4105
R4730 VGND.n1808 VGND.n1807 3.4105
R4731 VGND.n1390 VGND.n1389 3.4105
R4732 VGND.n2367 VGND.n305 3.4105
R4733 VGND.n1912 VGND.n1911 3.4105
R4734 VGND.n1910 VGND.n1909 3.4105
R4735 VGND.n1971 VGND.n408 3.4105
R4736 VGND.n2086 VGND.n2085 3.4105
R4737 VGND.n2084 VGND.n2083 3.4105
R4738 VGND.n2145 VGND.n341 3.4105
R4739 VGND.n2260 VGND.n2259 3.4105
R4740 VGND.n2258 VGND.n2257 3.4105
R4741 VGND.n2500 VGND.n216 3.4105
R4742 VGND.n2800 VGND.n2799 3.4105
R4743 VGND.n1797 VGND.n464 3.4105
R4744 VGND.n1798 VGND.n468 3.4105
R4745 VGND.n1799 VGND.n472 3.4105
R4746 VGND.n1800 VGND.n476 3.4105
R4747 VGND.n1801 VGND.n480 3.4105
R4748 VGND.n1802 VGND.n484 3.4105
R4749 VGND.n1803 VGND.n488 3.4105
R4750 VGND.n1804 VGND.n492 3.4105
R4751 VGND.n1806 VGND.n1805 3.4105
R4752 VGND.n1372 VGND.n574 3.4105
R4753 VGND.n1781 VGND.n511 3.4105
R4754 VGND.n1796 VGND.n460 3.4105
R4755 VGND.n1928 VGND.n1927 3.4105
R4756 VGND.n1930 VGND.n1929 3.4105
R4757 VGND.n1970 VGND.n404 3.4105
R4758 VGND.n2102 VGND.n2101 3.4105
R4759 VGND.n2104 VGND.n2103 3.4105
R4760 VGND.n2144 VGND.n337 3.4105
R4761 VGND.n2276 VGND.n2275 3.4105
R4762 VGND.n2278 VGND.n2277 3.4105
R4763 VGND.n2499 VGND.n219 3.4105
R4764 VGND.n2798 VGND.n2797 3.4105
R4765 VGND.n1756 VGND.n1755 3.4105
R4766 VGND.n1736 VGND.n1735 3.4105
R4767 VGND.n1725 VGND.n1724 3.4105
R4768 VGND.n1710 VGND.n1709 3.4105
R4769 VGND.n1699 VGND.n1698 3.4105
R4770 VGND.n1684 VGND.n1683 3.4105
R4771 VGND.n1673 VGND.n1672 3.4105
R4772 VGND.n1658 VGND.n1657 3.4105
R4773 VGND.n1647 VGND.n1646 3.4105
R4774 VGND.n1530 VGND.n496 3.4105
R4775 VGND.n1533 VGND.n1532 3.4105
R4776 VGND.n1778 VGND.n512 3.4105
R4777 VGND.n2377 VGND.n2376 3.4105
R4778 VGND.n1795 VGND.n297 3.4105
R4779 VGND.n2354 VGND.n2353 3.4105
R4780 VGND.n2352 VGND.n2351 3.4105
R4781 VGND.n1969 VGND.n309 3.4105
R4782 VGND.n2329 VGND.n2328 3.4105
R4783 VGND.n2327 VGND.n2326 3.4105
R4784 VGND.n2143 VGND.n321 3.4105
R4785 VGND.n2304 VGND.n2303 3.4105
R4786 VGND.n2302 VGND.n2301 3.4105
R4787 VGND.n2498 VGND.n222 3.4105
R4788 VGND.n2794 VGND.n2793 3.4105
R4789 VGND.n2379 VGND.n2378 3.4105
R4790 VGND.n1754 VGND.n1753 3.4105
R4791 VGND.n1738 VGND.n1737 3.4105
R4792 VGND.n1723 VGND.n1722 3.4105
R4793 VGND.n1712 VGND.n1711 3.4105
R4794 VGND.n1697 VGND.n1696 3.4105
R4795 VGND.n1686 VGND.n1685 3.4105
R4796 VGND.n1671 VGND.n1670 3.4105
R4797 VGND.n1660 VGND.n1659 3.4105
R4798 VGND.n1645 VGND.n1644 3.4105
R4799 VGND.n1634 VGND.n1633 3.4105
R4800 VGND.n1535 VGND.n1534 3.4105
R4801 VGND.n2392 VGND.n292 3.4105
R4802 VGND.n2380 VGND.n285 3.4105
R4803 VGND.n2375 VGND.n2374 3.4105
R4804 VGND.n2373 VGND.n2372 3.4105
R4805 VGND.n2355 VGND.n300 3.4105
R4806 VGND.n2350 VGND.n2349 3.4105
R4807 VGND.n2348 VGND.n2347 3.4105
R4808 VGND.n2330 VGND.n312 3.4105
R4809 VGND.n2325 VGND.n2324 3.4105
R4810 VGND.n2323 VGND.n2322 3.4105
R4811 VGND.n2305 VGND.n324 3.4105
R4812 VGND.n2300 VGND.n2299 3.4105
R4813 VGND.n2497 VGND.n225 3.4105
R4814 VGND.n2792 VGND.n2791 3.4105
R4815 VGND.n2398 VGND.n2397 3.4105
R4816 VGND.n1621 VGND.n296 3.4105
R4817 VGND.n1622 VGND.n516 3.4105
R4818 VGND.n1623 VGND.n520 3.4105
R4819 VGND.n1624 VGND.n524 3.4105
R4820 VGND.n1625 VGND.n528 3.4105
R4821 VGND.n1626 VGND.n532 3.4105
R4822 VGND.n1627 VGND.n536 3.4105
R4823 VGND.n1628 VGND.n540 3.4105
R4824 VGND.n1629 VGND.n544 3.4105
R4825 VGND.n1630 VGND.n548 3.4105
R4826 VGND.n1632 VGND.n1631 3.4105
R4827 VGND.n1302 VGND.n573 3.4105
R4828 VGND.n1607 VGND.n1606 3.4105
R4829 VGND.n2396 VGND.n2395 3.4105
R4830 VGND.n2394 VGND.n2393 3.4105
R4831 VGND.n514 VGND.n290 3.4105
R4832 VGND.n2371 VGND.n2370 3.4105
R4833 VGND.n2369 VGND.n2368 3.4105
R4834 VGND.n458 VGND.n303 3.4105
R4835 VGND.n2346 VGND.n2345 3.4105
R4836 VGND.n2344 VGND.n2343 3.4105
R4837 VGND.n402 VGND.n315 3.4105
R4838 VGND.n2321 VGND.n2320 3.4105
R4839 VGND.n2319 VGND.n2318 3.4105
R4840 VGND.n2298 VGND.n327 3.4105
R4841 VGND.n2496 VGND.n228 3.4105
R4842 VGND.n2788 VGND.n2787 3.4105
R4843 VGND.n289 VGND.n288 3.4105
R4844 VGND.n2400 VGND.n2399 3.4105
R4845 VGND.n1246 VGND.n1245 3.4105
R4846 VGND.n1248 VGND.n1247 3.4105
R4847 VGND.n1254 VGND.n1253 3.4105
R4848 VGND.n1256 VGND.n1255 3.4105
R4849 VGND.n1262 VGND.n1261 3.4105
R4850 VGND.n1264 VGND.n1263 3.4105
R4851 VGND.n1270 VGND.n1269 3.4105
R4852 VGND.n1272 VGND.n1271 3.4105
R4853 VGND.n1278 VGND.n1277 3.4105
R4854 VGND.n1280 VGND.n1279 3.4105
R4855 VGND.n898 VGND.n552 3.4105
R4856 VGND.n901 VGND.n900 3.4105
R4857 VGND.n2412 VGND.n281 3.4105
R4858 VGND.n899 VGND.n566 3.4105
R4859 VGND.n1548 VGND.n1547 3.4105
R4860 VGND.n1546 VGND.n1545 3.4105
R4861 VGND.n1531 VGND.n567 3.4105
R4862 VGND.n1371 VGND.n1370 3.4105
R4863 VGND.n1388 VGND.n666 3.4105
R4864 VGND.n1410 VGND.n1409 3.4105
R4865 VGND.n1412 VGND.n1411 3.4105
R4866 VGND.n660 VGND.n635 3.4105
R4867 VGND.n1503 VGND.n1502 3.4105
R4868 VGND.n1501 VGND.n1500 3.4105
R4869 VGND.n1436 VGND.n187 3.4105
R4870 VGND.n2830 VGND.n2829 3.4105
R4871 VGND.n2828 VGND.n2827 3.4105
R4872 VGND.n2717 VGND.n188 3.4105
R4873 VGND.n1239 VGND.n788 3.4105
R4874 VGND.n1225 VGND.n1224 3.4105
R4875 VGND.n1216 VGND.n718 3.4105
R4876 VGND.n1206 VGND.n715 3.4105
R4877 VGND.n1188 VGND.n712 3.4105
R4878 VGND.n1193 VGND.n709 3.4105
R4879 VGND.n1184 VGND.n706 3.4105
R4880 VGND.n1174 VGND.n703 3.4105
R4881 VGND.n1156 VGND.n700 3.4105
R4882 VGND.n1161 VGND.n697 3.4105
R4883 VGND.n1152 VGND.n694 3.4105
R4884 VGND.n1142 VGND.n691 3.4105
R4885 VGND.n1285 VGND.n685 3.4105
R4886 VGND.n1286 VGND.n684 3.4105
R4887 VGND.n1238 VGND.n1237 3.4105
R4888 VGND.n1221 VGND.n1220 3.4105
R4889 VGND.n1223 VGND.n1222 3.4105
R4890 VGND.n1218 VGND.n1217 3.4105
R4891 VGND.n1205 VGND.n794 3.4105
R4892 VGND.n1190 VGND.n1189 3.4105
R4893 VGND.n1192 VGND.n1191 3.4105
R4894 VGND.n1186 VGND.n1185 3.4105
R4895 VGND.n1173 VGND.n802 3.4105
R4896 VGND.n1158 VGND.n1157 3.4105
R4897 VGND.n1160 VGND.n1159 3.4105
R4898 VGND.n1154 VGND.n1153 3.4105
R4899 VGND.n1141 VGND.n810 3.4105
R4900 VGND.n822 VGND.n821 3.4105
R4901 VGND.n825 VGND.n824 3.4105
R4902 VGND.n1124 VGND.n1123 3.4105
R4903 VGND.n1241 VGND.n1240 3.4105
R4904 VGND.n1242 VGND.n284 3.4105
R4905 VGND.n1244 VGND.n1243 3.4105
R4906 VGND.n1250 VGND.n1249 3.4105
R4907 VGND.n1252 VGND.n1251 3.4105
R4908 VGND.n1258 VGND.n1257 3.4105
R4909 VGND.n1260 VGND.n1259 3.4105
R4910 VGND.n1266 VGND.n1265 3.4105
R4911 VGND.n1268 VGND.n1267 3.4105
R4912 VGND.n1274 VGND.n1273 3.4105
R4913 VGND.n1276 VGND.n1275 3.4105
R4914 VGND.n1282 VGND.n1281 3.4105
R4915 VGND.n1284 VGND.n1283 3.4105
R4916 VGND.n1288 VGND.n1287 3.4105
R4917 VGND.n1122 VGND.n1121 3.4105
R4918 VGND.n2415 VGND.n278 3.4105
R4919 VGND.n984 VGND.n973 3.01226
R4920 VGND.n78 VGND.n77 3.01226
R4921 VGND.n968 VGND.n903 2.63579
R4922 VGND.n2527 VGND 2.52282
R4923 VGND.n2530 VGND 2.52282
R4924 VGND.n2533 VGND 2.52282
R4925 VGND.n2536 VGND 2.52282
R4926 VGND.n2539 VGND 2.52282
R4927 VGND.n2542 VGND 2.52282
R4928 VGND.n2545 VGND 2.52282
R4929 VGND.n2548 VGND 2.52282
R4930 VGND.n2551 VGND 2.52282
R4931 VGND.n2554 VGND 2.52282
R4932 VGND.n2557 VGND 2.52282
R4933 VGND.n2560 VGND 2.52282
R4934 VGND.n2563 VGND 2.52282
R4935 VGND.n2566 VGND 2.52282
R4936 VGND.n2569 VGND 2.52282
R4937 VGND.n989 VGND.n988 2.25932
R4938 VGND.n109 VGND.n108 2.25932
R4939 VGND.n2864 VGND.n2863 2.25932
R4940 VGND.n2896 VGND.n2895 2.25932
R4941 VGND.n87 VGND.n66 2.25932
R4942 VGND.n83 VGND.n82 2.25932
R4943 VGND.n3033 VGND.n3032 2.19479
R4944 VGND.n139 VGND.n127 1.88285
R4945 VGND.n607 VGND.n595 1.88285
R4946 VGND.n169 VGND.n157 1.88285
R4947 VGND.n3022 VGND.n3021 1.8605
R4948 VGND.n3032 VGND.n3031 1.8605
R4949 VGND.n2570 VGND 1.79514
R4950 VGND.n1118 VGND.n279 1.76378
R4951 VGND.n2570 VGND 1.57193
R4952 VGND.n3004 VGND.n3003 1.54254
R4953 VGND.n3001 VGND.n33 1.54254
R4954 VGND.n2495 VGND.n2436 1.54254
R4955 VGND.n2435 VGND.n2434 1.54254
R4956 VGND.n2317 VGND.n263 1.54254
R4957 VGND.n2129 VGND.n2128 1.54254
R4958 VGND.n2127 VGND.n2126 1.54254
R4959 VGND.n2342 VGND.n318 1.54254
R4960 VGND.n1955 VGND.n1954 1.54254
R4961 VGND.n1953 VGND.n1952 1.54254
R4962 VGND.n2367 VGND.n306 1.54254
R4963 VGND.n1781 VGND.n1780 1.54254
R4964 VGND.n1779 VGND.n1778 1.54254
R4965 VGND.n2392 VGND.n293 1.54254
R4966 VGND.n1607 VGND.n280 1.54254
R4967 VGND.n2413 VGND.n2412 1.54254
R4968 VGND.n1238 VGND.n279 1.54254
R4969 VGND.n2415 VGND.n2414 1.54254
R4970 VGND.n996 VGND.n902 1.50638
R4971 VGND.n2915 VGND.n2914 1.50638
R4972 VGND VGND.n2524 1.3946
R4973 VGND.n2523 VGND 1.3946
R4974 VGND.n2522 VGND 1.3946
R4975 VGND VGND.n241 1.3946
R4976 VGND VGND.n1421 1.3946
R4977 VGND.n1420 VGND 1.3946
R4978 VGND.n1419 VGND 1.3946
R4979 VGND.n1417 VGND 1.3946
R4980 VGND VGND.n645 1.3946
R4981 VGND VGND.n1392 1.3946
R4982 VGND.n1391 VGND 1.3946
R4983 VGND.n1373 VGND 1.3946
R4984 VGND.n1305 VGND 1.3946
R4985 VGND.n1304 VGND 1.3946
R4986 VGND.n1303 VGND 1.3946
R4987 VGND VGND.n673 1.3946
R4988 VGND.n1119 VGND 1.3946
R4989 VGND VGND.n1120 1.3946
R4990 VGND.n1118 VGND.n1117 1.04899
R4991 VGND.n2712 VGND.n2573 1.00149
R4992 VGND.n2629 VGND.n2628 1.00149
R4993 VGND.n2625 VGND.n196 1.00149
R4994 VGND.n2622 VGND.n197 1.00149
R4995 VGND.n2619 VGND.n202 1.00149
R4996 VGND.n2616 VGND.n203 1.00149
R4997 VGND.n2613 VGND.n208 1.00149
R4998 VGND.n2610 VGND.n209 1.00149
R4999 VGND.n2607 VGND.n214 1.00149
R5000 VGND.n2604 VGND.n215 1.00149
R5001 VGND.n2601 VGND.n220 1.00149
R5002 VGND.n2598 VGND.n221 1.00149
R5003 VGND.n2595 VGND.n226 1.00149
R5004 VGND.n2592 VGND.n227 1.00149
R5005 VGND.n2590 VGND.n34 1.00149
R5006 VGND.n824 VGND.n684 1.00149
R5007 VGND.n821 VGND.n685 1.00149
R5008 VGND.n1142 VGND.n1141 1.00149
R5009 VGND.n1153 VGND.n1152 1.00149
R5010 VGND.n1161 VGND.n1160 1.00149
R5011 VGND.n1157 VGND.n1156 1.00149
R5012 VGND.n1174 VGND.n1173 1.00149
R5013 VGND.n1185 VGND.n1184 1.00149
R5014 VGND.n1193 VGND.n1192 1.00149
R5015 VGND.n1189 VGND.n1188 1.00149
R5016 VGND.n1206 VGND.n1205 1.00149
R5017 VGND.n1217 VGND.n1216 1.00149
R5018 VGND.n1225 VGND.n1223 1.00149
R5019 VGND.n1220 VGND.n788 1.00149
R5020 VGND.n1237 VGND.n790 1.00149
R5021 VGND.n1124 VGND.n827 1.00149
R5022 VGND.n2587 VGND.n2571 0.973133
R5023 VGND.n101 VGND.n97 0.929432
R5024 VGND.n2856 VGND.n2852 0.929432
R5025 VGND.n2888 VGND.n2884 0.929432
R5026 VGND.n74 VGND.n72 0.929432
R5027 VGND.n63 VGND.n1 0.916608
R5028 VGND VGND.n2527 0.839786
R5029 VGND VGND.n2530 0.839786
R5030 VGND VGND.n2533 0.839786
R5031 VGND VGND.n2536 0.839786
R5032 VGND VGND.n2539 0.839786
R5033 VGND VGND.n2542 0.839786
R5034 VGND VGND.n2545 0.839786
R5035 VGND VGND.n2548 0.839786
R5036 VGND VGND.n2551 0.839786
R5037 VGND VGND.n2554 0.839786
R5038 VGND VGND.n2557 0.839786
R5039 VGND VGND.n2560 0.839786
R5040 VGND VGND.n2563 0.839786
R5041 VGND VGND.n2566 0.839786
R5042 VGND VGND.n2569 0.839786
R5043 VGND.n121 VGND.n119 0.753441
R5044 VGND.n20 VGND.n18 0.753441
R5045 VGND.n49 VGND.n47 0.753441
R5046 VGND.n2868 VGND.n2845 0.753441
R5047 VGND.n2931 VGND.n2928 0.753441
R5048 VGND.n2973 VGND.n2971 0.753441
R5049 VGND.n3034 VGND.n3033 0.669548
R5050 VGND VGND.n0 0.542567
R5051 VGND.n3034 VGND.n1 0.507317
R5052 VGND.n3005 VGND.n3004 0.404308
R5053 VGND.n1100 VGND.n1097 0.376971
R5054 VGND.n1072 VGND.n1068 0.376971
R5055 VGND.n996 VGND.n995 0.376971
R5056 VGND.n1010 VGND.n1006 0.376971
R5057 VGND.n1041 VGND.n1037 0.376971
R5058 VGND.n88 VGND.n87 0.376971
R5059 VGND.n2914 VGND.n65 0.376971
R5060 VGND VGND.n3034 0.37415
R5061 VGND.n281 VGND.n278 0.362676
R5062 VGND.n1606 VGND.n281 0.362676
R5063 VGND.n1606 VGND.n292 0.362676
R5064 VGND.n512 VGND.n292 0.362676
R5065 VGND.n512 VGND.n511 0.362676
R5066 VGND.n511 VGND.n305 0.362676
R5067 VGND.n456 VGND.n305 0.362676
R5068 VGND.n456 VGND.n455 0.362676
R5069 VGND.n455 VGND.n317 0.362676
R5070 VGND.n400 VGND.n317 0.362676
R5071 VGND.n400 VGND.n399 0.362676
R5072 VGND.n399 VGND.n329 0.362676
R5073 VGND.n329 VGND.n264 0.362676
R5074 VGND.n264 VGND.n35 0.362676
R5075 VGND.n3002 VGND.n35 0.362676
R5076 VGND.n1122 VGND.n901 0.362676
R5077 VGND.n901 VGND.n573 0.362676
R5078 VGND.n1534 VGND.n573 0.362676
R5079 VGND.n1534 VGND.n1533 0.362676
R5080 VGND.n1533 VGND.n574 0.362676
R5081 VGND.n1389 VGND.n574 0.362676
R5082 VGND.n1389 VGND.n661 0.362676
R5083 VGND.n1414 VGND.n661 0.362676
R5084 VGND.n1415 VGND.n1414 0.362676
R5085 VGND.n1415 VGND.n642 0.362676
R5086 VGND.n1439 VGND.n642 0.362676
R5087 VGND.n1439 VGND.n1438 0.362676
R5088 VGND.n1438 VGND.n644 0.362676
R5089 VGND.n644 VGND.n240 0.362676
R5090 VGND.n2715 VGND.n240 0.362676
R5091 VGND.n1284 VGND.n552 0.362676
R5092 VGND.n1632 VGND.n552 0.362676
R5093 VGND.n1633 VGND.n1632 0.362676
R5094 VGND.n1633 VGND.n496 0.362676
R5095 VGND.n1806 VGND.n496 0.362676
R5096 VGND.n1807 VGND.n1806 0.362676
R5097 VGND.n1807 VGND.n440 0.362676
R5098 VGND.n1980 VGND.n440 0.362676
R5099 VGND.n1981 VGND.n1980 0.362676
R5100 VGND.n1981 VGND.n384 0.362676
R5101 VGND.n2154 VGND.n384 0.362676
R5102 VGND.n2155 VGND.n2154 0.362676
R5103 VGND.n2155 VGND.n191 0.362676
R5104 VGND.n2825 VGND.n191 0.362676
R5105 VGND.n2825 VGND.n2824 0.362676
R5106 VGND.n1281 VGND.n1280 0.362676
R5107 VGND.n1280 VGND.n548 0.362676
R5108 VGND.n1645 VGND.n548 0.362676
R5109 VGND.n1646 VGND.n1645 0.362676
R5110 VGND.n1646 VGND.n492 0.362676
R5111 VGND.n1819 VGND.n492 0.362676
R5112 VGND.n1820 VGND.n1819 0.362676
R5113 VGND.n1820 VGND.n436 0.362676
R5114 VGND.n1993 VGND.n436 0.362676
R5115 VGND.n1994 VGND.n1993 0.362676
R5116 VGND.n1994 VGND.n380 0.362676
R5117 VGND.n2167 VGND.n380 0.362676
R5118 VGND.n2168 VGND.n2167 0.362676
R5119 VGND.n2168 VGND.n195 0.362676
R5120 VGND.n2821 VGND.n195 0.362676
R5121 VGND.n1277 VGND.n1276 0.362676
R5122 VGND.n1277 VGND.n544 0.362676
R5123 VGND.n1659 VGND.n544 0.362676
R5124 VGND.n1659 VGND.n1658 0.362676
R5125 VGND.n1658 VGND.n488 0.362676
R5126 VGND.n1833 VGND.n488 0.362676
R5127 VGND.n1833 VGND.n1832 0.362676
R5128 VGND.n1832 VGND.n432 0.362676
R5129 VGND.n2007 VGND.n432 0.362676
R5130 VGND.n2007 VGND.n2006 0.362676
R5131 VGND.n2006 VGND.n365 0.362676
R5132 VGND.n2181 VGND.n365 0.362676
R5133 VGND.n2181 VGND.n2180 0.362676
R5134 VGND.n2180 VGND.n198 0.362676
R5135 VGND.n2818 VGND.n198 0.362676
R5136 VGND.n1273 VGND.n1272 0.362676
R5137 VGND.n1272 VGND.n540 0.362676
R5138 VGND.n1671 VGND.n540 0.362676
R5139 VGND.n1672 VGND.n1671 0.362676
R5140 VGND.n1672 VGND.n484 0.362676
R5141 VGND.n1845 VGND.n484 0.362676
R5142 VGND.n1846 VGND.n1845 0.362676
R5143 VGND.n1846 VGND.n428 0.362676
R5144 VGND.n2019 VGND.n428 0.362676
R5145 VGND.n2020 VGND.n2019 0.362676
R5146 VGND.n2020 VGND.n361 0.362676
R5147 VGND.n2193 VGND.n361 0.362676
R5148 VGND.n2194 VGND.n2193 0.362676
R5149 VGND.n2194 VGND.n201 0.362676
R5150 VGND.n2815 VGND.n201 0.362676
R5151 VGND.n1269 VGND.n1268 0.362676
R5152 VGND.n1269 VGND.n536 0.362676
R5153 VGND.n1685 VGND.n536 0.362676
R5154 VGND.n1685 VGND.n1684 0.362676
R5155 VGND.n1684 VGND.n480 0.362676
R5156 VGND.n1859 VGND.n480 0.362676
R5157 VGND.n1859 VGND.n1858 0.362676
R5158 VGND.n1858 VGND.n424 0.362676
R5159 VGND.n2033 VGND.n424 0.362676
R5160 VGND.n2033 VGND.n2032 0.362676
R5161 VGND.n2032 VGND.n357 0.362676
R5162 VGND.n2207 VGND.n357 0.362676
R5163 VGND.n2207 VGND.n2206 0.362676
R5164 VGND.n2206 VGND.n204 0.362676
R5165 VGND.n2812 VGND.n204 0.362676
R5166 VGND.n1265 VGND.n1264 0.362676
R5167 VGND.n1264 VGND.n532 0.362676
R5168 VGND.n1697 VGND.n532 0.362676
R5169 VGND.n1698 VGND.n1697 0.362676
R5170 VGND.n1698 VGND.n476 0.362676
R5171 VGND.n1871 VGND.n476 0.362676
R5172 VGND.n1872 VGND.n1871 0.362676
R5173 VGND.n1872 VGND.n420 0.362676
R5174 VGND.n2045 VGND.n420 0.362676
R5175 VGND.n2046 VGND.n2045 0.362676
R5176 VGND.n2046 VGND.n353 0.362676
R5177 VGND.n2219 VGND.n353 0.362676
R5178 VGND.n2220 VGND.n2219 0.362676
R5179 VGND.n2220 VGND.n207 0.362676
R5180 VGND.n2809 VGND.n207 0.362676
R5181 VGND.n1261 VGND.n1260 0.362676
R5182 VGND.n1261 VGND.n528 0.362676
R5183 VGND.n1711 VGND.n528 0.362676
R5184 VGND.n1711 VGND.n1710 0.362676
R5185 VGND.n1710 VGND.n472 0.362676
R5186 VGND.n1885 VGND.n472 0.362676
R5187 VGND.n1885 VGND.n1884 0.362676
R5188 VGND.n1884 VGND.n416 0.362676
R5189 VGND.n2059 VGND.n416 0.362676
R5190 VGND.n2059 VGND.n2058 0.362676
R5191 VGND.n2058 VGND.n349 0.362676
R5192 VGND.n2233 VGND.n349 0.362676
R5193 VGND.n2233 VGND.n2232 0.362676
R5194 VGND.n2232 VGND.n210 0.362676
R5195 VGND.n2806 VGND.n210 0.362676
R5196 VGND.n1257 VGND.n1256 0.362676
R5197 VGND.n1256 VGND.n524 0.362676
R5198 VGND.n1723 VGND.n524 0.362676
R5199 VGND.n1724 VGND.n1723 0.362676
R5200 VGND.n1724 VGND.n468 0.362676
R5201 VGND.n1897 VGND.n468 0.362676
R5202 VGND.n1898 VGND.n1897 0.362676
R5203 VGND.n1898 VGND.n412 0.362676
R5204 VGND.n2071 VGND.n412 0.362676
R5205 VGND.n2072 VGND.n2071 0.362676
R5206 VGND.n2072 VGND.n345 0.362676
R5207 VGND.n2245 VGND.n345 0.362676
R5208 VGND.n2246 VGND.n2245 0.362676
R5209 VGND.n2246 VGND.n213 0.362676
R5210 VGND.n2803 VGND.n213 0.362676
R5211 VGND.n1253 VGND.n1252 0.362676
R5212 VGND.n1253 VGND.n520 0.362676
R5213 VGND.n1737 VGND.n520 0.362676
R5214 VGND.n1737 VGND.n1736 0.362676
R5215 VGND.n1736 VGND.n464 0.362676
R5216 VGND.n1911 VGND.n464 0.362676
R5217 VGND.n1911 VGND.n1910 0.362676
R5218 VGND.n1910 VGND.n408 0.362676
R5219 VGND.n2085 VGND.n408 0.362676
R5220 VGND.n2085 VGND.n2084 0.362676
R5221 VGND.n2084 VGND.n341 0.362676
R5222 VGND.n2259 VGND.n341 0.362676
R5223 VGND.n2259 VGND.n2258 0.362676
R5224 VGND.n2258 VGND.n216 0.362676
R5225 VGND.n2800 VGND.n216 0.362676
R5226 VGND.n1249 VGND.n1248 0.362676
R5227 VGND.n1248 VGND.n516 0.362676
R5228 VGND.n1754 VGND.n516 0.362676
R5229 VGND.n1755 VGND.n1754 0.362676
R5230 VGND.n1755 VGND.n460 0.362676
R5231 VGND.n1928 VGND.n460 0.362676
R5232 VGND.n1929 VGND.n1928 0.362676
R5233 VGND.n1929 VGND.n404 0.362676
R5234 VGND.n2102 VGND.n404 0.362676
R5235 VGND.n2103 VGND.n2102 0.362676
R5236 VGND.n2103 VGND.n337 0.362676
R5237 VGND.n2276 VGND.n337 0.362676
R5238 VGND.n2277 VGND.n2276 0.362676
R5239 VGND.n2277 VGND.n219 0.362676
R5240 VGND.n2797 VGND.n219 0.362676
R5241 VGND.n1245 VGND.n1244 0.362676
R5242 VGND.n1245 VGND.n296 0.362676
R5243 VGND.n2378 VGND.n296 0.362676
R5244 VGND.n2378 VGND.n2377 0.362676
R5245 VGND.n2377 VGND.n297 0.362676
R5246 VGND.n2353 VGND.n297 0.362676
R5247 VGND.n2353 VGND.n2352 0.362676
R5248 VGND.n2352 VGND.n309 0.362676
R5249 VGND.n2328 VGND.n309 0.362676
R5250 VGND.n2328 VGND.n2327 0.362676
R5251 VGND.n2327 VGND.n321 0.362676
R5252 VGND.n2303 VGND.n321 0.362676
R5253 VGND.n2303 VGND.n2302 0.362676
R5254 VGND.n2302 VGND.n222 0.362676
R5255 VGND.n2794 VGND.n222 0.362676
R5256 VGND.n2399 VGND.n284 0.362676
R5257 VGND.n2399 VGND.n2398 0.362676
R5258 VGND.n2398 VGND.n285 0.362676
R5259 VGND.n2374 VGND.n285 0.362676
R5260 VGND.n2374 VGND.n2373 0.362676
R5261 VGND.n2373 VGND.n300 0.362676
R5262 VGND.n2349 VGND.n300 0.362676
R5263 VGND.n2349 VGND.n2348 0.362676
R5264 VGND.n2348 VGND.n312 0.362676
R5265 VGND.n2324 VGND.n312 0.362676
R5266 VGND.n2324 VGND.n2323 0.362676
R5267 VGND.n2323 VGND.n324 0.362676
R5268 VGND.n2299 VGND.n324 0.362676
R5269 VGND.n2299 VGND.n225 0.362676
R5270 VGND.n2791 VGND.n225 0.362676
R5271 VGND.n1240 VGND.n289 0.362676
R5272 VGND.n2395 VGND.n289 0.362676
R5273 VGND.n2395 VGND.n2394 0.362676
R5274 VGND.n2394 VGND.n290 0.362676
R5275 VGND.n2370 VGND.n290 0.362676
R5276 VGND.n2370 VGND.n2369 0.362676
R5277 VGND.n2369 VGND.n303 0.362676
R5278 VGND.n2345 VGND.n303 0.362676
R5279 VGND.n2345 VGND.n2344 0.362676
R5280 VGND.n2344 VGND.n315 0.362676
R5281 VGND.n2320 VGND.n315 0.362676
R5282 VGND.n2320 VGND.n2319 0.362676
R5283 VGND.n2319 VGND.n327 0.362676
R5284 VGND.n327 VGND.n228 0.362676
R5285 VGND.n2788 VGND.n228 0.362676
R5286 VGND.n1287 VGND.n566 0.362676
R5287 VGND.n1547 VGND.n566 0.362676
R5288 VGND.n1547 VGND.n1546 0.362676
R5289 VGND.n1546 VGND.n567 0.362676
R5290 VGND.n1370 VGND.n567 0.362676
R5291 VGND.n1370 VGND.n666 0.362676
R5292 VGND.n1410 VGND.n666 0.362676
R5293 VGND.n1411 VGND.n1410 0.362676
R5294 VGND.n1411 VGND.n635 0.362676
R5295 VGND.n1502 VGND.n635 0.362676
R5296 VGND.n1502 VGND.n1501 0.362676
R5297 VGND.n1501 VGND.n187 0.362676
R5298 VGND.n2829 VGND.n187 0.362676
R5299 VGND.n2829 VGND.n2828 0.362676
R5300 VGND.n2828 VGND.n188 0.362676
R5301 VGND.n2627 VGND.n2588 0.349144
R5302 VGND.n2627 VGND.n2626 0.349144
R5303 VGND.n2626 VGND.n2623 0.349144
R5304 VGND.n2623 VGND.n2620 0.349144
R5305 VGND.n2620 VGND.n2617 0.349144
R5306 VGND.n2617 VGND.n2614 0.349144
R5307 VGND.n2614 VGND.n2611 0.349144
R5308 VGND.n2611 VGND.n2608 0.349144
R5309 VGND.n2608 VGND.n2605 0.349144
R5310 VGND.n2605 VGND.n2602 0.349144
R5311 VGND.n2602 VGND.n2599 0.349144
R5312 VGND.n2599 VGND.n2596 0.349144
R5313 VGND.n2596 VGND.n2593 0.349144
R5314 VGND.n1222 VGND.n1221 0.349144
R5315 VGND.n1222 VGND.n1218 0.349144
R5316 VGND.n1218 VGND.n794 0.349144
R5317 VGND.n1190 VGND.n794 0.349144
R5318 VGND.n1191 VGND.n1190 0.349144
R5319 VGND.n1191 VGND.n1186 0.349144
R5320 VGND.n1186 VGND.n802 0.349144
R5321 VGND.n1158 VGND.n802 0.349144
R5322 VGND.n1159 VGND.n1158 0.349144
R5323 VGND.n1159 VGND.n1154 0.349144
R5324 VGND.n1154 VGND.n810 0.349144
R5325 VGND.n822 VGND.n810 0.349144
R5326 VGND.n825 VGND.n822 0.349144
R5327 VGND.n2659 VGND.n2654 0.327628
R5328 VGND.n2663 VGND.n2662 0.327628
R5329 VGND.n2667 VGND.n2650 0.327628
R5330 VGND.n2671 VGND.n2670 0.327628
R5331 VGND.n2675 VGND.n2646 0.327628
R5332 VGND.n2679 VGND.n2678 0.327628
R5333 VGND.n2683 VGND.n2642 0.327628
R5334 VGND.n2687 VGND.n2686 0.327628
R5335 VGND.n2691 VGND.n2638 0.327628
R5336 VGND.n2695 VGND.n2694 0.327628
R5337 VGND.n2699 VGND.n2634 0.327628
R5338 VGND.n2703 VGND.n2702 0.327628
R5339 VGND.n2707 VGND.n2630 0.327628
R5340 VGND.n2711 VGND.n2710 0.327628
R5341 VGND.n2581 VGND.n2579 0.327628
R5342 VGND.n2786 VGND.n2785 0.327628
R5343 VGND.n2782 VGND.n224 0.327628
R5344 VGND.n2777 VGND.n223 0.327628
R5345 VGND.n2772 VGND.n218 0.327628
R5346 VGND.n2767 VGND.n217 0.327628
R5347 VGND.n2762 VGND.n212 0.327628
R5348 VGND.n2757 VGND.n211 0.327628
R5349 VGND.n2752 VGND.n206 0.327628
R5350 VGND.n2747 VGND.n205 0.327628
R5351 VGND.n2742 VGND.n200 0.327628
R5352 VGND.n2737 VGND.n199 0.327628
R5353 VGND.n2732 VGND.n194 0.327628
R5354 VGND.n2727 VGND.n193 0.327628
R5355 VGND.n2722 VGND.n2718 0.327628
R5356 VGND.n239 VGND.n238 0.327628
R5357 VGND.n2491 VGND.n262 0.327628
R5358 VGND.n2486 VGND.n261 0.327628
R5359 VGND.n2481 VGND.n260 0.327628
R5360 VGND.n2476 VGND.n259 0.327628
R5361 VGND.n2471 VGND.n258 0.327628
R5362 VGND.n2466 VGND.n257 0.327628
R5363 VGND.n2461 VGND.n256 0.327628
R5364 VGND.n2456 VGND.n255 0.327628
R5365 VGND.n2451 VGND.n254 0.327628
R5366 VGND.n2446 VGND.n253 0.327628
R5367 VGND.n2441 VGND.n252 0.327628
R5368 VGND.n2508 VGND.n248 0.327628
R5369 VGND.n2511 VGND.n190 0.327628
R5370 VGND.n2516 VGND.n189 0.327628
R5371 VGND.n2520 VGND.n2519 0.327628
R5372 VGND.n2297 VGND.n2296 0.327628
R5373 VGND.n2293 VGND.n333 0.327628
R5374 VGND.n2288 VGND.n332 0.327628
R5375 VGND.n2283 VGND.n2279 0.327628
R5376 VGND.n2256 VGND.n2255 0.327628
R5377 VGND.n2252 VGND.n2248 0.327628
R5378 VGND.n2230 VGND.n2229 0.327628
R5379 VGND.n2226 VGND.n2222 0.327628
R5380 VGND.n2204 VGND.n2203 0.327628
R5381 VGND.n2200 VGND.n2196 0.327628
R5382 VGND.n2178 VGND.n2177 0.327628
R5383 VGND.n2174 VGND.n2170 0.327628
R5384 VGND.n378 VGND.n377 0.327628
R5385 VGND.n2831 VGND.n186 0.327628
R5386 VGND.n2834 VGND.n184 0.327628
R5387 VGND.n2313 VGND.n328 0.327628
R5388 VGND.n2310 VGND.n2306 0.327628
R5389 VGND.n2270 VGND.n331 0.327628
R5390 VGND.n2274 VGND.n2273 0.327628
R5391 VGND.n2265 VGND.n2261 0.327628
R5392 VGND.n2243 VGND.n2242 0.327628
R5393 VGND.n2239 VGND.n2235 0.327628
R5394 VGND.n2217 VGND.n2216 0.327628
R5395 VGND.n2213 VGND.n2209 0.327628
R5396 VGND.n2191 VGND.n2190 0.327628
R5397 VGND.n2187 VGND.n2183 0.327628
R5398 VGND.n2165 VGND.n2164 0.327628
R5399 VGND.n2161 VGND.n2157 0.327628
R5400 VGND.n1435 VGND.n1434 0.327628
R5401 VGND.n1431 VGND.n1424 0.327628
R5402 VGND.n2133 VGND.n326 0.327628
R5403 VGND.n2138 VGND.n325 0.327628
R5404 VGND.n2142 VGND.n2141 0.327628
R5405 VGND.n1450 VGND.n394 0.327628
R5406 VGND.n1455 VGND.n393 0.327628
R5407 VGND.n1460 VGND.n392 0.327628
R5408 VGND.n1465 VGND.n391 0.327628
R5409 VGND.n1470 VGND.n390 0.327628
R5410 VGND.n1475 VGND.n389 0.327628
R5411 VGND.n1480 VGND.n388 0.327628
R5412 VGND.n1485 VGND.n387 0.327628
R5413 VGND.n1490 VGND.n386 0.327628
R5414 VGND.n1495 VGND.n385 0.327628
R5415 VGND.n1499 VGND.n1498 0.327628
R5416 VGND.n1445 VGND.n1441 0.327628
R5417 VGND.n2122 VGND.n403 0.327628
R5418 VGND.n2119 VGND.n323 0.327628
R5419 VGND.n2114 VGND.n322 0.327628
R5420 VGND.n2109 VGND.n2105 0.327628
R5421 VGND.n2082 VGND.n2081 0.327628
R5422 VGND.n2078 VGND.n2074 0.327628
R5423 VGND.n2056 VGND.n2055 0.327628
R5424 VGND.n2052 VGND.n2048 0.327628
R5425 VGND.n2030 VGND.n2029 0.327628
R5426 VGND.n2026 VGND.n2022 0.327628
R5427 VGND.n2004 VGND.n2003 0.327628
R5428 VGND.n2000 VGND.n1996 0.327628
R5429 VGND.n633 VGND.n632 0.327628
R5430 VGND.n1504 VGND.n623 0.327628
R5431 VGND.n1507 VGND.n621 0.327628
R5432 VGND.n2338 VGND.n316 0.327628
R5433 VGND.n2335 VGND.n2331 0.327628
R5434 VGND.n2096 VGND.n320 0.327628
R5435 VGND.n2100 VGND.n2099 0.327628
R5436 VGND.n2091 VGND.n2087 0.327628
R5437 VGND.n2069 VGND.n2068 0.327628
R5438 VGND.n2065 VGND.n2061 0.327628
R5439 VGND.n2043 VGND.n2042 0.327628
R5440 VGND.n2039 VGND.n2035 0.327628
R5441 VGND.n2017 VGND.n2016 0.327628
R5442 VGND.n2013 VGND.n2009 0.327628
R5443 VGND.n1991 VGND.n1990 0.327628
R5444 VGND.n1987 VGND.n1983 0.327628
R5445 VGND.n659 VGND.n658 0.327628
R5446 VGND.n655 VGND.n648 0.327628
R5447 VGND.n1959 VGND.n314 0.327628
R5448 VGND.n1964 VGND.n313 0.327628
R5449 VGND.n1968 VGND.n1967 0.327628
R5450 VGND.n907 VGND.n450 0.327628
R5451 VGND.n912 VGND.n449 0.327628
R5452 VGND.n917 VGND.n448 0.327628
R5453 VGND.n922 VGND.n447 0.327628
R5454 VGND.n927 VGND.n446 0.327628
R5455 VGND.n932 VGND.n445 0.327628
R5456 VGND.n937 VGND.n444 0.327628
R5457 VGND.n942 VGND.n443 0.327628
R5458 VGND.n947 VGND.n442 0.327628
R5459 VGND.n952 VGND.n441 0.327628
R5460 VGND.n957 VGND.n665 0.327628
R5461 VGND.n962 VGND.n664 0.327628
R5462 VGND.n1948 VGND.n459 0.327628
R5463 VGND.n1945 VGND.n311 0.327628
R5464 VGND.n1940 VGND.n310 0.327628
R5465 VGND.n1935 VGND.n1931 0.327628
R5466 VGND.n1908 VGND.n1907 0.327628
R5467 VGND.n1904 VGND.n1900 0.327628
R5468 VGND.n1882 VGND.n1881 0.327628
R5469 VGND.n1878 VGND.n1874 0.327628
R5470 VGND.n1856 VGND.n1855 0.327628
R5471 VGND.n1852 VGND.n1848 0.327628
R5472 VGND.n1830 VGND.n1829 0.327628
R5473 VGND.n1826 VGND.n1822 0.327628
R5474 VGND.n1407 VGND.n1406 0.327628
R5475 VGND.n1403 VGND.n667 0.327628
R5476 VGND.n1398 VGND.n1394 0.327628
R5477 VGND.n2363 VGND.n304 0.327628
R5478 VGND.n2360 VGND.n2356 0.327628
R5479 VGND.n1922 VGND.n308 0.327628
R5480 VGND.n1926 VGND.n1925 0.327628
R5481 VGND.n1917 VGND.n1913 0.327628
R5482 VGND.n1895 VGND.n1894 0.327628
R5483 VGND.n1891 VGND.n1887 0.327628
R5484 VGND.n1869 VGND.n1868 0.327628
R5485 VGND.n1865 VGND.n1861 0.327628
R5486 VGND.n1843 VGND.n1842 0.327628
R5487 VGND.n1839 VGND.n1835 0.327628
R5488 VGND.n1817 VGND.n1816 0.327628
R5489 VGND.n1813 VGND.n1809 0.327628
R5490 VGND.n1387 VGND.n1386 0.327628
R5491 VGND.n1383 VGND.n1376 0.327628
R5492 VGND.n1785 VGND.n302 0.327628
R5493 VGND.n1790 VGND.n301 0.327628
R5494 VGND.n1794 VGND.n1793 0.327628
R5495 VGND.n1320 VGND.n506 0.327628
R5496 VGND.n1325 VGND.n505 0.327628
R5497 VGND.n1330 VGND.n504 0.327628
R5498 VGND.n1335 VGND.n503 0.327628
R5499 VGND.n1340 VGND.n502 0.327628
R5500 VGND.n1345 VGND.n501 0.327628
R5501 VGND.n1350 VGND.n500 0.327628
R5502 VGND.n1355 VGND.n499 0.327628
R5503 VGND.n1360 VGND.n498 0.327628
R5504 VGND.n1365 VGND.n497 0.327628
R5505 VGND.n1369 VGND.n1368 0.327628
R5506 VGND.n1315 VGND.n1308 0.327628
R5507 VGND.n1774 VGND.n515 0.327628
R5508 VGND.n1771 VGND.n299 0.327628
R5509 VGND.n1766 VGND.n298 0.327628
R5510 VGND.n1761 VGND.n1757 0.327628
R5511 VGND.n1734 VGND.n1733 0.327628
R5512 VGND.n1730 VGND.n1726 0.327628
R5513 VGND.n1708 VGND.n1707 0.327628
R5514 VGND.n1704 VGND.n1700 0.327628
R5515 VGND.n1682 VGND.n1681 0.327628
R5516 VGND.n1678 VGND.n1674 0.327628
R5517 VGND.n1656 VGND.n1655 0.327628
R5518 VGND.n1652 VGND.n1648 0.327628
R5519 VGND.n1529 VGND.n1528 0.327628
R5520 VGND.n1525 VGND.n578 0.327628
R5521 VGND.n1520 VGND.n577 0.327628
R5522 VGND.n2388 VGND.n291 0.327628
R5523 VGND.n2385 VGND.n2381 0.327628
R5524 VGND.n1748 VGND.n295 0.327628
R5525 VGND.n1752 VGND.n1751 0.327628
R5526 VGND.n1743 VGND.n1739 0.327628
R5527 VGND.n1721 VGND.n1720 0.327628
R5528 VGND.n1717 VGND.n1713 0.327628
R5529 VGND.n1695 VGND.n1694 0.327628
R5530 VGND.n1691 VGND.n1687 0.327628
R5531 VGND.n1669 VGND.n1668 0.327628
R5532 VGND.n1665 VGND.n1661 0.327628
R5533 VGND.n1643 VGND.n1642 0.327628
R5534 VGND.n1639 VGND.n1635 0.327628
R5535 VGND.n1544 VGND.n1543 0.327628
R5536 VGND.n1540 VGND.n1536 0.327628
R5537 VGND.n1611 VGND.n287 0.327628
R5538 VGND.n1616 VGND.n286 0.327628
R5539 VGND.n1620 VGND.n1619 0.327628
R5540 VGND.n1603 VGND.n562 0.327628
R5541 VGND.n1598 VGND.n561 0.327628
R5542 VGND.n1593 VGND.n560 0.327628
R5543 VGND.n1588 VGND.n559 0.327628
R5544 VGND.n1583 VGND.n558 0.327628
R5545 VGND.n1578 VGND.n557 0.327628
R5546 VGND.n1573 VGND.n556 0.327628
R5547 VGND.n1568 VGND.n555 0.327628
R5548 VGND.n1563 VGND.n554 0.327628
R5549 VGND.n1558 VGND.n553 0.327628
R5550 VGND.n1553 VGND.n1549 0.327628
R5551 VGND.n1301 VGND.n1300 0.327628
R5552 VGND.n2408 VGND.n283 0.327628
R5553 VGND.n2405 VGND.n2401 0.327628
R5554 VGND.n848 VGND.n717 0.327628
R5555 VGND.n853 VGND.n716 0.327628
R5556 VGND.n858 VGND.n711 0.327628
R5557 VGND.n863 VGND.n710 0.327628
R5558 VGND.n868 VGND.n705 0.327628
R5559 VGND.n873 VGND.n704 0.327628
R5560 VGND.n878 VGND.n699 0.327628
R5561 VGND.n883 VGND.n698 0.327628
R5562 VGND.n888 VGND.n693 0.327628
R5563 VGND.n893 VGND.n692 0.327628
R5564 VGND.n897 VGND.n896 0.327628
R5565 VGND.n843 VGND.n831 0.327628
R5566 VGND.n838 VGND.n830 0.327628
R5567 VGND.n1127 VGND.n1125 0.327628
R5568 VGND.n1134 VGND.n1130 0.327628
R5569 VGND.n1137 VGND.n816 0.327628
R5570 VGND.n1147 VGND.n1143 0.327628
R5571 VGND.n1151 VGND.n1150 0.327628
R5572 VGND.n1166 VGND.n1162 0.327628
R5573 VGND.n1169 VGND.n808 0.327628
R5574 VGND.n1179 VGND.n1175 0.327628
R5575 VGND.n1183 VGND.n1182 0.327628
R5576 VGND.n1198 VGND.n1194 0.327628
R5577 VGND.n1201 VGND.n800 0.327628
R5578 VGND.n1211 VGND.n1207 0.327628
R5579 VGND.n1215 VGND.n1214 0.327628
R5580 VGND.n1230 VGND.n1226 0.327628
R5581 VGND.n1233 VGND.n792 0.327628
R5582 VGND.n787 VGND.n786 0.327628
R5583 VGND.n783 VGND.n720 0.327628
R5584 VGND.n778 VGND.n719 0.327628
R5585 VGND.n773 VGND.n714 0.327628
R5586 VGND.n768 VGND.n713 0.327628
R5587 VGND.n763 VGND.n708 0.327628
R5588 VGND.n758 VGND.n707 0.327628
R5589 VGND.n753 VGND.n702 0.327628
R5590 VGND.n748 VGND.n701 0.327628
R5591 VGND.n743 VGND.n696 0.327628
R5592 VGND.n738 VGND.n695 0.327628
R5593 VGND.n733 VGND.n690 0.327628
R5594 VGND.n728 VGND.n689 0.327628
R5595 VGND.n1289 VGND.n683 0.327628
R5596 VGND.n1292 VGND.n681 0.327628
R5597 VGND.n2919 VGND.n63 0.213567
R5598 VGND.n2952 VGND.n2919 0.213567
R5599 VGND.n2953 VGND.n2952 0.213567
R5600 VGND.n2953 VGND.n32 0.213567
R5601 VGND.n1117 VGND.n1094 0.213567
R5602 VGND.n1094 VGND.n1064 0.213567
R5603 VGND.n1064 VGND.n1033 0.213567
R5604 VGND.n1033 VGND.n1002 0.213567
R5605 VGND.n1002 VGND.n0 0.213567
R5606 VGND.n3005 VGND.n32 0.2073
R5607 VGND.n1119 VGND.n1118 0.175967
R5608 VGND.n2714 VGND 0.169807
R5609 VGND.n2713 VGND 0.169807
R5610 VGND VGND.n192 0.169807
R5611 VGND.n2820 VGND 0.169807
R5612 VGND.n2819 VGND 0.169807
R5613 VGND.n2814 VGND 0.169807
R5614 VGND.n2813 VGND 0.169807
R5615 VGND.n2808 VGND 0.169807
R5616 VGND.n2807 VGND 0.169807
R5617 VGND.n2802 VGND 0.169807
R5618 VGND.n2801 VGND 0.169807
R5619 VGND.n2796 VGND 0.169807
R5620 VGND.n2795 VGND 0.169807
R5621 VGND.n2790 VGND 0.169807
R5622 VGND.n2789 VGND 0.169807
R5623 VGND VGND.n2716 0.169807
R5624 VGND.n2717 VGND 0.169807
R5625 VGND.n2823 VGND 0.169807
R5626 VGND.n2822 VGND 0.169807
R5627 VGND.n2817 VGND 0.169807
R5628 VGND.n2816 VGND 0.169807
R5629 VGND.n2811 VGND 0.169807
R5630 VGND.n2810 VGND 0.169807
R5631 VGND.n2805 VGND 0.169807
R5632 VGND.n2804 VGND 0.169807
R5633 VGND.n2799 VGND 0.169807
R5634 VGND.n2798 VGND 0.169807
R5635 VGND.n2793 VGND 0.169807
R5636 VGND.n2792 VGND 0.169807
R5637 VGND.n2787 VGND 0.169807
R5638 VGND.n2521 VGND 0.169807
R5639 VGND.n2827 VGND 0.169807
R5640 VGND.n2826 VGND 0.169807
R5641 VGND.n2507 VGND 0.169807
R5642 VGND.n2506 VGND 0.169807
R5643 VGND.n2505 VGND 0.169807
R5644 VGND.n2504 VGND 0.169807
R5645 VGND.n2503 VGND 0.169807
R5646 VGND.n2502 VGND 0.169807
R5647 VGND.n2501 VGND 0.169807
R5648 VGND.n2500 VGND 0.169807
R5649 VGND.n2499 VGND 0.169807
R5650 VGND.n2498 VGND 0.169807
R5651 VGND.n2497 VGND 0.169807
R5652 VGND.n2496 VGND 0.169807
R5653 VGND.n643 VGND 0.169807
R5654 VGND.n2830 VGND 0.169807
R5655 VGND VGND.n379 0.169807
R5656 VGND.n2169 VGND 0.169807
R5657 VGND.n2179 VGND 0.169807
R5658 VGND.n2195 VGND 0.169807
R5659 VGND.n2205 VGND 0.169807
R5660 VGND.n2221 VGND 0.169807
R5661 VGND.n2231 VGND 0.169807
R5662 VGND.n2247 VGND 0.169807
R5663 VGND.n2257 VGND 0.169807
R5664 VGND.n2278 VGND 0.169807
R5665 VGND.n2301 VGND 0.169807
R5666 VGND.n2300 VGND 0.169807
R5667 VGND.n2298 VGND 0.169807
R5668 VGND.n1437 VGND 0.169807
R5669 VGND.n1436 VGND 0.169807
R5670 VGND.n2156 VGND 0.169807
R5671 VGND.n2166 VGND 0.169807
R5672 VGND.n2182 VGND 0.169807
R5673 VGND.n2192 VGND 0.169807
R5674 VGND.n2208 VGND 0.169807
R5675 VGND.n2218 VGND 0.169807
R5676 VGND.n2234 VGND 0.169807
R5677 VGND.n2244 VGND 0.169807
R5678 VGND.n2260 VGND 0.169807
R5679 VGND.n2275 VGND 0.169807
R5680 VGND VGND.n2304 0.169807
R5681 VGND.n2305 VGND 0.169807
R5682 VGND.n2318 VGND 0.169807
R5683 VGND.n1440 VGND 0.169807
R5684 VGND.n1500 VGND 0.169807
R5685 VGND.n2153 VGND 0.169807
R5686 VGND.n2152 VGND 0.169807
R5687 VGND.n2151 VGND 0.169807
R5688 VGND.n2150 VGND 0.169807
R5689 VGND.n2149 VGND 0.169807
R5690 VGND.n2148 VGND 0.169807
R5691 VGND.n2147 VGND 0.169807
R5692 VGND.n2146 VGND 0.169807
R5693 VGND.n2145 VGND 0.169807
R5694 VGND.n2144 VGND 0.169807
R5695 VGND.n2143 VGND 0.169807
R5696 VGND.n2322 VGND 0.169807
R5697 VGND.n2321 VGND 0.169807
R5698 VGND.n1418 VGND 0.169807
R5699 VGND.n1503 VGND 0.169807
R5700 VGND.n634 VGND 0.169807
R5701 VGND.n1995 VGND 0.169807
R5702 VGND.n2005 VGND 0.169807
R5703 VGND.n2021 VGND 0.169807
R5704 VGND.n2031 VGND 0.169807
R5705 VGND.n2047 VGND 0.169807
R5706 VGND.n2057 VGND 0.169807
R5707 VGND.n2073 VGND 0.169807
R5708 VGND.n2083 VGND 0.169807
R5709 VGND.n2104 VGND 0.169807
R5710 VGND.n2326 VGND 0.169807
R5711 VGND.n2325 VGND 0.169807
R5712 VGND.n402 VGND 0.169807
R5713 VGND.n1416 VGND 0.169807
R5714 VGND.n660 VGND 0.169807
R5715 VGND.n1982 VGND 0.169807
R5716 VGND.n1992 VGND 0.169807
R5717 VGND.n2008 VGND 0.169807
R5718 VGND.n2018 VGND 0.169807
R5719 VGND.n2034 VGND 0.169807
R5720 VGND.n2044 VGND 0.169807
R5721 VGND.n2060 VGND 0.169807
R5722 VGND.n2070 VGND 0.169807
R5723 VGND.n2086 VGND 0.169807
R5724 VGND.n2101 VGND 0.169807
R5725 VGND VGND.n2329 0.169807
R5726 VGND.n2330 VGND 0.169807
R5727 VGND.n2343 VGND 0.169807
R5728 VGND.n1413 VGND 0.169807
R5729 VGND.n1412 VGND 0.169807
R5730 VGND.n1979 VGND 0.169807
R5731 VGND.n1978 VGND 0.169807
R5732 VGND.n1977 VGND 0.169807
R5733 VGND.n1976 VGND 0.169807
R5734 VGND.n1975 VGND 0.169807
R5735 VGND.n1974 VGND 0.169807
R5736 VGND.n1973 VGND 0.169807
R5737 VGND.n1972 VGND 0.169807
R5738 VGND.n1971 VGND 0.169807
R5739 VGND.n1970 VGND 0.169807
R5740 VGND.n1969 VGND 0.169807
R5741 VGND.n2347 VGND 0.169807
R5742 VGND.n2346 VGND 0.169807
R5743 VGND.n1393 VGND 0.169807
R5744 VGND.n1409 VGND 0.169807
R5745 VGND.n1408 VGND 0.169807
R5746 VGND.n1821 VGND 0.169807
R5747 VGND.n1831 VGND 0.169807
R5748 VGND.n1847 VGND 0.169807
R5749 VGND.n1857 VGND 0.169807
R5750 VGND.n1873 VGND 0.169807
R5751 VGND.n1883 VGND 0.169807
R5752 VGND.n1899 VGND 0.169807
R5753 VGND.n1909 VGND 0.169807
R5754 VGND.n1930 VGND 0.169807
R5755 VGND.n2351 VGND 0.169807
R5756 VGND.n2350 VGND 0.169807
R5757 VGND.n458 VGND 0.169807
R5758 VGND.n1390 VGND 0.169807
R5759 VGND.n1388 VGND 0.169807
R5760 VGND.n1808 VGND 0.169807
R5761 VGND.n1818 VGND 0.169807
R5762 VGND.n1834 VGND 0.169807
R5763 VGND.n1844 VGND 0.169807
R5764 VGND.n1860 VGND 0.169807
R5765 VGND.n1870 VGND 0.169807
R5766 VGND.n1886 VGND 0.169807
R5767 VGND.n1896 VGND 0.169807
R5768 VGND.n1912 VGND 0.169807
R5769 VGND.n1927 VGND 0.169807
R5770 VGND VGND.n2354 0.169807
R5771 VGND.n2355 VGND 0.169807
R5772 VGND.n2368 VGND 0.169807
R5773 VGND.n1372 VGND 0.169807
R5774 VGND.n1371 VGND 0.169807
R5775 VGND.n1805 VGND 0.169807
R5776 VGND.n1804 VGND 0.169807
R5777 VGND.n1803 VGND 0.169807
R5778 VGND.n1802 VGND 0.169807
R5779 VGND.n1801 VGND 0.169807
R5780 VGND.n1800 VGND 0.169807
R5781 VGND.n1799 VGND 0.169807
R5782 VGND.n1798 VGND 0.169807
R5783 VGND.n1797 VGND 0.169807
R5784 VGND.n1796 VGND 0.169807
R5785 VGND.n1795 VGND 0.169807
R5786 VGND.n2372 VGND 0.169807
R5787 VGND.n2371 VGND 0.169807
R5788 VGND.n1532 VGND 0.169807
R5789 VGND.n1531 VGND 0.169807
R5790 VGND.n1530 VGND 0.169807
R5791 VGND.n1647 VGND 0.169807
R5792 VGND.n1657 VGND 0.169807
R5793 VGND.n1673 VGND 0.169807
R5794 VGND.n1683 VGND 0.169807
R5795 VGND.n1699 VGND 0.169807
R5796 VGND.n1709 VGND 0.169807
R5797 VGND.n1725 VGND 0.169807
R5798 VGND.n1735 VGND 0.169807
R5799 VGND.n1756 VGND 0.169807
R5800 VGND.n2376 VGND 0.169807
R5801 VGND.n2375 VGND 0.169807
R5802 VGND.n514 VGND 0.169807
R5803 VGND.n1535 VGND 0.169807
R5804 VGND.n1545 VGND 0.169807
R5805 VGND.n1634 VGND 0.169807
R5806 VGND.n1644 VGND 0.169807
R5807 VGND.n1660 VGND 0.169807
R5808 VGND.n1670 VGND 0.169807
R5809 VGND.n1686 VGND 0.169807
R5810 VGND.n1696 VGND 0.169807
R5811 VGND.n1712 VGND 0.169807
R5812 VGND.n1722 VGND 0.169807
R5813 VGND.n1738 VGND 0.169807
R5814 VGND.n1753 VGND 0.169807
R5815 VGND VGND.n2379 0.169807
R5816 VGND.n2380 VGND 0.169807
R5817 VGND.n2393 VGND 0.169807
R5818 VGND.n1302 VGND 0.169807
R5819 VGND.n1548 VGND 0.169807
R5820 VGND.n1631 VGND 0.169807
R5821 VGND.n1630 VGND 0.169807
R5822 VGND.n1629 VGND 0.169807
R5823 VGND.n1628 VGND 0.169807
R5824 VGND.n1627 VGND 0.169807
R5825 VGND.n1626 VGND 0.169807
R5826 VGND.n1625 VGND 0.169807
R5827 VGND.n1624 VGND 0.169807
R5828 VGND.n1623 VGND 0.169807
R5829 VGND.n1622 VGND 0.169807
R5830 VGND.n1621 VGND 0.169807
R5831 VGND.n2397 VGND 0.169807
R5832 VGND.n2396 VGND 0.169807
R5833 VGND.n900 VGND 0.169807
R5834 VGND.n899 VGND 0.169807
R5835 VGND.n898 VGND 0.169807
R5836 VGND.n1279 VGND 0.169807
R5837 VGND.n1278 VGND 0.169807
R5838 VGND.n1271 VGND 0.169807
R5839 VGND.n1270 VGND 0.169807
R5840 VGND.n1263 VGND 0.169807
R5841 VGND.n1262 VGND 0.169807
R5842 VGND.n1255 VGND 0.169807
R5843 VGND.n1254 VGND 0.169807
R5844 VGND.n1247 VGND 0.169807
R5845 VGND.n1246 VGND 0.169807
R5846 VGND.n2400 VGND 0.169807
R5847 VGND.n288 VGND 0.169807
R5848 VGND.n1123 VGND 0.169807
R5849 VGND.n1286 VGND 0.169807
R5850 VGND.n1285 VGND 0.169807
R5851 VGND VGND.n691 0.169807
R5852 VGND VGND.n694 0.169807
R5853 VGND VGND.n697 0.169807
R5854 VGND VGND.n700 0.169807
R5855 VGND VGND.n703 0.169807
R5856 VGND VGND.n706 0.169807
R5857 VGND VGND.n709 0.169807
R5858 VGND VGND.n712 0.169807
R5859 VGND VGND.n715 0.169807
R5860 VGND VGND.n718 0.169807
R5861 VGND.n1224 VGND 0.169807
R5862 VGND.n1239 VGND 0.169807
R5863 VGND.n1121 VGND 0.169807
R5864 VGND.n1288 VGND 0.169807
R5865 VGND.n1283 VGND 0.169807
R5866 VGND.n1282 VGND 0.169807
R5867 VGND.n1275 VGND 0.169807
R5868 VGND.n1274 VGND 0.169807
R5869 VGND.n1267 VGND 0.169807
R5870 VGND.n1266 VGND 0.169807
R5871 VGND.n1259 VGND 0.169807
R5872 VGND.n1258 VGND 0.169807
R5873 VGND.n1251 VGND 0.169807
R5874 VGND.n1250 VGND 0.169807
R5875 VGND.n1243 VGND 0.169807
R5876 VGND.n1242 VGND 0.169807
R5877 VGND.n1241 VGND 0.169807
R5878 VGND.n113 VGND 0.159538
R5879 VGND.n2870 VGND 0.159538
R5880 VGND.n2414 VGND.n279 0.154425
R5881 VGND.n2414 VGND.n2413 0.154425
R5882 VGND.n2413 VGND.n280 0.154425
R5883 VGND.n293 VGND.n280 0.154425
R5884 VGND.n1779 VGND.n293 0.154425
R5885 VGND.n1780 VGND.n1779 0.154425
R5886 VGND.n1780 VGND.n306 0.154425
R5887 VGND.n1953 VGND.n306 0.154425
R5888 VGND.n1954 VGND.n1953 0.154425
R5889 VGND.n1954 VGND.n318 0.154425
R5890 VGND.n2127 VGND.n318 0.154425
R5891 VGND.n2128 VGND.n2127 0.154425
R5892 VGND.n2128 VGND.n263 0.154425
R5893 VGND.n2435 VGND.n263 0.154425
R5894 VGND.n2436 VGND.n2435 0.154425
R5895 VGND.n2436 VGND.n33 0.154425
R5896 VGND.n3004 VGND.n33 0.154425
R5897 VGND.n1120 VGND.n1119 0.154425
R5898 VGND.n1120 VGND.n673 0.154425
R5899 VGND.n1303 VGND.n673 0.154425
R5900 VGND.n1304 VGND.n1303 0.154425
R5901 VGND.n1305 VGND.n1304 0.154425
R5902 VGND.n1373 VGND.n1305 0.154425
R5903 VGND.n1391 VGND.n1373 0.154425
R5904 VGND.n1392 VGND.n1391 0.154425
R5905 VGND.n1392 VGND.n645 0.154425
R5906 VGND.n1417 VGND.n645 0.154425
R5907 VGND.n1419 VGND.n1417 0.154425
R5908 VGND.n1420 VGND.n1419 0.154425
R5909 VGND.n1421 VGND.n1420 0.154425
R5910 VGND.n1421 VGND.n241 0.154425
R5911 VGND.n2522 VGND.n241 0.154425
R5912 VGND.n2523 VGND.n2522 0.154425
R5913 VGND.n2524 VGND.n2523 0.154425
R5914 VGND.n1104 VGND.n1098 0.144904
R5915 VGND.n1077 VGND.n1069 0.144904
R5916 VGND.n1015 VGND.n1007 0.144904
R5917 VGND.n1046 VGND.n1038 0.144904
R5918 VGND.n2571 VGND.n2570 0.138284
R5919 VGND.n2659 VGND.n2658 0.13638
R5920 VGND.n2662 VGND.n2651 0.13638
R5921 VGND.n2667 VGND.n2666 0.13638
R5922 VGND.n2670 VGND.n2647 0.13638
R5923 VGND.n2675 VGND.n2674 0.13638
R5924 VGND.n2678 VGND.n2643 0.13638
R5925 VGND.n2683 VGND.n2682 0.13638
R5926 VGND.n2686 VGND.n2639 0.13638
R5927 VGND.n2691 VGND.n2690 0.13638
R5928 VGND.n2694 VGND.n2635 0.13638
R5929 VGND.n2699 VGND.n2698 0.13638
R5930 VGND.n2702 VGND.n2631 0.13638
R5931 VGND.n2707 VGND.n2706 0.13638
R5932 VGND.n2710 VGND.n2576 0.13638
R5933 VGND.n2581 VGND.n2580 0.13638
R5934 VGND.n2785 VGND.n231 0.13638
R5935 VGND.n2782 VGND.n2781 0.13638
R5936 VGND.n2777 VGND.n2776 0.13638
R5937 VGND.n2772 VGND.n2771 0.13638
R5938 VGND.n2767 VGND.n2766 0.13638
R5939 VGND.n2762 VGND.n2761 0.13638
R5940 VGND.n2757 VGND.n2756 0.13638
R5941 VGND.n2752 VGND.n2751 0.13638
R5942 VGND.n2747 VGND.n2746 0.13638
R5943 VGND.n2742 VGND.n2741 0.13638
R5944 VGND.n2737 VGND.n2736 0.13638
R5945 VGND.n2732 VGND.n2731 0.13638
R5946 VGND.n2727 VGND.n2726 0.13638
R5947 VGND.n2722 VGND.n2721 0.13638
R5948 VGND.n238 VGND.n236 0.13638
R5949 VGND.n2491 VGND.n2490 0.13638
R5950 VGND.n2486 VGND.n2485 0.13638
R5951 VGND.n2481 VGND.n2480 0.13638
R5952 VGND.n2476 VGND.n2475 0.13638
R5953 VGND.n2471 VGND.n2470 0.13638
R5954 VGND.n2466 VGND.n2465 0.13638
R5955 VGND.n2461 VGND.n2460 0.13638
R5956 VGND.n2456 VGND.n2455 0.13638
R5957 VGND.n2451 VGND.n2450 0.13638
R5958 VGND.n2446 VGND.n2445 0.13638
R5959 VGND.n2441 VGND.n2440 0.13638
R5960 VGND.n250 VGND.n248 0.13638
R5961 VGND.n2511 VGND.n2510 0.13638
R5962 VGND.n2516 VGND.n2515 0.13638
R5963 VGND.n2519 VGND.n246 0.13638
R5964 VGND.n2296 VGND.n336 0.13638
R5965 VGND.n2293 VGND.n2292 0.13638
R5966 VGND.n2288 VGND.n2287 0.13638
R5967 VGND.n2283 VGND.n2282 0.13638
R5968 VGND.n2255 VGND.n344 0.13638
R5969 VGND.n2252 VGND.n2251 0.13638
R5970 VGND.n2229 VGND.n352 0.13638
R5971 VGND.n2226 VGND.n2225 0.13638
R5972 VGND.n2203 VGND.n360 0.13638
R5973 VGND.n2200 VGND.n2199 0.13638
R5974 VGND.n2177 VGND.n368 0.13638
R5975 VGND.n2174 VGND.n2173 0.13638
R5976 VGND.n377 VGND.n374 0.13638
R5977 VGND.n370 VGND.n186 0.13638
R5978 VGND.n2834 VGND.n2833 0.13638
R5979 VGND.n2314 VGND.n2313 0.13638
R5980 VGND.n2310 VGND.n2309 0.13638
R5981 VGND.n2270 VGND.n2269 0.13638
R5982 VGND.n2273 VGND.n340 0.13638
R5983 VGND.n2265 VGND.n2264 0.13638
R5984 VGND.n2242 VGND.n348 0.13638
R5985 VGND.n2239 VGND.n2238 0.13638
R5986 VGND.n2216 VGND.n356 0.13638
R5987 VGND.n2213 VGND.n2212 0.13638
R5988 VGND.n2190 VGND.n364 0.13638
R5989 VGND.n2187 VGND.n2186 0.13638
R5990 VGND.n2164 VGND.n383 0.13638
R5991 VGND.n2161 VGND.n2160 0.13638
R5992 VGND.n1434 VGND.n1427 0.13638
R5993 VGND.n1431 VGND.n1430 0.13638
R5994 VGND.n2133 VGND.n2132 0.13638
R5995 VGND.n2138 VGND.n2137 0.13638
R5996 VGND.n2141 VGND.n397 0.13638
R5997 VGND.n1450 VGND.n1449 0.13638
R5998 VGND.n1455 VGND.n1454 0.13638
R5999 VGND.n1460 VGND.n1459 0.13638
R6000 VGND.n1465 VGND.n1464 0.13638
R6001 VGND.n1470 VGND.n1469 0.13638
R6002 VGND.n1475 VGND.n1474 0.13638
R6003 VGND.n1480 VGND.n1479 0.13638
R6004 VGND.n1485 VGND.n1484 0.13638
R6005 VGND.n1490 VGND.n1489 0.13638
R6006 VGND.n1495 VGND.n1494 0.13638
R6007 VGND.n1498 VGND.n638 0.13638
R6008 VGND.n1445 VGND.n1444 0.13638
R6009 VGND.n2123 VGND.n2122 0.13638
R6010 VGND.n2119 VGND.n2118 0.13638
R6011 VGND.n2114 VGND.n2113 0.13638
R6012 VGND.n2109 VGND.n2108 0.13638
R6013 VGND.n2081 VGND.n411 0.13638
R6014 VGND.n2078 VGND.n2077 0.13638
R6015 VGND.n2055 VGND.n419 0.13638
R6016 VGND.n2052 VGND.n2051 0.13638
R6017 VGND.n2029 VGND.n427 0.13638
R6018 VGND.n2026 VGND.n2025 0.13638
R6019 VGND.n2003 VGND.n435 0.13638
R6020 VGND.n2000 VGND.n1999 0.13638
R6021 VGND.n632 VGND.n629 0.13638
R6022 VGND.n625 VGND.n623 0.13638
R6023 VGND.n1507 VGND.n1506 0.13638
R6024 VGND.n2339 VGND.n2338 0.13638
R6025 VGND.n2335 VGND.n2334 0.13638
R6026 VGND.n2096 VGND.n2095 0.13638
R6027 VGND.n2099 VGND.n407 0.13638
R6028 VGND.n2091 VGND.n2090 0.13638
R6029 VGND.n2068 VGND.n415 0.13638
R6030 VGND.n2065 VGND.n2064 0.13638
R6031 VGND.n2042 VGND.n423 0.13638
R6032 VGND.n2039 VGND.n2038 0.13638
R6033 VGND.n2016 VGND.n431 0.13638
R6034 VGND.n2013 VGND.n2012 0.13638
R6035 VGND.n1990 VGND.n439 0.13638
R6036 VGND.n1987 VGND.n1986 0.13638
R6037 VGND.n658 VGND.n651 0.13638
R6038 VGND.n655 VGND.n654 0.13638
R6039 VGND.n1959 VGND.n1958 0.13638
R6040 VGND.n1964 VGND.n1963 0.13638
R6041 VGND.n1967 VGND.n453 0.13638
R6042 VGND.n907 VGND.n906 0.13638
R6043 VGND.n912 VGND.n911 0.13638
R6044 VGND.n917 VGND.n916 0.13638
R6045 VGND.n922 VGND.n921 0.13638
R6046 VGND.n927 VGND.n926 0.13638
R6047 VGND.n932 VGND.n931 0.13638
R6048 VGND.n937 VGND.n936 0.13638
R6049 VGND.n942 VGND.n941 0.13638
R6050 VGND.n947 VGND.n946 0.13638
R6051 VGND.n952 VGND.n951 0.13638
R6052 VGND.n957 VGND.n956 0.13638
R6053 VGND.n962 VGND.n961 0.13638
R6054 VGND.n1949 VGND.n1948 0.13638
R6055 VGND.n1945 VGND.n1944 0.13638
R6056 VGND.n1940 VGND.n1939 0.13638
R6057 VGND.n1935 VGND.n1934 0.13638
R6058 VGND.n1907 VGND.n467 0.13638
R6059 VGND.n1904 VGND.n1903 0.13638
R6060 VGND.n1881 VGND.n475 0.13638
R6061 VGND.n1878 VGND.n1877 0.13638
R6062 VGND.n1855 VGND.n483 0.13638
R6063 VGND.n1852 VGND.n1851 0.13638
R6064 VGND.n1829 VGND.n491 0.13638
R6065 VGND.n1826 VGND.n1825 0.13638
R6066 VGND.n1406 VGND.n670 0.13638
R6067 VGND.n1403 VGND.n1402 0.13638
R6068 VGND.n1398 VGND.n1397 0.13638
R6069 VGND.n2364 VGND.n2363 0.13638
R6070 VGND.n2360 VGND.n2359 0.13638
R6071 VGND.n1922 VGND.n1921 0.13638
R6072 VGND.n1925 VGND.n463 0.13638
R6073 VGND.n1917 VGND.n1916 0.13638
R6074 VGND.n1894 VGND.n471 0.13638
R6075 VGND.n1891 VGND.n1890 0.13638
R6076 VGND.n1868 VGND.n479 0.13638
R6077 VGND.n1865 VGND.n1864 0.13638
R6078 VGND.n1842 VGND.n487 0.13638
R6079 VGND.n1839 VGND.n1838 0.13638
R6080 VGND.n1816 VGND.n495 0.13638
R6081 VGND.n1813 VGND.n1812 0.13638
R6082 VGND.n1386 VGND.n1379 0.13638
R6083 VGND.n1383 VGND.n1382 0.13638
R6084 VGND.n1785 VGND.n1784 0.13638
R6085 VGND.n1790 VGND.n1789 0.13638
R6086 VGND.n1793 VGND.n509 0.13638
R6087 VGND.n1320 VGND.n1319 0.13638
R6088 VGND.n1325 VGND.n1324 0.13638
R6089 VGND.n1330 VGND.n1329 0.13638
R6090 VGND.n1335 VGND.n1334 0.13638
R6091 VGND.n1340 VGND.n1339 0.13638
R6092 VGND.n1345 VGND.n1344 0.13638
R6093 VGND.n1350 VGND.n1349 0.13638
R6094 VGND.n1355 VGND.n1354 0.13638
R6095 VGND.n1360 VGND.n1359 0.13638
R6096 VGND.n1365 VGND.n1364 0.13638
R6097 VGND.n1368 VGND.n1311 0.13638
R6098 VGND.n1315 VGND.n1314 0.13638
R6099 VGND.n1775 VGND.n1774 0.13638
R6100 VGND.n1771 VGND.n1770 0.13638
R6101 VGND.n1766 VGND.n1765 0.13638
R6102 VGND.n1761 VGND.n1760 0.13638
R6103 VGND.n1733 VGND.n523 0.13638
R6104 VGND.n1730 VGND.n1729 0.13638
R6105 VGND.n1707 VGND.n531 0.13638
R6106 VGND.n1704 VGND.n1703 0.13638
R6107 VGND.n1681 VGND.n539 0.13638
R6108 VGND.n1678 VGND.n1677 0.13638
R6109 VGND.n1655 VGND.n547 0.13638
R6110 VGND.n1652 VGND.n1651 0.13638
R6111 VGND.n1528 VGND.n581 0.13638
R6112 VGND.n1525 VGND.n1524 0.13638
R6113 VGND.n1520 VGND.n1519 0.13638
R6114 VGND.n2389 VGND.n2388 0.13638
R6115 VGND.n2385 VGND.n2384 0.13638
R6116 VGND.n1748 VGND.n1747 0.13638
R6117 VGND.n1751 VGND.n519 0.13638
R6118 VGND.n1743 VGND.n1742 0.13638
R6119 VGND.n1720 VGND.n527 0.13638
R6120 VGND.n1717 VGND.n1716 0.13638
R6121 VGND.n1694 VGND.n535 0.13638
R6122 VGND.n1691 VGND.n1690 0.13638
R6123 VGND.n1668 VGND.n543 0.13638
R6124 VGND.n1665 VGND.n1664 0.13638
R6125 VGND.n1642 VGND.n551 0.13638
R6126 VGND.n1639 VGND.n1638 0.13638
R6127 VGND.n1543 VGND.n570 0.13638
R6128 VGND.n1540 VGND.n1539 0.13638
R6129 VGND.n1611 VGND.n1610 0.13638
R6130 VGND.n1616 VGND.n1615 0.13638
R6131 VGND.n1619 VGND.n565 0.13638
R6132 VGND.n1603 VGND.n1602 0.13638
R6133 VGND.n1598 VGND.n1597 0.13638
R6134 VGND.n1593 VGND.n1592 0.13638
R6135 VGND.n1588 VGND.n1587 0.13638
R6136 VGND.n1583 VGND.n1582 0.13638
R6137 VGND.n1578 VGND.n1577 0.13638
R6138 VGND.n1573 VGND.n1572 0.13638
R6139 VGND.n1568 VGND.n1567 0.13638
R6140 VGND.n1563 VGND.n1562 0.13638
R6141 VGND.n1558 VGND.n1557 0.13638
R6142 VGND.n1553 VGND.n1552 0.13638
R6143 VGND.n1300 VGND.n678 0.13638
R6144 VGND.n2409 VGND.n2408 0.13638
R6145 VGND.n2405 VGND.n2404 0.13638
R6146 VGND.n848 VGND.n847 0.13638
R6147 VGND.n853 VGND.n852 0.13638
R6148 VGND.n858 VGND.n857 0.13638
R6149 VGND.n863 VGND.n862 0.13638
R6150 VGND.n868 VGND.n867 0.13638
R6151 VGND.n873 VGND.n872 0.13638
R6152 VGND.n878 VGND.n877 0.13638
R6153 VGND.n883 VGND.n882 0.13638
R6154 VGND.n888 VGND.n887 0.13638
R6155 VGND.n893 VGND.n892 0.13638
R6156 VGND.n896 VGND.n834 0.13638
R6157 VGND.n843 VGND.n842 0.13638
R6158 VGND.n838 VGND.n837 0.13638
R6159 VGND.n1128 VGND.n1127 0.13638
R6160 VGND.n1134 VGND.n1133 0.13638
R6161 VGND.n1138 VGND.n1137 0.13638
R6162 VGND.n1147 VGND.n1146 0.13638
R6163 VGND.n1150 VGND.n814 0.13638
R6164 VGND.n1166 VGND.n1165 0.13638
R6165 VGND.n1170 VGND.n1169 0.13638
R6166 VGND.n1179 VGND.n1178 0.13638
R6167 VGND.n1182 VGND.n806 0.13638
R6168 VGND.n1198 VGND.n1197 0.13638
R6169 VGND.n1202 VGND.n1201 0.13638
R6170 VGND.n1211 VGND.n1210 0.13638
R6171 VGND.n1214 VGND.n798 0.13638
R6172 VGND.n1230 VGND.n1229 0.13638
R6173 VGND.n1234 VGND.n1233 0.13638
R6174 VGND.n786 VGND.n723 0.13638
R6175 VGND.n783 VGND.n782 0.13638
R6176 VGND.n778 VGND.n777 0.13638
R6177 VGND.n773 VGND.n772 0.13638
R6178 VGND.n768 VGND.n767 0.13638
R6179 VGND.n763 VGND.n762 0.13638
R6180 VGND.n758 VGND.n757 0.13638
R6181 VGND.n753 VGND.n752 0.13638
R6182 VGND.n748 VGND.n747 0.13638
R6183 VGND.n743 VGND.n742 0.13638
R6184 VGND.n738 VGND.n737 0.13638
R6185 VGND.n733 VGND.n732 0.13638
R6186 VGND.n728 VGND.n727 0.13638
R6187 VGND.n687 VGND.n683 0.13638
R6188 VGND.n1292 VGND.n1291 0.13638
R6189 VGND VGND.n113 0.120838
R6190 VGND.n1112 VGND.n1111 0.120292
R6191 VGND.n1111 VGND.n1110 0.120292
R6192 VGND.n1110 VGND.n1096 0.120292
R6193 VGND.n1106 VGND.n1096 0.120292
R6194 VGND.n1106 VGND.n1105 0.120292
R6195 VGND.n1105 VGND.n1104 0.120292
R6196 VGND.n1090 VGND.n1089 0.120292
R6197 VGND.n1085 VGND.n1084 0.120292
R6198 VGND.n1084 VGND.n1083 0.120292
R6199 VGND.n1083 VGND.n1067 0.120292
R6200 VGND.n1079 VGND.n1067 0.120292
R6201 VGND.n1079 VGND.n1078 0.120292
R6202 VGND.n1078 VGND.n1077 0.120292
R6203 VGND.n147 VGND.n124 0.120292
R6204 VGND.n141 VGND.n124 0.120292
R6205 VGND.n141 VGND.n140 0.120292
R6206 VGND.n140 VGND.n128 0.120292
R6207 VGND.n133 VGND.n128 0.120292
R6208 VGND.n133 VGND.n132 0.120292
R6209 VGND.n132 VGND.n131 0.120292
R6210 VGND.n590 VGND.n587 0.120292
R6211 VGND.n591 VGND.n590 0.120292
R6212 VGND.n615 VGND.n592 0.120292
R6213 VGND.n609 VGND.n592 0.120292
R6214 VGND.n609 VGND.n608 0.120292
R6215 VGND.n608 VGND.n596 0.120292
R6216 VGND.n601 VGND.n596 0.120292
R6217 VGND.n601 VGND.n600 0.120292
R6218 VGND.n600 VGND.n599 0.120292
R6219 VGND.n998 VGND.n997 0.120292
R6220 VGND.n991 VGND.n967 0.120292
R6221 VGND.n986 VGND.n967 0.120292
R6222 VGND.n986 VGND.n985 0.120292
R6223 VGND.n982 VGND.n981 0.120292
R6224 VGND.n981 VGND.n976 0.120292
R6225 VGND.n977 VGND.n976 0.120292
R6226 VGND.n1028 VGND.n1027 0.120292
R6227 VGND.n1023 VGND.n1022 0.120292
R6228 VGND.n1022 VGND.n1021 0.120292
R6229 VGND.n1021 VGND.n1005 0.120292
R6230 VGND.n1017 VGND.n1005 0.120292
R6231 VGND.n1017 VGND.n1016 0.120292
R6232 VGND.n1016 VGND.n1015 0.120292
R6233 VGND.n1059 VGND.n1058 0.120292
R6234 VGND.n1054 VGND.n1053 0.120292
R6235 VGND.n1053 VGND.n1052 0.120292
R6236 VGND.n1052 VGND.n1036 0.120292
R6237 VGND.n1048 VGND.n1036 0.120292
R6238 VGND.n1048 VGND.n1047 0.120292
R6239 VGND.n1047 VGND.n1046 0.120292
R6240 VGND.n177 VGND.n154 0.120292
R6241 VGND.n171 VGND.n154 0.120292
R6242 VGND.n171 VGND.n170 0.120292
R6243 VGND.n170 VGND.n158 0.120292
R6244 VGND.n163 VGND.n158 0.120292
R6245 VGND.n163 VGND.n162 0.120292
R6246 VGND.n162 VGND.n161 0.120292
R6247 VGND.n19 VGND.n15 0.120292
R6248 VGND.n24 VGND.n15 0.120292
R6249 VGND.n25 VGND.n24 0.120292
R6250 VGND.n26 VGND.n25 0.120292
R6251 VGND.n26 VGND.n13 0.120292
R6252 VGND.n30 VGND.n13 0.120292
R6253 VGND.n31 VGND.n30 0.120292
R6254 VGND.n105 VGND.n97 0.120292
R6255 VGND.n106 VGND.n105 0.120292
R6256 VGND.n106 VGND.n91 0.120292
R6257 VGND.n111 VGND.n91 0.120292
R6258 VGND.n112 VGND.n111 0.120292
R6259 VGND.n2860 VGND.n2852 0.120292
R6260 VGND.n2861 VGND.n2860 0.120292
R6261 VGND.n2861 VGND.n2846 0.120292
R6262 VGND.n2866 VGND.n2846 0.120292
R6263 VGND.n2867 VGND.n2866 0.120292
R6264 VGND.n2892 VGND.n2884 0.120292
R6265 VGND.n2893 VGND.n2892 0.120292
R6266 VGND.n2893 VGND.n2878 0.120292
R6267 VGND.n2898 VGND.n2878 0.120292
R6268 VGND.n2899 VGND.n2898 0.120292
R6269 VGND.n2903 VGND.n2900 0.120292
R6270 VGND.n79 VGND.n72 0.120292
R6271 VGND.n80 VGND.n79 0.120292
R6272 VGND.n80 VGND.n67 0.120292
R6273 VGND.n85 VGND.n67 0.120292
R6274 VGND.n86 VGND.n85 0.120292
R6275 VGND.n2918 VGND.n64 0.120292
R6276 VGND.n2933 VGND.n2932 0.120292
R6277 VGND.n2933 VGND.n2925 0.120292
R6278 VGND.n2938 VGND.n2925 0.120292
R6279 VGND.n2939 VGND.n2938 0.120292
R6280 VGND.n2940 VGND.n2939 0.120292
R6281 VGND.n2940 VGND.n2923 0.120292
R6282 VGND.n2944 VGND.n2923 0.120292
R6283 VGND.n2946 VGND.n2920 0.120292
R6284 VGND.n2951 VGND.n2920 0.120292
R6285 VGND.n48 VGND.n42 0.120292
R6286 VGND.n53 VGND.n42 0.120292
R6287 VGND.n54 VGND.n53 0.120292
R6288 VGND.n55 VGND.n54 0.120292
R6289 VGND.n55 VGND.n40 0.120292
R6290 VGND.n59 VGND.n40 0.120292
R6291 VGND.n60 VGND.n59 0.120292
R6292 VGND.n2958 VGND.n2957 0.120292
R6293 VGND.n2957 VGND.n2956 0.120292
R6294 VGND.n2972 VGND.n2966 0.120292
R6295 VGND.n2977 VGND.n2966 0.120292
R6296 VGND.n2978 VGND.n2977 0.120292
R6297 VGND.n2979 VGND.n2978 0.120292
R6298 VGND.n2979 VGND.n2964 0.120292
R6299 VGND.n2983 VGND.n2964 0.120292
R6300 VGND.n2984 VGND.n2983 0.120292
R6301 VGND.n2990 VGND.n2989 0.120292
R6302 VGND.n2989 VGND.n2988 0.120292
R6303 VGND VGND.n2870 0.119536
R6304 VGND.n1098 VGND 0.117202
R6305 VGND.n1069 VGND 0.117202
R6306 VGND.n1007 VGND 0.117202
R6307 VGND.n1038 VGND 0.117202
R6308 VGND.n231 VGND.n230 0.110872
R6309 VGND.n2781 VGND.n2780 0.110872
R6310 VGND.n2776 VGND.n2775 0.110872
R6311 VGND.n2771 VGND.n2770 0.110872
R6312 VGND.n2766 VGND.n2765 0.110872
R6313 VGND.n2761 VGND.n2760 0.110872
R6314 VGND.n2756 VGND.n2755 0.110872
R6315 VGND.n2751 VGND.n2750 0.110872
R6316 VGND.n2746 VGND.n2745 0.110872
R6317 VGND.n2741 VGND.n2740 0.110872
R6318 VGND.n2736 VGND.n2735 0.110872
R6319 VGND.n2731 VGND.n2730 0.110872
R6320 VGND.n2726 VGND.n2725 0.110872
R6321 VGND.n2721 VGND.n2720 0.110872
R6322 VGND.n236 VGND.n235 0.110872
R6323 VGND.n2490 VGND.n2489 0.110872
R6324 VGND.n2485 VGND.n2484 0.110872
R6325 VGND.n2480 VGND.n2479 0.110872
R6326 VGND.n2475 VGND.n2474 0.110872
R6327 VGND.n2470 VGND.n2469 0.110872
R6328 VGND.n2465 VGND.n2464 0.110872
R6329 VGND.n2460 VGND.n2459 0.110872
R6330 VGND.n2455 VGND.n2454 0.110872
R6331 VGND.n2450 VGND.n2449 0.110872
R6332 VGND.n2445 VGND.n2444 0.110872
R6333 VGND.n2440 VGND.n2439 0.110872
R6334 VGND.n251 VGND.n250 0.110872
R6335 VGND.n2510 VGND.n2509 0.110872
R6336 VGND.n2515 VGND.n2514 0.110872
R6337 VGND.n246 VGND.n245 0.110872
R6338 VGND.n336 VGND.n335 0.110872
R6339 VGND.n2292 VGND.n2291 0.110872
R6340 VGND.n2287 VGND.n2286 0.110872
R6341 VGND.n2282 VGND.n2281 0.110872
R6342 VGND.n344 VGND.n343 0.110872
R6343 VGND.n2251 VGND.n2250 0.110872
R6344 VGND.n352 VGND.n351 0.110872
R6345 VGND.n2225 VGND.n2224 0.110872
R6346 VGND.n360 VGND.n359 0.110872
R6347 VGND.n2199 VGND.n2198 0.110872
R6348 VGND.n368 VGND.n367 0.110872
R6349 VGND.n2173 VGND.n2172 0.110872
R6350 VGND.n374 VGND.n373 0.110872
R6351 VGND.n371 VGND.n370 0.110872
R6352 VGND.n2833 VGND.n2832 0.110872
R6353 VGND.n2315 VGND.n2314 0.110872
R6354 VGND.n2309 VGND.n2308 0.110872
R6355 VGND.n2269 VGND.n2268 0.110872
R6356 VGND.n340 VGND.n339 0.110872
R6357 VGND.n2264 VGND.n2263 0.110872
R6358 VGND.n348 VGND.n347 0.110872
R6359 VGND.n2238 VGND.n2237 0.110872
R6360 VGND.n356 VGND.n355 0.110872
R6361 VGND.n2212 VGND.n2211 0.110872
R6362 VGND.n364 VGND.n363 0.110872
R6363 VGND.n2186 VGND.n2185 0.110872
R6364 VGND.n383 VGND.n382 0.110872
R6365 VGND.n2160 VGND.n2159 0.110872
R6366 VGND.n1427 VGND.n1426 0.110872
R6367 VGND.n1430 VGND.n1429 0.110872
R6368 VGND.n2132 VGND.n2131 0.110872
R6369 VGND.n2137 VGND.n2136 0.110872
R6370 VGND.n397 VGND.n396 0.110872
R6371 VGND.n1449 VGND.n1448 0.110872
R6372 VGND.n1454 VGND.n1453 0.110872
R6373 VGND.n1459 VGND.n1458 0.110872
R6374 VGND.n1464 VGND.n1463 0.110872
R6375 VGND.n1469 VGND.n1468 0.110872
R6376 VGND.n1474 VGND.n1473 0.110872
R6377 VGND.n1479 VGND.n1478 0.110872
R6378 VGND.n1484 VGND.n1483 0.110872
R6379 VGND.n1489 VGND.n1488 0.110872
R6380 VGND.n1494 VGND.n1493 0.110872
R6381 VGND.n638 VGND.n637 0.110872
R6382 VGND.n1444 VGND.n1443 0.110872
R6383 VGND.n2124 VGND.n2123 0.110872
R6384 VGND.n2118 VGND.n2117 0.110872
R6385 VGND.n2113 VGND.n2112 0.110872
R6386 VGND.n2108 VGND.n2107 0.110872
R6387 VGND.n411 VGND.n410 0.110872
R6388 VGND.n2077 VGND.n2076 0.110872
R6389 VGND.n419 VGND.n418 0.110872
R6390 VGND.n2051 VGND.n2050 0.110872
R6391 VGND.n427 VGND.n426 0.110872
R6392 VGND.n2025 VGND.n2024 0.110872
R6393 VGND.n435 VGND.n434 0.110872
R6394 VGND.n1999 VGND.n1998 0.110872
R6395 VGND.n629 VGND.n628 0.110872
R6396 VGND.n626 VGND.n625 0.110872
R6397 VGND.n1506 VGND.n1505 0.110872
R6398 VGND.n2340 VGND.n2339 0.110872
R6399 VGND.n2334 VGND.n2333 0.110872
R6400 VGND.n2095 VGND.n2094 0.110872
R6401 VGND.n407 VGND.n406 0.110872
R6402 VGND.n2090 VGND.n2089 0.110872
R6403 VGND.n415 VGND.n414 0.110872
R6404 VGND.n2064 VGND.n2063 0.110872
R6405 VGND.n423 VGND.n422 0.110872
R6406 VGND.n2038 VGND.n2037 0.110872
R6407 VGND.n431 VGND.n430 0.110872
R6408 VGND.n2012 VGND.n2011 0.110872
R6409 VGND.n439 VGND.n438 0.110872
R6410 VGND.n1986 VGND.n1985 0.110872
R6411 VGND.n651 VGND.n650 0.110872
R6412 VGND.n654 VGND.n653 0.110872
R6413 VGND.n1958 VGND.n1957 0.110872
R6414 VGND.n1963 VGND.n1962 0.110872
R6415 VGND.n453 VGND.n452 0.110872
R6416 VGND.n906 VGND.n905 0.110872
R6417 VGND.n911 VGND.n910 0.110872
R6418 VGND.n916 VGND.n915 0.110872
R6419 VGND.n921 VGND.n920 0.110872
R6420 VGND.n926 VGND.n925 0.110872
R6421 VGND.n931 VGND.n930 0.110872
R6422 VGND.n936 VGND.n935 0.110872
R6423 VGND.n941 VGND.n940 0.110872
R6424 VGND.n946 VGND.n945 0.110872
R6425 VGND.n951 VGND.n950 0.110872
R6426 VGND.n956 VGND.n955 0.110872
R6427 VGND.n961 VGND.n960 0.110872
R6428 VGND.n1950 VGND.n1949 0.110872
R6429 VGND.n1944 VGND.n1943 0.110872
R6430 VGND.n1939 VGND.n1938 0.110872
R6431 VGND.n1934 VGND.n1933 0.110872
R6432 VGND.n467 VGND.n466 0.110872
R6433 VGND.n1903 VGND.n1902 0.110872
R6434 VGND.n475 VGND.n474 0.110872
R6435 VGND.n1877 VGND.n1876 0.110872
R6436 VGND.n483 VGND.n482 0.110872
R6437 VGND.n1851 VGND.n1850 0.110872
R6438 VGND.n491 VGND.n490 0.110872
R6439 VGND.n1825 VGND.n1824 0.110872
R6440 VGND.n670 VGND.n669 0.110872
R6441 VGND.n1402 VGND.n1401 0.110872
R6442 VGND.n1397 VGND.n1396 0.110872
R6443 VGND.n2365 VGND.n2364 0.110872
R6444 VGND.n2359 VGND.n2358 0.110872
R6445 VGND.n1921 VGND.n1920 0.110872
R6446 VGND.n463 VGND.n462 0.110872
R6447 VGND.n1916 VGND.n1915 0.110872
R6448 VGND.n471 VGND.n470 0.110872
R6449 VGND.n1890 VGND.n1889 0.110872
R6450 VGND.n479 VGND.n478 0.110872
R6451 VGND.n1864 VGND.n1863 0.110872
R6452 VGND.n487 VGND.n486 0.110872
R6453 VGND.n1838 VGND.n1837 0.110872
R6454 VGND.n495 VGND.n494 0.110872
R6455 VGND.n1812 VGND.n1811 0.110872
R6456 VGND.n1379 VGND.n1378 0.110872
R6457 VGND.n1382 VGND.n1381 0.110872
R6458 VGND.n1784 VGND.n1783 0.110872
R6459 VGND.n1789 VGND.n1788 0.110872
R6460 VGND.n509 VGND.n508 0.110872
R6461 VGND.n1319 VGND.n1318 0.110872
R6462 VGND.n1324 VGND.n1323 0.110872
R6463 VGND.n1329 VGND.n1328 0.110872
R6464 VGND.n1334 VGND.n1333 0.110872
R6465 VGND.n1339 VGND.n1338 0.110872
R6466 VGND.n1344 VGND.n1343 0.110872
R6467 VGND.n1349 VGND.n1348 0.110872
R6468 VGND.n1354 VGND.n1353 0.110872
R6469 VGND.n1359 VGND.n1358 0.110872
R6470 VGND.n1364 VGND.n1363 0.110872
R6471 VGND.n1311 VGND.n1310 0.110872
R6472 VGND.n1314 VGND.n1313 0.110872
R6473 VGND.n1776 VGND.n1775 0.110872
R6474 VGND.n1770 VGND.n1769 0.110872
R6475 VGND.n1765 VGND.n1764 0.110872
R6476 VGND.n1760 VGND.n1759 0.110872
R6477 VGND.n523 VGND.n522 0.110872
R6478 VGND.n1729 VGND.n1728 0.110872
R6479 VGND.n531 VGND.n530 0.110872
R6480 VGND.n1703 VGND.n1702 0.110872
R6481 VGND.n539 VGND.n538 0.110872
R6482 VGND.n1677 VGND.n1676 0.110872
R6483 VGND.n547 VGND.n546 0.110872
R6484 VGND.n1651 VGND.n1650 0.110872
R6485 VGND.n581 VGND.n580 0.110872
R6486 VGND.n1524 VGND.n1523 0.110872
R6487 VGND.n1519 VGND.n1518 0.110872
R6488 VGND.n2390 VGND.n2389 0.110872
R6489 VGND.n2384 VGND.n2383 0.110872
R6490 VGND.n1747 VGND.n1746 0.110872
R6491 VGND.n519 VGND.n518 0.110872
R6492 VGND.n1742 VGND.n1741 0.110872
R6493 VGND.n527 VGND.n526 0.110872
R6494 VGND.n1716 VGND.n1715 0.110872
R6495 VGND.n535 VGND.n534 0.110872
R6496 VGND.n1690 VGND.n1689 0.110872
R6497 VGND.n543 VGND.n542 0.110872
R6498 VGND.n1664 VGND.n1663 0.110872
R6499 VGND.n551 VGND.n550 0.110872
R6500 VGND.n1638 VGND.n1637 0.110872
R6501 VGND.n570 VGND.n569 0.110872
R6502 VGND.n1539 VGND.n1538 0.110872
R6503 VGND.n1610 VGND.n1609 0.110872
R6504 VGND.n1615 VGND.n1614 0.110872
R6505 VGND.n565 VGND.n564 0.110872
R6506 VGND.n1602 VGND.n1601 0.110872
R6507 VGND.n1597 VGND.n1596 0.110872
R6508 VGND.n1592 VGND.n1591 0.110872
R6509 VGND.n1587 VGND.n1586 0.110872
R6510 VGND.n1582 VGND.n1581 0.110872
R6511 VGND.n1577 VGND.n1576 0.110872
R6512 VGND.n1572 VGND.n1571 0.110872
R6513 VGND.n1567 VGND.n1566 0.110872
R6514 VGND.n1562 VGND.n1561 0.110872
R6515 VGND.n1557 VGND.n1556 0.110872
R6516 VGND.n1552 VGND.n1551 0.110872
R6517 VGND.n678 VGND.n677 0.110872
R6518 VGND.n2410 VGND.n2409 0.110872
R6519 VGND.n2404 VGND.n2403 0.110872
R6520 VGND.n847 VGND.n846 0.110872
R6521 VGND.n852 VGND.n851 0.110872
R6522 VGND.n857 VGND.n856 0.110872
R6523 VGND.n862 VGND.n861 0.110872
R6524 VGND.n867 VGND.n866 0.110872
R6525 VGND.n872 VGND.n871 0.110872
R6526 VGND.n877 VGND.n876 0.110872
R6527 VGND.n882 VGND.n881 0.110872
R6528 VGND.n887 VGND.n886 0.110872
R6529 VGND.n892 VGND.n891 0.110872
R6530 VGND.n834 VGND.n833 0.110872
R6531 VGND.n842 VGND.n841 0.110872
R6532 VGND.n837 VGND.n836 0.110872
R6533 VGND.n1129 VGND.n1128 0.110872
R6534 VGND.n1133 VGND.n1132 0.110872
R6535 VGND.n1139 VGND.n1138 0.110872
R6536 VGND.n1146 VGND.n1145 0.110872
R6537 VGND.n814 VGND.n813 0.110872
R6538 VGND.n1165 VGND.n1164 0.110872
R6539 VGND.n1171 VGND.n1170 0.110872
R6540 VGND.n1178 VGND.n1177 0.110872
R6541 VGND.n806 VGND.n805 0.110872
R6542 VGND.n1197 VGND.n1196 0.110872
R6543 VGND.n1203 VGND.n1202 0.110872
R6544 VGND.n1210 VGND.n1209 0.110872
R6545 VGND.n798 VGND.n797 0.110872
R6546 VGND.n1229 VGND.n1228 0.110872
R6547 VGND.n1235 VGND.n1234 0.110872
R6548 VGND.n723 VGND.n722 0.110872
R6549 VGND.n782 VGND.n781 0.110872
R6550 VGND.n777 VGND.n776 0.110872
R6551 VGND.n772 VGND.n771 0.110872
R6552 VGND.n767 VGND.n766 0.110872
R6553 VGND.n762 VGND.n761 0.110872
R6554 VGND.n757 VGND.n756 0.110872
R6555 VGND.n752 VGND.n751 0.110872
R6556 VGND.n747 VGND.n746 0.110872
R6557 VGND.n742 VGND.n741 0.110872
R6558 VGND.n737 VGND.n736 0.110872
R6559 VGND.n732 VGND.n731 0.110872
R6560 VGND.n727 VGND.n726 0.110872
R6561 VGND.n688 VGND.n687 0.110872
R6562 VGND.n1291 VGND.n1290 0.110872
R6563 VGND.n1090 VGND 0.0981562
R6564 VGND.n998 VGND 0.0981562
R6565 VGND.n1059 VGND 0.0981562
R6566 VGND VGND.n147 0.0968542
R6567 VGND VGND.n615 0.0968542
R6568 VGND VGND.n991 0.0968542
R6569 VGND.n1028 VGND 0.0968542
R6570 VGND VGND.n177 0.0968542
R6571 VGND.n19 VGND 0.0968542
R6572 VGND VGND.n2903 0.0968542
R6573 VGND VGND.n64 0.0968542
R6574 VGND.n2932 VGND 0.0968542
R6575 VGND.n48 VGND 0.0968542
R6576 VGND.n2972 VGND 0.0968542
R6577 VGND.n2524 VGND 0.088625
R6578 VGND.n2714 VGND 0.0790114
R6579 VGND VGND.n2713 0.0790114
R6580 VGND VGND.n192 0.0790114
R6581 VGND.n2820 VGND 0.0790114
R6582 VGND VGND.n2819 0.0790114
R6583 VGND.n2814 VGND 0.0790114
R6584 VGND VGND.n2813 0.0790114
R6585 VGND.n2808 VGND 0.0790114
R6586 VGND VGND.n2807 0.0790114
R6587 VGND.n2802 VGND 0.0790114
R6588 VGND VGND.n2801 0.0790114
R6589 VGND.n2796 VGND 0.0790114
R6590 VGND VGND.n2795 0.0790114
R6591 VGND.n2790 VGND 0.0790114
R6592 VGND VGND.n2789 0.0790114
R6593 VGND.n3003 VGND 0.0790114
R6594 VGND.n2716 VGND 0.0790114
R6595 VGND.n2717 VGND 0.0790114
R6596 VGND.n2823 VGND 0.0790114
R6597 VGND VGND.n2822 0.0790114
R6598 VGND.n2817 VGND 0.0790114
R6599 VGND VGND.n2816 0.0790114
R6600 VGND.n2811 VGND 0.0790114
R6601 VGND VGND.n2810 0.0790114
R6602 VGND.n2805 VGND 0.0790114
R6603 VGND VGND.n2804 0.0790114
R6604 VGND.n2799 VGND 0.0790114
R6605 VGND VGND.n2798 0.0790114
R6606 VGND.n2793 VGND 0.0790114
R6607 VGND VGND.n2792 0.0790114
R6608 VGND.n2787 VGND 0.0790114
R6609 VGND.n3001 VGND 0.0790114
R6610 VGND VGND.n2521 0.0790114
R6611 VGND.n2827 VGND 0.0790114
R6612 VGND VGND.n2826 0.0790114
R6613 VGND.n2507 VGND 0.0790114
R6614 VGND VGND.n2506 0.0790114
R6615 VGND VGND.n2505 0.0790114
R6616 VGND VGND.n2504 0.0790114
R6617 VGND VGND.n2503 0.0790114
R6618 VGND VGND.n2502 0.0790114
R6619 VGND VGND.n2501 0.0790114
R6620 VGND VGND.n2500 0.0790114
R6621 VGND VGND.n2499 0.0790114
R6622 VGND VGND.n2498 0.0790114
R6623 VGND VGND.n2497 0.0790114
R6624 VGND VGND.n2496 0.0790114
R6625 VGND VGND.n2495 0.0790114
R6626 VGND.n643 VGND 0.0790114
R6627 VGND.n2830 VGND 0.0790114
R6628 VGND.n379 VGND 0.0790114
R6629 VGND.n2169 VGND 0.0790114
R6630 VGND.n2179 VGND 0.0790114
R6631 VGND.n2195 VGND 0.0790114
R6632 VGND.n2205 VGND 0.0790114
R6633 VGND.n2221 VGND 0.0790114
R6634 VGND.n2231 VGND 0.0790114
R6635 VGND.n2247 VGND 0.0790114
R6636 VGND.n2257 VGND 0.0790114
R6637 VGND.n2278 VGND 0.0790114
R6638 VGND.n2301 VGND 0.0790114
R6639 VGND VGND.n2300 0.0790114
R6640 VGND VGND.n2298 0.0790114
R6641 VGND.n2434 VGND 0.0790114
R6642 VGND.n1437 VGND 0.0790114
R6643 VGND VGND.n1436 0.0790114
R6644 VGND.n2156 VGND 0.0790114
R6645 VGND.n2166 VGND 0.0790114
R6646 VGND.n2182 VGND 0.0790114
R6647 VGND.n2192 VGND 0.0790114
R6648 VGND.n2208 VGND 0.0790114
R6649 VGND.n2218 VGND 0.0790114
R6650 VGND.n2234 VGND 0.0790114
R6651 VGND.n2244 VGND 0.0790114
R6652 VGND.n2260 VGND 0.0790114
R6653 VGND.n2275 VGND 0.0790114
R6654 VGND.n2304 VGND 0.0790114
R6655 VGND.n2305 VGND 0.0790114
R6656 VGND.n2318 VGND 0.0790114
R6657 VGND VGND.n2317 0.0790114
R6658 VGND.n1440 VGND 0.0790114
R6659 VGND.n1500 VGND 0.0790114
R6660 VGND.n2153 VGND 0.0790114
R6661 VGND VGND.n2152 0.0790114
R6662 VGND VGND.n2151 0.0790114
R6663 VGND VGND.n2150 0.0790114
R6664 VGND VGND.n2149 0.0790114
R6665 VGND VGND.n2148 0.0790114
R6666 VGND VGND.n2147 0.0790114
R6667 VGND VGND.n2146 0.0790114
R6668 VGND VGND.n2145 0.0790114
R6669 VGND VGND.n2144 0.0790114
R6670 VGND VGND.n2143 0.0790114
R6671 VGND.n2322 VGND 0.0790114
R6672 VGND VGND.n2321 0.0790114
R6673 VGND.n2129 VGND 0.0790114
R6674 VGND VGND.n1418 0.0790114
R6675 VGND.n1503 VGND 0.0790114
R6676 VGND VGND.n634 0.0790114
R6677 VGND.n1995 VGND 0.0790114
R6678 VGND.n2005 VGND 0.0790114
R6679 VGND.n2021 VGND 0.0790114
R6680 VGND.n2031 VGND 0.0790114
R6681 VGND.n2047 VGND 0.0790114
R6682 VGND.n2057 VGND 0.0790114
R6683 VGND.n2073 VGND 0.0790114
R6684 VGND.n2083 VGND 0.0790114
R6685 VGND.n2104 VGND 0.0790114
R6686 VGND.n2326 VGND 0.0790114
R6687 VGND VGND.n2325 0.0790114
R6688 VGND.n402 VGND 0.0790114
R6689 VGND.n2126 VGND 0.0790114
R6690 VGND VGND.n1416 0.0790114
R6691 VGND VGND.n660 0.0790114
R6692 VGND.n1982 VGND 0.0790114
R6693 VGND.n1992 VGND 0.0790114
R6694 VGND.n2008 VGND 0.0790114
R6695 VGND.n2018 VGND 0.0790114
R6696 VGND.n2034 VGND 0.0790114
R6697 VGND.n2044 VGND 0.0790114
R6698 VGND.n2060 VGND 0.0790114
R6699 VGND.n2070 VGND 0.0790114
R6700 VGND.n2086 VGND 0.0790114
R6701 VGND.n2101 VGND 0.0790114
R6702 VGND.n2329 VGND 0.0790114
R6703 VGND.n2330 VGND 0.0790114
R6704 VGND.n2343 VGND 0.0790114
R6705 VGND VGND.n2342 0.0790114
R6706 VGND.n1413 VGND 0.0790114
R6707 VGND VGND.n1412 0.0790114
R6708 VGND.n1979 VGND 0.0790114
R6709 VGND VGND.n1978 0.0790114
R6710 VGND VGND.n1977 0.0790114
R6711 VGND VGND.n1976 0.0790114
R6712 VGND VGND.n1975 0.0790114
R6713 VGND VGND.n1974 0.0790114
R6714 VGND VGND.n1973 0.0790114
R6715 VGND VGND.n1972 0.0790114
R6716 VGND VGND.n1971 0.0790114
R6717 VGND VGND.n1970 0.0790114
R6718 VGND VGND.n1969 0.0790114
R6719 VGND.n2347 VGND 0.0790114
R6720 VGND VGND.n2346 0.0790114
R6721 VGND.n1955 VGND 0.0790114
R6722 VGND.n1393 VGND 0.0790114
R6723 VGND.n1409 VGND 0.0790114
R6724 VGND VGND.n1408 0.0790114
R6725 VGND.n1821 VGND 0.0790114
R6726 VGND.n1831 VGND 0.0790114
R6727 VGND.n1847 VGND 0.0790114
R6728 VGND.n1857 VGND 0.0790114
R6729 VGND.n1873 VGND 0.0790114
R6730 VGND.n1883 VGND 0.0790114
R6731 VGND.n1899 VGND 0.0790114
R6732 VGND.n1909 VGND 0.0790114
R6733 VGND.n1930 VGND 0.0790114
R6734 VGND.n2351 VGND 0.0790114
R6735 VGND VGND.n2350 0.0790114
R6736 VGND.n458 VGND 0.0790114
R6737 VGND.n1952 VGND 0.0790114
R6738 VGND VGND.n1390 0.0790114
R6739 VGND VGND.n1388 0.0790114
R6740 VGND.n1808 VGND 0.0790114
R6741 VGND.n1818 VGND 0.0790114
R6742 VGND.n1834 VGND 0.0790114
R6743 VGND.n1844 VGND 0.0790114
R6744 VGND.n1860 VGND 0.0790114
R6745 VGND.n1870 VGND 0.0790114
R6746 VGND.n1886 VGND 0.0790114
R6747 VGND.n1896 VGND 0.0790114
R6748 VGND.n1912 VGND 0.0790114
R6749 VGND.n1927 VGND 0.0790114
R6750 VGND.n2354 VGND 0.0790114
R6751 VGND.n2355 VGND 0.0790114
R6752 VGND.n2368 VGND 0.0790114
R6753 VGND VGND.n2367 0.0790114
R6754 VGND VGND.n1372 0.0790114
R6755 VGND VGND.n1371 0.0790114
R6756 VGND.n1805 VGND 0.0790114
R6757 VGND VGND.n1804 0.0790114
R6758 VGND VGND.n1803 0.0790114
R6759 VGND VGND.n1802 0.0790114
R6760 VGND VGND.n1801 0.0790114
R6761 VGND VGND.n1800 0.0790114
R6762 VGND VGND.n1799 0.0790114
R6763 VGND VGND.n1798 0.0790114
R6764 VGND VGND.n1797 0.0790114
R6765 VGND VGND.n1796 0.0790114
R6766 VGND VGND.n1795 0.0790114
R6767 VGND.n2372 VGND 0.0790114
R6768 VGND VGND.n2371 0.0790114
R6769 VGND.n1781 VGND 0.0790114
R6770 VGND.n1532 VGND 0.0790114
R6771 VGND VGND.n1531 0.0790114
R6772 VGND VGND.n1530 0.0790114
R6773 VGND.n1647 VGND 0.0790114
R6774 VGND.n1657 VGND 0.0790114
R6775 VGND.n1673 VGND 0.0790114
R6776 VGND.n1683 VGND 0.0790114
R6777 VGND.n1699 VGND 0.0790114
R6778 VGND.n1709 VGND 0.0790114
R6779 VGND.n1725 VGND 0.0790114
R6780 VGND.n1735 VGND 0.0790114
R6781 VGND.n1756 VGND 0.0790114
R6782 VGND.n2376 VGND 0.0790114
R6783 VGND VGND.n2375 0.0790114
R6784 VGND.n514 VGND 0.0790114
R6785 VGND.n1778 VGND 0.0790114
R6786 VGND.n1535 VGND 0.0790114
R6787 VGND.n1545 VGND 0.0790114
R6788 VGND.n1634 VGND 0.0790114
R6789 VGND.n1644 VGND 0.0790114
R6790 VGND.n1660 VGND 0.0790114
R6791 VGND.n1670 VGND 0.0790114
R6792 VGND.n1686 VGND 0.0790114
R6793 VGND.n1696 VGND 0.0790114
R6794 VGND.n1712 VGND 0.0790114
R6795 VGND.n1722 VGND 0.0790114
R6796 VGND.n1738 VGND 0.0790114
R6797 VGND.n1753 VGND 0.0790114
R6798 VGND.n2379 VGND 0.0790114
R6799 VGND.n2380 VGND 0.0790114
R6800 VGND.n2393 VGND 0.0790114
R6801 VGND VGND.n2392 0.0790114
R6802 VGND VGND.n1302 0.0790114
R6803 VGND.n1548 VGND 0.0790114
R6804 VGND.n1631 VGND 0.0790114
R6805 VGND VGND.n1630 0.0790114
R6806 VGND VGND.n1629 0.0790114
R6807 VGND VGND.n1628 0.0790114
R6808 VGND VGND.n1627 0.0790114
R6809 VGND VGND.n1626 0.0790114
R6810 VGND VGND.n1625 0.0790114
R6811 VGND VGND.n1624 0.0790114
R6812 VGND VGND.n1623 0.0790114
R6813 VGND VGND.n1622 0.0790114
R6814 VGND VGND.n1621 0.0790114
R6815 VGND.n2397 VGND 0.0790114
R6816 VGND VGND.n2396 0.0790114
R6817 VGND.n1607 VGND 0.0790114
R6818 VGND.n900 VGND 0.0790114
R6819 VGND VGND.n899 0.0790114
R6820 VGND VGND.n898 0.0790114
R6821 VGND.n1279 VGND 0.0790114
R6822 VGND VGND.n1278 0.0790114
R6823 VGND.n1271 VGND 0.0790114
R6824 VGND VGND.n1270 0.0790114
R6825 VGND.n1263 VGND 0.0790114
R6826 VGND VGND.n1262 0.0790114
R6827 VGND.n1255 VGND 0.0790114
R6828 VGND VGND.n1254 0.0790114
R6829 VGND.n1247 VGND 0.0790114
R6830 VGND VGND.n1246 0.0790114
R6831 VGND.n2400 VGND 0.0790114
R6832 VGND.n288 VGND 0.0790114
R6833 VGND.n2412 VGND 0.0790114
R6834 VGND.n1123 VGND 0.0790114
R6835 VGND.n1286 VGND 0.0790114
R6836 VGND VGND.n1285 0.0790114
R6837 VGND.n691 VGND 0.0790114
R6838 VGND.n694 VGND 0.0790114
R6839 VGND.n697 VGND 0.0790114
R6840 VGND.n700 VGND 0.0790114
R6841 VGND.n703 VGND 0.0790114
R6842 VGND.n706 VGND 0.0790114
R6843 VGND.n709 VGND 0.0790114
R6844 VGND.n712 VGND 0.0790114
R6845 VGND.n715 VGND 0.0790114
R6846 VGND.n718 VGND 0.0790114
R6847 VGND.n1224 VGND 0.0790114
R6848 VGND.n1239 VGND 0.0790114
R6849 VGND VGND.n1238 0.0790114
R6850 VGND.n1121 VGND 0.0790114
R6851 VGND.n1288 VGND 0.0790114
R6852 VGND.n1283 VGND 0.0790114
R6853 VGND VGND.n1282 0.0790114
R6854 VGND.n1275 VGND 0.0790114
R6855 VGND VGND.n1274 0.0790114
R6856 VGND.n1267 VGND 0.0790114
R6857 VGND VGND.n1266 0.0790114
R6858 VGND.n1259 VGND 0.0790114
R6859 VGND VGND.n1258 0.0790114
R6860 VGND.n1251 VGND 0.0790114
R6861 VGND VGND.n1250 0.0790114
R6862 VGND.n1243 VGND 0.0790114
R6863 VGND VGND.n1242 0.0790114
R6864 VGND VGND.n1241 0.0790114
R6865 VGND.n2415 VGND 0.0790114
R6866 VGND.n2658 VGND.n2657 0.0656596
R6867 VGND.n2653 VGND.n2651 0.0656596
R6868 VGND.n2666 VGND.n2665 0.0656596
R6869 VGND.n2649 VGND.n2647 0.0656596
R6870 VGND.n2674 VGND.n2673 0.0656596
R6871 VGND.n2645 VGND.n2643 0.0656596
R6872 VGND.n2682 VGND.n2681 0.0656596
R6873 VGND.n2641 VGND.n2639 0.0656596
R6874 VGND.n2690 VGND.n2689 0.0656596
R6875 VGND.n2637 VGND.n2635 0.0656596
R6876 VGND.n2698 VGND.n2697 0.0656596
R6877 VGND.n2633 VGND.n2631 0.0656596
R6878 VGND.n2706 VGND.n2705 0.0656596
R6879 VGND.n2584 VGND.n2576 0.0656596
R6880 VGND.n2580 VGND.n2575 0.0656596
R6881 VGND.n2568 VGND 0.063
R6882 VGND.n2565 VGND 0.063
R6883 VGND.n2562 VGND 0.063
R6884 VGND.n2559 VGND 0.063
R6885 VGND.n2556 VGND 0.063
R6886 VGND.n2553 VGND 0.063
R6887 VGND.n2550 VGND 0.063
R6888 VGND.n2547 VGND 0.063
R6889 VGND.n2544 VGND 0.063
R6890 VGND.n2541 VGND 0.063
R6891 VGND.n2538 VGND 0.063
R6892 VGND.n2535 VGND 0.063
R6893 VGND.n2532 VGND 0.063
R6894 VGND.n2529 VGND 0.063
R6895 VGND.n2526 VGND 0.063
R6896 VGND.n1112 VGND 0.0603958
R6897 VGND.n1089 VGND 0.0603958
R6898 VGND VGND.n1088 0.0603958
R6899 VGND.n1085 VGND 0.0603958
R6900 VGND.n149 VGND 0.0603958
R6901 VGND VGND.n148 0.0603958
R6902 VGND.n131 VGND 0.0603958
R6903 VGND.n617 VGND 0.0603958
R6904 VGND VGND.n616 0.0603958
R6905 VGND.n599 VGND 0.0603958
R6906 VGND.n993 VGND 0.0603958
R6907 VGND VGND.n992 0.0603958
R6908 VGND.n985 VGND 0.0603958
R6909 VGND.n982 VGND 0.0603958
R6910 VGND.n977 VGND 0.0603958
R6911 VGND.n1027 VGND 0.0603958
R6912 VGND VGND.n1026 0.0603958
R6913 VGND.n1023 VGND 0.0603958
R6914 VGND.n1058 VGND 0.0603958
R6915 VGND VGND.n1057 0.0603958
R6916 VGND.n1054 VGND 0.0603958
R6917 VGND.n179 VGND 0.0603958
R6918 VGND VGND.n178 0.0603958
R6919 VGND.n161 VGND 0.0603958
R6920 VGND VGND.n31 0.0603958
R6921 VGND.n3006 VGND 0.0603958
R6922 VGND.n115 VGND 0.0603958
R6923 VGND VGND.n114 0.0603958
R6924 VGND.n2872 VGND 0.0603958
R6925 VGND VGND.n2871 0.0603958
R6926 VGND.n2905 VGND 0.0603958
R6927 VGND VGND.n2904 0.0603958
R6928 VGND.n2900 VGND 0.0603958
R6929 VGND.n2912 VGND 0.0603958
R6930 VGND.n2913 VGND 0.0603958
R6931 VGND VGND.n2944 0.0603958
R6932 VGND.n2945 VGND 0.0603958
R6933 VGND.n2946 VGND 0.0603958
R6934 VGND VGND.n60 0.0603958
R6935 VGND.n61 VGND 0.0603958
R6936 VGND.n2958 VGND 0.0603958
R6937 VGND VGND.n2984 0.0603958
R6938 VGND.n2985 VGND 0.0603958
R6939 VGND.n2990 VGND 0.0603958
R6940 VGND.n2657 VGND 0.0574853
R6941 VGND.n2653 VGND 0.0574853
R6942 VGND.n2665 VGND 0.0574853
R6943 VGND.n2649 VGND 0.0574853
R6944 VGND.n2673 VGND 0.0574853
R6945 VGND.n2645 VGND 0.0574853
R6946 VGND.n2681 VGND 0.0574853
R6947 VGND.n2641 VGND 0.0574853
R6948 VGND.n2689 VGND 0.0574853
R6949 VGND.n2637 VGND 0.0574853
R6950 VGND.n2697 VGND 0.0574853
R6951 VGND.n2633 VGND 0.0574853
R6952 VGND.n2705 VGND 0.0574853
R6953 VGND.n2584 VGND 0.0574853
R6954 VGND.n2575 VGND 0.0574853
R6955 VGND.n826 VGND 0.0489375
R6956 VGND.n789 VGND 0.0489375
R6957 VGND.n2589 VGND 0.0489375
R6958 VGND.n2586 VGND 0.0489375
R6959 VGND.n2572 VGND 0.0489375
R6960 VGND.n2585 VGND 0.0489375
R6961 VGND.n2624 VGND 0.0489375
R6962 VGND.n2621 VGND 0.0489375
R6963 VGND.n2618 VGND 0.0489375
R6964 VGND.n2615 VGND 0.0489375
R6965 VGND.n2612 VGND 0.0489375
R6966 VGND.n2609 VGND 0.0489375
R6967 VGND.n2606 VGND 0.0489375
R6968 VGND.n2603 VGND 0.0489375
R6969 VGND.n2600 VGND 0.0489375
R6970 VGND.n2597 VGND 0.0489375
R6971 VGND.n2594 VGND 0.0489375
R6972 VGND.n2591 VGND 0.0489375
R6973 VGND.n823 VGND 0.0489375
R6974 VGND.n820 VGND 0.0489375
R6975 VGND.n1140 VGND 0.0489375
R6976 VGND.n811 VGND 0.0489375
R6977 VGND.n809 VGND 0.0489375
R6978 VGND.n1155 VGND 0.0489375
R6979 VGND.n1172 VGND 0.0489375
R6980 VGND.n803 VGND 0.0489375
R6981 VGND.n801 VGND 0.0489375
R6982 VGND.n1187 VGND 0.0489375
R6983 VGND.n1204 VGND 0.0489375
R6984 VGND.n795 VGND 0.0489375
R6985 VGND.n793 VGND 0.0489375
R6986 VGND.n1219 VGND 0.0489375
R6987 VGND.n2 VGND 0.0445
R6988 VGND.n3032 VGND.n2 0.043
R6989 VGND VGND.n2578 0.037734
R6990 VGND.n230 VGND 0.037734
R6991 VGND.n2780 VGND 0.037734
R6992 VGND.n2775 VGND 0.037734
R6993 VGND.n2770 VGND 0.037734
R6994 VGND.n2765 VGND 0.037734
R6995 VGND.n2760 VGND 0.037734
R6996 VGND.n2755 VGND 0.037734
R6997 VGND.n2750 VGND 0.037734
R6998 VGND.n2745 VGND 0.037734
R6999 VGND.n2740 VGND 0.037734
R7000 VGND.n2735 VGND 0.037734
R7001 VGND.n2730 VGND 0.037734
R7002 VGND.n2725 VGND 0.037734
R7003 VGND.n2720 VGND 0.037734
R7004 VGND.n235 VGND 0.037734
R7005 VGND VGND.n233 0.037734
R7006 VGND.n2489 VGND 0.037734
R7007 VGND.n2484 VGND 0.037734
R7008 VGND.n2479 VGND 0.037734
R7009 VGND.n2474 VGND 0.037734
R7010 VGND.n2469 VGND 0.037734
R7011 VGND.n2464 VGND 0.037734
R7012 VGND.n2459 VGND 0.037734
R7013 VGND.n2454 VGND 0.037734
R7014 VGND.n2449 VGND 0.037734
R7015 VGND.n2444 VGND 0.037734
R7016 VGND.n2439 VGND 0.037734
R7017 VGND VGND.n251 0.037734
R7018 VGND.n2509 VGND 0.037734
R7019 VGND.n2514 VGND 0.037734
R7020 VGND.n245 VGND 0.037734
R7021 VGND VGND.n243 0.037734
R7022 VGND.n335 VGND 0.037734
R7023 VGND.n2291 VGND 0.037734
R7024 VGND.n2286 VGND 0.037734
R7025 VGND.n2281 VGND 0.037734
R7026 VGND.n343 VGND 0.037734
R7027 VGND.n2250 VGND 0.037734
R7028 VGND.n351 VGND 0.037734
R7029 VGND.n2224 VGND 0.037734
R7030 VGND.n359 VGND 0.037734
R7031 VGND.n2198 VGND 0.037734
R7032 VGND.n367 VGND 0.037734
R7033 VGND.n2172 VGND 0.037734
R7034 VGND.n373 VGND 0.037734
R7035 VGND VGND.n371 0.037734
R7036 VGND.n2832 VGND 0.037734
R7037 VGND VGND.n183 0.037734
R7038 VGND VGND.n2315 0.037734
R7039 VGND.n2308 VGND 0.037734
R7040 VGND.n2268 VGND 0.037734
R7041 VGND.n339 VGND 0.037734
R7042 VGND.n2263 VGND 0.037734
R7043 VGND.n347 VGND 0.037734
R7044 VGND.n2237 VGND 0.037734
R7045 VGND.n355 VGND 0.037734
R7046 VGND.n2211 VGND 0.037734
R7047 VGND.n363 VGND 0.037734
R7048 VGND.n2185 VGND 0.037734
R7049 VGND.n382 VGND 0.037734
R7050 VGND.n2159 VGND 0.037734
R7051 VGND.n1426 VGND 0.037734
R7052 VGND.n1429 VGND 0.037734
R7053 VGND VGND.n1423 0.037734
R7054 VGND.n2131 VGND 0.037734
R7055 VGND.n2136 VGND 0.037734
R7056 VGND.n396 VGND 0.037734
R7057 VGND.n1448 VGND 0.037734
R7058 VGND.n1453 VGND 0.037734
R7059 VGND.n1458 VGND 0.037734
R7060 VGND.n1463 VGND 0.037734
R7061 VGND.n1468 VGND 0.037734
R7062 VGND.n1473 VGND 0.037734
R7063 VGND.n1478 VGND 0.037734
R7064 VGND.n1483 VGND 0.037734
R7065 VGND.n1488 VGND 0.037734
R7066 VGND.n1493 VGND 0.037734
R7067 VGND.n637 VGND 0.037734
R7068 VGND.n1443 VGND 0.037734
R7069 VGND VGND.n641 0.037734
R7070 VGND VGND.n2124 0.037734
R7071 VGND.n2117 VGND 0.037734
R7072 VGND.n2112 VGND 0.037734
R7073 VGND.n2107 VGND 0.037734
R7074 VGND.n410 VGND 0.037734
R7075 VGND.n2076 VGND 0.037734
R7076 VGND.n418 VGND 0.037734
R7077 VGND.n2050 VGND 0.037734
R7078 VGND.n426 VGND 0.037734
R7079 VGND.n2024 VGND 0.037734
R7080 VGND.n434 VGND 0.037734
R7081 VGND.n1998 VGND 0.037734
R7082 VGND.n628 VGND 0.037734
R7083 VGND VGND.n626 0.037734
R7084 VGND.n1505 VGND 0.037734
R7085 VGND VGND.n620 0.037734
R7086 VGND VGND.n2340 0.037734
R7087 VGND.n2333 VGND 0.037734
R7088 VGND.n2094 VGND 0.037734
R7089 VGND.n406 VGND 0.037734
R7090 VGND.n2089 VGND 0.037734
R7091 VGND.n414 VGND 0.037734
R7092 VGND.n2063 VGND 0.037734
R7093 VGND.n422 VGND 0.037734
R7094 VGND.n2037 VGND 0.037734
R7095 VGND.n430 VGND 0.037734
R7096 VGND.n2011 VGND 0.037734
R7097 VGND.n438 VGND 0.037734
R7098 VGND.n1985 VGND 0.037734
R7099 VGND.n650 VGND 0.037734
R7100 VGND.n653 VGND 0.037734
R7101 VGND VGND.n647 0.037734
R7102 VGND.n1957 VGND 0.037734
R7103 VGND.n1962 VGND 0.037734
R7104 VGND.n452 VGND 0.037734
R7105 VGND.n905 VGND 0.037734
R7106 VGND.n910 VGND 0.037734
R7107 VGND.n915 VGND 0.037734
R7108 VGND.n920 VGND 0.037734
R7109 VGND.n925 VGND 0.037734
R7110 VGND.n930 VGND 0.037734
R7111 VGND.n935 VGND 0.037734
R7112 VGND.n940 VGND 0.037734
R7113 VGND.n945 VGND 0.037734
R7114 VGND.n950 VGND 0.037734
R7115 VGND.n955 VGND 0.037734
R7116 VGND.n960 VGND 0.037734
R7117 VGND VGND.n663 0.037734
R7118 VGND VGND.n1950 0.037734
R7119 VGND.n1943 VGND 0.037734
R7120 VGND.n1938 VGND 0.037734
R7121 VGND.n1933 VGND 0.037734
R7122 VGND.n466 VGND 0.037734
R7123 VGND.n1902 VGND 0.037734
R7124 VGND.n474 VGND 0.037734
R7125 VGND.n1876 VGND 0.037734
R7126 VGND.n482 VGND 0.037734
R7127 VGND.n1850 VGND 0.037734
R7128 VGND.n490 VGND 0.037734
R7129 VGND.n1824 VGND 0.037734
R7130 VGND.n669 VGND 0.037734
R7131 VGND.n1401 VGND 0.037734
R7132 VGND.n1396 VGND 0.037734
R7133 VGND VGND.n672 0.037734
R7134 VGND VGND.n2365 0.037734
R7135 VGND.n2358 VGND 0.037734
R7136 VGND.n1920 VGND 0.037734
R7137 VGND.n462 VGND 0.037734
R7138 VGND.n1915 VGND 0.037734
R7139 VGND.n470 VGND 0.037734
R7140 VGND.n1889 VGND 0.037734
R7141 VGND.n478 VGND 0.037734
R7142 VGND.n1863 VGND 0.037734
R7143 VGND.n486 VGND 0.037734
R7144 VGND.n1837 VGND 0.037734
R7145 VGND.n494 VGND 0.037734
R7146 VGND.n1811 VGND 0.037734
R7147 VGND.n1378 VGND 0.037734
R7148 VGND.n1381 VGND 0.037734
R7149 VGND VGND.n1375 0.037734
R7150 VGND.n1783 VGND 0.037734
R7151 VGND.n1788 VGND 0.037734
R7152 VGND.n508 VGND 0.037734
R7153 VGND.n1318 VGND 0.037734
R7154 VGND.n1323 VGND 0.037734
R7155 VGND.n1328 VGND 0.037734
R7156 VGND.n1333 VGND 0.037734
R7157 VGND.n1338 VGND 0.037734
R7158 VGND.n1343 VGND 0.037734
R7159 VGND.n1348 VGND 0.037734
R7160 VGND.n1353 VGND 0.037734
R7161 VGND.n1358 VGND 0.037734
R7162 VGND.n1363 VGND 0.037734
R7163 VGND.n1310 VGND 0.037734
R7164 VGND.n1313 VGND 0.037734
R7165 VGND VGND.n1307 0.037734
R7166 VGND VGND.n1776 0.037734
R7167 VGND.n1769 VGND 0.037734
R7168 VGND.n1764 VGND 0.037734
R7169 VGND.n1759 VGND 0.037734
R7170 VGND.n522 VGND 0.037734
R7171 VGND.n1728 VGND 0.037734
R7172 VGND.n530 VGND 0.037734
R7173 VGND.n1702 VGND 0.037734
R7174 VGND.n538 VGND 0.037734
R7175 VGND.n1676 VGND 0.037734
R7176 VGND.n546 VGND 0.037734
R7177 VGND.n1650 VGND 0.037734
R7178 VGND.n580 VGND 0.037734
R7179 VGND.n1523 VGND 0.037734
R7180 VGND.n1518 VGND 0.037734
R7181 VGND VGND.n576 0.037734
R7182 VGND VGND.n2390 0.037734
R7183 VGND.n2383 VGND 0.037734
R7184 VGND.n1746 VGND 0.037734
R7185 VGND.n518 VGND 0.037734
R7186 VGND.n1741 VGND 0.037734
R7187 VGND.n526 VGND 0.037734
R7188 VGND.n1715 VGND 0.037734
R7189 VGND.n534 VGND 0.037734
R7190 VGND.n1689 VGND 0.037734
R7191 VGND.n542 VGND 0.037734
R7192 VGND.n1663 VGND 0.037734
R7193 VGND.n550 VGND 0.037734
R7194 VGND.n1637 VGND 0.037734
R7195 VGND.n569 VGND 0.037734
R7196 VGND.n1538 VGND 0.037734
R7197 VGND VGND.n572 0.037734
R7198 VGND.n1609 VGND 0.037734
R7199 VGND.n1614 VGND 0.037734
R7200 VGND.n564 VGND 0.037734
R7201 VGND.n1601 VGND 0.037734
R7202 VGND.n1596 VGND 0.037734
R7203 VGND.n1591 VGND 0.037734
R7204 VGND.n1586 VGND 0.037734
R7205 VGND.n1581 VGND 0.037734
R7206 VGND.n1576 VGND 0.037734
R7207 VGND.n1571 VGND 0.037734
R7208 VGND.n1566 VGND 0.037734
R7209 VGND.n1561 VGND 0.037734
R7210 VGND.n1556 VGND 0.037734
R7211 VGND.n1551 VGND 0.037734
R7212 VGND.n677 VGND 0.037734
R7213 VGND VGND.n675 0.037734
R7214 VGND VGND.n2410 0.037734
R7215 VGND.n2403 VGND 0.037734
R7216 VGND.n846 VGND 0.037734
R7217 VGND.n851 VGND 0.037734
R7218 VGND.n856 VGND 0.037734
R7219 VGND.n861 VGND 0.037734
R7220 VGND.n866 VGND 0.037734
R7221 VGND.n871 VGND 0.037734
R7222 VGND.n876 VGND 0.037734
R7223 VGND.n881 VGND 0.037734
R7224 VGND.n886 VGND 0.037734
R7225 VGND.n891 VGND 0.037734
R7226 VGND.n833 VGND 0.037734
R7227 VGND.n841 VGND 0.037734
R7228 VGND.n836 VGND 0.037734
R7229 VGND VGND.n829 0.037734
R7230 VGND VGND.n819 0.037734
R7231 VGND VGND.n1129 0.037734
R7232 VGND.n1132 VGND 0.037734
R7233 VGND VGND.n1139 0.037734
R7234 VGND.n1145 VGND 0.037734
R7235 VGND.n813 VGND 0.037734
R7236 VGND.n1164 VGND 0.037734
R7237 VGND VGND.n1171 0.037734
R7238 VGND.n1177 VGND 0.037734
R7239 VGND.n805 VGND 0.037734
R7240 VGND.n1196 VGND 0.037734
R7241 VGND VGND.n1203 0.037734
R7242 VGND.n1209 VGND 0.037734
R7243 VGND.n797 VGND 0.037734
R7244 VGND.n1228 VGND 0.037734
R7245 VGND VGND.n1235 0.037734
R7246 VGND.n722 VGND 0.037734
R7247 VGND.n781 VGND 0.037734
R7248 VGND.n776 VGND 0.037734
R7249 VGND.n771 VGND 0.037734
R7250 VGND.n766 VGND 0.037734
R7251 VGND.n761 VGND 0.037734
R7252 VGND.n756 VGND 0.037734
R7253 VGND.n751 VGND 0.037734
R7254 VGND.n746 VGND 0.037734
R7255 VGND.n741 VGND 0.037734
R7256 VGND.n736 VGND 0.037734
R7257 VGND.n731 VGND 0.037734
R7258 VGND.n726 VGND 0.037734
R7259 VGND VGND.n688 0.037734
R7260 VGND.n1290 VGND 0.037734
R7261 VGND VGND.n680 0.037734
R7262 VGND.n1116 VGND 0.0343542
R7263 VGND.n1088 VGND 0.0343542
R7264 VGND.n149 VGND 0.0343542
R7265 VGND.n617 VGND 0.0343542
R7266 VGND.n993 VGND 0.0343542
R7267 VGND.n1026 VGND 0.0343542
R7268 VGND.n1057 VGND 0.0343542
R7269 VGND.n179 VGND 0.0343542
R7270 VGND.n3006 VGND 0.0330521
R7271 VGND.n115 VGND 0.0330521
R7272 VGND.n2872 VGND 0.0330521
R7273 VGND.n2905 VGND 0.0330521
R7274 VGND VGND.n2912 0.0330521
R7275 VGND VGND.n2945 0.0330521
R7276 VGND VGND.n61 0.0330521
R7277 VGND VGND.n2985 0.0330521
R7278 VGND.n3005 VGND 0.024
R7279 VGND.n1 VGND 0.024
R7280 VGND.n148 VGND 0.0239375
R7281 VGND.n616 VGND 0.0239375
R7282 VGND.n178 VGND 0.0239375
R7283 VGND.n2904 VGND 0.0239375
R7284 VGND.n2913 VGND 0.0239375
R7285 VGND.n1093 VGND 0.0226354
R7286 VGND VGND.n123 0.0226354
R7287 VGND.n1001 VGND 0.0226354
R7288 VGND.n992 VGND 0.0226354
R7289 VGND.n1032 VGND 0.0226354
R7290 VGND VGND.n2918 0.0226354
R7291 VGND.n2956 VGND 0.0226354
R7292 VGND.n2988 VGND 0.0226354
R7293 VGND VGND.n591 0.0213333
R7294 VGND.n997 VGND 0.0213333
R7295 VGND.n1063 VGND 0.0213333
R7296 VGND VGND.n112 0.0213333
R7297 VGND.n114 VGND 0.0213333
R7298 VGND VGND.n2867 0.0213333
R7299 VGND.n2871 VGND 0.0213333
R7300 VGND VGND.n2899 0.0213333
R7301 VGND.n86 VGND 0.0213333
R7302 VGND VGND.n2951 0.0213333
R7303 VGND.n3005 VGND 0.0161667
R7304 VGND.n3021 VGND 0.0144286
R7305 VGND.n2579 VGND 0.00980851
R7306 VGND.n3000 VGND 0.00980851
R7307 VGND.n2786 VGND 0.00980851
R7308 VGND VGND.n224 0.00980851
R7309 VGND VGND.n223 0.00980851
R7310 VGND VGND.n218 0.00980851
R7311 VGND VGND.n217 0.00980851
R7312 VGND VGND.n212 0.00980851
R7313 VGND VGND.n211 0.00980851
R7314 VGND VGND.n206 0.00980851
R7315 VGND VGND.n205 0.00980851
R7316 VGND VGND.n200 0.00980851
R7317 VGND VGND.n199 0.00980851
R7318 VGND VGND.n194 0.00980851
R7319 VGND VGND.n193 0.00980851
R7320 VGND.n2718 VGND 0.00980851
R7321 VGND.n239 VGND 0.00980851
R7322 VGND.n2494 VGND 0.00980851
R7323 VGND VGND.n262 0.00980851
R7324 VGND VGND.n261 0.00980851
R7325 VGND VGND.n260 0.00980851
R7326 VGND VGND.n259 0.00980851
R7327 VGND VGND.n258 0.00980851
R7328 VGND VGND.n257 0.00980851
R7329 VGND VGND.n256 0.00980851
R7330 VGND VGND.n255 0.00980851
R7331 VGND VGND.n254 0.00980851
R7332 VGND VGND.n253 0.00980851
R7333 VGND.n252 VGND 0.00980851
R7334 VGND VGND.n2508 0.00980851
R7335 VGND VGND.n190 0.00980851
R7336 VGND VGND.n189 0.00980851
R7337 VGND.n2520 VGND 0.00980851
R7338 VGND.n2433 VGND 0.00980851
R7339 VGND.n2297 VGND 0.00980851
R7340 VGND VGND.n333 0.00980851
R7341 VGND VGND.n332 0.00980851
R7342 VGND.n2279 VGND 0.00980851
R7343 VGND.n2256 VGND 0.00980851
R7344 VGND.n2248 VGND 0.00980851
R7345 VGND.n2230 VGND 0.00980851
R7346 VGND.n2222 VGND 0.00980851
R7347 VGND.n2204 VGND 0.00980851
R7348 VGND.n2196 VGND 0.00980851
R7349 VGND.n2178 VGND 0.00980851
R7350 VGND.n2170 VGND 0.00980851
R7351 VGND.n378 VGND 0.00980851
R7352 VGND VGND.n2831 0.00980851
R7353 VGND.n184 VGND 0.00980851
R7354 VGND.n2316 VGND 0.00980851
R7355 VGND VGND.n328 0.00980851
R7356 VGND.n2306 VGND 0.00980851
R7357 VGND VGND.n331 0.00980851
R7358 VGND.n2274 VGND 0.00980851
R7359 VGND.n2261 VGND 0.00980851
R7360 VGND.n2243 VGND 0.00980851
R7361 VGND.n2235 VGND 0.00980851
R7362 VGND.n2217 VGND 0.00980851
R7363 VGND.n2209 VGND 0.00980851
R7364 VGND.n2191 VGND 0.00980851
R7365 VGND.n2183 VGND 0.00980851
R7366 VGND.n2165 VGND 0.00980851
R7367 VGND.n2157 VGND 0.00980851
R7368 VGND.n1435 VGND 0.00980851
R7369 VGND.n1424 VGND 0.00980851
R7370 VGND VGND.n2130 0.00980851
R7371 VGND VGND.n326 0.00980851
R7372 VGND VGND.n325 0.00980851
R7373 VGND.n2142 VGND 0.00980851
R7374 VGND VGND.n394 0.00980851
R7375 VGND VGND.n393 0.00980851
R7376 VGND VGND.n392 0.00980851
R7377 VGND VGND.n391 0.00980851
R7378 VGND VGND.n390 0.00980851
R7379 VGND VGND.n389 0.00980851
R7380 VGND VGND.n388 0.00980851
R7381 VGND VGND.n387 0.00980851
R7382 VGND VGND.n386 0.00980851
R7383 VGND VGND.n385 0.00980851
R7384 VGND.n1499 VGND 0.00980851
R7385 VGND.n1441 VGND 0.00980851
R7386 VGND.n2125 VGND 0.00980851
R7387 VGND VGND.n403 0.00980851
R7388 VGND VGND.n323 0.00980851
R7389 VGND VGND.n322 0.00980851
R7390 VGND.n2105 VGND 0.00980851
R7391 VGND.n2082 VGND 0.00980851
R7392 VGND.n2074 VGND 0.00980851
R7393 VGND.n2056 VGND 0.00980851
R7394 VGND.n2048 VGND 0.00980851
R7395 VGND.n2030 VGND 0.00980851
R7396 VGND.n2022 VGND 0.00980851
R7397 VGND.n2004 VGND 0.00980851
R7398 VGND.n1996 VGND 0.00980851
R7399 VGND.n633 VGND 0.00980851
R7400 VGND VGND.n1504 0.00980851
R7401 VGND.n621 VGND 0.00980851
R7402 VGND.n2341 VGND 0.00980851
R7403 VGND VGND.n316 0.00980851
R7404 VGND.n2331 VGND 0.00980851
R7405 VGND VGND.n320 0.00980851
R7406 VGND.n2100 VGND 0.00980851
R7407 VGND.n2087 VGND 0.00980851
R7408 VGND.n2069 VGND 0.00980851
R7409 VGND.n2061 VGND 0.00980851
R7410 VGND.n2043 VGND 0.00980851
R7411 VGND.n2035 VGND 0.00980851
R7412 VGND.n2017 VGND 0.00980851
R7413 VGND.n2009 VGND 0.00980851
R7414 VGND.n1991 VGND 0.00980851
R7415 VGND.n1983 VGND 0.00980851
R7416 VGND.n659 VGND 0.00980851
R7417 VGND.n648 VGND 0.00980851
R7418 VGND VGND.n1956 0.00980851
R7419 VGND VGND.n314 0.00980851
R7420 VGND VGND.n313 0.00980851
R7421 VGND.n1968 VGND 0.00980851
R7422 VGND VGND.n450 0.00980851
R7423 VGND VGND.n449 0.00980851
R7424 VGND VGND.n448 0.00980851
R7425 VGND VGND.n447 0.00980851
R7426 VGND VGND.n446 0.00980851
R7427 VGND VGND.n445 0.00980851
R7428 VGND VGND.n444 0.00980851
R7429 VGND VGND.n443 0.00980851
R7430 VGND VGND.n442 0.00980851
R7431 VGND VGND.n441 0.00980851
R7432 VGND VGND.n665 0.00980851
R7433 VGND.n664 VGND 0.00980851
R7434 VGND.n1951 VGND 0.00980851
R7435 VGND VGND.n459 0.00980851
R7436 VGND VGND.n311 0.00980851
R7437 VGND VGND.n310 0.00980851
R7438 VGND.n1931 VGND 0.00980851
R7439 VGND.n1908 VGND 0.00980851
R7440 VGND.n1900 VGND 0.00980851
R7441 VGND.n1882 VGND 0.00980851
R7442 VGND.n1874 VGND 0.00980851
R7443 VGND.n1856 VGND 0.00980851
R7444 VGND.n1848 VGND 0.00980851
R7445 VGND.n1830 VGND 0.00980851
R7446 VGND.n1822 VGND 0.00980851
R7447 VGND.n1407 VGND 0.00980851
R7448 VGND VGND.n667 0.00980851
R7449 VGND.n1394 VGND 0.00980851
R7450 VGND.n2366 VGND 0.00980851
R7451 VGND VGND.n304 0.00980851
R7452 VGND.n2356 VGND 0.00980851
R7453 VGND VGND.n308 0.00980851
R7454 VGND.n1926 VGND 0.00980851
R7455 VGND.n1913 VGND 0.00980851
R7456 VGND.n1895 VGND 0.00980851
R7457 VGND.n1887 VGND 0.00980851
R7458 VGND.n1869 VGND 0.00980851
R7459 VGND.n1861 VGND 0.00980851
R7460 VGND.n1843 VGND 0.00980851
R7461 VGND.n1835 VGND 0.00980851
R7462 VGND.n1817 VGND 0.00980851
R7463 VGND.n1809 VGND 0.00980851
R7464 VGND.n1387 VGND 0.00980851
R7465 VGND.n1376 VGND 0.00980851
R7466 VGND VGND.n1782 0.00980851
R7467 VGND VGND.n302 0.00980851
R7468 VGND VGND.n301 0.00980851
R7469 VGND.n1794 VGND 0.00980851
R7470 VGND VGND.n506 0.00980851
R7471 VGND VGND.n505 0.00980851
R7472 VGND VGND.n504 0.00980851
R7473 VGND VGND.n503 0.00980851
R7474 VGND VGND.n502 0.00980851
R7475 VGND VGND.n501 0.00980851
R7476 VGND VGND.n500 0.00980851
R7477 VGND VGND.n499 0.00980851
R7478 VGND VGND.n498 0.00980851
R7479 VGND VGND.n497 0.00980851
R7480 VGND.n1369 VGND 0.00980851
R7481 VGND.n1308 VGND 0.00980851
R7482 VGND.n1777 VGND 0.00980851
R7483 VGND VGND.n515 0.00980851
R7484 VGND VGND.n299 0.00980851
R7485 VGND VGND.n298 0.00980851
R7486 VGND.n1757 VGND 0.00980851
R7487 VGND.n1734 VGND 0.00980851
R7488 VGND.n1726 VGND 0.00980851
R7489 VGND.n1708 VGND 0.00980851
R7490 VGND.n1700 VGND 0.00980851
R7491 VGND.n1682 VGND 0.00980851
R7492 VGND.n1674 VGND 0.00980851
R7493 VGND.n1656 VGND 0.00980851
R7494 VGND.n1648 VGND 0.00980851
R7495 VGND.n1529 VGND 0.00980851
R7496 VGND VGND.n578 0.00980851
R7497 VGND.n577 VGND 0.00980851
R7498 VGND.n2391 VGND 0.00980851
R7499 VGND VGND.n291 0.00980851
R7500 VGND.n2381 VGND 0.00980851
R7501 VGND VGND.n295 0.00980851
R7502 VGND.n1752 VGND 0.00980851
R7503 VGND.n1739 VGND 0.00980851
R7504 VGND.n1721 VGND 0.00980851
R7505 VGND.n1713 VGND 0.00980851
R7506 VGND.n1695 VGND 0.00980851
R7507 VGND.n1687 VGND 0.00980851
R7508 VGND.n1669 VGND 0.00980851
R7509 VGND.n1661 VGND 0.00980851
R7510 VGND.n1643 VGND 0.00980851
R7511 VGND.n1635 VGND 0.00980851
R7512 VGND.n1544 VGND 0.00980851
R7513 VGND.n1536 VGND 0.00980851
R7514 VGND VGND.n1608 0.00980851
R7515 VGND VGND.n287 0.00980851
R7516 VGND VGND.n286 0.00980851
R7517 VGND.n1620 VGND 0.00980851
R7518 VGND VGND.n562 0.00980851
R7519 VGND VGND.n561 0.00980851
R7520 VGND VGND.n560 0.00980851
R7521 VGND VGND.n559 0.00980851
R7522 VGND VGND.n558 0.00980851
R7523 VGND VGND.n557 0.00980851
R7524 VGND VGND.n556 0.00980851
R7525 VGND VGND.n555 0.00980851
R7526 VGND VGND.n554 0.00980851
R7527 VGND VGND.n553 0.00980851
R7528 VGND.n1549 VGND 0.00980851
R7529 VGND.n1301 VGND 0.00980851
R7530 VGND.n2411 VGND 0.00980851
R7531 VGND VGND.n283 0.00980851
R7532 VGND.n2401 VGND 0.00980851
R7533 VGND VGND.n717 0.00980851
R7534 VGND VGND.n716 0.00980851
R7535 VGND VGND.n711 0.00980851
R7536 VGND VGND.n710 0.00980851
R7537 VGND VGND.n705 0.00980851
R7538 VGND VGND.n704 0.00980851
R7539 VGND VGND.n699 0.00980851
R7540 VGND VGND.n698 0.00980851
R7541 VGND VGND.n693 0.00980851
R7542 VGND VGND.n692 0.00980851
R7543 VGND.n897 VGND 0.00980851
R7544 VGND VGND.n831 0.00980851
R7545 VGND.n830 VGND 0.00980851
R7546 VGND.n1125 VGND 0.00980851
R7547 VGND.n1130 VGND 0.00980851
R7548 VGND VGND.n816 0.00980851
R7549 VGND.n1143 VGND 0.00980851
R7550 VGND.n1151 VGND 0.00980851
R7551 VGND.n1162 VGND 0.00980851
R7552 VGND VGND.n808 0.00980851
R7553 VGND.n1175 VGND 0.00980851
R7554 VGND.n1183 VGND 0.00980851
R7555 VGND.n1194 VGND 0.00980851
R7556 VGND VGND.n800 0.00980851
R7557 VGND.n1207 VGND 0.00980851
R7558 VGND.n1215 VGND 0.00980851
R7559 VGND.n1226 VGND 0.00980851
R7560 VGND VGND.n792 0.00980851
R7561 VGND.n1236 VGND 0.00980851
R7562 VGND.n2416 VGND 0.00980851
R7563 VGND.n787 VGND 0.00980851
R7564 VGND VGND.n720 0.00980851
R7565 VGND VGND.n719 0.00980851
R7566 VGND VGND.n714 0.00980851
R7567 VGND VGND.n713 0.00980851
R7568 VGND VGND.n708 0.00980851
R7569 VGND VGND.n707 0.00980851
R7570 VGND VGND.n702 0.00980851
R7571 VGND VGND.n701 0.00980851
R7572 VGND VGND.n696 0.00980851
R7573 VGND VGND.n695 0.00980851
R7574 VGND VGND.n690 0.00980851
R7575 VGND.n689 VGND 0.00980851
R7576 VGND VGND.n1289 0.00980851
R7577 VGND.n681 VGND 0.00980851
R7578 VGND.n3033 VGND 0.00835714
R7579 VGND.n2657 VGND.n2655 0.00182979
R7580 VGND.n2654 VGND.n2653 0.00182979
R7581 VGND.n2665 VGND.n2663 0.00182979
R7582 VGND.n2650 VGND.n2649 0.00182979
R7583 VGND.n2673 VGND.n2671 0.00182979
R7584 VGND.n2646 VGND.n2645 0.00182979
R7585 VGND.n2681 VGND.n2679 0.00182979
R7586 VGND.n2642 VGND.n2641 0.00182979
R7587 VGND.n2689 VGND.n2687 0.00182979
R7588 VGND.n2638 VGND.n2637 0.00182979
R7589 VGND.n2697 VGND.n2695 0.00182979
R7590 VGND.n2634 VGND.n2633 0.00182979
R7591 VGND.n2705 VGND.n2703 0.00182979
R7592 VGND.n2630 VGND.n2584 0.00182979
R7593 VGND.n2711 VGND.n2575 0.00182979
R7594 XThR.Tn[2].n2 XThR.Tn[2].n1 332.332
R7595 XThR.Tn[2].n2 XThR.Tn[2].n0 296.493
R7596 XThR.Tn[2] XThR.Tn[2].n82 161.363
R7597 XThR.Tn[2] XThR.Tn[2].n77 161.363
R7598 XThR.Tn[2] XThR.Tn[2].n72 161.363
R7599 XThR.Tn[2] XThR.Tn[2].n67 161.363
R7600 XThR.Tn[2] XThR.Tn[2].n62 161.363
R7601 XThR.Tn[2] XThR.Tn[2].n57 161.363
R7602 XThR.Tn[2] XThR.Tn[2].n52 161.363
R7603 XThR.Tn[2] XThR.Tn[2].n47 161.363
R7604 XThR.Tn[2] XThR.Tn[2].n42 161.363
R7605 XThR.Tn[2] XThR.Tn[2].n37 161.363
R7606 XThR.Tn[2] XThR.Tn[2].n32 161.363
R7607 XThR.Tn[2] XThR.Tn[2].n27 161.363
R7608 XThR.Tn[2] XThR.Tn[2].n22 161.363
R7609 XThR.Tn[2] XThR.Tn[2].n17 161.363
R7610 XThR.Tn[2] XThR.Tn[2].n12 161.363
R7611 XThR.Tn[2] XThR.Tn[2].n10 161.363
R7612 XThR.Tn[2].n84 XThR.Tn[2].n83 161.3
R7613 XThR.Tn[2].n79 XThR.Tn[2].n78 161.3
R7614 XThR.Tn[2].n74 XThR.Tn[2].n73 161.3
R7615 XThR.Tn[2].n69 XThR.Tn[2].n68 161.3
R7616 XThR.Tn[2].n64 XThR.Tn[2].n63 161.3
R7617 XThR.Tn[2].n59 XThR.Tn[2].n58 161.3
R7618 XThR.Tn[2].n54 XThR.Tn[2].n53 161.3
R7619 XThR.Tn[2].n49 XThR.Tn[2].n48 161.3
R7620 XThR.Tn[2].n44 XThR.Tn[2].n43 161.3
R7621 XThR.Tn[2].n39 XThR.Tn[2].n38 161.3
R7622 XThR.Tn[2].n34 XThR.Tn[2].n33 161.3
R7623 XThR.Tn[2].n29 XThR.Tn[2].n28 161.3
R7624 XThR.Tn[2].n24 XThR.Tn[2].n23 161.3
R7625 XThR.Tn[2].n19 XThR.Tn[2].n18 161.3
R7626 XThR.Tn[2].n14 XThR.Tn[2].n13 161.3
R7627 XThR.Tn[2].n82 XThR.Tn[2].t65 161.106
R7628 XThR.Tn[2].n77 XThR.Tn[2].t72 161.106
R7629 XThR.Tn[2].n72 XThR.Tn[2].t51 161.106
R7630 XThR.Tn[2].n67 XThR.Tn[2].t36 161.106
R7631 XThR.Tn[2].n62 XThR.Tn[2].t64 161.106
R7632 XThR.Tn[2].n57 XThR.Tn[2].t26 161.106
R7633 XThR.Tn[2].n52 XThR.Tn[2].t69 161.106
R7634 XThR.Tn[2].n47 XThR.Tn[2].t49 161.106
R7635 XThR.Tn[2].n42 XThR.Tn[2].t35 161.106
R7636 XThR.Tn[2].n37 XThR.Tn[2].t41 161.106
R7637 XThR.Tn[2].n32 XThR.Tn[2].t25 161.106
R7638 XThR.Tn[2].n27 XThR.Tn[2].t50 161.106
R7639 XThR.Tn[2].n22 XThR.Tn[2].t23 161.106
R7640 XThR.Tn[2].n17 XThR.Tn[2].t67 161.106
R7641 XThR.Tn[2].n12 XThR.Tn[2].t31 161.106
R7642 XThR.Tn[2].n10 XThR.Tn[2].t14 161.106
R7643 XThR.Tn[2].n83 XThR.Tn[2].t38 159.978
R7644 XThR.Tn[2].n78 XThR.Tn[2].t46 159.978
R7645 XThR.Tn[2].n73 XThR.Tn[2].t29 159.978
R7646 XThR.Tn[2].n68 XThR.Tn[2].t13 159.978
R7647 XThR.Tn[2].n63 XThR.Tn[2].t37 159.978
R7648 XThR.Tn[2].n58 XThR.Tn[2].t63 159.978
R7649 XThR.Tn[2].n53 XThR.Tn[2].t45 159.978
R7650 XThR.Tn[2].n48 XThR.Tn[2].t27 159.978
R7651 XThR.Tn[2].n43 XThR.Tn[2].t12 159.978
R7652 XThR.Tn[2].n38 XThR.Tn[2].t20 159.978
R7653 XThR.Tn[2].n33 XThR.Tn[2].t62 159.978
R7654 XThR.Tn[2].n28 XThR.Tn[2].t28 159.978
R7655 XThR.Tn[2].n23 XThR.Tn[2].t60 159.978
R7656 XThR.Tn[2].n18 XThR.Tn[2].t43 159.978
R7657 XThR.Tn[2].n13 XThR.Tn[2].t66 159.978
R7658 XThR.Tn[2].n82 XThR.Tn[2].t53 145.038
R7659 XThR.Tn[2].n77 XThR.Tn[2].t19 145.038
R7660 XThR.Tn[2].n72 XThR.Tn[2].t59 145.038
R7661 XThR.Tn[2].n67 XThR.Tn[2].t42 145.038
R7662 XThR.Tn[2].n62 XThR.Tn[2].t73 145.038
R7663 XThR.Tn[2].n57 XThR.Tn[2].t52 145.038
R7664 XThR.Tn[2].n52 XThR.Tn[2].t61 145.038
R7665 XThR.Tn[2].n47 XThR.Tn[2].t44 145.038
R7666 XThR.Tn[2].n42 XThR.Tn[2].t39 145.038
R7667 XThR.Tn[2].n37 XThR.Tn[2].t70 145.038
R7668 XThR.Tn[2].n32 XThR.Tn[2].t34 145.038
R7669 XThR.Tn[2].n27 XThR.Tn[2].t58 145.038
R7670 XThR.Tn[2].n22 XThR.Tn[2].t32 145.038
R7671 XThR.Tn[2].n17 XThR.Tn[2].t15 145.038
R7672 XThR.Tn[2].n12 XThR.Tn[2].t40 145.038
R7673 XThR.Tn[2].n10 XThR.Tn[2].t21 145.038
R7674 XThR.Tn[2].n83 XThR.Tn[2].t71 143.911
R7675 XThR.Tn[2].n78 XThR.Tn[2].t33 143.911
R7676 XThR.Tn[2].n73 XThR.Tn[2].t17 143.911
R7677 XThR.Tn[2].n68 XThR.Tn[2].t56 143.911
R7678 XThR.Tn[2].n63 XThR.Tn[2].t24 143.911
R7679 XThR.Tn[2].n58 XThR.Tn[2].t68 143.911
R7680 XThR.Tn[2].n53 XThR.Tn[2].t18 143.911
R7681 XThR.Tn[2].n48 XThR.Tn[2].t57 143.911
R7682 XThR.Tn[2].n43 XThR.Tn[2].t54 143.911
R7683 XThR.Tn[2].n38 XThR.Tn[2].t22 143.911
R7684 XThR.Tn[2].n33 XThR.Tn[2].t48 143.911
R7685 XThR.Tn[2].n28 XThR.Tn[2].t16 143.911
R7686 XThR.Tn[2].n23 XThR.Tn[2].t47 143.911
R7687 XThR.Tn[2].n18 XThR.Tn[2].t30 143.911
R7688 XThR.Tn[2].n13 XThR.Tn[2].t55 143.911
R7689 XThR.Tn[2].n7 XThR.Tn[2].n5 135.249
R7690 XThR.Tn[2].n9 XThR.Tn[2].n3 98.982
R7691 XThR.Tn[2].n8 XThR.Tn[2].n4 98.982
R7692 XThR.Tn[2].n7 XThR.Tn[2].n6 98.982
R7693 XThR.Tn[2].n9 XThR.Tn[2].n8 36.2672
R7694 XThR.Tn[2].n8 XThR.Tn[2].n7 36.2672
R7695 XThR.Tn[2].n88 XThR.Tn[2].n9 32.6405
R7696 XThR.Tn[2].n1 XThR.Tn[2].t6 26.5955
R7697 XThR.Tn[2].n1 XThR.Tn[2].t2 26.5955
R7698 XThR.Tn[2].n0 XThR.Tn[2].t5 26.5955
R7699 XThR.Tn[2].n0 XThR.Tn[2].t3 26.5955
R7700 XThR.Tn[2].n3 XThR.Tn[2].t1 24.9236
R7701 XThR.Tn[2].n3 XThR.Tn[2].t8 24.9236
R7702 XThR.Tn[2].n4 XThR.Tn[2].t4 24.9236
R7703 XThR.Tn[2].n4 XThR.Tn[2].t10 24.9236
R7704 XThR.Tn[2].n5 XThR.Tn[2].t7 24.9236
R7705 XThR.Tn[2].n5 XThR.Tn[2].t9 24.9236
R7706 XThR.Tn[2].n6 XThR.Tn[2].t0 24.9236
R7707 XThR.Tn[2].n6 XThR.Tn[2].t11 24.9236
R7708 XThR.Tn[2] XThR.Tn[2].n2 23.3605
R7709 XThR.Tn[2] XThR.Tn[2].n88 6.7205
R7710 XThR.Tn[2].n88 XThR.Tn[2] 6.30883
R7711 XThR.Tn[2] XThR.Tn[2].n11 5.34038
R7712 XThR.Tn[2].n16 XThR.Tn[2].n15 4.5005
R7713 XThR.Tn[2].n21 XThR.Tn[2].n20 4.5005
R7714 XThR.Tn[2].n26 XThR.Tn[2].n25 4.5005
R7715 XThR.Tn[2].n31 XThR.Tn[2].n30 4.5005
R7716 XThR.Tn[2].n36 XThR.Tn[2].n35 4.5005
R7717 XThR.Tn[2].n41 XThR.Tn[2].n40 4.5005
R7718 XThR.Tn[2].n46 XThR.Tn[2].n45 4.5005
R7719 XThR.Tn[2].n51 XThR.Tn[2].n50 4.5005
R7720 XThR.Tn[2].n56 XThR.Tn[2].n55 4.5005
R7721 XThR.Tn[2].n61 XThR.Tn[2].n60 4.5005
R7722 XThR.Tn[2].n66 XThR.Tn[2].n65 4.5005
R7723 XThR.Tn[2].n71 XThR.Tn[2].n70 4.5005
R7724 XThR.Tn[2].n76 XThR.Tn[2].n75 4.5005
R7725 XThR.Tn[2].n81 XThR.Tn[2].n80 4.5005
R7726 XThR.Tn[2].n86 XThR.Tn[2].n85 4.5005
R7727 XThR.Tn[2].n87 XThR.Tn[2] 3.70586
R7728 XThR.Tn[2].n16 XThR.Tn[2] 2.52282
R7729 XThR.Tn[2].n21 XThR.Tn[2] 2.52282
R7730 XThR.Tn[2].n26 XThR.Tn[2] 2.52282
R7731 XThR.Tn[2].n31 XThR.Tn[2] 2.52282
R7732 XThR.Tn[2].n36 XThR.Tn[2] 2.52282
R7733 XThR.Tn[2].n41 XThR.Tn[2] 2.52282
R7734 XThR.Tn[2].n46 XThR.Tn[2] 2.52282
R7735 XThR.Tn[2].n51 XThR.Tn[2] 2.52282
R7736 XThR.Tn[2].n56 XThR.Tn[2] 2.52282
R7737 XThR.Tn[2].n61 XThR.Tn[2] 2.52282
R7738 XThR.Tn[2].n66 XThR.Tn[2] 2.52282
R7739 XThR.Tn[2].n71 XThR.Tn[2] 2.52282
R7740 XThR.Tn[2].n76 XThR.Tn[2] 2.52282
R7741 XThR.Tn[2].n81 XThR.Tn[2] 2.52282
R7742 XThR.Tn[2].n86 XThR.Tn[2] 2.52282
R7743 XThR.Tn[2].n84 XThR.Tn[2] 1.08677
R7744 XThR.Tn[2].n79 XThR.Tn[2] 1.08677
R7745 XThR.Tn[2].n74 XThR.Tn[2] 1.08677
R7746 XThR.Tn[2].n69 XThR.Tn[2] 1.08677
R7747 XThR.Tn[2].n64 XThR.Tn[2] 1.08677
R7748 XThR.Tn[2].n59 XThR.Tn[2] 1.08677
R7749 XThR.Tn[2].n54 XThR.Tn[2] 1.08677
R7750 XThR.Tn[2].n49 XThR.Tn[2] 1.08677
R7751 XThR.Tn[2].n44 XThR.Tn[2] 1.08677
R7752 XThR.Tn[2].n39 XThR.Tn[2] 1.08677
R7753 XThR.Tn[2].n34 XThR.Tn[2] 1.08677
R7754 XThR.Tn[2].n29 XThR.Tn[2] 1.08677
R7755 XThR.Tn[2].n24 XThR.Tn[2] 1.08677
R7756 XThR.Tn[2].n19 XThR.Tn[2] 1.08677
R7757 XThR.Tn[2].n14 XThR.Tn[2] 1.08677
R7758 XThR.Tn[2] XThR.Tn[2].n16 0.839786
R7759 XThR.Tn[2] XThR.Tn[2].n21 0.839786
R7760 XThR.Tn[2] XThR.Tn[2].n26 0.839786
R7761 XThR.Tn[2] XThR.Tn[2].n31 0.839786
R7762 XThR.Tn[2] XThR.Tn[2].n36 0.839786
R7763 XThR.Tn[2] XThR.Tn[2].n41 0.839786
R7764 XThR.Tn[2] XThR.Tn[2].n46 0.839786
R7765 XThR.Tn[2] XThR.Tn[2].n51 0.839786
R7766 XThR.Tn[2] XThR.Tn[2].n56 0.839786
R7767 XThR.Tn[2] XThR.Tn[2].n61 0.839786
R7768 XThR.Tn[2] XThR.Tn[2].n66 0.839786
R7769 XThR.Tn[2] XThR.Tn[2].n71 0.839786
R7770 XThR.Tn[2] XThR.Tn[2].n76 0.839786
R7771 XThR.Tn[2] XThR.Tn[2].n81 0.839786
R7772 XThR.Tn[2] XThR.Tn[2].n86 0.839786
R7773 XThR.Tn[2].n11 XThR.Tn[2] 0.499542
R7774 XThR.Tn[2].n85 XThR.Tn[2] 0.063
R7775 XThR.Tn[2].n80 XThR.Tn[2] 0.063
R7776 XThR.Tn[2].n75 XThR.Tn[2] 0.063
R7777 XThR.Tn[2].n70 XThR.Tn[2] 0.063
R7778 XThR.Tn[2].n65 XThR.Tn[2] 0.063
R7779 XThR.Tn[2].n60 XThR.Tn[2] 0.063
R7780 XThR.Tn[2].n55 XThR.Tn[2] 0.063
R7781 XThR.Tn[2].n50 XThR.Tn[2] 0.063
R7782 XThR.Tn[2].n45 XThR.Tn[2] 0.063
R7783 XThR.Tn[2].n40 XThR.Tn[2] 0.063
R7784 XThR.Tn[2].n35 XThR.Tn[2] 0.063
R7785 XThR.Tn[2].n30 XThR.Tn[2] 0.063
R7786 XThR.Tn[2].n25 XThR.Tn[2] 0.063
R7787 XThR.Tn[2].n20 XThR.Tn[2] 0.063
R7788 XThR.Tn[2].n15 XThR.Tn[2] 0.063
R7789 XThR.Tn[2].n87 XThR.Tn[2] 0.0540714
R7790 XThR.Tn[2] XThR.Tn[2].n87 0.038
R7791 XThR.Tn[2].n11 XThR.Tn[2] 0.0143889
R7792 XThR.Tn[2].n85 XThR.Tn[2].n84 0.00771154
R7793 XThR.Tn[2].n80 XThR.Tn[2].n79 0.00771154
R7794 XThR.Tn[2].n75 XThR.Tn[2].n74 0.00771154
R7795 XThR.Tn[2].n70 XThR.Tn[2].n69 0.00771154
R7796 XThR.Tn[2].n65 XThR.Tn[2].n64 0.00771154
R7797 XThR.Tn[2].n60 XThR.Tn[2].n59 0.00771154
R7798 XThR.Tn[2].n55 XThR.Tn[2].n54 0.00771154
R7799 XThR.Tn[2].n50 XThR.Tn[2].n49 0.00771154
R7800 XThR.Tn[2].n45 XThR.Tn[2].n44 0.00771154
R7801 XThR.Tn[2].n40 XThR.Tn[2].n39 0.00771154
R7802 XThR.Tn[2].n35 XThR.Tn[2].n34 0.00771154
R7803 XThR.Tn[2].n30 XThR.Tn[2].n29 0.00771154
R7804 XThR.Tn[2].n25 XThR.Tn[2].n24 0.00771154
R7805 XThR.Tn[2].n20 XThR.Tn[2].n19 0.00771154
R7806 XThR.Tn[2].n15 XThR.Tn[2].n14 0.00771154
R7807 VPWR.n2840 VPWR.n29 3532.94
R7808 VPWR.n2840 VPWR.n30 3532.94
R7809 VPWR.n2849 VPWR.n29 3532.94
R7810 VPWR.n2849 VPWR.n30 3532.94
R7811 VPWR.n2838 VPWR.n27 3532.94
R7812 VPWR.n2838 VPWR.n28 3532.94
R7813 VPWR.n2851 VPWR.n27 3532.94
R7814 VPWR.n2851 VPWR.n28 3532.94
R7815 VPWR.n2399 VPWR.t1561 1005.7
R7816 VPWR.t1779 VPWR.n504 1005.7
R7817 VPWR.t1628 VPWR.n2229 1005.7
R7818 VPWR.n658 VPWR.t1739 1005.7
R7819 VPWR.n2203 VPWR.t1462 1005.7
R7820 VPWR.t1569 VPWR.n696 1005.7
R7821 VPWR.t1529 VPWR.n2033 1005.7
R7822 VPWR.n850 VPWR.t1634 1005.7
R7823 VPWR.n2007 VPWR.t1454 1005.7
R7824 VPWR.t1641 VPWR.n888 1005.7
R7825 VPWR.n466 VPWR.t1446 1005.7
R7826 VPWR.t1749 VPWR.n1837 1005.7
R7827 VPWR.t1734 VPWR.n2425 1005.7
R7828 VPWR.n1042 VPWR.t1601 1005.7
R7829 VPWR.t1771 VPWR.n312 1005.7
R7830 VPWR.n1811 VPWR.t1718 1005.7
R7831 VPWR.n2610 VPWR.t1663 1005.7
R7832 VPWR.n1081 VPWR.t1547 1005.7
R7833 VPWR.t498 VPWR.n2328 983.14
R7834 VPWR.n2329 VPWR.t1918 983.14
R7835 VPWR.t1093 VPWR.n2338 983.14
R7836 VPWR.n2339 VPWR.t405 983.14
R7837 VPWR.t1263 VPWR.n2348 983.14
R7838 VPWR.n2349 VPWR.t858 983.14
R7839 VPWR.t454 VPWR.n2358 983.14
R7840 VPWR.n2359 VPWR.t952 983.14
R7841 VPWR.t653 VPWR.n2368 983.14
R7842 VPWR.n2369 VPWR.t334 983.14
R7843 VPWR.t1201 VPWR.n2378 983.14
R7844 VPWR.n2379 VPWR.t1867 983.14
R7845 VPWR.t193 VPWR.n2388 983.14
R7846 VPWR.n2389 VPWR.t1005 983.14
R7847 VPWR.t20 VPWR.n2398 983.14
R7848 VPWR.n561 VPWR.t839 983.14
R7849 VPWR.n560 VPWR.t1269 983.14
R7850 VPWR.n556 VPWR.t1069 983.14
R7851 VPWR.n552 VPWR.t6 983.14
R7852 VPWR.n548 VPWR.t1210 983.14
R7853 VPWR.n544 VPWR.t849 983.14
R7854 VPWR.n540 VPWR.t1911 983.14
R7855 VPWR.n536 VPWR.t541 983.14
R7856 VPWR.n532 VPWR.t665 983.14
R7857 VPWR.n528 VPWR.t385 983.14
R7858 VPWR.n524 VPWR.t476 983.14
R7859 VPWR.n520 VPWR.t66 983.14
R7860 VPWR.n516 VPWR.t1304 983.14
R7861 VPWR.n512 VPWR.t983 983.14
R7862 VPWR.n508 VPWR.t1253 983.14
R7863 VPWR.n2300 VPWR.t735 983.14
R7864 VPWR.n2299 VPWR.t1188 983.14
R7865 VPWR.n2290 VPWR.t1047 983.14
R7866 VPWR.n2289 VPWR.t681 983.14
R7867 VPWR.n2280 VPWR.t144 983.14
R7868 VPWR.n2279 VPWR.t52 983.14
R7869 VPWR.n2270 VPWR.t714 983.14
R7870 VPWR.n2269 VPWR.t930 983.14
R7871 VPWR.n2260 VPWR.t46 983.14
R7872 VPWR.n2259 VPWR.t322 983.14
R7873 VPWR.n2250 VPWR.t780 983.14
R7874 VPWR.n2249 VPWR.t1873 983.14
R7875 VPWR.n2240 VPWR.t179 983.14
R7876 VPWR.n2239 VPWR.t530 983.14
R7877 VPWR.n2230 VPWR.t1233 983.14
R7878 VPWR.t782 VPWR.n601 983.14
R7879 VPWR.t1114 VPWR.n605 983.14
R7880 VPWR.t1061 VPWR.n609 983.14
R7881 VPWR.t749 VPWR.n613 983.14
R7882 VPWR.t903 VPWR.n617 983.14
R7883 VPWR.t1823 VPWR.n621 983.14
R7884 VPWR.t1384 VPWR.n625 983.14
R7885 VPWR.t236 VPWR.n629 983.14
R7886 VPWR.t1281 VPWR.n633 983.14
R7887 VPWR.t354 VPWR.n637 983.14
R7888 VPWR.t486 VPWR.n641 983.14
R7889 VPWR.t630 VPWR.n645 983.14
R7890 VPWR.t1312 VPWR.n649 983.14
R7891 VPWR.t601 VPWR.n653 983.14
R7892 VPWR.t823 VPWR.n657 983.14
R7893 VPWR.t70 VPWR.n2132 983.14
R7894 VPWR.n2133 VPWR.t1151 983.14
R7895 VPWR.t1081 VPWR.n2142 983.14
R7896 VPWR.n2143 VPWR.t417 983.14
R7897 VPWR.t1323 VPWR.n2152 983.14
R7898 VPWR.n2153 VPWR.t1099 983.14
R7899 VPWR.t1899 VPWR.n2162 983.14
R7900 VPWR.n2163 VPWR.t222 983.14
R7901 VPWR.t794 VPWR.n2172 983.14
R7902 VPWR.n2173 VPWR.t346 983.14
R7903 VPWR.t1409 VPWR.n2182 983.14
R7904 VPWR.n2183 VPWR.t1163 983.14
R7905 VPWR.t254 VPWR.n2192 983.14
R7906 VPWR.n2193 VPWR.t999 983.14
R7907 VPWR.t16 VPWR.n2202 983.14
R7908 VPWR.n753 VPWR.t293 983.14
R7909 VPWR.n752 VPWR.t1916 983.14
R7910 VPWR.n748 VPWR.t1095 983.14
R7911 VPWR.n744 VPWR.t1402 983.14
R7912 VPWR.n740 VPWR.t1261 983.14
R7913 VPWR.n736 VPWR.t64 983.14
R7914 VPWR.n732 VPWR.t452 983.14
R7915 VPWR.n728 VPWR.t950 983.14
R7916 VPWR.n724 VPWR.t651 983.14
R7917 VPWR.n720 VPWR.t332 983.14
R7918 VPWR.n716 VPWR.t558 983.14
R7919 VPWR.n712 VPWR.t1865 983.14
R7920 VPWR.n708 VPWR.t191 983.14
R7921 VPWR.n704 VPWR.t1003 983.14
R7922 VPWR.n700 VPWR.t18 983.14
R7923 VPWR.n2104 VPWR.t642 983.14
R7924 VPWR.n2103 VPWR.t506 983.14
R7925 VPWR.n2094 VPWR.t1089 983.14
R7926 VPWR.n2093 VPWR.t407 983.14
R7927 VPWR.n2084 VPWR.t445 983.14
R7928 VPWR.n2083 VPWR.t864 983.14
R7929 VPWR.n2074 VPWR.t460 983.14
R7930 VPWR.n2073 VPWR.t226 983.14
R7931 VPWR.n2064 VPWR.t562 983.14
R7932 VPWR.n2063 VPWR.t340 983.14
R7933 VPWR.n2054 VPWR.t532 983.14
R7934 VPWR.n2053 VPWR.t1019 983.14
R7935 VPWR.n2044 VPWR.t244 983.14
R7936 VPWR.n2043 VPWR.t1011 983.14
R7937 VPWR.n2034 VPWR.t22 983.14
R7938 VPWR.t733 VPWR.n793 983.14
R7939 VPWR.t1186 VPWR.n797 983.14
R7940 VPWR.t1049 VPWR.n801 983.14
R7941 VPWR.t677 VPWR.n805 983.14
R7942 VPWR.t142 VPWR.n809 983.14
R7943 VPWR.t50 VPWR.n813 983.14
R7944 VPWR.t712 VPWR.n817 983.14
R7945 VPWR.t610 VPWR.n821 983.14
R7946 VPWR.t44 VPWR.n825 983.14
R7947 VPWR.t2 VPWR.n829 983.14
R7948 VPWR.t778 VPWR.n833 983.14
R7949 VPWR.t1871 VPWR.n837 983.14
R7950 VPWR.t976 VPWR.n841 983.14
R7951 VPWR.t40 VPWR.n845 983.14
R7952 VPWR.t1229 VPWR.n849 983.14
R7953 VPWR.t72 VPWR.n1936 983.14
R7954 VPWR.n1937 VPWR.t1153 983.14
R7955 VPWR.t1079 VPWR.n1946 983.14
R7956 VPWR.n1947 VPWR.t685 983.14
R7957 VPWR.t1325 VPWR.n1956 983.14
R7958 VPWR.n1957 VPWR.t1101 983.14
R7959 VPWR.t1901 VPWR.n1966 983.14
R7960 VPWR.n1967 VPWR.t224 983.14
R7961 VPWR.t796 VPWR.n1976 983.14
R7962 VPWR.n1977 VPWR.t348 983.14
R7963 VPWR.t1411 VPWR.n1986 983.14
R7964 VPWR.n1987 VPWR.t1805 983.14
R7965 VPWR.t256 VPWR.n1996 983.14
R7966 VPWR.n1997 VPWR.t1001 983.14
R7967 VPWR.t1243 VPWR.n2006 983.14
R7968 VPWR.n945 VPWR.t731 983.14
R7969 VPWR.n944 VPWR.t1184 983.14
R7970 VPWR.n940 VPWR.t1051 983.14
R7971 VPWR.n936 VPWR.t675 983.14
R7972 VPWR.n932 VPWR.t928 983.14
R7973 VPWR.n928 VPWR.t48 983.14
R7974 VPWR.n924 VPWR.t710 983.14
R7975 VPWR.n920 VPWR.t606 983.14
R7976 VPWR.n916 VPWR.t42 983.14
R7977 VPWR.n912 VPWR.t0 983.14
R7978 VPWR.n908 VPWR.t776 983.14
R7979 VPWR.n904 VPWR.t1869 983.14
R7980 VPWR.n900 VPWR.t972 983.14
R7981 VPWR.n896 VPWR.t38 983.14
R7982 VPWR.n892 VPWR.t1227 983.14
R7983 VPWR.t74 VPWR.n409 983.14
R7984 VPWR.t1155 VPWR.n413 983.14
R7985 VPWR.t1077 VPWR.n417 983.14
R7986 VPWR.t689 VPWR.n421 983.14
R7987 VPWR.t1327 VPWR.n425 983.14
R7988 VPWR.t1103 VPWR.n429 983.14
R7989 VPWR.t1903 VPWR.n433 983.14
R7990 VPWR.t1925 VPWR.n437 983.14
R7991 VPWR.t798 VPWR.n441 983.14
R7992 VPWR.t350 VPWR.n445 983.14
R7993 VPWR.t1120 VPWR.n449 983.14
R7994 VPWR.t1807 VPWR.n453 983.14
R7995 VPWR.t258 VPWR.n457 983.14
R7996 VPWR.t1193 VPWR.n461 983.14
R7997 VPWR.t1247 VPWR.n465 983.14
R7998 VPWR.n1908 VPWR.t1128 983.14
R7999 VPWR.n1907 VPWR.t1275 983.14
R8000 VPWR.n1898 VPWR.t1063 983.14
R8001 VPWR.n1897 VPWR.t10 983.14
R8002 VPWR.n1888 VPWR.t899 983.14
R8003 VPWR.n1887 VPWR.t1819 983.14
R8004 VPWR.n1878 VPWR.t1380 983.14
R8005 VPWR.n1877 VPWR.t234 983.14
R8006 VPWR.n1868 VPWR.t1277 983.14
R8007 VPWR.n1867 VPWR.t389 983.14
R8008 VPWR.n1858 VPWR.t482 983.14
R8009 VPWR.n1857 VPWR.t628 983.14
R8010 VPWR.n1848 VPWR.t1310 983.14
R8011 VPWR.n1847 VPWR.t599 983.14
R8012 VPWR.n1838 VPWR.t821 983.14
R8013 VPWR.n2496 VPWR.t784 983.14
R8014 VPWR.n2495 VPWR.t1116 983.14
R8015 VPWR.n2486 VPWR.t1059 983.14
R8016 VPWR.n2485 VPWR.t753 983.14
R8017 VPWR.n2476 VPWR.t905 983.14
R8018 VPWR.n2475 VPWR.t1825 983.14
R8019 VPWR.n2466 VPWR.t1386 983.14
R8020 VPWR.n2465 VPWR.t238 983.14
R8021 VPWR.n2456 VPWR.t1283 983.14
R8022 VPWR.n2455 VPWR.t356 983.14
R8023 VPWR.n2446 VPWR.t488 983.14
R8024 VPWR.n2445 VPWR.t632 983.14
R8025 VPWR.n2436 VPWR.t1314 983.14
R8026 VPWR.n2435 VPWR.t987 983.14
R8027 VPWR.n2426 VPWR.t827 983.14
R8028 VPWR.t285 VPWR.n985 983.14
R8029 VPWR.t514 VPWR.n989 983.14
R8030 VPWR.t1041 VPWR.n993 983.14
R8031 VPWR.t1398 VPWR.n997 983.14
R8032 VPWR.t150 VPWR.n1001 983.14
R8033 VPWR.t58 VPWR.n1005 983.14
R8034 VPWR.t720 VPWR.n1009 983.14
R8035 VPWR.t934 VPWR.n1013 983.14
R8036 VPWR.t524 VPWR.n1017 983.14
R8037 VPWR.t324 VPWR.n1021 983.14
R8038 VPWR.t552 VPWR.n1025 983.14
R8039 VPWR.t1875 VPWR.n1029 983.14
R8040 VPWR.t183 VPWR.n1033 983.14
R8041 VPWR.t634 VPWR.n1037 983.14
R8042 VPWR.t1239 VPWR.n1041 983.14
R8043 VPWR.n369 VPWR.t841 983.14
R8044 VPWR.n368 VPWR.t1271 983.14
R8045 VPWR.n364 VPWR.t1067 983.14
R8046 VPWR.n360 VPWR.t8 983.14
R8047 VPWR.n356 VPWR.t1212 983.14
R8048 VPWR.n352 VPWR.t1815 983.14
R8049 VPWR.n348 VPWR.t1376 983.14
R8050 VPWR.n344 VPWR.t545 983.14
R8051 VPWR.n340 VPWR.t667 983.14
R8052 VPWR.n336 VPWR.t387 983.14
R8053 VPWR.n332 VPWR.t478 983.14
R8054 VPWR.n328 VPWR.t68 983.14
R8055 VPWR.n324 VPWR.t1308 983.14
R8056 VPWR.n320 VPWR.t985 983.14
R8057 VPWR.n316 VPWR.t1255 983.14
R8058 VPWR.t1674 VPWR.n1487 983.14
R8059 VPWR.t1784 VPWR.n1494 983.14
R8060 VPWR.t1555 VPWR.n1500 983.14
R8061 VPWR.t1657 VPWR.n1511 983.14
R8062 VPWR.n1512 VPWR.t1682 983.14
R8063 VPWR.t1430 VPWR.n1525 983.14
R8064 VPWR.n1526 VPWR.t1552 983.14
R8065 VPWR.t1693 VPWR.n1539 983.14
R8066 VPWR.n1540 VPWR.t1715 983.14
R8067 VPWR.n1555 VPWR.t1449 983.14
R8068 VPWR.n1554 VPWR.t1582 983.14
R8069 VPWR.n1780 VPWR.t1623 983.14
R8070 VPWR.n1779 VPWR.t1459 983.14
R8071 VPWR.n1768 VPWR.t1496 983.14
R8072 VPWR.t1604 VPWR.n1810 983.14
R8073 VPWR.t1610 VPWR.n2525 983.14
R8074 VPWR.n2526 VPWR.t1725 983.14
R8075 VPWR.t1487 VPWR.n2537 983.14
R8076 VPWR.n2538 VPWR.t1595 983.14
R8077 VPWR.t1607 VPWR.n2549 983.14
R8078 VPWR.n2550 VPWR.t1763 983.14
R8079 VPWR.t1484 VPWR.n2561 983.14
R8080 VPWR.n2562 VPWR.t1644 983.14
R8081 VPWR.t1660 VPWR.n2573 983.14
R8082 VPWR.n2574 VPWR.t1790 983.14
R8083 VPWR.t1534 VPWR.n2585 983.14
R8084 VPWR.n2586 VPWR.t1564 983.14
R8085 VPWR.t1414 VPWR.n2597 983.14
R8086 VPWR.n2598 VPWR.t1433 983.14
R8087 VPWR.t1558 VPWR.n2609 983.14
R8088 VPWR.n1613 VPWR.t1493 983.14
R8089 VPWR.n1612 VPWR.t1598 983.14
R8090 VPWR.t1760 VPWR.n1201 983.14
R8091 VPWR.t1478 VPWR.n1204 983.14
R8092 VPWR.n1239 VPWR.t1490 983.14
R8093 VPWR.n1238 VPWR.t1649 983.14
R8094 VPWR.n1235 VPWR.t1752 983.14
R8095 VPWR.n1232 VPWR.t1518 983.14
R8096 VPWR.n1224 VPWR.t1544 983.14
R8097 VPWR.n1221 VPWR.t1666 983.14
R8098 VPWR.n1218 VPWR.t1417 983.14
R8099 VPWR.n1210 VPWR.t1438 983.14
R8100 VPWR.n1207 VPWR.t1679 983.14
R8101 VPWR.n1759 VPWR.t1710 983.14
R8102 VPWR.n1758 VPWR.t1424 983.14
R8103 VPWR.n1327 VPWR.t1348 877.144
R8104 VPWR.n2742 VPWR.t196 877.144
R8105 VPWR.n1141 VPWR.t1729 738.074
R8106 VPWR.n118 VPWR.t1466 738.074
R8107 VPWR.n309 VPWR.t584 738.074
R8108 VPWR.n87 VPWR.t1535 738.074
R8109 VPWR.n365 VPWR.t842 738.074
R8110 VPWR.n117 VPWR.t1611 738.074
R8111 VPWR.n982 VPWR.t567 738.074
R8112 VPWR.n375 VPWR.t578 738.074
R8113 VPWR.n376 VPWR.t785 738.074
R8114 VPWR.n337 VPWR.t546 738.074
R8115 VPWR.n94 VPWR.t1645 738.074
R8116 VPWR.n990 VPWR.t515 738.074
R8117 VPWR.n388 VPWR.t1387 738.074
R8118 VPWR.n341 VPWR.t1377 738.074
R8119 VPWR.n99 VPWR.t1485 738.074
R8120 VPWR.n951 VPWR.t582 738.074
R8121 VPWR.n952 VPWR.t1129 738.074
R8122 VPWR.n955 VPWR.t1276 738.074
R8123 VPWR.n406 VPWR.t588 738.074
R8124 VPWR.n410 VPWR.t75 738.074
R8125 VPWR.n414 VPWR.t1156 738.074
R8126 VPWR.n384 VPWR.t906 738.074
R8127 VPWR.n349 VPWR.t1213 738.074
R8128 VPWR.n105 VPWR.t1608 738.074
R8129 VPWR.n956 VPWR.t1064 738.074
R8130 VPWR.n422 VPWR.t690 738.074
R8131 VPWR.n383 VPWR.t754 738.074
R8132 VPWR.n353 VPWR.t9 738.074
R8133 VPWR.n106 VPWR.t1596 738.074
R8134 VPWR.n500 VPWR.t596 738.074
R8135 VPWR.n499 VPWR.t499 738.074
R8136 VPWR.n496 VPWR.t1919 738.074
R8137 VPWR.n495 VPWR.t1094 738.074
R8138 VPWR.n491 VPWR.t1264 738.074
R8139 VPWR.n488 VPWR.t859 738.074
R8140 VPWR.n487 VPWR.t455 738.074
R8141 VPWR.n484 VPWR.t953 738.074
R8142 VPWR.n483 VPWR.t654 738.074
R8143 VPWR.n480 VPWR.t335 738.074
R8144 VPWR.n479 VPWR.t1202 738.074
R8145 VPWR.n476 VPWR.t1868 738.074
R8146 VPWR.n475 VPWR.t194 738.074
R8147 VPWR.n472 VPWR.t1006 738.074
R8148 VPWR.n471 VPWR.t21 738.074
R8149 VPWR.n492 VPWR.t406 738.074
R8150 VPWR.n501 VPWR.t586 738.074
R8151 VPWR.n557 VPWR.t840 738.074
R8152 VPWR.n553 VPWR.t1270 738.074
R8153 VPWR.n549 VPWR.t1070 738.074
R8154 VPWR.n541 VPWR.t1211 738.074
R8155 VPWR.n537 VPWR.t850 738.074
R8156 VPWR.n533 VPWR.t1912 738.074
R8157 VPWR.n529 VPWR.t542 738.074
R8158 VPWR.n525 VPWR.t666 738.074
R8159 VPWR.n521 VPWR.t386 738.074
R8160 VPWR.n517 VPWR.t477 738.074
R8161 VPWR.n513 VPWR.t67 738.074
R8162 VPWR.n509 VPWR.t1305 738.074
R8163 VPWR.n505 VPWR.t984 738.074
R8164 VPWR.n502 VPWR.t1254 738.074
R8165 VPWR.n545 VPWR.t7 738.074
R8166 VPWR.n567 VPWR.t572 738.074
R8167 VPWR.n568 VPWR.t736 738.074
R8168 VPWR.n571 VPWR.t1189 738.074
R8169 VPWR.n572 VPWR.t1048 738.074
R8170 VPWR.n576 VPWR.t145 738.074
R8171 VPWR.n579 VPWR.t53 738.074
R8172 VPWR.n580 VPWR.t715 738.074
R8173 VPWR.n583 VPWR.t931 738.074
R8174 VPWR.n584 VPWR.t47 738.074
R8175 VPWR.n587 VPWR.t323 738.074
R8176 VPWR.n588 VPWR.t781 738.074
R8177 VPWR.n591 VPWR.t1874 738.074
R8178 VPWR.n592 VPWR.t180 738.074
R8179 VPWR.n595 VPWR.t531 738.074
R8180 VPWR.n596 VPWR.t1234 738.074
R8181 VPWR.n575 VPWR.t682 738.074
R8182 VPWR.n598 VPWR.t580 738.074
R8183 VPWR.n602 VPWR.t783 738.074
R8184 VPWR.n606 VPWR.t1115 738.074
R8185 VPWR.n610 VPWR.t1062 738.074
R8186 VPWR.n618 VPWR.t904 738.074
R8187 VPWR.n622 VPWR.t1824 738.074
R8188 VPWR.n626 VPWR.t1385 738.074
R8189 VPWR.n630 VPWR.t237 738.074
R8190 VPWR.n634 VPWR.t1282 738.074
R8191 VPWR.n638 VPWR.t355 738.074
R8192 VPWR.n642 VPWR.t487 738.074
R8193 VPWR.n646 VPWR.t631 738.074
R8194 VPWR.n650 VPWR.t1313 738.074
R8195 VPWR.n654 VPWR.t602 738.074
R8196 VPWR.n597 VPWR.t824 738.074
R8197 VPWR.n614 VPWR.t750 738.074
R8198 VPWR.n692 VPWR.t592 738.074
R8199 VPWR.n691 VPWR.t71 738.074
R8200 VPWR.n688 VPWR.t1152 738.074
R8201 VPWR.n687 VPWR.t1082 738.074
R8202 VPWR.n683 VPWR.t1324 738.074
R8203 VPWR.n680 VPWR.t1100 738.074
R8204 VPWR.n679 VPWR.t1900 738.074
R8205 VPWR.n676 VPWR.t223 738.074
R8206 VPWR.n675 VPWR.t795 738.074
R8207 VPWR.n672 VPWR.t347 738.074
R8208 VPWR.n671 VPWR.t1410 738.074
R8209 VPWR.n668 VPWR.t1164 738.074
R8210 VPWR.n667 VPWR.t255 738.074
R8211 VPWR.n664 VPWR.t1000 738.074
R8212 VPWR.n663 VPWR.t17 738.074
R8213 VPWR.n684 VPWR.t418 738.074
R8214 VPWR.n693 VPWR.t598 738.074
R8215 VPWR.n749 VPWR.t294 738.074
R8216 VPWR.n745 VPWR.t1917 738.074
R8217 VPWR.n741 VPWR.t1096 738.074
R8218 VPWR.n733 VPWR.t1262 738.074
R8219 VPWR.n729 VPWR.t65 738.074
R8220 VPWR.n725 VPWR.t453 738.074
R8221 VPWR.n721 VPWR.t951 738.074
R8222 VPWR.n717 VPWR.t652 738.074
R8223 VPWR.n713 VPWR.t333 738.074
R8224 VPWR.n709 VPWR.t559 738.074
R8225 VPWR.n705 VPWR.t1866 738.074
R8226 VPWR.n701 VPWR.t192 738.074
R8227 VPWR.n697 VPWR.t1004 738.074
R8228 VPWR.n694 VPWR.t19 738.074
R8229 VPWR.n737 VPWR.t1403 738.074
R8230 VPWR.n759 VPWR.t594 738.074
R8231 VPWR.n760 VPWR.t643 738.074
R8232 VPWR.n763 VPWR.t507 738.074
R8233 VPWR.n764 VPWR.t1090 738.074
R8234 VPWR.n768 VPWR.t446 738.074
R8235 VPWR.n771 VPWR.t865 738.074
R8236 VPWR.n772 VPWR.t461 738.074
R8237 VPWR.n775 VPWR.t227 738.074
R8238 VPWR.n776 VPWR.t563 738.074
R8239 VPWR.n779 VPWR.t341 738.074
R8240 VPWR.n780 VPWR.t533 738.074
R8241 VPWR.n783 VPWR.t1020 738.074
R8242 VPWR.n784 VPWR.t245 738.074
R8243 VPWR.n787 VPWR.t1012 738.074
R8244 VPWR.n788 VPWR.t23 738.074
R8245 VPWR.n767 VPWR.t408 738.074
R8246 VPWR.n790 VPWR.t574 738.074
R8247 VPWR.n794 VPWR.t734 738.074
R8248 VPWR.n798 VPWR.t1187 738.074
R8249 VPWR.n802 VPWR.t1050 738.074
R8250 VPWR.n810 VPWR.t143 738.074
R8251 VPWR.n814 VPWR.t51 738.074
R8252 VPWR.n818 VPWR.t713 738.074
R8253 VPWR.n822 VPWR.t611 738.074
R8254 VPWR.n826 VPWR.t45 738.074
R8255 VPWR.n830 VPWR.t3 738.074
R8256 VPWR.n834 VPWR.t779 738.074
R8257 VPWR.n838 VPWR.t1872 738.074
R8258 VPWR.n842 VPWR.t977 738.074
R8259 VPWR.n846 VPWR.t41 738.074
R8260 VPWR.n789 VPWR.t1230 738.074
R8261 VPWR.n806 VPWR.t678 738.074
R8262 VPWR.n884 VPWR.t590 738.074
R8263 VPWR.n883 VPWR.t73 738.074
R8264 VPWR.n880 VPWR.t1154 738.074
R8265 VPWR.n879 VPWR.t1080 738.074
R8266 VPWR.n875 VPWR.t1326 738.074
R8267 VPWR.n872 VPWR.t1102 738.074
R8268 VPWR.n871 VPWR.t1902 738.074
R8269 VPWR.n868 VPWR.t225 738.074
R8270 VPWR.n867 VPWR.t797 738.074
R8271 VPWR.n864 VPWR.t349 738.074
R8272 VPWR.n863 VPWR.t1412 738.074
R8273 VPWR.n860 VPWR.t1806 738.074
R8274 VPWR.n859 VPWR.t257 738.074
R8275 VPWR.n856 VPWR.t1002 738.074
R8276 VPWR.n855 VPWR.t1244 738.074
R8277 VPWR.n876 VPWR.t686 738.074
R8278 VPWR.n885 VPWR.t576 738.074
R8279 VPWR.n941 VPWR.t732 738.074
R8280 VPWR.n937 VPWR.t1185 738.074
R8281 VPWR.n933 VPWR.t1052 738.074
R8282 VPWR.n925 VPWR.t929 738.074
R8283 VPWR.n921 VPWR.t49 738.074
R8284 VPWR.n917 VPWR.t711 738.074
R8285 VPWR.n913 VPWR.t607 738.074
R8286 VPWR.n909 VPWR.t43 738.074
R8287 VPWR.n905 VPWR.t1 738.074
R8288 VPWR.n901 VPWR.t777 738.074
R8289 VPWR.n897 VPWR.t1870 738.074
R8290 VPWR.n893 VPWR.t973 738.074
R8291 VPWR.n889 VPWR.t39 738.074
R8292 VPWR.n886 VPWR.t1228 738.074
R8293 VPWR.n929 VPWR.t676 738.074
R8294 VPWR.n959 VPWR.t11 738.074
R8295 VPWR.n998 VPWR.t1399 738.074
R8296 VPWR.n1198 VPWR.t1479 738.074
R8297 VPWR.n418 VPWR.t1078 738.074
R8298 VPWR.n380 VPWR.t1060 738.074
R8299 VPWR.n357 VPWR.t1068 738.074
R8300 VPWR.n111 VPWR.t1488 738.074
R8301 VPWR.n994 VPWR.t1042 738.074
R8302 VPWR.n1202 VPWR.t1761 738.074
R8303 VPWR.n960 VPWR.t900 738.074
R8304 VPWR.n1002 VPWR.t151 738.074
R8305 VPWR.n1236 VPWR.t1491 738.074
R8306 VPWR.n426 VPWR.t1328 738.074
R8307 VPWR.n434 VPWR.t1904 738.074
R8308 VPWR.n438 VPWR.t1926 738.074
R8309 VPWR.n442 VPWR.t799 738.074
R8310 VPWR.n446 VPWR.t351 738.074
R8311 VPWR.n450 VPWR.t1121 738.074
R8312 VPWR.n454 VPWR.t1808 738.074
R8313 VPWR.n458 VPWR.t259 738.074
R8314 VPWR.n462 VPWR.t1194 738.074
R8315 VPWR.n405 VPWR.t1248 738.074
R8316 VPWR.n430 VPWR.t1104 738.074
R8317 VPWR.n387 VPWR.t1826 738.074
R8318 VPWR.n345 VPWR.t1816 738.074
R8319 VPWR.n100 VPWR.t1764 738.074
R8320 VPWR.n1006 VPWR.t59 738.074
R8321 VPWR.n1233 VPWR.t1650 738.074
R8322 VPWR.n963 VPWR.t1820 738.074
R8323 VPWR.n967 VPWR.t235 738.074
R8324 VPWR.n968 VPWR.t1278 738.074
R8325 VPWR.n971 VPWR.t390 738.074
R8326 VPWR.n972 VPWR.t483 738.074
R8327 VPWR.n975 VPWR.t629 738.074
R8328 VPWR.n976 VPWR.t1311 738.074
R8329 VPWR.n979 VPWR.t600 738.074
R8330 VPWR.n980 VPWR.t822 738.074
R8331 VPWR.n964 VPWR.t1381 738.074
R8332 VPWR.n1010 VPWR.t721 738.074
R8333 VPWR.n1225 VPWR.t1753 738.074
R8334 VPWR.n379 VPWR.t1117 738.074
R8335 VPWR.n361 VPWR.t1272 738.074
R8336 VPWR.n112 VPWR.t1726 738.074
R8337 VPWR.n1199 VPWR.t1599 738.074
R8338 VPWR.n1014 VPWR.t935 738.074
R8339 VPWR.n1222 VPWR.t1519 738.074
R8340 VPWR.n391 VPWR.t239 738.074
R8341 VPWR.n395 VPWR.t357 738.074
R8342 VPWR.n396 VPWR.t489 738.074
R8343 VPWR.n399 VPWR.t633 738.074
R8344 VPWR.n400 VPWR.t1315 738.074
R8345 VPWR.n403 VPWR.t988 738.074
R8346 VPWR.n404 VPWR.t828 738.074
R8347 VPWR.n392 VPWR.t1284 738.074
R8348 VPWR.n333 VPWR.t668 738.074
R8349 VPWR.n93 VPWR.t1661 738.074
R8350 VPWR.n1219 VPWR.t1545 738.074
R8351 VPWR.n1018 VPWR.t525 738.074
R8352 VPWR.n1022 VPWR.t325 738.074
R8353 VPWR.n1026 VPWR.t553 738.074
R8354 VPWR.n1030 VPWR.t1876 738.074
R8355 VPWR.n1034 VPWR.t184 738.074
R8356 VPWR.n1038 VPWR.t635 738.074
R8357 VPWR.n981 VPWR.t1240 738.074
R8358 VPWR.n986 VPWR.t286 738.074
R8359 VPWR.n1142 VPWR.t1494 738.074
R8360 VPWR.n329 VPWR.t388 738.074
R8361 VPWR.n88 VPWR.t1791 738.074
R8362 VPWR.n1211 VPWR.t1667 738.074
R8363 VPWR.n1208 VPWR.t1418 738.074
R8364 VPWR.n325 VPWR.t479 738.074
R8365 VPWR.n321 VPWR.t69 738.074
R8366 VPWR.n313 VPWR.t986 738.074
R8367 VPWR.n310 VPWR.t1256 738.074
R8368 VPWR.n317 VPWR.t1309 738.074
R8369 VPWR.n1077 VPWR.t1680 738.074
R8370 VPWR.n1205 VPWR.t1439 738.074
R8371 VPWR.n82 VPWR.t1565 738.074
R8372 VPWR.n81 VPWR.t1415 738.074
R8373 VPWR.n76 VPWR.t1434 738.074
R8374 VPWR.n75 VPWR.t1559 738.074
R8375 VPWR.n1078 VPWR.t1711 738.074
R8376 VPWR.n1080 VPWR.t1425 738.074
R8377 VPWR.n1080 VPWR.t1548 646.071
R8378 VPWR.n1141 VPWR.t1444 646.071
R8379 VPWR.n1078 VPWR.t1703 646.071
R8380 VPWR.n75 VPWR.t1664 646.071
R8381 VPWR.n81 VPWR.t1788 646.071
R8382 VPWR.n118 VPWR.t1573 646.071
R8383 VPWR.n1072 VPWR.t190 646.071
R8384 VPWR.n1250 VPWR.t664 646.071
R8385 VPWR.n317 VPWR.t992 646.071
R8386 VPWR.n309 VPWR.t789 646.071
R8387 VPWR.n325 VPWR.t1026 646.071
R8388 VPWR.n87 VPWR.t1527 646.071
R8389 VPWR.n1172 VPWR.t1846 646.071
R8390 VPWR.n365 VPWR.t1113 646.071
R8391 VPWR.n117 VPWR.t1708 646.071
R8392 VPWR.n986 VPWR.t519 646.071
R8393 VPWR.n982 VPWR.t501 646.071
R8394 VPWR.n1018 VPWR.t337 646.071
R8395 VPWR.n392 VPWR.t367 646.071
R8396 VPWR.n375 VPWR.t662 646.071
R8397 VPWR.n376 VPWR.t1335 646.071
R8398 VPWR.n391 VPWR.t296 646.071
R8399 VPWR.n337 VPWR.t1280 646.071
R8400 VPWR.n94 VPWR.t1632 646.071
R8401 VPWR.n990 VPWR.t1076 646.071
R8402 VPWR.n388 VPWR.t939 646.071
R8403 VPWR.n341 VPWR.t613 646.071
R8404 VPWR.n99 VPWR.t1504 646.071
R8405 VPWR.n964 VPWR.t933 646.071
R8406 VPWR.n951 VPWR.t791 646.071
R8407 VPWR.n952 VPWR.t1119 646.071
R8408 VPWR.n955 VPWR.t1040 646.071
R8409 VPWR.n963 VPWR.t1389 646.071
R8410 VPWR.n430 VPWR.t1910 646.071
R8411 VPWR.n406 VPWR.t838 646.071
R8412 VPWR.n410 VPWR.t709 646.071
R8413 VPWR.n414 VPWR.t1054 646.071
R8414 VPWR.n426 VPWR.t848 646.071
R8415 VPWR.n384 VPWR.t1802 646.071
R8416 VPWR.n349 VPWR.t1822 646.071
R8417 VPWR.n105 VPWR.t1745 646.071
R8418 VPWR.n956 VPWR.t680 646.071
R8419 VPWR.n422 VPWR.t1183 646.071
R8420 VPWR.n383 VPWR.t1146 646.071
R8421 VPWR.n353 VPWR.t902 646.071
R8422 VPWR.n106 VPWR.t1590 646.071
R8423 VPWR.n492 VPWR.t444 646.071
R8424 VPWR.n500 VPWR.t645 646.071
R8425 VPWR.n499 VPWR.t505 646.071
R8426 VPWR.n496 VPWR.t1072 646.071
R8427 VPWR.n495 VPWR.t692 646.071
R8428 VPWR.n491 VPWR.t863 646.071
R8429 VPWR.n488 VPWR.t459 646.071
R8430 VPWR.n487 VPWR.t1930 646.071
R8431 VPWR.n484 VPWR.t561 646.071
R8432 VPWR.n483 VPWR.t343 646.071
R8433 VPWR.n480 VPWR.t1206 646.071
R8434 VPWR.n479 VPWR.t1022 646.071
R8435 VPWR.n476 VPWR.t1303 646.071
R8436 VPWR.n475 VPWR.t1014 646.071
R8437 VPWR.n472 VPWR.t1250 646.071
R8438 VPWR.n471 VPWR.t1562 646.071
R8439 VPWR.n545 VPWR.t898 646.071
R8440 VPWR.n501 VPWR.t787 646.071
R8441 VPWR.n557 VPWR.t1274 646.071
R8442 VPWR.n553 VPWR.t1046 646.071
R8443 VPWR.n549 VPWR.t672 646.071
R8444 VPWR.n541 VPWR.t1818 646.071
R8445 VPWR.n537 VPWR.t1379 646.071
R8446 VPWR.n533 VPWR.t609 646.071
R8447 VPWR.n529 VPWR.t670 646.071
R8448 VPWR.n525 VPWR.t359 646.071
R8449 VPWR.n521 VPWR.t481 646.071
R8450 VPWR.n517 VPWR.t1024 646.071
R8451 VPWR.n513 VPWR.t975 646.071
R8452 VPWR.n509 VPWR.t990 646.071
R8453 VPWR.n505 VPWR.t1224 646.071
R8454 VPWR.n502 VPWR.t1780 646.071
R8455 VPWR.n575 VPWR.t153 646.071
R8456 VPWR.n567 VPWR.t292 646.071
R8457 VPWR.n568 VPWR.t517 646.071
R8458 VPWR.n571 VPWR.t1084 646.071
R8459 VPWR.n572 VPWR.t414 646.071
R8460 VPWR.n576 VPWR.t61 646.071
R8461 VPWR.n579 VPWR.t723 646.071
R8462 VPWR.n580 VPWR.t219 646.071
R8463 VPWR.n583 VPWR.t527 646.071
R8464 VPWR.n584 VPWR.t331 646.071
R8465 VPWR.n587 VPWR.t555 646.071
R8466 VPWR.n588 VPWR.t1864 646.071
R8467 VPWR.n591 VPWR.t251 646.071
R8468 VPWR.n592 VPWR.t641 646.071
R8469 VPWR.n595 VPWR.t13 646.071
R8470 VPWR.n596 VPWR.t1629 646.071
R8471 VPWR.n614 VPWR.t1144 646.071
R8472 VPWR.n598 VPWR.t793 646.071
R8473 VPWR.n602 VPWR.t910 646.071
R8474 VPWR.n606 VPWR.t1038 646.071
R8475 VPWR.n610 VPWR.t684 646.071
R8476 VPWR.n618 VPWR.t1800 646.071
R8477 VPWR.n622 VPWR.t1391 646.071
R8478 VPWR.n626 VPWR.t937 646.071
R8479 VPWR.n630 VPWR.t1288 646.071
R8480 VPWR.n634 VPWR.t365 646.071
R8481 VPWR.n638 VPWR.t1842 646.071
R8482 VPWR.n642 VPWR.t1030 646.071
R8483 VPWR.n646 VPWR.t186 646.071
R8484 VPWR.n650 VPWR.t996 646.071
R8485 VPWR.n654 VPWR.t1236 646.071
R8486 VPWR.n597 VPWR.t1740 646.071
R8487 VPWR.n684 VPWR.t1179 646.071
R8488 VPWR.n692 VPWR.t649 646.071
R8489 VPWR.n691 VPWR.t1158 646.071
R8490 VPWR.n688 VPWR.t1058 646.071
R8491 VPWR.n687 VPWR.t752 646.071
R8492 VPWR.n683 VPWR.t844 646.071
R8493 VPWR.n680 VPWR.t1906 646.071
R8494 VPWR.n679 VPWR.t241 646.071
R8495 VPWR.n676 VPWR.t801 646.071
R8496 VPWR.n675 VPWR.t353 646.071
R8497 VPWR.n672 VPWR.t1123 646.071
R8498 VPWR.n671 VPWR.t1810 646.071
R8499 VPWR.n668 VPWR.t1317 646.071
R8500 VPWR.n667 VPWR.t1196 646.071
R8501 VPWR.n664 VPWR.t826 646.071
R8502 VPWR.n663 VPWR.t1463 646.071
R8503 VPWR.n737 VPWR.t442 646.071
R8504 VPWR.n693 VPWR.t503 646.071
R8505 VPWR.n749 VPWR.t1921 646.071
R8506 VPWR.n745 VPWR.t1074 646.071
R8507 VPWR.n741 VPWR.t688 646.071
R8508 VPWR.n733 VPWR.t861 646.071
R8509 VPWR.n729 VPWR.t457 646.071
R8510 VPWR.n725 VPWR.t1928 646.071
R8511 VPWR.n721 VPWR.t656 646.071
R8512 VPWR.n717 VPWR.t339 646.071
R8513 VPWR.n713 VPWR.t1204 646.071
R8514 VPWR.n709 VPWR.t1018 646.071
R8515 VPWR.n705 VPWR.t1301 646.071
R8516 VPWR.n701 VPWR.t1010 646.071
R8517 VPWR.n697 VPWR.t1246 646.071
R8518 VPWR.n694 VPWR.t1570 646.071
R8519 VPWR.n767 VPWR.t448 646.071
R8520 VPWR.n759 VPWR.t647 646.071
R8521 VPWR.n760 VPWR.t509 646.071
R8522 VPWR.n763 VPWR.t1066 646.071
R8523 VPWR.n764 VPWR.t5 646.071
R8524 VPWR.n768 VPWR.t1098 646.071
R8525 VPWR.n771 VPWR.t463 646.071
R8526 VPWR.n772 VPWR.t544 646.071
R8527 VPWR.n775 VPWR.t565 646.071
R8528 VPWR.n776 VPWR.t345 646.071
R8529 VPWR.n779 VPWR.t1408 646.071
R8530 VPWR.n780 VPWR.t1162 646.071
R8531 VPWR.n783 VPWR.t1307 646.071
R8532 VPWR.n784 VPWR.t998 646.071
R8533 VPWR.n787 VPWR.t1252 646.071
R8534 VPWR.n788 VPWR.t1530 646.071
R8535 VPWR.n806 VPWR.t149 646.071
R8536 VPWR.n790 VPWR.t290 646.071
R8537 VPWR.n794 VPWR.t513 646.071
R8538 VPWR.n798 VPWR.t1086 646.071
R8539 VPWR.n802 VPWR.t412 646.071
R8540 VPWR.n810 VPWR.t57 646.071
R8541 VPWR.n814 VPWR.t719 646.071
R8542 VPWR.n818 VPWR.t231 646.071
R8543 VPWR.n822 VPWR.t523 646.071
R8544 VPWR.n826 VPWR.t329 646.071
R8545 VPWR.n830 VPWR.t551 646.071
R8546 VPWR.n834 VPWR.t1862 646.071
R8547 VPWR.n838 VPWR.t249 646.071
R8548 VPWR.n842 VPWR.t639 646.071
R8549 VPWR.n846 VPWR.t27 646.071
R8550 VPWR.n789 VPWR.t1635 646.071
R8551 VPWR.n876 VPWR.t1181 646.071
R8552 VPWR.n884 VPWR.t836 646.071
R8553 VPWR.n883 VPWR.t1160 646.071
R8554 VPWR.n880 VPWR.t1056 646.071
R8555 VPWR.n879 VPWR.t756 646.071
R8556 VPWR.n875 VPWR.t846 646.071
R8557 VPWR.n872 VPWR.t1908 646.071
R8558 VPWR.n871 VPWR.t243 646.071
R8559 VPWR.n868 VPWR.t803 646.071
R8560 VPWR.n867 VPWR.t382 646.071
R8561 VPWR.n864 VPWR.t1125 646.071
R8562 VPWR.n863 VPWR.t1812 646.071
R8563 VPWR.n860 VPWR.t398 646.071
R8564 VPWR.n859 VPWR.t1198 646.071
R8565 VPWR.n856 VPWR.t830 646.071
R8566 VPWR.n855 VPWR.t1455 646.071
R8567 VPWR.n929 VPWR.t147 646.071
R8568 VPWR.n885 VPWR.t288 646.071
R8569 VPWR.n941 VPWR.t511 646.071
R8570 VPWR.n937 VPWR.t1088 646.071
R8571 VPWR.n933 VPWR.t410 646.071
R8572 VPWR.n925 VPWR.t55 646.071
R8573 VPWR.n921 VPWR.t717 646.071
R8574 VPWR.n917 VPWR.t229 646.071
R8575 VPWR.n913 VPWR.t521 646.071
R8576 VPWR.n909 VPWR.t327 646.071
R8577 VPWR.n905 VPWR.t549 646.071
R8578 VPWR.n901 VPWR.t1860 646.071
R8579 VPWR.n897 VPWR.t247 646.071
R8580 VPWR.n893 VPWR.t637 646.071
R8581 VPWR.n889 VPWR.t25 646.071
R8582 VPWR.n886 VPWR.t1642 646.071
R8583 VPWR.n959 VPWR.t908 646.071
R8584 VPWR.n998 VPWR.t1260 646.071
R8585 VPWR.n1246 VPWR.t1148 646.071
R8586 VPWR.n1198 VPWR.t1474 646.071
R8587 VPWR.n418 VPWR.t758 646.071
R8588 VPWR.n380 VPWR.t1397 646.071
R8589 VPWR.n357 VPWR.t674 646.071
R8590 VPWR.n111 VPWR.t1482 646.071
R8591 VPWR.n994 VPWR.t416 646.071
R8592 VPWR.n1504 VPWR.t1401 646.071
R8593 VPWR.n1202 VPWR.t1756 646.071
R8594 VPWR.n960 VPWR.t1828 646.071
R8595 VPWR.n1002 VPWR.t63 646.071
R8596 VPWR.n1192 VPWR.t1804 646.071
R8597 VPWR.n1236 VPWR.t1621 646.071
R8598 VPWR.n434 VPWR.t233 646.071
R8599 VPWR.n438 VPWR.t157 646.071
R8600 VPWR.n442 VPWR.t384 646.071
R8601 VPWR.n446 VPWR.t1127 646.071
R8602 VPWR.n450 VPWR.t1814 646.071
R8603 VPWR.n454 VPWR.t400 646.071
R8604 VPWR.n458 VPWR.t1200 646.071
R8605 VPWR.n462 VPWR.t832 646.071
R8606 VPWR.n405 VPWR.t1447 646.071
R8607 VPWR.n387 VPWR.t1393 646.071
R8608 VPWR.n345 VPWR.t1383 646.071
R8609 VPWR.n100 VPWR.t1469 646.071
R8610 VPWR.n1006 VPWR.t725 646.071
R8611 VPWR.n1188 VPWR.t1395 646.071
R8612 VPWR.n1233 VPWR.t1732 646.071
R8613 VPWR.n967 VPWR.t1286 646.071
R8614 VPWR.n968 VPWR.t363 646.071
R8615 VPWR.n971 VPWR.t1840 646.071
R8616 VPWR.n972 VPWR.t1028 646.071
R8617 VPWR.n975 VPWR.t182 646.071
R8618 VPWR.n976 VPWR.t994 646.071
R8619 VPWR.n979 VPWR.t1232 646.071
R8620 VPWR.n980 VPWR.t1750 646.071
R8621 VPWR.n1010 VPWR.t221 646.071
R8622 VPWR.n1182 VPWR.t949 646.071
R8623 VPWR.n1225 VPWR.t1769 646.071
R8624 VPWR.n379 VPWR.t1036 646.071
R8625 VPWR.n361 VPWR.t1044 646.071
R8626 VPWR.n112 VPWR.t1700 646.071
R8627 VPWR.n1498 VPWR.t1092 646.071
R8628 VPWR.n1199 VPWR.t1593 646.071
R8629 VPWR.n1014 VPWR.t529 646.071
R8630 VPWR.n1178 VPWR.t298 646.071
R8631 VPWR.n1222 VPWR.t1514 646.071
R8632 VPWR.n395 VPWR.t1844 646.071
R8633 VPWR.n396 VPWR.t1885 646.071
R8634 VPWR.n399 VPWR.t188 646.071
R8635 VPWR.n400 VPWR.t980 646.071
R8636 VPWR.n403 VPWR.t1238 646.071
R8637 VPWR.n404 VPWR.t1735 646.071
R8638 VPWR.n333 VPWR.t361 646.071
R8639 VPWR.n93 VPWR.t1697 646.071
R8640 VPWR.n1168 VPWR.t369 646.071
R8641 VPWR.n1219 VPWR.t1618 646.071
R8642 VPWR.n1022 VPWR.t557 646.071
R8643 VPWR.n1026 VPWR.t1016 646.071
R8644 VPWR.n1030 VPWR.t253 646.071
R8645 VPWR.n1034 VPWR.t1008 646.071
R8646 VPWR.n1038 VPWR.t15 646.071
R8647 VPWR.n981 VPWR.t1602 646.071
R8648 VPWR.n1491 VPWR.t1337 646.071
R8649 VPWR.n1142 VPWR.t1580 646.071
R8650 VPWR.n329 VPWR.t485 646.071
R8651 VPWR.n88 VPWR.t1509 646.071
R8652 VPWR.n1211 VPWR.t1777 646.071
R8653 VPWR.n1068 VPWR.t1887 646.071
R8654 VPWR.n1208 VPWR.t1796 646.071
R8655 VPWR.n321 VPWR.t178 646.071
R8656 VPWR.n313 VPWR.t1226 646.071
R8657 VPWR.n310 VPWR.t1772 646.071
R8658 VPWR.n1077 VPWR.t1672 646.071
R8659 VPWR.n1767 VPWR.t982 646.071
R8660 VPWR.n1055 VPWR.t1242 646.071
R8661 VPWR.n1051 VPWR.t1719 646.071
R8662 VPWR.n1205 VPWR.t1540 646.071
R8663 VPWR.n82 VPWR.t1655 646.071
R8664 VPWR.n76 VPWR.t1428 646.071
R8665 VPWR.n1249 VPWR.t1522 642.13
R8666 VPWR.n1171 VPWR.t1450 642.13
R8667 VPWR.n1245 VPWR.t1658 642.13
R8668 VPWR.n1503 VPWR.t1556 642.13
R8669 VPWR.n1191 VPWR.t1683 642.13
R8670 VPWR.n1187 VPWR.t1431 642.13
R8671 VPWR.n1181 VPWR.t1553 642.13
R8672 VPWR.n1497 VPWR.t1785 642.13
R8673 VPWR.n1177 VPWR.t1694 642.13
R8674 VPWR.n1167 VPWR.t1716 642.13
R8675 VPWR.n1490 VPWR.t1675 642.13
R8676 VPWR.n1067 VPWR.t1583 642.13
R8677 VPWR.n1766 VPWR.t1460 642.13
R8678 VPWR.n1054 VPWR.t1497 642.13
R8679 VPWR.n1050 VPWR.t1605 642.13
R8680 VPWR.n1071 VPWR.t1624 642.13
R8681 VPWR.n2328 VPWR.t644 629.652
R8682 VPWR.n2329 VPWR.t504 629.652
R8683 VPWR.n2338 VPWR.t1071 629.652
R8684 VPWR.n2339 VPWR.t691 629.652
R8685 VPWR.n2348 VPWR.t443 629.652
R8686 VPWR.n2349 VPWR.t862 629.652
R8687 VPWR.n2358 VPWR.t458 629.652
R8688 VPWR.n2359 VPWR.t1929 629.652
R8689 VPWR.n2368 VPWR.t560 629.652
R8690 VPWR.n2369 VPWR.t342 629.652
R8691 VPWR.n2378 VPWR.t1205 629.652
R8692 VPWR.n2379 VPWR.t1021 629.652
R8693 VPWR.n2388 VPWR.t1302 629.652
R8694 VPWR.n2389 VPWR.t1013 629.652
R8695 VPWR.n2398 VPWR.t1249 629.652
R8696 VPWR.n561 VPWR.t786 629.652
R8697 VPWR.t1273 VPWR.n560 629.652
R8698 VPWR.t1045 VPWR.n556 629.652
R8699 VPWR.t671 VPWR.n552 629.652
R8700 VPWR.t897 VPWR.n548 629.652
R8701 VPWR.t1817 VPWR.n544 629.652
R8702 VPWR.t1378 VPWR.n540 629.652
R8703 VPWR.t608 VPWR.n536 629.652
R8704 VPWR.t669 VPWR.n532 629.652
R8705 VPWR.t358 VPWR.n528 629.652
R8706 VPWR.t480 VPWR.n524 629.652
R8707 VPWR.t1023 VPWR.n520 629.652
R8708 VPWR.t974 VPWR.n516 629.652
R8709 VPWR.t989 VPWR.n512 629.652
R8710 VPWR.t1223 VPWR.n508 629.652
R8711 VPWR.n2300 VPWR.t291 629.652
R8712 VPWR.t516 VPWR.n2299 629.652
R8713 VPWR.n2290 VPWR.t1083 629.652
R8714 VPWR.t413 VPWR.n2289 629.652
R8715 VPWR.n2280 VPWR.t152 629.652
R8716 VPWR.t60 VPWR.n2279 629.652
R8717 VPWR.n2270 VPWR.t722 629.652
R8718 VPWR.t218 VPWR.n2269 629.652
R8719 VPWR.n2260 VPWR.t526 629.652
R8720 VPWR.t330 VPWR.n2259 629.652
R8721 VPWR.n2250 VPWR.t554 629.652
R8722 VPWR.t1863 VPWR.n2249 629.652
R8723 VPWR.n2240 VPWR.t250 629.652
R8724 VPWR.t640 VPWR.n2239 629.652
R8725 VPWR.n2230 VPWR.t12 629.652
R8726 VPWR.n601 VPWR.t792 629.652
R8727 VPWR.n605 VPWR.t909 629.652
R8728 VPWR.n609 VPWR.t1037 629.652
R8729 VPWR.n613 VPWR.t683 629.652
R8730 VPWR.n617 VPWR.t1143 629.652
R8731 VPWR.n621 VPWR.t1799 629.652
R8732 VPWR.n625 VPWR.t1390 629.652
R8733 VPWR.n629 VPWR.t936 629.652
R8734 VPWR.n633 VPWR.t1287 629.652
R8735 VPWR.n637 VPWR.t364 629.652
R8736 VPWR.n641 VPWR.t1841 629.652
R8737 VPWR.n645 VPWR.t1029 629.652
R8738 VPWR.n649 VPWR.t185 629.652
R8739 VPWR.n653 VPWR.t995 629.652
R8740 VPWR.n657 VPWR.t1235 629.652
R8741 VPWR.n2132 VPWR.t648 629.652
R8742 VPWR.n2133 VPWR.t1157 629.652
R8743 VPWR.n2142 VPWR.t1057 629.652
R8744 VPWR.n2143 VPWR.t751 629.652
R8745 VPWR.n2152 VPWR.t1178 629.652
R8746 VPWR.n2153 VPWR.t843 629.652
R8747 VPWR.n2162 VPWR.t1905 629.652
R8748 VPWR.n2163 VPWR.t240 629.652
R8749 VPWR.n2172 VPWR.t800 629.652
R8750 VPWR.n2173 VPWR.t352 629.652
R8751 VPWR.n2182 VPWR.t1122 629.652
R8752 VPWR.n2183 VPWR.t1809 629.652
R8753 VPWR.n2192 VPWR.t1316 629.652
R8754 VPWR.n2193 VPWR.t1195 629.652
R8755 VPWR.n2202 VPWR.t825 629.652
R8756 VPWR.n753 VPWR.t502 629.652
R8757 VPWR.t1920 VPWR.n752 629.652
R8758 VPWR.t1073 VPWR.n748 629.652
R8759 VPWR.t687 VPWR.n744 629.652
R8760 VPWR.t441 VPWR.n740 629.652
R8761 VPWR.t860 VPWR.n736 629.652
R8762 VPWR.t456 VPWR.n732 629.652
R8763 VPWR.t1927 VPWR.n728 629.652
R8764 VPWR.t655 VPWR.n724 629.652
R8765 VPWR.t338 VPWR.n720 629.652
R8766 VPWR.t1203 VPWR.n716 629.652
R8767 VPWR.t1017 VPWR.n712 629.652
R8768 VPWR.t1300 VPWR.n708 629.652
R8769 VPWR.t1009 VPWR.n704 629.652
R8770 VPWR.t1245 VPWR.n700 629.652
R8771 VPWR.n2104 VPWR.t646 629.652
R8772 VPWR.t508 VPWR.n2103 629.652
R8773 VPWR.n2094 VPWR.t1065 629.652
R8774 VPWR.t4 VPWR.n2093 629.652
R8775 VPWR.n2084 VPWR.t447 629.652
R8776 VPWR.t1097 VPWR.n2083 629.652
R8777 VPWR.n2074 VPWR.t462 629.652
R8778 VPWR.t543 VPWR.n2073 629.652
R8779 VPWR.n2064 VPWR.t564 629.652
R8780 VPWR.t344 VPWR.n2063 629.652
R8781 VPWR.n2054 VPWR.t1407 629.652
R8782 VPWR.t1161 VPWR.n2053 629.652
R8783 VPWR.n2044 VPWR.t1306 629.652
R8784 VPWR.t997 VPWR.n2043 629.652
R8785 VPWR.n2034 VPWR.t1251 629.652
R8786 VPWR.n793 VPWR.t289 629.652
R8787 VPWR.n797 VPWR.t512 629.652
R8788 VPWR.n801 VPWR.t1085 629.652
R8789 VPWR.n805 VPWR.t411 629.652
R8790 VPWR.n809 VPWR.t148 629.652
R8791 VPWR.n813 VPWR.t56 629.652
R8792 VPWR.n817 VPWR.t718 629.652
R8793 VPWR.n821 VPWR.t230 629.652
R8794 VPWR.n825 VPWR.t522 629.652
R8795 VPWR.n829 VPWR.t328 629.652
R8796 VPWR.n833 VPWR.t550 629.652
R8797 VPWR.n837 VPWR.t1861 629.652
R8798 VPWR.n841 VPWR.t248 629.652
R8799 VPWR.n845 VPWR.t638 629.652
R8800 VPWR.n849 VPWR.t26 629.652
R8801 VPWR.n1936 VPWR.t835 629.652
R8802 VPWR.n1937 VPWR.t1159 629.652
R8803 VPWR.n1946 VPWR.t1055 629.652
R8804 VPWR.n1947 VPWR.t755 629.652
R8805 VPWR.n1956 VPWR.t1180 629.652
R8806 VPWR.n1957 VPWR.t845 629.652
R8807 VPWR.n1966 VPWR.t1907 629.652
R8808 VPWR.n1967 VPWR.t242 629.652
R8809 VPWR.n1976 VPWR.t802 629.652
R8810 VPWR.n1977 VPWR.t381 629.652
R8811 VPWR.n1986 VPWR.t1124 629.652
R8812 VPWR.n1987 VPWR.t1811 629.652
R8813 VPWR.n1996 VPWR.t397 629.652
R8814 VPWR.n1997 VPWR.t1197 629.652
R8815 VPWR.n2006 VPWR.t829 629.652
R8816 VPWR.n945 VPWR.t287 629.652
R8817 VPWR.t510 VPWR.n944 629.652
R8818 VPWR.t1087 VPWR.n940 629.652
R8819 VPWR.t409 VPWR.n936 629.652
R8820 VPWR.t146 VPWR.n932 629.652
R8821 VPWR.t54 VPWR.n928 629.652
R8822 VPWR.t716 VPWR.n924 629.652
R8823 VPWR.t228 VPWR.n920 629.652
R8824 VPWR.t520 VPWR.n916 629.652
R8825 VPWR.t326 VPWR.n912 629.652
R8826 VPWR.t548 VPWR.n908 629.652
R8827 VPWR.t1859 VPWR.n904 629.652
R8828 VPWR.t246 VPWR.n900 629.652
R8829 VPWR.t636 VPWR.n896 629.652
R8830 VPWR.t24 VPWR.n892 629.652
R8831 VPWR.n409 VPWR.t837 629.652
R8832 VPWR.n413 VPWR.t708 629.652
R8833 VPWR.n417 VPWR.t1053 629.652
R8834 VPWR.n421 VPWR.t757 629.652
R8835 VPWR.n425 VPWR.t1182 629.652
R8836 VPWR.n429 VPWR.t847 629.652
R8837 VPWR.n433 VPWR.t1909 629.652
R8838 VPWR.n437 VPWR.t232 629.652
R8839 VPWR.n441 VPWR.t156 629.652
R8840 VPWR.n445 VPWR.t383 629.652
R8841 VPWR.n449 VPWR.t1126 629.652
R8842 VPWR.n453 VPWR.t1813 629.652
R8843 VPWR.n457 VPWR.t399 629.652
R8844 VPWR.n461 VPWR.t1199 629.652
R8845 VPWR.n465 VPWR.t831 629.652
R8846 VPWR.n1908 VPWR.t790 629.652
R8847 VPWR.t1118 VPWR.n1907 629.652
R8848 VPWR.n1898 VPWR.t1039 629.652
R8849 VPWR.t679 VPWR.n1897 629.652
R8850 VPWR.n1888 VPWR.t907 629.652
R8851 VPWR.t1827 VPWR.n1887 629.652
R8852 VPWR.n1878 VPWR.t1388 629.652
R8853 VPWR.t932 VPWR.n1877 629.652
R8854 VPWR.n1868 VPWR.t1285 629.652
R8855 VPWR.t362 VPWR.n1867 629.652
R8856 VPWR.n1858 VPWR.t1839 629.652
R8857 VPWR.t1027 VPWR.n1857 629.652
R8858 VPWR.n1848 VPWR.t181 629.652
R8859 VPWR.t993 VPWR.n1847 629.652
R8860 VPWR.n1838 VPWR.t1231 629.652
R8861 VPWR.n2496 VPWR.t661 629.652
R8862 VPWR.t1334 VPWR.n2495 629.652
R8863 VPWR.n2486 VPWR.t1035 629.652
R8864 VPWR.t1396 VPWR.n2485 629.652
R8865 VPWR.n2476 VPWR.t1145 629.652
R8866 VPWR.t1801 VPWR.n2475 629.652
R8867 VPWR.n2466 VPWR.t1392 629.652
R8868 VPWR.t938 VPWR.n2465 629.652
R8869 VPWR.n2456 VPWR.t295 629.652
R8870 VPWR.t366 VPWR.n2455 629.652
R8871 VPWR.n2446 VPWR.t1843 629.652
R8872 VPWR.t1884 VPWR.n2445 629.652
R8873 VPWR.n2436 VPWR.t187 629.652
R8874 VPWR.t979 VPWR.n2435 629.652
R8875 VPWR.n2426 VPWR.t1237 629.652
R8876 VPWR.n985 VPWR.t500 629.652
R8877 VPWR.n989 VPWR.t518 629.652
R8878 VPWR.n993 VPWR.t1075 629.652
R8879 VPWR.n997 VPWR.t415 629.652
R8880 VPWR.n1001 VPWR.t1259 629.652
R8881 VPWR.n1005 VPWR.t62 629.652
R8882 VPWR.n1009 VPWR.t724 629.652
R8883 VPWR.n1013 VPWR.t220 629.652
R8884 VPWR.n1017 VPWR.t528 629.652
R8885 VPWR.n1021 VPWR.t336 629.652
R8886 VPWR.n1025 VPWR.t556 629.652
R8887 VPWR.n1029 VPWR.t1015 629.652
R8888 VPWR.n1033 VPWR.t252 629.652
R8889 VPWR.n1037 VPWR.t1007 629.652
R8890 VPWR.n1041 VPWR.t14 629.652
R8891 VPWR.n369 VPWR.t788 629.652
R8892 VPWR.t1112 VPWR.n368 629.652
R8893 VPWR.t1043 VPWR.n364 629.652
R8894 VPWR.t673 VPWR.n360 629.652
R8895 VPWR.t901 VPWR.n356 629.652
R8896 VPWR.t1821 VPWR.n352 629.652
R8897 VPWR.t1382 VPWR.n348 629.652
R8898 VPWR.t612 VPWR.n344 629.652
R8899 VPWR.t1279 VPWR.n340 629.652
R8900 VPWR.t360 VPWR.n336 629.652
R8901 VPWR.t484 VPWR.n332 629.652
R8902 VPWR.t1025 VPWR.n328 629.652
R8903 VPWR.t177 VPWR.n324 629.652
R8904 VPWR.t991 VPWR.n320 629.652
R8905 VPWR.t1225 VPWR.n316 629.652
R8906 VPWR.n1487 VPWR.t663 629.652
R8907 VPWR.n1494 VPWR.t1336 629.652
R8908 VPWR.n1500 VPWR.t1091 629.652
R8909 VPWR.n1511 VPWR.t1400 629.652
R8910 VPWR.n1512 VPWR.t1147 629.652
R8911 VPWR.n1525 VPWR.t1803 629.652
R8912 VPWR.n1526 VPWR.t1394 629.652
R8913 VPWR.n1539 VPWR.t948 629.652
R8914 VPWR.n1540 VPWR.t297 629.652
R8915 VPWR.n1555 VPWR.t368 629.652
R8916 VPWR.t1845 VPWR.n1554 629.652
R8917 VPWR.n1780 VPWR.t1886 629.652
R8918 VPWR.t189 VPWR.n1779 629.652
R8919 VPWR.n1768 VPWR.t981 629.652
R8920 VPWR.n1810 VPWR.t1241 629.652
R8921 VPWR.n2525 VPWR.t1572 629.652
R8922 VPWR.n2526 VPWR.t1707 629.652
R8923 VPWR.n2537 VPWR.t1699 629.652
R8924 VPWR.n2538 VPWR.t1481 629.652
R8925 VPWR.n2549 VPWR.t1589 629.652
R8926 VPWR.n2550 VPWR.t1744 629.652
R8927 VPWR.n2561 VPWR.t1468 629.652
R8928 VPWR.n2562 VPWR.t1503 629.652
R8929 VPWR.n2573 VPWR.t1631 629.652
R8930 VPWR.n2574 VPWR.t1696 629.652
R8931 VPWR.n2585 VPWR.t1508 629.652
R8932 VPWR.n2586 VPWR.t1526 629.652
R8933 VPWR.n2597 VPWR.t1654 629.652
R8934 VPWR.n2598 VPWR.t1787 629.652
R8935 VPWR.n2609 VPWR.t1427 629.652
R8936 VPWR.n1613 VPWR.t1443 629.652
R8937 VPWR.t1579 VPWR.n1612 629.652
R8938 VPWR.n1201 VPWR.t1592 629.652
R8939 VPWR.n1204 VPWR.t1755 629.652
R8940 VPWR.n1239 VPWR.t1473 629.652
R8941 VPWR.t1620 VPWR.n1238 629.652
R8942 VPWR.t1731 VPWR.n1235 629.652
R8943 VPWR.t1768 VPWR.n1232 629.652
R8944 VPWR.t1513 VPWR.n1224 629.652
R8945 VPWR.t1617 VPWR.n1221 629.652
R8946 VPWR.t1776 VPWR.n1218 629.652
R8947 VPWR.t1795 VPWR.n1210 629.652
R8948 VPWR.t1539 VPWR.n1207 629.652
R8949 VPWR.n1759 VPWR.t1671 629.652
R8950 VPWR.t1702 VPWR.n1758 629.652
R8951 VPWR.t644 VPWR.t138 486.048
R8952 VPWR.t504 VPWR.t1321 486.048
R8953 VPWR.t770 VPWR.t1071 486.048
R8954 VPWR.t691 VPWR.t141 486.048
R8955 VPWR.t1838 VPWR.t443 486.048
R8956 VPWR.t862 VPWR.t775 486.048
R8957 VPWR.t774 VPWR.t458 486.048
R8958 VPWR.t1929 VPWR.t1837 486.048
R8959 VPWR.t650 VPWR.t560 486.048
R8960 VPWR.t342 VPWR.t1320 486.048
R8961 VPWR.t140 VPWR.t1205 486.048
R8962 VPWR.t1021 VPWR.t139 486.048
R8963 VPWR.t773 VPWR.t1302 486.048
R8964 VPWR.t1013 VPWR.t772 486.048
R8965 VPWR.t771 VPWR.t1249 486.048
R8966 VPWR.t1561 VPWR.t1322 486.048
R8967 VPWR.t786 VPWR.t1879 486.048
R8968 VPWR.t1220 VPWR.t1273 486.048
R8969 VPWR.t852 VPWR.t1045 486.048
R8970 VPWR.t851 VPWR.t671 486.048
R8971 VPWR.t1878 VPWR.t897 486.048
R8972 VPWR.t1332 VPWR.t1817 486.048
R8973 VPWR.t1331 VPWR.t1378 486.048
R8974 VPWR.t1877 VPWR.t608 486.048
R8975 VPWR.t1222 VPWR.t669 486.048
R8976 VPWR.t1333 VPWR.t358 486.048
R8977 VPWR.t1881 VPWR.t480 486.048
R8978 VPWR.t1880 VPWR.t1023 486.048
R8979 VPWR.t1330 VPWR.t974 486.048
R8980 VPWR.t1329 VPWR.t989 486.048
R8981 VPWR.t853 VPWR.t1223 486.048
R8982 VPWR.t1221 VPWR.t1779 486.048
R8983 VPWR.t291 VPWR.t1353 486.048
R8984 VPWR.t1345 VPWR.t516 486.048
R8985 VPWR.t1083 VPWR.t1338 486.048
R8986 VPWR.t868 VPWR.t413 486.048
R8987 VPWR.t152 VPWR.t1352 486.048
R8988 VPWR.t1343 VPWR.t60 486.048
R8989 VPWR.t722 VPWR.t1342 486.048
R8990 VPWR.t1351 VPWR.t218 486.048
R8991 VPWR.t526 VPWR.t1350 486.048
R8992 VPWR.t1344 VPWR.t330 486.048
R8993 VPWR.t554 VPWR.t867 486.048
R8994 VPWR.t866 VPWR.t1863 486.048
R8995 VPWR.t250 VPWR.t1341 486.048
R8996 VPWR.t1340 VPWR.t640 486.048
R8997 VPWR.t12 VPWR.t1339 486.048
R8998 VPWR.t1349 VPWR.t1628 486.048
R8999 VPWR.t792 VPWR.t303 486.048
R9000 VPWR.t909 VPWR.t437 486.048
R9001 VPWR.t1037 VPWR.t440 486.048
R9002 VPWR.t683 VPWR.t439 486.048
R9003 VPWR.t1143 VPWR.t302 486.048
R9004 VPWR.t1799 VPWR.t435 486.048
R9005 VPWR.t1390 VPWR.t434 486.048
R9006 VPWR.t936 VPWR.t301 486.048
R9007 VPWR.t1287 VPWR.t300 486.048
R9008 VPWR.t364 VPWR.t436 486.048
R9009 VPWR.t1841 VPWR.t305 486.048
R9010 VPWR.t1029 VPWR.t304 486.048
R9011 VPWR.t185 VPWR.t433 486.048
R9012 VPWR.t995 VPWR.t432 486.048
R9013 VPWR.t1235 VPWR.t431 486.048
R9014 VPWR.t1739 VPWR.t438 486.048
R9015 VPWR.t648 VPWR.t702 486.048
R9016 VPWR.t1157 VPWR.t1257 486.048
R9017 VPWR.t603 VPWR.t1057 486.048
R9018 VPWR.t751 VPWR.t497 486.048
R9019 VPWR.t701 VPWR.t1178 486.048
R9020 VPWR.t843 VPWR.t1141 486.048
R9021 VPWR.t1140 VPWR.t1905 486.048
R9022 VPWR.t240 VPWR.t700 486.048
R9023 VPWR.t699 VPWR.t800 486.048
R9024 VPWR.t352 VPWR.t1142 486.048
R9025 VPWR.t496 VPWR.t1122 486.048
R9026 VPWR.t1809 VPWR.t495 486.048
R9027 VPWR.t1139 VPWR.t1316 486.048
R9028 VPWR.t1195 VPWR.t1138 486.048
R9029 VPWR.t604 VPWR.t825 486.048
R9030 VPWR.t1462 VPWR.t1258 486.048
R9031 VPWR.t502 VPWR.t1265 486.048
R9032 VPWR.t1191 VPWR.t1920 486.048
R9033 VPWR.t1374 VPWR.t1073 486.048
R9034 VPWR.t1373 VPWR.t687 486.048
R9035 VPWR.t1150 VPWR.t441 486.048
R9036 VPWR.t872 VPWR.t860 486.048
R9037 VPWR.t871 VPWR.t456 486.048
R9038 VPWR.t1149 VPWR.t1927 486.048
R9039 VPWR.t547 VPWR.t655 486.048
R9040 VPWR.t873 VPWR.t338 486.048
R9041 VPWR.t1267 VPWR.t1203 486.048
R9042 VPWR.t1266 VPWR.t1017 486.048
R9043 VPWR.t870 VPWR.t1300 486.048
R9044 VPWR.t869 VPWR.t1009 486.048
R9045 VPWR.t1375 VPWR.t1245 486.048
R9046 VPWR.t1192 VPWR.t1569 486.048
R9047 VPWR.t646 VPWR.t808 486.048
R9048 VPWR.t1034 VPWR.t508 486.048
R9049 VPWR.t1065 VPWR.t968 486.048
R9050 VPWR.t967 VPWR.t4 486.048
R9051 VPWR.t447 VPWR.t807 486.048
R9052 VPWR.t1032 VPWR.t1097 486.048
R9053 VPWR.t462 VPWR.t1031 486.048
R9054 VPWR.t806 VPWR.t543 486.048
R9055 VPWR.t564 VPWR.t805 486.048
R9056 VPWR.t1033 VPWR.t344 486.048
R9057 VPWR.t1407 VPWR.t966 486.048
R9058 VPWR.t965 VPWR.t1161 486.048
R9059 VPWR.t1306 VPWR.t971 486.048
R9060 VPWR.t970 VPWR.t997 486.048
R9061 VPWR.t1251 VPWR.t969 486.048
R9062 VPWR.t804 VPWR.t1529 486.048
R9063 VPWR.t289 VPWR.t396 486.048
R9064 VPWR.t512 VPWR.t391 486.048
R9065 VPWR.t1085 VPWR.t1849 486.048
R9066 VPWR.t411 VPWR.t1848 486.048
R9067 VPWR.t148 VPWR.t395 486.048
R9068 VPWR.t56 VPWR.t1854 486.048
R9069 VPWR.t718 VPWR.t1853 486.048
R9070 VPWR.t230 VPWR.t394 486.048
R9071 VPWR.t522 VPWR.t393 486.048
R9072 VPWR.t328 VPWR.t1855 486.048
R9073 VPWR.t550 VPWR.t1847 486.048
R9074 VPWR.t1861 VPWR.t321 486.048
R9075 VPWR.t248 VPWR.t1852 486.048
R9076 VPWR.t638 VPWR.t1851 486.048
R9077 VPWR.t26 VPWR.t1850 486.048
R9078 VPWR.t1634 VPWR.t392 486.048
R9079 VPWR.t835 VPWR.t538 486.048
R9080 VPWR.t1159 VPWR.t451 486.048
R9081 VPWR.t814 VPWR.t1055 486.048
R9082 VPWR.t755 VPWR.t813 486.048
R9083 VPWR.t537 VPWR.t1180 486.048
R9084 VPWR.t845 VPWR.t819 486.048
R9085 VPWR.t818 VPWR.t1907 486.048
R9086 VPWR.t242 VPWR.t536 486.048
R9087 VPWR.t535 VPWR.t802 486.048
R9088 VPWR.t381 VPWR.t820 486.048
R9089 VPWR.t540 VPWR.t1124 486.048
R9090 VPWR.t1811 VPWR.t539 486.048
R9091 VPWR.t817 VPWR.t397 486.048
R9092 VPWR.t1197 VPWR.t816 486.048
R9093 VPWR.t815 VPWR.t829 486.048
R9094 VPWR.t1454 VPWR.t534 486.048
R9095 VPWR.t287 VPWR.t217 486.048
R9096 VPWR.t212 VPWR.t510 486.048
R9097 VPWR.t954 VPWR.t1087 486.048
R9098 VPWR.t1915 VPWR.t409 486.048
R9099 VPWR.t216 VPWR.t146 486.048
R9100 VPWR.t959 VPWR.t54 486.048
R9101 VPWR.t958 VPWR.t716 486.048
R9102 VPWR.t215 VPWR.t228 486.048
R9103 VPWR.t214 VPWR.t520 486.048
R9104 VPWR.t960 VPWR.t326 486.048
R9105 VPWR.t1914 VPWR.t548 486.048
R9106 VPWR.t1913 VPWR.t1859 486.048
R9107 VPWR.t957 VPWR.t246 486.048
R9108 VPWR.t956 VPWR.t636 486.048
R9109 VPWR.t955 VPWR.t24 486.048
R9110 VPWR.t213 VPWR.t1641 486.048
R9111 VPWR.t837 VPWR.t923 486.048
R9112 VPWR.t708 VPWR.t1190 486.048
R9113 VPWR.t1053 VPWR.t706 486.048
R9114 VPWR.t757 VPWR.t705 486.048
R9115 VPWR.t1182 VPWR.t922 486.048
R9116 VPWR.t847 VPWR.t915 486.048
R9117 VPWR.t1909 VPWR.t914 486.048
R9118 VPWR.t232 VPWR.t921 486.048
R9119 VPWR.t156 VPWR.t920 486.048
R9120 VPWR.t383 VPWR.t916 486.048
R9121 VPWR.t1126 VPWR.t704 486.048
R9122 VPWR.t1813 VPWR.t703 486.048
R9123 VPWR.t399 VPWR.t913 486.048
R9124 VPWR.t1199 VPWR.t912 486.048
R9125 VPWR.t831 VPWR.t911 486.048
R9126 VPWR.t1446 VPWR.t919 486.048
R9127 VPWR.t790 VPWR.t1133 486.048
R9128 VPWR.t1355 VPWR.t1118 486.048
R9129 VPWR.t1039 VPWR.t1137 486.048
R9130 VPWR.t1136 VPWR.t679 486.048
R9131 VPWR.t907 VPWR.t1132 486.048
R9132 VPWR.t174 VPWR.t1827 486.048
R9133 VPWR.t1388 VPWR.t173 486.048
R9134 VPWR.t1358 VPWR.t932 486.048
R9135 VPWR.t1285 VPWR.t1357 486.048
R9136 VPWR.t1354 VPWR.t362 486.048
R9137 VPWR.t1839 VPWR.t1135 486.048
R9138 VPWR.t1134 VPWR.t1027 486.048
R9139 VPWR.t181 VPWR.t172 486.048
R9140 VPWR.t171 VPWR.t993 486.048
R9141 VPWR.t1231 VPWR.t170 486.048
R9142 VPWR.t1356 VPWR.t1749 486.048
R9143 VPWR.t661 VPWR.t1362 486.048
R9144 VPWR.t1364 VPWR.t1334 486.048
R9145 VPWR.t1035 VPWR.t883 486.048
R9146 VPWR.t1209 VPWR.t1396 486.048
R9147 VPWR.t1145 VPWR.t1361 486.048
R9148 VPWR.t888 VPWR.t1801 486.048
R9149 VPWR.t1392 VPWR.t887 486.048
R9150 VPWR.t1360 VPWR.t938 486.048
R9151 VPWR.t295 VPWR.t1359 486.048
R9152 VPWR.t1363 VPWR.t366 486.048
R9153 VPWR.t1843 VPWR.t1208 486.048
R9154 VPWR.t1207 VPWR.t1884 486.048
R9155 VPWR.t187 VPWR.t886 486.048
R9156 VPWR.t885 VPWR.t979 486.048
R9157 VPWR.t1237 VPWR.t884 486.048
R9158 VPWR.t1365 VPWR.t1734 486.048
R9159 VPWR.t500 VPWR.t1292 486.048
R9160 VPWR.t518 VPWR.t1289 486.048
R9161 VPWR.t1075 VPWR.t96 486.048
R9162 VPWR.t415 VPWR.t95 486.048
R9163 VPWR.t1259 VPWR.t492 486.048
R9164 VPWR.t62 VPWR.t1298 486.048
R9165 VPWR.t724 VPWR.t1297 486.048
R9166 VPWR.t220 VPWR.t491 486.048
R9167 VPWR.t528 VPWR.t1291 486.048
R9168 VPWR.t336 VPWR.t1299 486.048
R9169 VPWR.t556 VPWR.t94 486.048
R9170 VPWR.t1015 VPWR.t1293 486.048
R9171 VPWR.t252 VPWR.t1296 486.048
R9172 VPWR.t1007 VPWR.t1295 486.048
R9173 VPWR.t14 VPWR.t97 486.048
R9174 VPWR.t1601 VPWR.t1290 486.048
R9175 VPWR.t788 VPWR.t1218 486.048
R9176 VPWR.t746 VPWR.t1112 486.048
R9177 VPWR.t811 VPWR.t1043 486.048
R9178 VPWR.t810 VPWR.t673 486.048
R9179 VPWR.t1217 VPWR.t901 486.048
R9180 VPWR.t744 VPWR.t1821 486.048
R9181 VPWR.t743 VPWR.t1382 486.048
R9182 VPWR.t1216 VPWR.t612 486.048
R9183 VPWR.t1215 VPWR.t1279 486.048
R9184 VPWR.t745 VPWR.t360 486.048
R9185 VPWR.t809 VPWR.t484 486.048
R9186 VPWR.t1219 VPWR.t1025 486.048
R9187 VPWR.t742 VPWR.t177 486.048
R9188 VPWR.t741 VPWR.t991 486.048
R9189 VPWR.t812 VPWR.t1225 486.048
R9190 VPWR.t1214 VPWR.t1771 486.048
R9191 VPWR.t663 VPWR.t1506 486.048
R9192 VPWR.t1336 VPWR.t1637 486.048
R9193 VPWR.t1091 VPWR.t1766 486.048
R9194 VPWR.t1400 VPWR.t1422 486.048
R9195 VPWR.t1147 VPWR.t1532 486.048
R9196 VPWR.t1687 VPWR.t1803 486.048
R9197 VPWR.t1394 VPWR.t1689 486.048
R9198 VPWR.t1537 VPWR.t948 486.048
R9199 VPWR.t297 VPWR.t1567 486.048
R9200 VPWR.t1685 VPWR.t368 486.048
R9201 VPWR.t1436 VPWR.t1845 486.048
R9202 VPWR.t1452 VPWR.t1886 486.048
R9203 VPWR.t1705 VPWR.t189 486.048
R9204 VPWR.t981 VPWR.t1723 486.048
R9205 VPWR.t1758 VPWR.t1241 486.048
R9206 VPWR.t1718 VPWR.t1587 486.048
R9207 VPWR.t1572 VPWR.t1441 486.048
R9208 VPWR.t1707 VPWR.t1577 486.048
R9209 VPWR.t1713 VPWR.t1699 486.048
R9210 VPWR.t1481 VPWR.t1747 486.048
R9211 VPWR.t1471 VPWR.t1589 486.048
R9212 VPWR.t1744 VPWR.t1615 486.048
R9213 VPWR.t1639 VPWR.t1468 486.048
R9214 VPWR.t1503 VPWR.t1476 486.048
R9215 VPWR.t1511 VPWR.t1631 486.048
R9216 VPWR.t1696 VPWR.t1613 486.048
R9217 VPWR.t1774 VPWR.t1508 486.048
R9218 VPWR.t1526 VPWR.t1793 486.048
R9219 VPWR.t1647 VPWR.t1654 486.048
R9220 VPWR.t1787 VPWR.t1669 486.048
R9221 VPWR.t1691 VPWR.t1427 486.048
R9222 VPWR.t1663 VPWR.t1542 486.048
R9223 VPWR.t1443 VPWR.t1721 486.048
R9224 VPWR.t1457 VPWR.t1579 486.048
R9225 VPWR.t1592 VPWR.t1585 486.048
R9226 VPWR.t1755 VPWR.t1626 486.048
R9227 VPWR.t1473 VPWR.t1737 486.048
R9228 VPWR.t1501 VPWR.t1620 486.048
R9229 VPWR.t1516 VPWR.t1731 486.048
R9230 VPWR.t1742 VPWR.t1768 486.048
R9231 VPWR.t1782 VPWR.t1513 486.048
R9232 VPWR.t1499 VPWR.t1617 486.048
R9233 VPWR.t1652 VPWR.t1776 486.048
R9234 VPWR.t1677 VPWR.t1795 486.048
R9235 VPWR.t1524 VPWR.t1539 486.048
R9236 VPWR.t1550 VPWR.t1671 486.048
R9237 VPWR.t1575 VPWR.t1702 486.048
R9238 VPWR.t1547 VPWR.t1420 486.048
R9239 VPWR.t138 VPWR.t595 463.954
R9240 VPWR.t1321 VPWR.t498 463.954
R9241 VPWR.t1918 VPWR.t770 463.954
R9242 VPWR.t141 VPWR.t1093 463.954
R9243 VPWR.t405 VPWR.t1838 463.954
R9244 VPWR.t775 VPWR.t1263 463.954
R9245 VPWR.t858 VPWR.t774 463.954
R9246 VPWR.t1837 VPWR.t454 463.954
R9247 VPWR.t952 VPWR.t650 463.954
R9248 VPWR.t1320 VPWR.t653 463.954
R9249 VPWR.t334 VPWR.t140 463.954
R9250 VPWR.t139 VPWR.t1201 463.954
R9251 VPWR.t1867 VPWR.t773 463.954
R9252 VPWR.t772 VPWR.t193 463.954
R9253 VPWR.t1005 VPWR.t771 463.954
R9254 VPWR.t1322 VPWR.t20 463.954
R9255 VPWR.t1879 VPWR.t585 463.954
R9256 VPWR.t839 VPWR.t1220 463.954
R9257 VPWR.t1269 VPWR.t852 463.954
R9258 VPWR.t1069 VPWR.t851 463.954
R9259 VPWR.t6 VPWR.t1878 463.954
R9260 VPWR.t1210 VPWR.t1332 463.954
R9261 VPWR.t849 VPWR.t1331 463.954
R9262 VPWR.t1911 VPWR.t1877 463.954
R9263 VPWR.t541 VPWR.t1222 463.954
R9264 VPWR.t665 VPWR.t1333 463.954
R9265 VPWR.t385 VPWR.t1881 463.954
R9266 VPWR.t476 VPWR.t1880 463.954
R9267 VPWR.t66 VPWR.t1330 463.954
R9268 VPWR.t1304 VPWR.t1329 463.954
R9269 VPWR.t983 VPWR.t853 463.954
R9270 VPWR.t1253 VPWR.t1221 463.954
R9271 VPWR.t1353 VPWR.t571 463.954
R9272 VPWR.t735 VPWR.t1345 463.954
R9273 VPWR.t1338 VPWR.t1188 463.954
R9274 VPWR.t1047 VPWR.t868 463.954
R9275 VPWR.t1352 VPWR.t681 463.954
R9276 VPWR.t144 VPWR.t1343 463.954
R9277 VPWR.t1342 VPWR.t52 463.954
R9278 VPWR.t714 VPWR.t1351 463.954
R9279 VPWR.t1350 VPWR.t930 463.954
R9280 VPWR.t46 VPWR.t1344 463.954
R9281 VPWR.t867 VPWR.t322 463.954
R9282 VPWR.t780 VPWR.t866 463.954
R9283 VPWR.t1341 VPWR.t1873 463.954
R9284 VPWR.t179 VPWR.t1340 463.954
R9285 VPWR.t1339 VPWR.t530 463.954
R9286 VPWR.t1233 VPWR.t1349 463.954
R9287 VPWR.t303 VPWR.t579 463.954
R9288 VPWR.t437 VPWR.t782 463.954
R9289 VPWR.t440 VPWR.t1114 463.954
R9290 VPWR.t439 VPWR.t1061 463.954
R9291 VPWR.t302 VPWR.t749 463.954
R9292 VPWR.t435 VPWR.t903 463.954
R9293 VPWR.t434 VPWR.t1823 463.954
R9294 VPWR.t301 VPWR.t1384 463.954
R9295 VPWR.t300 VPWR.t236 463.954
R9296 VPWR.t436 VPWR.t1281 463.954
R9297 VPWR.t305 VPWR.t354 463.954
R9298 VPWR.t304 VPWR.t486 463.954
R9299 VPWR.t433 VPWR.t630 463.954
R9300 VPWR.t432 VPWR.t1312 463.954
R9301 VPWR.t431 VPWR.t601 463.954
R9302 VPWR.t438 VPWR.t823 463.954
R9303 VPWR.t702 VPWR.t591 463.954
R9304 VPWR.t1257 VPWR.t70 463.954
R9305 VPWR.t1151 VPWR.t603 463.954
R9306 VPWR.t497 VPWR.t1081 463.954
R9307 VPWR.t417 VPWR.t701 463.954
R9308 VPWR.t1141 VPWR.t1323 463.954
R9309 VPWR.t1099 VPWR.t1140 463.954
R9310 VPWR.t700 VPWR.t1899 463.954
R9311 VPWR.t222 VPWR.t699 463.954
R9312 VPWR.t1142 VPWR.t794 463.954
R9313 VPWR.t346 VPWR.t496 463.954
R9314 VPWR.t495 VPWR.t1409 463.954
R9315 VPWR.t1163 VPWR.t1139 463.954
R9316 VPWR.t1138 VPWR.t254 463.954
R9317 VPWR.t999 VPWR.t604 463.954
R9318 VPWR.t1258 VPWR.t16 463.954
R9319 VPWR.t1265 VPWR.t597 463.954
R9320 VPWR.t293 VPWR.t1191 463.954
R9321 VPWR.t1916 VPWR.t1374 463.954
R9322 VPWR.t1095 VPWR.t1373 463.954
R9323 VPWR.t1402 VPWR.t1150 463.954
R9324 VPWR.t1261 VPWR.t872 463.954
R9325 VPWR.t64 VPWR.t871 463.954
R9326 VPWR.t452 VPWR.t1149 463.954
R9327 VPWR.t950 VPWR.t547 463.954
R9328 VPWR.t651 VPWR.t873 463.954
R9329 VPWR.t332 VPWR.t1267 463.954
R9330 VPWR.t558 VPWR.t1266 463.954
R9331 VPWR.t1865 VPWR.t870 463.954
R9332 VPWR.t191 VPWR.t869 463.954
R9333 VPWR.t1003 VPWR.t1375 463.954
R9334 VPWR.t18 VPWR.t1192 463.954
R9335 VPWR.t808 VPWR.t593 463.954
R9336 VPWR.t642 VPWR.t1034 463.954
R9337 VPWR.t968 VPWR.t506 463.954
R9338 VPWR.t1089 VPWR.t967 463.954
R9339 VPWR.t807 VPWR.t407 463.954
R9340 VPWR.t445 VPWR.t1032 463.954
R9341 VPWR.t1031 VPWR.t864 463.954
R9342 VPWR.t460 VPWR.t806 463.954
R9343 VPWR.t805 VPWR.t226 463.954
R9344 VPWR.t562 VPWR.t1033 463.954
R9345 VPWR.t966 VPWR.t340 463.954
R9346 VPWR.t532 VPWR.t965 463.954
R9347 VPWR.t971 VPWR.t1019 463.954
R9348 VPWR.t244 VPWR.t970 463.954
R9349 VPWR.t969 VPWR.t1011 463.954
R9350 VPWR.t22 VPWR.t804 463.954
R9351 VPWR.t396 VPWR.t573 463.954
R9352 VPWR.t391 VPWR.t733 463.954
R9353 VPWR.t1849 VPWR.t1186 463.954
R9354 VPWR.t1848 VPWR.t1049 463.954
R9355 VPWR.t395 VPWR.t677 463.954
R9356 VPWR.t1854 VPWR.t142 463.954
R9357 VPWR.t1853 VPWR.t50 463.954
R9358 VPWR.t394 VPWR.t712 463.954
R9359 VPWR.t393 VPWR.t610 463.954
R9360 VPWR.t1855 VPWR.t44 463.954
R9361 VPWR.t1847 VPWR.t2 463.954
R9362 VPWR.t321 VPWR.t778 463.954
R9363 VPWR.t1852 VPWR.t1871 463.954
R9364 VPWR.t1851 VPWR.t976 463.954
R9365 VPWR.t1850 VPWR.t40 463.954
R9366 VPWR.t392 VPWR.t1229 463.954
R9367 VPWR.t538 VPWR.t589 463.954
R9368 VPWR.t451 VPWR.t72 463.954
R9369 VPWR.t1153 VPWR.t814 463.954
R9370 VPWR.t813 VPWR.t1079 463.954
R9371 VPWR.t685 VPWR.t537 463.954
R9372 VPWR.t819 VPWR.t1325 463.954
R9373 VPWR.t1101 VPWR.t818 463.954
R9374 VPWR.t536 VPWR.t1901 463.954
R9375 VPWR.t224 VPWR.t535 463.954
R9376 VPWR.t820 VPWR.t796 463.954
R9377 VPWR.t348 VPWR.t540 463.954
R9378 VPWR.t539 VPWR.t1411 463.954
R9379 VPWR.t1805 VPWR.t817 463.954
R9380 VPWR.t816 VPWR.t256 463.954
R9381 VPWR.t1001 VPWR.t815 463.954
R9382 VPWR.t534 VPWR.t1243 463.954
R9383 VPWR.t217 VPWR.t575 463.954
R9384 VPWR.t731 VPWR.t212 463.954
R9385 VPWR.t1184 VPWR.t954 463.954
R9386 VPWR.t1051 VPWR.t1915 463.954
R9387 VPWR.t675 VPWR.t216 463.954
R9388 VPWR.t928 VPWR.t959 463.954
R9389 VPWR.t48 VPWR.t958 463.954
R9390 VPWR.t710 VPWR.t215 463.954
R9391 VPWR.t606 VPWR.t214 463.954
R9392 VPWR.t42 VPWR.t960 463.954
R9393 VPWR.t0 VPWR.t1914 463.954
R9394 VPWR.t776 VPWR.t1913 463.954
R9395 VPWR.t1869 VPWR.t957 463.954
R9396 VPWR.t972 VPWR.t956 463.954
R9397 VPWR.t38 VPWR.t955 463.954
R9398 VPWR.t1227 VPWR.t213 463.954
R9399 VPWR.t923 VPWR.t587 463.954
R9400 VPWR.t1190 VPWR.t74 463.954
R9401 VPWR.t706 VPWR.t1155 463.954
R9402 VPWR.t705 VPWR.t1077 463.954
R9403 VPWR.t922 VPWR.t689 463.954
R9404 VPWR.t915 VPWR.t1327 463.954
R9405 VPWR.t914 VPWR.t1103 463.954
R9406 VPWR.t921 VPWR.t1903 463.954
R9407 VPWR.t920 VPWR.t1925 463.954
R9408 VPWR.t916 VPWR.t798 463.954
R9409 VPWR.t704 VPWR.t350 463.954
R9410 VPWR.t703 VPWR.t1120 463.954
R9411 VPWR.t913 VPWR.t1807 463.954
R9412 VPWR.t912 VPWR.t258 463.954
R9413 VPWR.t911 VPWR.t1193 463.954
R9414 VPWR.t919 VPWR.t1247 463.954
R9415 VPWR.t1133 VPWR.t581 463.954
R9416 VPWR.t1128 VPWR.t1355 463.954
R9417 VPWR.t1137 VPWR.t1275 463.954
R9418 VPWR.t1063 VPWR.t1136 463.954
R9419 VPWR.t1132 VPWR.t10 463.954
R9420 VPWR.t899 VPWR.t174 463.954
R9421 VPWR.t173 VPWR.t1819 463.954
R9422 VPWR.t1380 VPWR.t1358 463.954
R9423 VPWR.t1357 VPWR.t234 463.954
R9424 VPWR.t1277 VPWR.t1354 463.954
R9425 VPWR.t1135 VPWR.t389 463.954
R9426 VPWR.t482 VPWR.t1134 463.954
R9427 VPWR.t172 VPWR.t628 463.954
R9428 VPWR.t1310 VPWR.t171 463.954
R9429 VPWR.t170 VPWR.t599 463.954
R9430 VPWR.t821 VPWR.t1356 463.954
R9431 VPWR.t1362 VPWR.t577 463.954
R9432 VPWR.t784 VPWR.t1364 463.954
R9433 VPWR.t883 VPWR.t1116 463.954
R9434 VPWR.t1059 VPWR.t1209 463.954
R9435 VPWR.t1361 VPWR.t753 463.954
R9436 VPWR.t905 VPWR.t888 463.954
R9437 VPWR.t887 VPWR.t1825 463.954
R9438 VPWR.t1386 VPWR.t1360 463.954
R9439 VPWR.t1359 VPWR.t238 463.954
R9440 VPWR.t1283 VPWR.t1363 463.954
R9441 VPWR.t1208 VPWR.t356 463.954
R9442 VPWR.t488 VPWR.t1207 463.954
R9443 VPWR.t886 VPWR.t632 463.954
R9444 VPWR.t1314 VPWR.t885 463.954
R9445 VPWR.t884 VPWR.t987 463.954
R9446 VPWR.t827 VPWR.t1365 463.954
R9447 VPWR.t1292 VPWR.t566 463.954
R9448 VPWR.t1289 VPWR.t285 463.954
R9449 VPWR.t96 VPWR.t514 463.954
R9450 VPWR.t95 VPWR.t1041 463.954
R9451 VPWR.t492 VPWR.t1398 463.954
R9452 VPWR.t1298 VPWR.t150 463.954
R9453 VPWR.t1297 VPWR.t58 463.954
R9454 VPWR.t491 VPWR.t720 463.954
R9455 VPWR.t1291 VPWR.t934 463.954
R9456 VPWR.t1299 VPWR.t524 463.954
R9457 VPWR.t94 VPWR.t324 463.954
R9458 VPWR.t1293 VPWR.t552 463.954
R9459 VPWR.t1296 VPWR.t1875 463.954
R9460 VPWR.t1295 VPWR.t183 463.954
R9461 VPWR.t97 VPWR.t634 463.954
R9462 VPWR.t1290 VPWR.t1239 463.954
R9463 VPWR.t1218 VPWR.t583 463.954
R9464 VPWR.t841 VPWR.t746 463.954
R9465 VPWR.t1271 VPWR.t811 463.954
R9466 VPWR.t1067 VPWR.t810 463.954
R9467 VPWR.t8 VPWR.t1217 463.954
R9468 VPWR.t1212 VPWR.t744 463.954
R9469 VPWR.t1815 VPWR.t743 463.954
R9470 VPWR.t1376 VPWR.t1216 463.954
R9471 VPWR.t545 VPWR.t1215 463.954
R9472 VPWR.t667 VPWR.t745 463.954
R9473 VPWR.t387 VPWR.t809 463.954
R9474 VPWR.t478 VPWR.t1219 463.954
R9475 VPWR.t68 VPWR.t742 463.954
R9476 VPWR.t1308 VPWR.t741 463.954
R9477 VPWR.t985 VPWR.t812 463.954
R9478 VPWR.t1255 VPWR.t1214 463.954
R9479 VPWR.t1506 VPWR.t1521 463.954
R9480 VPWR.t1637 VPWR.t1674 463.954
R9481 VPWR.t1766 VPWR.t1784 463.954
R9482 VPWR.t1422 VPWR.t1555 463.954
R9483 VPWR.t1532 VPWR.t1657 463.954
R9484 VPWR.t1682 VPWR.t1687 463.954
R9485 VPWR.t1689 VPWR.t1430 463.954
R9486 VPWR.t1552 VPWR.t1537 463.954
R9487 VPWR.t1567 VPWR.t1693 463.954
R9488 VPWR.t1715 VPWR.t1685 463.954
R9489 VPWR.t1449 VPWR.t1436 463.954
R9490 VPWR.t1582 VPWR.t1452 463.954
R9491 VPWR.t1623 VPWR.t1705 463.954
R9492 VPWR.t1723 VPWR.t1459 463.954
R9493 VPWR.t1496 VPWR.t1758 463.954
R9494 VPWR.t1587 VPWR.t1604 463.954
R9495 VPWR.t1441 VPWR.t1465 463.954
R9496 VPWR.t1577 VPWR.t1610 463.954
R9497 VPWR.t1725 VPWR.t1713 463.954
R9498 VPWR.t1747 VPWR.t1487 463.954
R9499 VPWR.t1595 VPWR.t1471 463.954
R9500 VPWR.t1615 VPWR.t1607 463.954
R9501 VPWR.t1763 VPWR.t1639 463.954
R9502 VPWR.t1476 VPWR.t1484 463.954
R9503 VPWR.t1644 VPWR.t1511 463.954
R9504 VPWR.t1613 VPWR.t1660 463.954
R9505 VPWR.t1790 VPWR.t1774 463.954
R9506 VPWR.t1793 VPWR.t1534 463.954
R9507 VPWR.t1564 VPWR.t1647 463.954
R9508 VPWR.t1669 VPWR.t1414 463.954
R9509 VPWR.t1433 VPWR.t1691 463.954
R9510 VPWR.t1542 VPWR.t1558 463.954
R9511 VPWR.t1721 VPWR.t1728 463.954
R9512 VPWR.t1493 VPWR.t1457 463.954
R9513 VPWR.t1585 VPWR.t1598 463.954
R9514 VPWR.t1626 VPWR.t1760 463.954
R9515 VPWR.t1737 VPWR.t1478 463.954
R9516 VPWR.t1490 VPWR.t1501 463.954
R9517 VPWR.t1649 VPWR.t1516 463.954
R9518 VPWR.t1752 VPWR.t1742 463.954
R9519 VPWR.t1518 VPWR.t1782 463.954
R9520 VPWR.t1544 VPWR.t1499 463.954
R9521 VPWR.t1666 VPWR.t1652 463.954
R9522 VPWR.t1417 VPWR.t1677 463.954
R9523 VPWR.t1438 VPWR.t1524 463.954
R9524 VPWR.t1679 VPWR.t1550 463.954
R9525 VPWR.t1710 VPWR.t1575 463.954
R9526 VPWR.t1420 VPWR.t1424 463.954
R9527 VPWR.n2645 VPWR.t122 428.822
R9528 VPWR.t568 VPWR.n2835 376.524
R9529 VPWR.n1614 VPWR.n1613 376.045
R9530 VPWR.n2525 VPWR.n2524 376.045
R9531 VPWR.n1487 VPWR.n1486 376.045
R9532 VPWR.n370 VPWR.n369 376.045
R9533 VPWR.n2587 VPWR.n2586 376.045
R9534 VPWR.n1554 VPWR.n1553 376.045
R9535 VPWR.n368 VPWR.n367 376.045
R9536 VPWR.n2527 VPWR.n2526 376.045
R9537 VPWR.n985 VPWR.n984 376.045
R9538 VPWR.n2497 VPWR.n2496 376.045
R9539 VPWR.n2495 VPWR.n2494 376.045
R9540 VPWR.n340 VPWR.n339 376.045
R9541 VPWR.n2573 VPWR.n2572 376.045
R9542 VPWR.n993 VPWR.n992 376.045
R9543 VPWR.n2465 VPWR.n2464 376.045
R9544 VPWR.n344 VPWR.n343 376.045
R9545 VPWR.n2563 VPWR.n2562 376.045
R9546 VPWR.n1909 VPWR.n1908 376.045
R9547 VPWR.n1907 VPWR.n1906 376.045
R9548 VPWR.n1899 VPWR.n1898 376.045
R9549 VPWR.n409 VPWR.n408 376.045
R9550 VPWR.n413 VPWR.n412 376.045
R9551 VPWR.n417 VPWR.n416 376.045
R9552 VPWR.n2475 VPWR.n2474 376.045
R9553 VPWR.n352 VPWR.n351 376.045
R9554 VPWR.n2551 VPWR.n2550 376.045
R9555 VPWR.n1897 VPWR.n1896 376.045
R9556 VPWR.n425 VPWR.n424 376.045
R9557 VPWR.n2477 VPWR.n2476 376.045
R9558 VPWR.n356 VPWR.n355 376.045
R9559 VPWR.n2549 VPWR.n2548 376.045
R9560 VPWR.n2328 VPWR.n2327 376.045
R9561 VPWR.n2330 VPWR.n2329 376.045
R9562 VPWR.n2338 VPWR.n2337 376.045
R9563 VPWR.n2340 VPWR.n2339 376.045
R9564 VPWR.n2350 VPWR.n2349 376.045
R9565 VPWR.n2358 VPWR.n2357 376.045
R9566 VPWR.n2360 VPWR.n2359 376.045
R9567 VPWR.n2368 VPWR.n2367 376.045
R9568 VPWR.n2370 VPWR.n2369 376.045
R9569 VPWR.n2378 VPWR.n2377 376.045
R9570 VPWR.n2380 VPWR.n2379 376.045
R9571 VPWR.n2388 VPWR.n2387 376.045
R9572 VPWR.n2390 VPWR.n2389 376.045
R9573 VPWR.n2398 VPWR.n2397 376.045
R9574 VPWR.n2348 VPWR.n2347 376.045
R9575 VPWR.n562 VPWR.n561 376.045
R9576 VPWR.n560 VPWR.n559 376.045
R9577 VPWR.n556 VPWR.n555 376.045
R9578 VPWR.n552 VPWR.n551 376.045
R9579 VPWR.n544 VPWR.n543 376.045
R9580 VPWR.n540 VPWR.n539 376.045
R9581 VPWR.n536 VPWR.n535 376.045
R9582 VPWR.n532 VPWR.n531 376.045
R9583 VPWR.n528 VPWR.n527 376.045
R9584 VPWR.n524 VPWR.n523 376.045
R9585 VPWR.n520 VPWR.n519 376.045
R9586 VPWR.n516 VPWR.n515 376.045
R9587 VPWR.n512 VPWR.n511 376.045
R9588 VPWR.n508 VPWR.n507 376.045
R9589 VPWR.n548 VPWR.n547 376.045
R9590 VPWR.n2301 VPWR.n2300 376.045
R9591 VPWR.n2299 VPWR.n2298 376.045
R9592 VPWR.n2291 VPWR.n2290 376.045
R9593 VPWR.n2289 VPWR.n2288 376.045
R9594 VPWR.n2279 VPWR.n2278 376.045
R9595 VPWR.n2271 VPWR.n2270 376.045
R9596 VPWR.n2269 VPWR.n2268 376.045
R9597 VPWR.n2261 VPWR.n2260 376.045
R9598 VPWR.n2259 VPWR.n2258 376.045
R9599 VPWR.n2251 VPWR.n2250 376.045
R9600 VPWR.n2249 VPWR.n2248 376.045
R9601 VPWR.n2241 VPWR.n2240 376.045
R9602 VPWR.n2239 VPWR.n2238 376.045
R9603 VPWR.n2231 VPWR.n2230 376.045
R9604 VPWR.n2281 VPWR.n2280 376.045
R9605 VPWR.n601 VPWR.n600 376.045
R9606 VPWR.n605 VPWR.n604 376.045
R9607 VPWR.n609 VPWR.n608 376.045
R9608 VPWR.n613 VPWR.n612 376.045
R9609 VPWR.n621 VPWR.n620 376.045
R9610 VPWR.n625 VPWR.n624 376.045
R9611 VPWR.n629 VPWR.n628 376.045
R9612 VPWR.n633 VPWR.n632 376.045
R9613 VPWR.n637 VPWR.n636 376.045
R9614 VPWR.n641 VPWR.n640 376.045
R9615 VPWR.n645 VPWR.n644 376.045
R9616 VPWR.n649 VPWR.n648 376.045
R9617 VPWR.n653 VPWR.n652 376.045
R9618 VPWR.n657 VPWR.n656 376.045
R9619 VPWR.n617 VPWR.n616 376.045
R9620 VPWR.n2132 VPWR.n2131 376.045
R9621 VPWR.n2134 VPWR.n2133 376.045
R9622 VPWR.n2142 VPWR.n2141 376.045
R9623 VPWR.n2144 VPWR.n2143 376.045
R9624 VPWR.n2154 VPWR.n2153 376.045
R9625 VPWR.n2162 VPWR.n2161 376.045
R9626 VPWR.n2164 VPWR.n2163 376.045
R9627 VPWR.n2172 VPWR.n2171 376.045
R9628 VPWR.n2174 VPWR.n2173 376.045
R9629 VPWR.n2182 VPWR.n2181 376.045
R9630 VPWR.n2184 VPWR.n2183 376.045
R9631 VPWR.n2192 VPWR.n2191 376.045
R9632 VPWR.n2194 VPWR.n2193 376.045
R9633 VPWR.n2202 VPWR.n2201 376.045
R9634 VPWR.n2152 VPWR.n2151 376.045
R9635 VPWR.n754 VPWR.n753 376.045
R9636 VPWR.n752 VPWR.n751 376.045
R9637 VPWR.n748 VPWR.n747 376.045
R9638 VPWR.n744 VPWR.n743 376.045
R9639 VPWR.n736 VPWR.n735 376.045
R9640 VPWR.n732 VPWR.n731 376.045
R9641 VPWR.n728 VPWR.n727 376.045
R9642 VPWR.n724 VPWR.n723 376.045
R9643 VPWR.n720 VPWR.n719 376.045
R9644 VPWR.n716 VPWR.n715 376.045
R9645 VPWR.n712 VPWR.n711 376.045
R9646 VPWR.n708 VPWR.n707 376.045
R9647 VPWR.n704 VPWR.n703 376.045
R9648 VPWR.n700 VPWR.n699 376.045
R9649 VPWR.n740 VPWR.n739 376.045
R9650 VPWR.n2105 VPWR.n2104 376.045
R9651 VPWR.n2103 VPWR.n2102 376.045
R9652 VPWR.n2095 VPWR.n2094 376.045
R9653 VPWR.n2093 VPWR.n2092 376.045
R9654 VPWR.n2083 VPWR.n2082 376.045
R9655 VPWR.n2075 VPWR.n2074 376.045
R9656 VPWR.n2073 VPWR.n2072 376.045
R9657 VPWR.n2065 VPWR.n2064 376.045
R9658 VPWR.n2063 VPWR.n2062 376.045
R9659 VPWR.n2055 VPWR.n2054 376.045
R9660 VPWR.n2053 VPWR.n2052 376.045
R9661 VPWR.n2045 VPWR.n2044 376.045
R9662 VPWR.n2043 VPWR.n2042 376.045
R9663 VPWR.n2035 VPWR.n2034 376.045
R9664 VPWR.n2085 VPWR.n2084 376.045
R9665 VPWR.n793 VPWR.n792 376.045
R9666 VPWR.n797 VPWR.n796 376.045
R9667 VPWR.n801 VPWR.n800 376.045
R9668 VPWR.n805 VPWR.n804 376.045
R9669 VPWR.n813 VPWR.n812 376.045
R9670 VPWR.n817 VPWR.n816 376.045
R9671 VPWR.n821 VPWR.n820 376.045
R9672 VPWR.n825 VPWR.n824 376.045
R9673 VPWR.n829 VPWR.n828 376.045
R9674 VPWR.n833 VPWR.n832 376.045
R9675 VPWR.n837 VPWR.n836 376.045
R9676 VPWR.n841 VPWR.n840 376.045
R9677 VPWR.n845 VPWR.n844 376.045
R9678 VPWR.n849 VPWR.n848 376.045
R9679 VPWR.n809 VPWR.n808 376.045
R9680 VPWR.n1936 VPWR.n1935 376.045
R9681 VPWR.n1938 VPWR.n1937 376.045
R9682 VPWR.n1946 VPWR.n1945 376.045
R9683 VPWR.n1948 VPWR.n1947 376.045
R9684 VPWR.n1958 VPWR.n1957 376.045
R9685 VPWR.n1966 VPWR.n1965 376.045
R9686 VPWR.n1968 VPWR.n1967 376.045
R9687 VPWR.n1976 VPWR.n1975 376.045
R9688 VPWR.n1978 VPWR.n1977 376.045
R9689 VPWR.n1986 VPWR.n1985 376.045
R9690 VPWR.n1988 VPWR.n1987 376.045
R9691 VPWR.n1996 VPWR.n1995 376.045
R9692 VPWR.n1998 VPWR.n1997 376.045
R9693 VPWR.n2006 VPWR.n2005 376.045
R9694 VPWR.n1956 VPWR.n1955 376.045
R9695 VPWR.n946 VPWR.n945 376.045
R9696 VPWR.n944 VPWR.n943 376.045
R9697 VPWR.n940 VPWR.n939 376.045
R9698 VPWR.n936 VPWR.n935 376.045
R9699 VPWR.n928 VPWR.n927 376.045
R9700 VPWR.n924 VPWR.n923 376.045
R9701 VPWR.n920 VPWR.n919 376.045
R9702 VPWR.n916 VPWR.n915 376.045
R9703 VPWR.n912 VPWR.n911 376.045
R9704 VPWR.n908 VPWR.n907 376.045
R9705 VPWR.n904 VPWR.n903 376.045
R9706 VPWR.n900 VPWR.n899 376.045
R9707 VPWR.n896 VPWR.n895 376.045
R9708 VPWR.n892 VPWR.n891 376.045
R9709 VPWR.n932 VPWR.n931 376.045
R9710 VPWR.n1889 VPWR.n1888 376.045
R9711 VPWR.n1001 VPWR.n1000 376.045
R9712 VPWR.n1513 VPWR.n1512 376.045
R9713 VPWR.n1240 VPWR.n1239 376.045
R9714 VPWR.n421 VPWR.n420 376.045
R9715 VPWR.n2485 VPWR.n2484 376.045
R9716 VPWR.n360 VPWR.n359 376.045
R9717 VPWR.n2539 VPWR.n2538 376.045
R9718 VPWR.n997 VPWR.n996 376.045
R9719 VPWR.n1511 VPWR.n1510 376.045
R9720 VPWR.n1204 VPWR.n1203 376.045
R9721 VPWR.n1887 VPWR.n1886 376.045
R9722 VPWR.n1005 VPWR.n1004 376.045
R9723 VPWR.n1525 VPWR.n1524 376.045
R9724 VPWR.n1238 VPWR.n1237 376.045
R9725 VPWR.n429 VPWR.n428 376.045
R9726 VPWR.n437 VPWR.n436 376.045
R9727 VPWR.n441 VPWR.n440 376.045
R9728 VPWR.n445 VPWR.n444 376.045
R9729 VPWR.n449 VPWR.n448 376.045
R9730 VPWR.n453 VPWR.n452 376.045
R9731 VPWR.n457 VPWR.n456 376.045
R9732 VPWR.n461 VPWR.n460 376.045
R9733 VPWR.n465 VPWR.n464 376.045
R9734 VPWR.n433 VPWR.n432 376.045
R9735 VPWR.n2467 VPWR.n2466 376.045
R9736 VPWR.n348 VPWR.n347 376.045
R9737 VPWR.n2561 VPWR.n2560 376.045
R9738 VPWR.n1009 VPWR.n1008 376.045
R9739 VPWR.n1527 VPWR.n1526 376.045
R9740 VPWR.n1235 VPWR.n1234 376.045
R9741 VPWR.n1879 VPWR.n1878 376.045
R9742 VPWR.n1869 VPWR.n1868 376.045
R9743 VPWR.n1867 VPWR.n1866 376.045
R9744 VPWR.n1859 VPWR.n1858 376.045
R9745 VPWR.n1857 VPWR.n1856 376.045
R9746 VPWR.n1849 VPWR.n1848 376.045
R9747 VPWR.n1847 VPWR.n1846 376.045
R9748 VPWR.n1839 VPWR.n1838 376.045
R9749 VPWR.n1877 VPWR.n1876 376.045
R9750 VPWR.n1013 VPWR.n1012 376.045
R9751 VPWR.n1539 VPWR.n1538 376.045
R9752 VPWR.n1232 VPWR.n1231 376.045
R9753 VPWR.n2487 VPWR.n2486 376.045
R9754 VPWR.n364 VPWR.n363 376.045
R9755 VPWR.n2537 VPWR.n2536 376.045
R9756 VPWR.n1500 VPWR.n1499 376.045
R9757 VPWR.n1201 VPWR.n1200 376.045
R9758 VPWR.n1017 VPWR.n1016 376.045
R9759 VPWR.n1541 VPWR.n1540 376.045
R9760 VPWR.n1224 VPWR.n1223 376.045
R9761 VPWR.n2457 VPWR.n2456 376.045
R9762 VPWR.n2447 VPWR.n2446 376.045
R9763 VPWR.n2445 VPWR.n2444 376.045
R9764 VPWR.n2437 VPWR.n2436 376.045
R9765 VPWR.n2435 VPWR.n2434 376.045
R9766 VPWR.n2427 VPWR.n2426 376.045
R9767 VPWR.n2455 VPWR.n2454 376.045
R9768 VPWR.n336 VPWR.n335 376.045
R9769 VPWR.n2575 VPWR.n2574 376.045
R9770 VPWR.n1556 VPWR.n1555 376.045
R9771 VPWR.n1221 VPWR.n1220 376.045
R9772 VPWR.n1021 VPWR.n1020 376.045
R9773 VPWR.n1025 VPWR.n1024 376.045
R9774 VPWR.n1029 VPWR.n1028 376.045
R9775 VPWR.n1033 VPWR.n1032 376.045
R9776 VPWR.n1037 VPWR.n1036 376.045
R9777 VPWR.n1041 VPWR.n1040 376.045
R9778 VPWR.n989 VPWR.n988 376.045
R9779 VPWR.n1494 VPWR.n1493 376.045
R9780 VPWR.n1612 VPWR.n1611 376.045
R9781 VPWR.n332 VPWR.n331 376.045
R9782 VPWR.n2585 VPWR.n2584 376.045
R9783 VPWR.n1218 VPWR.n1217 376.045
R9784 VPWR.n1781 VPWR.n1780 376.045
R9785 VPWR.n1210 VPWR.n1209 376.045
R9786 VPWR.n328 VPWR.n327 376.045
R9787 VPWR.n324 VPWR.n323 376.045
R9788 VPWR.n316 VPWR.n315 376.045
R9789 VPWR.n320 VPWR.n319 376.045
R9790 VPWR.n1760 VPWR.n1759 376.045
R9791 VPWR.n1769 VPWR.n1768 376.045
R9792 VPWR.n1810 VPWR.n1809 376.045
R9793 VPWR.n1779 VPWR.n1778 376.045
R9794 VPWR.n1207 VPWR.n1206 376.045
R9795 VPWR.n2597 VPWR.n2596 376.045
R9796 VPWR.n2599 VPWR.n2598 376.045
R9797 VPWR.n2609 VPWR.n2608 376.045
R9798 VPWR.n1758 VPWR.n1757 376.045
R9799 VPWR.n2842 VPWR.n2834 350.719
R9800 VPWR.n2842 VPWR.n2841 350.719
R9801 VPWR.n2837 VPWR.n25 350.719
R9802 VPWR.n2837 VPWR.n2836 350.719
R9803 VPWR.n1358 VPWR.t37 342.841
R9804 VPWR.n1397 VPWR.t161 342.841
R9805 VPWR.n1434 VPWR.t118 342.841
R9806 VPWR.n2712 VPWR.t1922 342.841
R9807 VPWR.n2675 VPWR.t1894 342.841
R9808 VPWR.n2618 VPWR.t942 342.841
R9809 VPWR.n1358 VPWR.t108 342.839
R9810 VPWR.n1397 VPWR.t659 342.839
R9811 VPWR.n1434 VPWR.t764 342.839
R9812 VPWR.n2712 VPWR.t1171 342.839
R9813 VPWR.n2675 VPWR.t89 342.839
R9814 VPWR.n2618 VPWR.t123 342.839
R9815 VPWR.n1325 VPWR.t450 338.488
R9816 VPWR.n2748 VPWR.t619 338.488
R9817 VPWR.n1334 VPWR.n1333 327.377
R9818 VPWR.n1327 VPWR.n1326 327.377
R9819 VPWR.n1341 VPWR.n1340 327.377
R9820 VPWR.n1371 VPWR.n1369 327.377
R9821 VPWR.n1364 VPWR.n1362 327.377
R9822 VPWR.n1379 VPWR.n1377 327.377
R9823 VPWR.n1410 VPWR.n1408 327.377
R9824 VPWR.n1403 VPWR.n1401 327.377
R9825 VPWR.n1418 VPWR.n1416 327.377
R9826 VPWR.n1447 VPWR.n1445 327.377
R9827 VPWR.n1440 VPWR.n1438 327.377
R9828 VPWR.n1455 VPWR.n1453 327.377
R9829 VPWR.n1343 VPWR.n1342 327.375
R9830 VPWR.n1371 VPWR.n1370 327.375
R9831 VPWR.n1364 VPWR.n1363 327.375
R9832 VPWR.n1379 VPWR.n1378 327.375
R9833 VPWR.n1410 VPWR.n1409 327.375
R9834 VPWR.n1403 VPWR.n1402 327.375
R9835 VPWR.n1418 VPWR.n1417 327.375
R9836 VPWR.n1447 VPWR.n1446 327.375
R9837 VPWR.n1440 VPWR.n1439 327.375
R9838 VPWR.n1455 VPWR.n1454 327.375
R9839 VPWR.n2848 VPWR.t1797 326.106
R9840 VPWR.n2852 VPWR.t494 326.106
R9841 VPWR.n2837 VPWR.t569 326.106
R9842 VPWR.n2842 VPWR.t570 326.106
R9843 VPWR.n1 VPWR 325.546
R9844 VPWR.n2686 VPWR.t1170 322.262
R9845 VPWR.n2649 VPWR.t88 322.262
R9846 VPWR.n2824 VPWR.n2823 321.642
R9847 VPWR.n2741 VPWR.n2731 320.976
R9848 VPWR.n2735 VPWR.n2734 320.976
R9849 VPWR.n2729 VPWR.n2728 320.976
R9850 VPWR.n2699 VPWR.n2698 320.976
R9851 VPWR.n2705 VPWR.n2694 320.976
R9852 VPWR.n2691 VPWR.n2690 320.976
R9853 VPWR.n2662 VPWR.n2661 320.976
R9854 VPWR.n2668 VPWR.n2657 320.976
R9855 VPWR.n2654 VPWR.n2653 320.976
R9856 VPWR.n2629 VPWR.n2625 320.976
R9857 VPWR.n2633 VPWR.n2632 320.976
R9858 VPWR.n2639 VPWR.n2621 320.976
R9859 VPWR.n2746 VPWR.n2727 320.976
R9860 VPWR.n2699 VPWR.n2697 320.976
R9861 VPWR.n2705 VPWR.n2693 320.976
R9862 VPWR.n2691 VPWR.n2689 320.976
R9863 VPWR.n2662 VPWR.n2660 320.976
R9864 VPWR.n2668 VPWR.n2656 320.976
R9865 VPWR.n2654 VPWR.n2652 320.976
R9866 VPWR.n2629 VPWR.n2624 320.976
R9867 VPWR.n2633 VPWR.n2631 320.976
R9868 VPWR.n2639 VPWR.n2620 320.976
R9869 VPWR.n2820 VPWR 319.627
R9870 VPWR.n6 VPWR.n5 316.245
R9871 VPWR.n1260 VPWR.n1258 316.245
R9872 VPWR.n1283 VPWR.n1281 316.245
R9873 VPWR.n1307 VPWR.n1305 316.245
R9874 VPWR.n2803 VPWR.n2802 316.245
R9875 VPWR.n2783 VPWR.n2782 316.245
R9876 VPWR.n2764 VPWR.n2763 316.245
R9877 VPWR.n1260 VPWR.n1259 316.245
R9878 VPWR.n1283 VPWR.n1282 316.245
R9879 VPWR.n1307 VPWR.n1306 316.245
R9880 VPWR.n2803 VPWR.n2801 316.245
R9881 VPWR.n2783 VPWR.n2781 316.245
R9882 VPWR.n2764 VPWR.n2762 316.245
R9883 VPWR.n2649 VPWR.t168 313.87
R9884 VPWR.n10 VPWR.n4 310.502
R9885 VPWR.n1265 VPWR.n1257 310.502
R9886 VPWR.n1288 VPWR.n1280 310.502
R9887 VPWR.n1312 VPWR.n1304 310.502
R9888 VPWR.n2822 VPWR.n2821 310.502
R9889 VPWR.n2807 VPWR.n2806 310.502
R9890 VPWR.n2787 VPWR.n2786 310.502
R9891 VPWR.n2768 VPWR.n2767 310.502
R9892 VPWR.n1265 VPWR.n1264 310.5
R9893 VPWR.n1288 VPWR.n1287 310.5
R9894 VPWR.n1312 VPWR.n1311 310.5
R9895 VPWR.n2807 VPWR.n2805 310.5
R9896 VPWR.n2787 VPWR.n2785 310.5
R9897 VPWR.n2768 VPWR.n2766 310.5
R9898 VPWR.t833 VPWR.t747 297.909
R9899 VPWR.n2855 VPWR.n2854 292.5
R9900 VPWR.n33 VPWR.n32 292.5
R9901 VPWR.n2839 VPWR.t568 272.257
R9902 VPWR.n2853 VPWR.n2852 256.226
R9903 VPWR.n2848 VPWR.n31 256.226
R9904 VPWR.n1431 VPWR.t707 255.905
R9905 VPWR.n2682 VPWR.t1798 255.905
R9906 VPWR.n1294 VPWR.t730 255.904
R9907 VPWR.n1431 VPWR.t1268 255.904
R9908 VPWR.n2793 VPWR.t879 255.904
R9909 VPWR.n2682 VPWR.t169 255.904
R9910 VPWR.n26 VPWR.n24 255.653
R9911 VPWR.n2847 VPWR.n35 255.653
R9912 VPWR.n1322 VPWR.t471 254.019
R9913 VPWR.n2754 VPWR.t740 254.019
R9914 VPWR.n1354 VPWR.t469 252.948
R9915 VPWR.n2756 VPWR.t738 252.948
R9916 VPWR.n1392 VPWR.t1318 250.722
R9917 VPWR.n2719 VPWR.t155 250.722
R9918 VPWR.n1329 VPWR.t1371 249.901
R9919 VPWR.n1365 VPWR.t891 249.901
R9920 VPWR.n1404 VPWR.t401 249.901
R9921 VPWR.n1441 VPWR.t893 249.901
R9922 VPWR.n2733 VPWR.t379 249.901
R9923 VPWR.n2696 VPWR.t420 249.901
R9924 VPWR.n2659 VPWR.t695 249.901
R9925 VPWR.n2626 VPWR.t274 249.901
R9926 VPWR.n1365 VPWR.t474 249.901
R9927 VPWR.n1404 VPWR.t269 249.901
R9928 VPWR.n1441 VPWR.t430 249.901
R9929 VPWR.n2696 VPWR.t696 249.901
R9930 VPWR.n2659 VPWR.t276 249.901
R9931 VPWR.n2626 VPWR.t199 249.901
R9932 VPWR.n1272 VPWR.t1405 249.363
R9933 VPWR.n1357 VPWR.t605 249.363
R9934 VPWR.n2830 VPWR.t925 249.363
R9935 VPWR.n2814 VPWR.t1889 249.363
R9936 VPWR.n2717 VPWR.t1109 249.363
R9937 VPWR.n17 VPWR.t761 249.362
R9938 VPWR.n1272 VPWR.t1882 249.362
R9939 VPWR.n2814 VPWR.t964 249.362
R9940 VPWR.t726 VPWR.t760 248.599
R9941 VPWR.t626 VPWR.t1829 248.599
R9942 VPWR.t1829 VPWR.t1833 248.599
R9943 VPWR.t1833 VPWR.t622 248.599
R9944 VPWR.t622 VPWR.t1346 248.599
R9945 VPWR.t1346 VPWR.t1366 248.599
R9946 VPWR.t1366 VPWR.t890 248.599
R9947 VPWR.t890 VPWR.t895 248.599
R9948 VPWR.t319 VPWR.t472 248.599
R9949 VPWR.t472 VPWR.t1370 248.599
R9950 VPWR.t693 VPWR.t427 248.599
R9951 VPWR.t309 VPWR.t693 248.599
R9952 VPWR.t1857 VPWR.t309 248.599
R9953 VPWR.t616 VPWR.t1857 248.599
R9954 VPWR.t1130 VPWR.t616 248.599
R9955 VPWR.t854 VPWR.t1130 248.599
R9956 VPWR.t175 VPWR.t854 248.599
R9957 VPWR.t880 VPWR.t924 248.599
R9958 VPWR.t283 VPWR.t378 248.599
R9959 VPWR.t372 VPWR.t283 248.599
R9960 VPWR.n15 VPWR.t727 247.394
R9961 VPWR.n1270 VPWR.t729 247.394
R9962 VPWR.n2828 VPWR.t881 247.394
R9963 VPWR.n2812 VPWR.t875 247.394
R9964 VPWR.n1270 VPWR.t728 247.394
R9965 VPWR.n2812 VPWR.t877 247.394
R9966 VPWR.n1323 VPWR.t264 244.737
R9967 VPWR.n2749 VPWR.t467 244.737
R9968 VPWR.n1393 VPWR.t1404 243.886
R9969 VPWR.n2720 VPWR.t93 243.886
R9970 VPWR.n1296 VPWR.t759 243.512
R9971 VPWR.n1319 VPWR.t1406 243.512
R9972 VPWR.n1322 VPWR.t918 243.512
R9973 VPWR.n2795 VPWR.t927 243.512
R9974 VPWR.n2775 VPWR.t1890 243.512
R9975 VPWR.n2754 VPWR.t99 243.512
R9976 VPWR.n1319 VPWR.t1883 243.512
R9977 VPWR.n2775 VPWR.t962 243.512
R9978 VPWR.n1348 VPWR.t470 238.339
R9979 VPWR.n2724 VPWR.t739 238.339
R9980 VPWR.n2686 VPWR.t1108 234.982
R9981 VPWR.t317 VPWR.t319 228.101
R9982 VPWR.t203 VPWR.t372 228.101
R9983 VPWR.n2820 VPWR 224.923
R9984 VPWR.n1 VPWR 219.004
R9985 VPWR.n1463 VPWR.n1462 214.613
R9986 VPWR.n1463 VPWR.n1461 214.613
R9987 VPWR.n1255 VPWR.n1254 214.326
R9988 VPWR.n1278 VPWR.n1277 214.326
R9989 VPWR.n1302 VPWR.n1301 214.326
R9990 VPWR.n1387 VPWR.n1386 214.326
R9991 VPWR.n1426 VPWR.n1425 214.326
R9992 VPWR.n1255 VPWR.n1253 214.326
R9993 VPWR.n1278 VPWR.n1276 214.326
R9994 VPWR.n1302 VPWR.n1300 214.326
R9995 VPWR.n1387 VPWR.n1385 214.326
R9996 VPWR.n1426 VPWR.n1424 214.326
R9997 VPWR.n2 VPWR.n1 213.119
R9998 VPWR.n2827 VPWR.n2820 213.119
R9999 VPWR VPWR.t726 207.166
R10000 VPWR VPWR.t175 201.246
R10001 VPWR.t747 VPWR.t493 200.262
R10002 VPWR.t1370 VPWR 189.409
R10003 VPWR.n2760 VPWR 184.63
R10004 VPWR.n1348 VPWR 182.952
R10005 VPWR.n2779 VPWR 182.952
R10006 VPWR.n2799 VPWR 181.273
R10007 VPWR.t168 VPWR 177.916
R10008 VPWR.n1789 VPWR.n1787 161.365
R10009 VPWR.n1060 VPWR.n1058 161.365
R10010 VPWR.n1564 VPWR.n1562 161.365
R10011 VPWR.n1569 VPWR.n1567 161.365
R10012 VPWR.n1574 VPWR.n1572 161.365
R10013 VPWR.n1579 VPWR.n1577 161.365
R10014 VPWR.n1584 VPWR.n1582 161.365
R10015 VPWR.n1589 VPWR.n1587 161.365
R10016 VPWR.n1594 VPWR.n1592 161.365
R10017 VPWR.n1599 VPWR.n1597 161.365
R10018 VPWR.n1154 VPWR.n1152 161.365
R10019 VPWR.n1479 VPWR.n1477 161.365
R10020 VPWR.n1474 VPWR.n1472 161.365
R10021 VPWR.n1794 VPWR.n1792 161.365
R10022 VPWR.n1802 VPWR.n1800 161.365
R10023 VPWR.n1798 VPWR.n1796 161.365
R10024 VPWR VPWR.n72 161.363
R10025 VPWR VPWR.n70 161.363
R10026 VPWR VPWR.n68 161.363
R10027 VPWR VPWR.n66 161.363
R10028 VPWR VPWR.n64 161.363
R10029 VPWR VPWR.n62 161.363
R10030 VPWR VPWR.n60 161.363
R10031 VPWR VPWR.n58 161.363
R10032 VPWR VPWR.n56 161.363
R10033 VPWR VPWR.n54 161.363
R10034 VPWR VPWR.n52 161.363
R10035 VPWR VPWR.n50 161.363
R10036 VPWR VPWR.n48 161.363
R10037 VPWR VPWR.n46 161.363
R10038 VPWR VPWR.n44 161.363
R10039 VPWR VPWR.n42 161.363
R10040 VPWR.n1134 VPWR.n1133 161.303
R10041 VPWR.n126 VPWR.n125 161.303
R10042 VPWR.n1139 VPWR.n1138 161.3
R10043 VPWR.n1618 VPWR.n1617 161.3
R10044 VPWR.n1621 VPWR.n1620 161.3
R10045 VPWR.n1130 VPWR.n1129 161.3
R10046 VPWR.n1145 VPWR.n1144 161.3
R10047 VPWR.n1126 VPWR.n1125 161.3
R10048 VPWR.n1631 VPWR.n1630 161.3
R10049 VPWR.n1634 VPWR.n1633 161.3
R10050 VPWR.n1637 VPWR.n1636 161.3
R10051 VPWR.n1642 VPWR.n1641 161.3
R10052 VPWR.n1645 VPWR.n1644 161.3
R10053 VPWR.n1648 VPWR.n1647 161.3
R10054 VPWR.n1120 VPWR.n1119 161.3
R10055 VPWR.n1196 VPWR.n1195 161.3
R10056 VPWR.n1116 VPWR.n1115 161.3
R10057 VPWR.n1658 VPWR.n1657 161.3
R10058 VPWR.n1661 VPWR.n1660 161.3
R10059 VPWR.n1664 VPWR.n1663 161.3
R10060 VPWR.n1669 VPWR.n1668 161.3
R10061 VPWR.n1672 VPWR.n1671 161.3
R10062 VPWR.n1675 VPWR.n1674 161.3
R10063 VPWR.n1110 VPWR.n1109 161.3
R10064 VPWR.n1228 VPWR.n1227 161.3
R10065 VPWR.n1106 VPWR.n1105 161.3
R10066 VPWR.n1685 VPWR.n1684 161.3
R10067 VPWR.n1688 VPWR.n1687 161.3
R10068 VPWR.n1691 VPWR.n1690 161.3
R10069 VPWR.n1696 VPWR.n1695 161.3
R10070 VPWR.n1699 VPWR.n1698 161.3
R10071 VPWR.n1702 VPWR.n1701 161.3
R10072 VPWR.n1100 VPWR.n1099 161.3
R10073 VPWR.n1214 VPWR.n1213 161.3
R10074 VPWR.n1096 VPWR.n1095 161.3
R10075 VPWR.n1712 VPWR.n1711 161.3
R10076 VPWR.n1715 VPWR.n1714 161.3
R10077 VPWR.n1718 VPWR.n1717 161.3
R10078 VPWR.n1723 VPWR.n1722 161.3
R10079 VPWR.n1726 VPWR.n1725 161.3
R10080 VPWR.n1729 VPWR.n1728 161.3
R10081 VPWR.n1089 VPWR.n1088 161.3
R10082 VPWR.n1738 VPWR.n1737 161.3
R10083 VPWR.n1741 VPWR.n1740 161.3
R10084 VPWR.n1736 VPWR.n1735 161.3
R10085 VPWR.n1753 VPWR.n1752 161.3
R10086 VPWR.n1136 VPWR.n1135 161.3
R10087 VPWR.n1750 VPWR.n1749 161.3
R10088 VPWR.n1084 VPWR.n1083 161.3
R10089 VPWR.n145 VPWR.n144 161.3
R10090 VPWR.n136 VPWR.n135 161.3
R10091 VPWR.n139 VPWR.n138 161.3
R10092 VPWR.n134 VPWR.n133 161.3
R10093 VPWR.n157 VPWR.n156 161.3
R10094 VPWR.n147 VPWR.n146 161.3
R10095 VPWR.n128 VPWR.n127 161.3
R10096 VPWR.n124 VPWR.n123 161.3
R10097 VPWR.n307 VPWR.n306 161.3
R10098 VPWR.n304 VPWR.n303 161.3
R10099 VPWR.n120 VPWR.n119 161.3
R10100 VPWR.n291 VPWR.n290 161.3
R10101 VPWR.n294 VPWR.n293 161.3
R10102 VPWR.n289 VPWR.n288 161.3
R10103 VPWR.n279 VPWR.n278 161.3
R10104 VPWR.n282 VPWR.n281 161.3
R10105 VPWR.n277 VPWR.n276 161.3
R10106 VPWR.n267 VPWR.n266 161.3
R10107 VPWR.n270 VPWR.n269 161.3
R10108 VPWR.n265 VPWR.n264 161.3
R10109 VPWR.n255 VPWR.n254 161.3
R10110 VPWR.n258 VPWR.n257 161.3
R10111 VPWR.n253 VPWR.n252 161.3
R10112 VPWR.n243 VPWR.n242 161.3
R10113 VPWR.n246 VPWR.n245 161.3
R10114 VPWR.n241 VPWR.n240 161.3
R10115 VPWR.n231 VPWR.n230 161.3
R10116 VPWR.n234 VPWR.n233 161.3
R10117 VPWR.n229 VPWR.n228 161.3
R10118 VPWR.n219 VPWR.n218 161.3
R10119 VPWR.n222 VPWR.n221 161.3
R10120 VPWR.n217 VPWR.n216 161.3
R10121 VPWR.n207 VPWR.n206 161.3
R10122 VPWR.n210 VPWR.n209 161.3
R10123 VPWR.n205 VPWR.n204 161.3
R10124 VPWR.n195 VPWR.n194 161.3
R10125 VPWR.n198 VPWR.n197 161.3
R10126 VPWR.n193 VPWR.n192 161.3
R10127 VPWR.n183 VPWR.n182 161.3
R10128 VPWR.n186 VPWR.n185 161.3
R10129 VPWR.n181 VPWR.n180 161.3
R10130 VPWR.n171 VPWR.n170 161.3
R10131 VPWR.n174 VPWR.n173 161.3
R10132 VPWR.n169 VPWR.n168 161.3
R10133 VPWR.n159 VPWR.n158 161.3
R10134 VPWR.n162 VPWR.n161 161.3
R10135 VPWR.n150 VPWR.n149 161.3
R10136 VPWR.n1620 VPWR.t1456 161.202
R10137 VPWR.n1125 VPWR.t1584 161.202
R10138 VPWR.n1636 VPWR.t1625 161.202
R10139 VPWR.n1647 VPWR.t1736 161.202
R10140 VPWR.n1115 VPWR.t1500 161.202
R10141 VPWR.n1663 VPWR.t1515 161.202
R10142 VPWR.n1674 VPWR.t1741 161.202
R10143 VPWR.n1105 VPWR.t1781 161.202
R10144 VPWR.n1690 VPWR.t1498 161.202
R10145 VPWR.n1701 VPWR.t1651 161.202
R10146 VPWR.n1095 VPWR.t1676 161.202
R10147 VPWR.n1717 VPWR.t1523 161.202
R10148 VPWR.n1728 VPWR.t1549 161.202
R10149 VPWR.n1740 VPWR.t1574 161.202
R10150 VPWR.n1135 VPWR.t1720 161.202
R10151 VPWR.n1749 VPWR.t1419 161.202
R10152 VPWR.n138 VPWR.t1541 161.202
R10153 VPWR.n127 VPWR.t1440 161.202
R10154 VPWR.n303 VPWR.t1576 161.202
R10155 VPWR.n293 VPWR.t1712 161.202
R10156 VPWR.n281 VPWR.t1746 161.202
R10157 VPWR.n269 VPWR.t1470 161.202
R10158 VPWR.n257 VPWR.t1614 161.202
R10159 VPWR.n245 VPWR.t1638 161.202
R10160 VPWR.n233 VPWR.t1475 161.202
R10161 VPWR.n221 VPWR.t1510 161.202
R10162 VPWR.n209 VPWR.t1612 161.202
R10163 VPWR.n197 VPWR.t1773 161.202
R10164 VPWR.n185 VPWR.t1792 161.202
R10165 VPWR.n173 VPWR.t1646 161.202
R10166 VPWR.n1787 VPWR.t1704 161.202
R10167 VPWR.n1058 VPWR.t1451 161.202
R10168 VPWR.n1562 VPWR.t1435 161.202
R10169 VPWR.n1567 VPWR.t1684 161.202
R10170 VPWR.n1572 VPWR.t1566 161.202
R10171 VPWR.n1577 VPWR.t1536 161.202
R10172 VPWR.n1582 VPWR.t1688 161.202
R10173 VPWR.n1587 VPWR.t1686 161.202
R10174 VPWR.n1592 VPWR.t1531 161.202
R10175 VPWR.n1597 VPWR.t1421 161.202
R10176 VPWR.n1152 VPWR.t1765 161.202
R10177 VPWR.n1477 VPWR.t1636 161.202
R10178 VPWR.n1472 VPWR.t1505 161.202
R10179 VPWR.n1792 VPWR.t1722 161.202
R10180 VPWR.n1800 VPWR.t1757 161.202
R10181 VPWR.n1796 VPWR.t1586 161.202
R10182 VPWR.n161 VPWR.t1668 161.202
R10183 VPWR.n149 VPWR.t1690 161.202
R10184 VPWR.n1138 VPWR.t1442 161.106
R10185 VPWR.n1129 VPWR.t1578 161.106
R10186 VPWR.n1630 VPWR.t1591 161.106
R10187 VPWR.n1641 VPWR.t1754 161.106
R10188 VPWR.n1119 VPWR.t1472 161.106
R10189 VPWR.n1657 VPWR.t1619 161.106
R10190 VPWR.n1668 VPWR.t1730 161.106
R10191 VPWR.n1109 VPWR.t1767 161.106
R10192 VPWR.n1684 VPWR.t1512 161.106
R10193 VPWR.n1695 VPWR.t1616 161.106
R10194 VPWR.n1099 VPWR.t1775 161.106
R10195 VPWR.n1711 VPWR.t1794 161.106
R10196 VPWR.n1722 VPWR.t1538 161.106
R10197 VPWR.n1088 VPWR.t1670 161.106
R10198 VPWR.n1735 VPWR.t1701 161.106
R10199 VPWR.n1083 VPWR.t1546 161.106
R10200 VPWR.n144 VPWR.t1426 161.106
R10201 VPWR.n133 VPWR.t1662 161.106
R10202 VPWR.n156 VPWR.t1786 161.106
R10203 VPWR.n123 VPWR.t1571 161.106
R10204 VPWR.n119 VPWR.t1706 161.106
R10205 VPWR.n288 VPWR.t1698 161.106
R10206 VPWR.n276 VPWR.t1480 161.106
R10207 VPWR.n264 VPWR.t1588 161.106
R10208 VPWR.n252 VPWR.t1743 161.106
R10209 VPWR.n240 VPWR.t1467 161.106
R10210 VPWR.n228 VPWR.t1502 161.106
R10211 VPWR.n216 VPWR.t1630 161.106
R10212 VPWR.n204 VPWR.t1695 161.106
R10213 VPWR.n192 VPWR.t1507 161.106
R10214 VPWR.n180 VPWR.t1525 161.106
R10215 VPWR.n168 VPWR.t1653 161.106
R10216 VPWR.n72 VPWR.t1770 161.106
R10217 VPWR.n70 VPWR.t1733 161.106
R10218 VPWR.n68 VPWR.t1445 161.106
R10219 VPWR.n66 VPWR.t1560 161.106
R10220 VPWR.n64 VPWR.t1778 161.106
R10221 VPWR.n62 VPWR.t1627 161.106
R10222 VPWR.n60 VPWR.t1738 161.106
R10223 VPWR.n58 VPWR.t1461 161.106
R10224 VPWR.n56 VPWR.t1568 161.106
R10225 VPWR.n54 VPWR.t1528 161.106
R10226 VPWR.n52 VPWR.t1633 161.106
R10227 VPWR.n50 VPWR.t1453 161.106
R10228 VPWR.n48 VPWR.t1640 161.106
R10229 VPWR.n46 VPWR.t1748 161.106
R10230 VPWR.n44 VPWR.t1600 161.106
R10231 VPWR.n42 VPWR.t1717 161.106
R10232 VPWR.n1617 VPWR.t1492 159.978
R10233 VPWR.n1144 VPWR.t1597 159.978
R10234 VPWR.n1633 VPWR.t1759 159.978
R10235 VPWR.n1644 VPWR.t1477 159.978
R10236 VPWR.n1195 VPWR.t1489 159.978
R10237 VPWR.n1660 VPWR.t1648 159.978
R10238 VPWR.n1671 VPWR.t1751 159.978
R10239 VPWR.n1227 VPWR.t1517 159.978
R10240 VPWR.n1687 VPWR.t1543 159.978
R10241 VPWR.n1698 VPWR.t1665 159.978
R10242 VPWR.n1213 VPWR.t1416 159.978
R10243 VPWR.n1714 VPWR.t1437 159.978
R10244 VPWR.n1725 VPWR.t1678 159.978
R10245 VPWR.n1737 VPWR.t1709 159.978
R10246 VPWR.n1752 VPWR.t1423 159.978
R10247 VPWR.n1133 VPWR.t1727 159.978
R10248 VPWR.n135 VPWR.t1557 159.978
R10249 VPWR.n146 VPWR.t1432 159.978
R10250 VPWR.n125 VPWR.t1464 159.978
R10251 VPWR.n306 VPWR.t1609 159.978
R10252 VPWR.n290 VPWR.t1724 159.978
R10253 VPWR.n278 VPWR.t1486 159.978
R10254 VPWR.n266 VPWR.t1594 159.978
R10255 VPWR.n254 VPWR.t1606 159.978
R10256 VPWR.n242 VPWR.t1762 159.978
R10257 VPWR.n230 VPWR.t1483 159.978
R10258 VPWR.n218 VPWR.t1643 159.978
R10259 VPWR.n206 VPWR.t1659 159.978
R10260 VPWR.n194 VPWR.t1789 159.978
R10261 VPWR.n182 VPWR.t1533 159.978
R10262 VPWR.n170 VPWR.t1563 159.978
R10263 VPWR.n1247 VPWR.t1520 159.978
R10264 VPWR.n1169 VPWR.t1448 159.978
R10265 VPWR.n1243 VPWR.t1656 159.978
R10266 VPWR.n1501 VPWR.t1554 159.978
R10267 VPWR.n1189 VPWR.t1681 159.978
R10268 VPWR.n1185 VPWR.t1429 159.978
R10269 VPWR.n1179 VPWR.t1551 159.978
R10270 VPWR.n1495 VPWR.t1783 159.978
R10271 VPWR.n1175 VPWR.t1692 159.978
R10272 VPWR.n1165 VPWR.t1714 159.978
R10273 VPWR.n1488 VPWR.t1673 159.978
R10274 VPWR.n1065 VPWR.t1581 159.978
R10275 VPWR.n1764 VPWR.t1458 159.978
R10276 VPWR.n1052 VPWR.t1495 159.978
R10277 VPWR.n1048 VPWR.t1603 159.978
R10278 VPWR.n1069 VPWR.t1622 159.978
R10279 VPWR.n158 VPWR.t1413 159.978
R10280 VPWR.n1248 VPWR.n1247 152
R10281 VPWR.n1170 VPWR.n1169 152
R10282 VPWR.n1244 VPWR.n1243 152
R10283 VPWR.n1502 VPWR.n1501 152
R10284 VPWR.n1190 VPWR.n1189 152
R10285 VPWR.n1186 VPWR.n1185 152
R10286 VPWR.n1180 VPWR.n1179 152
R10287 VPWR.n1496 VPWR.n1495 152
R10288 VPWR.n1176 VPWR.n1175 152
R10289 VPWR.n1166 VPWR.n1165 152
R10290 VPWR.n1489 VPWR.n1488 152
R10291 VPWR.n1066 VPWR.n1065 152
R10292 VPWR.n1765 VPWR.n1764 152
R10293 VPWR.n1053 VPWR.n1052 152
R10294 VPWR.n1049 VPWR.n1048 152
R10295 VPWR.n1070 VPWR.n1069 152
R10296 VPWR.n2850 VPWR.t493 148.127
R10297 VPWR.n1620 VPWR.t2068 145.137
R10298 VPWR.n1125 VPWR.t2019 145.137
R10299 VPWR.n1636 VPWR.t2005 145.137
R10300 VPWR.n1647 VPWR.t1967 145.137
R10301 VPWR.n1115 VPWR.t2054 145.137
R10302 VPWR.n1663 VPWR.t2047 145.137
R10303 VPWR.n1674 VPWR.t1964 145.137
R10304 VPWR.n1105 VPWR.t1950 145.137
R10305 VPWR.n1690 VPWR.t2055 145.137
R10306 VPWR.n1701 VPWR.t1998 145.137
R10307 VPWR.n1095 VPWR.t1993 145.137
R10308 VPWR.n1717 VPWR.t2045 145.137
R10309 VPWR.n1728 VPWR.t2038 145.137
R10310 VPWR.n1740 VPWR.t2024 145.137
R10311 VPWR.n1135 VPWR.t1974 145.137
R10312 VPWR.n1749 VPWR.t1942 145.137
R10313 VPWR.n138 VPWR.t2053 145.137
R10314 VPWR.n127 VPWR.t1939 145.137
R10315 VPWR.n303 VPWR.t2035 145.137
R10316 VPWR.n293 VPWR.t1988 145.137
R10317 VPWR.n281 VPWR.t1976 145.137
R10318 VPWR.n269 VPWR.t1935 145.137
R10319 VPWR.n257 VPWR.t2021 145.137
R10320 VPWR.n245 VPWR.t2013 145.137
R10321 VPWR.n233 VPWR.t1933 145.137
R10322 VPWR.n221 VPWR.t2062 145.137
R10323 VPWR.n209 VPWR.t2022 145.137
R10324 VPWR.n197 VPWR.t1966 145.137
R10325 VPWR.n185 VPWR.t1957 145.137
R10326 VPWR.n173 VPWR.t2012 145.137
R10327 VPWR.n1787 VPWR.t1981 145.137
R10328 VPWR.n1058 VPWR.t2070 145.137
R10329 VPWR.n1562 VPWR.t1934 145.137
R10330 VPWR.n1567 VPWR.t1991 145.137
R10331 VPWR.n1572 VPWR.t2030 145.137
R10332 VPWR.n1577 VPWR.t2042 145.137
R10333 VPWR.n1582 VPWR.t1984 145.137
R10334 VPWR.n1587 VPWR.t1990 145.137
R10335 VPWR.n1592 VPWR.t2044 145.137
R10336 VPWR.n1597 VPWR.t1941 145.137
R10337 VPWR.n1152 VPWR.t1955 145.137
R10338 VPWR.n1477 VPWR.t2001 145.137
R10339 VPWR.n1472 VPWR.t2050 145.137
R10340 VPWR.n1792 VPWR.t1973 145.137
R10341 VPWR.n1800 VPWR.t1958 145.137
R10342 VPWR.n1796 VPWR.t2018 145.137
R10343 VPWR.n161 VPWR.t2004 145.137
R10344 VPWR.n149 VPWR.t1995 145.137
R10345 VPWR.n1138 VPWR.t2072 145.038
R10346 VPWR.n1129 VPWR.t2023 145.038
R10347 VPWR.n1630 VPWR.t2015 145.038
R10348 VPWR.n1641 VPWR.t1960 145.038
R10349 VPWR.n1119 VPWR.t2064 145.038
R10350 VPWR.n1657 VPWR.t2007 145.038
R10351 VPWR.n1668 VPWR.t1969 145.038
R10352 VPWR.n1109 VPWR.t1954 145.038
R10353 VPWR.n1684 VPWR.t2048 145.038
R10354 VPWR.n1695 VPWR.t2008 145.038
R10355 VPWR.n1099 VPWR.t1952 145.038
R10356 VPWR.n1711 VPWR.t1944 145.038
R10357 VPWR.n1722 VPWR.t2041 145.038
R10358 VPWR.n1088 VPWR.t1994 145.038
R10359 VPWR.n1735 VPWR.t1982 145.038
R10360 VPWR.n1083 VPWR.t2039 145.038
R10361 VPWR.n144 VPWR.t1945 145.038
R10362 VPWR.n133 VPWR.t2006 145.038
R10363 VPWR.n156 VPWR.t1959 145.038
R10364 VPWR.n123 VPWR.t2037 145.038
R10365 VPWR.n119 VPWR.t1992 145.038
R10366 VPWR.n288 VPWR.t1985 145.038
R10367 VPWR.n276 VPWR.t2073 145.038
R10368 VPWR.n264 VPWR.t2032 145.038
R10369 VPWR.n252 VPWR.t1977 145.038
R10370 VPWR.n240 VPWR.t1936 145.038
R10371 VPWR.n228 VPWR.t2065 145.038
R10372 VPWR.n216 VPWR.t2014 145.038
R10373 VPWR.n204 VPWR.t1978 145.038
R10374 VPWR.n192 VPWR.t2063 145.038
R10375 VPWR.n180 VPWR.t2057 145.038
R10376 VPWR.n168 VPWR.t2009 145.038
R10377 VPWR.n72 VPWR.t2058 145.038
R10378 VPWR.n70 VPWR.t1968 145.038
R10379 VPWR.n68 VPWR.t2071 145.038
R10380 VPWR.n66 VPWR.t2031 145.038
R10381 VPWR.n64 VPWR.t1951 145.038
R10382 VPWR.n62 VPWR.t2056 145.038
R10383 VPWR.n60 VPWR.t2074 145.038
R10384 VPWR.n58 VPWR.t2033 145.038
R10385 VPWR.n56 VPWR.t2027 145.038
R10386 VPWR.n54 VPWR.t1948 145.038
R10387 VPWR.n52 VPWR.t2002 145.038
R10388 VPWR.n50 VPWR.t2069 145.038
R10389 VPWR.n48 VPWR.t2000 145.038
R10390 VPWR.n46 VPWR.t1961 145.038
R10391 VPWR.n44 VPWR.t2026 145.038
R10392 VPWR.n42 VPWR.t1975 145.038
R10393 VPWR.n1617 VPWR.t1971 143.911
R10394 VPWR.n1144 VPWR.t2067 143.911
R10395 VPWR.n1633 VPWR.t2052 143.911
R10396 VPWR.n1644 VPWR.t1970 143.911
R10397 VPWR.n1195 VPWR.t1963 143.911
R10398 VPWR.n1660 VPWR.t1949 143.911
R10399 VPWR.n1671 VPWR.t2010 143.911
R10400 VPWR.n1227 VPWR.t1997 143.911
R10401 VPWR.n1687 VPWR.t1946 143.911
R10402 VPWR.n1698 VPWR.t2043 143.911
R10403 VPWR.n1213 VPWR.t2036 143.911
R10404 VPWR.n1714 VPWR.t1983 143.911
R10405 VPWR.n1725 VPWR.t1940 143.911
R10406 VPWR.n1737 VPWR.t2029 143.911
R10407 VPWR.n1752 VPWR.t1989 143.911
R10408 VPWR.n1133 VPWR.t2017 143.911
R10409 VPWR.n135 VPWR.t1956 143.911
R10410 VPWR.n146 VPWR.t1996 143.911
R10411 VPWR.n125 VPWR.t1986 143.911
R10412 VPWR.n306 VPWR.t1938 143.911
R10413 VPWR.n290 VPWR.t2034 143.911
R10414 VPWR.n278 VPWR.t2020 143.911
R10415 VPWR.n266 VPWR.t1937 143.911
R10416 VPWR.n254 VPWR.t1931 143.911
R10417 VPWR.n242 VPWR.t2061 143.911
R10418 VPWR.n230 VPWR.t1979 143.911
R10419 VPWR.n218 VPWR.t1965 143.911
R10420 VPWR.n206 VPWR.t2059 143.911
R10421 VPWR.n194 VPWR.t2011 143.911
R10422 VPWR.n182 VPWR.t2003 143.911
R10423 VPWR.n170 VPWR.t1947 143.911
R10424 VPWR.n1247 VPWR.t1953 143.911
R10425 VPWR.n1169 VPWR.t1980 143.911
R10426 VPWR.n1243 VPWR.t2046 143.911
R10427 VPWR.n1501 VPWR.t1987 143.911
R10428 VPWR.n1189 VPWR.t2040 143.911
R10429 VPWR.n1185 VPWR.t2028 143.911
R10430 VPWR.n1179 VPWR.t1943 143.911
R10431 VPWR.n1495 VPWR.t1999 143.911
R10432 VPWR.n1175 VPWR.t1932 143.911
R10433 VPWR.n1165 VPWR.t2025 143.911
R10434 VPWR.n1488 VPWR.t2049 143.911
R10435 VPWR.n1065 VPWR.t1972 143.911
R10436 VPWR.n1764 VPWR.t2016 143.911
R10437 VPWR.n1052 VPWR.t1962 143.911
R10438 VPWR.n1048 VPWR.t2066 143.911
R10439 VPWR.n1069 VPWR.t2060 143.911
R10440 VPWR.n158 VPWR.t2051 143.911
R10441 VPWR.t1835 VPWR.t317 140.989
R10442 VPWR.t197 VPWR.t370 140.989
R10443 VPWR.t421 VPWR.t197 140.989
R10444 VPWR.t270 VPWR.t421 140.989
R10445 VPWR.t1176 VPWR.t270 140.989
R10446 VPWR.t1110 VPWR.t1176 140.989
R10447 VPWR.t136 VPWR.t1110 140.989
R10448 VPWR.t1166 VPWR.t136 140.989
R10449 VPWR.t874 VPWR.t963 140.989
R10450 VPWR.t371 VPWR.t308 140.989
R10451 VPWR.t279 VPWR.t371 140.989
R10452 VPWR.t698 VPWR.t279 140.989
R10453 VPWR.t80 VPWR.t698 140.989
R10454 VPWR.t90 VPWR.t80 140.989
R10455 VPWR.t82 VPWR.t90 140.989
R10456 VPWR.t84 VPWR.t82 140.989
R10457 VPWR.t464 VPWR.t422 140.989
R10458 VPWR.t202 VPWR.t464 140.989
R10459 VPWR.t282 VPWR.t202 140.989
R10460 VPWR.t130 VPWR.t282 140.989
R10461 VPWR.t124 VPWR.t130 140.989
R10462 VPWR.t132 VPWR.t124 140.989
R10463 VPWR.t134 VPWR.t132 140.989
R10464 VPWR.t614 VPWR.t203 140.989
R10465 VPWR.t312 VPWR.t419 140.989
R10466 VPWR.t374 VPWR.t312 140.989
R10467 VPWR.t205 VPWR.t374 140.989
R10468 VPWR.t657 VPWR.t205 140.989
R10469 VPWR.t1168 VPWR.t657 140.989
R10470 VPWR.t1174 VPWR.t1168 140.989
R10471 VPWR.t1170 VPWR.t1174 140.989
R10472 VPWR.t310 VPWR.t275 140.989
R10473 VPWR.t271 VPWR.t310 140.989
R10474 VPWR.t376 VPWR.t271 140.989
R10475 VPWR.t76 VPWR.t376 140.989
R10476 VPWR.t86 VPWR.t76 140.989
R10477 VPWR.t78 VPWR.t86 140.989
R10478 VPWR.t88 VPWR.t78 140.989
R10479 VPWR.t314 VPWR.t198 140.989
R10480 VPWR.t306 VPWR.t314 140.989
R10481 VPWR.t200 VPWR.t306 140.989
R10482 VPWR.t126 VPWR.t200 140.989
R10483 VPWR.t120 VPWR.t126 140.989
R10484 VPWR.t128 VPWR.t120 140.989
R10485 VPWR.t122 VPWR.t128 140.989
R10486 VPWR VPWR.n1461 133.312
R10487 VPWR.n2799 VPWR 127.562
R10488 VPWR.n2779 VPWR 127.562
R10489 VPWR.n2760 VPWR 127.562
R10490 VPWR VPWR.t466 125.883
R10491 VPWR.n2724 VPWR 125.883
R10492 VPWR.t876 VPWR.t961 120.849
R10493 VPWR.t917 VPWR.t468 117.492
R10494 VPWR.t98 VPWR.t737 117.492
R10495 VPWR.t92 VPWR 115.814
R10496 VPWR VPWR.t1166 114.135
R10497 VPWR VPWR.t84 114.135
R10498 VPWR VPWR.t134 114.135
R10499 VPWR.t490 VPWR 107.421
R10500 VPWR.n1349 VPWR.n1348 106.561
R10501 VPWR.n2800 VPWR.n2799 106.561
R10502 VPWR.n2780 VPWR.n2779 106.561
R10503 VPWR.n2761 VPWR.n2760 106.561
R10504 VPWR.n2725 VPWR.n2724 106.561
R10505 VPWR.n2687 VPWR.n2686 106.561
R10506 VPWR.n2650 VPWR.n2649 106.561
R10507 VPWR VPWR.t880 106.543
R10508 VPWR VPWR.n1253 104.8
R10509 VPWR VPWR.n1276 104.8
R10510 VPWR VPWR.n1300 104.8
R10511 VPWR VPWR.n1385 104.8
R10512 VPWR VPWR.n1424 104.8
R10513 VPWR.n1462 VPWR 100.883
R10514 VPWR VPWR.t626 100.624
R10515 VPWR.n1250 VPWR.n1249 91.8492
R10516 VPWR.n1172 VPWR.n1171 91.8492
R10517 VPWR.n1246 VPWR.n1245 91.8492
R10518 VPWR.n1504 VPWR.n1503 91.8492
R10519 VPWR.n1192 VPWR.n1191 91.8492
R10520 VPWR.n1188 VPWR.n1187 91.8492
R10521 VPWR.n1182 VPWR.n1181 91.8492
R10522 VPWR.n1498 VPWR.n1497 91.8492
R10523 VPWR.n1178 VPWR.n1177 91.8492
R10524 VPWR.n1168 VPWR.n1167 91.8492
R10525 VPWR.n1491 VPWR.n1490 91.8492
R10526 VPWR.n1068 VPWR.n1067 91.8492
R10527 VPWR.n1767 VPWR.n1766 91.8492
R10528 VPWR.n1055 VPWR.n1054 91.8492
R10529 VPWR.n1051 VPWR.n1050 91.8492
R10530 VPWR.n1072 VPWR.n1071 91.8492
R10531 VPWR.t378 VPWR 88.7855
R10532 VPWR.n2855 VPWR.n2853 83.2005
R10533 VPWR.n33 VPWR.n31 83.2005
R10534 VPWR.n2856 VPWR.n24 82.4894
R10535 VPWR.n35 VPWR.n34 82.4894
R10536 VPWR.n2841 VPWR.n35 80.9417
R10537 VPWR.n2853 VPWR.n25 80.9417
R10538 VPWR.n2836 VPWR.n24 80.9417
R10539 VPWR.n2834 VPWR.n31 80.9417
R10540 VPWR.n1254 VPWR 79.407
R10541 VPWR.n1277 VPWR 79.407
R10542 VPWR.n1301 VPWR 79.407
R10543 VPWR.n1386 VPWR 79.407
R10544 VPWR.n1425 VPWR 79.407
R10545 VPWR.t1108 VPWR.t154 78.8874
R10546 VPWR.t263 VPWR.t449 70.4952
R10547 VPWR.t449 VPWR.t265 70.4952
R10548 VPWR.t265 VPWR.t1831 70.4952
R10549 VPWR.t1831 VPWR.t428 70.4952
R10550 VPWR.t428 VPWR.t624 70.4952
R10551 VPWR.t624 VPWR.t1347 70.4952
R10552 VPWR.t1347 VPWR.t1835 70.4952
R10553 VPWR.t195 VPWR.t614 70.4952
R10554 VPWR.t620 VPWR.t195 70.4952
R10555 VPWR.t280 VPWR.t620 70.4952
R10556 VPWR.t856 VPWR.t280 70.4952
R10557 VPWR.t424 VPWR.t856 70.4952
R10558 VPWR.t618 VPWR.t424 70.4952
R10559 VPWR.t466 VPWR.t618 70.4952
R10560 VPWR VPWR.t263 68.8168
R10561 VPWR.t882 VPWR.t878 68.8168
R10562 VPWR.t154 VPWR.t92 62.103
R10563 VPWR VPWR.t874 60.4245
R10564 VPWR.t878 VPWR.t926 52.0323
R10565 VPWR.t299 VPWR 50.3539
R10566 VPWR VPWR.t882 50.3539
R10567 VPWR VPWR.t876 50.3539
R10568 VPWR.t419 VPWR 50.3539
R10569 VPWR.t275 VPWR 50.3539
R10570 VPWR.t198 VPWR 50.3539
R10571 VPWR.n2842 VPWR.n2840 37.0005
R10572 VPWR.n2840 VPWR.n2839 37.0005
R10573 VPWR.n2838 VPWR.n2837 37.0005
R10574 VPWR.n2839 VPWR.n2838 37.0005
R10575 VPWR.n2852 VPWR.n2851 37.0005
R10576 VPWR.n2851 VPWR.n2850 37.0005
R10577 VPWR.n2849 VPWR.n2848 37.0005
R10578 VPWR.n2850 VPWR.n2849 37.0005
R10579 VPWR.n32 VPWR.t1294 34.7652
R10580 VPWR.n32 VPWR.t748 34.7652
R10581 VPWR.n2854 VPWR.t834 34.7652
R10582 VPWR.n2854 VPWR.t978 34.7652
R10583 VPWR.n1249 VPWR.n1248 34.7473
R10584 VPWR.n1171 VPWR.n1170 34.7473
R10585 VPWR.n1245 VPWR.n1244 34.7473
R10586 VPWR.n1503 VPWR.n1502 34.7473
R10587 VPWR.n1191 VPWR.n1190 34.7473
R10588 VPWR.n1187 VPWR.n1186 34.7473
R10589 VPWR.n1181 VPWR.n1180 34.7473
R10590 VPWR.n1497 VPWR.n1496 34.7473
R10591 VPWR.n1177 VPWR.n1176 34.7473
R10592 VPWR.n1167 VPWR.n1166 34.7473
R10593 VPWR.n1490 VPWR.n1489 34.7473
R10594 VPWR.n1067 VPWR.n1066 34.7473
R10595 VPWR.n1766 VPWR.n1765 34.7473
R10596 VPWR.n1054 VPWR.n1053 34.7473
R10597 VPWR.n1050 VPWR.n1049 34.7473
R10598 VPWR.n1071 VPWR.n1070 34.7473
R10599 VPWR.n1318 VPWR.n1317 34.6358
R10600 VPWR.n1376 VPWR.n1360 34.6358
R10601 VPWR.n1381 VPWR.n1380 34.6358
R10602 VPWR.n1415 VPWR.n1399 34.6358
R10603 VPWR.n1420 VPWR.n1419 34.6358
R10604 VPWR.n1430 VPWR.n1396 34.6358
R10605 VPWR.n1452 VPWR.n1436 34.6358
R10606 VPWR.n1457 VPWR.n1456 34.6358
R10607 VPWR.n2774 VPWR.n2773 34.6358
R10608 VPWR.n2740 VPWR.n2732 34.6358
R10609 VPWR.n2747 VPWR.n2746 34.6358
R10610 VPWR.n2704 VPWR.n2695 34.6358
R10611 VPWR.n2707 VPWR.n2706 34.6358
R10612 VPWR.n2711 VPWR.n2710 34.6358
R10613 VPWR.n2667 VPWR.n2658 34.6358
R10614 VPWR.n2670 VPWR.n2669 34.6358
R10615 VPWR.n2674 VPWR.n2673 34.6358
R10616 VPWR.n2681 VPWR.n2680 34.6358
R10617 VPWR.n2634 VPWR.n2630 34.6358
R10618 VPWR.n2638 VPWR.n2622 34.6358
R10619 VPWR.n2641 VPWR.n2640 34.6358
R10620 VPWR.n1335 VPWR.n1334 32.0005
R10621 VPWR.n1372 VPWR.n1371 32.0005
R10622 VPWR.n1411 VPWR.n1410 32.0005
R10623 VPWR.n1448 VPWR.n1447 32.0005
R10624 VPWR.n2736 VPWR.n2735 30.8711
R10625 VPWR.n2700 VPWR.n2699 30.8711
R10626 VPWR.n2663 VPWR.n2662 30.8711
R10627 VPWR.n2629 VPWR.n2628 30.8711
R10628 VPWR.n1344 VPWR.n1343 28.2358
R10629 VPWR.n5 VPWR.t1834 26.5955
R10630 VPWR.n5 VPWR.t623 26.5955
R10631 VPWR.n4 VPWR.t627 26.5955
R10632 VPWR.n4 VPWR.t1830 26.5955
R10633 VPWR.n1259 VPWR.t106 26.5955
R10634 VPWR.n1259 VPWR.t105 26.5955
R10635 VPWR.n1258 VPWR.t36 26.5955
R10636 VPWR.n1258 VPWR.t29 26.5955
R10637 VPWR.n1264 VPWR.t101 26.5955
R10638 VPWR.n1264 VPWR.t107 26.5955
R10639 VPWR.n1257 VPWR.t32 26.5955
R10640 VPWR.n1257 VPWR.t35 26.5955
R10641 VPWR.n1282 VPWR.t208 26.5955
R10642 VPWR.n1282 VPWR.t209 26.5955
R10643 VPWR.n1281 VPWR.t162 26.5955
R10644 VPWR.n1281 VPWR.t159 26.5955
R10645 VPWR.n1287 VPWR.t1107 26.5955
R10646 VPWR.n1287 VPWR.t660 26.5955
R10647 VPWR.n1280 VPWR.t165 26.5955
R10648 VPWR.n1280 VPWR.t163 26.5955
R10649 VPWR.n1306 VPWR.t762 26.5955
R10650 VPWR.n1306 VPWR.t769 26.5955
R10651 VPWR.n1305 VPWR.t116 26.5955
R10652 VPWR.n1305 VPWR.t115 26.5955
R10653 VPWR.n1311 VPWR.t766 26.5955
R10654 VPWR.n1311 VPWR.t763 26.5955
R10655 VPWR.n1304 VPWR.t119 26.5955
R10656 VPWR.n1304 VPWR.t117 26.5955
R10657 VPWR.n1333 VPWR.t320 26.5955
R10658 VPWR.n1333 VPWR.t473 26.5955
R10659 VPWR.n1326 VPWR.t1836 26.5955
R10660 VPWR.n1326 VPWR.t318 26.5955
R10661 VPWR.n1340 VPWR.t1832 26.5955
R10662 VPWR.n1340 VPWR.t625 26.5955
R10663 VPWR.n1342 VPWR.t266 26.5955
R10664 VPWR.n1342 VPWR.t429 26.5955
R10665 VPWR.n1370 VPWR.t894 26.5955
R10666 VPWR.n1370 VPWR.t277 26.5955
R10667 VPWR.n1369 VPWR.t260 26.5955
R10668 VPWR.n1369 VPWR.t1367 26.5955
R10669 VPWR.n1363 VPWR.t109 26.5955
R10670 VPWR.n1363 VPWR.t889 26.5955
R10671 VPWR.n1362 VPWR.t33 26.5955
R10672 VPWR.n1362 VPWR.t403 26.5955
R10673 VPWR.n1378 VPWR.t104 26.5955
R10674 VPWR.n1378 VPWR.t103 26.5955
R10675 VPWR.n1377 VPWR.t31 26.5955
R10676 VPWR.n1377 VPWR.t34 26.5955
R10677 VPWR.n1409 VPWR.t402 26.5955
R10678 VPWR.n1409 VPWR.t262 26.5955
R10679 VPWR.n1408 VPWR.t896 26.5955
R10680 VPWR.n1408 VPWR.t278 26.5955
R10681 VPWR.n1402 VPWR.t1105 26.5955
R10682 VPWR.n1402 VPWR.t475 26.5955
R10683 VPWR.n1401 VPWR.t166 26.5955
R10684 VPWR.n1401 VPWR.t892 26.5955
R10685 VPWR.n1417 VPWR.t211 26.5955
R10686 VPWR.n1417 VPWR.t1106 26.5955
R10687 VPWR.n1416 VPWR.t167 26.5955
R10688 VPWR.n1416 VPWR.t164 26.5955
R10689 VPWR.n1446 VPWR.t1372 26.5955
R10690 VPWR.n1446 VPWR.t268 26.5955
R10691 VPWR.n1445 VPWR.t261 26.5955
R10692 VPWR.n1445 VPWR.t1368 26.5955
R10693 VPWR.n1439 VPWR.t765 26.5955
R10694 VPWR.n1439 VPWR.t1369 26.5955
R10695 VPWR.n1438 VPWR.t112 26.5955
R10696 VPWR.n1438 VPWR.t404 26.5955
R10697 VPWR.n1454 VPWR.t768 26.5955
R10698 VPWR.n1454 VPWR.t767 26.5955
R10699 VPWR.n1453 VPWR.t113 26.5955
R10700 VPWR.n1453 VPWR.t111 26.5955
R10701 VPWR.n2821 VPWR.t855 26.5955
R10702 VPWR.n2821 VPWR.t176 26.5955
R10703 VPWR.n2823 VPWR.t617 26.5955
R10704 VPWR.n2823 VPWR.t1131 26.5955
R10705 VPWR.n2801 VPWR.t1177 26.5955
R10706 VPWR.n2801 VPWR.t1172 26.5955
R10707 VPWR.n2802 VPWR.t1888 26.5955
R10708 VPWR.n2802 VPWR.t1111 26.5955
R10709 VPWR.n2805 VPWR.t1165 26.5955
R10710 VPWR.n2805 VPWR.t1167 26.5955
R10711 VPWR.n2806 VPWR.t137 26.5955
R10712 VPWR.n2806 VPWR.t1924 26.5955
R10713 VPWR.n2781 VPWR.t81 26.5955
R10714 VPWR.n2781 VPWR.t91 26.5955
R10715 VPWR.n2782 VPWR.t1891 26.5955
R10716 VPWR.n2782 VPWR.t1897 26.5955
R10717 VPWR.n2785 VPWR.t83 26.5955
R10718 VPWR.n2785 VPWR.t85 26.5955
R10719 VPWR.n2786 VPWR.t1893 26.5955
R10720 VPWR.n2786 VPWR.t1895 26.5955
R10721 VPWR.n2762 VPWR.t131 26.5955
R10722 VPWR.n2762 VPWR.t125 26.5955
R10723 VPWR.n2763 VPWR.t944 26.5955
R10724 VPWR.n2763 VPWR.t943 26.5955
R10725 VPWR.n2766 VPWR.t133 26.5955
R10726 VPWR.n2766 VPWR.t135 26.5955
R10727 VPWR.n2767 VPWR.t946 26.5955
R10728 VPWR.n2767 VPWR.t940 26.5955
R10729 VPWR.n2727 VPWR.t281 26.5955
R10730 VPWR.n2727 VPWR.t425 26.5955
R10731 VPWR.n2731 VPWR.t204 26.5955
R10732 VPWR.n2731 VPWR.t615 26.5955
R10733 VPWR.n2734 VPWR.t284 26.5955
R10734 VPWR.n2734 VPWR.t373 26.5955
R10735 VPWR.n2728 VPWR.t621 26.5955
R10736 VPWR.n2728 VPWR.t857 26.5955
R10737 VPWR.n2698 VPWR.t1856 26.5955
R10738 VPWR.n2698 VPWR.t375 26.5955
R10739 VPWR.n2697 VPWR.t313 26.5955
R10740 VPWR.n2697 VPWR.t465 26.5955
R10741 VPWR.n2694 VPWR.t206 26.5955
R10742 VPWR.n2694 VPWR.t658 26.5955
R10743 VPWR.n2693 VPWR.t380 26.5955
R10744 VPWR.n2693 VPWR.t1173 26.5955
R10745 VPWR.n2690 VPWR.t1923 26.5955
R10746 VPWR.n2690 VPWR.t1319 26.5955
R10747 VPWR.n2689 VPWR.t1169 26.5955
R10748 VPWR.n2689 VPWR.t1175 26.5955
R10749 VPWR.n2661 VPWR.t311 26.5955
R10750 VPWR.n2661 VPWR.t1858 26.5955
R10751 VPWR.n2660 VPWR.t423 26.5955
R10752 VPWR.n2660 VPWR.t272 26.5955
R10753 VPWR.n2657 VPWR.t377 26.5955
R10754 VPWR.n2657 VPWR.t1896 26.5955
R10755 VPWR.n2656 VPWR.t694 26.5955
R10756 VPWR.n2656 VPWR.t77 26.5955
R10757 VPWR.n2653 VPWR.t1892 26.5955
R10758 VPWR.n2653 VPWR.t1898 26.5955
R10759 VPWR.n2652 VPWR.t87 26.5955
R10760 VPWR.n2652 VPWR.t79 26.5955
R10761 VPWR.n2625 VPWR.t315 26.5955
R10762 VPWR.n2625 VPWR.t307 26.5955
R10763 VPWR.n2624 VPWR.t697 26.5955
R10764 VPWR.n2624 VPWR.t426 26.5955
R10765 VPWR.n2632 VPWR.t201 26.5955
R10766 VPWR.n2632 VPWR.t945 26.5955
R10767 VPWR.n2631 VPWR.t273 26.5955
R10768 VPWR.n2631 VPWR.t127 26.5955
R10769 VPWR.n2621 VPWR.t947 26.5955
R10770 VPWR.n2621 VPWR.t941 26.5955
R10771 VPWR.n2620 VPWR.t121 26.5955
R10772 VPWR.n2620 VPWR.t129 26.5955
R10773 VPWR.n17 VPWR.n16 25.977
R10774 VPWR.n1272 VPWR.n1271 25.977
R10775 VPWR.n1332 VPWR.n1329 25.977
R10776 VPWR.n1368 VPWR.n1365 25.977
R10777 VPWR.n1391 VPWR.n1357 25.977
R10778 VPWR.n1407 VPWR.n1404 25.977
R10779 VPWR.n1444 VPWR.n1441 25.977
R10780 VPWR.n2830 VPWR.n2829 25.977
R10781 VPWR.n2814 VPWR.n2813 25.977
R10782 VPWR.n2736 VPWR.n2733 25.977
R10783 VPWR.n2700 VPWR.n2696 25.977
R10784 VPWR.n2718 VPWR.n2717 25.977
R10785 VPWR.n2663 VPWR.n2659 25.977
R10786 VPWR.n2628 VPWR.n2626 25.977
R10787 VPWR.n1354 VPWR.n1353 25.224
R10788 VPWR.n2756 VPWR.n2755 25.224
R10789 VPWR.n2741 VPWR.n2740 24.8476
R10790 VPWR.n2705 VPWR.n2704 24.8476
R10791 VPWR.n2668 VPWR.n2667 24.8476
R10792 VPWR.n2634 VPWR.n2633 24.8476
R10793 VPWR.n16 VPWR.n15 24.4711
R10794 VPWR.n1271 VPWR.n1270 24.4711
R10795 VPWR.n1334 VPWR.n1332 24.4711
R10796 VPWR.n1371 VPWR.n1368 24.4711
R10797 VPWR.n1410 VPWR.n1407 24.4711
R10798 VPWR.n1447 VPWR.n1444 24.4711
R10799 VPWR.n2829 VPWR.n2828 24.4711
R10800 VPWR.n2813 VPWR.n2812 24.4711
R10801 VPWR.n11 VPWR.n2 23.7181
R10802 VPWR.n1266 VPWR.n1255 23.7181
R10803 VPWR.n1289 VPWR.n1278 23.7181
R10804 VPWR.n1293 VPWR.n1278 23.7181
R10805 VPWR.n1313 VPWR.n1302 23.7181
R10806 VPWR.n1317 VPWR.n1302 23.7181
R10807 VPWR.n1349 VPWR.n1347 23.7181
R10808 VPWR.n1387 VPWR.n1384 23.7181
R10809 VPWR.n1426 VPWR.n1423 23.7181
R10810 VPWR.n1426 VPWR.n1396 23.7181
R10811 VPWR.n1463 VPWR.n1460 23.7181
R10812 VPWR.n2827 VPWR.n2826 23.7181
R10813 VPWR.n2808 VPWR.n2800 23.7181
R10814 VPWR.n2788 VPWR.n2780 23.7181
R10815 VPWR.n2792 VPWR.n2780 23.7181
R10816 VPWR.n2769 VPWR.n2761 23.7181
R10817 VPWR.n2773 VPWR.n2761 23.7181
R10818 VPWR.n2750 VPWR.n2725 23.7181
R10819 VPWR.n2713 VPWR.n2687 23.7181
R10820 VPWR.n2676 VPWR.n2650 23.7181
R10821 VPWR.n2680 VPWR.n2650 23.7181
R10822 VPWR.n2645 VPWR.n2644 23.7181
R10823 VPWR.t470 VPWR.t917 23.4987
R10824 VPWR.t739 VPWR.t98 23.4987
R10825 VPWR.n11 VPWR.n10 22.9652
R10826 VPWR.n1266 VPWR.n1265 22.9652
R10827 VPWR.n1289 VPWR.n1288 22.9652
R10828 VPWR.n1313 VPWR.n1312 22.9652
R10829 VPWR.n2826 VPWR.n2822 22.9652
R10830 VPWR.n2808 VPWR.n2807 22.9652
R10831 VPWR.n2788 VPWR.n2787 22.9652
R10832 VPWR.n2769 VPWR.n2768 22.9652
R10833 VPWR.n1339 VPWR.n1327 22.2123
R10834 VPWR.n2743 VPWR.n2742 22.2123
R10835 VPWR.n10 VPWR.n3 21.4593
R10836 VPWR.n1265 VPWR.n1256 21.4593
R10837 VPWR.n1288 VPWR.n1279 21.4593
R10838 VPWR.n1312 VPWR.n1303 21.4593
R10839 VPWR.n1461 VPWR.t110 20.5957
R10840 VPWR.n1462 VPWR.t267 20.5957
R10841 VPWR.n1296 VPWR.n1295 19.9534
R10842 VPWR.n1319 VPWR.n1318 19.9534
R10843 VPWR.n1353 VPWR.n1322 19.9534
R10844 VPWR.n2795 VPWR.n2794 19.9534
R10845 VPWR.n2775 VPWR.n2774 19.9534
R10846 VPWR.n2755 VPWR.n2754 19.9534
R10847 VPWR.n2743 VPWR.n2729 18.824
R10848 VPWR.n2707 VPWR.n2691 18.824
R10849 VPWR.n2670 VPWR.n2654 18.824
R10850 VPWR.n2639 VPWR.n2638 18.824
R10851 VPWR.n1335 VPWR.n1327 18.4476
R10852 VPWR.n1372 VPWR.n1364 18.4476
R10853 VPWR.n1392 VPWR.n1391 18.4476
R10854 VPWR.n1411 VPWR.n1403 18.4476
R10855 VPWR.n1448 VPWR.n1440 18.4476
R10856 VPWR.n2719 VPWR.n2718 18.4476
R10857 VPWR.n1432 VPWR.n1431 17.5829
R10858 VPWR.n2683 VPWR.n2682 17.5829
R10859 VPWR.n6 VPWR.n3 16.9417
R10860 VPWR.n1260 VPWR.n1256 16.9417
R10861 VPWR.n1283 VPWR.n1279 16.9417
R10862 VPWR.n1307 VPWR.n1303 16.9417
R10863 VPWR.n2749 VPWR.n2748 16.5652
R10864 VPWR.n1325 VPWR.n1323 16.1887
R10865 VPWR.n1393 VPWR.n1392 16.1887
R10866 VPWR.n2720 VPWR.n2719 16.1887
R10867 VPWR.n1254 VPWR.t100 16.0935
R10868 VPWR.n1277 VPWR.t207 16.0935
R10869 VPWR.n1301 VPWR.t316 16.0935
R10870 VPWR.n1386 VPWR.t102 16.0935
R10871 VPWR.n1425 VPWR.t210 16.0935
R10872 VPWR.n1253 VPWR.t28 16.0935
R10873 VPWR.n1276 VPWR.t158 16.0935
R10874 VPWR.n1300 VPWR.t114 16.0935
R10875 VPWR.n1385 VPWR.t30 16.0935
R10876 VPWR.n1424 VPWR.t160 16.0935
R10877 VPWR.n1344 VPWR.n1325 15.8123
R10878 VPWR.n2746 VPWR.n2729 15.8123
R10879 VPWR.n2748 VPWR.n2747 15.8123
R10880 VPWR.n2710 VPWR.n2691 15.8123
R10881 VPWR.n2673 VPWR.n2654 15.8123
R10882 VPWR.n2640 VPWR.n2639 15.8123
R10883 VPWR.n1349 VPWR.n1322 13.5534
R10884 VPWR.n2754 VPWR.n2725 13.5534
R10885 VPWR.n15 VPWR.n2 12.8005
R10886 VPWR.n1270 VPWR.n1255 12.8005
R10887 VPWR.n1387 VPWR.n1357 12.8005
R10888 VPWR.n2828 VPWR.n2827 12.8005
R10889 VPWR.n2812 VPWR.n2800 12.8005
R10890 VPWR.n2717 VPWR.n2687 12.8005
R10891 VPWR.n1341 VPWR.n1339 12.424
R10892 VPWR.n1379 VPWR.n1376 12.424
R10893 VPWR.n1418 VPWR.n1415 12.424
R10894 VPWR.n1455 VPWR.n1452 12.424
R10895 VPWR.n1295 VPWR.n1294 10.5417
R10896 VPWR.n1431 VPWR.n1430 10.5417
R10897 VPWR.n2794 VPWR.n2793 10.5417
R10898 VPWR.n2682 VPWR.n2681 10.5417
R10899 VPWR.n2706 VPWR.n2705 9.78874
R10900 VPWR.n2669 VPWR.n2668 9.78874
R10901 VPWR.n2633 VPWR.n2622 9.78874
R10902 VPWR.n1380 VPWR.n1379 9.41227
R10903 VPWR.n1384 VPWR.n1358 9.41227
R10904 VPWR.n1419 VPWR.n1418 9.41227
R10905 VPWR.n1423 VPWR.n1397 9.41227
R10906 VPWR.n1456 VPWR.n1455 9.41227
R10907 VPWR.n1460 VPWR.n1434 9.41227
R10908 VPWR.n2713 VPWR.n2712 9.41227
R10909 VPWR.n2676 VPWR.n2675 9.41227
R10910 VPWR.n2644 VPWR.n2618 9.41227
R10911 VPWR.n1248 VPWR 9.37021
R10912 VPWR.n1170 VPWR 9.37021
R10913 VPWR.n1244 VPWR 9.37021
R10914 VPWR.n1502 VPWR 9.37021
R10915 VPWR.n1190 VPWR 9.37021
R10916 VPWR.n1186 VPWR 9.37021
R10917 VPWR.n1180 VPWR 9.37021
R10918 VPWR.n1496 VPWR 9.37021
R10919 VPWR.n1176 VPWR 9.37021
R10920 VPWR.n1166 VPWR 9.37021
R10921 VPWR.n1489 VPWR 9.37021
R10922 VPWR.n1066 VPWR 9.37021
R10923 VPWR.n1765 VPWR 9.37021
R10924 VPWR.n1053 VPWR 9.37021
R10925 VPWR.n1049 VPWR 9.37021
R10926 VPWR.n1070 VPWR 9.37021
R10927 VPWR.n1486 VPWR.n1485 9.33404
R10928 VPWR.n371 VPWR.n370 9.33404
R10929 VPWR.n1553 VPWR.n1552 9.33404
R10930 VPWR.n367 VPWR.n366 9.33404
R10931 VPWR.n984 VPWR.n983 9.33404
R10932 VPWR.n2498 VPWR.n2497 9.33404
R10933 VPWR.n2494 VPWR.n2493 9.33404
R10934 VPWR.n339 VPWR.n338 9.33404
R10935 VPWR.n992 VPWR.n991 9.33404
R10936 VPWR.n2464 VPWR.n2463 9.33404
R10937 VPWR.n343 VPWR.n342 9.33404
R10938 VPWR.n1910 VPWR.n1909 9.33404
R10939 VPWR.n1906 VPWR.n1905 9.33404
R10940 VPWR.n1900 VPWR.n1899 9.33404
R10941 VPWR.n408 VPWR.n407 9.33404
R10942 VPWR.n412 VPWR.n411 9.33404
R10943 VPWR.n416 VPWR.n415 9.33404
R10944 VPWR.n2474 VPWR.n2473 9.33404
R10945 VPWR.n351 VPWR.n350 9.33404
R10946 VPWR.n1896 VPWR.n1895 9.33404
R10947 VPWR.n424 VPWR.n423 9.33404
R10948 VPWR.n2478 VPWR.n2477 9.33404
R10949 VPWR.n355 VPWR.n354 9.33404
R10950 VPWR.n2327 VPWR.n2326 9.33404
R10951 VPWR.n2331 VPWR.n2330 9.33404
R10952 VPWR.n2337 VPWR.n2336 9.33404
R10953 VPWR.n2341 VPWR.n2340 9.33404
R10954 VPWR.n2351 VPWR.n2350 9.33404
R10955 VPWR.n2357 VPWR.n2356 9.33404
R10956 VPWR.n2361 VPWR.n2360 9.33404
R10957 VPWR.n2367 VPWR.n2366 9.33404
R10958 VPWR.n2371 VPWR.n2370 9.33404
R10959 VPWR.n2377 VPWR.n2376 9.33404
R10960 VPWR.n2381 VPWR.n2380 9.33404
R10961 VPWR.n2387 VPWR.n2386 9.33404
R10962 VPWR.n2391 VPWR.n2390 9.33404
R10963 VPWR.n2397 VPWR.n2396 9.33404
R10964 VPWR.n2400 VPWR.n2399 9.33404
R10965 VPWR.n2347 VPWR.n2346 9.33404
R10966 VPWR.n563 VPWR.n562 9.33404
R10967 VPWR.n559 VPWR.n558 9.33404
R10968 VPWR.n555 VPWR.n554 9.33404
R10969 VPWR.n551 VPWR.n550 9.33404
R10970 VPWR.n543 VPWR.n542 9.33404
R10971 VPWR.n539 VPWR.n538 9.33404
R10972 VPWR.n535 VPWR.n534 9.33404
R10973 VPWR.n531 VPWR.n530 9.33404
R10974 VPWR.n527 VPWR.n526 9.33404
R10975 VPWR.n523 VPWR.n522 9.33404
R10976 VPWR.n519 VPWR.n518 9.33404
R10977 VPWR.n515 VPWR.n514 9.33404
R10978 VPWR.n511 VPWR.n510 9.33404
R10979 VPWR.n507 VPWR.n506 9.33404
R10980 VPWR.n504 VPWR.n503 9.33404
R10981 VPWR.n547 VPWR.n546 9.33404
R10982 VPWR.n2302 VPWR.n2301 9.33404
R10983 VPWR.n2298 VPWR.n2297 9.33404
R10984 VPWR.n2292 VPWR.n2291 9.33404
R10985 VPWR.n2288 VPWR.n2287 9.33404
R10986 VPWR.n2278 VPWR.n2277 9.33404
R10987 VPWR.n2272 VPWR.n2271 9.33404
R10988 VPWR.n2268 VPWR.n2267 9.33404
R10989 VPWR.n2262 VPWR.n2261 9.33404
R10990 VPWR.n2258 VPWR.n2257 9.33404
R10991 VPWR.n2252 VPWR.n2251 9.33404
R10992 VPWR.n2248 VPWR.n2247 9.33404
R10993 VPWR.n2242 VPWR.n2241 9.33404
R10994 VPWR.n2238 VPWR.n2237 9.33404
R10995 VPWR.n2232 VPWR.n2231 9.33404
R10996 VPWR.n2229 VPWR.n2228 9.33404
R10997 VPWR.n2282 VPWR.n2281 9.33404
R10998 VPWR.n600 VPWR.n599 9.33404
R10999 VPWR.n604 VPWR.n603 9.33404
R11000 VPWR.n608 VPWR.n607 9.33404
R11001 VPWR.n612 VPWR.n611 9.33404
R11002 VPWR.n620 VPWR.n619 9.33404
R11003 VPWR.n624 VPWR.n623 9.33404
R11004 VPWR.n628 VPWR.n627 9.33404
R11005 VPWR.n632 VPWR.n631 9.33404
R11006 VPWR.n636 VPWR.n635 9.33404
R11007 VPWR.n640 VPWR.n639 9.33404
R11008 VPWR.n644 VPWR.n643 9.33404
R11009 VPWR.n648 VPWR.n647 9.33404
R11010 VPWR.n652 VPWR.n651 9.33404
R11011 VPWR.n656 VPWR.n655 9.33404
R11012 VPWR.n659 VPWR.n658 9.33404
R11013 VPWR.n616 VPWR.n615 9.33404
R11014 VPWR.n2131 VPWR.n2130 9.33404
R11015 VPWR.n2135 VPWR.n2134 9.33404
R11016 VPWR.n2141 VPWR.n2140 9.33404
R11017 VPWR.n2145 VPWR.n2144 9.33404
R11018 VPWR.n2155 VPWR.n2154 9.33404
R11019 VPWR.n2161 VPWR.n2160 9.33404
R11020 VPWR.n2165 VPWR.n2164 9.33404
R11021 VPWR.n2171 VPWR.n2170 9.33404
R11022 VPWR.n2175 VPWR.n2174 9.33404
R11023 VPWR.n2181 VPWR.n2180 9.33404
R11024 VPWR.n2185 VPWR.n2184 9.33404
R11025 VPWR.n2191 VPWR.n2190 9.33404
R11026 VPWR.n2195 VPWR.n2194 9.33404
R11027 VPWR.n2201 VPWR.n2200 9.33404
R11028 VPWR.n2204 VPWR.n2203 9.33404
R11029 VPWR.n2151 VPWR.n2150 9.33404
R11030 VPWR.n755 VPWR.n754 9.33404
R11031 VPWR.n751 VPWR.n750 9.33404
R11032 VPWR.n747 VPWR.n746 9.33404
R11033 VPWR.n743 VPWR.n742 9.33404
R11034 VPWR.n735 VPWR.n734 9.33404
R11035 VPWR.n731 VPWR.n730 9.33404
R11036 VPWR.n727 VPWR.n726 9.33404
R11037 VPWR.n723 VPWR.n722 9.33404
R11038 VPWR.n719 VPWR.n718 9.33404
R11039 VPWR.n715 VPWR.n714 9.33404
R11040 VPWR.n711 VPWR.n710 9.33404
R11041 VPWR.n707 VPWR.n706 9.33404
R11042 VPWR.n703 VPWR.n702 9.33404
R11043 VPWR.n699 VPWR.n698 9.33404
R11044 VPWR.n696 VPWR.n695 9.33404
R11045 VPWR.n739 VPWR.n738 9.33404
R11046 VPWR.n2106 VPWR.n2105 9.33404
R11047 VPWR.n2102 VPWR.n2101 9.33404
R11048 VPWR.n2096 VPWR.n2095 9.33404
R11049 VPWR.n2092 VPWR.n2091 9.33404
R11050 VPWR.n2082 VPWR.n2081 9.33404
R11051 VPWR.n2076 VPWR.n2075 9.33404
R11052 VPWR.n2072 VPWR.n2071 9.33404
R11053 VPWR.n2066 VPWR.n2065 9.33404
R11054 VPWR.n2062 VPWR.n2061 9.33404
R11055 VPWR.n2056 VPWR.n2055 9.33404
R11056 VPWR.n2052 VPWR.n2051 9.33404
R11057 VPWR.n2046 VPWR.n2045 9.33404
R11058 VPWR.n2042 VPWR.n2041 9.33404
R11059 VPWR.n2036 VPWR.n2035 9.33404
R11060 VPWR.n2033 VPWR.n2032 9.33404
R11061 VPWR.n2086 VPWR.n2085 9.33404
R11062 VPWR.n792 VPWR.n791 9.33404
R11063 VPWR.n796 VPWR.n795 9.33404
R11064 VPWR.n800 VPWR.n799 9.33404
R11065 VPWR.n804 VPWR.n803 9.33404
R11066 VPWR.n812 VPWR.n811 9.33404
R11067 VPWR.n816 VPWR.n815 9.33404
R11068 VPWR.n820 VPWR.n819 9.33404
R11069 VPWR.n824 VPWR.n823 9.33404
R11070 VPWR.n828 VPWR.n827 9.33404
R11071 VPWR.n832 VPWR.n831 9.33404
R11072 VPWR.n836 VPWR.n835 9.33404
R11073 VPWR.n840 VPWR.n839 9.33404
R11074 VPWR.n844 VPWR.n843 9.33404
R11075 VPWR.n848 VPWR.n847 9.33404
R11076 VPWR.n851 VPWR.n850 9.33404
R11077 VPWR.n808 VPWR.n807 9.33404
R11078 VPWR.n1935 VPWR.n1934 9.33404
R11079 VPWR.n1939 VPWR.n1938 9.33404
R11080 VPWR.n1945 VPWR.n1944 9.33404
R11081 VPWR.n1949 VPWR.n1948 9.33404
R11082 VPWR.n1959 VPWR.n1958 9.33404
R11083 VPWR.n1965 VPWR.n1964 9.33404
R11084 VPWR.n1969 VPWR.n1968 9.33404
R11085 VPWR.n1975 VPWR.n1974 9.33404
R11086 VPWR.n1979 VPWR.n1978 9.33404
R11087 VPWR.n1985 VPWR.n1984 9.33404
R11088 VPWR.n1989 VPWR.n1988 9.33404
R11089 VPWR.n1995 VPWR.n1994 9.33404
R11090 VPWR.n1999 VPWR.n1998 9.33404
R11091 VPWR.n2005 VPWR.n2004 9.33404
R11092 VPWR.n2008 VPWR.n2007 9.33404
R11093 VPWR.n1955 VPWR.n1954 9.33404
R11094 VPWR.n947 VPWR.n946 9.33404
R11095 VPWR.n943 VPWR.n942 9.33404
R11096 VPWR.n939 VPWR.n938 9.33404
R11097 VPWR.n935 VPWR.n934 9.33404
R11098 VPWR.n927 VPWR.n926 9.33404
R11099 VPWR.n923 VPWR.n922 9.33404
R11100 VPWR.n919 VPWR.n918 9.33404
R11101 VPWR.n915 VPWR.n914 9.33404
R11102 VPWR.n911 VPWR.n910 9.33404
R11103 VPWR.n907 VPWR.n906 9.33404
R11104 VPWR.n903 VPWR.n902 9.33404
R11105 VPWR.n899 VPWR.n898 9.33404
R11106 VPWR.n895 VPWR.n894 9.33404
R11107 VPWR.n891 VPWR.n890 9.33404
R11108 VPWR.n888 VPWR.n887 9.33404
R11109 VPWR.n931 VPWR.n930 9.33404
R11110 VPWR.n1890 VPWR.n1889 9.33404
R11111 VPWR.n1000 VPWR.n999 9.33404
R11112 VPWR.n1514 VPWR.n1513 9.33404
R11113 VPWR.n420 VPWR.n419 9.33404
R11114 VPWR.n2484 VPWR.n2483 9.33404
R11115 VPWR.n359 VPWR.n358 9.33404
R11116 VPWR.n996 VPWR.n995 9.33404
R11117 VPWR.n1510 VPWR.n1509 9.33404
R11118 VPWR.n1886 VPWR.n1885 9.33404
R11119 VPWR.n1004 VPWR.n1003 9.33404
R11120 VPWR.n1524 VPWR.n1523 9.33404
R11121 VPWR.n428 VPWR.n427 9.33404
R11122 VPWR.n436 VPWR.n435 9.33404
R11123 VPWR.n440 VPWR.n439 9.33404
R11124 VPWR.n444 VPWR.n443 9.33404
R11125 VPWR.n448 VPWR.n447 9.33404
R11126 VPWR.n452 VPWR.n451 9.33404
R11127 VPWR.n456 VPWR.n455 9.33404
R11128 VPWR.n460 VPWR.n459 9.33404
R11129 VPWR.n464 VPWR.n463 9.33404
R11130 VPWR.n467 VPWR.n466 9.33404
R11131 VPWR.n432 VPWR.n431 9.33404
R11132 VPWR.n2468 VPWR.n2467 9.33404
R11133 VPWR.n347 VPWR.n346 9.33404
R11134 VPWR.n1008 VPWR.n1007 9.33404
R11135 VPWR.n1528 VPWR.n1527 9.33404
R11136 VPWR.n1880 VPWR.n1879 9.33404
R11137 VPWR.n1870 VPWR.n1869 9.33404
R11138 VPWR.n1866 VPWR.n1865 9.33404
R11139 VPWR.n1860 VPWR.n1859 9.33404
R11140 VPWR.n1856 VPWR.n1855 9.33404
R11141 VPWR.n1850 VPWR.n1849 9.33404
R11142 VPWR.n1846 VPWR.n1845 9.33404
R11143 VPWR.n1840 VPWR.n1839 9.33404
R11144 VPWR.n1837 VPWR.n1836 9.33404
R11145 VPWR.n1876 VPWR.n1875 9.33404
R11146 VPWR.n1012 VPWR.n1011 9.33404
R11147 VPWR.n1538 VPWR.n1537 9.33404
R11148 VPWR.n2488 VPWR.n2487 9.33404
R11149 VPWR.n363 VPWR.n362 9.33404
R11150 VPWR.n1499 VPWR.n1149 9.33404
R11151 VPWR.n1016 VPWR.n1015 9.33404
R11152 VPWR.n1542 VPWR.n1541 9.33404
R11153 VPWR.n2458 VPWR.n2457 9.33404
R11154 VPWR.n2448 VPWR.n2447 9.33404
R11155 VPWR.n2444 VPWR.n2443 9.33404
R11156 VPWR.n2438 VPWR.n2437 9.33404
R11157 VPWR.n2434 VPWR.n2433 9.33404
R11158 VPWR.n2428 VPWR.n2427 9.33404
R11159 VPWR.n2425 VPWR.n2424 9.33404
R11160 VPWR.n2454 VPWR.n2453 9.33404
R11161 VPWR.n335 VPWR.n334 9.33404
R11162 VPWR.n1557 VPWR.n1556 9.33404
R11163 VPWR.n1020 VPWR.n1019 9.33404
R11164 VPWR.n1024 VPWR.n1023 9.33404
R11165 VPWR.n1028 VPWR.n1027 9.33404
R11166 VPWR.n1032 VPWR.n1031 9.33404
R11167 VPWR.n1036 VPWR.n1035 9.33404
R11168 VPWR.n1040 VPWR.n1039 9.33404
R11169 VPWR.n1043 VPWR.n1042 9.33404
R11170 VPWR.n988 VPWR.n987 9.33404
R11171 VPWR.n1493 VPWR.n1492 9.33404
R11172 VPWR.n331 VPWR.n330 9.33404
R11173 VPWR.n1782 VPWR.n1781 9.33404
R11174 VPWR.n327 VPWR.n326 9.33404
R11175 VPWR.n323 VPWR.n322 9.33404
R11176 VPWR.n315 VPWR.n314 9.33404
R11177 VPWR.n312 VPWR.n311 9.33404
R11178 VPWR.n319 VPWR.n318 9.33404
R11179 VPWR.n1770 VPWR.n1769 9.33404
R11180 VPWR.n1809 VPWR.n1808 9.33404
R11181 VPWR.n1812 VPWR.n1811 9.33404
R11182 VPWR.n1778 VPWR.n1777 9.33404
R11183 VPWR.n2733 VPWR 9.32394
R11184 VPWR.n2696 VPWR 9.32394
R11185 VPWR.n2659 VPWR 9.32394
R11186 VPWR VPWR.n2626 9.32394
R11187 VPWR.n18 VPWR.n17 9.3005
R11188 VPWR.n15 VPWR.n14 9.3005
R11189 VPWR.n13 VPWR.n2 9.3005
R11190 VPWR.n10 VPWR.n9 9.3005
R11191 VPWR.n8 VPWR.n3 9.3005
R11192 VPWR.n12 VPWR.n11 9.3005
R11193 VPWR.n16 VPWR.n0 9.3005
R11194 VPWR.n1273 VPWR.n1272 9.3005
R11195 VPWR.n1270 VPWR.n1269 9.3005
R11196 VPWR.n1268 VPWR.n1255 9.3005
R11197 VPWR.n1265 VPWR.n1263 9.3005
R11198 VPWR.n1262 VPWR.n1256 9.3005
R11199 VPWR.n1267 VPWR.n1266 9.3005
R11200 VPWR.n1271 VPWR.n1252 9.3005
R11201 VPWR.n1297 VPWR.n1296 9.3005
R11202 VPWR.n1291 VPWR.n1278 9.3005
R11203 VPWR.n1288 VPWR.n1286 9.3005
R11204 VPWR.n1285 VPWR.n1279 9.3005
R11205 VPWR.n1290 VPWR.n1289 9.3005
R11206 VPWR.n1293 VPWR.n1292 9.3005
R11207 VPWR.n1295 VPWR.n1275 9.3005
R11208 VPWR.n1320 VPWR.n1319 9.3005
R11209 VPWR.n1315 VPWR.n1302 9.3005
R11210 VPWR.n1312 VPWR.n1310 9.3005
R11211 VPWR.n1309 VPWR.n1303 9.3005
R11212 VPWR.n1314 VPWR.n1313 9.3005
R11213 VPWR.n1317 VPWR.n1316 9.3005
R11214 VPWR.n1318 VPWR.n1299 9.3005
R11215 VPWR.n1351 VPWR.n1322 9.3005
R11216 VPWR.n1350 VPWR.n1349 9.3005
R11217 VPWR.n1330 VPWR.n1329 9.3005
R11218 VPWR.n1332 VPWR.n1331 9.3005
R11219 VPWR.n1334 VPWR.n1328 9.3005
R11220 VPWR.n1336 VPWR.n1335 9.3005
R11221 VPWR.n1337 VPWR.n1327 9.3005
R11222 VPWR.n1339 VPWR.n1338 9.3005
R11223 VPWR.n1343 VPWR.n1324 9.3005
R11224 VPWR.n1345 VPWR.n1344 9.3005
R11225 VPWR.n1347 VPWR.n1346 9.3005
R11226 VPWR.n1353 VPWR.n1352 9.3005
R11227 VPWR.n1355 VPWR.n1354 9.3005
R11228 VPWR.n1394 VPWR.n1393 9.3005
R11229 VPWR.n1389 VPWR.n1357 9.3005
R11230 VPWR.n1388 VPWR.n1387 9.3005
R11231 VPWR.n1366 VPWR.n1365 9.3005
R11232 VPWR.n1368 VPWR.n1367 9.3005
R11233 VPWR.n1371 VPWR.n1361 9.3005
R11234 VPWR.n1373 VPWR.n1372 9.3005
R11235 VPWR.n1374 VPWR.n1360 9.3005
R11236 VPWR.n1376 VPWR.n1375 9.3005
R11237 VPWR.n1380 VPWR.n1359 9.3005
R11238 VPWR.n1382 VPWR.n1381 9.3005
R11239 VPWR.n1384 VPWR.n1383 9.3005
R11240 VPWR.n1391 VPWR.n1390 9.3005
R11241 VPWR.n1427 VPWR.n1426 9.3005
R11242 VPWR.n1405 VPWR.n1404 9.3005
R11243 VPWR.n1407 VPWR.n1406 9.3005
R11244 VPWR.n1410 VPWR.n1400 9.3005
R11245 VPWR.n1412 VPWR.n1411 9.3005
R11246 VPWR.n1413 VPWR.n1399 9.3005
R11247 VPWR.n1415 VPWR.n1414 9.3005
R11248 VPWR.n1419 VPWR.n1398 9.3005
R11249 VPWR.n1421 VPWR.n1420 9.3005
R11250 VPWR.n1423 VPWR.n1422 9.3005
R11251 VPWR.n1428 VPWR.n1396 9.3005
R11252 VPWR.n1430 VPWR.n1429 9.3005
R11253 VPWR.n1464 VPWR.n1463 9.3005
R11254 VPWR.n1442 VPWR.n1441 9.3005
R11255 VPWR.n1444 VPWR.n1443 9.3005
R11256 VPWR.n1447 VPWR.n1437 9.3005
R11257 VPWR.n1449 VPWR.n1448 9.3005
R11258 VPWR.n1450 VPWR.n1436 9.3005
R11259 VPWR.n1452 VPWR.n1451 9.3005
R11260 VPWR.n1456 VPWR.n1435 9.3005
R11261 VPWR.n1458 VPWR.n1457 9.3005
R11262 VPWR.n1460 VPWR.n1459 9.3005
R11263 VPWR.n2826 VPWR.n2825 9.3005
R11264 VPWR.n2827 VPWR.n2819 9.3005
R11265 VPWR.n2828 VPWR.n2818 9.3005
R11266 VPWR.n2829 VPWR.n2817 9.3005
R11267 VPWR.n2831 VPWR.n2830 9.3005
R11268 VPWR.n2815 VPWR.n2814 9.3005
R11269 VPWR.n2809 VPWR.n2808 9.3005
R11270 VPWR.n2810 VPWR.n2800 9.3005
R11271 VPWR.n2812 VPWR.n2811 9.3005
R11272 VPWR.n2813 VPWR.n2798 9.3005
R11273 VPWR.n2796 VPWR.n2795 9.3005
R11274 VPWR.n2794 VPWR.n2778 9.3005
R11275 VPWR.n2789 VPWR.n2788 9.3005
R11276 VPWR.n2790 VPWR.n2780 9.3005
R11277 VPWR.n2792 VPWR.n2791 9.3005
R11278 VPWR.n2776 VPWR.n2775 9.3005
R11279 VPWR.n2770 VPWR.n2769 9.3005
R11280 VPWR.n2771 VPWR.n2761 9.3005
R11281 VPWR.n2773 VPWR.n2772 9.3005
R11282 VPWR.n2774 VPWR.n2759 9.3005
R11283 VPWR.n2757 VPWR.n2756 9.3005
R11284 VPWR.n2737 VPWR.n2736 9.3005
R11285 VPWR.n2738 VPWR.n2732 9.3005
R11286 VPWR.n2740 VPWR.n2739 9.3005
R11287 VPWR.n2742 VPWR.n2730 9.3005
R11288 VPWR.n2744 VPWR.n2743 9.3005
R11289 VPWR.n2746 VPWR.n2745 9.3005
R11290 VPWR.n2747 VPWR.n2726 9.3005
R11291 VPWR.n2751 VPWR.n2750 9.3005
R11292 VPWR.n2752 VPWR.n2725 9.3005
R11293 VPWR.n2754 VPWR.n2753 9.3005
R11294 VPWR.n2755 VPWR.n2723 9.3005
R11295 VPWR.n2721 VPWR.n2720 9.3005
R11296 VPWR.n2701 VPWR.n2700 9.3005
R11297 VPWR.n2702 VPWR.n2695 9.3005
R11298 VPWR.n2704 VPWR.n2703 9.3005
R11299 VPWR.n2706 VPWR.n2692 9.3005
R11300 VPWR.n2708 VPWR.n2707 9.3005
R11301 VPWR.n2710 VPWR.n2709 9.3005
R11302 VPWR.n2711 VPWR.n2688 9.3005
R11303 VPWR.n2714 VPWR.n2713 9.3005
R11304 VPWR.n2715 VPWR.n2687 9.3005
R11305 VPWR.n2717 VPWR.n2716 9.3005
R11306 VPWR.n2718 VPWR.n2685 9.3005
R11307 VPWR.n2664 VPWR.n2663 9.3005
R11308 VPWR.n2665 VPWR.n2658 9.3005
R11309 VPWR.n2667 VPWR.n2666 9.3005
R11310 VPWR.n2669 VPWR.n2655 9.3005
R11311 VPWR.n2671 VPWR.n2670 9.3005
R11312 VPWR.n2673 VPWR.n2672 9.3005
R11313 VPWR.n2674 VPWR.n2651 9.3005
R11314 VPWR.n2677 VPWR.n2676 9.3005
R11315 VPWR.n2678 VPWR.n2650 9.3005
R11316 VPWR.n2680 VPWR.n2679 9.3005
R11317 VPWR.n2681 VPWR.n2648 9.3005
R11318 VPWR.n2646 VPWR.n2645 9.3005
R11319 VPWR.n2628 VPWR.n2627 9.3005
R11320 VPWR.n2630 VPWR.n2623 9.3005
R11321 VPWR.n2635 VPWR.n2634 9.3005
R11322 VPWR.n2636 VPWR.n2622 9.3005
R11323 VPWR.n2638 VPWR.n2637 9.3005
R11324 VPWR.n2640 VPWR.n2619 9.3005
R11325 VPWR.n2642 VPWR.n2641 9.3005
R11326 VPWR.n2644 VPWR.n2643 9.3005
R11327 VPWR.n2524 VPWR.n2523 9.3005
R11328 VPWR.n2588 VPWR.n2587 9.3005
R11329 VPWR.n2528 VPWR.n2527 9.3005
R11330 VPWR.n2572 VPWR.n2571 9.3005
R11331 VPWR.n2564 VPWR.n2563 9.3005
R11332 VPWR.n2552 VPWR.n2551 9.3005
R11333 VPWR.n2548 VPWR.n2547 9.3005
R11334 VPWR.n1241 VPWR.n1240 9.3005
R11335 VPWR.n2540 VPWR.n2539 9.3005
R11336 VPWR.n1203 VPWR.n1121 9.3005
R11337 VPWR.n1237 VPWR.n1113 9.3005
R11338 VPWR.n2560 VPWR.n2559 9.3005
R11339 VPWR.n1234 VPWR.n1111 9.3005
R11340 VPWR.n1231 VPWR.n1230 9.3005
R11341 VPWR.n2536 VPWR.n2535 9.3005
R11342 VPWR.n1200 VPWR.n1123 9.3005
R11343 VPWR.n1223 VPWR.n1103 9.3005
R11344 VPWR.n2576 VPWR.n2575 9.3005
R11345 VPWR.n1220 VPWR.n1101 9.3005
R11346 VPWR.n1611 VPWR.n1610 9.3005
R11347 VPWR.n2584 VPWR.n2583 9.3005
R11348 VPWR.n1217 VPWR.n1216 9.3005
R11349 VPWR.n1209 VPWR.n1093 9.3005
R11350 VPWR.n1761 VPWR.n1760 9.3005
R11351 VPWR.n1206 VPWR.n1090 9.3005
R11352 VPWR.n2596 VPWR.n2595 9.3005
R11353 VPWR.n2600 VPWR.n2599 9.3005
R11354 VPWR.n2611 VPWR.n2610 9.3005
R11355 VPWR.n2608 VPWR.n2607 9.3005
R11356 VPWR.n1757 VPWR.n1756 9.3005
R11357 VPWR.n1082 VPWR.n1081 9.3005
R11358 VPWR.n1615 VPWR.n1614 9.3005
R11359 VPWR.n2841 VPWR.n30 8.40959
R11360 VPWR.n2835 VPWR.n30 8.40959
R11361 VPWR.n28 VPWR.n25 8.40959
R11362 VPWR.n2835 VPWR.n28 8.40959
R11363 VPWR.n2836 VPWR.n27 8.40959
R11364 VPWR.n2835 VPWR.n27 8.40959
R11365 VPWR.n2834 VPWR.n29 8.40959
R11366 VPWR.n2835 VPWR.n29 8.40959
R11367 VPWR.n1294 VPWR.n1293 8.28285
R11368 VPWR.n2793 VPWR.n2792 8.28285
R11369 VPWR.n1626 VPWR.n1128 8.25914
R11370 VPWR.n1747 VPWR.n1746 8.25914
R11371 VPWR.n300 VPWR.n132 8.25914
R11372 VPWR.n155 VPWR.n143 8.25914
R11373 VPWR.n1799 VPWR.n1798 7.91351
R11374 VPWR.n1790 VPWR.n1789 7.9105
R11375 VPWR.n1061 VPWR.n1060 7.9105
R11376 VPWR.n1565 VPWR.n1564 7.9105
R11377 VPWR.n1570 VPWR.n1569 7.9105
R11378 VPWR.n1575 VPWR.n1574 7.9105
R11379 VPWR.n1580 VPWR.n1579 7.9105
R11380 VPWR.n1585 VPWR.n1584 7.9105
R11381 VPWR.n1590 VPWR.n1589 7.9105
R11382 VPWR.n1595 VPWR.n1594 7.9105
R11383 VPWR.n1600 VPWR.n1599 7.9105
R11384 VPWR.n1155 VPWR.n1154 7.9105
R11385 VPWR.n1480 VPWR.n1479 7.9105
R11386 VPWR.n1475 VPWR.n1474 7.9105
R11387 VPWR.n1795 VPWR.n1794 7.9105
R11388 VPWR.n1803 VPWR.n1802 7.9105
R11389 VPWR.n301 VPWR.n300 7.9105
R11390 VPWR.n299 VPWR.n298 7.9105
R11391 VPWR.n287 VPWR.n286 7.9105
R11392 VPWR.n275 VPWR.n274 7.9105
R11393 VPWR.n263 VPWR.n262 7.9105
R11394 VPWR.n251 VPWR.n250 7.9105
R11395 VPWR.n239 VPWR.n238 7.9105
R11396 VPWR.n227 VPWR.n226 7.9105
R11397 VPWR.n215 VPWR.n214 7.9105
R11398 VPWR.n203 VPWR.n202 7.9105
R11399 VPWR.n191 VPWR.n190 7.9105
R11400 VPWR.n179 VPWR.n178 7.9105
R11401 VPWR.n167 VPWR.n166 7.9105
R11402 VPWR.n155 VPWR.n154 7.9105
R11403 VPWR.n1746 VPWR.n1745 7.9105
R11404 VPWR.n1734 VPWR.n1733 7.9105
R11405 VPWR.n1720 VPWR.n1087 7.9105
R11406 VPWR.n1709 VPWR.n1708 7.9105
R11407 VPWR.n1707 VPWR.n1706 7.9105
R11408 VPWR.n1693 VPWR.n1098 7.9105
R11409 VPWR.n1682 VPWR.n1681 7.9105
R11410 VPWR.n1680 VPWR.n1679 7.9105
R11411 VPWR.n1666 VPWR.n1108 7.9105
R11412 VPWR.n1655 VPWR.n1654 7.9105
R11413 VPWR.n1653 VPWR.n1652 7.9105
R11414 VPWR.n1639 VPWR.n1118 7.9105
R11415 VPWR.n1628 VPWR.n1627 7.9105
R11416 VPWR.n1626 VPWR.n1625 7.9105
R11417 VPWR.n45 VPWR.n43 7.8627
R11418 VPWR.n7 VPWR.n6 7.56315
R11419 VPWR.n1261 VPWR.n1260 7.56315
R11420 VPWR.n1284 VPWR.n1283 7.56315
R11421 VPWR.n1308 VPWR.n1307 7.56315
R11422 VPWR.n2844 VPWR.n2843 7.0697
R11423 VPWR.n2860 VPWR.n2859 6.57193
R11424 VPWR.n2824 VPWR.n2822 6.4511
R11425 VPWR.n2807 VPWR.n2804 6.4511
R11426 VPWR.n2787 VPWR.n2784 6.4511
R11427 VPWR.n2768 VPWR.n2765 6.4511
R11428 VPWR.n1381 VPWR.n1358 6.4005
R11429 VPWR.n1420 VPWR.n1397 6.4005
R11430 VPWR.n1457 VPWR.n1434 6.4005
R11431 VPWR.n2742 VPWR.n2741 6.4005
R11432 VPWR.n2712 VPWR.n2711 6.4005
R11433 VPWR.n2675 VPWR.n2674 6.4005
R11434 VPWR.n2641 VPWR.n2618 6.4005
R11435 VPWR.n1614 VPWR.n1141 6.04494
R11436 VPWR.n2524 VPWR.n118 6.04494
R11437 VPWR.n1486 VPWR.n1250 6.04494
R11438 VPWR.n370 VPWR.n309 6.04494
R11439 VPWR.n2587 VPWR.n87 6.04494
R11440 VPWR.n1553 VPWR.n1172 6.04494
R11441 VPWR.n367 VPWR.n365 6.04494
R11442 VPWR.n2527 VPWR.n117 6.04494
R11443 VPWR.n984 VPWR.n982 6.04494
R11444 VPWR.n2497 VPWR.n375 6.04494
R11445 VPWR.n2494 VPWR.n376 6.04494
R11446 VPWR.n339 VPWR.n337 6.04494
R11447 VPWR.n2572 VPWR.n94 6.04494
R11448 VPWR.n992 VPWR.n990 6.04494
R11449 VPWR.n2464 VPWR.n388 6.04494
R11450 VPWR.n343 VPWR.n341 6.04494
R11451 VPWR.n2563 VPWR.n99 6.04494
R11452 VPWR.n1909 VPWR.n951 6.04494
R11453 VPWR.n1906 VPWR.n952 6.04494
R11454 VPWR.n1899 VPWR.n955 6.04494
R11455 VPWR.n408 VPWR.n406 6.04494
R11456 VPWR.n412 VPWR.n410 6.04494
R11457 VPWR.n416 VPWR.n414 6.04494
R11458 VPWR.n2474 VPWR.n384 6.04494
R11459 VPWR.n351 VPWR.n349 6.04494
R11460 VPWR.n2551 VPWR.n105 6.04494
R11461 VPWR.n1896 VPWR.n956 6.04494
R11462 VPWR.n424 VPWR.n422 6.04494
R11463 VPWR.n2477 VPWR.n383 6.04494
R11464 VPWR.n355 VPWR.n353 6.04494
R11465 VPWR.n2548 VPWR.n106 6.04494
R11466 VPWR.n2327 VPWR.n500 6.04494
R11467 VPWR.n2330 VPWR.n499 6.04494
R11468 VPWR.n2337 VPWR.n496 6.04494
R11469 VPWR.n2340 VPWR.n495 6.04494
R11470 VPWR.n2350 VPWR.n491 6.04494
R11471 VPWR.n2357 VPWR.n488 6.04494
R11472 VPWR.n2360 VPWR.n487 6.04494
R11473 VPWR.n2367 VPWR.n484 6.04494
R11474 VPWR.n2370 VPWR.n483 6.04494
R11475 VPWR.n2377 VPWR.n480 6.04494
R11476 VPWR.n2380 VPWR.n479 6.04494
R11477 VPWR.n2387 VPWR.n476 6.04494
R11478 VPWR.n2390 VPWR.n475 6.04494
R11479 VPWR.n2397 VPWR.n472 6.04494
R11480 VPWR.n2399 VPWR.n471 6.04494
R11481 VPWR.n2347 VPWR.n492 6.04494
R11482 VPWR.n562 VPWR.n501 6.04494
R11483 VPWR.n559 VPWR.n557 6.04494
R11484 VPWR.n555 VPWR.n553 6.04494
R11485 VPWR.n551 VPWR.n549 6.04494
R11486 VPWR.n543 VPWR.n541 6.04494
R11487 VPWR.n539 VPWR.n537 6.04494
R11488 VPWR.n535 VPWR.n533 6.04494
R11489 VPWR.n531 VPWR.n529 6.04494
R11490 VPWR.n527 VPWR.n525 6.04494
R11491 VPWR.n523 VPWR.n521 6.04494
R11492 VPWR.n519 VPWR.n517 6.04494
R11493 VPWR.n515 VPWR.n513 6.04494
R11494 VPWR.n511 VPWR.n509 6.04494
R11495 VPWR.n507 VPWR.n505 6.04494
R11496 VPWR.n504 VPWR.n502 6.04494
R11497 VPWR.n547 VPWR.n545 6.04494
R11498 VPWR.n2301 VPWR.n567 6.04494
R11499 VPWR.n2298 VPWR.n568 6.04494
R11500 VPWR.n2291 VPWR.n571 6.04494
R11501 VPWR.n2288 VPWR.n572 6.04494
R11502 VPWR.n2278 VPWR.n576 6.04494
R11503 VPWR.n2271 VPWR.n579 6.04494
R11504 VPWR.n2268 VPWR.n580 6.04494
R11505 VPWR.n2261 VPWR.n583 6.04494
R11506 VPWR.n2258 VPWR.n584 6.04494
R11507 VPWR.n2251 VPWR.n587 6.04494
R11508 VPWR.n2248 VPWR.n588 6.04494
R11509 VPWR.n2241 VPWR.n591 6.04494
R11510 VPWR.n2238 VPWR.n592 6.04494
R11511 VPWR.n2231 VPWR.n595 6.04494
R11512 VPWR.n2229 VPWR.n596 6.04494
R11513 VPWR.n2281 VPWR.n575 6.04494
R11514 VPWR.n600 VPWR.n598 6.04494
R11515 VPWR.n604 VPWR.n602 6.04494
R11516 VPWR.n608 VPWR.n606 6.04494
R11517 VPWR.n612 VPWR.n610 6.04494
R11518 VPWR.n620 VPWR.n618 6.04494
R11519 VPWR.n624 VPWR.n622 6.04494
R11520 VPWR.n628 VPWR.n626 6.04494
R11521 VPWR.n632 VPWR.n630 6.04494
R11522 VPWR.n636 VPWR.n634 6.04494
R11523 VPWR.n640 VPWR.n638 6.04494
R11524 VPWR.n644 VPWR.n642 6.04494
R11525 VPWR.n648 VPWR.n646 6.04494
R11526 VPWR.n652 VPWR.n650 6.04494
R11527 VPWR.n656 VPWR.n654 6.04494
R11528 VPWR.n658 VPWR.n597 6.04494
R11529 VPWR.n616 VPWR.n614 6.04494
R11530 VPWR.n2131 VPWR.n692 6.04494
R11531 VPWR.n2134 VPWR.n691 6.04494
R11532 VPWR.n2141 VPWR.n688 6.04494
R11533 VPWR.n2144 VPWR.n687 6.04494
R11534 VPWR.n2154 VPWR.n683 6.04494
R11535 VPWR.n2161 VPWR.n680 6.04494
R11536 VPWR.n2164 VPWR.n679 6.04494
R11537 VPWR.n2171 VPWR.n676 6.04494
R11538 VPWR.n2174 VPWR.n675 6.04494
R11539 VPWR.n2181 VPWR.n672 6.04494
R11540 VPWR.n2184 VPWR.n671 6.04494
R11541 VPWR.n2191 VPWR.n668 6.04494
R11542 VPWR.n2194 VPWR.n667 6.04494
R11543 VPWR.n2201 VPWR.n664 6.04494
R11544 VPWR.n2203 VPWR.n663 6.04494
R11545 VPWR.n2151 VPWR.n684 6.04494
R11546 VPWR.n754 VPWR.n693 6.04494
R11547 VPWR.n751 VPWR.n749 6.04494
R11548 VPWR.n747 VPWR.n745 6.04494
R11549 VPWR.n743 VPWR.n741 6.04494
R11550 VPWR.n735 VPWR.n733 6.04494
R11551 VPWR.n731 VPWR.n729 6.04494
R11552 VPWR.n727 VPWR.n725 6.04494
R11553 VPWR.n723 VPWR.n721 6.04494
R11554 VPWR.n719 VPWR.n717 6.04494
R11555 VPWR.n715 VPWR.n713 6.04494
R11556 VPWR.n711 VPWR.n709 6.04494
R11557 VPWR.n707 VPWR.n705 6.04494
R11558 VPWR.n703 VPWR.n701 6.04494
R11559 VPWR.n699 VPWR.n697 6.04494
R11560 VPWR.n696 VPWR.n694 6.04494
R11561 VPWR.n739 VPWR.n737 6.04494
R11562 VPWR.n2105 VPWR.n759 6.04494
R11563 VPWR.n2102 VPWR.n760 6.04494
R11564 VPWR.n2095 VPWR.n763 6.04494
R11565 VPWR.n2092 VPWR.n764 6.04494
R11566 VPWR.n2082 VPWR.n768 6.04494
R11567 VPWR.n2075 VPWR.n771 6.04494
R11568 VPWR.n2072 VPWR.n772 6.04494
R11569 VPWR.n2065 VPWR.n775 6.04494
R11570 VPWR.n2062 VPWR.n776 6.04494
R11571 VPWR.n2055 VPWR.n779 6.04494
R11572 VPWR.n2052 VPWR.n780 6.04494
R11573 VPWR.n2045 VPWR.n783 6.04494
R11574 VPWR.n2042 VPWR.n784 6.04494
R11575 VPWR.n2035 VPWR.n787 6.04494
R11576 VPWR.n2033 VPWR.n788 6.04494
R11577 VPWR.n2085 VPWR.n767 6.04494
R11578 VPWR.n792 VPWR.n790 6.04494
R11579 VPWR.n796 VPWR.n794 6.04494
R11580 VPWR.n800 VPWR.n798 6.04494
R11581 VPWR.n804 VPWR.n802 6.04494
R11582 VPWR.n812 VPWR.n810 6.04494
R11583 VPWR.n816 VPWR.n814 6.04494
R11584 VPWR.n820 VPWR.n818 6.04494
R11585 VPWR.n824 VPWR.n822 6.04494
R11586 VPWR.n828 VPWR.n826 6.04494
R11587 VPWR.n832 VPWR.n830 6.04494
R11588 VPWR.n836 VPWR.n834 6.04494
R11589 VPWR.n840 VPWR.n838 6.04494
R11590 VPWR.n844 VPWR.n842 6.04494
R11591 VPWR.n848 VPWR.n846 6.04494
R11592 VPWR.n850 VPWR.n789 6.04494
R11593 VPWR.n808 VPWR.n806 6.04494
R11594 VPWR.n1935 VPWR.n884 6.04494
R11595 VPWR.n1938 VPWR.n883 6.04494
R11596 VPWR.n1945 VPWR.n880 6.04494
R11597 VPWR.n1948 VPWR.n879 6.04494
R11598 VPWR.n1958 VPWR.n875 6.04494
R11599 VPWR.n1965 VPWR.n872 6.04494
R11600 VPWR.n1968 VPWR.n871 6.04494
R11601 VPWR.n1975 VPWR.n868 6.04494
R11602 VPWR.n1978 VPWR.n867 6.04494
R11603 VPWR.n1985 VPWR.n864 6.04494
R11604 VPWR.n1988 VPWR.n863 6.04494
R11605 VPWR.n1995 VPWR.n860 6.04494
R11606 VPWR.n1998 VPWR.n859 6.04494
R11607 VPWR.n2005 VPWR.n856 6.04494
R11608 VPWR.n2007 VPWR.n855 6.04494
R11609 VPWR.n1955 VPWR.n876 6.04494
R11610 VPWR.n946 VPWR.n885 6.04494
R11611 VPWR.n943 VPWR.n941 6.04494
R11612 VPWR.n939 VPWR.n937 6.04494
R11613 VPWR.n935 VPWR.n933 6.04494
R11614 VPWR.n927 VPWR.n925 6.04494
R11615 VPWR.n923 VPWR.n921 6.04494
R11616 VPWR.n919 VPWR.n917 6.04494
R11617 VPWR.n915 VPWR.n913 6.04494
R11618 VPWR.n911 VPWR.n909 6.04494
R11619 VPWR.n907 VPWR.n905 6.04494
R11620 VPWR.n903 VPWR.n901 6.04494
R11621 VPWR.n899 VPWR.n897 6.04494
R11622 VPWR.n895 VPWR.n893 6.04494
R11623 VPWR.n891 VPWR.n889 6.04494
R11624 VPWR.n888 VPWR.n886 6.04494
R11625 VPWR.n931 VPWR.n929 6.04494
R11626 VPWR.n1889 VPWR.n959 6.04494
R11627 VPWR.n1000 VPWR.n998 6.04494
R11628 VPWR.n1513 VPWR.n1246 6.04494
R11629 VPWR.n1240 VPWR.n1198 6.04494
R11630 VPWR.n420 VPWR.n418 6.04494
R11631 VPWR.n2484 VPWR.n380 6.04494
R11632 VPWR.n359 VPWR.n357 6.04494
R11633 VPWR.n2539 VPWR.n111 6.04494
R11634 VPWR.n996 VPWR.n994 6.04494
R11635 VPWR.n1510 VPWR.n1504 6.04494
R11636 VPWR.n1203 VPWR.n1202 6.04494
R11637 VPWR.n1886 VPWR.n960 6.04494
R11638 VPWR.n1004 VPWR.n1002 6.04494
R11639 VPWR.n1524 VPWR.n1192 6.04494
R11640 VPWR.n1237 VPWR.n1236 6.04494
R11641 VPWR.n428 VPWR.n426 6.04494
R11642 VPWR.n436 VPWR.n434 6.04494
R11643 VPWR.n440 VPWR.n438 6.04494
R11644 VPWR.n444 VPWR.n442 6.04494
R11645 VPWR.n448 VPWR.n446 6.04494
R11646 VPWR.n452 VPWR.n450 6.04494
R11647 VPWR.n456 VPWR.n454 6.04494
R11648 VPWR.n460 VPWR.n458 6.04494
R11649 VPWR.n464 VPWR.n462 6.04494
R11650 VPWR.n466 VPWR.n405 6.04494
R11651 VPWR.n432 VPWR.n430 6.04494
R11652 VPWR.n2467 VPWR.n387 6.04494
R11653 VPWR.n347 VPWR.n345 6.04494
R11654 VPWR.n2560 VPWR.n100 6.04494
R11655 VPWR.n1008 VPWR.n1006 6.04494
R11656 VPWR.n1527 VPWR.n1188 6.04494
R11657 VPWR.n1234 VPWR.n1233 6.04494
R11658 VPWR.n1879 VPWR.n963 6.04494
R11659 VPWR.n1869 VPWR.n967 6.04494
R11660 VPWR.n1866 VPWR.n968 6.04494
R11661 VPWR.n1859 VPWR.n971 6.04494
R11662 VPWR.n1856 VPWR.n972 6.04494
R11663 VPWR.n1849 VPWR.n975 6.04494
R11664 VPWR.n1846 VPWR.n976 6.04494
R11665 VPWR.n1839 VPWR.n979 6.04494
R11666 VPWR.n1837 VPWR.n980 6.04494
R11667 VPWR.n1876 VPWR.n964 6.04494
R11668 VPWR.n1012 VPWR.n1010 6.04494
R11669 VPWR.n1538 VPWR.n1182 6.04494
R11670 VPWR.n1231 VPWR.n1225 6.04494
R11671 VPWR.n2487 VPWR.n379 6.04494
R11672 VPWR.n363 VPWR.n361 6.04494
R11673 VPWR.n2536 VPWR.n112 6.04494
R11674 VPWR.n1499 VPWR.n1498 6.04494
R11675 VPWR.n1200 VPWR.n1199 6.04494
R11676 VPWR.n1016 VPWR.n1014 6.04494
R11677 VPWR.n1541 VPWR.n1178 6.04494
R11678 VPWR.n1223 VPWR.n1222 6.04494
R11679 VPWR.n2457 VPWR.n391 6.04494
R11680 VPWR.n2447 VPWR.n395 6.04494
R11681 VPWR.n2444 VPWR.n396 6.04494
R11682 VPWR.n2437 VPWR.n399 6.04494
R11683 VPWR.n2434 VPWR.n400 6.04494
R11684 VPWR.n2427 VPWR.n403 6.04494
R11685 VPWR.n2425 VPWR.n404 6.04494
R11686 VPWR.n2454 VPWR.n392 6.04494
R11687 VPWR.n335 VPWR.n333 6.04494
R11688 VPWR.n2575 VPWR.n93 6.04494
R11689 VPWR.n1556 VPWR.n1168 6.04494
R11690 VPWR.n1220 VPWR.n1219 6.04494
R11691 VPWR.n1020 VPWR.n1018 6.04494
R11692 VPWR.n1024 VPWR.n1022 6.04494
R11693 VPWR.n1028 VPWR.n1026 6.04494
R11694 VPWR.n1032 VPWR.n1030 6.04494
R11695 VPWR.n1036 VPWR.n1034 6.04494
R11696 VPWR.n1040 VPWR.n1038 6.04494
R11697 VPWR.n1042 VPWR.n981 6.04494
R11698 VPWR.n988 VPWR.n986 6.04494
R11699 VPWR.n1493 VPWR.n1491 6.04494
R11700 VPWR.n1611 VPWR.n1142 6.04494
R11701 VPWR.n331 VPWR.n329 6.04494
R11702 VPWR.n2584 VPWR.n88 6.04494
R11703 VPWR.n1217 VPWR.n1211 6.04494
R11704 VPWR.n1781 VPWR.n1068 6.04494
R11705 VPWR.n1209 VPWR.n1208 6.04494
R11706 VPWR.n327 VPWR.n325 6.04494
R11707 VPWR.n323 VPWR.n321 6.04494
R11708 VPWR.n315 VPWR.n313 6.04494
R11709 VPWR.n312 VPWR.n310 6.04494
R11710 VPWR.n319 VPWR.n317 6.04494
R11711 VPWR.n1760 VPWR.n1077 6.04494
R11712 VPWR.n1769 VPWR.n1767 6.04494
R11713 VPWR.n1809 VPWR.n1055 6.04494
R11714 VPWR.n1811 VPWR.n1051 6.04494
R11715 VPWR.n1778 VPWR.n1072 6.04494
R11716 VPWR.n1206 VPWR.n1205 6.04494
R11717 VPWR.n2596 VPWR.n82 6.04494
R11718 VPWR.n2599 VPWR.n81 6.04494
R11719 VPWR.n2608 VPWR.n76 6.04494
R11720 VPWR.n2610 VPWR.n75 6.04494
R11721 VPWR.n1757 VPWR.n1078 6.04494
R11722 VPWR.n1081 VPWR.n1080 6.04494
R11723 VPWR.n2858 VPWR.n20 5.59663
R11724 VPWR.n2861 VPWR.n2860 5.59663
R11725 VPWR.n2859 VPWR.n22 5.59425
R11726 VPWR.n2845 VPWR.n2844 5.59425
R11727 VPWR.n2804 VPWR.n2803 5.39628
R11728 VPWR.n2784 VPWR.n2783 5.39628
R11729 VPWR.n2765 VPWR.n2764 5.39628
R11730 VPWR.n2844 VPWR.n23 4.9938
R11731 VPWR VPWR.n2833 4.94464
R11732 VPWR.n73 VPWR 4.72593
R11733 VPWR.n71 VPWR 4.72593
R11734 VPWR.n69 VPWR 4.72593
R11735 VPWR.n67 VPWR 4.72593
R11736 VPWR.n65 VPWR 4.72593
R11737 VPWR.n63 VPWR 4.72593
R11738 VPWR.n61 VPWR 4.72593
R11739 VPWR.n59 VPWR 4.72593
R11740 VPWR.n57 VPWR 4.72593
R11741 VPWR.n55 VPWR 4.72593
R11742 VPWR.n53 VPWR 4.72593
R11743 VPWR.n51 VPWR 4.72593
R11744 VPWR.n49 VPWR 4.72593
R11745 VPWR.n47 VPWR 4.72593
R11746 VPWR.n45 VPWR 4.72593
R11747 VPWR.n36 VPWR.n26 4.6505
R11748 VPWR.n2847 VPWR.n2846 4.6505
R11749 VPWR.n34 VPWR.n23 4.6505
R11750 VPWR.n2857 VPWR.n2856 4.6505
R11751 VPWR.n2843 VPWR.n2842 4.6505
R11752 VPWR.n2837 VPWR.n21 4.6505
R11753 VPWR.n1465 VPWR.n1464 4.55954
R11754 VPWR.n2859 VPWR.n2858 4.5005
R11755 VPWR.n2590 VPWR.n2589 4.5005
R11756 VPWR.n2530 VPWR.n2529 4.5005
R11757 VPWR.n2570 VPWR.n2569 4.5005
R11758 VPWR.n338 VPWR.n96 4.5005
R11759 VPWR.n2566 VPWR.n2565 4.5005
R11760 VPWR.n342 VPWR.n97 4.5005
R11761 VPWR.n2554 VPWR.n2553 4.5005
R11762 VPWR.n350 VPWR.n103 4.5005
R11763 VPWR.n2473 VPWR.n2472 4.5005
R11764 VPWR.n2546 VPWR.n2545 4.5005
R11765 VPWR.n354 VPWR.n108 4.5005
R11766 VPWR.n2479 VPWR.n2478 4.5005
R11767 VPWR.n1517 VPWR.n1242 4.5005
R11768 VPWR.n1516 VPWR.n1514 4.5005
R11769 VPWR.n999 VPWR.n958 4.5005
R11770 VPWR.n1891 VPWR.n1890 4.5005
R11771 VPWR.n930 VPWR.n877 4.5005
R11772 VPWR.n1954 VPWR.n1953 4.5005
R11773 VPWR.n807 VPWR.n766 4.5005
R11774 VPWR.n2087 VPWR.n2086 4.5005
R11775 VPWR.n738 VPWR.n685 4.5005
R11776 VPWR.n2150 VPWR.n2149 4.5005
R11777 VPWR.n615 VPWR.n574 4.5005
R11778 VPWR.n2283 VPWR.n2282 4.5005
R11779 VPWR.n546 VPWR.n493 4.5005
R11780 VPWR.n2346 VPWR.n2345 4.5005
R11781 VPWR.n423 VPWR.n382 4.5005
R11782 VPWR.n2542 VPWR.n2541 4.5005
R11783 VPWR.n358 VPWR.n109 4.5005
R11784 VPWR.n2483 VPWR.n2482 4.5005
R11785 VPWR.n419 VPWR.n381 4.5005
R11786 VPWR.n2342 VPWR.n2341 4.5005
R11787 VPWR.n550 VPWR.n494 4.5005
R11788 VPWR.n2287 VPWR.n2286 4.5005
R11789 VPWR.n611 VPWR.n573 4.5005
R11790 VPWR.n2146 VPWR.n2145 4.5005
R11791 VPWR.n742 VPWR.n686 4.5005
R11792 VPWR.n2091 VPWR.n2090 4.5005
R11793 VPWR.n803 VPWR.n765 4.5005
R11794 VPWR.n1950 VPWR.n1949 4.5005
R11795 VPWR.n934 VPWR.n878 4.5005
R11796 VPWR.n1507 VPWR.n1505 4.5005
R11797 VPWR.n1509 VPWR.n1508 4.5005
R11798 VPWR.n995 VPWR.n957 4.5005
R11799 VPWR.n1895 VPWR.n1894 4.5005
R11800 VPWR.n1520 VPWR.n1193 4.5005
R11801 VPWR.n1523 VPWR.n1522 4.5005
R11802 VPWR.n1003 VPWR.n961 4.5005
R11803 VPWR.n1885 VPWR.n1884 4.5005
R11804 VPWR.n926 VPWR.n874 4.5005
R11805 VPWR.n1960 VPWR.n1959 4.5005
R11806 VPWR.n811 VPWR.n769 4.5005
R11807 VPWR.n2081 VPWR.n2080 4.5005
R11808 VPWR.n734 VPWR.n682 4.5005
R11809 VPWR.n2156 VPWR.n2155 4.5005
R11810 VPWR.n619 VPWR.n577 4.5005
R11811 VPWR.n2277 VPWR.n2276 4.5005
R11812 VPWR.n542 VPWR.n490 4.5005
R11813 VPWR.n2352 VPWR.n2351 4.5005
R11814 VPWR.n427 VPWR.n385 4.5005
R11815 VPWR.n2558 VPWR.n2557 4.5005
R11816 VPWR.n346 VPWR.n102 4.5005
R11817 VPWR.n2469 VPWR.n2468 4.5005
R11818 VPWR.n431 VPWR.n386 4.5005
R11819 VPWR.n2356 VPWR.n2355 4.5005
R11820 VPWR.n538 VPWR.n489 4.5005
R11821 VPWR.n2273 VPWR.n2272 4.5005
R11822 VPWR.n623 VPWR.n578 4.5005
R11823 VPWR.n2160 VPWR.n2159 4.5005
R11824 VPWR.n730 VPWR.n681 4.5005
R11825 VPWR.n2077 VPWR.n2076 4.5005
R11826 VPWR.n815 VPWR.n770 4.5005
R11827 VPWR.n1964 VPWR.n1963 4.5005
R11828 VPWR.n922 VPWR.n873 4.5005
R11829 VPWR.n1531 VPWR.n1184 4.5005
R11830 VPWR.n1530 VPWR.n1528 4.5005
R11831 VPWR.n1007 VPWR.n962 4.5005
R11832 VPWR.n1881 VPWR.n1880 4.5005
R11833 VPWR.n1534 VPWR.n1183 4.5005
R11834 VPWR.n1537 VPWR.n1536 4.5005
R11835 VPWR.n1011 VPWR.n965 4.5005
R11836 VPWR.n1875 VPWR.n1874 4.5005
R11837 VPWR.n918 VPWR.n870 4.5005
R11838 VPWR.n1970 VPWR.n1969 4.5005
R11839 VPWR.n819 VPWR.n773 4.5005
R11840 VPWR.n2071 VPWR.n2070 4.5005
R11841 VPWR.n726 VPWR.n678 4.5005
R11842 VPWR.n2166 VPWR.n2165 4.5005
R11843 VPWR.n627 VPWR.n581 4.5005
R11844 VPWR.n2267 VPWR.n2266 4.5005
R11845 VPWR.n534 VPWR.n486 4.5005
R11846 VPWR.n2362 VPWR.n2361 4.5005
R11847 VPWR.n435 VPWR.n389 4.5005
R11848 VPWR.n2463 VPWR.n2462 4.5005
R11849 VPWR.n2534 VPWR.n2533 4.5005
R11850 VPWR.n362 VPWR.n114 4.5005
R11851 VPWR.n2489 VPWR.n2488 4.5005
R11852 VPWR.n415 VPWR.n378 4.5005
R11853 VPWR.n2336 VPWR.n2335 4.5005
R11854 VPWR.n554 VPWR.n497 4.5005
R11855 VPWR.n2293 VPWR.n2292 4.5005
R11856 VPWR.n607 VPWR.n570 4.5005
R11857 VPWR.n2140 VPWR.n2139 4.5005
R11858 VPWR.n746 VPWR.n689 4.5005
R11859 VPWR.n2097 VPWR.n2096 4.5005
R11860 VPWR.n799 VPWR.n762 4.5005
R11861 VPWR.n1944 VPWR.n1943 4.5005
R11862 VPWR.n938 VPWR.n881 4.5005
R11863 VPWR.n1901 VPWR.n1900 4.5005
R11864 VPWR.n1605 VPWR.n1148 4.5005
R11865 VPWR.n1604 VPWR.n1149 4.5005
R11866 VPWR.n991 VPWR.n954 4.5005
R11867 VPWR.n1545 VPWR.n1174 4.5005
R11868 VPWR.n1544 VPWR.n1542 4.5005
R11869 VPWR.n1015 VPWR.n966 4.5005
R11870 VPWR.n1871 VPWR.n1870 4.5005
R11871 VPWR.n914 VPWR.n869 4.5005
R11872 VPWR.n1974 VPWR.n1973 4.5005
R11873 VPWR.n823 VPWR.n774 4.5005
R11874 VPWR.n2067 VPWR.n2066 4.5005
R11875 VPWR.n722 VPWR.n677 4.5005
R11876 VPWR.n2170 VPWR.n2169 4.5005
R11877 VPWR.n631 VPWR.n582 4.5005
R11878 VPWR.n2263 VPWR.n2262 4.5005
R11879 VPWR.n530 VPWR.n485 4.5005
R11880 VPWR.n2366 VPWR.n2365 4.5005
R11881 VPWR.n439 VPWR.n390 4.5005
R11882 VPWR.n2459 VPWR.n2458 4.5005
R11883 VPWR.n2578 VPWR.n2577 4.5005
R11884 VPWR.n334 VPWR.n91 4.5005
R11885 VPWR.n2453 VPWR.n2452 4.5005
R11886 VPWR.n443 VPWR.n393 4.5005
R11887 VPWR.n2372 VPWR.n2371 4.5005
R11888 VPWR.n526 VPWR.n482 4.5005
R11889 VPWR.n2257 VPWR.n2256 4.5005
R11890 VPWR.n635 VPWR.n585 4.5005
R11891 VPWR.n2176 VPWR.n2175 4.5005
R11892 VPWR.n718 VPWR.n674 4.5005
R11893 VPWR.n2061 VPWR.n2060 4.5005
R11894 VPWR.n827 VPWR.n777 4.5005
R11895 VPWR.n1980 VPWR.n1979 4.5005
R11896 VPWR.n910 VPWR.n866 4.5005
R11897 VPWR.n1865 VPWR.n1864 4.5005
R11898 VPWR.n1164 VPWR.n1163 4.5005
R11899 VPWR.n1558 VPWR.n1557 4.5005
R11900 VPWR.n1019 VPWR.n969 4.5005
R11901 VPWR.n1609 VPWR.n1608 4.5005
R11902 VPWR.n1492 VPWR.n1147 4.5005
R11903 VPWR.n987 VPWR.n953 4.5005
R11904 VPWR.n1905 VPWR.n1904 4.5005
R11905 VPWR.n942 VPWR.n882 4.5005
R11906 VPWR.n1940 VPWR.n1939 4.5005
R11907 VPWR.n795 VPWR.n761 4.5005
R11908 VPWR.n2101 VPWR.n2100 4.5005
R11909 VPWR.n750 VPWR.n690 4.5005
R11910 VPWR.n2136 VPWR.n2135 4.5005
R11911 VPWR.n603 VPWR.n569 4.5005
R11912 VPWR.n2297 VPWR.n2296 4.5005
R11913 VPWR.n558 VPWR.n498 4.5005
R11914 VPWR.n2332 VPWR.n2331 4.5005
R11915 VPWR.n411 VPWR.n377 4.5005
R11916 VPWR.n2493 VPWR.n2492 4.5005
R11917 VPWR.n366 VPWR.n115 4.5005
R11918 VPWR.n2582 VPWR.n2581 4.5005
R11919 VPWR.n330 VPWR.n90 4.5005
R11920 VPWR.n2449 VPWR.n2448 4.5005
R11921 VPWR.n447 VPWR.n394 4.5005
R11922 VPWR.n2376 VPWR.n2375 4.5005
R11923 VPWR.n522 VPWR.n481 4.5005
R11924 VPWR.n2253 VPWR.n2252 4.5005
R11925 VPWR.n639 VPWR.n586 4.5005
R11926 VPWR.n2180 VPWR.n2179 4.5005
R11927 VPWR.n714 VPWR.n673 4.5005
R11928 VPWR.n2057 VPWR.n2056 4.5005
R11929 VPWR.n831 VPWR.n778 4.5005
R11930 VPWR.n1984 VPWR.n1983 4.5005
R11931 VPWR.n906 VPWR.n865 4.5005
R11932 VPWR.n1861 VPWR.n1860 4.5005
R11933 VPWR.n1023 VPWR.n970 4.5005
R11934 VPWR.n1550 VPWR.n1173 4.5005
R11935 VPWR.n1552 VPWR.n1551 4.5005
R11936 VPWR.n1092 VPWR.n1064 4.5005
R11937 VPWR.n1783 VPWR.n1782 4.5005
R11938 VPWR.n1027 VPWR.n973 4.5005
R11939 VPWR.n1855 VPWR.n1854 4.5005
R11940 VPWR.n902 VPWR.n862 4.5005
R11941 VPWR.n1990 VPWR.n1989 4.5005
R11942 VPWR.n835 VPWR.n781 4.5005
R11943 VPWR.n2051 VPWR.n2050 4.5005
R11944 VPWR.n710 VPWR.n670 4.5005
R11945 VPWR.n2186 VPWR.n2185 4.5005
R11946 VPWR.n643 VPWR.n589 4.5005
R11947 VPWR.n2247 VPWR.n2246 4.5005
R11948 VPWR.n518 VPWR.n478 4.5005
R11949 VPWR.n2382 VPWR.n2381 4.5005
R11950 VPWR.n451 VPWR.n397 4.5005
R11951 VPWR.n2443 VPWR.n2442 4.5005
R11952 VPWR.n326 VPWR.n85 4.5005
R11953 VPWR.n318 VPWR.n79 4.5005
R11954 VPWR.n2433 VPWR.n2432 4.5005
R11955 VPWR.n459 VPWR.n401 4.5005
R11956 VPWR.n2392 VPWR.n2391 4.5005
R11957 VPWR.n510 VPWR.n474 4.5005
R11958 VPWR.n2237 VPWR.n2236 4.5005
R11959 VPWR.n651 VPWR.n593 4.5005
R11960 VPWR.n2196 VPWR.n2195 4.5005
R11961 VPWR.n702 VPWR.n666 4.5005
R11962 VPWR.n2041 VPWR.n2040 4.5005
R11963 VPWR.n843 VPWR.n785 4.5005
R11964 VPWR.n2000 VPWR.n1999 4.5005
R11965 VPWR.n894 VPWR.n858 4.5005
R11966 VPWR.n1845 VPWR.n1844 4.5005
R11967 VPWR.n1035 VPWR.n977 4.5005
R11968 VPWR.n1772 VPWR.n1762 4.5005
R11969 VPWR.n1771 VPWR.n1770 4.5005
R11970 VPWR.n1775 VPWR.n1073 4.5005
R11971 VPWR.n1777 VPWR.n1776 4.5005
R11972 VPWR.n1031 VPWR.n974 4.5005
R11973 VPWR.n1851 VPWR.n1850 4.5005
R11974 VPWR.n898 VPWR.n861 4.5005
R11975 VPWR.n1994 VPWR.n1993 4.5005
R11976 VPWR.n839 VPWR.n782 4.5005
R11977 VPWR.n2047 VPWR.n2046 4.5005
R11978 VPWR.n706 VPWR.n669 4.5005
R11979 VPWR.n2190 VPWR.n2189 4.5005
R11980 VPWR.n647 VPWR.n590 4.5005
R11981 VPWR.n2243 VPWR.n2242 4.5005
R11982 VPWR.n514 VPWR.n477 4.5005
R11983 VPWR.n2386 VPWR.n2385 4.5005
R11984 VPWR.n455 VPWR.n398 4.5005
R11985 VPWR.n2439 VPWR.n2438 4.5005
R11986 VPWR.n322 VPWR.n84 4.5005
R11987 VPWR.n2594 VPWR.n2593 4.5005
R11988 VPWR.n2602 VPWR.n2601 4.5005
R11989 VPWR.n2606 VPWR.n2605 4.5005
R11990 VPWR.n314 VPWR.n78 4.5005
R11991 VPWR.n2429 VPWR.n2428 4.5005
R11992 VPWR.n463 VPWR.n402 4.5005
R11993 VPWR.n2396 VPWR.n2395 4.5005
R11994 VPWR.n506 VPWR.n473 4.5005
R11995 VPWR.n2233 VPWR.n2232 4.5005
R11996 VPWR.n655 VPWR.n594 4.5005
R11997 VPWR.n2200 VPWR.n2199 4.5005
R11998 VPWR.n698 VPWR.n665 4.5005
R11999 VPWR.n2037 VPWR.n2036 4.5005
R12000 VPWR.n847 VPWR.n786 4.5005
R12001 VPWR.n2004 VPWR.n2003 4.5005
R12002 VPWR.n890 VPWR.n857 4.5005
R12003 VPWR.n1841 VPWR.n1840 4.5005
R12004 VPWR.n1039 VPWR.n978 4.5005
R12005 VPWR.n1808 VPWR.n1807 4.5005
R12006 VPWR.n1755 VPWR.n1056 4.5005
R12007 VPWR.n1251 VPWR.n1140 4.5005
R12008 VPWR.n1485 VPWR.n1484 4.5005
R12009 VPWR.n983 VPWR.n950 4.5005
R12010 VPWR.n1911 VPWR.n1910 4.5005
R12011 VPWR.n948 VPWR.n947 4.5005
R12012 VPWR.n1934 VPWR.n1933 4.5005
R12013 VPWR.n791 VPWR.n758 4.5005
R12014 VPWR.n2107 VPWR.n2106 4.5005
R12015 VPWR.n756 VPWR.n755 4.5005
R12016 VPWR.n2130 VPWR.n2129 4.5005
R12017 VPWR.n599 VPWR.n566 4.5005
R12018 VPWR.n2303 VPWR.n2302 4.5005
R12019 VPWR.n564 VPWR.n563 4.5005
R12020 VPWR.n2326 VPWR.n2325 4.5005
R12021 VPWR.n407 VPWR.n374 4.5005
R12022 VPWR.n2499 VPWR.n2498 4.5005
R12023 VPWR.n372 VPWR.n371 4.5005
R12024 VPWR.n2522 VPWR.n2521 4.5005
R12025 VPWR.n2613 VPWR.n2612 4.5005
R12026 VPWR.n311 VPWR.n41 4.5005
R12027 VPWR.n2424 VPWR.n2423 4.5005
R12028 VPWR.n468 VPWR.n467 4.5005
R12029 VPWR.n2401 VPWR.n2400 4.5005
R12030 VPWR.n503 VPWR.n470 4.5005
R12031 VPWR.n2228 VPWR.n2227 4.5005
R12032 VPWR.n660 VPWR.n659 4.5005
R12033 VPWR.n2205 VPWR.n2204 4.5005
R12034 VPWR.n695 VPWR.n662 4.5005
R12035 VPWR.n2032 VPWR.n2031 4.5005
R12036 VPWR.n852 VPWR.n851 4.5005
R12037 VPWR.n2009 VPWR.n2008 4.5005
R12038 VPWR.n887 VPWR.n854 4.5005
R12039 VPWR.n1836 VPWR.n1835 4.5005
R12040 VPWR.n1044 VPWR.n1043 4.5005
R12041 VPWR.n1813 VPWR.n1812 4.5005
R12042 VPWR.n1079 VPWR.n1047 4.5005
R12043 VPWR.n2647 VPWR 4.49965
R12044 VPWR.n19 VPWR.n18 4.20017
R12045 VPWR.n1274 VPWR.n1273 4.20017
R12046 VPWR.n1298 VPWR.n1297 4.20017
R12047 VPWR.n1321 VPWR.n1320 4.20017
R12048 VPWR.n1356 VPWR.n1355 4.20017
R12049 VPWR.n1395 VPWR.n1394 4.20017
R12050 VPWR.n1433 VPWR.n1432 4.20017
R12051 VPWR.n2832 VPWR 4.14027
R12052 VPWR.n2816 VPWR 4.14027
R12053 VPWR.n2797 VPWR 4.14027
R12054 VPWR.n2777 VPWR 4.14027
R12055 VPWR.n2758 VPWR 4.14027
R12056 VPWR.n2722 VPWR 4.14027
R12057 VPWR.n2684 VPWR 4.14027
R12058 VPWR.n74 VPWR.n73 4.0005
R12059 VPWR.n2735 VPWR.n2732 3.76521
R12060 VPWR.n2699 VPWR.n2695 3.76521
R12061 VPWR.n2662 VPWR.n2658 3.76521
R12062 VPWR.n2630 VPWR.n2629 3.76521
R12063 VPWR.n37 VPWR 3.57245
R12064 VPWR.n1925 VPWR.n877 3.4105
R12065 VPWR.n1953 VPWR.n1952 3.4105
R12066 VPWR.n2016 VPWR.n766 3.4105
R12067 VPWR.n2088 VPWR.n2087 3.4105
R12068 VPWR.n2121 VPWR.n685 3.4105
R12069 VPWR.n2149 VPWR.n2148 3.4105
R12070 VPWR.n2212 VPWR.n574 3.4105
R12071 VPWR.n2284 VPWR.n2283 3.4105
R12072 VPWR.n2317 VPWR.n493 3.4105
R12073 VPWR.n2345 VPWR.n2344 3.4105
R12074 VPWR.n2408 VPWR.n382 3.4105
R12075 VPWR.n2407 VPWR.n381 3.4105
R12076 VPWR.n2343 VPWR.n2342 3.4105
R12077 VPWR.n2318 VPWR.n494 3.4105
R12078 VPWR.n2286 VPWR.n2285 3.4105
R12079 VPWR.n2211 VPWR.n573 3.4105
R12080 VPWR.n2147 VPWR.n2146 3.4105
R12081 VPWR.n2122 VPWR.n686 3.4105
R12082 VPWR.n2090 VPWR.n2089 3.4105
R12083 VPWR.n2015 VPWR.n765 3.4105
R12084 VPWR.n1951 VPWR.n1950 3.4105
R12085 VPWR.n1926 VPWR.n878 3.4105
R12086 VPWR.n1894 VPWR.n1893 3.4105
R12087 VPWR.n1892 VPWR.n1891 3.4105
R12088 VPWR.n1884 VPWR.n1883 3.4105
R12089 VPWR.n1924 VPWR.n874 3.4105
R12090 VPWR.n1961 VPWR.n1960 3.4105
R12091 VPWR.n2017 VPWR.n769 3.4105
R12092 VPWR.n2080 VPWR.n2079 3.4105
R12093 VPWR.n2120 VPWR.n682 3.4105
R12094 VPWR.n2157 VPWR.n2156 3.4105
R12095 VPWR.n2213 VPWR.n577 3.4105
R12096 VPWR.n2276 VPWR.n2275 3.4105
R12097 VPWR.n2316 VPWR.n490 3.4105
R12098 VPWR.n2353 VPWR.n2352 3.4105
R12099 VPWR.n2409 VPWR.n385 3.4105
R12100 VPWR.n2410 VPWR.n386 3.4105
R12101 VPWR.n2355 VPWR.n2354 3.4105
R12102 VPWR.n2315 VPWR.n489 3.4105
R12103 VPWR.n2274 VPWR.n2273 3.4105
R12104 VPWR.n2214 VPWR.n578 3.4105
R12105 VPWR.n2159 VPWR.n2158 3.4105
R12106 VPWR.n2119 VPWR.n681 3.4105
R12107 VPWR.n2078 VPWR.n2077 3.4105
R12108 VPWR.n2018 VPWR.n770 3.4105
R12109 VPWR.n1963 VPWR.n1962 3.4105
R12110 VPWR.n1923 VPWR.n873 3.4105
R12111 VPWR.n1882 VPWR.n1881 3.4105
R12112 VPWR.n1874 VPWR.n1873 3.4105
R12113 VPWR.n1922 VPWR.n870 3.4105
R12114 VPWR.n1971 VPWR.n1970 3.4105
R12115 VPWR.n2019 VPWR.n773 3.4105
R12116 VPWR.n2070 VPWR.n2069 3.4105
R12117 VPWR.n2118 VPWR.n678 3.4105
R12118 VPWR.n2167 VPWR.n2166 3.4105
R12119 VPWR.n2215 VPWR.n581 3.4105
R12120 VPWR.n2266 VPWR.n2265 3.4105
R12121 VPWR.n2314 VPWR.n486 3.4105
R12122 VPWR.n2363 VPWR.n2362 3.4105
R12123 VPWR.n2411 VPWR.n389 3.4105
R12124 VPWR.n2462 VPWR.n2461 3.4105
R12125 VPWR.n2470 VPWR.n2469 3.4105
R12126 VPWR.n2472 VPWR.n2471 3.4105
R12127 VPWR.n2480 VPWR.n2479 3.4105
R12128 VPWR.n2482 VPWR.n2481 3.4105
R12129 VPWR.n2490 VPWR.n2489 3.4105
R12130 VPWR.n2406 VPWR.n378 3.4105
R12131 VPWR.n2335 VPWR.n2334 3.4105
R12132 VPWR.n2319 VPWR.n497 3.4105
R12133 VPWR.n2294 VPWR.n2293 3.4105
R12134 VPWR.n2210 VPWR.n570 3.4105
R12135 VPWR.n2139 VPWR.n2138 3.4105
R12136 VPWR.n2123 VPWR.n689 3.4105
R12137 VPWR.n2098 VPWR.n2097 3.4105
R12138 VPWR.n2014 VPWR.n762 3.4105
R12139 VPWR.n1943 VPWR.n1942 3.4105
R12140 VPWR.n1927 VPWR.n881 3.4105
R12141 VPWR.n1902 VPWR.n1901 3.4105
R12142 VPWR.n1818 VPWR.n954 3.4105
R12143 VPWR.n1819 VPWR.n957 3.4105
R12144 VPWR.n1820 VPWR.n958 3.4105
R12145 VPWR.n1821 VPWR.n961 3.4105
R12146 VPWR.n1822 VPWR.n962 3.4105
R12147 VPWR.n1823 VPWR.n965 3.4105
R12148 VPWR.n1824 VPWR.n966 3.4105
R12149 VPWR.n1872 VPWR.n1871 3.4105
R12150 VPWR.n1921 VPWR.n869 3.4105
R12151 VPWR.n1973 VPWR.n1972 3.4105
R12152 VPWR.n2020 VPWR.n774 3.4105
R12153 VPWR.n2068 VPWR.n2067 3.4105
R12154 VPWR.n2117 VPWR.n677 3.4105
R12155 VPWR.n2169 VPWR.n2168 3.4105
R12156 VPWR.n2216 VPWR.n582 3.4105
R12157 VPWR.n2264 VPWR.n2263 3.4105
R12158 VPWR.n2313 VPWR.n485 3.4105
R12159 VPWR.n2365 VPWR.n2364 3.4105
R12160 VPWR.n2412 VPWR.n390 3.4105
R12161 VPWR.n2460 VPWR.n2459 3.4105
R12162 VPWR.n2452 VPWR.n2451 3.4105
R12163 VPWR.n2413 VPWR.n393 3.4105
R12164 VPWR.n2373 VPWR.n2372 3.4105
R12165 VPWR.n2312 VPWR.n482 3.4105
R12166 VPWR.n2256 VPWR.n2255 3.4105
R12167 VPWR.n2217 VPWR.n585 3.4105
R12168 VPWR.n2177 VPWR.n2176 3.4105
R12169 VPWR.n2116 VPWR.n674 3.4105
R12170 VPWR.n2060 VPWR.n2059 3.4105
R12171 VPWR.n2021 VPWR.n777 3.4105
R12172 VPWR.n1981 VPWR.n1980 3.4105
R12173 VPWR.n1920 VPWR.n866 3.4105
R12174 VPWR.n1864 VPWR.n1863 3.4105
R12175 VPWR.n1825 VPWR.n969 3.4105
R12176 VPWR.n1817 VPWR.n953 3.4105
R12177 VPWR.n1904 VPWR.n1903 3.4105
R12178 VPWR.n1928 VPWR.n882 3.4105
R12179 VPWR.n1941 VPWR.n1940 3.4105
R12180 VPWR.n2013 VPWR.n761 3.4105
R12181 VPWR.n2100 VPWR.n2099 3.4105
R12182 VPWR.n2124 VPWR.n690 3.4105
R12183 VPWR.n2137 VPWR.n2136 3.4105
R12184 VPWR.n2209 VPWR.n569 3.4105
R12185 VPWR.n2296 VPWR.n2295 3.4105
R12186 VPWR.n2320 VPWR.n498 3.4105
R12187 VPWR.n2333 VPWR.n2332 3.4105
R12188 VPWR.n2405 VPWR.n377 3.4105
R12189 VPWR.n2492 VPWR.n2491 3.4105
R12190 VPWR.n2516 VPWR.n115 3.4105
R12191 VPWR.n2515 VPWR.n114 3.4105
R12192 VPWR.n2514 VPWR.n109 3.4105
R12193 VPWR.n2513 VPWR.n108 3.4105
R12194 VPWR.n2512 VPWR.n103 3.4105
R12195 VPWR.n2511 VPWR.n102 3.4105
R12196 VPWR.n2510 VPWR.n97 3.4105
R12197 VPWR.n2509 VPWR.n96 3.4105
R12198 VPWR.n2508 VPWR.n91 3.4105
R12199 VPWR.n2507 VPWR.n90 3.4105
R12200 VPWR.n2450 VPWR.n2449 3.4105
R12201 VPWR.n2414 VPWR.n394 3.4105
R12202 VPWR.n2375 VPWR.n2374 3.4105
R12203 VPWR.n2311 VPWR.n481 3.4105
R12204 VPWR.n2254 VPWR.n2253 3.4105
R12205 VPWR.n2218 VPWR.n586 3.4105
R12206 VPWR.n2179 VPWR.n2178 3.4105
R12207 VPWR.n2115 VPWR.n673 3.4105
R12208 VPWR.n2058 VPWR.n2057 3.4105
R12209 VPWR.n2022 VPWR.n778 3.4105
R12210 VPWR.n1983 VPWR.n1982 3.4105
R12211 VPWR.n1919 VPWR.n865 3.4105
R12212 VPWR.n1862 VPWR.n1861 3.4105
R12213 VPWR.n1826 VPWR.n970 3.4105
R12214 VPWR.n1551 VPWR.n1162 3.4105
R12215 VPWR.n1559 VPWR.n1558 3.4105
R12216 VPWR.n1544 VPWR.n1543 3.4105
R12217 VPWR.n1536 VPWR.n1535 3.4105
R12218 VPWR.n1530 VPWR.n1529 3.4105
R12219 VPWR.n1522 VPWR.n1521 3.4105
R12220 VPWR.n1516 VPWR.n1515 3.4105
R12221 VPWR.n1508 VPWR.n1151 3.4105
R12222 VPWR.n1604 VPWR.n1603 3.4105
R12223 VPWR.n1471 VPWR.n1147 3.4105
R12224 VPWR.n1784 VPWR.n1783 3.4105
R12225 VPWR.n1827 VPWR.n973 3.4105
R12226 VPWR.n1854 VPWR.n1853 3.4105
R12227 VPWR.n1918 VPWR.n862 3.4105
R12228 VPWR.n1991 VPWR.n1990 3.4105
R12229 VPWR.n2023 VPWR.n781 3.4105
R12230 VPWR.n2050 VPWR.n2049 3.4105
R12231 VPWR.n2114 VPWR.n670 3.4105
R12232 VPWR.n2187 VPWR.n2186 3.4105
R12233 VPWR.n2219 VPWR.n589 3.4105
R12234 VPWR.n2246 VPWR.n2245 3.4105
R12235 VPWR.n2310 VPWR.n478 3.4105
R12236 VPWR.n2383 VPWR.n2382 3.4105
R12237 VPWR.n2415 VPWR.n397 3.4105
R12238 VPWR.n2442 VPWR.n2441 3.4105
R12239 VPWR.n2506 VPWR.n85 3.4105
R12240 VPWR.n2504 VPWR.n79 3.4105
R12241 VPWR.n2432 VPWR.n2431 3.4105
R12242 VPWR.n2417 VPWR.n401 3.4105
R12243 VPWR.n2393 VPWR.n2392 3.4105
R12244 VPWR.n2308 VPWR.n474 3.4105
R12245 VPWR.n2236 VPWR.n2235 3.4105
R12246 VPWR.n2221 VPWR.n593 3.4105
R12247 VPWR.n2197 VPWR.n2196 3.4105
R12248 VPWR.n2112 VPWR.n666 3.4105
R12249 VPWR.n2040 VPWR.n2039 3.4105
R12250 VPWR.n2025 VPWR.n785 3.4105
R12251 VPWR.n2001 VPWR.n2000 3.4105
R12252 VPWR.n1916 VPWR.n858 3.4105
R12253 VPWR.n1844 VPWR.n1843 3.4105
R12254 VPWR.n1829 VPWR.n977 3.4105
R12255 VPWR.n1771 VPWR.n1763 3.4105
R12256 VPWR.n1776 VPWR.n1062 3.4105
R12257 VPWR.n1828 VPWR.n974 3.4105
R12258 VPWR.n1852 VPWR.n1851 3.4105
R12259 VPWR.n1917 VPWR.n861 3.4105
R12260 VPWR.n1993 VPWR.n1992 3.4105
R12261 VPWR.n2024 VPWR.n782 3.4105
R12262 VPWR.n2048 VPWR.n2047 3.4105
R12263 VPWR.n2113 VPWR.n669 3.4105
R12264 VPWR.n2189 VPWR.n2188 3.4105
R12265 VPWR.n2220 VPWR.n590 3.4105
R12266 VPWR.n2244 VPWR.n2243 3.4105
R12267 VPWR.n2309 VPWR.n477 3.4105
R12268 VPWR.n2385 VPWR.n2384 3.4105
R12269 VPWR.n2416 VPWR.n398 3.4105
R12270 VPWR.n2440 VPWR.n2439 3.4105
R12271 VPWR.n2505 VPWR.n84 3.4105
R12272 VPWR.n2503 VPWR.n78 3.4105
R12273 VPWR.n2430 VPWR.n2429 3.4105
R12274 VPWR.n2418 VPWR.n402 3.4105
R12275 VPWR.n2395 VPWR.n2394 3.4105
R12276 VPWR.n2307 VPWR.n473 3.4105
R12277 VPWR.n2234 VPWR.n2233 3.4105
R12278 VPWR.n2222 VPWR.n594 3.4105
R12279 VPWR.n2199 VPWR.n2198 3.4105
R12280 VPWR.n2111 VPWR.n665 3.4105
R12281 VPWR.n2038 VPWR.n2037 3.4105
R12282 VPWR.n2026 VPWR.n786 3.4105
R12283 VPWR.n2003 VPWR.n2002 3.4105
R12284 VPWR.n1915 VPWR.n857 3.4105
R12285 VPWR.n1842 VPWR.n1841 3.4105
R12286 VPWR.n1830 VPWR.n978 3.4105
R12287 VPWR.n1807 VPWR.n1806 3.4105
R12288 VPWR.n1484 VPWR.n1483 3.4105
R12289 VPWR.n1816 VPWR.n950 3.4105
R12290 VPWR.n1912 VPWR.n1911 3.4105
R12291 VPWR.n1929 VPWR.n948 3.4105
R12292 VPWR.n1933 VPWR.n1932 3.4105
R12293 VPWR.n2012 VPWR.n758 3.4105
R12294 VPWR.n2108 VPWR.n2107 3.4105
R12295 VPWR.n2125 VPWR.n756 3.4105
R12296 VPWR.n2129 VPWR.n2128 3.4105
R12297 VPWR.n2208 VPWR.n566 3.4105
R12298 VPWR.n2304 VPWR.n2303 3.4105
R12299 VPWR.n2321 VPWR.n564 3.4105
R12300 VPWR.n2325 VPWR.n2324 3.4105
R12301 VPWR.n2404 VPWR.n374 3.4105
R12302 VPWR.n2500 VPWR.n2499 3.4105
R12303 VPWR.n2517 VPWR.n372 3.4105
R12304 VPWR.n2521 VPWR.n2520 3.4105
R12305 VPWR.n2531 VPWR.n2530 3.4105
R12306 VPWR.n2533 VPWR.n2532 3.4105
R12307 VPWR.n2543 VPWR.n2542 3.4105
R12308 VPWR.n2545 VPWR.n2544 3.4105
R12309 VPWR.n2555 VPWR.n2554 3.4105
R12310 VPWR.n2557 VPWR.n2556 3.4105
R12311 VPWR.n2567 VPWR.n2566 3.4105
R12312 VPWR.n2569 VPWR.n2568 3.4105
R12313 VPWR.n2579 VPWR.n2578 3.4105
R12314 VPWR.n2581 VPWR.n2580 3.4105
R12315 VPWR.n2591 VPWR.n2590 3.4105
R12316 VPWR.n2593 VPWR.n2592 3.4105
R12317 VPWR.n2603 VPWR.n2602 3.4105
R12318 VPWR.n2605 VPWR.n2604 3.4105
R12319 VPWR.n2614 VPWR.n2613 3.4105
R12320 VPWR.n2502 VPWR.n41 3.4105
R12321 VPWR.n2423 VPWR.n2422 3.4105
R12322 VPWR.n2419 VPWR.n468 3.4105
R12323 VPWR.n2402 VPWR.n2401 3.4105
R12324 VPWR.n2306 VPWR.n470 3.4105
R12325 VPWR.n2227 VPWR.n2226 3.4105
R12326 VPWR.n2223 VPWR.n660 3.4105
R12327 VPWR.n2206 VPWR.n2205 3.4105
R12328 VPWR.n2110 VPWR.n662 3.4105
R12329 VPWR.n2031 VPWR.n2030 3.4105
R12330 VPWR.n2027 VPWR.n852 3.4105
R12331 VPWR.n2010 VPWR.n2009 3.4105
R12332 VPWR.n1914 VPWR.n854 3.4105
R12333 VPWR.n1835 VPWR.n1834 3.4105
R12334 VPWR.n1831 VPWR.n1044 3.4105
R12335 VPWR.n1814 VPWR.n1813 3.4105
R12336 VPWR.n1074 VPWR.n1047 3.4105
R12337 VPWR.n1075 VPWR.n1056 3.4105
R12338 VPWR.n1773 VPWR.n1772 3.4105
R12339 VPWR.n1775 VPWR.n1774 3.4105
R12340 VPWR.n1548 VPWR.n1064 3.4105
R12341 VPWR.n1550 VPWR.n1549 3.4105
R12342 VPWR.n1547 VPWR.n1164 3.4105
R12343 VPWR.n1546 VPWR.n1545 3.4105
R12344 VPWR.n1534 VPWR.n1533 3.4105
R12345 VPWR.n1532 VPWR.n1531 3.4105
R12346 VPWR.n1520 VPWR.n1519 3.4105
R12347 VPWR.n1518 VPWR.n1517 3.4105
R12348 VPWR.n1507 VPWR.n1506 3.4105
R12349 VPWR.n1606 VPWR.n1605 3.4105
R12350 VPWR.n1608 VPWR.n1607 3.4105
R12351 VPWR.n1467 VPWR.n1251 3.4105
R12352 VPWR.n1364 VPWR.n1360 3.38874
R12353 VPWR.n1403 VPWR.n1399 3.38874
R12354 VPWR.n1440 VPWR.n1436 3.38874
R12355 VPWR.n47 VPWR.n45 3.36211
R12356 VPWR.n49 VPWR.n47 3.36211
R12357 VPWR.n51 VPWR.n49 3.36211
R12358 VPWR.n53 VPWR.n51 3.36211
R12359 VPWR.n55 VPWR.n53 3.36211
R12360 VPWR.n57 VPWR.n55 3.36211
R12361 VPWR.n59 VPWR.n57 3.36211
R12362 VPWR.n61 VPWR.n59 3.36211
R12363 VPWR.n63 VPWR.n61 3.36211
R12364 VPWR.n65 VPWR.n63 3.36211
R12365 VPWR.n67 VPWR.n65 3.36211
R12366 VPWR.n69 VPWR.n67 3.36211
R12367 VPWR.n71 VPWR.n69 3.36211
R12368 VPWR.n73 VPWR.n71 3.36211
R12369 VPWR.t468 VPWR.t299 3.35739
R12370 VPWR.t737 VPWR.t490 3.35739
R12371 VPWR.n2590 VPWR.n85 3.28012
R12372 VPWR.n2530 VPWR.n115 3.28012
R12373 VPWR.n2569 VPWR.n96 3.28012
R12374 VPWR.n2459 VPWR.n96 3.28012
R12375 VPWR.n2566 VPWR.n97 3.28012
R12376 VPWR.n2462 VPWR.n97 3.28012
R12377 VPWR.n2554 VPWR.n103 3.28012
R12378 VPWR.n2472 VPWR.n103 3.28012
R12379 VPWR.n2472 VPWR.n385 3.28012
R12380 VPWR.n2545 VPWR.n108 3.28012
R12381 VPWR.n2479 VPWR.n108 3.28012
R12382 VPWR.n2479 VPWR.n382 3.28012
R12383 VPWR.n1517 VPWR.n1516 3.28012
R12384 VPWR.n1516 VPWR.n958 3.28012
R12385 VPWR.n1891 VPWR.n958 3.28012
R12386 VPWR.n1891 VPWR.n877 3.28012
R12387 VPWR.n1953 VPWR.n877 3.28012
R12388 VPWR.n1953 VPWR.n766 3.28012
R12389 VPWR.n2087 VPWR.n766 3.28012
R12390 VPWR.n2087 VPWR.n685 3.28012
R12391 VPWR.n2149 VPWR.n685 3.28012
R12392 VPWR.n2149 VPWR.n574 3.28012
R12393 VPWR.n2283 VPWR.n574 3.28012
R12394 VPWR.n2283 VPWR.n493 3.28012
R12395 VPWR.n2345 VPWR.n493 3.28012
R12396 VPWR.n2345 VPWR.n382 3.28012
R12397 VPWR.n2542 VPWR.n109 3.28012
R12398 VPWR.n2482 VPWR.n109 3.28012
R12399 VPWR.n2482 VPWR.n381 3.28012
R12400 VPWR.n2342 VPWR.n381 3.28012
R12401 VPWR.n2342 VPWR.n494 3.28012
R12402 VPWR.n2286 VPWR.n494 3.28012
R12403 VPWR.n2286 VPWR.n573 3.28012
R12404 VPWR.n2146 VPWR.n573 3.28012
R12405 VPWR.n2146 VPWR.n686 3.28012
R12406 VPWR.n2090 VPWR.n686 3.28012
R12407 VPWR.n2090 VPWR.n765 3.28012
R12408 VPWR.n1950 VPWR.n765 3.28012
R12409 VPWR.n1950 VPWR.n878 3.28012
R12410 VPWR.n1894 VPWR.n878 3.28012
R12411 VPWR.n1508 VPWR.n1507 3.28012
R12412 VPWR.n1508 VPWR.n957 3.28012
R12413 VPWR.n1894 VPWR.n957 3.28012
R12414 VPWR.n1522 VPWR.n1520 3.28012
R12415 VPWR.n1522 VPWR.n961 3.28012
R12416 VPWR.n1884 VPWR.n961 3.28012
R12417 VPWR.n1884 VPWR.n874 3.28012
R12418 VPWR.n1960 VPWR.n874 3.28012
R12419 VPWR.n1960 VPWR.n769 3.28012
R12420 VPWR.n2080 VPWR.n769 3.28012
R12421 VPWR.n2080 VPWR.n682 3.28012
R12422 VPWR.n2156 VPWR.n682 3.28012
R12423 VPWR.n2156 VPWR.n577 3.28012
R12424 VPWR.n2276 VPWR.n577 3.28012
R12425 VPWR.n2276 VPWR.n490 3.28012
R12426 VPWR.n2352 VPWR.n490 3.28012
R12427 VPWR.n2352 VPWR.n385 3.28012
R12428 VPWR.n2557 VPWR.n102 3.28012
R12429 VPWR.n2469 VPWR.n102 3.28012
R12430 VPWR.n2469 VPWR.n386 3.28012
R12431 VPWR.n2355 VPWR.n386 3.28012
R12432 VPWR.n2355 VPWR.n489 3.28012
R12433 VPWR.n2273 VPWR.n489 3.28012
R12434 VPWR.n2273 VPWR.n578 3.28012
R12435 VPWR.n2159 VPWR.n578 3.28012
R12436 VPWR.n2159 VPWR.n681 3.28012
R12437 VPWR.n2077 VPWR.n681 3.28012
R12438 VPWR.n2077 VPWR.n770 3.28012
R12439 VPWR.n1963 VPWR.n770 3.28012
R12440 VPWR.n1963 VPWR.n873 3.28012
R12441 VPWR.n1881 VPWR.n873 3.28012
R12442 VPWR.n1531 VPWR.n1530 3.28012
R12443 VPWR.n1530 VPWR.n962 3.28012
R12444 VPWR.n1881 VPWR.n962 3.28012
R12445 VPWR.n1536 VPWR.n1534 3.28012
R12446 VPWR.n1536 VPWR.n965 3.28012
R12447 VPWR.n1874 VPWR.n965 3.28012
R12448 VPWR.n1874 VPWR.n870 3.28012
R12449 VPWR.n1970 VPWR.n870 3.28012
R12450 VPWR.n1970 VPWR.n773 3.28012
R12451 VPWR.n2070 VPWR.n773 3.28012
R12452 VPWR.n2070 VPWR.n678 3.28012
R12453 VPWR.n2166 VPWR.n678 3.28012
R12454 VPWR.n2166 VPWR.n581 3.28012
R12455 VPWR.n2266 VPWR.n581 3.28012
R12456 VPWR.n2266 VPWR.n486 3.28012
R12457 VPWR.n2362 VPWR.n486 3.28012
R12458 VPWR.n2362 VPWR.n389 3.28012
R12459 VPWR.n2462 VPWR.n389 3.28012
R12460 VPWR.n2533 VPWR.n114 3.28012
R12461 VPWR.n2489 VPWR.n114 3.28012
R12462 VPWR.n2489 VPWR.n378 3.28012
R12463 VPWR.n2335 VPWR.n378 3.28012
R12464 VPWR.n2335 VPWR.n497 3.28012
R12465 VPWR.n2293 VPWR.n497 3.28012
R12466 VPWR.n2293 VPWR.n570 3.28012
R12467 VPWR.n2139 VPWR.n570 3.28012
R12468 VPWR.n2139 VPWR.n689 3.28012
R12469 VPWR.n2097 VPWR.n689 3.28012
R12470 VPWR.n2097 VPWR.n762 3.28012
R12471 VPWR.n1943 VPWR.n762 3.28012
R12472 VPWR.n1943 VPWR.n881 3.28012
R12473 VPWR.n1901 VPWR.n881 3.28012
R12474 VPWR.n1901 VPWR.n954 3.28012
R12475 VPWR.n1605 VPWR.n1604 3.28012
R12476 VPWR.n1604 VPWR.n954 3.28012
R12477 VPWR.n1545 VPWR.n1544 3.28012
R12478 VPWR.n1544 VPWR.n966 3.28012
R12479 VPWR.n1871 VPWR.n966 3.28012
R12480 VPWR.n1871 VPWR.n869 3.28012
R12481 VPWR.n1973 VPWR.n869 3.28012
R12482 VPWR.n1973 VPWR.n774 3.28012
R12483 VPWR.n2067 VPWR.n774 3.28012
R12484 VPWR.n2067 VPWR.n677 3.28012
R12485 VPWR.n2169 VPWR.n677 3.28012
R12486 VPWR.n2169 VPWR.n582 3.28012
R12487 VPWR.n2263 VPWR.n582 3.28012
R12488 VPWR.n2263 VPWR.n485 3.28012
R12489 VPWR.n2365 VPWR.n485 3.28012
R12490 VPWR.n2365 VPWR.n390 3.28012
R12491 VPWR.n2459 VPWR.n390 3.28012
R12492 VPWR.n2578 VPWR.n91 3.28012
R12493 VPWR.n2452 VPWR.n91 3.28012
R12494 VPWR.n2452 VPWR.n393 3.28012
R12495 VPWR.n2372 VPWR.n393 3.28012
R12496 VPWR.n2372 VPWR.n482 3.28012
R12497 VPWR.n2256 VPWR.n482 3.28012
R12498 VPWR.n2256 VPWR.n585 3.28012
R12499 VPWR.n2176 VPWR.n585 3.28012
R12500 VPWR.n2176 VPWR.n674 3.28012
R12501 VPWR.n2060 VPWR.n674 3.28012
R12502 VPWR.n2060 VPWR.n777 3.28012
R12503 VPWR.n1980 VPWR.n777 3.28012
R12504 VPWR.n1980 VPWR.n866 3.28012
R12505 VPWR.n1864 VPWR.n866 3.28012
R12506 VPWR.n1864 VPWR.n969 3.28012
R12507 VPWR.n1558 VPWR.n1164 3.28012
R12508 VPWR.n1558 VPWR.n969 3.28012
R12509 VPWR.n1608 VPWR.n1147 3.28012
R12510 VPWR.n1147 VPWR.n953 3.28012
R12511 VPWR.n1904 VPWR.n953 3.28012
R12512 VPWR.n1904 VPWR.n882 3.28012
R12513 VPWR.n1940 VPWR.n882 3.28012
R12514 VPWR.n1940 VPWR.n761 3.28012
R12515 VPWR.n2100 VPWR.n761 3.28012
R12516 VPWR.n2100 VPWR.n690 3.28012
R12517 VPWR.n2136 VPWR.n690 3.28012
R12518 VPWR.n2136 VPWR.n569 3.28012
R12519 VPWR.n2296 VPWR.n569 3.28012
R12520 VPWR.n2296 VPWR.n498 3.28012
R12521 VPWR.n2332 VPWR.n498 3.28012
R12522 VPWR.n2332 VPWR.n377 3.28012
R12523 VPWR.n2492 VPWR.n377 3.28012
R12524 VPWR.n2492 VPWR.n115 3.28012
R12525 VPWR.n2581 VPWR.n90 3.28012
R12526 VPWR.n2449 VPWR.n90 3.28012
R12527 VPWR.n2449 VPWR.n394 3.28012
R12528 VPWR.n2375 VPWR.n394 3.28012
R12529 VPWR.n2375 VPWR.n481 3.28012
R12530 VPWR.n2253 VPWR.n481 3.28012
R12531 VPWR.n2253 VPWR.n586 3.28012
R12532 VPWR.n2179 VPWR.n586 3.28012
R12533 VPWR.n2179 VPWR.n673 3.28012
R12534 VPWR.n2057 VPWR.n673 3.28012
R12535 VPWR.n2057 VPWR.n778 3.28012
R12536 VPWR.n1983 VPWR.n778 3.28012
R12537 VPWR.n1983 VPWR.n865 3.28012
R12538 VPWR.n1861 VPWR.n865 3.28012
R12539 VPWR.n1861 VPWR.n970 3.28012
R12540 VPWR.n1551 VPWR.n970 3.28012
R12541 VPWR.n1551 VPWR.n1550 3.28012
R12542 VPWR.n1783 VPWR.n1064 3.28012
R12543 VPWR.n1783 VPWR.n973 3.28012
R12544 VPWR.n1854 VPWR.n973 3.28012
R12545 VPWR.n1854 VPWR.n862 3.28012
R12546 VPWR.n1990 VPWR.n862 3.28012
R12547 VPWR.n1990 VPWR.n781 3.28012
R12548 VPWR.n2050 VPWR.n781 3.28012
R12549 VPWR.n2050 VPWR.n670 3.28012
R12550 VPWR.n2186 VPWR.n670 3.28012
R12551 VPWR.n2186 VPWR.n589 3.28012
R12552 VPWR.n2246 VPWR.n589 3.28012
R12553 VPWR.n2246 VPWR.n478 3.28012
R12554 VPWR.n2382 VPWR.n478 3.28012
R12555 VPWR.n2382 VPWR.n397 3.28012
R12556 VPWR.n2442 VPWR.n397 3.28012
R12557 VPWR.n2442 VPWR.n85 3.28012
R12558 VPWR.n2602 VPWR.n79 3.28012
R12559 VPWR.n2432 VPWR.n79 3.28012
R12560 VPWR.n2432 VPWR.n401 3.28012
R12561 VPWR.n2392 VPWR.n401 3.28012
R12562 VPWR.n2392 VPWR.n474 3.28012
R12563 VPWR.n2236 VPWR.n474 3.28012
R12564 VPWR.n2236 VPWR.n593 3.28012
R12565 VPWR.n2196 VPWR.n593 3.28012
R12566 VPWR.n2196 VPWR.n666 3.28012
R12567 VPWR.n2040 VPWR.n666 3.28012
R12568 VPWR.n2040 VPWR.n785 3.28012
R12569 VPWR.n2000 VPWR.n785 3.28012
R12570 VPWR.n2000 VPWR.n858 3.28012
R12571 VPWR.n1844 VPWR.n858 3.28012
R12572 VPWR.n1844 VPWR.n977 3.28012
R12573 VPWR.n1771 VPWR.n977 3.28012
R12574 VPWR.n1772 VPWR.n1771 3.28012
R12575 VPWR.n1776 VPWR.n1775 3.28012
R12576 VPWR.n1776 VPWR.n974 3.28012
R12577 VPWR.n1851 VPWR.n974 3.28012
R12578 VPWR.n1851 VPWR.n861 3.28012
R12579 VPWR.n1993 VPWR.n861 3.28012
R12580 VPWR.n1993 VPWR.n782 3.28012
R12581 VPWR.n2047 VPWR.n782 3.28012
R12582 VPWR.n2047 VPWR.n669 3.28012
R12583 VPWR.n2189 VPWR.n669 3.28012
R12584 VPWR.n2189 VPWR.n590 3.28012
R12585 VPWR.n2243 VPWR.n590 3.28012
R12586 VPWR.n2243 VPWR.n477 3.28012
R12587 VPWR.n2385 VPWR.n477 3.28012
R12588 VPWR.n2385 VPWR.n398 3.28012
R12589 VPWR.n2439 VPWR.n398 3.28012
R12590 VPWR.n2439 VPWR.n84 3.28012
R12591 VPWR.n2593 VPWR.n84 3.28012
R12592 VPWR.n2605 VPWR.n78 3.28012
R12593 VPWR.n2429 VPWR.n78 3.28012
R12594 VPWR.n2429 VPWR.n402 3.28012
R12595 VPWR.n2395 VPWR.n402 3.28012
R12596 VPWR.n2395 VPWR.n473 3.28012
R12597 VPWR.n2233 VPWR.n473 3.28012
R12598 VPWR.n2233 VPWR.n594 3.28012
R12599 VPWR.n2199 VPWR.n594 3.28012
R12600 VPWR.n2199 VPWR.n665 3.28012
R12601 VPWR.n2037 VPWR.n665 3.28012
R12602 VPWR.n2037 VPWR.n786 3.28012
R12603 VPWR.n2003 VPWR.n786 3.28012
R12604 VPWR.n2003 VPWR.n857 3.28012
R12605 VPWR.n1841 VPWR.n857 3.28012
R12606 VPWR.n1841 VPWR.n978 3.28012
R12607 VPWR.n1807 VPWR.n978 3.28012
R12608 VPWR.n1807 VPWR.n1056 3.28012
R12609 VPWR.n1484 VPWR.n1251 3.28012
R12610 VPWR.n1484 VPWR.n950 3.28012
R12611 VPWR.n1911 VPWR.n950 3.28012
R12612 VPWR.n1911 VPWR.n948 3.28012
R12613 VPWR.n1933 VPWR.n948 3.28012
R12614 VPWR.n1933 VPWR.n758 3.28012
R12615 VPWR.n2107 VPWR.n758 3.28012
R12616 VPWR.n2107 VPWR.n756 3.28012
R12617 VPWR.n2129 VPWR.n756 3.28012
R12618 VPWR.n2129 VPWR.n566 3.28012
R12619 VPWR.n2303 VPWR.n566 3.28012
R12620 VPWR.n2303 VPWR.n564 3.28012
R12621 VPWR.n2325 VPWR.n564 3.28012
R12622 VPWR.n2325 VPWR.n374 3.28012
R12623 VPWR.n2499 VPWR.n374 3.28012
R12624 VPWR.n2499 VPWR.n372 3.28012
R12625 VPWR.n2521 VPWR.n372 3.28012
R12626 VPWR.n2423 VPWR.n41 3.28012
R12627 VPWR.n2423 VPWR.n468 3.28012
R12628 VPWR.n2401 VPWR.n468 3.28012
R12629 VPWR.n2401 VPWR.n470 3.28012
R12630 VPWR.n2227 VPWR.n470 3.28012
R12631 VPWR.n2227 VPWR.n660 3.28012
R12632 VPWR.n2205 VPWR.n660 3.28012
R12633 VPWR.n2205 VPWR.n662 3.28012
R12634 VPWR.n2031 VPWR.n662 3.28012
R12635 VPWR.n2031 VPWR.n852 3.28012
R12636 VPWR.n2009 VPWR.n852 3.28012
R12637 VPWR.n2009 VPWR.n854 3.28012
R12638 VPWR.n1835 VPWR.n854 3.28012
R12639 VPWR.n1835 VPWR.n1044 3.28012
R12640 VPWR.n1813 VPWR.n1044 3.28012
R12641 VPWR.n1813 VPWR.n1047 3.28012
R12642 VPWR.n2613 VPWR.n41 3.26393
R12643 VPWR.n1343 VPWR.n1341 3.01226
R12644 VPWR.n1347 VPWR.n1323 2.63579
R12645 VPWR.n2835 VPWR.t833 2.48308
R12646 VPWR.n2750 VPWR.n2749 2.25932
R12647 VPWR.n1466 VPWR.n1465 2.06026
R12648 VPWR.n1466 VPWR.n1045 1.78803
R12649 VPWR.n2403 VPWR.n2402 1.32852
R12650 VPWR.n2306 VPWR.n469 1.32852
R12651 VPWR.n2226 VPWR.n2225 1.32852
R12652 VPWR.n2224 VPWR.n2223 1.32852
R12653 VPWR.n2207 VPWR.n2206 1.32852
R12654 VPWR.n2110 VPWR.n661 1.32852
R12655 VPWR.n2030 VPWR.n2029 1.32852
R12656 VPWR.n2028 VPWR.n2027 1.32852
R12657 VPWR.n2011 VPWR.n2010 1.32852
R12658 VPWR.n1914 VPWR.n853 1.32852
R12659 VPWR.n2420 VPWR.n2419 1.32852
R12660 VPWR.n1834 VPWR.n1833 1.32852
R12661 VPWR.n2422 VPWR.n2421 1.32852
R12662 VPWR.n1832 VPWR.n1831 1.32852
R12663 VPWR.n2502 VPWR.n40 1.32852
R12664 VPWR.n1815 VPWR.n1814 1.32852
R12665 VPWR.n2615 VPWR.n2614 1.32852
R12666 VPWR.n1074 VPWR.n1045 1.32852
R12667 VPWR.n2857 VPWR.n23 1.29068
R12668 VPWR.n2843 VPWR.n21 1.28175
R12669 VPWR.n2501 VPWR 1.25994
R12670 VPWR VPWR.n373 1.25994
R12671 VPWR VPWR.n2323 1.25994
R12672 VPWR.n2322 VPWR 1.25994
R12673 VPWR.n2305 VPWR 1.25994
R12674 VPWR VPWR.n565 1.25994
R12675 VPWR VPWR.n2127 1.25994
R12676 VPWR.n2126 VPWR 1.25994
R12677 VPWR.n2109 VPWR 1.25994
R12678 VPWR VPWR.n757 1.25994
R12679 VPWR VPWR.n1931 1.25994
R12680 VPWR.n1930 VPWR 1.25994
R12681 VPWR.n1913 VPWR 1.25994
R12682 VPWR VPWR.n949 1.25994
R12683 VPWR.n2518 VPWR 1.25994
R12684 VPWR VPWR.n1469 1.25994
R12685 VPWR VPWR.n2519 1.25994
R12686 VPWR.n1468 VPWR 1.25994
R12687 VPWR.n2616 VPWR.n2615 1.144
R12688 VPWR.n2611 VPWR 0.925943
R12689 VPWR VPWR.n1082 0.925943
R12690 VPWR.n2588 VPWR.n86 0.904391
R12691 VPWR.n2528 VPWR.n116 0.904391
R12692 VPWR.n2571 VPWR.n95 0.904391
R12693 VPWR.n2564 VPWR.n98 0.904391
R12694 VPWR.n2552 VPWR.n104 0.904391
R12695 VPWR.n2547 VPWR.n107 0.904391
R12696 VPWR.n1241 VPWR.n1197 0.904391
R12697 VPWR.n2540 VPWR.n110 0.904391
R12698 VPWR.n1643 VPWR.n1121 0.904391
R12699 VPWR.n1659 VPWR.n1113 0.904391
R12700 VPWR.n2559 VPWR.n101 0.904391
R12701 VPWR.n1670 VPWR.n1111 0.904391
R12702 VPWR.n1230 VPWR.n1229 0.904391
R12703 VPWR.n2535 VPWR.n113 0.904391
R12704 VPWR.n1632 VPWR.n1123 0.904391
R12705 VPWR.n1686 VPWR.n1103 0.904391
R12706 VPWR.n2576 VPWR.n92 0.904391
R12707 VPWR.n1697 VPWR.n1101 0.904391
R12708 VPWR.n1610 VPWR.n1146 0.904391
R12709 VPWR.n2583 VPWR.n89 0.904391
R12710 VPWR.n1216 VPWR.n1215 0.904391
R12711 VPWR.n1713 VPWR.n1093 0.904391
R12712 VPWR.n1761 VPWR.n1076 0.904391
R12713 VPWR.n1724 VPWR.n1090 0.904391
R12714 VPWR.n2600 VPWR.n80 0.904391
R12715 VPWR.n2607 VPWR.n77 0.904391
R12716 VPWR.n1756 VPWR.n1754 0.904391
R12717 VPWR.n1616 VPWR.n1615 0.904391
R12718 VPWR.n2523 VPWR.n308 0.904391
R12719 VPWR.n2595 VPWR.n83 0.904391
R12720 VPWR.n2856 VPWR.n2855 0.711611
R12721 VPWR.n34 VPWR.n33 0.711611
R12722 VPWR.n159 VPWR.n83 0.675548
R12723 VPWR.n171 VPWR.n86 0.675548
R12724 VPWR.n183 VPWR.n89 0.675548
R12725 VPWR.n195 VPWR.n92 0.675548
R12726 VPWR.n207 VPWR.n95 0.675548
R12727 VPWR.n219 VPWR.n98 0.675548
R12728 VPWR.n231 VPWR.n101 0.675548
R12729 VPWR.n243 VPWR.n104 0.675548
R12730 VPWR.n255 VPWR.n107 0.675548
R12731 VPWR.n267 VPWR.n110 0.675548
R12732 VPWR.n279 VPWR.n113 0.675548
R12733 VPWR.n291 VPWR.n116 0.675548
R12734 VPWR.n308 VPWR.n307 0.675548
R12735 VPWR.n147 VPWR.n80 0.675548
R12736 VPWR.n136 VPWR.n77 0.675548
R12737 VPWR.n1754 VPWR.n1753 0.675548
R12738 VPWR.n1738 VPWR.n1076 0.675548
R12739 VPWR.n1726 VPWR.n1724 0.675548
R12740 VPWR.n1715 VPWR.n1713 0.675548
R12741 VPWR.n1215 VPWR.n1214 0.675548
R12742 VPWR.n1699 VPWR.n1697 0.675548
R12743 VPWR.n1688 VPWR.n1686 0.675548
R12744 VPWR.n1229 VPWR.n1228 0.675548
R12745 VPWR.n1672 VPWR.n1670 0.675548
R12746 VPWR.n1661 VPWR.n1659 0.675548
R12747 VPWR.n1197 VPWR.n1196 0.675548
R12748 VPWR.n1645 VPWR.n1643 0.675548
R12749 VPWR.n1634 VPWR.n1632 0.675548
R12750 VPWR.n1146 VPWR.n1145 0.675548
R12751 VPWR.n1618 VPWR.n1616 0.675548
R12752 VPWR.n2825 VPWR.n2824 0.672385
R12753 VPWR.n2809 VPWR.n2804 0.672385
R12754 VPWR.n2789 VPWR.n2784 0.672385
R12755 VPWR.n2770 VPWR.n2765 0.672385
R12756 VPWR.n2846 VPWR.n36 0.654518
R12757 VPWR.n7 VPWR 0.63497
R12758 VPWR.n1261 VPWR 0.63497
R12759 VPWR.n1284 VPWR 0.63497
R12760 VPWR.n1308 VPWR 0.63497
R12761 VPWR.n2852 VPWR.n26 0.573634
R12762 VPWR.n2848 VPWR.n2847 0.573634
R12763 VPWR VPWR.n2861 0.541783
R12764 VPWR.n43 VPWR 0.499542
R12765 VPWR.n2860 VPWR.n21 0.498268
R12766 VPWR.n2858 VPWR.n2857 0.493804
R12767 VPWR.n1139 VPWR.n1137 0.404056
R12768 VPWR.n163 VPWR.n157 0.404056
R12769 VPWR.n175 VPWR.n169 0.404056
R12770 VPWR.n187 VPWR.n181 0.404056
R12771 VPWR.n199 VPWR.n193 0.404056
R12772 VPWR.n211 VPWR.n205 0.404056
R12773 VPWR.n223 VPWR.n217 0.404056
R12774 VPWR.n235 VPWR.n229 0.404056
R12775 VPWR.n247 VPWR.n241 0.404056
R12776 VPWR.n259 VPWR.n253 0.404056
R12777 VPWR.n271 VPWR.n265 0.404056
R12778 VPWR.n283 VPWR.n277 0.404056
R12779 VPWR.n295 VPWR.n289 0.404056
R12780 VPWR.n302 VPWR.n120 0.404056
R12781 VPWR.n129 VPWR.n124 0.404056
R12782 VPWR.n151 VPWR.n145 0.404056
R12783 VPWR.n140 VPWR.n134 0.404056
R12784 VPWR.n1748 VPWR.n1084 0.404056
R12785 VPWR.n1742 VPWR.n1736 0.404056
R12786 VPWR.n1730 VPWR.n1089 0.404056
R12787 VPWR.n1723 VPWR.n1721 0.404056
R12788 VPWR.n1712 VPWR.n1710 0.404056
R12789 VPWR.n1703 VPWR.n1100 0.404056
R12790 VPWR.n1696 VPWR.n1694 0.404056
R12791 VPWR.n1685 VPWR.n1683 0.404056
R12792 VPWR.n1676 VPWR.n1110 0.404056
R12793 VPWR.n1669 VPWR.n1667 0.404056
R12794 VPWR.n1658 VPWR.n1656 0.404056
R12795 VPWR.n1649 VPWR.n1120 0.404056
R12796 VPWR.n1642 VPWR.n1640 0.404056
R12797 VPWR.n1631 VPWR.n1629 0.404056
R12798 VPWR.n1622 VPWR.n1130 0.404056
R12799 VPWR.n1627 VPWR.n1626 0.349144
R12800 VPWR.n1627 VPWR.n1118 0.349144
R12801 VPWR.n1653 VPWR.n1118 0.349144
R12802 VPWR.n1654 VPWR.n1653 0.349144
R12803 VPWR.n1654 VPWR.n1108 0.349144
R12804 VPWR.n1680 VPWR.n1108 0.349144
R12805 VPWR.n1681 VPWR.n1680 0.349144
R12806 VPWR.n1681 VPWR.n1098 0.349144
R12807 VPWR.n1707 VPWR.n1098 0.349144
R12808 VPWR.n1708 VPWR.n1707 0.349144
R12809 VPWR.n1708 VPWR.n1087 0.349144
R12810 VPWR.n1734 VPWR.n1087 0.349144
R12811 VPWR.n1746 VPWR.n1734 0.349144
R12812 VPWR.n300 VPWR.n299 0.349144
R12813 VPWR.n299 VPWR.n287 0.349144
R12814 VPWR.n287 VPWR.n275 0.349144
R12815 VPWR.n275 VPWR.n263 0.349144
R12816 VPWR.n263 VPWR.n251 0.349144
R12817 VPWR.n251 VPWR.n239 0.349144
R12818 VPWR.n239 VPWR.n227 0.349144
R12819 VPWR.n227 VPWR.n215 0.349144
R12820 VPWR.n215 VPWR.n203 0.349144
R12821 VPWR.n203 VPWR.n191 0.349144
R12822 VPWR.n191 VPWR.n179 0.349144
R12823 VPWR.n179 VPWR.n167 0.349144
R12824 VPWR.n167 VPWR.n155 0.349144
R12825 VPWR.n1481 VPWR.n1475 0.346131
R12826 VPWR.n1480 VPWR.n1476 0.346131
R12827 VPWR.n1601 VPWR.n1155 0.346131
R12828 VPWR.n1600 VPWR.n1596 0.346131
R12829 VPWR.n1595 VPWR.n1591 0.346131
R12830 VPWR.n1590 VPWR.n1586 0.346131
R12831 VPWR.n1585 VPWR.n1581 0.346131
R12832 VPWR.n1580 VPWR.n1576 0.346131
R12833 VPWR.n1575 VPWR.n1571 0.346131
R12834 VPWR.n1570 VPWR.n1566 0.346131
R12835 VPWR.n1565 VPWR.n1561 0.346131
R12836 VPWR.n1786 VPWR.n1061 0.346131
R12837 VPWR.n1803 VPWR.n1799 0.346131
R12838 VPWR.n1804 VPWR.n1795 0.346131
R12839 VPWR.n1791 VPWR.n1790 0.346131
R12840 VPWR.n2613 VPWR.n74 0.300179
R12841 VPWR.n2833 VPWR.n38 0.298167
R12842 VPWR.n1137 VPWR.n1132 0.286958
R12843 VPWR.n164 VPWR.n163 0.286958
R12844 VPWR.n176 VPWR.n175 0.286958
R12845 VPWR.n188 VPWR.n187 0.286958
R12846 VPWR.n200 VPWR.n199 0.286958
R12847 VPWR.n212 VPWR.n211 0.286958
R12848 VPWR.n224 VPWR.n223 0.286958
R12849 VPWR.n236 VPWR.n235 0.286958
R12850 VPWR.n248 VPWR.n247 0.286958
R12851 VPWR.n260 VPWR.n259 0.286958
R12852 VPWR.n272 VPWR.n271 0.286958
R12853 VPWR.n284 VPWR.n283 0.286958
R12854 VPWR.n296 VPWR.n295 0.286958
R12855 VPWR.n302 VPWR.n121 0.286958
R12856 VPWR.n130 VPWR.n129 0.286958
R12857 VPWR.n152 VPWR.n151 0.286958
R12858 VPWR.n141 VPWR.n140 0.286958
R12859 VPWR.n1748 VPWR.n1085 0.286958
R12860 VPWR.n1743 VPWR.n1742 0.286958
R12861 VPWR.n1731 VPWR.n1730 0.286958
R12862 VPWR.n1721 VPWR.n1091 0.286958
R12863 VPWR.n1710 VPWR.n1094 0.286958
R12864 VPWR.n1704 VPWR.n1703 0.286958
R12865 VPWR.n1694 VPWR.n1102 0.286958
R12866 VPWR.n1683 VPWR.n1104 0.286958
R12867 VPWR.n1677 VPWR.n1676 0.286958
R12868 VPWR.n1667 VPWR.n1112 0.286958
R12869 VPWR.n1656 VPWR.n1114 0.286958
R12870 VPWR.n1650 VPWR.n1649 0.286958
R12871 VPWR.n1640 VPWR.n1122 0.286958
R12872 VPWR.n1629 VPWR.n1124 0.286958
R12873 VPWR.n1623 VPWR.n1622 0.286958
R12874 VPWR.n74 VPWR 0.2505
R12875 VPWR VPWR.n2500 0.249238
R12876 VPWR.n2491 VPWR 0.249238
R12877 VPWR VPWR.n2490 0.249238
R12878 VPWR.n2404 VPWR 0.249238
R12879 VPWR.n2405 VPWR 0.249238
R12880 VPWR.n2406 VPWR 0.249238
R12881 VPWR.n2407 VPWR 0.249238
R12882 VPWR.n2324 VPWR 0.249238
R12883 VPWR.n2333 VPWR 0.249238
R12884 VPWR.n2334 VPWR 0.249238
R12885 VPWR.n2343 VPWR 0.249238
R12886 VPWR.n2344 VPWR 0.249238
R12887 VPWR.n2402 VPWR 0.249238
R12888 VPWR.n2394 VPWR 0.249238
R12889 VPWR.n2393 VPWR 0.249238
R12890 VPWR.n2384 VPWR 0.249238
R12891 VPWR.n2383 VPWR 0.249238
R12892 VPWR.n2374 VPWR 0.249238
R12893 VPWR.n2373 VPWR 0.249238
R12894 VPWR.n2364 VPWR 0.249238
R12895 VPWR.n2363 VPWR 0.249238
R12896 VPWR.n2354 VPWR 0.249238
R12897 VPWR.n2353 VPWR 0.249238
R12898 VPWR VPWR.n2321 0.249238
R12899 VPWR VPWR.n2320 0.249238
R12900 VPWR VPWR.n2319 0.249238
R12901 VPWR VPWR.n2318 0.249238
R12902 VPWR VPWR.n2317 0.249238
R12903 VPWR VPWR.n2306 0.249238
R12904 VPWR VPWR.n2307 0.249238
R12905 VPWR VPWR.n2308 0.249238
R12906 VPWR VPWR.n2309 0.249238
R12907 VPWR VPWR.n2310 0.249238
R12908 VPWR VPWR.n2311 0.249238
R12909 VPWR VPWR.n2312 0.249238
R12910 VPWR VPWR.n2313 0.249238
R12911 VPWR VPWR.n2314 0.249238
R12912 VPWR VPWR.n2315 0.249238
R12913 VPWR VPWR.n2316 0.249238
R12914 VPWR VPWR.n2304 0.249238
R12915 VPWR.n2295 VPWR 0.249238
R12916 VPWR VPWR.n2294 0.249238
R12917 VPWR.n2285 VPWR 0.249238
R12918 VPWR VPWR.n2284 0.249238
R12919 VPWR.n2226 VPWR 0.249238
R12920 VPWR VPWR.n2234 0.249238
R12921 VPWR.n2235 VPWR 0.249238
R12922 VPWR VPWR.n2244 0.249238
R12923 VPWR.n2245 VPWR 0.249238
R12924 VPWR VPWR.n2254 0.249238
R12925 VPWR.n2255 VPWR 0.249238
R12926 VPWR VPWR.n2264 0.249238
R12927 VPWR.n2265 VPWR 0.249238
R12928 VPWR VPWR.n2274 0.249238
R12929 VPWR.n2275 VPWR 0.249238
R12930 VPWR.n2208 VPWR 0.249238
R12931 VPWR.n2209 VPWR 0.249238
R12932 VPWR.n2210 VPWR 0.249238
R12933 VPWR.n2211 VPWR 0.249238
R12934 VPWR.n2212 VPWR 0.249238
R12935 VPWR.n2223 VPWR 0.249238
R12936 VPWR.n2222 VPWR 0.249238
R12937 VPWR.n2221 VPWR 0.249238
R12938 VPWR.n2220 VPWR 0.249238
R12939 VPWR.n2219 VPWR 0.249238
R12940 VPWR.n2218 VPWR 0.249238
R12941 VPWR.n2217 VPWR 0.249238
R12942 VPWR.n2216 VPWR 0.249238
R12943 VPWR.n2215 VPWR 0.249238
R12944 VPWR.n2214 VPWR 0.249238
R12945 VPWR.n2213 VPWR 0.249238
R12946 VPWR.n2128 VPWR 0.249238
R12947 VPWR.n2137 VPWR 0.249238
R12948 VPWR.n2138 VPWR 0.249238
R12949 VPWR.n2147 VPWR 0.249238
R12950 VPWR.n2148 VPWR 0.249238
R12951 VPWR.n2206 VPWR 0.249238
R12952 VPWR.n2198 VPWR 0.249238
R12953 VPWR.n2197 VPWR 0.249238
R12954 VPWR.n2188 VPWR 0.249238
R12955 VPWR.n2187 VPWR 0.249238
R12956 VPWR.n2178 VPWR 0.249238
R12957 VPWR.n2177 VPWR 0.249238
R12958 VPWR.n2168 VPWR 0.249238
R12959 VPWR.n2167 VPWR 0.249238
R12960 VPWR.n2158 VPWR 0.249238
R12961 VPWR.n2157 VPWR 0.249238
R12962 VPWR VPWR.n2125 0.249238
R12963 VPWR VPWR.n2124 0.249238
R12964 VPWR VPWR.n2123 0.249238
R12965 VPWR VPWR.n2122 0.249238
R12966 VPWR VPWR.n2121 0.249238
R12967 VPWR VPWR.n2110 0.249238
R12968 VPWR VPWR.n2111 0.249238
R12969 VPWR VPWR.n2112 0.249238
R12970 VPWR VPWR.n2113 0.249238
R12971 VPWR VPWR.n2114 0.249238
R12972 VPWR VPWR.n2115 0.249238
R12973 VPWR VPWR.n2116 0.249238
R12974 VPWR VPWR.n2117 0.249238
R12975 VPWR VPWR.n2118 0.249238
R12976 VPWR VPWR.n2119 0.249238
R12977 VPWR VPWR.n2120 0.249238
R12978 VPWR VPWR.n2108 0.249238
R12979 VPWR.n2099 VPWR 0.249238
R12980 VPWR VPWR.n2098 0.249238
R12981 VPWR.n2089 VPWR 0.249238
R12982 VPWR VPWR.n2088 0.249238
R12983 VPWR.n2030 VPWR 0.249238
R12984 VPWR VPWR.n2038 0.249238
R12985 VPWR.n2039 VPWR 0.249238
R12986 VPWR VPWR.n2048 0.249238
R12987 VPWR.n2049 VPWR 0.249238
R12988 VPWR VPWR.n2058 0.249238
R12989 VPWR.n2059 VPWR 0.249238
R12990 VPWR VPWR.n2068 0.249238
R12991 VPWR.n2069 VPWR 0.249238
R12992 VPWR VPWR.n2078 0.249238
R12993 VPWR.n2079 VPWR 0.249238
R12994 VPWR.n2012 VPWR 0.249238
R12995 VPWR.n2013 VPWR 0.249238
R12996 VPWR.n2014 VPWR 0.249238
R12997 VPWR.n2015 VPWR 0.249238
R12998 VPWR.n2016 VPWR 0.249238
R12999 VPWR.n2027 VPWR 0.249238
R13000 VPWR.n2026 VPWR 0.249238
R13001 VPWR.n2025 VPWR 0.249238
R13002 VPWR.n2024 VPWR 0.249238
R13003 VPWR.n2023 VPWR 0.249238
R13004 VPWR.n2022 VPWR 0.249238
R13005 VPWR.n2021 VPWR 0.249238
R13006 VPWR.n2020 VPWR 0.249238
R13007 VPWR.n2019 VPWR 0.249238
R13008 VPWR.n2018 VPWR 0.249238
R13009 VPWR.n2017 VPWR 0.249238
R13010 VPWR.n1932 VPWR 0.249238
R13011 VPWR.n1941 VPWR 0.249238
R13012 VPWR.n1942 VPWR 0.249238
R13013 VPWR.n1951 VPWR 0.249238
R13014 VPWR.n1952 VPWR 0.249238
R13015 VPWR.n2010 VPWR 0.249238
R13016 VPWR.n2002 VPWR 0.249238
R13017 VPWR.n2001 VPWR 0.249238
R13018 VPWR.n1992 VPWR 0.249238
R13019 VPWR.n1991 VPWR 0.249238
R13020 VPWR.n1982 VPWR 0.249238
R13021 VPWR.n1981 VPWR 0.249238
R13022 VPWR.n1972 VPWR 0.249238
R13023 VPWR.n1971 VPWR 0.249238
R13024 VPWR.n1962 VPWR 0.249238
R13025 VPWR.n1961 VPWR 0.249238
R13026 VPWR VPWR.n1929 0.249238
R13027 VPWR VPWR.n1928 0.249238
R13028 VPWR VPWR.n1927 0.249238
R13029 VPWR VPWR.n1926 0.249238
R13030 VPWR VPWR.n1925 0.249238
R13031 VPWR VPWR.n1914 0.249238
R13032 VPWR VPWR.n1915 0.249238
R13033 VPWR VPWR.n1916 0.249238
R13034 VPWR VPWR.n1917 0.249238
R13035 VPWR VPWR.n1918 0.249238
R13036 VPWR VPWR.n1919 0.249238
R13037 VPWR VPWR.n1920 0.249238
R13038 VPWR VPWR.n1921 0.249238
R13039 VPWR VPWR.n1922 0.249238
R13040 VPWR VPWR.n1923 0.249238
R13041 VPWR VPWR.n1924 0.249238
R13042 VPWR.n2419 VPWR 0.249238
R13043 VPWR.n2418 VPWR 0.249238
R13044 VPWR.n2417 VPWR 0.249238
R13045 VPWR.n2416 VPWR 0.249238
R13046 VPWR.n2415 VPWR 0.249238
R13047 VPWR.n2414 VPWR 0.249238
R13048 VPWR.n2413 VPWR 0.249238
R13049 VPWR.n2412 VPWR 0.249238
R13050 VPWR.n2411 VPWR 0.249238
R13051 VPWR.n2410 VPWR 0.249238
R13052 VPWR.n2409 VPWR 0.249238
R13053 VPWR.n2408 VPWR 0.249238
R13054 VPWR VPWR.n1912 0.249238
R13055 VPWR.n1903 VPWR 0.249238
R13056 VPWR VPWR.n1902 0.249238
R13057 VPWR.n1893 VPWR 0.249238
R13058 VPWR VPWR.n1892 0.249238
R13059 VPWR.n1883 VPWR 0.249238
R13060 VPWR.n1834 VPWR 0.249238
R13061 VPWR VPWR.n1842 0.249238
R13062 VPWR.n1843 VPWR 0.249238
R13063 VPWR VPWR.n1852 0.249238
R13064 VPWR.n1853 VPWR 0.249238
R13065 VPWR VPWR.n1862 0.249238
R13066 VPWR.n1863 VPWR 0.249238
R13067 VPWR VPWR.n1872 0.249238
R13068 VPWR.n1873 VPWR 0.249238
R13069 VPWR VPWR.n1882 0.249238
R13070 VPWR.n2422 VPWR 0.249238
R13071 VPWR VPWR.n2430 0.249238
R13072 VPWR.n2431 VPWR 0.249238
R13073 VPWR VPWR.n2440 0.249238
R13074 VPWR.n2441 VPWR 0.249238
R13075 VPWR VPWR.n2450 0.249238
R13076 VPWR.n2451 VPWR 0.249238
R13077 VPWR VPWR.n2460 0.249238
R13078 VPWR.n2461 VPWR 0.249238
R13079 VPWR VPWR.n2470 0.249238
R13080 VPWR.n2471 VPWR 0.249238
R13081 VPWR VPWR.n2480 0.249238
R13082 VPWR.n2481 VPWR 0.249238
R13083 VPWR.n1816 VPWR 0.249238
R13084 VPWR.n1817 VPWR 0.249238
R13085 VPWR.n1818 VPWR 0.249238
R13086 VPWR.n1819 VPWR 0.249238
R13087 VPWR.n1820 VPWR 0.249238
R13088 VPWR.n1821 VPWR 0.249238
R13089 VPWR.n1822 VPWR 0.249238
R13090 VPWR.n1823 VPWR 0.249238
R13091 VPWR.n1824 VPWR 0.249238
R13092 VPWR.n1831 VPWR 0.249238
R13093 VPWR.n1830 VPWR 0.249238
R13094 VPWR.n1829 VPWR 0.249238
R13095 VPWR.n1828 VPWR 0.249238
R13096 VPWR.n1827 VPWR 0.249238
R13097 VPWR.n1826 VPWR 0.249238
R13098 VPWR.n1825 VPWR 0.249238
R13099 VPWR VPWR.n2517 0.249238
R13100 VPWR VPWR.n2516 0.249238
R13101 VPWR VPWR.n2515 0.249238
R13102 VPWR VPWR.n2514 0.249238
R13103 VPWR VPWR.n2513 0.249238
R13104 VPWR VPWR.n2512 0.249238
R13105 VPWR VPWR.n2511 0.249238
R13106 VPWR VPWR.n2510 0.249238
R13107 VPWR VPWR.n2509 0.249238
R13108 VPWR VPWR.n2508 0.249238
R13109 VPWR VPWR.n2507 0.249238
R13110 VPWR VPWR.n2502 0.249238
R13111 VPWR VPWR.n2503 0.249238
R13112 VPWR VPWR.n2504 0.249238
R13113 VPWR VPWR.n2505 0.249238
R13114 VPWR VPWR.n2506 0.249238
R13115 VPWR.n2520 VPWR 0.249238
R13116 VPWR.n2531 VPWR 0.249238
R13117 VPWR.n2532 VPWR 0.249238
R13118 VPWR.n2543 VPWR 0.249238
R13119 VPWR.n2544 VPWR 0.249238
R13120 VPWR.n2555 VPWR 0.249238
R13121 VPWR.n2556 VPWR 0.249238
R13122 VPWR.n2567 VPWR 0.249238
R13123 VPWR.n2568 VPWR 0.249238
R13124 VPWR.n2579 VPWR 0.249238
R13125 VPWR.n2580 VPWR 0.249238
R13126 VPWR.n2591 VPWR 0.249238
R13127 VPWR.n2592 VPWR 0.249238
R13128 VPWR.n2603 VPWR 0.249238
R13129 VPWR.n2604 VPWR 0.249238
R13130 VPWR.n2614 VPWR 0.249238
R13131 VPWR VPWR.n1074 0.249238
R13132 VPWR VPWR.n1075 0.249238
R13133 VPWR VPWR.n1773 0.249238
R13134 VPWR.n1774 VPWR 0.249238
R13135 VPWR VPWR.n1548 0.249238
R13136 VPWR.n1549 VPWR 0.249238
R13137 VPWR.n1547 VPWR 0.249238
R13138 VPWR.n1546 VPWR 0.249238
R13139 VPWR.n1533 VPWR 0.249238
R13140 VPWR.n1532 VPWR 0.249238
R13141 VPWR.n1519 VPWR 0.249238
R13142 VPWR.n1518 VPWR 0.249238
R13143 VPWR.n1506 VPWR 0.249238
R13144 VPWR VPWR.n1606 0.249238
R13145 VPWR.n1607 VPWR 0.249238
R13146 VPWR VPWR.n1467 0.249238
R13147 VPWR.n36 VPWR.n22 0.242688
R13148 VPWR.n2832 VPWR.n2816 0.213567
R13149 VPWR.n2816 VPWR.n2797 0.213567
R13150 VPWR.n2797 VPWR.n2777 0.213567
R13151 VPWR.n2777 VPWR.n2758 0.213567
R13152 VPWR.n2758 VPWR.n2722 0.213567
R13153 VPWR.n2722 VPWR.n2684 0.213567
R13154 VPWR.n2684 VPWR.n2647 0.213567
R13155 VPWR.n1465 VPWR.n1433 0.213567
R13156 VPWR.n1433 VPWR.n1395 0.213567
R13157 VPWR.n1395 VPWR.n1356 0.213567
R13158 VPWR.n1356 VPWR.n1321 0.213567
R13159 VPWR.n1321 VPWR.n1298 0.213567
R13160 VPWR.n1298 VPWR.n1274 0.213567
R13161 VPWR.n1274 VPWR.n19 0.213567
R13162 VPWR.n2846 VPWR.n2845 0.189116
R13163 VPWR.n2861 VPWR.n20 0.182233
R13164 VPWR.n1468 VPWR.n1466 0.179202
R13165 VPWR.n1469 VPWR.n1468 0.154425
R13166 VPWR.n1469 VPWR.n949 0.154425
R13167 VPWR.n1913 VPWR.n949 0.154425
R13168 VPWR.n1930 VPWR.n1913 0.154425
R13169 VPWR.n1931 VPWR.n1930 0.154425
R13170 VPWR.n1931 VPWR.n757 0.154425
R13171 VPWR.n2109 VPWR.n757 0.154425
R13172 VPWR.n2126 VPWR.n2109 0.154425
R13173 VPWR.n2127 VPWR.n2126 0.154425
R13174 VPWR.n2127 VPWR.n565 0.154425
R13175 VPWR.n2305 VPWR.n565 0.154425
R13176 VPWR.n2322 VPWR.n2305 0.154425
R13177 VPWR.n2323 VPWR.n2322 0.154425
R13178 VPWR.n2323 VPWR.n373 0.154425
R13179 VPWR.n2501 VPWR.n373 0.154425
R13180 VPWR.n2518 VPWR.n2501 0.154425
R13181 VPWR.n2519 VPWR.n2518 0.154425
R13182 VPWR.n1815 VPWR.n1045 0.154425
R13183 VPWR.n1832 VPWR.n1815 0.154425
R13184 VPWR.n1833 VPWR.n1832 0.154425
R13185 VPWR.n1833 VPWR.n853 0.154425
R13186 VPWR.n2011 VPWR.n853 0.154425
R13187 VPWR.n2028 VPWR.n2011 0.154425
R13188 VPWR.n2029 VPWR.n2028 0.154425
R13189 VPWR.n2029 VPWR.n661 0.154425
R13190 VPWR.n2207 VPWR.n661 0.154425
R13191 VPWR.n2224 VPWR.n2207 0.154425
R13192 VPWR.n2225 VPWR.n2224 0.154425
R13193 VPWR.n2225 VPWR.n469 0.154425
R13194 VPWR.n2403 VPWR.n469 0.154425
R13195 VPWR.n2420 VPWR.n2403 0.154425
R13196 VPWR.n2421 VPWR.n2420 0.154425
R13197 VPWR.n2421 VPWR.n40 0.154425
R13198 VPWR.n2615 VPWR.n40 0.154425
R13199 VPWR.n8 VPWR.n7 0.147771
R13200 VPWR.n1262 VPWR.n1261 0.147771
R13201 VPWR.n1285 VPWR.n1284 0.147771
R13202 VPWR.n1309 VPWR.n1308 0.147771
R13203 VPWR.n2833 VPWR.n2832 0.145025
R13204 VPWR.n1132 VPWR 0.135917
R13205 VPWR.n164 VPWR 0.135917
R13206 VPWR.n176 VPWR 0.135917
R13207 VPWR.n188 VPWR 0.135917
R13208 VPWR.n200 VPWR 0.135917
R13209 VPWR.n212 VPWR 0.135917
R13210 VPWR.n224 VPWR 0.135917
R13211 VPWR.n236 VPWR 0.135917
R13212 VPWR.n248 VPWR 0.135917
R13213 VPWR.n260 VPWR 0.135917
R13214 VPWR.n272 VPWR 0.135917
R13215 VPWR.n284 VPWR 0.135917
R13216 VPWR.n296 VPWR 0.135917
R13217 VPWR.n121 VPWR 0.135917
R13218 VPWR.n130 VPWR 0.135917
R13219 VPWR.n152 VPWR 0.135917
R13220 VPWR.n141 VPWR 0.135917
R13221 VPWR.n1085 VPWR 0.135917
R13222 VPWR.n1743 VPWR 0.135917
R13223 VPWR.n1731 VPWR 0.135917
R13224 VPWR.n1091 VPWR 0.135917
R13225 VPWR.n1094 VPWR 0.135917
R13226 VPWR.n1704 VPWR 0.135917
R13227 VPWR.n1102 VPWR 0.135917
R13228 VPWR.n1104 VPWR 0.135917
R13229 VPWR.n1677 VPWR 0.135917
R13230 VPWR.n1112 VPWR 0.135917
R13231 VPWR.n1114 VPWR 0.135917
R13232 VPWR.n1650 VPWR 0.135917
R13233 VPWR.n1122 VPWR 0.135917
R13234 VPWR.n1124 VPWR 0.135917
R13235 VPWR.n1623 VPWR 0.135917
R13236 VPWR.n38 VPWR.n37 0.123287
R13237 VPWR.n18 VPWR.n0 0.120292
R13238 VPWR.n14 VPWR.n0 0.120292
R13239 VPWR.n9 VPWR.n8 0.120292
R13240 VPWR.n1273 VPWR.n1252 0.120292
R13241 VPWR.n1269 VPWR.n1252 0.120292
R13242 VPWR.n1263 VPWR.n1262 0.120292
R13243 VPWR.n1297 VPWR.n1275 0.120292
R13244 VPWR.n1292 VPWR.n1275 0.120292
R13245 VPWR.n1286 VPWR.n1285 0.120292
R13246 VPWR.n1320 VPWR.n1299 0.120292
R13247 VPWR.n1316 VPWR.n1299 0.120292
R13248 VPWR.n1310 VPWR.n1309 0.120292
R13249 VPWR.n1352 VPWR.n1351 0.120292
R13250 VPWR.n1345 VPWR.n1324 0.120292
R13251 VPWR.n1338 VPWR.n1324 0.120292
R13252 VPWR.n1338 VPWR.n1337 0.120292
R13253 VPWR.n1336 VPWR.n1328 0.120292
R13254 VPWR.n1331 VPWR.n1328 0.120292
R13255 VPWR.n1331 VPWR.n1330 0.120292
R13256 VPWR.n1390 VPWR.n1389 0.120292
R13257 VPWR.n1383 VPWR.n1382 0.120292
R13258 VPWR.n1382 VPWR.n1359 0.120292
R13259 VPWR.n1375 VPWR.n1359 0.120292
R13260 VPWR.n1375 VPWR.n1374 0.120292
R13261 VPWR.n1374 VPWR.n1373 0.120292
R13262 VPWR.n1373 VPWR.n1361 0.120292
R13263 VPWR.n1367 VPWR.n1361 0.120292
R13264 VPWR.n1367 VPWR.n1366 0.120292
R13265 VPWR.n1429 VPWR.n1428 0.120292
R13266 VPWR.n1422 VPWR.n1421 0.120292
R13267 VPWR.n1421 VPWR.n1398 0.120292
R13268 VPWR.n1414 VPWR.n1398 0.120292
R13269 VPWR.n1414 VPWR.n1413 0.120292
R13270 VPWR.n1413 VPWR.n1412 0.120292
R13271 VPWR.n1412 VPWR.n1400 0.120292
R13272 VPWR.n1406 VPWR.n1400 0.120292
R13273 VPWR.n1406 VPWR.n1405 0.120292
R13274 VPWR.n1459 VPWR.n1458 0.120292
R13275 VPWR.n1458 VPWR.n1435 0.120292
R13276 VPWR.n1451 VPWR.n1435 0.120292
R13277 VPWR.n1451 VPWR.n1450 0.120292
R13278 VPWR.n1450 VPWR.n1449 0.120292
R13279 VPWR.n1449 VPWR.n1437 0.120292
R13280 VPWR.n1443 VPWR.n1437 0.120292
R13281 VPWR.n1443 VPWR.n1442 0.120292
R13282 VPWR.n2831 VPWR.n2817 0.120292
R13283 VPWR.n2815 VPWR.n2798 0.120292
R13284 VPWR.n2796 VPWR.n2778 0.120292
R13285 VPWR.n2776 VPWR.n2759 0.120292
R13286 VPWR.n2738 VPWR.n2737 0.120292
R13287 VPWR.n2739 VPWR.n2738 0.120292
R13288 VPWR.n2739 VPWR.n2730 0.120292
R13289 VPWR.n2744 VPWR.n2730 0.120292
R13290 VPWR.n2745 VPWR.n2744 0.120292
R13291 VPWR.n2745 VPWR.n2726 0.120292
R13292 VPWR.n2751 VPWR.n2726 0.120292
R13293 VPWR.n2753 VPWR.n2723 0.120292
R13294 VPWR.n2757 VPWR.n2723 0.120292
R13295 VPWR.n2702 VPWR.n2701 0.120292
R13296 VPWR.n2703 VPWR.n2702 0.120292
R13297 VPWR.n2703 VPWR.n2692 0.120292
R13298 VPWR.n2708 VPWR.n2692 0.120292
R13299 VPWR.n2709 VPWR.n2708 0.120292
R13300 VPWR.n2709 VPWR.n2688 0.120292
R13301 VPWR.n2714 VPWR.n2688 0.120292
R13302 VPWR.n2716 VPWR.n2685 0.120292
R13303 VPWR.n2721 VPWR.n2685 0.120292
R13304 VPWR.n2665 VPWR.n2664 0.120292
R13305 VPWR.n2666 VPWR.n2665 0.120292
R13306 VPWR.n2666 VPWR.n2655 0.120292
R13307 VPWR.n2671 VPWR.n2655 0.120292
R13308 VPWR.n2672 VPWR.n2671 0.120292
R13309 VPWR.n2672 VPWR.n2651 0.120292
R13310 VPWR.n2677 VPWR.n2651 0.120292
R13311 VPWR.n2679 VPWR.n2648 0.120292
R13312 VPWR.n2683 VPWR.n2648 0.120292
R13313 VPWR.n2627 VPWR.n2623 0.120292
R13314 VPWR.n2635 VPWR.n2623 0.120292
R13315 VPWR.n2636 VPWR.n2635 0.120292
R13316 VPWR.n2637 VPWR.n2636 0.120292
R13317 VPWR.n2637 VPWR.n2619 0.120292
R13318 VPWR.n2642 VPWR.n2619 0.120292
R13319 VPWR.n2643 VPWR.n2642 0.120292
R13320 VPWR.n1624 VPWR 0.118556
R13321 VPWR.n1127 VPWR 0.118556
R13322 VPWR.n1638 VPWR 0.118556
R13323 VPWR.n1651 VPWR 0.118556
R13324 VPWR.n1117 VPWR 0.118556
R13325 VPWR.n1665 VPWR 0.118556
R13326 VPWR.n1678 VPWR 0.118556
R13327 VPWR.n1107 VPWR 0.118556
R13328 VPWR.n1692 VPWR 0.118556
R13329 VPWR.n1705 VPWR 0.118556
R13330 VPWR.n1097 VPWR 0.118556
R13331 VPWR.n1719 VPWR 0.118556
R13332 VPWR.n1732 VPWR 0.118556
R13333 VPWR.n1744 VPWR 0.118556
R13334 VPWR VPWR.n1131 0.118556
R13335 VPWR.n1086 VPWR 0.118556
R13336 VPWR.n142 VPWR 0.118556
R13337 VPWR.n131 VPWR 0.118556
R13338 VPWR.n122 VPWR 0.118556
R13339 VPWR.n297 VPWR 0.118556
R13340 VPWR.n285 VPWR 0.118556
R13341 VPWR.n273 VPWR 0.118556
R13342 VPWR.n261 VPWR 0.118556
R13343 VPWR.n249 VPWR 0.118556
R13344 VPWR.n237 VPWR 0.118556
R13345 VPWR.n225 VPWR 0.118556
R13346 VPWR.n213 VPWR 0.118556
R13347 VPWR.n201 VPWR 0.118556
R13348 VPWR.n189 VPWR 0.118556
R13349 VPWR.n177 VPWR 0.118556
R13350 VPWR.n165 VPWR 0.118556
R13351 VPWR.n153 VPWR 0.118556
R13352 VPWR.n1784 VPWR.n1063 0.108238
R13353 VPWR.n1560 VPWR.n1162 0.108238
R13354 VPWR.n1559 VPWR.n1161 0.108238
R13355 VPWR.n1543 VPWR.n1160 0.108238
R13356 VPWR.n1535 VPWR.n1159 0.108238
R13357 VPWR.n1529 VPWR.n1158 0.108238
R13358 VPWR.n1521 VPWR.n1157 0.108238
R13359 VPWR.n1515 VPWR.n1156 0.108238
R13360 VPWR.n1602 VPWR.n1151 0.108238
R13361 VPWR.n1603 VPWR.n1150 0.108238
R13362 VPWR.n1482 VPWR.n1471 0.108238
R13363 VPWR.n1483 VPWR.n1470 0.108238
R13364 VPWR.n1814 VPWR.n1046 0.108238
R13365 VPWR.n1785 VPWR.n1062 0.108238
R13366 VPWR.n1763 VPWR.n1057 0.108238
R13367 VPWR.n1806 VPWR.n1805 0.108238
R13368 VPWR.n2500 VPWR 0.100405
R13369 VPWR.n2491 VPWR 0.100405
R13370 VPWR VPWR.n2404 0.100405
R13371 VPWR VPWR.n2405 0.100405
R13372 VPWR VPWR.n2406 0.100405
R13373 VPWR.n2324 VPWR 0.100405
R13374 VPWR VPWR.n2333 0.100405
R13375 VPWR.n2334 VPWR 0.100405
R13376 VPWR VPWR.n2343 0.100405
R13377 VPWR.n2394 VPWR 0.100405
R13378 VPWR VPWR.n2393 0.100405
R13379 VPWR.n2384 VPWR 0.100405
R13380 VPWR VPWR.n2383 0.100405
R13381 VPWR.n2374 VPWR 0.100405
R13382 VPWR VPWR.n2373 0.100405
R13383 VPWR.n2364 VPWR 0.100405
R13384 VPWR VPWR.n2363 0.100405
R13385 VPWR.n2354 VPWR 0.100405
R13386 VPWR VPWR.n2353 0.100405
R13387 VPWR.n2344 VPWR 0.100405
R13388 VPWR.n2321 VPWR 0.100405
R13389 VPWR.n2320 VPWR 0.100405
R13390 VPWR.n2319 VPWR 0.100405
R13391 VPWR.n2318 VPWR 0.100405
R13392 VPWR.n2307 VPWR 0.100405
R13393 VPWR.n2308 VPWR 0.100405
R13394 VPWR.n2309 VPWR 0.100405
R13395 VPWR.n2310 VPWR 0.100405
R13396 VPWR.n2311 VPWR 0.100405
R13397 VPWR.n2312 VPWR 0.100405
R13398 VPWR.n2313 VPWR 0.100405
R13399 VPWR.n2314 VPWR 0.100405
R13400 VPWR.n2315 VPWR 0.100405
R13401 VPWR.n2316 VPWR 0.100405
R13402 VPWR.n2317 VPWR 0.100405
R13403 VPWR.n2304 VPWR 0.100405
R13404 VPWR.n2295 VPWR 0.100405
R13405 VPWR.n2294 VPWR 0.100405
R13406 VPWR.n2285 VPWR 0.100405
R13407 VPWR.n2234 VPWR 0.100405
R13408 VPWR.n2235 VPWR 0.100405
R13409 VPWR.n2244 VPWR 0.100405
R13410 VPWR.n2245 VPWR 0.100405
R13411 VPWR.n2254 VPWR 0.100405
R13412 VPWR.n2255 VPWR 0.100405
R13413 VPWR.n2264 VPWR 0.100405
R13414 VPWR.n2265 VPWR 0.100405
R13415 VPWR.n2274 VPWR 0.100405
R13416 VPWR.n2275 VPWR 0.100405
R13417 VPWR.n2284 VPWR 0.100405
R13418 VPWR VPWR.n2208 0.100405
R13419 VPWR VPWR.n2209 0.100405
R13420 VPWR VPWR.n2210 0.100405
R13421 VPWR VPWR.n2211 0.100405
R13422 VPWR VPWR.n2222 0.100405
R13423 VPWR VPWR.n2221 0.100405
R13424 VPWR VPWR.n2220 0.100405
R13425 VPWR VPWR.n2219 0.100405
R13426 VPWR VPWR.n2218 0.100405
R13427 VPWR VPWR.n2217 0.100405
R13428 VPWR VPWR.n2216 0.100405
R13429 VPWR VPWR.n2215 0.100405
R13430 VPWR VPWR.n2214 0.100405
R13431 VPWR VPWR.n2213 0.100405
R13432 VPWR VPWR.n2212 0.100405
R13433 VPWR.n2128 VPWR 0.100405
R13434 VPWR VPWR.n2137 0.100405
R13435 VPWR.n2138 VPWR 0.100405
R13436 VPWR VPWR.n2147 0.100405
R13437 VPWR.n2198 VPWR 0.100405
R13438 VPWR VPWR.n2197 0.100405
R13439 VPWR.n2188 VPWR 0.100405
R13440 VPWR VPWR.n2187 0.100405
R13441 VPWR.n2178 VPWR 0.100405
R13442 VPWR VPWR.n2177 0.100405
R13443 VPWR.n2168 VPWR 0.100405
R13444 VPWR VPWR.n2167 0.100405
R13445 VPWR.n2158 VPWR 0.100405
R13446 VPWR VPWR.n2157 0.100405
R13447 VPWR.n2148 VPWR 0.100405
R13448 VPWR.n2125 VPWR 0.100405
R13449 VPWR.n2124 VPWR 0.100405
R13450 VPWR.n2123 VPWR 0.100405
R13451 VPWR.n2122 VPWR 0.100405
R13452 VPWR.n2111 VPWR 0.100405
R13453 VPWR.n2112 VPWR 0.100405
R13454 VPWR.n2113 VPWR 0.100405
R13455 VPWR.n2114 VPWR 0.100405
R13456 VPWR.n2115 VPWR 0.100405
R13457 VPWR.n2116 VPWR 0.100405
R13458 VPWR.n2117 VPWR 0.100405
R13459 VPWR.n2118 VPWR 0.100405
R13460 VPWR.n2119 VPWR 0.100405
R13461 VPWR.n2120 VPWR 0.100405
R13462 VPWR.n2121 VPWR 0.100405
R13463 VPWR.n2108 VPWR 0.100405
R13464 VPWR.n2099 VPWR 0.100405
R13465 VPWR.n2098 VPWR 0.100405
R13466 VPWR.n2089 VPWR 0.100405
R13467 VPWR.n2038 VPWR 0.100405
R13468 VPWR.n2039 VPWR 0.100405
R13469 VPWR.n2048 VPWR 0.100405
R13470 VPWR.n2049 VPWR 0.100405
R13471 VPWR.n2058 VPWR 0.100405
R13472 VPWR.n2059 VPWR 0.100405
R13473 VPWR.n2068 VPWR 0.100405
R13474 VPWR.n2069 VPWR 0.100405
R13475 VPWR.n2078 VPWR 0.100405
R13476 VPWR.n2079 VPWR 0.100405
R13477 VPWR.n2088 VPWR 0.100405
R13478 VPWR VPWR.n2012 0.100405
R13479 VPWR VPWR.n2013 0.100405
R13480 VPWR VPWR.n2014 0.100405
R13481 VPWR VPWR.n2015 0.100405
R13482 VPWR VPWR.n2026 0.100405
R13483 VPWR VPWR.n2025 0.100405
R13484 VPWR VPWR.n2024 0.100405
R13485 VPWR VPWR.n2023 0.100405
R13486 VPWR VPWR.n2022 0.100405
R13487 VPWR VPWR.n2021 0.100405
R13488 VPWR VPWR.n2020 0.100405
R13489 VPWR VPWR.n2019 0.100405
R13490 VPWR VPWR.n2018 0.100405
R13491 VPWR VPWR.n2017 0.100405
R13492 VPWR VPWR.n2016 0.100405
R13493 VPWR.n1932 VPWR 0.100405
R13494 VPWR VPWR.n1941 0.100405
R13495 VPWR.n1942 VPWR 0.100405
R13496 VPWR VPWR.n1951 0.100405
R13497 VPWR.n2002 VPWR 0.100405
R13498 VPWR VPWR.n2001 0.100405
R13499 VPWR.n1992 VPWR 0.100405
R13500 VPWR VPWR.n1991 0.100405
R13501 VPWR.n1982 VPWR 0.100405
R13502 VPWR VPWR.n1981 0.100405
R13503 VPWR.n1972 VPWR 0.100405
R13504 VPWR VPWR.n1971 0.100405
R13505 VPWR.n1962 VPWR 0.100405
R13506 VPWR VPWR.n1961 0.100405
R13507 VPWR.n1952 VPWR 0.100405
R13508 VPWR.n1929 VPWR 0.100405
R13509 VPWR.n1928 VPWR 0.100405
R13510 VPWR.n1927 VPWR 0.100405
R13511 VPWR.n1926 VPWR 0.100405
R13512 VPWR.n1915 VPWR 0.100405
R13513 VPWR.n1916 VPWR 0.100405
R13514 VPWR.n1917 VPWR 0.100405
R13515 VPWR.n1918 VPWR 0.100405
R13516 VPWR.n1919 VPWR 0.100405
R13517 VPWR.n1920 VPWR 0.100405
R13518 VPWR.n1921 VPWR 0.100405
R13519 VPWR.n1922 VPWR 0.100405
R13520 VPWR.n1923 VPWR 0.100405
R13521 VPWR.n1924 VPWR 0.100405
R13522 VPWR.n1925 VPWR 0.100405
R13523 VPWR VPWR.n2418 0.100405
R13524 VPWR VPWR.n2417 0.100405
R13525 VPWR VPWR.n2416 0.100405
R13526 VPWR VPWR.n2415 0.100405
R13527 VPWR VPWR.n2414 0.100405
R13528 VPWR VPWR.n2413 0.100405
R13529 VPWR VPWR.n2412 0.100405
R13530 VPWR VPWR.n2411 0.100405
R13531 VPWR VPWR.n2410 0.100405
R13532 VPWR VPWR.n2409 0.100405
R13533 VPWR VPWR.n2408 0.100405
R13534 VPWR VPWR.n2407 0.100405
R13535 VPWR.n1912 VPWR 0.100405
R13536 VPWR.n1903 VPWR 0.100405
R13537 VPWR.n1902 VPWR 0.100405
R13538 VPWR.n1893 VPWR 0.100405
R13539 VPWR.n1892 VPWR 0.100405
R13540 VPWR.n1842 VPWR 0.100405
R13541 VPWR.n1843 VPWR 0.100405
R13542 VPWR.n1852 VPWR 0.100405
R13543 VPWR.n1853 VPWR 0.100405
R13544 VPWR.n1862 VPWR 0.100405
R13545 VPWR.n1863 VPWR 0.100405
R13546 VPWR.n1872 VPWR 0.100405
R13547 VPWR.n1873 VPWR 0.100405
R13548 VPWR.n1882 VPWR 0.100405
R13549 VPWR.n1883 VPWR 0.100405
R13550 VPWR.n2430 VPWR 0.100405
R13551 VPWR.n2431 VPWR 0.100405
R13552 VPWR.n2440 VPWR 0.100405
R13553 VPWR.n2441 VPWR 0.100405
R13554 VPWR.n2450 VPWR 0.100405
R13555 VPWR.n2451 VPWR 0.100405
R13556 VPWR.n2460 VPWR 0.100405
R13557 VPWR.n2461 VPWR 0.100405
R13558 VPWR.n2470 VPWR 0.100405
R13559 VPWR.n2471 VPWR 0.100405
R13560 VPWR.n2480 VPWR 0.100405
R13561 VPWR.n2481 VPWR 0.100405
R13562 VPWR.n2490 VPWR 0.100405
R13563 VPWR VPWR.n1816 0.100405
R13564 VPWR VPWR.n1817 0.100405
R13565 VPWR VPWR.n1818 0.100405
R13566 VPWR VPWR.n1819 0.100405
R13567 VPWR VPWR.n1820 0.100405
R13568 VPWR VPWR.n1821 0.100405
R13569 VPWR VPWR.n1822 0.100405
R13570 VPWR VPWR.n1823 0.100405
R13571 VPWR VPWR.n1830 0.100405
R13572 VPWR VPWR.n1829 0.100405
R13573 VPWR VPWR.n1828 0.100405
R13574 VPWR VPWR.n1827 0.100405
R13575 VPWR VPWR.n1826 0.100405
R13576 VPWR VPWR.n1825 0.100405
R13577 VPWR VPWR.n1824 0.100405
R13578 VPWR.n2517 VPWR 0.100405
R13579 VPWR.n2516 VPWR 0.100405
R13580 VPWR.n2515 VPWR 0.100405
R13581 VPWR.n2514 VPWR 0.100405
R13582 VPWR.n2513 VPWR 0.100405
R13583 VPWR.n2512 VPWR 0.100405
R13584 VPWR.n2511 VPWR 0.100405
R13585 VPWR.n2510 VPWR 0.100405
R13586 VPWR.n2509 VPWR 0.100405
R13587 VPWR.n2508 VPWR 0.100405
R13588 VPWR.n2503 VPWR 0.100405
R13589 VPWR.n2504 VPWR 0.100405
R13590 VPWR.n2505 VPWR 0.100405
R13591 VPWR.n2506 VPWR 0.100405
R13592 VPWR.n2507 VPWR 0.100405
R13593 VPWR.n1162 VPWR 0.100405
R13594 VPWR VPWR.n1559 0.100405
R13595 VPWR.n1543 VPWR 0.100405
R13596 VPWR.n1535 VPWR 0.100405
R13597 VPWR.n1529 VPWR 0.100405
R13598 VPWR.n1521 VPWR 0.100405
R13599 VPWR.n1515 VPWR 0.100405
R13600 VPWR VPWR.n1151 0.100405
R13601 VPWR.n1603 VPWR 0.100405
R13602 VPWR.n1471 VPWR 0.100405
R13603 VPWR.n1483 VPWR 0.100405
R13604 VPWR.n1062 VPWR 0.100405
R13605 VPWR.n1763 VPWR 0.100405
R13606 VPWR.n1806 VPWR 0.100405
R13607 VPWR VPWR.n1784 0.100405
R13608 VPWR.n2520 VPWR 0.100405
R13609 VPWR VPWR.n2531 0.100405
R13610 VPWR.n2532 VPWR 0.100405
R13611 VPWR VPWR.n2543 0.100405
R13612 VPWR.n2544 VPWR 0.100405
R13613 VPWR VPWR.n2555 0.100405
R13614 VPWR.n2556 VPWR 0.100405
R13615 VPWR VPWR.n2567 0.100405
R13616 VPWR.n2568 VPWR 0.100405
R13617 VPWR VPWR.n2579 0.100405
R13618 VPWR.n2580 VPWR 0.100405
R13619 VPWR VPWR.n2591 0.100405
R13620 VPWR.n2592 VPWR 0.100405
R13621 VPWR VPWR.n2603 0.100405
R13622 VPWR.n2604 VPWR 0.100405
R13623 VPWR.n1075 VPWR 0.100405
R13624 VPWR.n1773 VPWR 0.100405
R13625 VPWR.n1774 VPWR 0.100405
R13626 VPWR.n1548 VPWR 0.100405
R13627 VPWR.n1549 VPWR 0.100405
R13628 VPWR VPWR.n1547 0.100405
R13629 VPWR VPWR.n1546 0.100405
R13630 VPWR.n1533 VPWR 0.100405
R13631 VPWR VPWR.n1532 0.100405
R13632 VPWR.n1519 VPWR 0.100405
R13633 VPWR VPWR.n1518 0.100405
R13634 VPWR.n1506 VPWR 0.100405
R13635 VPWR.n1606 VPWR 0.100405
R13636 VPWR.n1607 VPWR 0.100405
R13637 VPWR.n1467 VPWR 0.100405
R13638 VPWR VPWR.n2817 0.0994583
R13639 VPWR VPWR.n2798 0.0994583
R13640 VPWR VPWR.n1345 0.0981562
R13641 VPWR.n1390 VPWR 0.0981562
R13642 VPWR.n1429 VPWR 0.0981562
R13643 VPWR.n9 VPWR 0.0968542
R13644 VPWR.n1263 VPWR 0.0968542
R13645 VPWR.n1286 VPWR 0.0968542
R13646 VPWR.n1310 VPWR 0.0968542
R13647 VPWR.n1352 VPWR 0.0968542
R13648 VPWR VPWR.n2778 0.0968542
R13649 VPWR VPWR.n2759 0.0968542
R13650 VPWR.n2737 VPWR 0.0968542
R13651 VPWR.n2701 VPWR 0.0968542
R13652 VPWR.n2664 VPWR 0.0968542
R13653 VPWR.n2627 VPWR 0.0968542
R13654 VPWR VPWR.n1063 0.0945
R13655 VPWR.n1560 VPWR 0.0945
R13656 VPWR VPWR.n1161 0.0945
R13657 VPWR VPWR.n1160 0.0945
R13658 VPWR VPWR.n1159 0.0945
R13659 VPWR VPWR.n1158 0.0945
R13660 VPWR VPWR.n1157 0.0945
R13661 VPWR.n1156 VPWR 0.0945
R13662 VPWR VPWR.n1602 0.0945
R13663 VPWR VPWR.n1150 0.0945
R13664 VPWR VPWR.n1482 0.0945
R13665 VPWR.n1470 VPWR 0.0945
R13666 VPWR VPWR.n1057 0.0945
R13667 VPWR.n1805 VPWR 0.0945
R13668 VPWR VPWR.n1046 0.0945
R13669 VPWR.n1785 VPWR 0.0945
R13670 VPWR.n37 VPWR.n20 0.0939125
R13671 VPWR.n1136 VPWR 0.093504
R13672 VPWR.n128 VPWR 0.093504
R13673 VPWR.n162 VPWR 0.093504
R13674 VPWR.n174 VPWR 0.093504
R13675 VPWR.n186 VPWR 0.093504
R13676 VPWR.n198 VPWR 0.093504
R13677 VPWR.n210 VPWR 0.093504
R13678 VPWR.n222 VPWR 0.093504
R13679 VPWR.n234 VPWR 0.093504
R13680 VPWR.n246 VPWR 0.093504
R13681 VPWR.n258 VPWR 0.093504
R13682 VPWR.n270 VPWR 0.093504
R13683 VPWR.n282 VPWR 0.093504
R13684 VPWR.n294 VPWR 0.093504
R13685 VPWR VPWR.n304 0.093504
R13686 VPWR.n150 VPWR 0.093504
R13687 VPWR.n139 VPWR 0.093504
R13688 VPWR VPWR.n1750 0.093504
R13689 VPWR.n1741 VPWR 0.093504
R13690 VPWR.n1729 VPWR 0.093504
R13691 VPWR.n1718 VPWR 0.093504
R13692 VPWR VPWR.n1096 0.093504
R13693 VPWR.n1702 VPWR 0.093504
R13694 VPWR.n1691 VPWR 0.093504
R13695 VPWR VPWR.n1106 0.093504
R13696 VPWR.n1675 VPWR 0.093504
R13697 VPWR.n1664 VPWR 0.093504
R13698 VPWR VPWR.n1116 0.093504
R13699 VPWR.n1648 VPWR 0.093504
R13700 VPWR.n1637 VPWR 0.093504
R13701 VPWR VPWR.n1126 0.093504
R13702 VPWR.n1621 VPWR 0.093504
R13703 VPWR.n2617 VPWR 0.0849042
R13704 VPWR.n1131 VPWR.n1128 0.0845517
R13705 VPWR.n166 VPWR.n165 0.0845517
R13706 VPWR.n178 VPWR.n177 0.0845517
R13707 VPWR.n190 VPWR.n189 0.0845517
R13708 VPWR.n202 VPWR.n201 0.0845517
R13709 VPWR.n214 VPWR.n213 0.0845517
R13710 VPWR.n226 VPWR.n225 0.0845517
R13711 VPWR.n238 VPWR.n237 0.0845517
R13712 VPWR.n250 VPWR.n249 0.0845517
R13713 VPWR.n262 VPWR.n261 0.0845517
R13714 VPWR.n274 VPWR.n273 0.0845517
R13715 VPWR.n286 VPWR.n285 0.0845517
R13716 VPWR.n298 VPWR.n297 0.0845517
R13717 VPWR.n301 VPWR.n122 0.0845517
R13718 VPWR.n132 VPWR.n131 0.0845517
R13719 VPWR.n154 VPWR.n153 0.0845517
R13720 VPWR.n143 VPWR.n142 0.0845517
R13721 VPWR.n1747 VPWR.n1086 0.0845517
R13722 VPWR.n1745 VPWR.n1744 0.0845517
R13723 VPWR.n1733 VPWR.n1732 0.0845517
R13724 VPWR.n1720 VPWR.n1719 0.0845517
R13725 VPWR.n1709 VPWR.n1097 0.0845517
R13726 VPWR.n1706 VPWR.n1705 0.0845517
R13727 VPWR.n1693 VPWR.n1692 0.0845517
R13728 VPWR.n1682 VPWR.n1107 0.0845517
R13729 VPWR.n1679 VPWR.n1678 0.0845517
R13730 VPWR.n1666 VPWR.n1665 0.0845517
R13731 VPWR.n1655 VPWR.n1117 0.0845517
R13732 VPWR.n1652 VPWR.n1651 0.0845517
R13733 VPWR.n1639 VPWR.n1638 0.0845517
R13734 VPWR.n1628 VPWR.n1127 0.0845517
R13735 VPWR.n1625 VPWR.n1624 0.0845517
R13736 VPWR.n1475 VPWR.n1470 0.0740128
R13737 VPWR.n1561 VPWR.n1063 0.071
R13738 VPWR.n1566 VPWR.n1560 0.071
R13739 VPWR.n1571 VPWR.n1161 0.071
R13740 VPWR.n1576 VPWR.n1160 0.071
R13741 VPWR.n1581 VPWR.n1159 0.071
R13742 VPWR.n1586 VPWR.n1158 0.071
R13743 VPWR.n1591 VPWR.n1157 0.071
R13744 VPWR.n1596 VPWR.n1156 0.071
R13745 VPWR.n1602 VPWR.n1601 0.071
R13746 VPWR.n1476 VPWR.n1150 0.071
R13747 VPWR.n1482 VPWR.n1481 0.071
R13748 VPWR.n1791 VPWR.n1057 0.071
R13749 VPWR.n1805 VPWR.n1804 0.071
R13750 VPWR.n1799 VPWR.n1046 0.071
R13751 VPWR.n1786 VPWR.n1785 0.071
R13752 VPWR VPWR.n1134 0.0678077
R13753 VPWR VPWR.n126 0.0678077
R13754 VPWR VPWR.n160 0.0678077
R13755 VPWR VPWR.n172 0.0678077
R13756 VPWR VPWR.n184 0.0678077
R13757 VPWR VPWR.n196 0.0678077
R13758 VPWR VPWR.n208 0.0678077
R13759 VPWR VPWR.n220 0.0678077
R13760 VPWR VPWR.n232 0.0678077
R13761 VPWR VPWR.n244 0.0678077
R13762 VPWR VPWR.n256 0.0678077
R13763 VPWR VPWR.n268 0.0678077
R13764 VPWR VPWR.n280 0.0678077
R13765 VPWR VPWR.n292 0.0678077
R13766 VPWR.n305 VPWR 0.0678077
R13767 VPWR VPWR.n148 0.0678077
R13768 VPWR VPWR.n137 0.0678077
R13769 VPWR.n1751 VPWR 0.0678077
R13770 VPWR VPWR.n1739 0.0678077
R13771 VPWR VPWR.n1727 0.0678077
R13772 VPWR VPWR.n1716 0.0678077
R13773 VPWR.n1212 VPWR 0.0678077
R13774 VPWR VPWR.n1700 0.0678077
R13775 VPWR VPWR.n1689 0.0678077
R13776 VPWR.n1226 VPWR 0.0678077
R13777 VPWR VPWR.n1673 0.0678077
R13778 VPWR VPWR.n1662 0.0678077
R13779 VPWR.n1194 VPWR 0.0678077
R13780 VPWR VPWR.n1646 0.0678077
R13781 VPWR VPWR.n1635 0.0678077
R13782 VPWR.n1143 VPWR 0.0678077
R13783 VPWR VPWR.n1619 0.0678077
R13784 VPWR.n2845 VPWR 0.063
R13785 VPWR.n169 VPWR 0.063
R13786 VPWR.n181 VPWR 0.063
R13787 VPWR.n193 VPWR 0.063
R13788 VPWR.n205 VPWR 0.063
R13789 VPWR.n217 VPWR 0.063
R13790 VPWR.n229 VPWR 0.063
R13791 VPWR.n241 VPWR 0.063
R13792 VPWR.n253 VPWR 0.063
R13793 VPWR.n265 VPWR 0.063
R13794 VPWR.n277 VPWR 0.063
R13795 VPWR.n289 VPWR 0.063
R13796 VPWR.n120 VPWR 0.063
R13797 VPWR.n124 VPWR 0.063
R13798 VPWR.n157 VPWR 0.063
R13799 VPWR.n134 VPWR 0.063
R13800 VPWR.n145 VPWR 0.063
R13801 VPWR.n1084 VPWR 0.063
R13802 VPWR.n1736 VPWR 0.063
R13803 VPWR.n1089 VPWR 0.063
R13804 VPWR VPWR.n1723 0.063
R13805 VPWR VPWR.n1712 0.063
R13806 VPWR VPWR.n1100 0.063
R13807 VPWR VPWR.n1696 0.063
R13808 VPWR VPWR.n1685 0.063
R13809 VPWR VPWR.n1110 0.063
R13810 VPWR VPWR.n1669 0.063
R13811 VPWR VPWR.n1658 0.063
R13812 VPWR VPWR.n1120 0.063
R13813 VPWR VPWR.n1642 0.063
R13814 VPWR VPWR.n1631 0.063
R13815 VPWR VPWR.n1130 0.063
R13816 VPWR VPWR.n1139 0.063
R13817 VPWR.n1134 VPWR 0.0608448
R13818 VPWR.n126 VPWR 0.0608448
R13819 VPWR.n160 VPWR 0.0608448
R13820 VPWR.n172 VPWR 0.0608448
R13821 VPWR.n184 VPWR 0.0608448
R13822 VPWR.n196 VPWR 0.0608448
R13823 VPWR.n208 VPWR 0.0608448
R13824 VPWR.n220 VPWR 0.0608448
R13825 VPWR.n232 VPWR 0.0608448
R13826 VPWR.n244 VPWR 0.0608448
R13827 VPWR.n256 VPWR 0.0608448
R13828 VPWR.n268 VPWR 0.0608448
R13829 VPWR.n280 VPWR 0.0608448
R13830 VPWR.n292 VPWR 0.0608448
R13831 VPWR.n305 VPWR 0.0608448
R13832 VPWR.n148 VPWR 0.0608448
R13833 VPWR.n137 VPWR 0.0608448
R13834 VPWR.n1751 VPWR 0.0608448
R13835 VPWR.n1739 VPWR 0.0608448
R13836 VPWR.n1727 VPWR 0.0608448
R13837 VPWR.n1716 VPWR 0.0608448
R13838 VPWR.n1212 VPWR 0.0608448
R13839 VPWR.n1700 VPWR 0.0608448
R13840 VPWR.n1689 VPWR 0.0608448
R13841 VPWR.n1226 VPWR 0.0608448
R13842 VPWR.n1673 VPWR 0.0608448
R13843 VPWR.n1662 VPWR 0.0608448
R13844 VPWR.n1194 VPWR 0.0608448
R13845 VPWR.n1646 VPWR 0.0608448
R13846 VPWR.n1635 VPWR 0.0608448
R13847 VPWR.n1143 VPWR 0.0608448
R13848 VPWR.n1619 VPWR 0.0608448
R13849 VPWR VPWR.n13 0.0603958
R13850 VPWR VPWR.n12 0.0603958
R13851 VPWR VPWR.n1268 0.0603958
R13852 VPWR VPWR.n1267 0.0603958
R13853 VPWR VPWR.n1291 0.0603958
R13854 VPWR VPWR.n1290 0.0603958
R13855 VPWR VPWR.n1315 0.0603958
R13856 VPWR VPWR.n1314 0.0603958
R13857 VPWR.n1351 VPWR 0.0603958
R13858 VPWR VPWR.n1350 0.0603958
R13859 VPWR.n1346 VPWR 0.0603958
R13860 VPWR.n1337 VPWR 0.0603958
R13861 VPWR VPWR.n1336 0.0603958
R13862 VPWR.n1389 VPWR 0.0603958
R13863 VPWR VPWR.n1388 0.0603958
R13864 VPWR.n1383 VPWR 0.0603958
R13865 VPWR.n1428 VPWR 0.0603958
R13866 VPWR VPWR.n1427 0.0603958
R13867 VPWR.n1422 VPWR 0.0603958
R13868 VPWR.n1459 VPWR 0.0603958
R13869 VPWR VPWR.n2819 0.0603958
R13870 VPWR VPWR.n2818 0.0603958
R13871 VPWR VPWR.n2831 0.0603958
R13872 VPWR.n2810 VPWR 0.0603958
R13873 VPWR.n2811 VPWR 0.0603958
R13874 VPWR VPWR.n2815 0.0603958
R13875 VPWR.n2790 VPWR 0.0603958
R13876 VPWR.n2791 VPWR 0.0603958
R13877 VPWR VPWR.n2796 0.0603958
R13878 VPWR.n2771 VPWR 0.0603958
R13879 VPWR.n2772 VPWR 0.0603958
R13880 VPWR VPWR.n2776 0.0603958
R13881 VPWR.n2752 VPWR 0.0603958
R13882 VPWR.n2753 VPWR 0.0603958
R13883 VPWR VPWR.n2714 0.0603958
R13884 VPWR.n2715 VPWR 0.0603958
R13885 VPWR.n2716 VPWR 0.0603958
R13886 VPWR VPWR.n2677 0.0603958
R13887 VPWR.n2678 VPWR 0.0603958
R13888 VPWR.n2679 VPWR 0.0603958
R13889 VPWR.n2643 VPWR 0.0603958
R13890 VPWR.n2646 VPWR 0.0603958
R13891 VPWR.n1789 VPWR.n1788 0.0599512
R13892 VPWR.n1060 VPWR.n1059 0.0599512
R13893 VPWR.n1564 VPWR.n1563 0.0599512
R13894 VPWR.n1569 VPWR.n1568 0.0599512
R13895 VPWR.n1574 VPWR.n1573 0.0599512
R13896 VPWR.n1579 VPWR.n1578 0.0599512
R13897 VPWR.n1584 VPWR.n1583 0.0599512
R13898 VPWR.n1589 VPWR.n1588 0.0599512
R13899 VPWR.n1594 VPWR.n1593 0.0599512
R13900 VPWR.n1599 VPWR.n1598 0.0599512
R13901 VPWR.n1154 VPWR.n1153 0.0599512
R13902 VPWR.n1479 VPWR.n1478 0.0599512
R13903 VPWR.n1474 VPWR.n1473 0.0599512
R13904 VPWR.n1794 VPWR.n1793 0.0599512
R13905 VPWR.n1802 VPWR.n1801 0.0599512
R13906 VPWR.n1798 VPWR.n1797 0.0599512
R13907 VPWR.n1137 VPWR.n1136 0.0565345
R13908 VPWR.n1131 VPWR 0.0565345
R13909 VPWR.n163 VPWR.n162 0.0565345
R13910 VPWR.n165 VPWR 0.0565345
R13911 VPWR.n175 VPWR.n174 0.0565345
R13912 VPWR.n177 VPWR 0.0565345
R13913 VPWR.n187 VPWR.n186 0.0565345
R13914 VPWR.n189 VPWR 0.0565345
R13915 VPWR.n199 VPWR.n198 0.0565345
R13916 VPWR.n201 VPWR 0.0565345
R13917 VPWR.n211 VPWR.n210 0.0565345
R13918 VPWR.n213 VPWR 0.0565345
R13919 VPWR.n223 VPWR.n222 0.0565345
R13920 VPWR.n225 VPWR 0.0565345
R13921 VPWR.n235 VPWR.n234 0.0565345
R13922 VPWR.n237 VPWR 0.0565345
R13923 VPWR.n247 VPWR.n246 0.0565345
R13924 VPWR.n249 VPWR 0.0565345
R13925 VPWR.n259 VPWR.n258 0.0565345
R13926 VPWR.n261 VPWR 0.0565345
R13927 VPWR.n271 VPWR.n270 0.0565345
R13928 VPWR.n273 VPWR 0.0565345
R13929 VPWR.n283 VPWR.n282 0.0565345
R13930 VPWR.n285 VPWR 0.0565345
R13931 VPWR.n295 VPWR.n294 0.0565345
R13932 VPWR.n297 VPWR 0.0565345
R13933 VPWR.n304 VPWR.n302 0.0565345
R13934 VPWR.n122 VPWR 0.0565345
R13935 VPWR.n129 VPWR.n128 0.0565345
R13936 VPWR.n131 VPWR 0.0565345
R13937 VPWR.n151 VPWR.n150 0.0565345
R13938 VPWR.n153 VPWR 0.0565345
R13939 VPWR.n140 VPWR.n139 0.0565345
R13940 VPWR.n142 VPWR 0.0565345
R13941 VPWR.n1750 VPWR.n1748 0.0565345
R13942 VPWR.n1086 VPWR 0.0565345
R13943 VPWR.n1742 VPWR.n1741 0.0565345
R13944 VPWR.n1744 VPWR 0.0565345
R13945 VPWR.n1730 VPWR.n1729 0.0565345
R13946 VPWR.n1732 VPWR 0.0565345
R13947 VPWR.n1721 VPWR.n1718 0.0565345
R13948 VPWR.n1719 VPWR 0.0565345
R13949 VPWR.n1710 VPWR.n1096 0.0565345
R13950 VPWR.n1097 VPWR 0.0565345
R13951 VPWR.n1703 VPWR.n1702 0.0565345
R13952 VPWR.n1705 VPWR 0.0565345
R13953 VPWR.n1694 VPWR.n1691 0.0565345
R13954 VPWR.n1692 VPWR 0.0565345
R13955 VPWR.n1683 VPWR.n1106 0.0565345
R13956 VPWR.n1107 VPWR 0.0565345
R13957 VPWR.n1676 VPWR.n1675 0.0565345
R13958 VPWR.n1678 VPWR 0.0565345
R13959 VPWR.n1667 VPWR.n1664 0.0565345
R13960 VPWR.n1665 VPWR 0.0565345
R13961 VPWR.n1656 VPWR.n1116 0.0565345
R13962 VPWR.n1117 VPWR 0.0565345
R13963 VPWR.n1649 VPWR.n1648 0.0565345
R13964 VPWR.n1651 VPWR 0.0565345
R13965 VPWR.n1640 VPWR.n1637 0.0565345
R13966 VPWR.n1638 VPWR 0.0565345
R13967 VPWR.n1629 VPWR.n1126 0.0565345
R13968 VPWR.n1127 VPWR 0.0565345
R13969 VPWR.n1622 VPWR.n1621 0.0565345
R13970 VPWR.n1624 VPWR 0.0565345
R13971 VPWR.n1788 VPWR 0.0469286
R13972 VPWR.n1059 VPWR 0.0469286
R13973 VPWR.n1563 VPWR 0.0469286
R13974 VPWR.n1568 VPWR 0.0469286
R13975 VPWR.n1573 VPWR 0.0469286
R13976 VPWR.n1578 VPWR 0.0469286
R13977 VPWR.n1583 VPWR 0.0469286
R13978 VPWR.n1588 VPWR 0.0469286
R13979 VPWR.n1593 VPWR 0.0469286
R13980 VPWR.n1598 VPWR 0.0469286
R13981 VPWR.n1153 VPWR 0.0469286
R13982 VPWR.n1478 VPWR 0.0469286
R13983 VPWR.n1473 VPWR 0.0469286
R13984 VPWR.n1793 VPWR 0.0469286
R13985 VPWR.n1801 VPWR 0.0469286
R13986 VPWR.n1797 VPWR 0.0469286
R13987 VPWR.n1788 VPWR 0.0401341
R13988 VPWR.n1059 VPWR 0.0401341
R13989 VPWR.n1563 VPWR 0.0401341
R13990 VPWR.n1568 VPWR 0.0401341
R13991 VPWR.n1573 VPWR 0.0401341
R13992 VPWR.n1578 VPWR 0.0401341
R13993 VPWR.n1583 VPWR 0.0401341
R13994 VPWR.n1588 VPWR 0.0401341
R13995 VPWR.n1593 VPWR 0.0401341
R13996 VPWR.n1598 VPWR 0.0401341
R13997 VPWR.n1153 VPWR 0.0401341
R13998 VPWR.n1478 VPWR 0.0401341
R13999 VPWR.n1473 VPWR 0.0401341
R14000 VPWR.n1793 VPWR 0.0401341
R14001 VPWR.n1801 VPWR 0.0401341
R14002 VPWR.n1797 VPWR 0.0401341
R14003 VPWR.n13 VPWR 0.0382604
R14004 VPWR.n1268 VPWR 0.0382604
R14005 VPWR.n1291 VPWR 0.0382604
R14006 VPWR.n1315 VPWR 0.0382604
R14007 VPWR.n1350 VPWR 0.0382604
R14008 VPWR.n1388 VPWR 0.0382604
R14009 VPWR.n1427 VPWR 0.0382604
R14010 VPWR.n1464 VPWR 0.0382604
R14011 VPWR.n39 VPWR 0.0375125
R14012 VPWR.n39 VPWR 0.0373589
R14013 VPWR.n1137 VPWR.n1128 0.0349828
R14014 VPWR.n166 VPWR.n163 0.0349828
R14015 VPWR.n178 VPWR.n175 0.0349828
R14016 VPWR.n190 VPWR.n187 0.0349828
R14017 VPWR.n202 VPWR.n199 0.0349828
R14018 VPWR.n214 VPWR.n211 0.0349828
R14019 VPWR.n226 VPWR.n223 0.0349828
R14020 VPWR.n238 VPWR.n235 0.0349828
R14021 VPWR.n250 VPWR.n247 0.0349828
R14022 VPWR.n262 VPWR.n259 0.0349828
R14023 VPWR.n274 VPWR.n271 0.0349828
R14024 VPWR.n286 VPWR.n283 0.0349828
R14025 VPWR.n298 VPWR.n295 0.0349828
R14026 VPWR.n302 VPWR.n301 0.0349828
R14027 VPWR.n132 VPWR.n129 0.0349828
R14028 VPWR.n154 VPWR.n151 0.0349828
R14029 VPWR.n143 VPWR.n140 0.0349828
R14030 VPWR.n1748 VPWR.n1747 0.0349828
R14031 VPWR.n1745 VPWR.n1742 0.0349828
R14032 VPWR.n1733 VPWR.n1730 0.0349828
R14033 VPWR.n1721 VPWR.n1720 0.0349828
R14034 VPWR.n1710 VPWR.n1709 0.0349828
R14035 VPWR.n1706 VPWR.n1703 0.0349828
R14036 VPWR.n1694 VPWR.n1693 0.0349828
R14037 VPWR.n1683 VPWR.n1682 0.0349828
R14038 VPWR.n1679 VPWR.n1676 0.0349828
R14039 VPWR.n1667 VPWR.n1666 0.0349828
R14040 VPWR.n1656 VPWR.n1655 0.0349828
R14041 VPWR.n1652 VPWR.n1649 0.0349828
R14042 VPWR.n1640 VPWR.n1639 0.0349828
R14043 VPWR.n1629 VPWR.n1628 0.0349828
R14044 VPWR.n1625 VPWR.n1622 0.0349828
R14045 VPWR.n2523 VPWR.n2522 0.0340366
R14046 VPWR.n2589 VPWR.n2588 0.0340366
R14047 VPWR.n2529 VPWR.n2528 0.0340366
R14048 VPWR.n2571 VPWR.n2570 0.0340366
R14049 VPWR.n2565 VPWR.n2564 0.0340366
R14050 VPWR.n2553 VPWR.n2552 0.0340366
R14051 VPWR.n2547 VPWR.n2546 0.0340366
R14052 VPWR.n1242 VPWR.n1241 0.0340366
R14053 VPWR.n2541 VPWR.n2540 0.0340366
R14054 VPWR.n1505 VPWR.n1121 0.0340366
R14055 VPWR.n1193 VPWR.n1113 0.0340366
R14056 VPWR.n2559 VPWR.n2558 0.0340366
R14057 VPWR.n1184 VPWR.n1111 0.0340366
R14058 VPWR.n1230 VPWR.n1183 0.0340366
R14059 VPWR.n2535 VPWR.n2534 0.0340366
R14060 VPWR.n1148 VPWR.n1123 0.0340366
R14061 VPWR.n1174 VPWR.n1103 0.0340366
R14062 VPWR.n2577 VPWR.n2576 0.0340366
R14063 VPWR.n1163 VPWR.n1101 0.0340366
R14064 VPWR.n1610 VPWR.n1609 0.0340366
R14065 VPWR.n2583 VPWR.n2582 0.0340366
R14066 VPWR.n1216 VPWR.n1173 0.0340366
R14067 VPWR.n1093 VPWR.n1092 0.0340366
R14068 VPWR.n1762 VPWR.n1761 0.0340366
R14069 VPWR.n1090 VPWR.n1073 0.0340366
R14070 VPWR.n2595 VPWR.n2594 0.0340366
R14071 VPWR.n2601 VPWR.n2600 0.0340366
R14072 VPWR.n2612 VPWR.n2611 0.0340366
R14073 VPWR.n2607 VPWR.n2606 0.0340366
R14074 VPWR.n1756 VPWR.n1755 0.0340366
R14075 VPWR.n1082 VPWR.n1079 0.0340366
R14076 VPWR.n1615 VPWR.n1140 0.0340366
R14077 VPWR.n2647 VPWR.n2617 0.0320292
R14078 VPWR VPWR.n22 0.03175
R14079 VPWR.n2819 VPWR 0.03175
R14080 VPWR VPWR.n2810 0.03175
R14081 VPWR VPWR.n2790 0.03175
R14082 VPWR VPWR.n2771 0.03175
R14083 VPWR VPWR.n2752 0.03175
R14084 VPWR VPWR.n2715 0.03175
R14085 VPWR VPWR.n2678 0.03175
R14086 VPWR VPWR.n2646 0.03175
R14087 VPWR.n2617 VPWR.n2616 0.0240975
R14088 VPWR.n2616 VPWR.n39 0.0240975
R14089 VPWR.n38 VPWR 0.024
R14090 VPWR.n14 VPWR 0.0239375
R14091 VPWR.n12 VPWR 0.0239375
R14092 VPWR.n1269 VPWR 0.0239375
R14093 VPWR.n1267 VPWR 0.0239375
R14094 VPWR.n1290 VPWR 0.0239375
R14095 VPWR.n1314 VPWR 0.0239375
R14096 VPWR.n2772 VPWR 0.0239375
R14097 VPWR.n2522 VPWR 0.0233659
R14098 VPWR.n1485 VPWR 0.0233659
R14099 VPWR.n371 VPWR 0.0233659
R14100 VPWR.n2589 VPWR 0.0233659
R14101 VPWR.n1552 VPWR 0.0233659
R14102 VPWR.n366 VPWR 0.0233659
R14103 VPWR.n2529 VPWR 0.0233659
R14104 VPWR.n983 VPWR 0.0233659
R14105 VPWR.n2498 VPWR 0.0233659
R14106 VPWR.n2493 VPWR 0.0233659
R14107 VPWR.n338 VPWR 0.0233659
R14108 VPWR.n2570 VPWR 0.0233659
R14109 VPWR.n991 VPWR 0.0233659
R14110 VPWR.n2463 VPWR 0.0233659
R14111 VPWR.n342 VPWR 0.0233659
R14112 VPWR.n2565 VPWR 0.0233659
R14113 VPWR.n1910 VPWR 0.0233659
R14114 VPWR.n1905 VPWR 0.0233659
R14115 VPWR.n1900 VPWR 0.0233659
R14116 VPWR.n407 VPWR 0.0233659
R14117 VPWR.n411 VPWR 0.0233659
R14118 VPWR.n415 VPWR 0.0233659
R14119 VPWR.n2473 VPWR 0.0233659
R14120 VPWR.n350 VPWR 0.0233659
R14121 VPWR.n2553 VPWR 0.0233659
R14122 VPWR.n1895 VPWR 0.0233659
R14123 VPWR.n423 VPWR 0.0233659
R14124 VPWR.n2478 VPWR 0.0233659
R14125 VPWR.n354 VPWR 0.0233659
R14126 VPWR.n2546 VPWR 0.0233659
R14127 VPWR.n2326 VPWR 0.0233659
R14128 VPWR.n2331 VPWR 0.0233659
R14129 VPWR.n2336 VPWR 0.0233659
R14130 VPWR.n2341 VPWR 0.0233659
R14131 VPWR.n2351 VPWR 0.0233659
R14132 VPWR.n2356 VPWR 0.0233659
R14133 VPWR.n2361 VPWR 0.0233659
R14134 VPWR.n2366 VPWR 0.0233659
R14135 VPWR.n2371 VPWR 0.0233659
R14136 VPWR.n2376 VPWR 0.0233659
R14137 VPWR.n2381 VPWR 0.0233659
R14138 VPWR.n2386 VPWR 0.0233659
R14139 VPWR.n2391 VPWR 0.0233659
R14140 VPWR.n2396 VPWR 0.0233659
R14141 VPWR.n2400 VPWR 0.0233659
R14142 VPWR.n2346 VPWR 0.0233659
R14143 VPWR.n563 VPWR 0.0233659
R14144 VPWR.n558 VPWR 0.0233659
R14145 VPWR.n554 VPWR 0.0233659
R14146 VPWR.n550 VPWR 0.0233659
R14147 VPWR.n542 VPWR 0.0233659
R14148 VPWR.n538 VPWR 0.0233659
R14149 VPWR.n534 VPWR 0.0233659
R14150 VPWR.n530 VPWR 0.0233659
R14151 VPWR.n526 VPWR 0.0233659
R14152 VPWR.n522 VPWR 0.0233659
R14153 VPWR.n518 VPWR 0.0233659
R14154 VPWR.n514 VPWR 0.0233659
R14155 VPWR.n510 VPWR 0.0233659
R14156 VPWR.n506 VPWR 0.0233659
R14157 VPWR.n503 VPWR 0.0233659
R14158 VPWR.n546 VPWR 0.0233659
R14159 VPWR.n2302 VPWR 0.0233659
R14160 VPWR.n2297 VPWR 0.0233659
R14161 VPWR.n2292 VPWR 0.0233659
R14162 VPWR.n2287 VPWR 0.0233659
R14163 VPWR.n2277 VPWR 0.0233659
R14164 VPWR.n2272 VPWR 0.0233659
R14165 VPWR.n2267 VPWR 0.0233659
R14166 VPWR.n2262 VPWR 0.0233659
R14167 VPWR.n2257 VPWR 0.0233659
R14168 VPWR.n2252 VPWR 0.0233659
R14169 VPWR.n2247 VPWR 0.0233659
R14170 VPWR.n2242 VPWR 0.0233659
R14171 VPWR.n2237 VPWR 0.0233659
R14172 VPWR.n2232 VPWR 0.0233659
R14173 VPWR.n2228 VPWR 0.0233659
R14174 VPWR.n2282 VPWR 0.0233659
R14175 VPWR.n599 VPWR 0.0233659
R14176 VPWR.n603 VPWR 0.0233659
R14177 VPWR.n607 VPWR 0.0233659
R14178 VPWR.n611 VPWR 0.0233659
R14179 VPWR.n619 VPWR 0.0233659
R14180 VPWR.n623 VPWR 0.0233659
R14181 VPWR.n627 VPWR 0.0233659
R14182 VPWR.n631 VPWR 0.0233659
R14183 VPWR.n635 VPWR 0.0233659
R14184 VPWR.n639 VPWR 0.0233659
R14185 VPWR.n643 VPWR 0.0233659
R14186 VPWR.n647 VPWR 0.0233659
R14187 VPWR.n651 VPWR 0.0233659
R14188 VPWR.n655 VPWR 0.0233659
R14189 VPWR.n659 VPWR 0.0233659
R14190 VPWR.n615 VPWR 0.0233659
R14191 VPWR.n2130 VPWR 0.0233659
R14192 VPWR.n2135 VPWR 0.0233659
R14193 VPWR.n2140 VPWR 0.0233659
R14194 VPWR.n2145 VPWR 0.0233659
R14195 VPWR.n2155 VPWR 0.0233659
R14196 VPWR.n2160 VPWR 0.0233659
R14197 VPWR.n2165 VPWR 0.0233659
R14198 VPWR.n2170 VPWR 0.0233659
R14199 VPWR.n2175 VPWR 0.0233659
R14200 VPWR.n2180 VPWR 0.0233659
R14201 VPWR.n2185 VPWR 0.0233659
R14202 VPWR.n2190 VPWR 0.0233659
R14203 VPWR.n2195 VPWR 0.0233659
R14204 VPWR.n2200 VPWR 0.0233659
R14205 VPWR.n2204 VPWR 0.0233659
R14206 VPWR.n2150 VPWR 0.0233659
R14207 VPWR.n755 VPWR 0.0233659
R14208 VPWR.n750 VPWR 0.0233659
R14209 VPWR.n746 VPWR 0.0233659
R14210 VPWR.n742 VPWR 0.0233659
R14211 VPWR.n734 VPWR 0.0233659
R14212 VPWR.n730 VPWR 0.0233659
R14213 VPWR.n726 VPWR 0.0233659
R14214 VPWR.n722 VPWR 0.0233659
R14215 VPWR.n718 VPWR 0.0233659
R14216 VPWR.n714 VPWR 0.0233659
R14217 VPWR.n710 VPWR 0.0233659
R14218 VPWR.n706 VPWR 0.0233659
R14219 VPWR.n702 VPWR 0.0233659
R14220 VPWR.n698 VPWR 0.0233659
R14221 VPWR.n695 VPWR 0.0233659
R14222 VPWR.n738 VPWR 0.0233659
R14223 VPWR.n2106 VPWR 0.0233659
R14224 VPWR.n2101 VPWR 0.0233659
R14225 VPWR.n2096 VPWR 0.0233659
R14226 VPWR.n2091 VPWR 0.0233659
R14227 VPWR.n2081 VPWR 0.0233659
R14228 VPWR.n2076 VPWR 0.0233659
R14229 VPWR.n2071 VPWR 0.0233659
R14230 VPWR.n2066 VPWR 0.0233659
R14231 VPWR.n2061 VPWR 0.0233659
R14232 VPWR.n2056 VPWR 0.0233659
R14233 VPWR.n2051 VPWR 0.0233659
R14234 VPWR.n2046 VPWR 0.0233659
R14235 VPWR.n2041 VPWR 0.0233659
R14236 VPWR.n2036 VPWR 0.0233659
R14237 VPWR.n2032 VPWR 0.0233659
R14238 VPWR.n2086 VPWR 0.0233659
R14239 VPWR.n791 VPWR 0.0233659
R14240 VPWR.n795 VPWR 0.0233659
R14241 VPWR.n799 VPWR 0.0233659
R14242 VPWR.n803 VPWR 0.0233659
R14243 VPWR.n811 VPWR 0.0233659
R14244 VPWR.n815 VPWR 0.0233659
R14245 VPWR.n819 VPWR 0.0233659
R14246 VPWR.n823 VPWR 0.0233659
R14247 VPWR.n827 VPWR 0.0233659
R14248 VPWR.n831 VPWR 0.0233659
R14249 VPWR.n835 VPWR 0.0233659
R14250 VPWR.n839 VPWR 0.0233659
R14251 VPWR.n843 VPWR 0.0233659
R14252 VPWR.n847 VPWR 0.0233659
R14253 VPWR.n851 VPWR 0.0233659
R14254 VPWR.n807 VPWR 0.0233659
R14255 VPWR.n1934 VPWR 0.0233659
R14256 VPWR.n1939 VPWR 0.0233659
R14257 VPWR.n1944 VPWR 0.0233659
R14258 VPWR.n1949 VPWR 0.0233659
R14259 VPWR.n1959 VPWR 0.0233659
R14260 VPWR.n1964 VPWR 0.0233659
R14261 VPWR.n1969 VPWR 0.0233659
R14262 VPWR.n1974 VPWR 0.0233659
R14263 VPWR.n1979 VPWR 0.0233659
R14264 VPWR.n1984 VPWR 0.0233659
R14265 VPWR.n1989 VPWR 0.0233659
R14266 VPWR.n1994 VPWR 0.0233659
R14267 VPWR.n1999 VPWR 0.0233659
R14268 VPWR.n2004 VPWR 0.0233659
R14269 VPWR.n2008 VPWR 0.0233659
R14270 VPWR.n1954 VPWR 0.0233659
R14271 VPWR.n947 VPWR 0.0233659
R14272 VPWR.n942 VPWR 0.0233659
R14273 VPWR.n938 VPWR 0.0233659
R14274 VPWR.n934 VPWR 0.0233659
R14275 VPWR.n926 VPWR 0.0233659
R14276 VPWR.n922 VPWR 0.0233659
R14277 VPWR.n918 VPWR 0.0233659
R14278 VPWR.n914 VPWR 0.0233659
R14279 VPWR.n910 VPWR 0.0233659
R14280 VPWR.n906 VPWR 0.0233659
R14281 VPWR.n902 VPWR 0.0233659
R14282 VPWR.n898 VPWR 0.0233659
R14283 VPWR.n894 VPWR 0.0233659
R14284 VPWR.n890 VPWR 0.0233659
R14285 VPWR.n887 VPWR 0.0233659
R14286 VPWR.n930 VPWR 0.0233659
R14287 VPWR.n1890 VPWR 0.0233659
R14288 VPWR.n999 VPWR 0.0233659
R14289 VPWR.n1514 VPWR 0.0233659
R14290 VPWR.n1242 VPWR 0.0233659
R14291 VPWR.n419 VPWR 0.0233659
R14292 VPWR.n2483 VPWR 0.0233659
R14293 VPWR.n358 VPWR 0.0233659
R14294 VPWR.n2541 VPWR 0.0233659
R14295 VPWR.n995 VPWR 0.0233659
R14296 VPWR.n1509 VPWR 0.0233659
R14297 VPWR.n1505 VPWR 0.0233659
R14298 VPWR.n1885 VPWR 0.0233659
R14299 VPWR.n1003 VPWR 0.0233659
R14300 VPWR.n1523 VPWR 0.0233659
R14301 VPWR.n1193 VPWR 0.0233659
R14302 VPWR.n427 VPWR 0.0233659
R14303 VPWR.n435 VPWR 0.0233659
R14304 VPWR.n439 VPWR 0.0233659
R14305 VPWR.n443 VPWR 0.0233659
R14306 VPWR.n447 VPWR 0.0233659
R14307 VPWR.n451 VPWR 0.0233659
R14308 VPWR.n455 VPWR 0.0233659
R14309 VPWR.n459 VPWR 0.0233659
R14310 VPWR.n463 VPWR 0.0233659
R14311 VPWR.n467 VPWR 0.0233659
R14312 VPWR.n431 VPWR 0.0233659
R14313 VPWR.n2468 VPWR 0.0233659
R14314 VPWR.n346 VPWR 0.0233659
R14315 VPWR.n2558 VPWR 0.0233659
R14316 VPWR.n1007 VPWR 0.0233659
R14317 VPWR.n1528 VPWR 0.0233659
R14318 VPWR.n1184 VPWR 0.0233659
R14319 VPWR.n1880 VPWR 0.0233659
R14320 VPWR.n1870 VPWR 0.0233659
R14321 VPWR.n1865 VPWR 0.0233659
R14322 VPWR.n1860 VPWR 0.0233659
R14323 VPWR.n1855 VPWR 0.0233659
R14324 VPWR.n1850 VPWR 0.0233659
R14325 VPWR.n1845 VPWR 0.0233659
R14326 VPWR.n1840 VPWR 0.0233659
R14327 VPWR.n1836 VPWR 0.0233659
R14328 VPWR.n1875 VPWR 0.0233659
R14329 VPWR.n1011 VPWR 0.0233659
R14330 VPWR.n1537 VPWR 0.0233659
R14331 VPWR.n1183 VPWR 0.0233659
R14332 VPWR.n2488 VPWR 0.0233659
R14333 VPWR.n362 VPWR 0.0233659
R14334 VPWR.n2534 VPWR 0.0233659
R14335 VPWR.n1149 VPWR 0.0233659
R14336 VPWR.n1148 VPWR 0.0233659
R14337 VPWR.n1015 VPWR 0.0233659
R14338 VPWR.n1542 VPWR 0.0233659
R14339 VPWR.n1174 VPWR 0.0233659
R14340 VPWR.n2458 VPWR 0.0233659
R14341 VPWR.n2448 VPWR 0.0233659
R14342 VPWR.n2443 VPWR 0.0233659
R14343 VPWR.n2438 VPWR 0.0233659
R14344 VPWR.n2433 VPWR 0.0233659
R14345 VPWR.n2428 VPWR 0.0233659
R14346 VPWR.n2424 VPWR 0.0233659
R14347 VPWR.n2453 VPWR 0.0233659
R14348 VPWR.n334 VPWR 0.0233659
R14349 VPWR.n2577 VPWR 0.0233659
R14350 VPWR.n1557 VPWR 0.0233659
R14351 VPWR.n1163 VPWR 0.0233659
R14352 VPWR.n1019 VPWR 0.0233659
R14353 VPWR.n1023 VPWR 0.0233659
R14354 VPWR.n1027 VPWR 0.0233659
R14355 VPWR.n1031 VPWR 0.0233659
R14356 VPWR.n1035 VPWR 0.0233659
R14357 VPWR.n1039 VPWR 0.0233659
R14358 VPWR.n1043 VPWR 0.0233659
R14359 VPWR.n987 VPWR 0.0233659
R14360 VPWR.n1492 VPWR 0.0233659
R14361 VPWR.n1609 VPWR 0.0233659
R14362 VPWR.n330 VPWR 0.0233659
R14363 VPWR.n2582 VPWR 0.0233659
R14364 VPWR.n1173 VPWR 0.0233659
R14365 VPWR.n1782 VPWR 0.0233659
R14366 VPWR.n1092 VPWR 0.0233659
R14367 VPWR.n326 VPWR 0.0233659
R14368 VPWR.n322 VPWR 0.0233659
R14369 VPWR.n314 VPWR 0.0233659
R14370 VPWR.n311 VPWR 0.0233659
R14371 VPWR.n318 VPWR 0.0233659
R14372 VPWR.n1762 VPWR 0.0233659
R14373 VPWR.n1770 VPWR 0.0233659
R14374 VPWR.n1808 VPWR 0.0233659
R14375 VPWR.n1812 VPWR 0.0233659
R14376 VPWR.n1777 VPWR 0.0233659
R14377 VPWR.n1073 VPWR 0.0233659
R14378 VPWR.n2594 VPWR 0.0233659
R14379 VPWR.n2601 VPWR 0.0233659
R14380 VPWR.n2612 VPWR 0.0233659
R14381 VPWR.n2606 VPWR 0.0233659
R14382 VPWR.n1755 VPWR 0.0233659
R14383 VPWR.n1079 VPWR 0.0233659
R14384 VPWR.n1140 VPWR 0.0233659
R14385 VPWR.n1355 VPWR 0.0226354
R14386 VPWR.n1346 VPWR 0.0226354
R14387 VPWR.n1432 VPWR 0.0226354
R14388 VPWR.n2791 VPWR 0.0226354
R14389 VPWR VPWR.n2751 0.0226354
R14390 VPWR VPWR.n2721 0.0226354
R14391 VPWR VPWR.n2683 0.0226354
R14392 VPWR VPWR.n83 0.0220517
R14393 VPWR VPWR.n86 0.0220517
R14394 VPWR VPWR.n89 0.0220517
R14395 VPWR VPWR.n92 0.0220517
R14396 VPWR VPWR.n95 0.0220517
R14397 VPWR VPWR.n98 0.0220517
R14398 VPWR VPWR.n101 0.0220517
R14399 VPWR VPWR.n104 0.0220517
R14400 VPWR VPWR.n107 0.0220517
R14401 VPWR VPWR.n110 0.0220517
R14402 VPWR VPWR.n113 0.0220517
R14403 VPWR VPWR.n116 0.0220517
R14404 VPWR.n308 VPWR 0.0220517
R14405 VPWR VPWR.n80 0.0220517
R14406 VPWR VPWR.n77 0.0220517
R14407 VPWR.n1754 VPWR 0.0220517
R14408 VPWR VPWR.n1076 0.0220517
R14409 VPWR.n1724 VPWR 0.0220517
R14410 VPWR.n1713 VPWR 0.0220517
R14411 VPWR.n1215 VPWR 0.0220517
R14412 VPWR.n1697 VPWR 0.0220517
R14413 VPWR.n1686 VPWR 0.0220517
R14414 VPWR.n1229 VPWR 0.0220517
R14415 VPWR.n1670 VPWR 0.0220517
R14416 VPWR.n1659 VPWR 0.0220517
R14417 VPWR.n1197 VPWR 0.0220517
R14418 VPWR.n1643 VPWR 0.0220517
R14419 VPWR.n1632 VPWR 0.0220517
R14420 VPWR.n1146 VPWR 0.0220517
R14421 VPWR.n1616 VPWR 0.0220517
R14422 VPWR.n1292 VPWR 0.0213333
R14423 VPWR.n1316 VPWR 0.0213333
R14424 VPWR.n1330 VPWR 0.0213333
R14425 VPWR.n1394 VPWR 0.0213333
R14426 VPWR.n1366 VPWR 0.0213333
R14427 VPWR.n1405 VPWR 0.0213333
R14428 VPWR.n1442 VPWR 0.0213333
R14429 VPWR.n2825 VPWR 0.0213333
R14430 VPWR.n2818 VPWR 0.0213333
R14431 VPWR VPWR.n2809 0.0213333
R14432 VPWR.n2811 VPWR 0.0213333
R14433 VPWR VPWR.n2789 0.0213333
R14434 VPWR VPWR.n2770 0.0213333
R14435 VPWR VPWR.n2757 0.0213333
R14436 VPWR.n2519 VPWR 0.0196917
R14437 VPWR.n43 VPWR 0.0143889
R14438 VPWR VPWR.n19 0.0099
R14439 VPWR VPWR.n1623 0.00397222
R14440 VPWR VPWR.n1124 0.00397222
R14441 VPWR VPWR.n1122 0.00397222
R14442 VPWR VPWR.n1650 0.00397222
R14443 VPWR VPWR.n1114 0.00397222
R14444 VPWR VPWR.n1112 0.00397222
R14445 VPWR VPWR.n1677 0.00397222
R14446 VPWR VPWR.n1104 0.00397222
R14447 VPWR VPWR.n1102 0.00397222
R14448 VPWR VPWR.n1704 0.00397222
R14449 VPWR VPWR.n1094 0.00397222
R14450 VPWR VPWR.n1091 0.00397222
R14451 VPWR VPWR.n1731 0.00397222
R14452 VPWR VPWR.n1743 0.00397222
R14453 VPWR.n1132 VPWR 0.00397222
R14454 VPWR VPWR.n1085 0.00397222
R14455 VPWR VPWR.n141 0.00397222
R14456 VPWR VPWR.n130 0.00397222
R14457 VPWR VPWR.n121 0.00397222
R14458 VPWR VPWR.n296 0.00397222
R14459 VPWR VPWR.n284 0.00397222
R14460 VPWR VPWR.n272 0.00397222
R14461 VPWR VPWR.n260 0.00397222
R14462 VPWR VPWR.n248 0.00397222
R14463 VPWR VPWR.n236 0.00397222
R14464 VPWR VPWR.n224 0.00397222
R14465 VPWR VPWR.n212 0.00397222
R14466 VPWR VPWR.n200 0.00397222
R14467 VPWR VPWR.n188 0.00397222
R14468 VPWR VPWR.n176 0.00397222
R14469 VPWR VPWR.n164 0.00397222
R14470 VPWR VPWR.n152 0.00397222
R14471 VPWR.n1481 VPWR.n1480 0.00351282
R14472 VPWR.n1476 VPWR.n1155 0.00351282
R14473 VPWR.n1601 VPWR.n1600 0.00351282
R14474 VPWR.n1596 VPWR.n1595 0.00351282
R14475 VPWR.n1591 VPWR.n1590 0.00351282
R14476 VPWR.n1586 VPWR.n1585 0.00351282
R14477 VPWR.n1581 VPWR.n1580 0.00351282
R14478 VPWR.n1576 VPWR.n1575 0.00351282
R14479 VPWR.n1571 VPWR.n1570 0.00351282
R14480 VPWR.n1566 VPWR.n1565 0.00351282
R14481 VPWR.n1561 VPWR.n1061 0.00351282
R14482 VPWR.n1804 VPWR.n1803 0.00351282
R14483 VPWR.n1795 VPWR.n1791 0.00351282
R14484 VPWR.n1790 VPWR.n1786 0.00351282
R14485 VPWR.n160 VPWR.n159 0.00265517
R14486 VPWR.n172 VPWR.n171 0.00265517
R14487 VPWR.n184 VPWR.n183 0.00265517
R14488 VPWR.n196 VPWR.n195 0.00265517
R14489 VPWR.n208 VPWR.n207 0.00265517
R14490 VPWR.n220 VPWR.n219 0.00265517
R14491 VPWR.n232 VPWR.n231 0.00265517
R14492 VPWR.n244 VPWR.n243 0.00265517
R14493 VPWR.n256 VPWR.n255 0.00265517
R14494 VPWR.n268 VPWR.n267 0.00265517
R14495 VPWR.n280 VPWR.n279 0.00265517
R14496 VPWR.n292 VPWR.n291 0.00265517
R14497 VPWR.n307 VPWR.n305 0.00265517
R14498 VPWR.n148 VPWR.n147 0.00265517
R14499 VPWR.n137 VPWR.n136 0.00265517
R14500 VPWR.n1753 VPWR.n1751 0.00265517
R14501 VPWR.n1739 VPWR.n1738 0.00265517
R14502 VPWR.n1727 VPWR.n1726 0.00265517
R14503 VPWR.n1716 VPWR.n1715 0.00265517
R14504 VPWR.n1214 VPWR.n1212 0.00265517
R14505 VPWR.n1700 VPWR.n1699 0.00265517
R14506 VPWR.n1689 VPWR.n1688 0.00265517
R14507 VPWR.n1228 VPWR.n1226 0.00265517
R14508 VPWR.n1673 VPWR.n1672 0.00265517
R14509 VPWR.n1662 VPWR.n1661 0.00265517
R14510 VPWR.n1196 VPWR.n1194 0.00265517
R14511 VPWR.n1646 VPWR.n1645 0.00265517
R14512 VPWR.n1635 VPWR.n1634 0.00265517
R14513 VPWR.n1145 VPWR.n1143 0.00265517
R14514 VPWR.n1619 VPWR.n1618 0.00265517
R14515 Iout.n1020 Iout.t100 239.927
R14516 Iout.n509 Iout.t185 239.927
R14517 Iout.n513 Iout.t41 239.927
R14518 Iout.n507 Iout.t207 239.927
R14519 Iout.n504 Iout.t246 239.927
R14520 Iout.n500 Iout.t219 239.927
R14521 Iout.n192 Iout.t75 239.927
R14522 Iout.n195 Iout.t194 239.927
R14523 Iout.n199 Iout.t118 239.927
R14524 Iout.n202 Iout.t87 239.927
R14525 Iout.n206 Iout.t144 239.927
R14526 Iout.n210 Iout.t141 239.927
R14527 Iout.n214 Iout.t26 239.927
R14528 Iout.n218 Iout.t156 239.927
R14529 Iout.n222 Iout.t67 239.927
R14530 Iout.n226 Iout.t180 239.927
R14531 Iout.n232 Iout.t132 239.927
R14532 Iout.n235 Iout.t212 239.927
R14533 Iout.n238 Iout.t7 239.927
R14534 Iout.n241 Iout.t46 239.927
R14535 Iout.n244 Iout.t44 239.927
R14536 Iout.n247 Iout.t241 239.927
R14537 Iout.n250 Iout.t22 239.927
R14538 Iout.n255 Iout.t250 239.927
R14539 Iout.n252 Iout.t114 239.927
R14540 Iout.n489 Iout.t36 239.927
R14541 Iout.n494 Iout.t51 239.927
R14542 Iout.n491 Iout.t160 239.927
R14543 Iout.n519 Iout.t24 239.927
R14544 Iout.n149 Iout.t17 239.927
R14545 Iout.n146 Iout.t170 239.927
R14546 Iout.n1010 Iout.t203 239.927
R14547 Iout.n1007 Iout.t222 239.927
R14548 Iout.n140 Iout.t80 239.927
R14549 Iout.n143 Iout.t14 239.927
R14550 Iout.n525 Iout.t96 239.927
R14551 Iout.n480 Iout.t138 239.927
R14552 Iout.n483 Iout.t153 239.927
R14553 Iout.n478 Iout.t117 239.927
R14554 Iout.n259 Iout.t223 239.927
R14555 Iout.n186 Iout.t91 239.927
R14556 Iout.n271 Iout.t225 239.927
R14557 Iout.n180 Iout.t52 239.927
R14558 Iout.n283 Iout.t127 239.927
R14559 Iout.n174 Iout.t85 239.927
R14560 Iout.n168 Iout.t166 239.927
R14561 Iout.n301 Iout.t4 239.927
R14562 Iout.n289 Iout.t116 239.927
R14563 Iout.n177 Iout.t10 239.927
R14564 Iout.n277 Iout.t174 239.927
R14565 Iout.n183 Iout.t5 239.927
R14566 Iout.n265 Iout.t188 239.927
R14567 Iout.n189 Iout.t120 239.927
R14568 Iout.n472 Iout.t106 239.927
R14569 Iout.n469 Iout.t150 239.927
R14570 Iout.n156 Iout.t205 239.927
R14571 Iout.n531 Iout.t171 239.927
R14572 Iout.n534 Iout.t217 239.927
R14573 Iout.n536 Iout.t69 239.927
R14574 Iout.n133 Iout.t218 239.927
R14575 Iout.n136 Iout.t220 239.927
R14576 Iout.n542 Iout.t226 239.927
R14577 Iout.n460 Iout.t56 239.927
R14578 Iout.n463 Iout.t79 239.927
R14579 Iout.n458 Iout.t146 239.927
R14580 Iout.n305 Iout.t216 239.927
R14581 Iout.n308 Iout.t193 239.927
R14582 Iout.n311 Iout.t25 239.927
R14583 Iout.n314 Iout.t154 239.927
R14584 Iout.n317 Iout.t143 239.927
R14585 Iout.n320 Iout.t113 239.927
R14586 Iout.n392 Iout.t237 239.927
R14587 Iout.n378 Iout.t54 239.927
R14588 Iout.n376 Iout.t72 239.927
R14589 Iout.n394 Iout.t195 239.927
R14590 Iout.n408 Iout.t11 239.927
R14591 Iout.n410 Iout.t40 239.927
R14592 Iout.n424 Iout.t88 239.927
R14593 Iout.n426 Iout.t210 239.927
R14594 Iout.n447 Iout.t176 239.927
R14595 Iout.n452 Iout.t243 239.927
R14596 Iout.n449 Iout.t129 239.927
R14597 Iout.n548 Iout.t135 239.927
R14598 Iout.n130 Iout.t236 239.927
R14599 Iout.n559 Iout.t108 239.927
R14600 Iout.n557 Iout.t209 239.927
R14601 Iout.n554 Iout.t49 239.927
R14602 Iout.n434 Iout.t18 239.927
R14603 Iout.n438 Iout.t172 239.927
R14604 Iout.n441 Iout.t68 239.927
R14605 Iout.n432 Iout.t58 239.927
R14606 Iout.n418 Iout.t162 239.927
R14607 Iout.n416 Iout.t142 239.927
R14608 Iout.n402 Iout.t23 239.927
R14609 Iout.n357 Iout.t251 239.927
R14610 Iout.n360 Iout.t82 239.927
R14611 Iout.n363 Iout.t248 239.927
R14612 Iout.n366 Iout.t70 239.927
R14613 Iout.n354 Iout.t66 239.927
R14614 Iout.n351 Iout.t90 239.927
R14615 Iout.n348 Iout.t233 239.927
R14616 Iout.n345 Iout.t214 239.927
R14617 Iout.n342 Iout.t184 239.927
R14618 Iout.n339 Iout.t151 239.927
R14619 Iout.n336 Iout.t215 239.927
R14620 Iout.n333 Iout.t136 239.927
R14621 Iout.n117 Iout.t152 239.927
R14622 Iout.n582 Iout.t224 239.927
R14623 Iout.n111 Iout.t155 239.927
R14624 Iout.n594 Iout.t164 239.927
R14625 Iout.n105 Iout.t157 239.927
R14626 Iout.n606 Iout.t86 239.927
R14627 Iout.n99 Iout.t55 239.927
R14628 Iout.n618 Iout.t98 239.927
R14629 Iout.n624 Iout.t239 239.927
R14630 Iout.n90 Iout.t95 239.927
R14631 Iout.n636 Iout.t201 239.927
R14632 Iout.n81 Iout.t131 239.927
R14633 Iout.n648 Iout.t228 239.927
R14634 Iout.n96 Iout.t94 239.927
R14635 Iout.n612 Iout.t244 239.927
R14636 Iout.n102 Iout.t33 239.927
R14637 Iout.n600 Iout.t137 239.927
R14638 Iout.n108 Iout.t145 239.927
R14639 Iout.n588 Iout.t81 239.927
R14640 Iout.n687 Iout.t59 239.927
R14641 Iout.n684 Iout.t182 239.927
R14642 Iout.n681 Iout.t140 239.927
R14643 Iout.n678 Iout.t240 239.927
R14644 Iout.n675 Iout.t247 239.927
R14645 Iout.n672 Iout.t112 239.927
R14646 Iout.n747 Iout.t1 239.927
R14647 Iout.n50 Iout.t186 239.927
R14648 Iout.n759 Iout.t77 239.927
R14649 Iout.n44 Iout.t109 239.927
R14650 Iout.n771 Iout.t38 239.927
R14651 Iout.n42 Iout.t71 239.927
R14652 Iout.n56 Iout.t229 239.927
R14653 Iout.n735 Iout.t105 239.927
R14654 Iout.n62 Iout.t211 239.927
R14655 Iout.n723 Iout.t149 239.927
R14656 Iout.n717 Iout.t202 239.927
R14657 Iout.n65 Iout.t60 239.927
R14658 Iout.n729 Iout.t192 239.927
R14659 Iout.n59 Iout.t27 239.927
R14660 Iout.n805 Iout.t31 239.927
R14661 Iout.n808 Iout.t191 239.927
R14662 Iout.n811 Iout.t208 239.927
R14663 Iout.n814 Iout.t78 239.927
R14664 Iout.n817 Iout.t231 239.927
R14665 Iout.n820 Iout.t65 239.927
R14666 Iout.n823 Iout.t74 239.927
R14667 Iout.n802 Iout.t20 239.927
R14668 Iout.n799 Iout.t199 239.927
R14669 Iout.n890 Iout.t163 239.927
R14670 Iout.n888 Iout.t102 239.927
R14671 Iout.n881 Iout.t28 239.927
R14672 Iout.n869 Iout.t133 239.927
R14673 Iout.n867 Iout.t103 239.927
R14674 Iout.n855 Iout.t125 239.927
R14675 Iout.n853 Iout.t89 239.927
R14676 Iout.n841 Iout.t249 239.927
R14677 Iout.n839 Iout.t9 239.927
R14678 Iout.n827 Iout.t227 239.927
R14679 Iout.n883 Iout.t13 239.927
R14680 Iout.n895 Iout.t245 239.927
R14681 Iout.n897 Iout.t122 239.927
R14682 Iout.n909 Iout.t99 239.927
R14683 Iout.n911 Iout.t64 239.927
R14684 Iout.n923 Iout.t121 239.927
R14685 Iout.n926 Iout.t50 239.927
R14686 Iout.n22 Iout.t139 239.927
R14687 Iout.n876 Iout.t159 239.927
R14688 Iout.n874 Iout.t128 239.927
R14689 Iout.n862 Iout.t253 239.927
R14690 Iout.n860 Iout.t12 239.927
R14691 Iout.n848 Iout.t165 239.927
R14692 Iout.n846 Iout.t130 239.927
R14693 Iout.n834 Iout.t35 239.927
R14694 Iout.n832 Iout.t196 239.927
R14695 Iout.n902 Iout.t200 239.927
R14696 Iout.n904 Iout.t57 239.927
R14697 Iout.n916 Iout.t221 239.927
R14698 Iout.n918 Iout.t148 239.927
R14699 Iout.n931 Iout.t2 239.927
R14700 Iout.n934 Iout.t0 239.927
R14701 Iout.n796 Iout.t115 239.927
R14702 Iout.n793 Iout.t235 239.927
R14703 Iout.n790 Iout.t178 239.927
R14704 Iout.n787 Iout.t147 239.927
R14705 Iout.n784 Iout.t104 239.927
R14706 Iout.n781 Iout.t83 239.927
R14707 Iout.n938 Iout.t169 239.927
R14708 Iout.n741 Iout.t101 239.927
R14709 Iout.n53 Iout.t187 239.927
R14710 Iout.n753 Iout.t3 239.927
R14711 Iout.n47 Iout.t92 239.927
R14712 Iout.n765 Iout.t254 239.927
R14713 Iout.n38 Iout.t30 239.927
R14714 Iout.n777 Iout.t42 239.927
R14715 Iout.n71 Iout.t111 239.927
R14716 Iout.n705 Iout.t234 239.927
R14717 Iout.n77 Iout.t190 239.927
R14718 Iout.n944 Iout.t179 239.927
R14719 Iout.n19 Iout.t16 239.927
R14720 Iout.n68 Iout.t43 239.927
R14721 Iout.n711 Iout.t158 239.927
R14722 Iout.n74 Iout.t76 239.927
R14723 Iout.n699 Iout.t232 239.927
R14724 Iout.n950 Iout.t110 239.927
R14725 Iout.n953 Iout.t32 239.927
R14726 Iout.n669 Iout.t37 239.927
R14727 Iout.n666 Iout.t84 239.927
R14728 Iout.n663 Iout.t126 239.927
R14729 Iout.n660 Iout.t206 239.927
R14730 Iout.n657 Iout.t8 239.927
R14731 Iout.n654 Iout.t134 239.927
R14732 Iout.n690 Iout.t19 239.927
R14733 Iout.n695 Iout.t34 239.927
R14734 Iout.n692 Iout.t198 239.927
R14735 Iout.n957 Iout.t93 239.927
R14736 Iout.n114 Iout.t168 239.927
R14737 Iout.n576 Iout.t197 239.927
R14738 Iout.n573 Iout.t15 239.927
R14739 Iout.n963 Iout.t39 239.927
R14740 Iout.n14 Iout.t183 239.927
R14741 Iout.n93 Iout.t29 239.927
R14742 Iout.n630 Iout.t6 239.927
R14743 Iout.n87 Iout.t21 239.927
R14744 Iout.n642 Iout.t73 239.927
R14745 Iout.n85 Iout.t177 239.927
R14746 Iout.n563 Iout.t48 239.927
R14747 Iout.n969 Iout.t124 239.927
R14748 Iout.n972 Iout.t63 239.927
R14749 Iout.n569 Iout.t255 239.927
R14750 Iout.n123 Iout.t161 239.927
R14751 Iout.n120 Iout.t189 239.927
R14752 Iout.n976 Iout.t204 239.927
R14753 Iout.n400 Iout.t181 239.927
R14754 Iout.n386 Iout.t61 239.927
R14755 Iout.n384 Iout.t175 239.927
R14756 Iout.n370 Iout.t62 239.927
R14757 Iout.n982 Iout.t45 239.927
R14758 Iout.n9 Iout.t238 239.927
R14759 Iout.n127 Iout.t173 239.927
R14760 Iout.n988 Iout.t107 239.927
R14761 Iout.n991 Iout.t167 239.927
R14762 Iout.n323 Iout.t213 239.927
R14763 Iout.n326 Iout.t230 239.927
R14764 Iout.n329 Iout.t47 239.927
R14765 Iout.n995 Iout.t242 239.927
R14766 Iout.n1001 Iout.t123 239.927
R14767 Iout.n4 Iout.t119 239.927
R14768 Iout.n295 Iout.t252 239.927
R14769 Iout.n172 Iout.t53 239.927
R14770 Iout.n1014 Iout.t97 239.927
R14771 Iout.n1021 Iout.n1020 7.9105
R14772 Iout.n510 Iout.n509 7.9105
R14773 Iout.n514 Iout.n513 7.9105
R14774 Iout.n508 Iout.n507 7.9105
R14775 Iout.n505 Iout.n504 7.9105
R14776 Iout.n501 Iout.n500 7.9105
R14777 Iout.n193 Iout.n192 7.9105
R14778 Iout.n196 Iout.n195 7.9105
R14779 Iout.n200 Iout.n199 7.9105
R14780 Iout.n203 Iout.n202 7.9105
R14781 Iout.n207 Iout.n206 7.9105
R14782 Iout.n211 Iout.n210 7.9105
R14783 Iout.n215 Iout.n214 7.9105
R14784 Iout.n219 Iout.n218 7.9105
R14785 Iout.n223 Iout.n222 7.9105
R14786 Iout.n227 Iout.n226 7.9105
R14787 Iout.n233 Iout.n232 7.9105
R14788 Iout.n236 Iout.n235 7.9105
R14789 Iout.n239 Iout.n238 7.9105
R14790 Iout.n242 Iout.n241 7.9105
R14791 Iout.n245 Iout.n244 7.9105
R14792 Iout.n248 Iout.n247 7.9105
R14793 Iout.n251 Iout.n250 7.9105
R14794 Iout.n256 Iout.n255 7.9105
R14795 Iout.n253 Iout.n252 7.9105
R14796 Iout.n490 Iout.n489 7.9105
R14797 Iout.n495 Iout.n494 7.9105
R14798 Iout.n492 Iout.n491 7.9105
R14799 Iout.n520 Iout.n519 7.9105
R14800 Iout.n150 Iout.n149 7.9105
R14801 Iout.n147 Iout.n146 7.9105
R14802 Iout.n1011 Iout.n1010 7.9105
R14803 Iout.n1008 Iout.n1007 7.9105
R14804 Iout.n141 Iout.n140 7.9105
R14805 Iout.n144 Iout.n143 7.9105
R14806 Iout.n526 Iout.n525 7.9105
R14807 Iout.n481 Iout.n480 7.9105
R14808 Iout.n484 Iout.n483 7.9105
R14809 Iout.n479 Iout.n478 7.9105
R14810 Iout.n260 Iout.n259 7.9105
R14811 Iout.n187 Iout.n186 7.9105
R14812 Iout.n272 Iout.n271 7.9105
R14813 Iout.n181 Iout.n180 7.9105
R14814 Iout.n284 Iout.n283 7.9105
R14815 Iout.n175 Iout.n174 7.9105
R14816 Iout.n169 Iout.n168 7.9105
R14817 Iout.n302 Iout.n301 7.9105
R14818 Iout.n290 Iout.n289 7.9105
R14819 Iout.n178 Iout.n177 7.9105
R14820 Iout.n278 Iout.n277 7.9105
R14821 Iout.n184 Iout.n183 7.9105
R14822 Iout.n266 Iout.n265 7.9105
R14823 Iout.n190 Iout.n189 7.9105
R14824 Iout.n473 Iout.n472 7.9105
R14825 Iout.n470 Iout.n469 7.9105
R14826 Iout.n157 Iout.n156 7.9105
R14827 Iout.n532 Iout.n531 7.9105
R14828 Iout.n535 Iout.n534 7.9105
R14829 Iout.n537 Iout.n536 7.9105
R14830 Iout.n134 Iout.n133 7.9105
R14831 Iout.n137 Iout.n136 7.9105
R14832 Iout.n543 Iout.n542 7.9105
R14833 Iout.n461 Iout.n460 7.9105
R14834 Iout.n464 Iout.n463 7.9105
R14835 Iout.n459 Iout.n458 7.9105
R14836 Iout.n306 Iout.n305 7.9105
R14837 Iout.n309 Iout.n308 7.9105
R14838 Iout.n312 Iout.n311 7.9105
R14839 Iout.n315 Iout.n314 7.9105
R14840 Iout.n318 Iout.n317 7.9105
R14841 Iout.n321 Iout.n320 7.9105
R14842 Iout.n393 Iout.n392 7.9105
R14843 Iout.n379 Iout.n378 7.9105
R14844 Iout.n377 Iout.n376 7.9105
R14845 Iout.n395 Iout.n394 7.9105
R14846 Iout.n409 Iout.n408 7.9105
R14847 Iout.n411 Iout.n410 7.9105
R14848 Iout.n425 Iout.n424 7.9105
R14849 Iout.n427 Iout.n426 7.9105
R14850 Iout.n448 Iout.n447 7.9105
R14851 Iout.n453 Iout.n452 7.9105
R14852 Iout.n450 Iout.n449 7.9105
R14853 Iout.n549 Iout.n548 7.9105
R14854 Iout.n131 Iout.n130 7.9105
R14855 Iout.n560 Iout.n559 7.9105
R14856 Iout.n558 Iout.n557 7.9105
R14857 Iout.n555 Iout.n554 7.9105
R14858 Iout.n435 Iout.n434 7.9105
R14859 Iout.n439 Iout.n438 7.9105
R14860 Iout.n442 Iout.n441 7.9105
R14861 Iout.n433 Iout.n432 7.9105
R14862 Iout.n419 Iout.n418 7.9105
R14863 Iout.n417 Iout.n416 7.9105
R14864 Iout.n403 Iout.n402 7.9105
R14865 Iout.n358 Iout.n357 7.9105
R14866 Iout.n361 Iout.n360 7.9105
R14867 Iout.n364 Iout.n363 7.9105
R14868 Iout.n367 Iout.n366 7.9105
R14869 Iout.n355 Iout.n354 7.9105
R14870 Iout.n352 Iout.n351 7.9105
R14871 Iout.n349 Iout.n348 7.9105
R14872 Iout.n346 Iout.n345 7.9105
R14873 Iout.n343 Iout.n342 7.9105
R14874 Iout.n340 Iout.n339 7.9105
R14875 Iout.n337 Iout.n336 7.9105
R14876 Iout.n334 Iout.n333 7.9105
R14877 Iout.n118 Iout.n117 7.9105
R14878 Iout.n583 Iout.n582 7.9105
R14879 Iout.n112 Iout.n111 7.9105
R14880 Iout.n595 Iout.n594 7.9105
R14881 Iout.n106 Iout.n105 7.9105
R14882 Iout.n607 Iout.n606 7.9105
R14883 Iout.n100 Iout.n99 7.9105
R14884 Iout.n619 Iout.n618 7.9105
R14885 Iout.n625 Iout.n624 7.9105
R14886 Iout.n91 Iout.n90 7.9105
R14887 Iout.n637 Iout.n636 7.9105
R14888 Iout.n82 Iout.n81 7.9105
R14889 Iout.n649 Iout.n648 7.9105
R14890 Iout.n97 Iout.n96 7.9105
R14891 Iout.n613 Iout.n612 7.9105
R14892 Iout.n103 Iout.n102 7.9105
R14893 Iout.n601 Iout.n600 7.9105
R14894 Iout.n109 Iout.n108 7.9105
R14895 Iout.n589 Iout.n588 7.9105
R14896 Iout.n688 Iout.n687 7.9105
R14897 Iout.n685 Iout.n684 7.9105
R14898 Iout.n682 Iout.n681 7.9105
R14899 Iout.n679 Iout.n678 7.9105
R14900 Iout.n676 Iout.n675 7.9105
R14901 Iout.n673 Iout.n672 7.9105
R14902 Iout.n748 Iout.n747 7.9105
R14903 Iout.n51 Iout.n50 7.9105
R14904 Iout.n760 Iout.n759 7.9105
R14905 Iout.n45 Iout.n44 7.9105
R14906 Iout.n772 Iout.n771 7.9105
R14907 Iout.n43 Iout.n42 7.9105
R14908 Iout.n57 Iout.n56 7.9105
R14909 Iout.n736 Iout.n735 7.9105
R14910 Iout.n63 Iout.n62 7.9105
R14911 Iout.n724 Iout.n723 7.9105
R14912 Iout.n718 Iout.n717 7.9105
R14913 Iout.n66 Iout.n65 7.9105
R14914 Iout.n730 Iout.n729 7.9105
R14915 Iout.n60 Iout.n59 7.9105
R14916 Iout.n806 Iout.n805 7.9105
R14917 Iout.n809 Iout.n808 7.9105
R14918 Iout.n812 Iout.n811 7.9105
R14919 Iout.n815 Iout.n814 7.9105
R14920 Iout.n818 Iout.n817 7.9105
R14921 Iout.n821 Iout.n820 7.9105
R14922 Iout.n824 Iout.n823 7.9105
R14923 Iout.n803 Iout.n802 7.9105
R14924 Iout.n800 Iout.n799 7.9105
R14925 Iout.n891 Iout.n890 7.9105
R14926 Iout.n889 Iout.n888 7.9105
R14927 Iout.n882 Iout.n881 7.9105
R14928 Iout.n870 Iout.n869 7.9105
R14929 Iout.n868 Iout.n867 7.9105
R14930 Iout.n856 Iout.n855 7.9105
R14931 Iout.n854 Iout.n853 7.9105
R14932 Iout.n842 Iout.n841 7.9105
R14933 Iout.n840 Iout.n839 7.9105
R14934 Iout.n828 Iout.n827 7.9105
R14935 Iout.n884 Iout.n883 7.9105
R14936 Iout.n896 Iout.n895 7.9105
R14937 Iout.n898 Iout.n897 7.9105
R14938 Iout.n910 Iout.n909 7.9105
R14939 Iout.n912 Iout.n911 7.9105
R14940 Iout.n924 Iout.n923 7.9105
R14941 Iout.n927 Iout.n926 7.9105
R14942 Iout.n23 Iout.n22 7.9105
R14943 Iout.n877 Iout.n876 7.9105
R14944 Iout.n875 Iout.n874 7.9105
R14945 Iout.n863 Iout.n862 7.9105
R14946 Iout.n861 Iout.n860 7.9105
R14947 Iout.n849 Iout.n848 7.9105
R14948 Iout.n847 Iout.n846 7.9105
R14949 Iout.n835 Iout.n834 7.9105
R14950 Iout.n833 Iout.n832 7.9105
R14951 Iout.n903 Iout.n902 7.9105
R14952 Iout.n905 Iout.n904 7.9105
R14953 Iout.n917 Iout.n916 7.9105
R14954 Iout.n919 Iout.n918 7.9105
R14955 Iout.n932 Iout.n931 7.9105
R14956 Iout.n935 Iout.n934 7.9105
R14957 Iout.n797 Iout.n796 7.9105
R14958 Iout.n794 Iout.n793 7.9105
R14959 Iout.n791 Iout.n790 7.9105
R14960 Iout.n788 Iout.n787 7.9105
R14961 Iout.n785 Iout.n784 7.9105
R14962 Iout.n782 Iout.n781 7.9105
R14963 Iout.n939 Iout.n938 7.9105
R14964 Iout.n742 Iout.n741 7.9105
R14965 Iout.n54 Iout.n53 7.9105
R14966 Iout.n754 Iout.n753 7.9105
R14967 Iout.n48 Iout.n47 7.9105
R14968 Iout.n766 Iout.n765 7.9105
R14969 Iout.n39 Iout.n38 7.9105
R14970 Iout.n778 Iout.n777 7.9105
R14971 Iout.n72 Iout.n71 7.9105
R14972 Iout.n706 Iout.n705 7.9105
R14973 Iout.n78 Iout.n77 7.9105
R14974 Iout.n945 Iout.n944 7.9105
R14975 Iout.n20 Iout.n19 7.9105
R14976 Iout.n69 Iout.n68 7.9105
R14977 Iout.n712 Iout.n711 7.9105
R14978 Iout.n75 Iout.n74 7.9105
R14979 Iout.n700 Iout.n699 7.9105
R14980 Iout.n951 Iout.n950 7.9105
R14981 Iout.n954 Iout.n953 7.9105
R14982 Iout.n670 Iout.n669 7.9105
R14983 Iout.n667 Iout.n666 7.9105
R14984 Iout.n664 Iout.n663 7.9105
R14985 Iout.n661 Iout.n660 7.9105
R14986 Iout.n658 Iout.n657 7.9105
R14987 Iout.n655 Iout.n654 7.9105
R14988 Iout.n691 Iout.n690 7.9105
R14989 Iout.n696 Iout.n695 7.9105
R14990 Iout.n693 Iout.n692 7.9105
R14991 Iout.n958 Iout.n957 7.9105
R14992 Iout.n115 Iout.n114 7.9105
R14993 Iout.n577 Iout.n576 7.9105
R14994 Iout.n574 Iout.n573 7.9105
R14995 Iout.n964 Iout.n963 7.9105
R14996 Iout.n15 Iout.n14 7.9105
R14997 Iout.n94 Iout.n93 7.9105
R14998 Iout.n631 Iout.n630 7.9105
R14999 Iout.n88 Iout.n87 7.9105
R15000 Iout.n643 Iout.n642 7.9105
R15001 Iout.n86 Iout.n85 7.9105
R15002 Iout.n564 Iout.n563 7.9105
R15003 Iout.n970 Iout.n969 7.9105
R15004 Iout.n973 Iout.n972 7.9105
R15005 Iout.n570 Iout.n569 7.9105
R15006 Iout.n124 Iout.n123 7.9105
R15007 Iout.n121 Iout.n120 7.9105
R15008 Iout.n977 Iout.n976 7.9105
R15009 Iout.n401 Iout.n400 7.9105
R15010 Iout.n387 Iout.n386 7.9105
R15011 Iout.n385 Iout.n384 7.9105
R15012 Iout.n371 Iout.n370 7.9105
R15013 Iout.n983 Iout.n982 7.9105
R15014 Iout.n10 Iout.n9 7.9105
R15015 Iout.n128 Iout.n127 7.9105
R15016 Iout.n989 Iout.n988 7.9105
R15017 Iout.n992 Iout.n991 7.9105
R15018 Iout.n324 Iout.n323 7.9105
R15019 Iout.n327 Iout.n326 7.9105
R15020 Iout.n330 Iout.n329 7.9105
R15021 Iout.n996 Iout.n995 7.9105
R15022 Iout.n1002 Iout.n1001 7.9105
R15023 Iout.n5 Iout.n4 7.9105
R15024 Iout.n296 Iout.n295 7.9105
R15025 Iout.n173 Iout.n172 7.9105
R15026 Iout.n1015 Iout.n1014 7.9105
R15027 Iout.n886 Iout.n885 3.86101
R15028 Iout.n880 Iout.n879 3.86101
R15029 Iout.n894 Iout.n893 3.86101
R15030 Iout.n872 Iout.n871 3.86101
R15031 Iout.n900 Iout.n899 3.86101
R15032 Iout.n866 Iout.n865 3.86101
R15033 Iout.n908 Iout.n907 3.86101
R15034 Iout.n858 Iout.n857 3.86101
R15035 Iout.n914 Iout.n913 3.86101
R15036 Iout.n852 Iout.n851 3.86101
R15037 Iout.n922 Iout.n921 3.86101
R15038 Iout.n844 Iout.n843 3.86101
R15039 Iout.n929 Iout.n928 3.86101
R15040 Iout.n838 Iout.n837 3.86101
R15041 Iout.n925 Iout.n21 3.86101
R15042 Iout.n830 Iout.n829 3.86101
R15043 Iout.n879 Iout.n878 3.4105
R15044 Iout.n887 Iout.n886 3.4105
R15045 Iout.n893 Iout.n892 3.4105
R15046 Iout.n798 Iout.n28 3.4105
R15047 Iout.n801 Iout.n29 3.4105
R15048 Iout.n804 Iout.n30 3.4105
R15049 Iout.n807 Iout.n31 3.4105
R15050 Iout.n873 Iout.n872 3.4105
R15051 Iout.n744 Iout.n743 3.4105
R15052 Iout.n740 Iout.n739 3.4105
R15053 Iout.n732 Iout.n731 3.4105
R15054 Iout.n728 Iout.n727 3.4105
R15055 Iout.n720 Iout.n719 3.4105
R15056 Iout.n795 Iout.n27 3.4105
R15057 Iout.n901 Iout.n900 3.4105
R15058 Iout.n722 Iout.n721 3.4105
R15059 Iout.n726 Iout.n725 3.4105
R15060 Iout.n734 Iout.n733 3.4105
R15061 Iout.n738 Iout.n737 3.4105
R15062 Iout.n746 Iout.n745 3.4105
R15063 Iout.n750 Iout.n749 3.4105
R15064 Iout.n752 Iout.n751 3.4105
R15065 Iout.n810 Iout.n32 3.4105
R15066 Iout.n865 Iout.n864 3.4105
R15067 Iout.n668 Iout.n55 3.4105
R15068 Iout.n671 Iout.n58 3.4105
R15069 Iout.n674 Iout.n61 3.4105
R15070 Iout.n677 Iout.n64 3.4105
R15071 Iout.n680 Iout.n67 3.4105
R15072 Iout.n683 Iout.n70 3.4105
R15073 Iout.n686 Iout.n73 3.4105
R15074 Iout.n714 Iout.n713 3.4105
R15075 Iout.n716 Iout.n715 3.4105
R15076 Iout.n792 Iout.n26 3.4105
R15077 Iout.n907 Iout.n906 3.4105
R15078 Iout.n587 Iout.n586 3.4105
R15079 Iout.n591 Iout.n590 3.4105
R15080 Iout.n599 Iout.n598 3.4105
R15081 Iout.n603 Iout.n602 3.4105
R15082 Iout.n611 Iout.n610 3.4105
R15083 Iout.n615 Iout.n614 3.4105
R15084 Iout.n623 Iout.n622 3.4105
R15085 Iout.n627 Iout.n626 3.4105
R15086 Iout.n665 Iout.n52 3.4105
R15087 Iout.n758 Iout.n757 3.4105
R15088 Iout.n756 Iout.n755 3.4105
R15089 Iout.n813 Iout.n33 3.4105
R15090 Iout.n859 Iout.n858 3.4105
R15091 Iout.n629 Iout.n628 3.4105
R15092 Iout.n621 Iout.n620 3.4105
R15093 Iout.n617 Iout.n616 3.4105
R15094 Iout.n609 Iout.n608 3.4105
R15095 Iout.n605 Iout.n604 3.4105
R15096 Iout.n597 Iout.n596 3.4105
R15097 Iout.n593 Iout.n592 3.4105
R15098 Iout.n585 Iout.n584 3.4105
R15099 Iout.n581 Iout.n580 3.4105
R15100 Iout.n579 Iout.n578 3.4105
R15101 Iout.n689 Iout.n76 3.4105
R15102 Iout.n710 Iout.n709 3.4105
R15103 Iout.n708 Iout.n707 3.4105
R15104 Iout.n789 Iout.n25 3.4105
R15105 Iout.n915 Iout.n914 3.4105
R15106 Iout.n572 Iout.n571 3.4105
R15107 Iout.n335 Iout.n116 3.4105
R15108 Iout.n338 Iout.n113 3.4105
R15109 Iout.n341 Iout.n110 3.4105
R15110 Iout.n344 Iout.n107 3.4105
R15111 Iout.n347 Iout.n104 3.4105
R15112 Iout.n350 Iout.n101 3.4105
R15113 Iout.n353 Iout.n98 3.4105
R15114 Iout.n356 Iout.n95 3.4105
R15115 Iout.n359 Iout.n92 3.4105
R15116 Iout.n633 Iout.n632 3.4105
R15117 Iout.n635 Iout.n634 3.4105
R15118 Iout.n662 Iout.n49 3.4105
R15119 Iout.n762 Iout.n761 3.4105
R15120 Iout.n764 Iout.n763 3.4105
R15121 Iout.n816 Iout.n34 3.4105
R15122 Iout.n851 Iout.n850 3.4105
R15123 Iout.n399 Iout.n398 3.4105
R15124 Iout.n405 Iout.n404 3.4105
R15125 Iout.n415 Iout.n414 3.4105
R15126 Iout.n421 Iout.n420 3.4105
R15127 Iout.n431 Iout.n430 3.4105
R15128 Iout.n444 Iout.n443 3.4105
R15129 Iout.n440 Iout.n159 3.4105
R15130 Iout.n437 Iout.n436 3.4105
R15131 Iout.n553 Iout.n552 3.4105
R15132 Iout.n556 Iout.n119 3.4105
R15133 Iout.n562 Iout.n561 3.4105
R15134 Iout.n568 Iout.n567 3.4105
R15135 Iout.n566 Iout.n565 3.4105
R15136 Iout.n575 Iout.n79 3.4105
R15137 Iout.n698 Iout.n697 3.4105
R15138 Iout.n702 Iout.n701 3.4105
R15139 Iout.n704 Iout.n703 3.4105
R15140 Iout.n786 Iout.n24 3.4105
R15141 Iout.n921 Iout.n920 3.4105
R15142 Iout.n129 Iout.n125 3.4105
R15143 Iout.n547 Iout.n546 3.4105
R15144 Iout.n551 Iout.n550 3.4105
R15145 Iout.n451 Iout.n158 3.4105
R15146 Iout.n455 Iout.n454 3.4105
R15147 Iout.n446 Iout.n445 3.4105
R15148 Iout.n429 Iout.n428 3.4105
R15149 Iout.n423 Iout.n422 3.4105
R15150 Iout.n413 Iout.n412 3.4105
R15151 Iout.n407 Iout.n406 3.4105
R15152 Iout.n397 Iout.n396 3.4105
R15153 Iout.n391 Iout.n390 3.4105
R15154 Iout.n389 Iout.n388 3.4105
R15155 Iout.n362 Iout.n89 3.4105
R15156 Iout.n641 Iout.n640 3.4105
R15157 Iout.n639 Iout.n638 3.4105
R15158 Iout.n659 Iout.n46 3.4105
R15159 Iout.n770 Iout.n769 3.4105
R15160 Iout.n768 Iout.n767 3.4105
R15161 Iout.n819 Iout.n35 3.4105
R15162 Iout.n845 Iout.n844 3.4105
R15163 Iout.n325 Iout.n165 3.4105
R15164 Iout.n322 Iout.n164 3.4105
R15165 Iout.n319 Iout.n163 3.4105
R15166 Iout.n316 Iout.n162 3.4105
R15167 Iout.n313 Iout.n161 3.4105
R15168 Iout.n310 Iout.n160 3.4105
R15169 Iout.n307 Iout.n155 3.4105
R15170 Iout.n457 Iout.n456 3.4105
R15171 Iout.n466 Iout.n465 3.4105
R15172 Iout.n462 Iout.n126 3.4105
R15173 Iout.n545 Iout.n544 3.4105
R15174 Iout.n541 Iout.n540 3.4105
R15175 Iout.n135 Iout.n3 3.4105
R15176 Iout.n987 Iout.n986 3.4105
R15177 Iout.n985 Iout.n984 3.4105
R15178 Iout.n122 Iout.n8 3.4105
R15179 Iout.n968 Iout.n967 3.4105
R15180 Iout.n966 Iout.n965 3.4105
R15181 Iout.n694 Iout.n13 3.4105
R15182 Iout.n949 Iout.n948 3.4105
R15183 Iout.n947 Iout.n946 3.4105
R15184 Iout.n783 Iout.n18 3.4105
R15185 Iout.n930 Iout.n929 3.4105
R15186 Iout.n1004 Iout.n1003 3.4105
R15187 Iout.n539 Iout.n538 3.4105
R15188 Iout.n533 Iout.n132 3.4105
R15189 Iout.n530 Iout.n529 3.4105
R15190 Iout.n468 Iout.n467 3.4105
R15191 Iout.n471 Iout.n153 3.4105
R15192 Iout.n475 Iout.n474 3.4105
R15193 Iout.n264 Iout.n263 3.4105
R15194 Iout.n268 Iout.n267 3.4105
R15195 Iout.n276 Iout.n275 3.4105
R15196 Iout.n280 Iout.n279 3.4105
R15197 Iout.n288 Iout.n287 3.4105
R15198 Iout.n292 Iout.n291 3.4105
R15199 Iout.n300 Iout.n299 3.4105
R15200 Iout.n328 Iout.n166 3.4105
R15201 Iout.n381 Iout.n380 3.4105
R15202 Iout.n383 Iout.n382 3.4105
R15203 Iout.n365 Iout.n83 3.4105
R15204 Iout.n645 Iout.n644 3.4105
R15205 Iout.n647 Iout.n646 3.4105
R15206 Iout.n656 Iout.n40 3.4105
R15207 Iout.n774 Iout.n773 3.4105
R15208 Iout.n776 Iout.n775 3.4105
R15209 Iout.n822 Iout.n36 3.4105
R15210 Iout.n837 Iout.n836 3.4105
R15211 Iout.n298 Iout.n297 3.4105
R15212 Iout.n294 Iout.n293 3.4105
R15213 Iout.n286 Iout.n285 3.4105
R15214 Iout.n282 Iout.n281 3.4105
R15215 Iout.n274 Iout.n273 3.4105
R15216 Iout.n270 Iout.n269 3.4105
R15217 Iout.n262 Iout.n261 3.4105
R15218 Iout.n477 Iout.n476 3.4105
R15219 Iout.n486 Iout.n485 3.4105
R15220 Iout.n482 Iout.n151 3.4105
R15221 Iout.n528 Iout.n527 3.4105
R15222 Iout.n524 Iout.n523 3.4105
R15223 Iout.n142 Iout.n138 3.4105
R15224 Iout.n1006 Iout.n1005 3.4105
R15225 Iout.n1009 Iout.n0 3.4105
R15226 Iout.n1000 Iout.n999 3.4105
R15227 Iout.n998 Iout.n997 3.4105
R15228 Iout.n990 Iout.n6 3.4105
R15229 Iout.n981 Iout.n980 3.4105
R15230 Iout.n979 Iout.n978 3.4105
R15231 Iout.n971 Iout.n11 3.4105
R15232 Iout.n962 Iout.n961 3.4105
R15233 Iout.n960 Iout.n959 3.4105
R15234 Iout.n952 Iout.n16 3.4105
R15235 Iout.n943 Iout.n942 3.4105
R15236 Iout.n941 Iout.n940 3.4105
R15237 Iout.n933 Iout.n21 3.4105
R15238 Iout.n1017 Iout.n1016 3.4105
R15239 Iout.n148 Iout.n2 3.4105
R15240 Iout.n518 Iout.n517 3.4105
R15241 Iout.n522 Iout.n521 3.4105
R15242 Iout.n493 Iout.n139 3.4105
R15243 Iout.n497 Iout.n496 3.4105
R15244 Iout.n488 Iout.n487 3.4105
R15245 Iout.n254 Iout.n154 3.4105
R15246 Iout.n258 Iout.n257 3.4105
R15247 Iout.n249 Iout.n188 3.4105
R15248 Iout.n246 Iout.n185 3.4105
R15249 Iout.n243 Iout.n182 3.4105
R15250 Iout.n240 Iout.n179 3.4105
R15251 Iout.n237 Iout.n176 3.4105
R15252 Iout.n234 Iout.n170 3.4105
R15253 Iout.n231 Iout.n230 3.4105
R15254 Iout.n171 Iout.n167 3.4105
R15255 Iout.n304 Iout.n303 3.4105
R15256 Iout.n332 Iout.n331 3.4105
R15257 Iout.n375 Iout.n374 3.4105
R15258 Iout.n373 Iout.n372 3.4105
R15259 Iout.n369 Iout.n368 3.4105
R15260 Iout.n84 Iout.n80 3.4105
R15261 Iout.n651 Iout.n650 3.4105
R15262 Iout.n653 Iout.n652 3.4105
R15263 Iout.n41 Iout.n37 3.4105
R15264 Iout.n780 Iout.n779 3.4105
R15265 Iout.n826 Iout.n825 3.4105
R15266 Iout.n831 Iout.n830 3.4105
R15267 Iout.n229 Iout.n228 3.4105
R15268 Iout.n225 Iout.n224 3.4105
R15269 Iout.n221 Iout.n220 3.4105
R15270 Iout.n217 Iout.n216 3.4105
R15271 Iout.n213 Iout.n212 3.4105
R15272 Iout.n209 Iout.n208 3.4105
R15273 Iout.n205 Iout.n204 3.4105
R15274 Iout.n201 Iout.n191 3.4105
R15275 Iout.n198 Iout.n197 3.4105
R15276 Iout.n194 Iout.n152 3.4105
R15277 Iout.n499 Iout.n498 3.4105
R15278 Iout.n503 Iout.n502 3.4105
R15279 Iout.n506 Iout.n145 3.4105
R15280 Iout.n516 Iout.n515 3.4105
R15281 Iout.n512 Iout.n511 3.4105
R15282 Iout.n1019 Iout.n1018 3.4105
R15283 Iout.n936 Iout.n23 1.43848
R15284 Iout.n936 Iout.n935 1.34612
R15285 Iout.n939 Iout.n937 1.34612
R15286 Iout.n20 Iout.n17 1.34612
R15287 Iout.n955 Iout.n954 1.34612
R15288 Iout.n958 Iout.n956 1.34612
R15289 Iout.n15 Iout.n12 1.34612
R15290 Iout.n974 Iout.n973 1.34612
R15291 Iout.n977 Iout.n975 1.34612
R15292 Iout.n10 Iout.n7 1.34612
R15293 Iout.n993 Iout.n992 1.34612
R15294 Iout.n996 Iout.n994 1.34612
R15295 Iout.n5 Iout.n1 1.34612
R15296 Iout.n1012 Iout.n1011 1.34612
R15297 Iout.n1015 Iout.n1013 1.34612
R15298 Iout.n1022 Iout.n1021 1.34612
R15299 Iout.n197 Iout.n154 0.451012
R15300 Iout.n476 Iout.n154 0.451012
R15301 Iout.n476 Iout.n475 0.451012
R15302 Iout.n475 Iout.n155 0.451012
R15303 Iout.n445 Iout.n155 0.451012
R15304 Iout.n445 Iout.n444 0.451012
R15305 Iout.n444 Iout.n107 0.451012
R15306 Iout.n604 Iout.n107 0.451012
R15307 Iout.n604 Iout.n603 0.451012
R15308 Iout.n603 Iout.n64 0.451012
R15309 Iout.n733 Iout.n64 0.451012
R15310 Iout.n733 Iout.n732 0.451012
R15311 Iout.n732 Iout.n29 0.451012
R15312 Iout.n886 Iout.n29 0.451012
R15313 Iout.n258 Iout.n191 0.451012
R15314 Iout.n262 Iout.n258 0.451012
R15315 Iout.n263 Iout.n262 0.451012
R15316 Iout.n263 Iout.n160 0.451012
R15317 Iout.n429 Iout.n160 0.451012
R15318 Iout.n430 Iout.n429 0.451012
R15319 Iout.n430 Iout.n104 0.451012
R15320 Iout.n609 Iout.n104 0.451012
R15321 Iout.n610 Iout.n609 0.451012
R15322 Iout.n610 Iout.n61 0.451012
R15323 Iout.n738 Iout.n61 0.451012
R15324 Iout.n739 Iout.n738 0.451012
R15325 Iout.n739 Iout.n30 0.451012
R15326 Iout.n879 Iout.n30 0.451012
R15327 Iout.n487 Iout.n152 0.451012
R15328 Iout.n487 Iout.n486 0.451012
R15329 Iout.n486 Iout.n153 0.451012
R15330 Iout.n456 Iout.n153 0.451012
R15331 Iout.n456 Iout.n455 0.451012
R15332 Iout.n455 Iout.n159 0.451012
R15333 Iout.n159 Iout.n110 0.451012
R15334 Iout.n597 Iout.n110 0.451012
R15335 Iout.n598 Iout.n597 0.451012
R15336 Iout.n598 Iout.n67 0.451012
R15337 Iout.n726 Iout.n67 0.451012
R15338 Iout.n727 Iout.n726 0.451012
R15339 Iout.n727 Iout.n28 0.451012
R15340 Iout.n893 Iout.n28 0.451012
R15341 Iout.n204 Iout.n188 0.451012
R15342 Iout.n269 Iout.n188 0.451012
R15343 Iout.n269 Iout.n268 0.451012
R15344 Iout.n268 Iout.n161 0.451012
R15345 Iout.n422 Iout.n161 0.451012
R15346 Iout.n422 Iout.n421 0.451012
R15347 Iout.n421 Iout.n101 0.451012
R15348 Iout.n616 Iout.n101 0.451012
R15349 Iout.n616 Iout.n615 0.451012
R15350 Iout.n615 Iout.n58 0.451012
R15351 Iout.n745 Iout.n58 0.451012
R15352 Iout.n745 Iout.n744 0.451012
R15353 Iout.n744 Iout.n31 0.451012
R15354 Iout.n872 Iout.n31 0.451012
R15355 Iout.n498 Iout.n497 0.451012
R15356 Iout.n497 Iout.n151 0.451012
R15357 Iout.n467 Iout.n151 0.451012
R15358 Iout.n467 Iout.n466 0.451012
R15359 Iout.n466 Iout.n158 0.451012
R15360 Iout.n436 Iout.n158 0.451012
R15361 Iout.n436 Iout.n113 0.451012
R15362 Iout.n592 Iout.n113 0.451012
R15363 Iout.n592 Iout.n591 0.451012
R15364 Iout.n591 Iout.n70 0.451012
R15365 Iout.n721 Iout.n70 0.451012
R15366 Iout.n721 Iout.n720 0.451012
R15367 Iout.n720 Iout.n27 0.451012
R15368 Iout.n900 Iout.n27 0.451012
R15369 Iout.n208 Iout.n185 0.451012
R15370 Iout.n274 Iout.n185 0.451012
R15371 Iout.n275 Iout.n274 0.451012
R15372 Iout.n275 Iout.n162 0.451012
R15373 Iout.n413 Iout.n162 0.451012
R15374 Iout.n414 Iout.n413 0.451012
R15375 Iout.n414 Iout.n98 0.451012
R15376 Iout.n621 Iout.n98 0.451012
R15377 Iout.n622 Iout.n621 0.451012
R15378 Iout.n622 Iout.n55 0.451012
R15379 Iout.n750 Iout.n55 0.451012
R15380 Iout.n751 Iout.n750 0.451012
R15381 Iout.n751 Iout.n32 0.451012
R15382 Iout.n865 Iout.n32 0.451012
R15383 Iout.n502 Iout.n139 0.451012
R15384 Iout.n528 Iout.n139 0.451012
R15385 Iout.n529 Iout.n528 0.451012
R15386 Iout.n529 Iout.n126 0.451012
R15387 Iout.n551 Iout.n126 0.451012
R15388 Iout.n552 Iout.n551 0.451012
R15389 Iout.n552 Iout.n116 0.451012
R15390 Iout.n585 Iout.n116 0.451012
R15391 Iout.n586 Iout.n585 0.451012
R15392 Iout.n586 Iout.n73 0.451012
R15393 Iout.n714 Iout.n73 0.451012
R15394 Iout.n715 Iout.n714 0.451012
R15395 Iout.n715 Iout.n26 0.451012
R15396 Iout.n907 Iout.n26 0.451012
R15397 Iout.n212 Iout.n182 0.451012
R15398 Iout.n281 Iout.n182 0.451012
R15399 Iout.n281 Iout.n280 0.451012
R15400 Iout.n280 Iout.n163 0.451012
R15401 Iout.n406 Iout.n163 0.451012
R15402 Iout.n406 Iout.n405 0.451012
R15403 Iout.n405 Iout.n95 0.451012
R15404 Iout.n628 Iout.n95 0.451012
R15405 Iout.n628 Iout.n627 0.451012
R15406 Iout.n627 Iout.n52 0.451012
R15407 Iout.n757 Iout.n52 0.451012
R15408 Iout.n757 Iout.n756 0.451012
R15409 Iout.n756 Iout.n33 0.451012
R15410 Iout.n858 Iout.n33 0.451012
R15411 Iout.n522 Iout.n145 0.451012
R15412 Iout.n523 Iout.n522 0.451012
R15413 Iout.n523 Iout.n132 0.451012
R15414 Iout.n545 Iout.n132 0.451012
R15415 Iout.n546 Iout.n545 0.451012
R15416 Iout.n546 Iout.n119 0.451012
R15417 Iout.n572 Iout.n119 0.451012
R15418 Iout.n580 Iout.n572 0.451012
R15419 Iout.n580 Iout.n579 0.451012
R15420 Iout.n579 Iout.n76 0.451012
R15421 Iout.n709 Iout.n76 0.451012
R15422 Iout.n709 Iout.n708 0.451012
R15423 Iout.n708 Iout.n25 0.451012
R15424 Iout.n914 Iout.n25 0.451012
R15425 Iout.n216 Iout.n179 0.451012
R15426 Iout.n286 Iout.n179 0.451012
R15427 Iout.n287 Iout.n286 0.451012
R15428 Iout.n287 Iout.n164 0.451012
R15429 Iout.n397 Iout.n164 0.451012
R15430 Iout.n398 Iout.n397 0.451012
R15431 Iout.n398 Iout.n92 0.451012
R15432 Iout.n633 Iout.n92 0.451012
R15433 Iout.n634 Iout.n633 0.451012
R15434 Iout.n634 Iout.n49 0.451012
R15435 Iout.n762 Iout.n49 0.451012
R15436 Iout.n763 Iout.n762 0.451012
R15437 Iout.n763 Iout.n34 0.451012
R15438 Iout.n851 Iout.n34 0.451012
R15439 Iout.n517 Iout.n516 0.451012
R15440 Iout.n517 Iout.n138 0.451012
R15441 Iout.n539 Iout.n138 0.451012
R15442 Iout.n540 Iout.n539 0.451012
R15443 Iout.n540 Iout.n125 0.451012
R15444 Iout.n562 Iout.n125 0.451012
R15445 Iout.n567 Iout.n562 0.451012
R15446 Iout.n567 Iout.n566 0.451012
R15447 Iout.n566 Iout.n79 0.451012
R15448 Iout.n698 Iout.n79 0.451012
R15449 Iout.n702 Iout.n698 0.451012
R15450 Iout.n703 Iout.n702 0.451012
R15451 Iout.n703 Iout.n24 0.451012
R15452 Iout.n921 Iout.n24 0.451012
R15453 Iout.n220 Iout.n176 0.451012
R15454 Iout.n293 Iout.n176 0.451012
R15455 Iout.n293 Iout.n292 0.451012
R15456 Iout.n292 Iout.n165 0.451012
R15457 Iout.n390 Iout.n165 0.451012
R15458 Iout.n390 Iout.n389 0.451012
R15459 Iout.n389 Iout.n89 0.451012
R15460 Iout.n640 Iout.n89 0.451012
R15461 Iout.n640 Iout.n639 0.451012
R15462 Iout.n639 Iout.n46 0.451012
R15463 Iout.n769 Iout.n46 0.451012
R15464 Iout.n769 Iout.n768 0.451012
R15465 Iout.n768 Iout.n35 0.451012
R15466 Iout.n844 Iout.n35 0.451012
R15467 Iout.n511 Iout.n2 0.451012
R15468 Iout.n1005 Iout.n2 0.451012
R15469 Iout.n1005 Iout.n1004 0.451012
R15470 Iout.n1004 Iout.n3 0.451012
R15471 Iout.n986 Iout.n3 0.451012
R15472 Iout.n986 Iout.n985 0.451012
R15473 Iout.n985 Iout.n8 0.451012
R15474 Iout.n967 Iout.n8 0.451012
R15475 Iout.n967 Iout.n966 0.451012
R15476 Iout.n966 Iout.n13 0.451012
R15477 Iout.n948 Iout.n13 0.451012
R15478 Iout.n948 Iout.n947 0.451012
R15479 Iout.n947 Iout.n18 0.451012
R15480 Iout.n929 Iout.n18 0.451012
R15481 Iout.n224 Iout.n170 0.451012
R15482 Iout.n298 Iout.n170 0.451012
R15483 Iout.n299 Iout.n298 0.451012
R15484 Iout.n299 Iout.n166 0.451012
R15485 Iout.n381 Iout.n166 0.451012
R15486 Iout.n382 Iout.n381 0.451012
R15487 Iout.n382 Iout.n83 0.451012
R15488 Iout.n645 Iout.n83 0.451012
R15489 Iout.n646 Iout.n645 0.451012
R15490 Iout.n646 Iout.n40 0.451012
R15491 Iout.n774 Iout.n40 0.451012
R15492 Iout.n775 Iout.n774 0.451012
R15493 Iout.n775 Iout.n36 0.451012
R15494 Iout.n837 Iout.n36 0.451012
R15495 Iout.n1018 Iout.n1017 0.451012
R15496 Iout.n1017 Iout.n0 0.451012
R15497 Iout.n999 Iout.n0 0.451012
R15498 Iout.n999 Iout.n998 0.451012
R15499 Iout.n998 Iout.n6 0.451012
R15500 Iout.n980 Iout.n6 0.451012
R15501 Iout.n980 Iout.n979 0.451012
R15502 Iout.n979 Iout.n11 0.451012
R15503 Iout.n961 Iout.n11 0.451012
R15504 Iout.n961 Iout.n960 0.451012
R15505 Iout.n960 Iout.n16 0.451012
R15506 Iout.n942 Iout.n16 0.451012
R15507 Iout.n942 Iout.n941 0.451012
R15508 Iout.n941 Iout.n21 0.451012
R15509 Iout.n230 Iout.n229 0.451012
R15510 Iout.n230 Iout.n167 0.451012
R15511 Iout.n304 Iout.n167 0.451012
R15512 Iout.n332 Iout.n304 0.451012
R15513 Iout.n374 Iout.n332 0.451012
R15514 Iout.n374 Iout.n373 0.451012
R15515 Iout.n373 Iout.n369 0.451012
R15516 Iout.n369 Iout.n80 0.451012
R15517 Iout.n651 Iout.n80 0.451012
R15518 Iout.n652 Iout.n651 0.451012
R15519 Iout.n652 Iout.n37 0.451012
R15520 Iout.n780 Iout.n37 0.451012
R15521 Iout.n826 Iout.n780 0.451012
R15522 Iout.n830 Iout.n826 0.451012
R15523 Iout.n231 Iout 0.2919
R15524 Iout.n303 Iout 0.2919
R15525 Iout Iout.n300 0.2919
R15526 Iout.n375 Iout 0.2919
R15527 Iout.n380 Iout 0.2919
R15528 Iout.n391 Iout 0.2919
R15529 Iout.n368 Iout 0.2919
R15530 Iout Iout.n365 0.2919
R15531 Iout Iout.n362 0.2919
R15532 Iout Iout.n359 0.2919
R15533 Iout.n650 Iout 0.2919
R15534 Iout Iout.n647 0.2919
R15535 Iout.n638 Iout 0.2919
R15536 Iout Iout.n635 0.2919
R15537 Iout.n626 Iout 0.2919
R15538 Iout.n41 Iout 0.2919
R15539 Iout.n773 Iout 0.2919
R15540 Iout Iout.n770 0.2919
R15541 Iout.n761 Iout 0.2919
R15542 Iout Iout.n758 0.2919
R15543 Iout.n749 Iout 0.2919
R15544 Iout.n825 Iout 0.2919
R15545 Iout Iout.n822 0.2919
R15546 Iout Iout.n819 0.2919
R15547 Iout Iout.n816 0.2919
R15548 Iout Iout.n813 0.2919
R15549 Iout Iout.n810 0.2919
R15550 Iout Iout.n807 0.2919
R15551 Iout.n829 Iout 0.2919
R15552 Iout.n838 Iout 0.2919
R15553 Iout.n843 Iout 0.2919
R15554 Iout.n852 Iout 0.2919
R15555 Iout.n857 Iout 0.2919
R15556 Iout.n866 Iout 0.2919
R15557 Iout.n871 Iout 0.2919
R15558 Iout.n880 Iout 0.2919
R15559 Iout Iout.n925 0.2919
R15560 Iout.n928 Iout 0.2919
R15561 Iout.n922 Iout 0.2919
R15562 Iout.n913 Iout 0.2919
R15563 Iout.n908 Iout 0.2919
R15564 Iout.n899 Iout 0.2919
R15565 Iout.n894 Iout 0.2919
R15566 Iout.n885 Iout 0.2919
R15567 Iout.n831 Iout 0.2919
R15568 Iout.n836 Iout 0.2919
R15569 Iout.n845 Iout 0.2919
R15570 Iout.n850 Iout 0.2919
R15571 Iout.n859 Iout 0.2919
R15572 Iout.n864 Iout 0.2919
R15573 Iout.n873 Iout 0.2919
R15574 Iout.n878 Iout 0.2919
R15575 Iout.n887 Iout 0.2919
R15576 Iout.n892 Iout 0.2919
R15577 Iout.n933 Iout 0.2919
R15578 Iout.n930 Iout 0.2919
R15579 Iout.n920 Iout 0.2919
R15580 Iout.n915 Iout 0.2919
R15581 Iout.n906 Iout 0.2919
R15582 Iout.n901 Iout 0.2919
R15583 Iout.n940 Iout 0.2919
R15584 Iout Iout.n783 0.2919
R15585 Iout Iout.n786 0.2919
R15586 Iout Iout.n789 0.2919
R15587 Iout Iout.n792 0.2919
R15588 Iout Iout.n795 0.2919
R15589 Iout Iout.n798 0.2919
R15590 Iout Iout.n801 0.2919
R15591 Iout Iout.n804 0.2919
R15592 Iout.n779 Iout 0.2919
R15593 Iout Iout.n776 0.2919
R15594 Iout.n767 Iout 0.2919
R15595 Iout Iout.n764 0.2919
R15596 Iout.n755 Iout 0.2919
R15597 Iout Iout.n752 0.2919
R15598 Iout.n743 Iout 0.2919
R15599 Iout Iout.n740 0.2919
R15600 Iout.n731 Iout 0.2919
R15601 Iout Iout.n728 0.2919
R15602 Iout.n719 Iout 0.2919
R15603 Iout Iout.n943 0.2919
R15604 Iout.n946 Iout 0.2919
R15605 Iout Iout.n704 0.2919
R15606 Iout.n707 Iout 0.2919
R15607 Iout Iout.n716 0.2919
R15608 Iout.n952 Iout 0.2919
R15609 Iout.n949 Iout 0.2919
R15610 Iout.n701 Iout 0.2919
R15611 Iout Iout.n710 0.2919
R15612 Iout.n713 Iout 0.2919
R15613 Iout Iout.n722 0.2919
R15614 Iout.n725 Iout 0.2919
R15615 Iout Iout.n734 0.2919
R15616 Iout.n737 Iout 0.2919
R15617 Iout Iout.n746 0.2919
R15618 Iout.n653 Iout 0.2919
R15619 Iout.n656 Iout 0.2919
R15620 Iout.n659 Iout 0.2919
R15621 Iout.n662 Iout 0.2919
R15622 Iout.n665 Iout 0.2919
R15623 Iout.n668 Iout 0.2919
R15624 Iout.n671 Iout 0.2919
R15625 Iout.n674 Iout 0.2919
R15626 Iout.n677 Iout 0.2919
R15627 Iout.n680 Iout 0.2919
R15628 Iout.n683 Iout 0.2919
R15629 Iout.n686 Iout 0.2919
R15630 Iout.n959 Iout 0.2919
R15631 Iout Iout.n694 0.2919
R15632 Iout.n697 Iout 0.2919
R15633 Iout.n689 Iout 0.2919
R15634 Iout Iout.n962 0.2919
R15635 Iout.n965 Iout 0.2919
R15636 Iout Iout.n575 0.2919
R15637 Iout.n578 Iout 0.2919
R15638 Iout Iout.n587 0.2919
R15639 Iout.n590 Iout 0.2919
R15640 Iout Iout.n599 0.2919
R15641 Iout.n602 Iout 0.2919
R15642 Iout Iout.n611 0.2919
R15643 Iout.n614 Iout 0.2919
R15644 Iout Iout.n623 0.2919
R15645 Iout.n84 Iout 0.2919
R15646 Iout.n644 Iout 0.2919
R15647 Iout Iout.n641 0.2919
R15648 Iout.n632 Iout 0.2919
R15649 Iout Iout.n629 0.2919
R15650 Iout.n620 Iout 0.2919
R15651 Iout Iout.n617 0.2919
R15652 Iout.n608 Iout 0.2919
R15653 Iout Iout.n605 0.2919
R15654 Iout.n596 Iout 0.2919
R15655 Iout Iout.n593 0.2919
R15656 Iout.n584 Iout 0.2919
R15657 Iout Iout.n581 0.2919
R15658 Iout.n971 Iout 0.2919
R15659 Iout.n968 Iout 0.2919
R15660 Iout.n565 Iout 0.2919
R15661 Iout.n978 Iout 0.2919
R15662 Iout Iout.n122 0.2919
R15663 Iout Iout.n568 0.2919
R15664 Iout.n571 Iout 0.2919
R15665 Iout Iout.n335 0.2919
R15666 Iout Iout.n338 0.2919
R15667 Iout Iout.n341 0.2919
R15668 Iout Iout.n344 0.2919
R15669 Iout Iout.n347 0.2919
R15670 Iout Iout.n350 0.2919
R15671 Iout Iout.n353 0.2919
R15672 Iout Iout.n356 0.2919
R15673 Iout.n372 Iout 0.2919
R15674 Iout.n383 Iout 0.2919
R15675 Iout.n388 Iout 0.2919
R15676 Iout.n399 Iout 0.2919
R15677 Iout.n404 Iout 0.2919
R15678 Iout.n415 Iout 0.2919
R15679 Iout.n420 Iout 0.2919
R15680 Iout.n431 Iout 0.2919
R15681 Iout.n443 Iout 0.2919
R15682 Iout Iout.n440 0.2919
R15683 Iout Iout.n437 0.2919
R15684 Iout.n553 Iout 0.2919
R15685 Iout.n556 Iout 0.2919
R15686 Iout.n561 Iout 0.2919
R15687 Iout Iout.n981 0.2919
R15688 Iout.n984 Iout 0.2919
R15689 Iout.n990 Iout 0.2919
R15690 Iout.n987 Iout 0.2919
R15691 Iout Iout.n129 0.2919
R15692 Iout Iout.n547 0.2919
R15693 Iout.n550 Iout 0.2919
R15694 Iout Iout.n451 0.2919
R15695 Iout.n454 Iout 0.2919
R15696 Iout.n446 Iout 0.2919
R15697 Iout.n428 Iout 0.2919
R15698 Iout.n423 Iout 0.2919
R15699 Iout.n412 Iout 0.2919
R15700 Iout.n407 Iout 0.2919
R15701 Iout.n396 Iout 0.2919
R15702 Iout.n331 Iout 0.2919
R15703 Iout Iout.n328 0.2919
R15704 Iout Iout.n325 0.2919
R15705 Iout Iout.n322 0.2919
R15706 Iout Iout.n319 0.2919
R15707 Iout Iout.n316 0.2919
R15708 Iout Iout.n313 0.2919
R15709 Iout Iout.n310 0.2919
R15710 Iout Iout.n307 0.2919
R15711 Iout.n457 Iout 0.2919
R15712 Iout.n465 Iout 0.2919
R15713 Iout Iout.n462 0.2919
R15714 Iout.n544 Iout 0.2919
R15715 Iout Iout.n541 0.2919
R15716 Iout Iout.n135 0.2919
R15717 Iout.n997 Iout 0.2919
R15718 Iout Iout.n1000 0.2919
R15719 Iout.n1003 Iout 0.2919
R15720 Iout.n538 Iout 0.2919
R15721 Iout.n533 Iout 0.2919
R15722 Iout.n530 Iout 0.2919
R15723 Iout Iout.n468 0.2919
R15724 Iout Iout.n471 0.2919
R15725 Iout.n474 Iout 0.2919
R15726 Iout Iout.n264 0.2919
R15727 Iout.n267 Iout 0.2919
R15728 Iout Iout.n276 0.2919
R15729 Iout.n279 Iout 0.2919
R15730 Iout Iout.n288 0.2919
R15731 Iout.n291 Iout 0.2919
R15732 Iout.n171 Iout 0.2919
R15733 Iout.n297 Iout 0.2919
R15734 Iout Iout.n294 0.2919
R15735 Iout.n285 Iout 0.2919
R15736 Iout Iout.n282 0.2919
R15737 Iout.n273 Iout 0.2919
R15738 Iout Iout.n270 0.2919
R15739 Iout.n261 Iout 0.2919
R15740 Iout.n477 Iout 0.2919
R15741 Iout.n485 Iout 0.2919
R15742 Iout Iout.n482 0.2919
R15743 Iout.n527 Iout 0.2919
R15744 Iout Iout.n524 0.2919
R15745 Iout Iout.n142 0.2919
R15746 Iout.n1006 Iout 0.2919
R15747 Iout.n1009 Iout 0.2919
R15748 Iout.n1016 Iout 0.2919
R15749 Iout Iout.n148 0.2919
R15750 Iout Iout.n518 0.2919
R15751 Iout.n521 Iout 0.2919
R15752 Iout Iout.n493 0.2919
R15753 Iout.n496 Iout 0.2919
R15754 Iout.n488 Iout 0.2919
R15755 Iout Iout.n254 0.2919
R15756 Iout.n257 Iout 0.2919
R15757 Iout.n249 Iout 0.2919
R15758 Iout.n246 Iout 0.2919
R15759 Iout.n243 Iout 0.2919
R15760 Iout.n240 Iout 0.2919
R15761 Iout.n237 Iout 0.2919
R15762 Iout.n234 Iout 0.2919
R15763 Iout.n228 Iout 0.2919
R15764 Iout Iout.n225 0.2919
R15765 Iout Iout.n221 0.2919
R15766 Iout Iout.n217 0.2919
R15767 Iout Iout.n213 0.2919
R15768 Iout Iout.n209 0.2919
R15769 Iout Iout.n205 0.2919
R15770 Iout Iout.n201 0.2919
R15771 Iout Iout.n198 0.2919
R15772 Iout Iout.n194 0.2919
R15773 Iout.n499 Iout 0.2919
R15774 Iout.n503 Iout 0.2919
R15775 Iout.n506 Iout 0.2919
R15776 Iout.n515 Iout 0.2919
R15777 Iout Iout.n512 0.2919
R15778 Iout.n1019 Iout 0.2919
R15779 Iout.n1013 Iout.n1012 0.092855
R15780 Iout.n1012 Iout.n1 0.092855
R15781 Iout.n994 Iout.n1 0.092855
R15782 Iout.n994 Iout.n993 0.092855
R15783 Iout.n993 Iout.n7 0.092855
R15784 Iout.n975 Iout.n7 0.092855
R15785 Iout.n975 Iout.n974 0.092855
R15786 Iout.n974 Iout.n12 0.092855
R15787 Iout.n956 Iout.n12 0.092855
R15788 Iout.n956 Iout.n955 0.092855
R15789 Iout.n955 Iout.n17 0.092855
R15790 Iout.n937 Iout.n17 0.092855
R15791 Iout.n937 Iout.n936 0.092855
R15792 Iout.n197 Iout 0.0818902
R15793 Iout.n191 Iout 0.0818902
R15794 Iout.n152 Iout 0.0818902
R15795 Iout.n204 Iout 0.0818902
R15796 Iout.n498 Iout 0.0818902
R15797 Iout.n208 Iout 0.0818902
R15798 Iout.n502 Iout 0.0818902
R15799 Iout.n212 Iout 0.0818902
R15800 Iout.n145 Iout 0.0818902
R15801 Iout.n216 Iout 0.0818902
R15802 Iout.n516 Iout 0.0818902
R15803 Iout.n220 Iout 0.0818902
R15804 Iout.n511 Iout 0.0818902
R15805 Iout.n224 Iout 0.0818902
R15806 Iout.n1018 Iout 0.0818902
R15807 Iout.n229 Iout 0.0818902
R15808 Iout.n1013 Iout 0.072645
R15809 Iout.n302 Iout 0.0532071
R15810 Iout Iout.n377 0.0532071
R15811 Iout.n379 Iout 0.0532071
R15812 Iout.n367 Iout 0.0532071
R15813 Iout.n364 Iout 0.0532071
R15814 Iout.n361 Iout 0.0532071
R15815 Iout.n649 Iout 0.0532071
R15816 Iout Iout.n82 0.0532071
R15817 Iout.n637 Iout 0.0532071
R15818 Iout Iout.n91 0.0532071
R15819 Iout Iout.n43 0.0532071
R15820 Iout.n772 Iout 0.0532071
R15821 Iout Iout.n45 0.0532071
R15822 Iout.n760 Iout 0.0532071
R15823 Iout Iout.n51 0.0532071
R15824 Iout.n824 Iout 0.0532071
R15825 Iout.n821 Iout 0.0532071
R15826 Iout.n818 Iout 0.0532071
R15827 Iout.n815 Iout 0.0532071
R15828 Iout.n812 Iout 0.0532071
R15829 Iout.n809 Iout 0.0532071
R15830 Iout.n828 Iout 0.0532071
R15831 Iout Iout.n840 0.0532071
R15832 Iout.n842 Iout 0.0532071
R15833 Iout Iout.n854 0.0532071
R15834 Iout.n856 Iout 0.0532071
R15835 Iout Iout.n868 0.0532071
R15836 Iout.n870 Iout 0.0532071
R15837 Iout.n927 Iout 0.0532071
R15838 Iout Iout.n924 0.0532071
R15839 Iout.n912 Iout 0.0532071
R15840 Iout Iout.n910 0.0532071
R15841 Iout.n898 Iout 0.0532071
R15842 Iout Iout.n896 0.0532071
R15843 Iout.n884 Iout 0.0532071
R15844 Iout Iout.n882 0.0532071
R15845 Iout Iout.n833 0.0532071
R15846 Iout.n835 Iout 0.0532071
R15847 Iout Iout.n847 0.0532071
R15848 Iout.n849 Iout 0.0532071
R15849 Iout Iout.n861 0.0532071
R15850 Iout.n863 Iout 0.0532071
R15851 Iout Iout.n875 0.0532071
R15852 Iout.n877 Iout 0.0532071
R15853 Iout Iout.n889 0.0532071
R15854 Iout Iout.n932 0.0532071
R15855 Iout.n919 Iout 0.0532071
R15856 Iout Iout.n917 0.0532071
R15857 Iout.n905 Iout 0.0532071
R15858 Iout Iout.n903 0.0532071
R15859 Iout.n891 Iout 0.0532071
R15860 Iout.n782 Iout 0.0532071
R15861 Iout.n785 Iout 0.0532071
R15862 Iout.n788 Iout 0.0532071
R15863 Iout.n791 Iout 0.0532071
R15864 Iout.n794 Iout 0.0532071
R15865 Iout.n797 Iout 0.0532071
R15866 Iout.n800 Iout 0.0532071
R15867 Iout.n803 Iout 0.0532071
R15868 Iout.n806 Iout 0.0532071
R15869 Iout.n778 Iout 0.0532071
R15870 Iout Iout.n39 0.0532071
R15871 Iout.n766 Iout 0.0532071
R15872 Iout Iout.n48 0.0532071
R15873 Iout.n754 Iout 0.0532071
R15874 Iout Iout.n54 0.0532071
R15875 Iout.n742 Iout 0.0532071
R15876 Iout Iout.n60 0.0532071
R15877 Iout.n730 Iout 0.0532071
R15878 Iout Iout.n66 0.0532071
R15879 Iout.n945 Iout 0.0532071
R15880 Iout.n78 Iout 0.0532071
R15881 Iout.n706 Iout 0.0532071
R15882 Iout Iout.n72 0.0532071
R15883 Iout.n718 Iout 0.0532071
R15884 Iout Iout.n951 0.0532071
R15885 Iout.n700 Iout 0.0532071
R15886 Iout Iout.n75 0.0532071
R15887 Iout.n712 Iout 0.0532071
R15888 Iout Iout.n69 0.0532071
R15889 Iout.n724 Iout 0.0532071
R15890 Iout Iout.n63 0.0532071
R15891 Iout.n736 Iout 0.0532071
R15892 Iout Iout.n57 0.0532071
R15893 Iout.n748 Iout 0.0532071
R15894 Iout Iout.n655 0.0532071
R15895 Iout Iout.n658 0.0532071
R15896 Iout Iout.n661 0.0532071
R15897 Iout Iout.n664 0.0532071
R15898 Iout Iout.n667 0.0532071
R15899 Iout Iout.n670 0.0532071
R15900 Iout Iout.n673 0.0532071
R15901 Iout Iout.n676 0.0532071
R15902 Iout Iout.n679 0.0532071
R15903 Iout Iout.n682 0.0532071
R15904 Iout Iout.n685 0.0532071
R15905 Iout.n693 Iout 0.0532071
R15906 Iout.n696 Iout 0.0532071
R15907 Iout Iout.n691 0.0532071
R15908 Iout Iout.n688 0.0532071
R15909 Iout.n964 Iout 0.0532071
R15910 Iout.n574 Iout 0.0532071
R15911 Iout.n577 Iout 0.0532071
R15912 Iout Iout.n115 0.0532071
R15913 Iout.n589 Iout 0.0532071
R15914 Iout Iout.n109 0.0532071
R15915 Iout.n601 Iout 0.0532071
R15916 Iout Iout.n103 0.0532071
R15917 Iout.n613 Iout 0.0532071
R15918 Iout Iout.n97 0.0532071
R15919 Iout.n625 Iout 0.0532071
R15920 Iout Iout.n86 0.0532071
R15921 Iout.n643 Iout 0.0532071
R15922 Iout Iout.n88 0.0532071
R15923 Iout.n631 Iout 0.0532071
R15924 Iout Iout.n94 0.0532071
R15925 Iout.n619 Iout 0.0532071
R15926 Iout Iout.n100 0.0532071
R15927 Iout.n607 Iout 0.0532071
R15928 Iout Iout.n106 0.0532071
R15929 Iout.n595 Iout 0.0532071
R15930 Iout Iout.n112 0.0532071
R15931 Iout.n583 Iout 0.0532071
R15932 Iout Iout.n970 0.0532071
R15933 Iout.n564 Iout 0.0532071
R15934 Iout Iout.n118 0.0532071
R15935 Iout.n121 Iout 0.0532071
R15936 Iout.n124 Iout 0.0532071
R15937 Iout.n570 Iout 0.0532071
R15938 Iout.n334 Iout 0.0532071
R15939 Iout.n337 Iout 0.0532071
R15940 Iout.n340 Iout 0.0532071
R15941 Iout.n343 Iout 0.0532071
R15942 Iout.n346 Iout 0.0532071
R15943 Iout.n349 Iout 0.0532071
R15944 Iout.n352 Iout 0.0532071
R15945 Iout.n355 Iout 0.0532071
R15946 Iout.n358 Iout 0.0532071
R15947 Iout.n371 Iout 0.0532071
R15948 Iout Iout.n385 0.0532071
R15949 Iout.n387 Iout 0.0532071
R15950 Iout Iout.n401 0.0532071
R15951 Iout.n403 Iout 0.0532071
R15952 Iout Iout.n417 0.0532071
R15953 Iout.n419 Iout 0.0532071
R15954 Iout Iout.n433 0.0532071
R15955 Iout.n442 Iout 0.0532071
R15956 Iout.n439 Iout 0.0532071
R15957 Iout.n435 Iout 0.0532071
R15958 Iout Iout.n555 0.0532071
R15959 Iout Iout.n558 0.0532071
R15960 Iout.n983 Iout 0.0532071
R15961 Iout.n560 Iout 0.0532071
R15962 Iout Iout.n989 0.0532071
R15963 Iout.n128 Iout 0.0532071
R15964 Iout.n131 Iout 0.0532071
R15965 Iout.n549 Iout 0.0532071
R15966 Iout.n450 Iout 0.0532071
R15967 Iout.n453 Iout 0.0532071
R15968 Iout Iout.n448 0.0532071
R15969 Iout.n427 Iout 0.0532071
R15970 Iout Iout.n425 0.0532071
R15971 Iout.n411 Iout 0.0532071
R15972 Iout Iout.n409 0.0532071
R15973 Iout.n395 Iout 0.0532071
R15974 Iout Iout.n393 0.0532071
R15975 Iout.n330 Iout 0.0532071
R15976 Iout.n327 Iout 0.0532071
R15977 Iout.n324 Iout 0.0532071
R15978 Iout.n321 Iout 0.0532071
R15979 Iout.n318 Iout 0.0532071
R15980 Iout.n315 Iout 0.0532071
R15981 Iout.n312 Iout 0.0532071
R15982 Iout.n309 Iout 0.0532071
R15983 Iout.n306 Iout 0.0532071
R15984 Iout Iout.n459 0.0532071
R15985 Iout.n464 Iout 0.0532071
R15986 Iout.n461 Iout 0.0532071
R15987 Iout.n543 Iout 0.0532071
R15988 Iout.n137 Iout 0.0532071
R15989 Iout.n134 Iout 0.0532071
R15990 Iout.n1002 Iout 0.0532071
R15991 Iout.n537 Iout 0.0532071
R15992 Iout Iout.n535 0.0532071
R15993 Iout Iout.n532 0.0532071
R15994 Iout.n157 Iout 0.0532071
R15995 Iout.n470 Iout 0.0532071
R15996 Iout.n473 Iout 0.0532071
R15997 Iout.n190 Iout 0.0532071
R15998 Iout.n266 Iout 0.0532071
R15999 Iout Iout.n184 0.0532071
R16000 Iout.n278 Iout 0.0532071
R16001 Iout Iout.n178 0.0532071
R16002 Iout.n290 Iout 0.0532071
R16003 Iout Iout.n169 0.0532071
R16004 Iout Iout.n173 0.0532071
R16005 Iout.n296 Iout 0.0532071
R16006 Iout Iout.n175 0.0532071
R16007 Iout.n284 Iout 0.0532071
R16008 Iout Iout.n181 0.0532071
R16009 Iout.n272 Iout 0.0532071
R16010 Iout Iout.n187 0.0532071
R16011 Iout.n260 Iout 0.0532071
R16012 Iout Iout.n479 0.0532071
R16013 Iout.n484 Iout 0.0532071
R16014 Iout.n481 Iout 0.0532071
R16015 Iout.n526 Iout 0.0532071
R16016 Iout.n144 Iout 0.0532071
R16017 Iout.n141 Iout 0.0532071
R16018 Iout Iout.n1008 0.0532071
R16019 Iout.n147 Iout 0.0532071
R16020 Iout.n150 Iout 0.0532071
R16021 Iout.n520 Iout 0.0532071
R16022 Iout.n492 Iout 0.0532071
R16023 Iout.n495 Iout 0.0532071
R16024 Iout Iout.n490 0.0532071
R16025 Iout.n253 Iout 0.0532071
R16026 Iout.n256 Iout 0.0532071
R16027 Iout Iout.n251 0.0532071
R16028 Iout Iout.n248 0.0532071
R16029 Iout Iout.n245 0.0532071
R16030 Iout Iout.n242 0.0532071
R16031 Iout Iout.n239 0.0532071
R16032 Iout Iout.n236 0.0532071
R16033 Iout Iout.n233 0.0532071
R16034 Iout.n227 Iout 0.0532071
R16035 Iout.n223 Iout 0.0532071
R16036 Iout.n219 Iout 0.0532071
R16037 Iout.n215 Iout 0.0532071
R16038 Iout.n211 Iout 0.0532071
R16039 Iout.n207 Iout 0.0532071
R16040 Iout.n203 Iout 0.0532071
R16041 Iout.n200 Iout 0.0532071
R16042 Iout.n196 Iout 0.0532071
R16043 Iout.n193 Iout 0.0532071
R16044 Iout Iout.n501 0.0532071
R16045 Iout Iout.n505 0.0532071
R16046 Iout Iout.n508 0.0532071
R16047 Iout.n514 Iout 0.0532071
R16048 Iout.n510 Iout 0.0532071
R16049 Iout.n1020 Iout 0.03925
R16050 Iout.n509 Iout 0.03925
R16051 Iout.n513 Iout 0.03925
R16052 Iout.n507 Iout 0.03925
R16053 Iout.n504 Iout 0.03925
R16054 Iout.n500 Iout 0.03925
R16055 Iout.n192 Iout 0.03925
R16056 Iout.n195 Iout 0.03925
R16057 Iout.n199 Iout 0.03925
R16058 Iout.n202 Iout 0.03925
R16059 Iout.n206 Iout 0.03925
R16060 Iout.n210 Iout 0.03925
R16061 Iout.n214 Iout 0.03925
R16062 Iout.n218 Iout 0.03925
R16063 Iout.n222 Iout 0.03925
R16064 Iout.n226 Iout 0.03925
R16065 Iout.n232 Iout 0.03925
R16066 Iout.n235 Iout 0.03925
R16067 Iout.n238 Iout 0.03925
R16068 Iout.n241 Iout 0.03925
R16069 Iout.n244 Iout 0.03925
R16070 Iout.n247 Iout 0.03925
R16071 Iout.n250 Iout 0.03925
R16072 Iout.n255 Iout 0.03925
R16073 Iout.n252 Iout 0.03925
R16074 Iout.n489 Iout 0.03925
R16075 Iout.n494 Iout 0.03925
R16076 Iout.n491 Iout 0.03925
R16077 Iout.n519 Iout 0.03925
R16078 Iout.n149 Iout 0.03925
R16079 Iout.n146 Iout 0.03925
R16080 Iout.n1010 Iout 0.03925
R16081 Iout.n1007 Iout 0.03925
R16082 Iout.n140 Iout 0.03925
R16083 Iout.n143 Iout 0.03925
R16084 Iout.n525 Iout 0.03925
R16085 Iout.n480 Iout 0.03925
R16086 Iout.n483 Iout 0.03925
R16087 Iout.n478 Iout 0.03925
R16088 Iout.n259 Iout 0.03925
R16089 Iout.n186 Iout 0.03925
R16090 Iout.n271 Iout 0.03925
R16091 Iout.n180 Iout 0.03925
R16092 Iout.n283 Iout 0.03925
R16093 Iout.n174 Iout 0.03925
R16094 Iout.n168 Iout 0.03925
R16095 Iout.n301 Iout 0.03925
R16096 Iout.n289 Iout 0.03925
R16097 Iout.n177 Iout 0.03925
R16098 Iout.n277 Iout 0.03925
R16099 Iout.n183 Iout 0.03925
R16100 Iout.n265 Iout 0.03925
R16101 Iout.n189 Iout 0.03925
R16102 Iout.n472 Iout 0.03925
R16103 Iout.n469 Iout 0.03925
R16104 Iout.n156 Iout 0.03925
R16105 Iout.n531 Iout 0.03925
R16106 Iout.n534 Iout 0.03925
R16107 Iout.n536 Iout 0.03925
R16108 Iout.n133 Iout 0.03925
R16109 Iout.n136 Iout 0.03925
R16110 Iout.n542 Iout 0.03925
R16111 Iout.n460 Iout 0.03925
R16112 Iout.n463 Iout 0.03925
R16113 Iout.n458 Iout 0.03925
R16114 Iout.n305 Iout 0.03925
R16115 Iout.n308 Iout 0.03925
R16116 Iout.n311 Iout 0.03925
R16117 Iout.n314 Iout 0.03925
R16118 Iout.n317 Iout 0.03925
R16119 Iout.n320 Iout 0.03925
R16120 Iout.n392 Iout 0.03925
R16121 Iout.n378 Iout 0.03925
R16122 Iout.n376 Iout 0.03925
R16123 Iout.n394 Iout 0.03925
R16124 Iout.n408 Iout 0.03925
R16125 Iout.n410 Iout 0.03925
R16126 Iout.n424 Iout 0.03925
R16127 Iout.n426 Iout 0.03925
R16128 Iout.n447 Iout 0.03925
R16129 Iout.n452 Iout 0.03925
R16130 Iout.n449 Iout 0.03925
R16131 Iout.n548 Iout 0.03925
R16132 Iout.n130 Iout 0.03925
R16133 Iout.n559 Iout 0.03925
R16134 Iout.n557 Iout 0.03925
R16135 Iout.n554 Iout 0.03925
R16136 Iout.n434 Iout 0.03925
R16137 Iout.n438 Iout 0.03925
R16138 Iout.n441 Iout 0.03925
R16139 Iout.n432 Iout 0.03925
R16140 Iout.n418 Iout 0.03925
R16141 Iout.n416 Iout 0.03925
R16142 Iout.n402 Iout 0.03925
R16143 Iout.n357 Iout 0.03925
R16144 Iout.n360 Iout 0.03925
R16145 Iout.n363 Iout 0.03925
R16146 Iout.n366 Iout 0.03925
R16147 Iout.n354 Iout 0.03925
R16148 Iout.n351 Iout 0.03925
R16149 Iout.n348 Iout 0.03925
R16150 Iout.n345 Iout 0.03925
R16151 Iout.n342 Iout 0.03925
R16152 Iout.n339 Iout 0.03925
R16153 Iout.n336 Iout 0.03925
R16154 Iout.n333 Iout 0.03925
R16155 Iout.n117 Iout 0.03925
R16156 Iout.n582 Iout 0.03925
R16157 Iout.n111 Iout 0.03925
R16158 Iout.n594 Iout 0.03925
R16159 Iout.n105 Iout 0.03925
R16160 Iout.n606 Iout 0.03925
R16161 Iout.n99 Iout 0.03925
R16162 Iout.n618 Iout 0.03925
R16163 Iout.n624 Iout 0.03925
R16164 Iout.n90 Iout 0.03925
R16165 Iout.n636 Iout 0.03925
R16166 Iout.n81 Iout 0.03925
R16167 Iout.n648 Iout 0.03925
R16168 Iout.n96 Iout 0.03925
R16169 Iout.n612 Iout 0.03925
R16170 Iout.n102 Iout 0.03925
R16171 Iout.n600 Iout 0.03925
R16172 Iout.n108 Iout 0.03925
R16173 Iout.n588 Iout 0.03925
R16174 Iout.n687 Iout 0.03925
R16175 Iout.n684 Iout 0.03925
R16176 Iout.n681 Iout 0.03925
R16177 Iout.n678 Iout 0.03925
R16178 Iout.n675 Iout 0.03925
R16179 Iout.n672 Iout 0.03925
R16180 Iout.n747 Iout 0.03925
R16181 Iout.n50 Iout 0.03925
R16182 Iout.n759 Iout 0.03925
R16183 Iout.n44 Iout 0.03925
R16184 Iout.n771 Iout 0.03925
R16185 Iout.n42 Iout 0.03925
R16186 Iout.n56 Iout 0.03925
R16187 Iout.n735 Iout 0.03925
R16188 Iout.n62 Iout 0.03925
R16189 Iout.n723 Iout 0.03925
R16190 Iout.n717 Iout 0.03925
R16191 Iout.n65 Iout 0.03925
R16192 Iout.n729 Iout 0.03925
R16193 Iout.n59 Iout 0.03925
R16194 Iout.n805 Iout 0.03925
R16195 Iout.n808 Iout 0.03925
R16196 Iout.n811 Iout 0.03925
R16197 Iout.n814 Iout 0.03925
R16198 Iout.n817 Iout 0.03925
R16199 Iout.n820 Iout 0.03925
R16200 Iout.n823 Iout 0.03925
R16201 Iout.n802 Iout 0.03925
R16202 Iout.n799 Iout 0.03925
R16203 Iout.n890 Iout 0.03925
R16204 Iout.n888 Iout 0.03925
R16205 Iout.n881 Iout 0.03925
R16206 Iout.n869 Iout 0.03925
R16207 Iout.n867 Iout 0.03925
R16208 Iout.n855 Iout 0.03925
R16209 Iout.n853 Iout 0.03925
R16210 Iout.n841 Iout 0.03925
R16211 Iout.n839 Iout 0.03925
R16212 Iout.n827 Iout 0.03925
R16213 Iout.n883 Iout 0.03925
R16214 Iout.n895 Iout 0.03925
R16215 Iout.n897 Iout 0.03925
R16216 Iout.n909 Iout 0.03925
R16217 Iout.n911 Iout 0.03925
R16218 Iout.n923 Iout 0.03925
R16219 Iout.n926 Iout 0.03925
R16220 Iout.n22 Iout 0.03925
R16221 Iout.n876 Iout 0.03925
R16222 Iout.n874 Iout 0.03925
R16223 Iout.n862 Iout 0.03925
R16224 Iout.n860 Iout 0.03925
R16225 Iout.n848 Iout 0.03925
R16226 Iout.n846 Iout 0.03925
R16227 Iout.n834 Iout 0.03925
R16228 Iout.n832 Iout 0.03925
R16229 Iout.n902 Iout 0.03925
R16230 Iout.n904 Iout 0.03925
R16231 Iout.n916 Iout 0.03925
R16232 Iout.n918 Iout 0.03925
R16233 Iout.n931 Iout 0.03925
R16234 Iout.n934 Iout 0.03925
R16235 Iout.n796 Iout 0.03925
R16236 Iout.n793 Iout 0.03925
R16237 Iout.n790 Iout 0.03925
R16238 Iout.n787 Iout 0.03925
R16239 Iout.n784 Iout 0.03925
R16240 Iout.n781 Iout 0.03925
R16241 Iout.n938 Iout 0.03925
R16242 Iout.n741 Iout 0.03925
R16243 Iout.n53 Iout 0.03925
R16244 Iout.n753 Iout 0.03925
R16245 Iout.n47 Iout 0.03925
R16246 Iout.n765 Iout 0.03925
R16247 Iout.n38 Iout 0.03925
R16248 Iout.n777 Iout 0.03925
R16249 Iout.n71 Iout 0.03925
R16250 Iout.n705 Iout 0.03925
R16251 Iout.n77 Iout 0.03925
R16252 Iout.n944 Iout 0.03925
R16253 Iout.n19 Iout 0.03925
R16254 Iout.n68 Iout 0.03925
R16255 Iout.n711 Iout 0.03925
R16256 Iout.n74 Iout 0.03925
R16257 Iout.n699 Iout 0.03925
R16258 Iout.n950 Iout 0.03925
R16259 Iout.n953 Iout 0.03925
R16260 Iout.n669 Iout 0.03925
R16261 Iout.n666 Iout 0.03925
R16262 Iout.n663 Iout 0.03925
R16263 Iout.n660 Iout 0.03925
R16264 Iout.n657 Iout 0.03925
R16265 Iout.n654 Iout 0.03925
R16266 Iout.n690 Iout 0.03925
R16267 Iout.n695 Iout 0.03925
R16268 Iout.n692 Iout 0.03925
R16269 Iout.n957 Iout 0.03925
R16270 Iout.n114 Iout 0.03925
R16271 Iout.n576 Iout 0.03925
R16272 Iout.n573 Iout 0.03925
R16273 Iout.n963 Iout 0.03925
R16274 Iout.n14 Iout 0.03925
R16275 Iout.n93 Iout 0.03925
R16276 Iout.n630 Iout 0.03925
R16277 Iout.n87 Iout 0.03925
R16278 Iout.n642 Iout 0.03925
R16279 Iout.n85 Iout 0.03925
R16280 Iout.n563 Iout 0.03925
R16281 Iout.n969 Iout 0.03925
R16282 Iout.n972 Iout 0.03925
R16283 Iout.n569 Iout 0.03925
R16284 Iout.n123 Iout 0.03925
R16285 Iout.n120 Iout 0.03925
R16286 Iout.n976 Iout 0.03925
R16287 Iout.n400 Iout 0.03925
R16288 Iout.n386 Iout 0.03925
R16289 Iout.n384 Iout 0.03925
R16290 Iout.n370 Iout 0.03925
R16291 Iout.n982 Iout 0.03925
R16292 Iout.n9 Iout 0.03925
R16293 Iout.n127 Iout 0.03925
R16294 Iout.n988 Iout 0.03925
R16295 Iout.n991 Iout 0.03925
R16296 Iout.n323 Iout 0.03925
R16297 Iout.n326 Iout 0.03925
R16298 Iout.n329 Iout 0.03925
R16299 Iout.n995 Iout 0.03925
R16300 Iout.n1001 Iout 0.03925
R16301 Iout.n4 Iout 0.03925
R16302 Iout.n295 Iout 0.03925
R16303 Iout.n172 Iout 0.03925
R16304 Iout.n1014 Iout 0.03925
R16305 Iout.n1022 Iout 0.02071
R16306 Iout Iout.n1022 0.00379
R16307 Iout.n303 Iout.n302 0.00105952
R16308 Iout.n377 Iout.n375 0.00105952
R16309 Iout.n380 Iout.n379 0.00105952
R16310 Iout.n368 Iout.n367 0.00105952
R16311 Iout.n365 Iout.n364 0.00105952
R16312 Iout.n362 Iout.n361 0.00105952
R16313 Iout.n650 Iout.n649 0.00105952
R16314 Iout.n647 Iout.n82 0.00105952
R16315 Iout.n638 Iout.n637 0.00105952
R16316 Iout.n635 Iout.n91 0.00105952
R16317 Iout.n43 Iout.n41 0.00105952
R16318 Iout.n773 Iout.n772 0.00105952
R16319 Iout.n770 Iout.n45 0.00105952
R16320 Iout.n761 Iout.n760 0.00105952
R16321 Iout.n758 Iout.n51 0.00105952
R16322 Iout.n825 Iout.n824 0.00105952
R16323 Iout.n822 Iout.n821 0.00105952
R16324 Iout.n819 Iout.n818 0.00105952
R16325 Iout.n816 Iout.n815 0.00105952
R16326 Iout.n813 Iout.n812 0.00105952
R16327 Iout.n810 Iout.n809 0.00105952
R16328 Iout.n829 Iout.n828 0.00105952
R16329 Iout.n840 Iout.n838 0.00105952
R16330 Iout.n843 Iout.n842 0.00105952
R16331 Iout.n854 Iout.n852 0.00105952
R16332 Iout.n857 Iout.n856 0.00105952
R16333 Iout.n868 Iout.n866 0.00105952
R16334 Iout.n871 Iout.n870 0.00105952
R16335 Iout.n925 Iout.n23 0.00105952
R16336 Iout.n928 Iout.n927 0.00105952
R16337 Iout.n924 Iout.n922 0.00105952
R16338 Iout.n913 Iout.n912 0.00105952
R16339 Iout.n910 Iout.n908 0.00105952
R16340 Iout.n899 Iout.n898 0.00105952
R16341 Iout.n896 Iout.n894 0.00105952
R16342 Iout.n885 Iout.n884 0.00105952
R16343 Iout.n882 Iout.n880 0.00105952
R16344 Iout.n833 Iout.n831 0.00105952
R16345 Iout.n836 Iout.n835 0.00105952
R16346 Iout.n847 Iout.n845 0.00105952
R16347 Iout.n850 Iout.n849 0.00105952
R16348 Iout.n861 Iout.n859 0.00105952
R16349 Iout.n864 Iout.n863 0.00105952
R16350 Iout.n875 Iout.n873 0.00105952
R16351 Iout.n878 Iout.n877 0.00105952
R16352 Iout.n889 Iout.n887 0.00105952
R16353 Iout.n935 Iout.n933 0.00105952
R16354 Iout.n932 Iout.n930 0.00105952
R16355 Iout.n920 Iout.n919 0.00105952
R16356 Iout.n917 Iout.n915 0.00105952
R16357 Iout.n906 Iout.n905 0.00105952
R16358 Iout.n903 Iout.n901 0.00105952
R16359 Iout.n892 Iout.n891 0.00105952
R16360 Iout.n940 Iout.n939 0.00105952
R16361 Iout.n783 Iout.n782 0.00105952
R16362 Iout.n786 Iout.n785 0.00105952
R16363 Iout.n789 Iout.n788 0.00105952
R16364 Iout.n792 Iout.n791 0.00105952
R16365 Iout.n795 Iout.n794 0.00105952
R16366 Iout.n798 Iout.n797 0.00105952
R16367 Iout.n801 Iout.n800 0.00105952
R16368 Iout.n804 Iout.n803 0.00105952
R16369 Iout.n807 Iout.n806 0.00105952
R16370 Iout.n779 Iout.n778 0.00105952
R16371 Iout.n776 Iout.n39 0.00105952
R16372 Iout.n767 Iout.n766 0.00105952
R16373 Iout.n764 Iout.n48 0.00105952
R16374 Iout.n755 Iout.n754 0.00105952
R16375 Iout.n752 Iout.n54 0.00105952
R16376 Iout.n743 Iout.n742 0.00105952
R16377 Iout.n740 Iout.n60 0.00105952
R16378 Iout.n731 Iout.n730 0.00105952
R16379 Iout.n728 Iout.n66 0.00105952
R16380 Iout.n943 Iout.n20 0.00105952
R16381 Iout.n946 Iout.n945 0.00105952
R16382 Iout.n704 Iout.n78 0.00105952
R16383 Iout.n707 Iout.n706 0.00105952
R16384 Iout.n716 Iout.n72 0.00105952
R16385 Iout.n719 Iout.n718 0.00105952
R16386 Iout.n954 Iout.n952 0.00105952
R16387 Iout.n951 Iout.n949 0.00105952
R16388 Iout.n701 Iout.n700 0.00105952
R16389 Iout.n710 Iout.n75 0.00105952
R16390 Iout.n713 Iout.n712 0.00105952
R16391 Iout.n722 Iout.n69 0.00105952
R16392 Iout.n725 Iout.n724 0.00105952
R16393 Iout.n734 Iout.n63 0.00105952
R16394 Iout.n737 Iout.n736 0.00105952
R16395 Iout.n746 Iout.n57 0.00105952
R16396 Iout.n749 Iout.n748 0.00105952
R16397 Iout.n655 Iout.n653 0.00105952
R16398 Iout.n658 Iout.n656 0.00105952
R16399 Iout.n661 Iout.n659 0.00105952
R16400 Iout.n664 Iout.n662 0.00105952
R16401 Iout.n667 Iout.n665 0.00105952
R16402 Iout.n670 Iout.n668 0.00105952
R16403 Iout.n673 Iout.n671 0.00105952
R16404 Iout.n676 Iout.n674 0.00105952
R16405 Iout.n679 Iout.n677 0.00105952
R16406 Iout.n682 Iout.n680 0.00105952
R16407 Iout.n685 Iout.n683 0.00105952
R16408 Iout.n959 Iout.n958 0.00105952
R16409 Iout.n694 Iout.n693 0.00105952
R16410 Iout.n697 Iout.n696 0.00105952
R16411 Iout.n691 Iout.n689 0.00105952
R16412 Iout.n688 Iout.n686 0.00105952
R16413 Iout.n962 Iout.n15 0.00105952
R16414 Iout.n965 Iout.n964 0.00105952
R16415 Iout.n575 Iout.n574 0.00105952
R16416 Iout.n578 Iout.n577 0.00105952
R16417 Iout.n587 Iout.n115 0.00105952
R16418 Iout.n590 Iout.n589 0.00105952
R16419 Iout.n599 Iout.n109 0.00105952
R16420 Iout.n602 Iout.n601 0.00105952
R16421 Iout.n611 Iout.n103 0.00105952
R16422 Iout.n614 Iout.n613 0.00105952
R16423 Iout.n623 Iout.n97 0.00105952
R16424 Iout.n626 Iout.n625 0.00105952
R16425 Iout.n86 Iout.n84 0.00105952
R16426 Iout.n644 Iout.n643 0.00105952
R16427 Iout.n641 Iout.n88 0.00105952
R16428 Iout.n632 Iout.n631 0.00105952
R16429 Iout.n629 Iout.n94 0.00105952
R16430 Iout.n620 Iout.n619 0.00105952
R16431 Iout.n617 Iout.n100 0.00105952
R16432 Iout.n608 Iout.n607 0.00105952
R16433 Iout.n605 Iout.n106 0.00105952
R16434 Iout.n596 Iout.n595 0.00105952
R16435 Iout.n593 Iout.n112 0.00105952
R16436 Iout.n584 Iout.n583 0.00105952
R16437 Iout.n973 Iout.n971 0.00105952
R16438 Iout.n970 Iout.n968 0.00105952
R16439 Iout.n565 Iout.n564 0.00105952
R16440 Iout.n581 Iout.n118 0.00105952
R16441 Iout.n978 Iout.n977 0.00105952
R16442 Iout.n122 Iout.n121 0.00105952
R16443 Iout.n568 Iout.n124 0.00105952
R16444 Iout.n571 Iout.n570 0.00105952
R16445 Iout.n335 Iout.n334 0.00105952
R16446 Iout.n338 Iout.n337 0.00105952
R16447 Iout.n341 Iout.n340 0.00105952
R16448 Iout.n344 Iout.n343 0.00105952
R16449 Iout.n347 Iout.n346 0.00105952
R16450 Iout.n350 Iout.n349 0.00105952
R16451 Iout.n353 Iout.n352 0.00105952
R16452 Iout.n356 Iout.n355 0.00105952
R16453 Iout.n359 Iout.n358 0.00105952
R16454 Iout.n372 Iout.n371 0.00105952
R16455 Iout.n385 Iout.n383 0.00105952
R16456 Iout.n388 Iout.n387 0.00105952
R16457 Iout.n401 Iout.n399 0.00105952
R16458 Iout.n404 Iout.n403 0.00105952
R16459 Iout.n417 Iout.n415 0.00105952
R16460 Iout.n420 Iout.n419 0.00105952
R16461 Iout.n433 Iout.n431 0.00105952
R16462 Iout.n443 Iout.n442 0.00105952
R16463 Iout.n440 Iout.n439 0.00105952
R16464 Iout.n437 Iout.n435 0.00105952
R16465 Iout.n555 Iout.n553 0.00105952
R16466 Iout.n558 Iout.n556 0.00105952
R16467 Iout.n981 Iout.n10 0.00105952
R16468 Iout.n984 Iout.n983 0.00105952
R16469 Iout.n561 Iout.n560 0.00105952
R16470 Iout.n992 Iout.n990 0.00105952
R16471 Iout.n989 Iout.n987 0.00105952
R16472 Iout.n129 Iout.n128 0.00105952
R16473 Iout.n547 Iout.n131 0.00105952
R16474 Iout.n550 Iout.n549 0.00105952
R16475 Iout.n451 Iout.n450 0.00105952
R16476 Iout.n454 Iout.n453 0.00105952
R16477 Iout.n448 Iout.n446 0.00105952
R16478 Iout.n428 Iout.n427 0.00105952
R16479 Iout.n425 Iout.n423 0.00105952
R16480 Iout.n412 Iout.n411 0.00105952
R16481 Iout.n409 Iout.n407 0.00105952
R16482 Iout.n396 Iout.n395 0.00105952
R16483 Iout.n393 Iout.n391 0.00105952
R16484 Iout.n331 Iout.n330 0.00105952
R16485 Iout.n328 Iout.n327 0.00105952
R16486 Iout.n325 Iout.n324 0.00105952
R16487 Iout.n322 Iout.n321 0.00105952
R16488 Iout.n319 Iout.n318 0.00105952
R16489 Iout.n316 Iout.n315 0.00105952
R16490 Iout.n313 Iout.n312 0.00105952
R16491 Iout.n310 Iout.n309 0.00105952
R16492 Iout.n307 Iout.n306 0.00105952
R16493 Iout.n459 Iout.n457 0.00105952
R16494 Iout.n465 Iout.n464 0.00105952
R16495 Iout.n462 Iout.n461 0.00105952
R16496 Iout.n544 Iout.n543 0.00105952
R16497 Iout.n541 Iout.n137 0.00105952
R16498 Iout.n997 Iout.n996 0.00105952
R16499 Iout.n135 Iout.n134 0.00105952
R16500 Iout.n1000 Iout.n5 0.00105952
R16501 Iout.n1003 Iout.n1002 0.00105952
R16502 Iout.n538 Iout.n537 0.00105952
R16503 Iout.n535 Iout.n533 0.00105952
R16504 Iout.n532 Iout.n530 0.00105952
R16505 Iout.n468 Iout.n157 0.00105952
R16506 Iout.n471 Iout.n470 0.00105952
R16507 Iout.n474 Iout.n473 0.00105952
R16508 Iout.n264 Iout.n190 0.00105952
R16509 Iout.n267 Iout.n266 0.00105952
R16510 Iout.n276 Iout.n184 0.00105952
R16511 Iout.n279 Iout.n278 0.00105952
R16512 Iout.n288 Iout.n178 0.00105952
R16513 Iout.n291 Iout.n290 0.00105952
R16514 Iout.n300 Iout.n169 0.00105952
R16515 Iout.n173 Iout.n171 0.00105952
R16516 Iout.n297 Iout.n296 0.00105952
R16517 Iout.n294 Iout.n175 0.00105952
R16518 Iout.n285 Iout.n284 0.00105952
R16519 Iout.n282 Iout.n181 0.00105952
R16520 Iout.n273 Iout.n272 0.00105952
R16521 Iout.n270 Iout.n187 0.00105952
R16522 Iout.n261 Iout.n260 0.00105952
R16523 Iout.n479 Iout.n477 0.00105952
R16524 Iout.n485 Iout.n484 0.00105952
R16525 Iout.n482 Iout.n481 0.00105952
R16526 Iout.n527 Iout.n526 0.00105952
R16527 Iout.n524 Iout.n144 0.00105952
R16528 Iout.n142 Iout.n141 0.00105952
R16529 Iout.n1008 Iout.n1006 0.00105952
R16530 Iout.n1011 Iout.n1009 0.00105952
R16531 Iout.n1016 Iout.n1015 0.00105952
R16532 Iout.n148 Iout.n147 0.00105952
R16533 Iout.n518 Iout.n150 0.00105952
R16534 Iout.n521 Iout.n520 0.00105952
R16535 Iout.n493 Iout.n492 0.00105952
R16536 Iout.n496 Iout.n495 0.00105952
R16537 Iout.n490 Iout.n488 0.00105952
R16538 Iout.n254 Iout.n253 0.00105952
R16539 Iout.n257 Iout.n256 0.00105952
R16540 Iout.n251 Iout.n249 0.00105952
R16541 Iout.n248 Iout.n246 0.00105952
R16542 Iout.n245 Iout.n243 0.00105952
R16543 Iout.n242 Iout.n240 0.00105952
R16544 Iout.n239 Iout.n237 0.00105952
R16545 Iout.n236 Iout.n234 0.00105952
R16546 Iout.n233 Iout.n231 0.00105952
R16547 Iout.n228 Iout.n227 0.00105952
R16548 Iout.n225 Iout.n223 0.00105952
R16549 Iout.n221 Iout.n219 0.00105952
R16550 Iout.n217 Iout.n215 0.00105952
R16551 Iout.n213 Iout.n211 0.00105952
R16552 Iout.n209 Iout.n207 0.00105952
R16553 Iout.n205 Iout.n203 0.00105952
R16554 Iout.n201 Iout.n200 0.00105952
R16555 Iout.n198 Iout.n196 0.00105952
R16556 Iout.n194 Iout.n193 0.00105952
R16557 Iout.n501 Iout.n499 0.00105952
R16558 Iout.n505 Iout.n503 0.00105952
R16559 Iout.n508 Iout.n506 0.00105952
R16560 Iout.n515 Iout.n514 0.00105952
R16561 Iout.n512 Iout.n510 0.00105952
R16562 Iout.n1021 Iout.n1019 0.00105952
R16563 XThC.Tn[10].n55 XThC.Tn[10].n54 256.103
R16564 XThC.Tn[10].n59 XThC.Tn[10].n57 243.68
R16565 XThC.Tn[10].n2 XThC.Tn[10].n0 241.847
R16566 XThC.Tn[10].n59 XThC.Tn[10].n58 205.28
R16567 XThC.Tn[10].n55 XThC.Tn[10].n53 202.095
R16568 XThC.Tn[10].n2 XThC.Tn[10].n1 185
R16569 XThC.Tn[10].n5 XThC.Tn[10].n3 161.406
R16570 XThC.Tn[10].n8 XThC.Tn[10].n6 161.406
R16571 XThC.Tn[10].n11 XThC.Tn[10].n9 161.406
R16572 XThC.Tn[10].n14 XThC.Tn[10].n12 161.406
R16573 XThC.Tn[10].n17 XThC.Tn[10].n15 161.406
R16574 XThC.Tn[10].n20 XThC.Tn[10].n18 161.406
R16575 XThC.Tn[10].n23 XThC.Tn[10].n21 161.406
R16576 XThC.Tn[10].n26 XThC.Tn[10].n24 161.406
R16577 XThC.Tn[10].n29 XThC.Tn[10].n27 161.406
R16578 XThC.Tn[10].n32 XThC.Tn[10].n30 161.406
R16579 XThC.Tn[10].n35 XThC.Tn[10].n33 161.406
R16580 XThC.Tn[10].n38 XThC.Tn[10].n36 161.406
R16581 XThC.Tn[10].n41 XThC.Tn[10].n39 161.406
R16582 XThC.Tn[10].n44 XThC.Tn[10].n42 161.406
R16583 XThC.Tn[10].n47 XThC.Tn[10].n45 161.406
R16584 XThC.Tn[10].n50 XThC.Tn[10].n48 161.406
R16585 XThC.Tn[10].n3 XThC.Tn[10].t36 161.202
R16586 XThC.Tn[10].n6 XThC.Tn[10].t21 161.202
R16587 XThC.Tn[10].n9 XThC.Tn[10].t23 161.202
R16588 XThC.Tn[10].n12 XThC.Tn[10].t25 161.202
R16589 XThC.Tn[10].n15 XThC.Tn[10].t14 161.202
R16590 XThC.Tn[10].n18 XThC.Tn[10].t15 161.202
R16591 XThC.Tn[10].n21 XThC.Tn[10].t28 161.202
R16592 XThC.Tn[10].n24 XThC.Tn[10].t37 161.202
R16593 XThC.Tn[10].n27 XThC.Tn[10].t39 161.202
R16594 XThC.Tn[10].n30 XThC.Tn[10].t26 161.202
R16595 XThC.Tn[10].n33 XThC.Tn[10].t27 161.202
R16596 XThC.Tn[10].n36 XThC.Tn[10].t40 161.202
R16597 XThC.Tn[10].n39 XThC.Tn[10].t16 161.202
R16598 XThC.Tn[10].n42 XThC.Tn[10].t19 161.202
R16599 XThC.Tn[10].n45 XThC.Tn[10].t32 161.202
R16600 XThC.Tn[10].n48 XThC.Tn[10].t42 161.202
R16601 XThC.Tn[10].n3 XThC.Tn[10].t38 145.137
R16602 XThC.Tn[10].n6 XThC.Tn[10].t24 145.137
R16603 XThC.Tn[10].n9 XThC.Tn[10].t29 145.137
R16604 XThC.Tn[10].n12 XThC.Tn[10].t30 145.137
R16605 XThC.Tn[10].n15 XThC.Tn[10].t17 145.137
R16606 XThC.Tn[10].n18 XThC.Tn[10].t18 145.137
R16607 XThC.Tn[10].n21 XThC.Tn[10].t34 145.137
R16608 XThC.Tn[10].n24 XThC.Tn[10].t41 145.137
R16609 XThC.Tn[10].n27 XThC.Tn[10].t43 145.137
R16610 XThC.Tn[10].n30 XThC.Tn[10].t31 145.137
R16611 XThC.Tn[10].n33 XThC.Tn[10].t33 145.137
R16612 XThC.Tn[10].n36 XThC.Tn[10].t12 145.137
R16613 XThC.Tn[10].n39 XThC.Tn[10].t20 145.137
R16614 XThC.Tn[10].n42 XThC.Tn[10].t22 145.137
R16615 XThC.Tn[10].n45 XThC.Tn[10].t35 145.137
R16616 XThC.Tn[10].n48 XThC.Tn[10].t13 145.137
R16617 XThC.Tn[10].n53 XThC.Tn[10].t4 26.5955
R16618 XThC.Tn[10].n53 XThC.Tn[10].t3 26.5955
R16619 XThC.Tn[10].n57 XThC.Tn[10].t11 26.5955
R16620 XThC.Tn[10].n57 XThC.Tn[10].t10 26.5955
R16621 XThC.Tn[10].n58 XThC.Tn[10].t9 26.5955
R16622 XThC.Tn[10].n58 XThC.Tn[10].t8 26.5955
R16623 XThC.Tn[10].n54 XThC.Tn[10].t6 26.5955
R16624 XThC.Tn[10].n54 XThC.Tn[10].t0 26.5955
R16625 XThC.Tn[10].n1 XThC.Tn[10].t7 24.9236
R16626 XThC.Tn[10].n1 XThC.Tn[10].t2 24.9236
R16627 XThC.Tn[10].n0 XThC.Tn[10].t1 24.9236
R16628 XThC.Tn[10].n0 XThC.Tn[10].t5 24.9236
R16629 XThC.Tn[10] XThC.Tn[10].n59 22.9652
R16630 XThC.Tn[10] XThC.Tn[10].n2 22.9615
R16631 XThC.Tn[10].n56 XThC.Tn[10].n55 13.9299
R16632 XThC.Tn[10] XThC.Tn[10].n56 13.9299
R16633 XThC.Tn[10].n52 XThC.Tn[10].n51 5.13256
R16634 XThC.Tn[10].n56 XThC.Tn[10].n52 2.99115
R16635 XThC.Tn[10].n56 XThC.Tn[10] 2.87153
R16636 XThC.Tn[10].n52 XThC.Tn[10] 2.2734
R16637 XThC.Tn[10].n51 XThC.Tn[10] 2.26343
R16638 XThC.Tn[10].n8 XThC.Tn[10] 0.931056
R16639 XThC.Tn[10].n11 XThC.Tn[10] 0.931056
R16640 XThC.Tn[10].n14 XThC.Tn[10] 0.931056
R16641 XThC.Tn[10].n17 XThC.Tn[10] 0.931056
R16642 XThC.Tn[10].n20 XThC.Tn[10] 0.931056
R16643 XThC.Tn[10].n23 XThC.Tn[10] 0.931056
R16644 XThC.Tn[10].n26 XThC.Tn[10] 0.931056
R16645 XThC.Tn[10].n29 XThC.Tn[10] 0.931056
R16646 XThC.Tn[10].n32 XThC.Tn[10] 0.931056
R16647 XThC.Tn[10].n35 XThC.Tn[10] 0.931056
R16648 XThC.Tn[10].n38 XThC.Tn[10] 0.931056
R16649 XThC.Tn[10].n41 XThC.Tn[10] 0.931056
R16650 XThC.Tn[10].n44 XThC.Tn[10] 0.931056
R16651 XThC.Tn[10].n47 XThC.Tn[10] 0.931056
R16652 XThC.Tn[10].n50 XThC.Tn[10] 0.931056
R16653 XThC.Tn[10] XThC.Tn[10].n5 0.396333
R16654 XThC.Tn[10] XThC.Tn[10].n8 0.396333
R16655 XThC.Tn[10] XThC.Tn[10].n11 0.396333
R16656 XThC.Tn[10] XThC.Tn[10].n14 0.396333
R16657 XThC.Tn[10] XThC.Tn[10].n17 0.396333
R16658 XThC.Tn[10] XThC.Tn[10].n20 0.396333
R16659 XThC.Tn[10] XThC.Tn[10].n23 0.396333
R16660 XThC.Tn[10] XThC.Tn[10].n26 0.396333
R16661 XThC.Tn[10] XThC.Tn[10].n29 0.396333
R16662 XThC.Tn[10] XThC.Tn[10].n32 0.396333
R16663 XThC.Tn[10] XThC.Tn[10].n35 0.396333
R16664 XThC.Tn[10] XThC.Tn[10].n38 0.396333
R16665 XThC.Tn[10] XThC.Tn[10].n41 0.396333
R16666 XThC.Tn[10] XThC.Tn[10].n44 0.396333
R16667 XThC.Tn[10] XThC.Tn[10].n47 0.396333
R16668 XThC.Tn[10] XThC.Tn[10].n50 0.396333
R16669 XThC.Tn[10].n4 XThC.Tn[10] 0.104667
R16670 XThC.Tn[10].n7 XThC.Tn[10] 0.104667
R16671 XThC.Tn[10].n10 XThC.Tn[10] 0.104667
R16672 XThC.Tn[10].n13 XThC.Tn[10] 0.104667
R16673 XThC.Tn[10].n16 XThC.Tn[10] 0.104667
R16674 XThC.Tn[10].n19 XThC.Tn[10] 0.104667
R16675 XThC.Tn[10].n22 XThC.Tn[10] 0.104667
R16676 XThC.Tn[10].n25 XThC.Tn[10] 0.104667
R16677 XThC.Tn[10].n28 XThC.Tn[10] 0.104667
R16678 XThC.Tn[10].n31 XThC.Tn[10] 0.104667
R16679 XThC.Tn[10].n34 XThC.Tn[10] 0.104667
R16680 XThC.Tn[10].n37 XThC.Tn[10] 0.104667
R16681 XThC.Tn[10].n40 XThC.Tn[10] 0.104667
R16682 XThC.Tn[10].n43 XThC.Tn[10] 0.104667
R16683 XThC.Tn[10].n46 XThC.Tn[10] 0.104667
R16684 XThC.Tn[10].n49 XThC.Tn[10] 0.104667
R16685 XThC.Tn[10].n4 XThC.Tn[10] 0.0309878
R16686 XThC.Tn[10].n7 XThC.Tn[10] 0.0309878
R16687 XThC.Tn[10].n10 XThC.Tn[10] 0.0309878
R16688 XThC.Tn[10].n13 XThC.Tn[10] 0.0309878
R16689 XThC.Tn[10].n16 XThC.Tn[10] 0.0309878
R16690 XThC.Tn[10].n19 XThC.Tn[10] 0.0309878
R16691 XThC.Tn[10].n22 XThC.Tn[10] 0.0309878
R16692 XThC.Tn[10].n25 XThC.Tn[10] 0.0309878
R16693 XThC.Tn[10].n28 XThC.Tn[10] 0.0309878
R16694 XThC.Tn[10].n31 XThC.Tn[10] 0.0309878
R16695 XThC.Tn[10].n34 XThC.Tn[10] 0.0309878
R16696 XThC.Tn[10].n37 XThC.Tn[10] 0.0309878
R16697 XThC.Tn[10].n40 XThC.Tn[10] 0.0309878
R16698 XThC.Tn[10].n43 XThC.Tn[10] 0.0309878
R16699 XThC.Tn[10].n46 XThC.Tn[10] 0.0309878
R16700 XThC.Tn[10].n49 XThC.Tn[10] 0.0309878
R16701 XThC.Tn[10].n5 XThC.Tn[10].n4 0.027939
R16702 XThC.Tn[10].n8 XThC.Tn[10].n7 0.027939
R16703 XThC.Tn[10].n11 XThC.Tn[10].n10 0.027939
R16704 XThC.Tn[10].n14 XThC.Tn[10].n13 0.027939
R16705 XThC.Tn[10].n17 XThC.Tn[10].n16 0.027939
R16706 XThC.Tn[10].n20 XThC.Tn[10].n19 0.027939
R16707 XThC.Tn[10].n23 XThC.Tn[10].n22 0.027939
R16708 XThC.Tn[10].n26 XThC.Tn[10].n25 0.027939
R16709 XThC.Tn[10].n29 XThC.Tn[10].n28 0.027939
R16710 XThC.Tn[10].n32 XThC.Tn[10].n31 0.027939
R16711 XThC.Tn[10].n35 XThC.Tn[10].n34 0.027939
R16712 XThC.Tn[10].n38 XThC.Tn[10].n37 0.027939
R16713 XThC.Tn[10].n41 XThC.Tn[10].n40 0.027939
R16714 XThC.Tn[10].n44 XThC.Tn[10].n43 0.027939
R16715 XThC.Tn[10].n47 XThC.Tn[10].n46 0.027939
R16716 XThC.Tn[10].n50 XThC.Tn[10].n49 0.027939
R16717 XThC.Tn[10].n51 XThC.Tn[10] 0.00285068
R16718 XThR.XTBN.Y.n1 XThR.XTBN.Y.t60 212.081
R16719 XThR.XTBN.Y.n8 XThR.XTBN.Y.t12 212.081
R16720 XThR.XTBN.Y.n2 XThR.XTBN.Y.t81 212.081
R16721 XThR.XTBN.Y.n3 XThR.XTBN.Y.t121 212.081
R16722 XThR.XTBN.Y.n12 XThR.XTBN.Y.t115 212.081
R16723 XThR.XTBN.Y.n19 XThR.XTBN.Y.t65 212.081
R16724 XThR.XTBN.Y.n13 XThR.XTBN.Y.t21 212.081
R16725 XThR.XTBN.Y.n14 XThR.XTBN.Y.t57 212.081
R16726 XThR.XTBN.Y.n24 XThR.XTBN.Y.t27 212.081
R16727 XThR.XTBN.Y.n31 XThR.XTBN.Y.t96 212.081
R16728 XThR.XTBN.Y.n25 XThR.XTBN.Y.t46 212.081
R16729 XThR.XTBN.Y.n26 XThR.XTBN.Y.t89 212.081
R16730 XThR.XTBN.Y.n36 XThR.XTBN.Y.t80 212.081
R16731 XThR.XTBN.Y.n43 XThR.XTBN.Y.t31 212.081
R16732 XThR.XTBN.Y.n37 XThR.XTBN.Y.t102 212.081
R16733 XThR.XTBN.Y.n38 XThR.XTBN.Y.t25 212.081
R16734 XThR.XTBN.Y.n48 XThR.XTBN.Y.t85 212.081
R16735 XThR.XTBN.Y.n55 XThR.XTBN.Y.t33 212.081
R16736 XThR.XTBN.Y.n49 XThR.XTBN.Y.t105 212.081
R16737 XThR.XTBN.Y.n50 XThR.XTBN.Y.t26 212.081
R16738 XThR.XTBN.Y.n60 XThR.XTBN.Y.t54 212.081
R16739 XThR.XTBN.Y.n67 XThR.XTBN.Y.t5 212.081
R16740 XThR.XTBN.Y.n61 XThR.XTBN.Y.t73 212.081
R16741 XThR.XTBN.Y.n62 XThR.XTBN.Y.t114 212.081
R16742 XThR.XTBN.Y.n72 XThR.XTBN.Y.t49 212.081
R16743 XThR.XTBN.Y.n79 XThR.XTBN.Y.t119 212.081
R16744 XThR.XTBN.Y.n73 XThR.XTBN.Y.t69 212.081
R16745 XThR.XTBN.Y.n74 XThR.XTBN.Y.t108 212.081
R16746 XThR.XTBN.Y.n163 XThR.XTBN.Y.t41 212.081
R16747 XThR.XTBN.Y.n154 XThR.XTBN.Y.t113 212.081
R16748 XThR.XTBN.Y.n158 XThR.XTBN.Y.t34 212.081
R16749 XThR.XTBN.Y.n155 XThR.XTBN.Y.t72 212.081
R16750 XThR.XTBN.Y.n151 XThR.XTBN.Y.t19 212.081
R16751 XThR.XTBN.Y.n142 XThR.XTBN.Y.t86 212.081
R16752 XThR.XTBN.Y.n146 XThR.XTBN.Y.t6 212.081
R16753 XThR.XTBN.Y.n143 XThR.XTBN.Y.t43 212.081
R16754 XThR.XTBN.Y.n139 XThR.XTBN.Y.t45 212.081
R16755 XThR.XTBN.Y.n130 XThR.XTBN.Y.t117 212.081
R16756 XThR.XTBN.Y.n134 XThR.XTBN.Y.t36 212.081
R16757 XThR.XTBN.Y.n131 XThR.XTBN.Y.t75 212.081
R16758 XThR.XTBN.Y.n127 XThR.XTBN.Y.t100 212.081
R16759 XThR.XTBN.Y.n118 XThR.XTBN.Y.t50 212.081
R16760 XThR.XTBN.Y.n122 XThR.XTBN.Y.t92 212.081
R16761 XThR.XTBN.Y.n119 XThR.XTBN.Y.t13 212.081
R16762 XThR.XTBN.Y.n115 XThR.XTBN.Y.t15 212.081
R16763 XThR.XTBN.Y.n106 XThR.XTBN.Y.t83 212.081
R16764 XThR.XTBN.Y.n110 XThR.XTBN.Y.t123 212.081
R16765 XThR.XTBN.Y.n107 XThR.XTBN.Y.t39 212.081
R16766 XThR.XTBN.Y.n103 XThR.XTBN.Y.t66 212.081
R16767 XThR.XTBN.Y.n94 XThR.XTBN.Y.t23 212.081
R16768 XThR.XTBN.Y.n98 XThR.XTBN.Y.t59 212.081
R16769 XThR.XTBN.Y.n95 XThR.XTBN.Y.t97 212.081
R16770 XThR.XTBN.Y.n92 XThR.XTBN.Y.t99 212.081
R16771 XThR.XTBN.Y.n83 XThR.XTBN.Y.t87 212.081
R16772 XThR.XTBN.Y.n87 XThR.XTBN.Y.t77 212.081
R16773 XThR.XTBN.Y.n84 XThR.XTBN.Y.t68 212.081
R16774 XThR.XTBN.Y.n167 XThR.XTBN.Y.t63 212.081
R16775 XThR.XTBN.Y.n169 XThR.XTBN.Y.t106 212.081
R16776 XThR.XTBN.Y.n174 XThR.XTBN.Y.t56 212.081
R16777 XThR.XTBN.Y.n170 XThR.XTBN.Y.t7 212.081
R16778 XThR.XTBN.Y XThR.XTBN.Y.n180 203.923
R16779 XThR.XTBN.Y.n171 XThR.XTBN.Y.n170 188.516
R16780 XThR.XTBN.Y.n164 XThR.XTBN.Y.n163 180.482
R16781 XThR.XTBN.Y.n152 XThR.XTBN.Y.n151 180.482
R16782 XThR.XTBN.Y.n140 XThR.XTBN.Y.n139 180.482
R16783 XThR.XTBN.Y.n128 XThR.XTBN.Y.n127 180.482
R16784 XThR.XTBN.Y.n116 XThR.XTBN.Y.n115 180.482
R16785 XThR.XTBN.Y.n104 XThR.XTBN.Y.n103 180.482
R16786 XThR.XTBN.Y.n93 XThR.XTBN.Y.n92 180.482
R16787 XThR.XTBN.Y.n5 XThR.XTBN.Y.n4 173.761
R16788 XThR.XTBN.Y.n16 XThR.XTBN.Y.n15 173.761
R16789 XThR.XTBN.Y.n28 XThR.XTBN.Y.n27 173.761
R16790 XThR.XTBN.Y.n40 XThR.XTBN.Y.n39 173.761
R16791 XThR.XTBN.Y.n52 XThR.XTBN.Y.n51 173.761
R16792 XThR.XTBN.Y.n64 XThR.XTBN.Y.n63 173.761
R16793 XThR.XTBN.Y.n76 XThR.XTBN.Y.n75 173.761
R16794 XThR.XTBN.Y.n168 XThR.XTBN.Y 154.304
R16795 XThR.XTBN.Y.n10 XThR.XTBN.Y.n9 152
R16796 XThR.XTBN.Y.n7 XThR.XTBN.Y.n0 152
R16797 XThR.XTBN.Y.n6 XThR.XTBN.Y.n5 152
R16798 XThR.XTBN.Y.n17 XThR.XTBN.Y.n16 152
R16799 XThR.XTBN.Y.n18 XThR.XTBN.Y.n11 152
R16800 XThR.XTBN.Y.n21 XThR.XTBN.Y.n20 152
R16801 XThR.XTBN.Y.n29 XThR.XTBN.Y.n28 152
R16802 XThR.XTBN.Y.n30 XThR.XTBN.Y.n23 152
R16803 XThR.XTBN.Y.n33 XThR.XTBN.Y.n32 152
R16804 XThR.XTBN.Y.n41 XThR.XTBN.Y.n40 152
R16805 XThR.XTBN.Y.n42 XThR.XTBN.Y.n35 152
R16806 XThR.XTBN.Y.n45 XThR.XTBN.Y.n44 152
R16807 XThR.XTBN.Y.n53 XThR.XTBN.Y.n52 152
R16808 XThR.XTBN.Y.n54 XThR.XTBN.Y.n47 152
R16809 XThR.XTBN.Y.n57 XThR.XTBN.Y.n56 152
R16810 XThR.XTBN.Y.n65 XThR.XTBN.Y.n64 152
R16811 XThR.XTBN.Y.n66 XThR.XTBN.Y.n59 152
R16812 XThR.XTBN.Y.n69 XThR.XTBN.Y.n68 152
R16813 XThR.XTBN.Y.n77 XThR.XTBN.Y.n76 152
R16814 XThR.XTBN.Y.n78 XThR.XTBN.Y.n71 152
R16815 XThR.XTBN.Y.n81 XThR.XTBN.Y.n80 152
R16816 XThR.XTBN.Y.n157 XThR.XTBN.Y.n156 152
R16817 XThR.XTBN.Y.n160 XThR.XTBN.Y.n159 152
R16818 XThR.XTBN.Y.n162 XThR.XTBN.Y.n161 152
R16819 XThR.XTBN.Y.n145 XThR.XTBN.Y.n144 152
R16820 XThR.XTBN.Y.n148 XThR.XTBN.Y.n147 152
R16821 XThR.XTBN.Y.n150 XThR.XTBN.Y.n149 152
R16822 XThR.XTBN.Y.n133 XThR.XTBN.Y.n132 152
R16823 XThR.XTBN.Y.n136 XThR.XTBN.Y.n135 152
R16824 XThR.XTBN.Y.n138 XThR.XTBN.Y.n137 152
R16825 XThR.XTBN.Y.n121 XThR.XTBN.Y.n120 152
R16826 XThR.XTBN.Y.n124 XThR.XTBN.Y.n123 152
R16827 XThR.XTBN.Y.n126 XThR.XTBN.Y.n125 152
R16828 XThR.XTBN.Y.n109 XThR.XTBN.Y.n108 152
R16829 XThR.XTBN.Y.n112 XThR.XTBN.Y.n111 152
R16830 XThR.XTBN.Y.n114 XThR.XTBN.Y.n113 152
R16831 XThR.XTBN.Y.n97 XThR.XTBN.Y.n96 152
R16832 XThR.XTBN.Y.n100 XThR.XTBN.Y.n99 152
R16833 XThR.XTBN.Y.n102 XThR.XTBN.Y.n101 152
R16834 XThR.XTBN.Y.n86 XThR.XTBN.Y.n85 152
R16835 XThR.XTBN.Y.n89 XThR.XTBN.Y.n88 152
R16836 XThR.XTBN.Y.n91 XThR.XTBN.Y.n90 152
R16837 XThR.XTBN.Y.n173 XThR.XTBN.Y.n172 152
R16838 XThR.XTBN.Y.n176 XThR.XTBN.Y.n175 152
R16839 XThR.XTBN.Y.n1 XThR.XTBN.Y.t95 139.78
R16840 XThR.XTBN.Y.n8 XThR.XTBN.Y.t44 139.78
R16841 XThR.XTBN.Y.n2 XThR.XTBN.Y.t116 139.78
R16842 XThR.XTBN.Y.n3 XThR.XTBN.Y.t35 139.78
R16843 XThR.XTBN.Y.n12 XThR.XTBN.Y.t42 139.78
R16844 XThR.XTBN.Y.n19 XThR.XTBN.Y.t112 139.78
R16845 XThR.XTBN.Y.n13 XThR.XTBN.Y.t64 139.78
R16846 XThR.XTBN.Y.n14 XThR.XTBN.Y.t107 139.78
R16847 XThR.XTBN.Y.n24 XThR.XTBN.Y.t61 139.78
R16848 XThR.XTBN.Y.n31 XThR.XTBN.Y.t14 139.78
R16849 XThR.XTBN.Y.n25 XThR.XTBN.Y.t82 139.78
R16850 XThR.XTBN.Y.n26 XThR.XTBN.Y.t122 139.78
R16851 XThR.XTBN.Y.n36 XThR.XTBN.Y.t11 139.78
R16852 XThR.XTBN.Y.n43 XThR.XTBN.Y.t79 139.78
R16853 XThR.XTBN.Y.n37 XThR.XTBN.Y.t32 139.78
R16854 XThR.XTBN.Y.n38 XThR.XTBN.Y.t71 139.78
R16855 XThR.XTBN.Y.n48 XThR.XTBN.Y.t29 139.78
R16856 XThR.XTBN.Y.n55 XThR.XTBN.Y.t98 139.78
R16857 XThR.XTBN.Y.n49 XThR.XTBN.Y.t47 139.78
R16858 XThR.XTBN.Y.n50 XThR.XTBN.Y.t90 139.78
R16859 XThR.XTBN.Y.n60 XThR.XTBN.Y.t8 139.78
R16860 XThR.XTBN.Y.n67 XThR.XTBN.Y.t74 139.78
R16861 XThR.XTBN.Y.n61 XThR.XTBN.Y.t28 139.78
R16862 XThR.XTBN.Y.n62 XThR.XTBN.Y.t67 139.78
R16863 XThR.XTBN.Y.n72 XThR.XTBN.Y.t111 139.78
R16864 XThR.XTBN.Y.n79 XThR.XTBN.Y.t62 139.78
R16865 XThR.XTBN.Y.n73 XThR.XTBN.Y.t18 139.78
R16866 XThR.XTBN.Y.n74 XThR.XTBN.Y.t53 139.78
R16867 XThR.XTBN.Y.n163 XThR.XTBN.Y.t101 139.78
R16868 XThR.XTBN.Y.n154 XThR.XTBN.Y.t52 139.78
R16869 XThR.XTBN.Y.n158 XThR.XTBN.Y.t93 139.78
R16870 XThR.XTBN.Y.n155 XThR.XTBN.Y.t16 139.78
R16871 XThR.XTBN.Y.n151 XThR.XTBN.Y.t88 139.78
R16872 XThR.XTBN.Y.n142 XThR.XTBN.Y.t37 139.78
R16873 XThR.XTBN.Y.n146 XThR.XTBN.Y.t76 139.78
R16874 XThR.XTBN.Y.n143 XThR.XTBN.Y.t118 139.78
R16875 XThR.XTBN.Y.n139 XThR.XTBN.Y.t104 139.78
R16876 XThR.XTBN.Y.n130 XThR.XTBN.Y.t55 139.78
R16877 XThR.XTBN.Y.n134 XThR.XTBN.Y.t94 139.78
R16878 XThR.XTBN.Y.n131 XThR.XTBN.Y.t17 139.78
R16879 XThR.XTBN.Y.n127 XThR.XTBN.Y.t51 139.78
R16880 XThR.XTBN.Y.n118 XThR.XTBN.Y.t4 139.78
R16881 XThR.XTBN.Y.n122 XThR.XTBN.Y.t40 139.78
R16882 XThR.XTBN.Y.n119 XThR.XTBN.Y.t84 139.78
R16883 XThR.XTBN.Y.n115 XThR.XTBN.Y.t38 139.78
R16884 XThR.XTBN.Y.n106 XThR.XTBN.Y.t109 139.78
R16885 XThR.XTBN.Y.n110 XThR.XTBN.Y.t30 139.78
R16886 XThR.XTBN.Y.n107 XThR.XTBN.Y.t70 139.78
R16887 XThR.XTBN.Y.n103 XThR.XTBN.Y.t24 139.78
R16888 XThR.XTBN.Y.n94 XThR.XTBN.Y.t91 139.78
R16889 XThR.XTBN.Y.n98 XThR.XTBN.Y.t10 139.78
R16890 XThR.XTBN.Y.n95 XThR.XTBN.Y.t48 139.78
R16891 XThR.XTBN.Y.n92 XThR.XTBN.Y.t20 139.78
R16892 XThR.XTBN.Y.n83 XThR.XTBN.Y.t120 139.78
R16893 XThR.XTBN.Y.n87 XThR.XTBN.Y.t110 139.78
R16894 XThR.XTBN.Y.n84 XThR.XTBN.Y.t103 139.78
R16895 XThR.XTBN.Y.n167 XThR.XTBN.Y.t22 139.78
R16896 XThR.XTBN.Y.n169 XThR.XTBN.Y.t58 139.78
R16897 XThR.XTBN.Y.n174 XThR.XTBN.Y.t9 139.78
R16898 XThR.XTBN.Y.n170 XThR.XTBN.Y.t78 139.78
R16899 XThR.XTBN.Y.n184 XThR.XTBN.Y.n183 101.489
R16900 XThR.XTBN.Y.n179 XThR.XTBN.Y 58.2909
R16901 XThR.XTBN.Y.n7 XThR.XTBN.Y.n6 49.6611
R16902 XThR.XTBN.Y.n18 XThR.XTBN.Y.n17 49.6611
R16903 XThR.XTBN.Y.n30 XThR.XTBN.Y.n29 49.6611
R16904 XThR.XTBN.Y.n42 XThR.XTBN.Y.n41 49.6611
R16905 XThR.XTBN.Y.n54 XThR.XTBN.Y.n53 49.6611
R16906 XThR.XTBN.Y.n66 XThR.XTBN.Y.n65 49.6611
R16907 XThR.XTBN.Y.n78 XThR.XTBN.Y.n77 49.6611
R16908 XThR.XTBN.Y.n9 XThR.XTBN.Y.n8 44.549
R16909 XThR.XTBN.Y.n20 XThR.XTBN.Y.n19 44.549
R16910 XThR.XTBN.Y.n32 XThR.XTBN.Y.n31 44.549
R16911 XThR.XTBN.Y.n44 XThR.XTBN.Y.n43 44.549
R16912 XThR.XTBN.Y.n56 XThR.XTBN.Y.n55 44.549
R16913 XThR.XTBN.Y.n68 XThR.XTBN.Y.n67 44.549
R16914 XThR.XTBN.Y.n80 XThR.XTBN.Y.n79 44.549
R16915 XThR.XTBN.Y.n4 XThR.XTBN.Y.n2 43.0884
R16916 XThR.XTBN.Y.n15 XThR.XTBN.Y.n13 43.0884
R16917 XThR.XTBN.Y.n27 XThR.XTBN.Y.n25 43.0884
R16918 XThR.XTBN.Y.n39 XThR.XTBN.Y.n37 43.0884
R16919 XThR.XTBN.Y.n51 XThR.XTBN.Y.n49 43.0884
R16920 XThR.XTBN.Y.n63 XThR.XTBN.Y.n61 43.0884
R16921 XThR.XTBN.Y.n75 XThR.XTBN.Y.n73 43.0884
R16922 XThR.XTBN.Y.n163 XThR.XTBN.Y.n162 30.6732
R16923 XThR.XTBN.Y.n162 XThR.XTBN.Y.n154 30.6732
R16924 XThR.XTBN.Y.n159 XThR.XTBN.Y.n154 30.6732
R16925 XThR.XTBN.Y.n159 XThR.XTBN.Y.n158 30.6732
R16926 XThR.XTBN.Y.n158 XThR.XTBN.Y.n157 30.6732
R16927 XThR.XTBN.Y.n157 XThR.XTBN.Y.n155 30.6732
R16928 XThR.XTBN.Y.n151 XThR.XTBN.Y.n150 30.6732
R16929 XThR.XTBN.Y.n150 XThR.XTBN.Y.n142 30.6732
R16930 XThR.XTBN.Y.n147 XThR.XTBN.Y.n142 30.6732
R16931 XThR.XTBN.Y.n147 XThR.XTBN.Y.n146 30.6732
R16932 XThR.XTBN.Y.n146 XThR.XTBN.Y.n145 30.6732
R16933 XThR.XTBN.Y.n145 XThR.XTBN.Y.n143 30.6732
R16934 XThR.XTBN.Y.n139 XThR.XTBN.Y.n138 30.6732
R16935 XThR.XTBN.Y.n138 XThR.XTBN.Y.n130 30.6732
R16936 XThR.XTBN.Y.n135 XThR.XTBN.Y.n130 30.6732
R16937 XThR.XTBN.Y.n135 XThR.XTBN.Y.n134 30.6732
R16938 XThR.XTBN.Y.n134 XThR.XTBN.Y.n133 30.6732
R16939 XThR.XTBN.Y.n133 XThR.XTBN.Y.n131 30.6732
R16940 XThR.XTBN.Y.n127 XThR.XTBN.Y.n126 30.6732
R16941 XThR.XTBN.Y.n126 XThR.XTBN.Y.n118 30.6732
R16942 XThR.XTBN.Y.n123 XThR.XTBN.Y.n118 30.6732
R16943 XThR.XTBN.Y.n123 XThR.XTBN.Y.n122 30.6732
R16944 XThR.XTBN.Y.n122 XThR.XTBN.Y.n121 30.6732
R16945 XThR.XTBN.Y.n121 XThR.XTBN.Y.n119 30.6732
R16946 XThR.XTBN.Y.n115 XThR.XTBN.Y.n114 30.6732
R16947 XThR.XTBN.Y.n114 XThR.XTBN.Y.n106 30.6732
R16948 XThR.XTBN.Y.n111 XThR.XTBN.Y.n106 30.6732
R16949 XThR.XTBN.Y.n111 XThR.XTBN.Y.n110 30.6732
R16950 XThR.XTBN.Y.n110 XThR.XTBN.Y.n109 30.6732
R16951 XThR.XTBN.Y.n109 XThR.XTBN.Y.n107 30.6732
R16952 XThR.XTBN.Y.n103 XThR.XTBN.Y.n102 30.6732
R16953 XThR.XTBN.Y.n102 XThR.XTBN.Y.n94 30.6732
R16954 XThR.XTBN.Y.n99 XThR.XTBN.Y.n94 30.6732
R16955 XThR.XTBN.Y.n99 XThR.XTBN.Y.n98 30.6732
R16956 XThR.XTBN.Y.n98 XThR.XTBN.Y.n97 30.6732
R16957 XThR.XTBN.Y.n97 XThR.XTBN.Y.n95 30.6732
R16958 XThR.XTBN.Y.n92 XThR.XTBN.Y.n91 30.6732
R16959 XThR.XTBN.Y.n91 XThR.XTBN.Y.n83 30.6732
R16960 XThR.XTBN.Y.n88 XThR.XTBN.Y.n83 30.6732
R16961 XThR.XTBN.Y.n88 XThR.XTBN.Y.n87 30.6732
R16962 XThR.XTBN.Y.n87 XThR.XTBN.Y.n86 30.6732
R16963 XThR.XTBN.Y.n86 XThR.XTBN.Y.n84 30.6732
R16964 XThR.XTBN.Y.n168 XThR.XTBN.Y.n167 30.6732
R16965 XThR.XTBN.Y.n169 XThR.XTBN.Y.n168 30.6732
R16966 XThR.XTBN.Y.n175 XThR.XTBN.Y.n169 30.6732
R16967 XThR.XTBN.Y.n175 XThR.XTBN.Y.n174 30.6732
R16968 XThR.XTBN.Y.n174 XThR.XTBN.Y.n173 30.6732
R16969 XThR.XTBN.Y.n173 XThR.XTBN.Y.n170 30.6732
R16970 XThR.XTBN.Y.n180 XThR.XTBN.Y.t3 26.5955
R16971 XThR.XTBN.Y.n180 XThR.XTBN.Y.t2 26.5955
R16972 XThR.XTBN.Y.n183 XThR.XTBN.Y.t0 24.9236
R16973 XThR.XTBN.Y.n183 XThR.XTBN.Y.t1 24.9236
R16974 XThR.XTBN.Y.n10 XThR.XTBN.Y.n0 21.7605
R16975 XThR.XTBN.Y.n21 XThR.XTBN.Y.n11 21.7605
R16976 XThR.XTBN.Y.n33 XThR.XTBN.Y.n23 21.7605
R16977 XThR.XTBN.Y.n45 XThR.XTBN.Y.n35 21.7605
R16978 XThR.XTBN.Y.n57 XThR.XTBN.Y.n47 21.7605
R16979 XThR.XTBN.Y.n69 XThR.XTBN.Y.n59 21.7605
R16980 XThR.XTBN.Y.n81 XThR.XTBN.Y.n71 21.7605
R16981 XThR.XTBN.Y.n161 XThR.XTBN.Y 18.4325
R16982 XThR.XTBN.Y.n149 XThR.XTBN.Y 18.4325
R16983 XThR.XTBN.Y.n137 XThR.XTBN.Y 18.4325
R16984 XThR.XTBN.Y.n125 XThR.XTBN.Y 18.4325
R16985 XThR.XTBN.Y.n113 XThR.XTBN.Y 18.4325
R16986 XThR.XTBN.Y.n101 XThR.XTBN.Y 18.4325
R16987 XThR.XTBN.Y.n90 XThR.XTBN.Y 18.4325
R16988 XThR.XTBN.Y.n4 XThR.XTBN.Y.n3 18.2581
R16989 XThR.XTBN.Y.n15 XThR.XTBN.Y.n14 18.2581
R16990 XThR.XTBN.Y.n27 XThR.XTBN.Y.n26 18.2581
R16991 XThR.XTBN.Y.n39 XThR.XTBN.Y.n38 18.2581
R16992 XThR.XTBN.Y.n51 XThR.XTBN.Y.n50 18.2581
R16993 XThR.XTBN.Y.n63 XThR.XTBN.Y.n62 18.2581
R16994 XThR.XTBN.Y.n75 XThR.XTBN.Y.n74 18.2581
R16995 XThR.XTBN.Y.n5 XThR.XTBN.Y 17.6005
R16996 XThR.XTBN.Y.n16 XThR.XTBN.Y 17.6005
R16997 XThR.XTBN.Y.n28 XThR.XTBN.Y 17.6005
R16998 XThR.XTBN.Y.n40 XThR.XTBN.Y 17.6005
R16999 XThR.XTBN.Y.n52 XThR.XTBN.Y 17.6005
R17000 XThR.XTBN.Y.n64 XThR.XTBN.Y 17.6005
R17001 XThR.XTBN.Y.n76 XThR.XTBN.Y 17.6005
R17002 XThR.XTBN.Y.n22 XThR.XTBN.Y.n10 17.1655
R17003 XThR.XTBN.Y.n172 XThR.XTBN.Y 17.1525
R17004 XThR.XTBN.Y XThR.XTBN.Y.n171 17.1525
R17005 XThR.XTBN.Y.n105 XThR.XTBN.Y.n93 17.054
R17006 XThR.XTBN.Y.n9 XThR.XTBN.Y.n1 16.7975
R17007 XThR.XTBN.Y.n20 XThR.XTBN.Y.n12 16.7975
R17008 XThR.XTBN.Y.n32 XThR.XTBN.Y.n24 16.7975
R17009 XThR.XTBN.Y.n44 XThR.XTBN.Y.n36 16.7975
R17010 XThR.XTBN.Y.n56 XThR.XTBN.Y.n48 16.7975
R17011 XThR.XTBN.Y.n68 XThR.XTBN.Y.n60 16.7975
R17012 XThR.XTBN.Y.n80 XThR.XTBN.Y.n72 16.7975
R17013 XThR.XTBN.Y XThR.XTBN.Y.n160 16.3845
R17014 XThR.XTBN.Y XThR.XTBN.Y.n148 16.3845
R17015 XThR.XTBN.Y XThR.XTBN.Y.n136 16.3845
R17016 XThR.XTBN.Y XThR.XTBN.Y.n124 16.3845
R17017 XThR.XTBN.Y XThR.XTBN.Y.n112 16.3845
R17018 XThR.XTBN.Y XThR.XTBN.Y.n100 16.3845
R17019 XThR.XTBN.Y XThR.XTBN.Y.n89 16.3845
R17020 XThR.XTBN.Y.n22 XThR.XTBN.Y.n21 16.0405
R17021 XThR.XTBN.Y.n34 XThR.XTBN.Y.n33 16.0405
R17022 XThR.XTBN.Y.n46 XThR.XTBN.Y.n45 16.0405
R17023 XThR.XTBN.Y.n58 XThR.XTBN.Y.n57 16.0405
R17024 XThR.XTBN.Y.n70 XThR.XTBN.Y.n69 16.0405
R17025 XThR.XTBN.Y.n82 XThR.XTBN.Y.n81 16.0405
R17026 XThR.XTBN.Y.n165 XThR.XTBN.Y.n164 15.5925
R17027 XThR.XTBN.Y.n153 XThR.XTBN.Y.n152 15.5925
R17028 XThR.XTBN.Y.n141 XThR.XTBN.Y.n140 15.5925
R17029 XThR.XTBN.Y.n129 XThR.XTBN.Y.n128 15.5925
R17030 XThR.XTBN.Y.n117 XThR.XTBN.Y.n116 15.5925
R17031 XThR.XTBN.Y.n105 XThR.XTBN.Y.n104 15.5925
R17032 XThR.XTBN.Y.n156 XThR.XTBN.Y 14.3365
R17033 XThR.XTBN.Y.n144 XThR.XTBN.Y 14.3365
R17034 XThR.XTBN.Y.n132 XThR.XTBN.Y 14.3365
R17035 XThR.XTBN.Y.n120 XThR.XTBN.Y 14.3365
R17036 XThR.XTBN.Y.n108 XThR.XTBN.Y 14.3365
R17037 XThR.XTBN.Y.n96 XThR.XTBN.Y 14.3365
R17038 XThR.XTBN.Y.n85 XThR.XTBN.Y 14.3365
R17039 XThR.XTBN.Y XThR.XTBN.Y.n182 13.5685
R17040 XThR.XTBN.Y.n177 XThR.XTBN.Y.n176 12.2885
R17041 XThR.XTBN.Y XThR.XTBN.Y.n181 10.7525
R17042 XThR.XTBN.Y.n156 XThR.XTBN.Y 9.2165
R17043 XThR.XTBN.Y.n144 XThR.XTBN.Y 9.2165
R17044 XThR.XTBN.Y.n132 XThR.XTBN.Y 9.2165
R17045 XThR.XTBN.Y.n120 XThR.XTBN.Y 9.2165
R17046 XThR.XTBN.Y.n108 XThR.XTBN.Y 9.2165
R17047 XThR.XTBN.Y.n96 XThR.XTBN.Y 9.2165
R17048 XThR.XTBN.Y.n85 XThR.XTBN.Y 9.2165
R17049 XThR.XTBN.Y.n160 XThR.XTBN.Y 7.1685
R17050 XThR.XTBN.Y.n148 XThR.XTBN.Y 7.1685
R17051 XThR.XTBN.Y.n136 XThR.XTBN.Y 7.1685
R17052 XThR.XTBN.Y.n124 XThR.XTBN.Y 7.1685
R17053 XThR.XTBN.Y.n112 XThR.XTBN.Y 7.1685
R17054 XThR.XTBN.Y.n100 XThR.XTBN.Y 7.1685
R17055 XThR.XTBN.Y.n89 XThR.XTBN.Y 7.1685
R17056 XThR.XTBN.Y.n177 XThR.XTBN.Y 6.9125
R17057 XThR.XTBN.Y.n181 XThR.XTBN.Y 6.6565
R17058 XThR.XTBN.Y.n6 XThR.XTBN.Y.n2 6.57323
R17059 XThR.XTBN.Y.n17 XThR.XTBN.Y.n13 6.57323
R17060 XThR.XTBN.Y.n29 XThR.XTBN.Y.n25 6.57323
R17061 XThR.XTBN.Y.n41 XThR.XTBN.Y.n37 6.57323
R17062 XThR.XTBN.Y.n53 XThR.XTBN.Y.n49 6.57323
R17063 XThR.XTBN.Y.n65 XThR.XTBN.Y.n61 6.57323
R17064 XThR.XTBN.Y.n77 XThR.XTBN.Y.n73 6.57323
R17065 XThR.XTBN.Y.n172 XThR.XTBN.Y 6.4005
R17066 XThR.XTBN.Y.n171 XThR.XTBN.Y 6.4005
R17067 XThR.XTBN.Y.n179 XThR.XTBN.Y.n178 5.74665
R17068 XThR.XTBN.Y.n178 XThR.XTBN.Y.n166 5.74569
R17069 XThR.XTBN.Y.n161 XThR.XTBN.Y 5.1205
R17070 XThR.XTBN.Y.n149 XThR.XTBN.Y 5.1205
R17071 XThR.XTBN.Y.n137 XThR.XTBN.Y 5.1205
R17072 XThR.XTBN.Y.n125 XThR.XTBN.Y 5.1205
R17073 XThR.XTBN.Y.n113 XThR.XTBN.Y 5.1205
R17074 XThR.XTBN.Y.n101 XThR.XTBN.Y 5.1205
R17075 XThR.XTBN.Y.n90 XThR.XTBN.Y 5.1205
R17076 XThR.XTBN.Y.n8 XThR.XTBN.Y.n7 5.11262
R17077 XThR.XTBN.Y.n19 XThR.XTBN.Y.n18 5.11262
R17078 XThR.XTBN.Y.n31 XThR.XTBN.Y.n30 5.11262
R17079 XThR.XTBN.Y.n43 XThR.XTBN.Y.n42 5.11262
R17080 XThR.XTBN.Y.n55 XThR.XTBN.Y.n54 5.11262
R17081 XThR.XTBN.Y.n67 XThR.XTBN.Y.n66 5.11262
R17082 XThR.XTBN.Y.n79 XThR.XTBN.Y.n78 5.11262
R17083 XThR.XTBN.Y.n182 XThR.XTBN.Y.n179 5.06717
R17084 XThR.XTBN.Y.n181 XThR.XTBN.Y 5.04292
R17085 XThR.XTBN.Y.n178 XThR.XTBN.Y.n177 4.6505
R17086 XThR.XTBN.Y.n176 XThR.XTBN.Y 4.3525
R17087 XThR.XTBN.Y XThR.XTBN.Y.n0 4.1605
R17088 XThR.XTBN.Y XThR.XTBN.Y.n11 4.1605
R17089 XThR.XTBN.Y XThR.XTBN.Y.n23 4.1605
R17090 XThR.XTBN.Y XThR.XTBN.Y.n35 4.1605
R17091 XThR.XTBN.Y XThR.XTBN.Y.n47 4.1605
R17092 XThR.XTBN.Y XThR.XTBN.Y.n59 4.1605
R17093 XThR.XTBN.Y XThR.XTBN.Y.n71 4.1605
R17094 XThR.XTBN.Y.n182 XThR.XTBN.Y 3.8405
R17095 XThR.XTBN.Y.n184 XThR.XTBN.Y 2.5605
R17096 XThR.XTBN.Y.n164 XThR.XTBN.Y 2.3045
R17097 XThR.XTBN.Y.n152 XThR.XTBN.Y 2.3045
R17098 XThR.XTBN.Y.n140 XThR.XTBN.Y 2.3045
R17099 XThR.XTBN.Y.n128 XThR.XTBN.Y 2.3045
R17100 XThR.XTBN.Y.n116 XThR.XTBN.Y 2.3045
R17101 XThR.XTBN.Y.n104 XThR.XTBN.Y 2.3045
R17102 XThR.XTBN.Y.n93 XThR.XTBN.Y 2.3045
R17103 XThR.XTBN.Y XThR.XTBN.Y.n184 1.93989
R17104 XThR.XTBN.Y.n166 XThR.XTBN.Y.n82 1.53415
R17105 XThR.XTBN.Y.n34 XThR.XTBN.Y.n22 1.49088
R17106 XThR.XTBN.Y.n58 XThR.XTBN.Y.n46 1.49088
R17107 XThR.XTBN.Y.n82 XThR.XTBN.Y.n70 1.48608
R17108 XThR.XTBN.Y.n153 XThR.XTBN.Y.n141 1.46204
R17109 XThR.XTBN.Y.n129 XThR.XTBN.Y.n117 1.46204
R17110 XThR.XTBN.Y.n166 XThR.XTBN.Y.n165 1.20723
R17111 XThR.XTBN.Y.n165 XThR.XTBN.Y.n153 1.15435
R17112 XThR.XTBN.Y.n141 XThR.XTBN.Y.n129 1.15435
R17113 XThR.XTBN.Y.n117 XThR.XTBN.Y.n105 1.15435
R17114 XThR.XTBN.Y.n70 XThR.XTBN.Y.n58 1.13031
R17115 XThR.XTBN.Y.n46 XThR.XTBN.Y.n34 1.1255
R17116 XThR.Tn[6].n2 XThR.Tn[6].n0 332.332
R17117 XThR.Tn[6].n2 XThR.Tn[6].n1 296.493
R17118 XThR.Tn[6] XThR.Tn[6].n82 161.363
R17119 XThR.Tn[6] XThR.Tn[6].n77 161.363
R17120 XThR.Tn[6] XThR.Tn[6].n72 161.363
R17121 XThR.Tn[6] XThR.Tn[6].n67 161.363
R17122 XThR.Tn[6] XThR.Tn[6].n62 161.363
R17123 XThR.Tn[6] XThR.Tn[6].n57 161.363
R17124 XThR.Tn[6] XThR.Tn[6].n52 161.363
R17125 XThR.Tn[6] XThR.Tn[6].n47 161.363
R17126 XThR.Tn[6] XThR.Tn[6].n42 161.363
R17127 XThR.Tn[6] XThR.Tn[6].n37 161.363
R17128 XThR.Tn[6] XThR.Tn[6].n32 161.363
R17129 XThR.Tn[6] XThR.Tn[6].n27 161.363
R17130 XThR.Tn[6] XThR.Tn[6].n22 161.363
R17131 XThR.Tn[6] XThR.Tn[6].n17 161.363
R17132 XThR.Tn[6] XThR.Tn[6].n12 161.363
R17133 XThR.Tn[6] XThR.Tn[6].n10 161.363
R17134 XThR.Tn[6].n84 XThR.Tn[6].n83 161.3
R17135 XThR.Tn[6].n79 XThR.Tn[6].n78 161.3
R17136 XThR.Tn[6].n74 XThR.Tn[6].n73 161.3
R17137 XThR.Tn[6].n69 XThR.Tn[6].n68 161.3
R17138 XThR.Tn[6].n64 XThR.Tn[6].n63 161.3
R17139 XThR.Tn[6].n59 XThR.Tn[6].n58 161.3
R17140 XThR.Tn[6].n54 XThR.Tn[6].n53 161.3
R17141 XThR.Tn[6].n49 XThR.Tn[6].n48 161.3
R17142 XThR.Tn[6].n44 XThR.Tn[6].n43 161.3
R17143 XThR.Tn[6].n39 XThR.Tn[6].n38 161.3
R17144 XThR.Tn[6].n34 XThR.Tn[6].n33 161.3
R17145 XThR.Tn[6].n29 XThR.Tn[6].n28 161.3
R17146 XThR.Tn[6].n24 XThR.Tn[6].n23 161.3
R17147 XThR.Tn[6].n19 XThR.Tn[6].n18 161.3
R17148 XThR.Tn[6].n14 XThR.Tn[6].n13 161.3
R17149 XThR.Tn[6].n82 XThR.Tn[6].t46 161.106
R17150 XThR.Tn[6].n77 XThR.Tn[6].t52 161.106
R17151 XThR.Tn[6].n72 XThR.Tn[6].t32 161.106
R17152 XThR.Tn[6].n67 XThR.Tn[6].t18 161.106
R17153 XThR.Tn[6].n62 XThR.Tn[6].t44 161.106
R17154 XThR.Tn[6].n57 XThR.Tn[6].t69 161.106
R17155 XThR.Tn[6].n52 XThR.Tn[6].t50 161.106
R17156 XThR.Tn[6].n47 XThR.Tn[6].t30 161.106
R17157 XThR.Tn[6].n42 XThR.Tn[6].t17 161.106
R17158 XThR.Tn[6].n37 XThR.Tn[6].t22 161.106
R17159 XThR.Tn[6].n32 XThR.Tn[6].t67 161.106
R17160 XThR.Tn[6].n27 XThR.Tn[6].t31 161.106
R17161 XThR.Tn[6].n22 XThR.Tn[6].t66 161.106
R17162 XThR.Tn[6].n17 XThR.Tn[6].t49 161.106
R17163 XThR.Tn[6].n12 XThR.Tn[6].t72 161.106
R17164 XThR.Tn[6].n10 XThR.Tn[6].t56 161.106
R17165 XThR.Tn[6].n83 XThR.Tn[6].t42 159.978
R17166 XThR.Tn[6].n78 XThR.Tn[6].t48 159.978
R17167 XThR.Tn[6].n73 XThR.Tn[6].t28 159.978
R17168 XThR.Tn[6].n68 XThR.Tn[6].t15 159.978
R17169 XThR.Tn[6].n63 XThR.Tn[6].t39 159.978
R17170 XThR.Tn[6].n58 XThR.Tn[6].t65 159.978
R17171 XThR.Tn[6].n53 XThR.Tn[6].t47 159.978
R17172 XThR.Tn[6].n48 XThR.Tn[6].t25 159.978
R17173 XThR.Tn[6].n43 XThR.Tn[6].t12 159.978
R17174 XThR.Tn[6].n38 XThR.Tn[6].t19 159.978
R17175 XThR.Tn[6].n33 XThR.Tn[6].t64 159.978
R17176 XThR.Tn[6].n28 XThR.Tn[6].t27 159.978
R17177 XThR.Tn[6].n23 XThR.Tn[6].t63 159.978
R17178 XThR.Tn[6].n18 XThR.Tn[6].t45 159.978
R17179 XThR.Tn[6].n13 XThR.Tn[6].t68 159.978
R17180 XThR.Tn[6].n82 XThR.Tn[6].t34 145.038
R17181 XThR.Tn[6].n77 XThR.Tn[6].t58 145.038
R17182 XThR.Tn[6].n72 XThR.Tn[6].t38 145.038
R17183 XThR.Tn[6].n67 XThR.Tn[6].t23 145.038
R17184 XThR.Tn[6].n62 XThR.Tn[6].t53 145.038
R17185 XThR.Tn[6].n57 XThR.Tn[6].t33 145.038
R17186 XThR.Tn[6].n52 XThR.Tn[6].t40 145.038
R17187 XThR.Tn[6].n47 XThR.Tn[6].t24 145.038
R17188 XThR.Tn[6].n42 XThR.Tn[6].t21 145.038
R17189 XThR.Tn[6].n37 XThR.Tn[6].t51 145.038
R17190 XThR.Tn[6].n32 XThR.Tn[6].t13 145.038
R17191 XThR.Tn[6].n27 XThR.Tn[6].t35 145.038
R17192 XThR.Tn[6].n22 XThR.Tn[6].t73 145.038
R17193 XThR.Tn[6].n17 XThR.Tn[6].t57 145.038
R17194 XThR.Tn[6].n12 XThR.Tn[6].t20 145.038
R17195 XThR.Tn[6].n10 XThR.Tn[6].t62 145.038
R17196 XThR.Tn[6].n83 XThR.Tn[6].t55 143.911
R17197 XThR.Tn[6].n78 XThR.Tn[6].t16 143.911
R17198 XThR.Tn[6].n73 XThR.Tn[6].t60 143.911
R17199 XThR.Tn[6].n68 XThR.Tn[6].t41 143.911
R17200 XThR.Tn[6].n63 XThR.Tn[6].t71 143.911
R17201 XThR.Tn[6].n58 XThR.Tn[6].t54 143.911
R17202 XThR.Tn[6].n53 XThR.Tn[6].t61 143.911
R17203 XThR.Tn[6].n48 XThR.Tn[6].t43 143.911
R17204 XThR.Tn[6].n43 XThR.Tn[6].t37 143.911
R17205 XThR.Tn[6].n38 XThR.Tn[6].t70 143.911
R17206 XThR.Tn[6].n33 XThR.Tn[6].t29 143.911
R17207 XThR.Tn[6].n28 XThR.Tn[6].t59 143.911
R17208 XThR.Tn[6].n23 XThR.Tn[6].t26 143.911
R17209 XThR.Tn[6].n18 XThR.Tn[6].t14 143.911
R17210 XThR.Tn[6].n13 XThR.Tn[6].t36 143.911
R17211 XThR.Tn[6].n5 XThR.Tn[6].n3 135.249
R17212 XThR.Tn[6].n5 XThR.Tn[6].n4 98.982
R17213 XThR.Tn[6].n7 XThR.Tn[6].n6 98.982
R17214 XThR.Tn[6].n9 XThR.Tn[6].n8 98.982
R17215 XThR.Tn[6].n7 XThR.Tn[6].n5 36.2672
R17216 XThR.Tn[6].n9 XThR.Tn[6].n7 36.2672
R17217 XThR.Tn[6].n88 XThR.Tn[6].n9 32.6405
R17218 XThR.Tn[6].n0 XThR.Tn[6].t2 26.5955
R17219 XThR.Tn[6].n0 XThR.Tn[6].t1 26.5955
R17220 XThR.Tn[6].n1 XThR.Tn[6].t3 26.5955
R17221 XThR.Tn[6].n1 XThR.Tn[6].t0 26.5955
R17222 XThR.Tn[6].n3 XThR.Tn[6].t8 24.9236
R17223 XThR.Tn[6].n3 XThR.Tn[6].t9 24.9236
R17224 XThR.Tn[6].n4 XThR.Tn[6].t11 24.9236
R17225 XThR.Tn[6].n4 XThR.Tn[6].t10 24.9236
R17226 XThR.Tn[6].n6 XThR.Tn[6].t7 24.9236
R17227 XThR.Tn[6].n6 XThR.Tn[6].t6 24.9236
R17228 XThR.Tn[6].n8 XThR.Tn[6].t4 24.9236
R17229 XThR.Tn[6].n8 XThR.Tn[6].t5 24.9236
R17230 XThR.Tn[6] XThR.Tn[6].n2 23.3605
R17231 XThR.Tn[6] XThR.Tn[6].n88 6.7205
R17232 XThR.Tn[6].n88 XThR.Tn[6] 5.37828
R17233 XThR.Tn[6] XThR.Tn[6].n11 5.34038
R17234 XThR.Tn[6].n16 XThR.Tn[6].n15 4.5005
R17235 XThR.Tn[6].n21 XThR.Tn[6].n20 4.5005
R17236 XThR.Tn[6].n26 XThR.Tn[6].n25 4.5005
R17237 XThR.Tn[6].n31 XThR.Tn[6].n30 4.5005
R17238 XThR.Tn[6].n36 XThR.Tn[6].n35 4.5005
R17239 XThR.Tn[6].n41 XThR.Tn[6].n40 4.5005
R17240 XThR.Tn[6].n46 XThR.Tn[6].n45 4.5005
R17241 XThR.Tn[6].n51 XThR.Tn[6].n50 4.5005
R17242 XThR.Tn[6].n56 XThR.Tn[6].n55 4.5005
R17243 XThR.Tn[6].n61 XThR.Tn[6].n60 4.5005
R17244 XThR.Tn[6].n66 XThR.Tn[6].n65 4.5005
R17245 XThR.Tn[6].n71 XThR.Tn[6].n70 4.5005
R17246 XThR.Tn[6].n76 XThR.Tn[6].n75 4.5005
R17247 XThR.Tn[6].n81 XThR.Tn[6].n80 4.5005
R17248 XThR.Tn[6].n86 XThR.Tn[6].n85 4.5005
R17249 XThR.Tn[6].n87 XThR.Tn[6] 3.70586
R17250 XThR.Tn[6].n16 XThR.Tn[6] 2.52282
R17251 XThR.Tn[6].n21 XThR.Tn[6] 2.52282
R17252 XThR.Tn[6].n26 XThR.Tn[6] 2.52282
R17253 XThR.Tn[6].n31 XThR.Tn[6] 2.52282
R17254 XThR.Tn[6].n36 XThR.Tn[6] 2.52282
R17255 XThR.Tn[6].n41 XThR.Tn[6] 2.52282
R17256 XThR.Tn[6].n46 XThR.Tn[6] 2.52282
R17257 XThR.Tn[6].n51 XThR.Tn[6] 2.52282
R17258 XThR.Tn[6].n56 XThR.Tn[6] 2.52282
R17259 XThR.Tn[6].n61 XThR.Tn[6] 2.52282
R17260 XThR.Tn[6].n66 XThR.Tn[6] 2.52282
R17261 XThR.Tn[6].n71 XThR.Tn[6] 2.52282
R17262 XThR.Tn[6].n76 XThR.Tn[6] 2.52282
R17263 XThR.Tn[6].n81 XThR.Tn[6] 2.52282
R17264 XThR.Tn[6].n86 XThR.Tn[6] 2.52282
R17265 XThR.Tn[6].n84 XThR.Tn[6] 1.08677
R17266 XThR.Tn[6].n79 XThR.Tn[6] 1.08677
R17267 XThR.Tn[6].n74 XThR.Tn[6] 1.08677
R17268 XThR.Tn[6].n69 XThR.Tn[6] 1.08677
R17269 XThR.Tn[6].n64 XThR.Tn[6] 1.08677
R17270 XThR.Tn[6].n59 XThR.Tn[6] 1.08677
R17271 XThR.Tn[6].n54 XThR.Tn[6] 1.08677
R17272 XThR.Tn[6].n49 XThR.Tn[6] 1.08677
R17273 XThR.Tn[6].n44 XThR.Tn[6] 1.08677
R17274 XThR.Tn[6].n39 XThR.Tn[6] 1.08677
R17275 XThR.Tn[6].n34 XThR.Tn[6] 1.08677
R17276 XThR.Tn[6].n29 XThR.Tn[6] 1.08677
R17277 XThR.Tn[6].n24 XThR.Tn[6] 1.08677
R17278 XThR.Tn[6].n19 XThR.Tn[6] 1.08677
R17279 XThR.Tn[6].n14 XThR.Tn[6] 1.08677
R17280 XThR.Tn[6] XThR.Tn[6].n16 0.839786
R17281 XThR.Tn[6] XThR.Tn[6].n21 0.839786
R17282 XThR.Tn[6] XThR.Tn[6].n26 0.839786
R17283 XThR.Tn[6] XThR.Tn[6].n31 0.839786
R17284 XThR.Tn[6] XThR.Tn[6].n36 0.839786
R17285 XThR.Tn[6] XThR.Tn[6].n41 0.839786
R17286 XThR.Tn[6] XThR.Tn[6].n46 0.839786
R17287 XThR.Tn[6] XThR.Tn[6].n51 0.839786
R17288 XThR.Tn[6] XThR.Tn[6].n56 0.839786
R17289 XThR.Tn[6] XThR.Tn[6].n61 0.839786
R17290 XThR.Tn[6] XThR.Tn[6].n66 0.839786
R17291 XThR.Tn[6] XThR.Tn[6].n71 0.839786
R17292 XThR.Tn[6] XThR.Tn[6].n76 0.839786
R17293 XThR.Tn[6] XThR.Tn[6].n81 0.839786
R17294 XThR.Tn[6] XThR.Tn[6].n86 0.839786
R17295 XThR.Tn[6].n11 XThR.Tn[6] 0.499542
R17296 XThR.Tn[6].n85 XThR.Tn[6] 0.063
R17297 XThR.Tn[6].n80 XThR.Tn[6] 0.063
R17298 XThR.Tn[6].n75 XThR.Tn[6] 0.063
R17299 XThR.Tn[6].n70 XThR.Tn[6] 0.063
R17300 XThR.Tn[6].n65 XThR.Tn[6] 0.063
R17301 XThR.Tn[6].n60 XThR.Tn[6] 0.063
R17302 XThR.Tn[6].n55 XThR.Tn[6] 0.063
R17303 XThR.Tn[6].n50 XThR.Tn[6] 0.063
R17304 XThR.Tn[6].n45 XThR.Tn[6] 0.063
R17305 XThR.Tn[6].n40 XThR.Tn[6] 0.063
R17306 XThR.Tn[6].n35 XThR.Tn[6] 0.063
R17307 XThR.Tn[6].n30 XThR.Tn[6] 0.063
R17308 XThR.Tn[6].n25 XThR.Tn[6] 0.063
R17309 XThR.Tn[6].n20 XThR.Tn[6] 0.063
R17310 XThR.Tn[6].n15 XThR.Tn[6] 0.063
R17311 XThR.Tn[6].n87 XThR.Tn[6] 0.0540714
R17312 XThR.Tn[6] XThR.Tn[6].n87 0.038
R17313 XThR.Tn[6].n11 XThR.Tn[6] 0.0143889
R17314 XThR.Tn[6].n85 XThR.Tn[6].n84 0.00771154
R17315 XThR.Tn[6].n80 XThR.Tn[6].n79 0.00771154
R17316 XThR.Tn[6].n75 XThR.Tn[6].n74 0.00771154
R17317 XThR.Tn[6].n70 XThR.Tn[6].n69 0.00771154
R17318 XThR.Tn[6].n65 XThR.Tn[6].n64 0.00771154
R17319 XThR.Tn[6].n60 XThR.Tn[6].n59 0.00771154
R17320 XThR.Tn[6].n55 XThR.Tn[6].n54 0.00771154
R17321 XThR.Tn[6].n50 XThR.Tn[6].n49 0.00771154
R17322 XThR.Tn[6].n45 XThR.Tn[6].n44 0.00771154
R17323 XThR.Tn[6].n40 XThR.Tn[6].n39 0.00771154
R17324 XThR.Tn[6].n35 XThR.Tn[6].n34 0.00771154
R17325 XThR.Tn[6].n30 XThR.Tn[6].n29 0.00771154
R17326 XThR.Tn[6].n25 XThR.Tn[6].n24 0.00771154
R17327 XThR.Tn[6].n20 XThR.Tn[6].n19 0.00771154
R17328 XThR.Tn[6].n15 XThR.Tn[6].n14 0.00771154
R17329 XThR.Tn[14].n87 XThR.Tn[14].n86 256.103
R17330 XThR.Tn[14].n2 XThR.Tn[14].n0 243.68
R17331 XThR.Tn[14].n5 XThR.Tn[14].n3 241.847
R17332 XThR.Tn[14].n2 XThR.Tn[14].n1 205.28
R17333 XThR.Tn[14].n87 XThR.Tn[14].n85 202.095
R17334 XThR.Tn[14].n5 XThR.Tn[14].n4 185
R17335 XThR.Tn[14] XThR.Tn[14].n78 161.363
R17336 XThR.Tn[14] XThR.Tn[14].n73 161.363
R17337 XThR.Tn[14] XThR.Tn[14].n68 161.363
R17338 XThR.Tn[14] XThR.Tn[14].n63 161.363
R17339 XThR.Tn[14] XThR.Tn[14].n58 161.363
R17340 XThR.Tn[14] XThR.Tn[14].n53 161.363
R17341 XThR.Tn[14] XThR.Tn[14].n48 161.363
R17342 XThR.Tn[14] XThR.Tn[14].n43 161.363
R17343 XThR.Tn[14] XThR.Tn[14].n38 161.363
R17344 XThR.Tn[14] XThR.Tn[14].n33 161.363
R17345 XThR.Tn[14] XThR.Tn[14].n28 161.363
R17346 XThR.Tn[14] XThR.Tn[14].n23 161.363
R17347 XThR.Tn[14] XThR.Tn[14].n18 161.363
R17348 XThR.Tn[14] XThR.Tn[14].n13 161.363
R17349 XThR.Tn[14] XThR.Tn[14].n8 161.363
R17350 XThR.Tn[14] XThR.Tn[14].n6 161.363
R17351 XThR.Tn[14].n80 XThR.Tn[14].n79 161.3
R17352 XThR.Tn[14].n75 XThR.Tn[14].n74 161.3
R17353 XThR.Tn[14].n70 XThR.Tn[14].n69 161.3
R17354 XThR.Tn[14].n65 XThR.Tn[14].n64 161.3
R17355 XThR.Tn[14].n60 XThR.Tn[14].n59 161.3
R17356 XThR.Tn[14].n55 XThR.Tn[14].n54 161.3
R17357 XThR.Tn[14].n50 XThR.Tn[14].n49 161.3
R17358 XThR.Tn[14].n45 XThR.Tn[14].n44 161.3
R17359 XThR.Tn[14].n40 XThR.Tn[14].n39 161.3
R17360 XThR.Tn[14].n35 XThR.Tn[14].n34 161.3
R17361 XThR.Tn[14].n30 XThR.Tn[14].n29 161.3
R17362 XThR.Tn[14].n25 XThR.Tn[14].n24 161.3
R17363 XThR.Tn[14].n20 XThR.Tn[14].n19 161.3
R17364 XThR.Tn[14].n15 XThR.Tn[14].n14 161.3
R17365 XThR.Tn[14].n10 XThR.Tn[14].n9 161.3
R17366 XThR.Tn[14].n78 XThR.Tn[14].t51 161.106
R17367 XThR.Tn[14].n73 XThR.Tn[14].t58 161.106
R17368 XThR.Tn[14].n68 XThR.Tn[14].t39 161.106
R17369 XThR.Tn[14].n63 XThR.Tn[14].t22 161.106
R17370 XThR.Tn[14].n58 XThR.Tn[14].t49 161.106
R17371 XThR.Tn[14].n53 XThR.Tn[14].t12 161.106
R17372 XThR.Tn[14].n48 XThR.Tn[14].t56 161.106
R17373 XThR.Tn[14].n43 XThR.Tn[14].t36 161.106
R17374 XThR.Tn[14].n38 XThR.Tn[14].t19 161.106
R17375 XThR.Tn[14].n33 XThR.Tn[14].t25 161.106
R17376 XThR.Tn[14].n28 XThR.Tn[14].t73 161.106
R17377 XThR.Tn[14].n23 XThR.Tn[14].t38 161.106
R17378 XThR.Tn[14].n18 XThR.Tn[14].t72 161.106
R17379 XThR.Tn[14].n13 XThR.Tn[14].t54 161.106
R17380 XThR.Tn[14].n8 XThR.Tn[14].t13 161.106
R17381 XThR.Tn[14].n6 XThR.Tn[14].t62 161.106
R17382 XThR.Tn[14].n79 XThR.Tn[14].t32 159.978
R17383 XThR.Tn[14].n74 XThR.Tn[14].t37 159.978
R17384 XThR.Tn[14].n69 XThR.Tn[14].t20 159.978
R17385 XThR.Tn[14].n64 XThR.Tn[14].t68 159.978
R17386 XThR.Tn[14].n59 XThR.Tn[14].t30 159.978
R17387 XThR.Tn[14].n54 XThR.Tn[14].t55 159.978
R17388 XThR.Tn[14].n49 XThR.Tn[14].t35 159.978
R17389 XThR.Tn[14].n44 XThR.Tn[14].t16 159.978
R17390 XThR.Tn[14].n39 XThR.Tn[14].t66 159.978
R17391 XThR.Tn[14].n34 XThR.Tn[14].t71 159.978
R17392 XThR.Tn[14].n29 XThR.Tn[14].t53 159.978
R17393 XThR.Tn[14].n24 XThR.Tn[14].t18 159.978
R17394 XThR.Tn[14].n19 XThR.Tn[14].t52 159.978
R17395 XThR.Tn[14].n14 XThR.Tn[14].t34 159.978
R17396 XThR.Tn[14].n9 XThR.Tn[14].t60 159.978
R17397 XThR.Tn[14].n78 XThR.Tn[14].t41 145.038
R17398 XThR.Tn[14].n73 XThR.Tn[14].t65 145.038
R17399 XThR.Tn[14].n68 XThR.Tn[14].t45 145.038
R17400 XThR.Tn[14].n63 XThR.Tn[14].t26 145.038
R17401 XThR.Tn[14].n58 XThR.Tn[14].t59 145.038
R17402 XThR.Tn[14].n53 XThR.Tn[14].t40 145.038
R17403 XThR.Tn[14].n48 XThR.Tn[14].t46 145.038
R17404 XThR.Tn[14].n43 XThR.Tn[14].t27 145.038
R17405 XThR.Tn[14].n38 XThR.Tn[14].t23 145.038
R17406 XThR.Tn[14].n33 XThR.Tn[14].t57 145.038
R17407 XThR.Tn[14].n28 XThR.Tn[14].t15 145.038
R17408 XThR.Tn[14].n23 XThR.Tn[14].t44 145.038
R17409 XThR.Tn[14].n18 XThR.Tn[14].t14 145.038
R17410 XThR.Tn[14].n13 XThR.Tn[14].t64 145.038
R17411 XThR.Tn[14].n8 XThR.Tn[14].t24 145.038
R17412 XThR.Tn[14].n6 XThR.Tn[14].t69 145.038
R17413 XThR.Tn[14].n79 XThR.Tn[14].t43 143.911
R17414 XThR.Tn[14].n74 XThR.Tn[14].t70 143.911
R17415 XThR.Tn[14].n69 XThR.Tn[14].t48 143.911
R17416 XThR.Tn[14].n64 XThR.Tn[14].t31 143.911
R17417 XThR.Tn[14].n59 XThR.Tn[14].t63 143.911
R17418 XThR.Tn[14].n54 XThR.Tn[14].t42 143.911
R17419 XThR.Tn[14].n49 XThR.Tn[14].t50 143.911
R17420 XThR.Tn[14].n44 XThR.Tn[14].t33 143.911
R17421 XThR.Tn[14].n39 XThR.Tn[14].t29 143.911
R17422 XThR.Tn[14].n34 XThR.Tn[14].t61 143.911
R17423 XThR.Tn[14].n29 XThR.Tn[14].t21 143.911
R17424 XThR.Tn[14].n24 XThR.Tn[14].t47 143.911
R17425 XThR.Tn[14].n19 XThR.Tn[14].t17 143.911
R17426 XThR.Tn[14].n14 XThR.Tn[14].t67 143.911
R17427 XThR.Tn[14].n9 XThR.Tn[14].t28 143.911
R17428 XThR.Tn[14] XThR.Tn[14].n2 35.7652
R17429 XThR.Tn[14].n0 XThR.Tn[14].t0 26.5955
R17430 XThR.Tn[14].n0 XThR.Tn[14].t1 26.5955
R17431 XThR.Tn[14].n85 XThR.Tn[14].t10 26.5955
R17432 XThR.Tn[14].n85 XThR.Tn[14].t11 26.5955
R17433 XThR.Tn[14].n86 XThR.Tn[14].t8 26.5955
R17434 XThR.Tn[14].n86 XThR.Tn[14].t9 26.5955
R17435 XThR.Tn[14].n1 XThR.Tn[14].t2 26.5955
R17436 XThR.Tn[14].n1 XThR.Tn[14].t3 26.5955
R17437 XThR.Tn[14].n4 XThR.Tn[14].t4 24.9236
R17438 XThR.Tn[14].n4 XThR.Tn[14].t5 24.9236
R17439 XThR.Tn[14].n3 XThR.Tn[14].t6 24.9236
R17440 XThR.Tn[14].n3 XThR.Tn[14].t7 24.9236
R17441 XThR.Tn[14] XThR.Tn[14].n5 18.8943
R17442 XThR.Tn[14].n88 XThR.Tn[14].n87 13.5534
R17443 XThR.Tn[14].n84 XThR.Tn[14] 8.47191
R17444 XThR.Tn[14].n84 XThR.Tn[14] 6.34069
R17445 XThR.Tn[14] XThR.Tn[14].n7 5.34038
R17446 XThR.Tn[14].n12 XThR.Tn[14].n11 4.5005
R17447 XThR.Tn[14].n17 XThR.Tn[14].n16 4.5005
R17448 XThR.Tn[14].n22 XThR.Tn[14].n21 4.5005
R17449 XThR.Tn[14].n27 XThR.Tn[14].n26 4.5005
R17450 XThR.Tn[14].n32 XThR.Tn[14].n31 4.5005
R17451 XThR.Tn[14].n37 XThR.Tn[14].n36 4.5005
R17452 XThR.Tn[14].n42 XThR.Tn[14].n41 4.5005
R17453 XThR.Tn[14].n47 XThR.Tn[14].n46 4.5005
R17454 XThR.Tn[14].n52 XThR.Tn[14].n51 4.5005
R17455 XThR.Tn[14].n57 XThR.Tn[14].n56 4.5005
R17456 XThR.Tn[14].n62 XThR.Tn[14].n61 4.5005
R17457 XThR.Tn[14].n67 XThR.Tn[14].n66 4.5005
R17458 XThR.Tn[14].n72 XThR.Tn[14].n71 4.5005
R17459 XThR.Tn[14].n77 XThR.Tn[14].n76 4.5005
R17460 XThR.Tn[14].n82 XThR.Tn[14].n81 4.5005
R17461 XThR.Tn[14].n83 XThR.Tn[14] 3.70586
R17462 XThR.Tn[14].n12 XThR.Tn[14] 2.52282
R17463 XThR.Tn[14].n17 XThR.Tn[14] 2.52282
R17464 XThR.Tn[14].n22 XThR.Tn[14] 2.52282
R17465 XThR.Tn[14].n27 XThR.Tn[14] 2.52282
R17466 XThR.Tn[14].n32 XThR.Tn[14] 2.52282
R17467 XThR.Tn[14].n37 XThR.Tn[14] 2.52282
R17468 XThR.Tn[14].n42 XThR.Tn[14] 2.52282
R17469 XThR.Tn[14].n47 XThR.Tn[14] 2.52282
R17470 XThR.Tn[14].n52 XThR.Tn[14] 2.52282
R17471 XThR.Tn[14].n57 XThR.Tn[14] 2.52282
R17472 XThR.Tn[14].n62 XThR.Tn[14] 2.52282
R17473 XThR.Tn[14].n67 XThR.Tn[14] 2.52282
R17474 XThR.Tn[14].n72 XThR.Tn[14] 2.52282
R17475 XThR.Tn[14].n77 XThR.Tn[14] 2.52282
R17476 XThR.Tn[14].n82 XThR.Tn[14] 2.52282
R17477 XThR.Tn[14] XThR.Tn[14].n84 1.79489
R17478 XThR.Tn[14] XThR.Tn[14].n88 1.50638
R17479 XThR.Tn[14].n88 XThR.Tn[14] 1.19676
R17480 XThR.Tn[14].n80 XThR.Tn[14] 1.08677
R17481 XThR.Tn[14].n75 XThR.Tn[14] 1.08677
R17482 XThR.Tn[14].n70 XThR.Tn[14] 1.08677
R17483 XThR.Tn[14].n65 XThR.Tn[14] 1.08677
R17484 XThR.Tn[14].n60 XThR.Tn[14] 1.08677
R17485 XThR.Tn[14].n55 XThR.Tn[14] 1.08677
R17486 XThR.Tn[14].n50 XThR.Tn[14] 1.08677
R17487 XThR.Tn[14].n45 XThR.Tn[14] 1.08677
R17488 XThR.Tn[14].n40 XThR.Tn[14] 1.08677
R17489 XThR.Tn[14].n35 XThR.Tn[14] 1.08677
R17490 XThR.Tn[14].n30 XThR.Tn[14] 1.08677
R17491 XThR.Tn[14].n25 XThR.Tn[14] 1.08677
R17492 XThR.Tn[14].n20 XThR.Tn[14] 1.08677
R17493 XThR.Tn[14].n15 XThR.Tn[14] 1.08677
R17494 XThR.Tn[14].n10 XThR.Tn[14] 1.08677
R17495 XThR.Tn[14] XThR.Tn[14].n12 0.839786
R17496 XThR.Tn[14] XThR.Tn[14].n17 0.839786
R17497 XThR.Tn[14] XThR.Tn[14].n22 0.839786
R17498 XThR.Tn[14] XThR.Tn[14].n27 0.839786
R17499 XThR.Tn[14] XThR.Tn[14].n32 0.839786
R17500 XThR.Tn[14] XThR.Tn[14].n37 0.839786
R17501 XThR.Tn[14] XThR.Tn[14].n42 0.839786
R17502 XThR.Tn[14] XThR.Tn[14].n47 0.839786
R17503 XThR.Tn[14] XThR.Tn[14].n52 0.839786
R17504 XThR.Tn[14] XThR.Tn[14].n57 0.839786
R17505 XThR.Tn[14] XThR.Tn[14].n62 0.839786
R17506 XThR.Tn[14] XThR.Tn[14].n67 0.839786
R17507 XThR.Tn[14] XThR.Tn[14].n72 0.839786
R17508 XThR.Tn[14] XThR.Tn[14].n77 0.839786
R17509 XThR.Tn[14] XThR.Tn[14].n82 0.839786
R17510 XThR.Tn[14].n7 XThR.Tn[14] 0.499542
R17511 XThR.Tn[14].n81 XThR.Tn[14] 0.063
R17512 XThR.Tn[14].n76 XThR.Tn[14] 0.063
R17513 XThR.Tn[14].n71 XThR.Tn[14] 0.063
R17514 XThR.Tn[14].n66 XThR.Tn[14] 0.063
R17515 XThR.Tn[14].n61 XThR.Tn[14] 0.063
R17516 XThR.Tn[14].n56 XThR.Tn[14] 0.063
R17517 XThR.Tn[14].n51 XThR.Tn[14] 0.063
R17518 XThR.Tn[14].n46 XThR.Tn[14] 0.063
R17519 XThR.Tn[14].n41 XThR.Tn[14] 0.063
R17520 XThR.Tn[14].n36 XThR.Tn[14] 0.063
R17521 XThR.Tn[14].n31 XThR.Tn[14] 0.063
R17522 XThR.Tn[14].n26 XThR.Tn[14] 0.063
R17523 XThR.Tn[14].n21 XThR.Tn[14] 0.063
R17524 XThR.Tn[14].n16 XThR.Tn[14] 0.063
R17525 XThR.Tn[14].n11 XThR.Tn[14] 0.063
R17526 XThR.Tn[14].n83 XThR.Tn[14] 0.0540714
R17527 XThR.Tn[14] XThR.Tn[14].n83 0.038
R17528 XThR.Tn[14].n7 XThR.Tn[14] 0.0143889
R17529 XThR.Tn[14].n81 XThR.Tn[14].n80 0.00771154
R17530 XThR.Tn[14].n76 XThR.Tn[14].n75 0.00771154
R17531 XThR.Tn[14].n71 XThR.Tn[14].n70 0.00771154
R17532 XThR.Tn[14].n66 XThR.Tn[14].n65 0.00771154
R17533 XThR.Tn[14].n61 XThR.Tn[14].n60 0.00771154
R17534 XThR.Tn[14].n56 XThR.Tn[14].n55 0.00771154
R17535 XThR.Tn[14].n51 XThR.Tn[14].n50 0.00771154
R17536 XThR.Tn[14].n46 XThR.Tn[14].n45 0.00771154
R17537 XThR.Tn[14].n41 XThR.Tn[14].n40 0.00771154
R17538 XThR.Tn[14].n36 XThR.Tn[14].n35 0.00771154
R17539 XThR.Tn[14].n31 XThR.Tn[14].n30 0.00771154
R17540 XThR.Tn[14].n26 XThR.Tn[14].n25 0.00771154
R17541 XThR.Tn[14].n21 XThR.Tn[14].n20 0.00771154
R17542 XThR.Tn[14].n16 XThR.Tn[14].n15 0.00771154
R17543 XThR.Tn[14].n11 XThR.Tn[14].n10 0.00771154
R17544 XThR.Tn[12].n87 XThR.Tn[12].n86 256.103
R17545 XThR.Tn[12].n2 XThR.Tn[12].n1 243.679
R17546 XThR.Tn[12].n5 XThR.Tn[12].n3 241.847
R17547 XThR.Tn[12].n2 XThR.Tn[12].n0 205.28
R17548 XThR.Tn[12].n87 XThR.Tn[12].n85 202.095
R17549 XThR.Tn[12].n5 XThR.Tn[12].n4 185
R17550 XThR.Tn[12] XThR.Tn[12].n78 161.363
R17551 XThR.Tn[12] XThR.Tn[12].n73 161.363
R17552 XThR.Tn[12] XThR.Tn[12].n68 161.363
R17553 XThR.Tn[12] XThR.Tn[12].n63 161.363
R17554 XThR.Tn[12] XThR.Tn[12].n58 161.363
R17555 XThR.Tn[12] XThR.Tn[12].n53 161.363
R17556 XThR.Tn[12] XThR.Tn[12].n48 161.363
R17557 XThR.Tn[12] XThR.Tn[12].n43 161.363
R17558 XThR.Tn[12] XThR.Tn[12].n38 161.363
R17559 XThR.Tn[12] XThR.Tn[12].n33 161.363
R17560 XThR.Tn[12] XThR.Tn[12].n28 161.363
R17561 XThR.Tn[12] XThR.Tn[12].n23 161.363
R17562 XThR.Tn[12] XThR.Tn[12].n18 161.363
R17563 XThR.Tn[12] XThR.Tn[12].n13 161.363
R17564 XThR.Tn[12] XThR.Tn[12].n8 161.363
R17565 XThR.Tn[12] XThR.Tn[12].n6 161.363
R17566 XThR.Tn[12].n80 XThR.Tn[12].n79 161.3
R17567 XThR.Tn[12].n75 XThR.Tn[12].n74 161.3
R17568 XThR.Tn[12].n70 XThR.Tn[12].n69 161.3
R17569 XThR.Tn[12].n65 XThR.Tn[12].n64 161.3
R17570 XThR.Tn[12].n60 XThR.Tn[12].n59 161.3
R17571 XThR.Tn[12].n55 XThR.Tn[12].n54 161.3
R17572 XThR.Tn[12].n50 XThR.Tn[12].n49 161.3
R17573 XThR.Tn[12].n45 XThR.Tn[12].n44 161.3
R17574 XThR.Tn[12].n40 XThR.Tn[12].n39 161.3
R17575 XThR.Tn[12].n35 XThR.Tn[12].n34 161.3
R17576 XThR.Tn[12].n30 XThR.Tn[12].n29 161.3
R17577 XThR.Tn[12].n25 XThR.Tn[12].n24 161.3
R17578 XThR.Tn[12].n20 XThR.Tn[12].n19 161.3
R17579 XThR.Tn[12].n15 XThR.Tn[12].n14 161.3
R17580 XThR.Tn[12].n10 XThR.Tn[12].n9 161.3
R17581 XThR.Tn[12].n78 XThR.Tn[12].t18 161.106
R17582 XThR.Tn[12].n73 XThR.Tn[12].t24 161.106
R17583 XThR.Tn[12].n68 XThR.Tn[12].t67 161.106
R17584 XThR.Tn[12].n63 XThR.Tn[12].t52 161.106
R17585 XThR.Tn[12].n58 XThR.Tn[12].t16 161.106
R17586 XThR.Tn[12].n53 XThR.Tn[12].t40 161.106
R17587 XThR.Tn[12].n48 XThR.Tn[12].t22 161.106
R17588 XThR.Tn[12].n43 XThR.Tn[12].t65 161.106
R17589 XThR.Tn[12].n38 XThR.Tn[12].t51 161.106
R17590 XThR.Tn[12].n33 XThR.Tn[12].t56 161.106
R17591 XThR.Tn[12].n28 XThR.Tn[12].t39 161.106
R17592 XThR.Tn[12].n23 XThR.Tn[12].t66 161.106
R17593 XThR.Tn[12].n18 XThR.Tn[12].t38 161.106
R17594 XThR.Tn[12].n13 XThR.Tn[12].t20 161.106
R17595 XThR.Tn[12].n8 XThR.Tn[12].t43 161.106
R17596 XThR.Tn[12].n6 XThR.Tn[12].t28 161.106
R17597 XThR.Tn[12].n79 XThR.Tn[12].t58 159.978
R17598 XThR.Tn[12].n74 XThR.Tn[12].t62 159.978
R17599 XThR.Tn[12].n69 XThR.Tn[12].t47 159.978
R17600 XThR.Tn[12].n64 XThR.Tn[12].t31 159.978
R17601 XThR.Tn[12].n59 XThR.Tn[12].t55 159.978
R17602 XThR.Tn[12].n54 XThR.Tn[12].t19 159.978
R17603 XThR.Tn[12].n49 XThR.Tn[12].t61 159.978
R17604 XThR.Tn[12].n44 XThR.Tn[12].t44 159.978
R17605 XThR.Tn[12].n39 XThR.Tn[12].t29 159.978
R17606 XThR.Tn[12].n34 XThR.Tn[12].t37 159.978
R17607 XThR.Tn[12].n29 XThR.Tn[12].t17 159.978
R17608 XThR.Tn[12].n24 XThR.Tn[12].t46 159.978
R17609 XThR.Tn[12].n19 XThR.Tn[12].t15 159.978
R17610 XThR.Tn[12].n14 XThR.Tn[12].t60 159.978
R17611 XThR.Tn[12].n9 XThR.Tn[12].t21 159.978
R17612 XThR.Tn[12].n78 XThR.Tn[12].t69 145.038
R17613 XThR.Tn[12].n73 XThR.Tn[12].t32 145.038
R17614 XThR.Tn[12].n68 XThR.Tn[12].t73 145.038
R17615 XThR.Tn[12].n63 XThR.Tn[12].t57 145.038
R17616 XThR.Tn[12].n58 XThR.Tn[12].t25 145.038
R17617 XThR.Tn[12].n53 XThR.Tn[12].t68 145.038
R17618 XThR.Tn[12].n48 XThR.Tn[12].t12 145.038
R17619 XThR.Tn[12].n43 XThR.Tn[12].t59 145.038
R17620 XThR.Tn[12].n38 XThR.Tn[12].t54 145.038
R17621 XThR.Tn[12].n33 XThR.Tn[12].t23 145.038
R17622 XThR.Tn[12].n28 XThR.Tn[12].t48 145.038
R17623 XThR.Tn[12].n23 XThR.Tn[12].t70 145.038
R17624 XThR.Tn[12].n18 XThR.Tn[12].t45 145.038
R17625 XThR.Tn[12].n13 XThR.Tn[12].t30 145.038
R17626 XThR.Tn[12].n8 XThR.Tn[12].t53 145.038
R17627 XThR.Tn[12].n6 XThR.Tn[12].t36 145.038
R17628 XThR.Tn[12].n79 XThR.Tn[12].t27 143.911
R17629 XThR.Tn[12].n74 XThR.Tn[12].t50 143.911
R17630 XThR.Tn[12].n69 XThR.Tn[12].t34 143.911
R17631 XThR.Tn[12].n64 XThR.Tn[12].t13 143.911
R17632 XThR.Tn[12].n59 XThR.Tn[12].t42 143.911
R17633 XThR.Tn[12].n54 XThR.Tn[12].t26 143.911
R17634 XThR.Tn[12].n49 XThR.Tn[12].t35 143.911
R17635 XThR.Tn[12].n44 XThR.Tn[12].t14 143.911
R17636 XThR.Tn[12].n39 XThR.Tn[12].t72 143.911
R17637 XThR.Tn[12].n34 XThR.Tn[12].t41 143.911
R17638 XThR.Tn[12].n29 XThR.Tn[12].t64 143.911
R17639 XThR.Tn[12].n24 XThR.Tn[12].t33 143.911
R17640 XThR.Tn[12].n19 XThR.Tn[12].t63 143.911
R17641 XThR.Tn[12].n14 XThR.Tn[12].t49 143.911
R17642 XThR.Tn[12].n9 XThR.Tn[12].t71 143.911
R17643 XThR.Tn[12] XThR.Tn[12].n2 35.7652
R17644 XThR.Tn[12].n85 XThR.Tn[12].t10 26.5955
R17645 XThR.Tn[12].n85 XThR.Tn[12].t8 26.5955
R17646 XThR.Tn[12].n86 XThR.Tn[12].t11 26.5955
R17647 XThR.Tn[12].n86 XThR.Tn[12].t9 26.5955
R17648 XThR.Tn[12].n0 XThR.Tn[12].t0 26.5955
R17649 XThR.Tn[12].n0 XThR.Tn[12].t2 26.5955
R17650 XThR.Tn[12].n1 XThR.Tn[12].t3 26.5955
R17651 XThR.Tn[12].n1 XThR.Tn[12].t1 26.5955
R17652 XThR.Tn[12].n4 XThR.Tn[12].t6 24.9236
R17653 XThR.Tn[12].n4 XThR.Tn[12].t4 24.9236
R17654 XThR.Tn[12].n3 XThR.Tn[12].t7 24.9236
R17655 XThR.Tn[12].n3 XThR.Tn[12].t5 24.9236
R17656 XThR.Tn[12] XThR.Tn[12].n5 18.8943
R17657 XThR.Tn[12].n88 XThR.Tn[12].n87 13.5534
R17658 XThR.Tn[12].n84 XThR.Tn[12] 8.18715
R17659 XThR.Tn[12].n84 XThR.Tn[12] 6.34069
R17660 XThR.Tn[12] XThR.Tn[12].n7 5.34038
R17661 XThR.Tn[12].n12 XThR.Tn[12].n11 4.5005
R17662 XThR.Tn[12].n17 XThR.Tn[12].n16 4.5005
R17663 XThR.Tn[12].n22 XThR.Tn[12].n21 4.5005
R17664 XThR.Tn[12].n27 XThR.Tn[12].n26 4.5005
R17665 XThR.Tn[12].n32 XThR.Tn[12].n31 4.5005
R17666 XThR.Tn[12].n37 XThR.Tn[12].n36 4.5005
R17667 XThR.Tn[12].n42 XThR.Tn[12].n41 4.5005
R17668 XThR.Tn[12].n47 XThR.Tn[12].n46 4.5005
R17669 XThR.Tn[12].n52 XThR.Tn[12].n51 4.5005
R17670 XThR.Tn[12].n57 XThR.Tn[12].n56 4.5005
R17671 XThR.Tn[12].n62 XThR.Tn[12].n61 4.5005
R17672 XThR.Tn[12].n67 XThR.Tn[12].n66 4.5005
R17673 XThR.Tn[12].n72 XThR.Tn[12].n71 4.5005
R17674 XThR.Tn[12].n77 XThR.Tn[12].n76 4.5005
R17675 XThR.Tn[12].n82 XThR.Tn[12].n81 4.5005
R17676 XThR.Tn[12].n83 XThR.Tn[12] 3.70586
R17677 XThR.Tn[12].n12 XThR.Tn[12] 2.52282
R17678 XThR.Tn[12].n17 XThR.Tn[12] 2.52282
R17679 XThR.Tn[12].n22 XThR.Tn[12] 2.52282
R17680 XThR.Tn[12].n27 XThR.Tn[12] 2.52282
R17681 XThR.Tn[12].n32 XThR.Tn[12] 2.52282
R17682 XThR.Tn[12].n37 XThR.Tn[12] 2.52282
R17683 XThR.Tn[12].n42 XThR.Tn[12] 2.52282
R17684 XThR.Tn[12].n47 XThR.Tn[12] 2.52282
R17685 XThR.Tn[12].n52 XThR.Tn[12] 2.52282
R17686 XThR.Tn[12].n57 XThR.Tn[12] 2.52282
R17687 XThR.Tn[12].n62 XThR.Tn[12] 2.52282
R17688 XThR.Tn[12].n67 XThR.Tn[12] 2.52282
R17689 XThR.Tn[12].n72 XThR.Tn[12] 2.52282
R17690 XThR.Tn[12].n77 XThR.Tn[12] 2.52282
R17691 XThR.Tn[12].n82 XThR.Tn[12] 2.52282
R17692 XThR.Tn[12] XThR.Tn[12].n84 1.79489
R17693 XThR.Tn[12] XThR.Tn[12].n88 1.50638
R17694 XThR.Tn[12].n88 XThR.Tn[12] 1.19676
R17695 XThR.Tn[12].n80 XThR.Tn[12] 1.08677
R17696 XThR.Tn[12].n75 XThR.Tn[12] 1.08677
R17697 XThR.Tn[12].n70 XThR.Tn[12] 1.08677
R17698 XThR.Tn[12].n65 XThR.Tn[12] 1.08677
R17699 XThR.Tn[12].n60 XThR.Tn[12] 1.08677
R17700 XThR.Tn[12].n55 XThR.Tn[12] 1.08677
R17701 XThR.Tn[12].n50 XThR.Tn[12] 1.08677
R17702 XThR.Tn[12].n45 XThR.Tn[12] 1.08677
R17703 XThR.Tn[12].n40 XThR.Tn[12] 1.08677
R17704 XThR.Tn[12].n35 XThR.Tn[12] 1.08677
R17705 XThR.Tn[12].n30 XThR.Tn[12] 1.08677
R17706 XThR.Tn[12].n25 XThR.Tn[12] 1.08677
R17707 XThR.Tn[12].n20 XThR.Tn[12] 1.08677
R17708 XThR.Tn[12].n15 XThR.Tn[12] 1.08677
R17709 XThR.Tn[12].n10 XThR.Tn[12] 1.08677
R17710 XThR.Tn[12] XThR.Tn[12].n12 0.839786
R17711 XThR.Tn[12] XThR.Tn[12].n17 0.839786
R17712 XThR.Tn[12] XThR.Tn[12].n22 0.839786
R17713 XThR.Tn[12] XThR.Tn[12].n27 0.839786
R17714 XThR.Tn[12] XThR.Tn[12].n32 0.839786
R17715 XThR.Tn[12] XThR.Tn[12].n37 0.839786
R17716 XThR.Tn[12] XThR.Tn[12].n42 0.839786
R17717 XThR.Tn[12] XThR.Tn[12].n47 0.839786
R17718 XThR.Tn[12] XThR.Tn[12].n52 0.839786
R17719 XThR.Tn[12] XThR.Tn[12].n57 0.839786
R17720 XThR.Tn[12] XThR.Tn[12].n62 0.839786
R17721 XThR.Tn[12] XThR.Tn[12].n67 0.839786
R17722 XThR.Tn[12] XThR.Tn[12].n72 0.839786
R17723 XThR.Tn[12] XThR.Tn[12].n77 0.839786
R17724 XThR.Tn[12] XThR.Tn[12].n82 0.839786
R17725 XThR.Tn[12].n7 XThR.Tn[12] 0.499542
R17726 XThR.Tn[12].n81 XThR.Tn[12] 0.063
R17727 XThR.Tn[12].n76 XThR.Tn[12] 0.063
R17728 XThR.Tn[12].n71 XThR.Tn[12] 0.063
R17729 XThR.Tn[12].n66 XThR.Tn[12] 0.063
R17730 XThR.Tn[12].n61 XThR.Tn[12] 0.063
R17731 XThR.Tn[12].n56 XThR.Tn[12] 0.063
R17732 XThR.Tn[12].n51 XThR.Tn[12] 0.063
R17733 XThR.Tn[12].n46 XThR.Tn[12] 0.063
R17734 XThR.Tn[12].n41 XThR.Tn[12] 0.063
R17735 XThR.Tn[12].n36 XThR.Tn[12] 0.063
R17736 XThR.Tn[12].n31 XThR.Tn[12] 0.063
R17737 XThR.Tn[12].n26 XThR.Tn[12] 0.063
R17738 XThR.Tn[12].n21 XThR.Tn[12] 0.063
R17739 XThR.Tn[12].n16 XThR.Tn[12] 0.063
R17740 XThR.Tn[12].n11 XThR.Tn[12] 0.063
R17741 XThR.Tn[12].n83 XThR.Tn[12] 0.0540714
R17742 XThR.Tn[12] XThR.Tn[12].n83 0.038
R17743 XThR.Tn[12].n7 XThR.Tn[12] 0.0143889
R17744 XThR.Tn[12].n81 XThR.Tn[12].n80 0.00771154
R17745 XThR.Tn[12].n76 XThR.Tn[12].n75 0.00771154
R17746 XThR.Tn[12].n71 XThR.Tn[12].n70 0.00771154
R17747 XThR.Tn[12].n66 XThR.Tn[12].n65 0.00771154
R17748 XThR.Tn[12].n61 XThR.Tn[12].n60 0.00771154
R17749 XThR.Tn[12].n56 XThR.Tn[12].n55 0.00771154
R17750 XThR.Tn[12].n51 XThR.Tn[12].n50 0.00771154
R17751 XThR.Tn[12].n46 XThR.Tn[12].n45 0.00771154
R17752 XThR.Tn[12].n41 XThR.Tn[12].n40 0.00771154
R17753 XThR.Tn[12].n36 XThR.Tn[12].n35 0.00771154
R17754 XThR.Tn[12].n31 XThR.Tn[12].n30 0.00771154
R17755 XThR.Tn[12].n26 XThR.Tn[12].n25 0.00771154
R17756 XThR.Tn[12].n21 XThR.Tn[12].n20 0.00771154
R17757 XThR.Tn[12].n16 XThR.Tn[12].n15 0.00771154
R17758 XThR.Tn[12].n11 XThR.Tn[12].n10 0.00771154
R17759 XThC.XTBN.Y.n182 XThC.XTBN.Y.t9 212.081
R17760 XThC.XTBN.Y.n181 XThC.XTBN.Y.t75 212.081
R17761 XThC.XTBN.Y.n175 XThC.XTBN.Y.t33 212.081
R17762 XThC.XTBN.Y.n176 XThC.XTBN.Y.t27 212.081
R17763 XThC.XTBN.Y.n87 XThC.XTBN.Y.t25 212.081
R17764 XThC.XTBN.Y.n78 XThC.XTBN.Y.t100 212.081
R17765 XThC.XTBN.Y.n82 XThC.XTBN.Y.t93 212.081
R17766 XThC.XTBN.Y.n80 XThC.XTBN.Y.t90 212.081
R17767 XThC.XTBN.Y.n61 XThC.XTBN.Y.t47 212.081
R17768 XThC.XTBN.Y.n52 XThC.XTBN.Y.t17 212.081
R17769 XThC.XTBN.Y.n56 XThC.XTBN.Y.t116 212.081
R17770 XThC.XTBN.Y.n54 XThC.XTBN.Y.t111 212.081
R17771 XThC.XTBN.Y.n35 XThC.XTBN.Y.t106 212.081
R17772 XThC.XTBN.Y.n26 XThC.XTBN.Y.t70 212.081
R17773 XThC.XTBN.Y.n30 XThC.XTBN.Y.t56 212.081
R17774 XThC.XTBN.Y.n28 XThC.XTBN.Y.t48 212.081
R17775 XThC.XTBN.Y.n10 XThC.XTBN.Y.t50 212.081
R17776 XThC.XTBN.Y.n1 XThC.XTBN.Y.t18 212.081
R17777 XThC.XTBN.Y.n5 XThC.XTBN.Y.t120 212.081
R17778 XThC.XTBN.Y.n3 XThC.XTBN.Y.t114 212.081
R17779 XThC.XTBN.Y.n74 XThC.XTBN.Y.t101 212.081
R17780 XThC.XTBN.Y.n65 XThC.XTBN.Y.t63 212.081
R17781 XThC.XTBN.Y.n69 XThC.XTBN.Y.t52 212.081
R17782 XThC.XTBN.Y.n67 XThC.XTBN.Y.t44 212.081
R17783 XThC.XTBN.Y.n48 XThC.XTBN.Y.t39 212.081
R17784 XThC.XTBN.Y.n39 XThC.XTBN.Y.t122 212.081
R17785 XThC.XTBN.Y.n43 XThC.XTBN.Y.t109 212.081
R17786 XThC.XTBN.Y.n41 XThC.XTBN.Y.t102 212.081
R17787 XThC.XTBN.Y.n22 XThC.XTBN.Y.t79 212.081
R17788 XThC.XTBN.Y.n13 XThC.XTBN.Y.t36 212.081
R17789 XThC.XTBN.Y.n17 XThC.XTBN.Y.t26 212.081
R17790 XThC.XTBN.Y.n15 XThC.XTBN.Y.t21 212.081
R17791 XThC.XTBN.Y.n99 XThC.XTBN.Y.t54 212.081
R17792 XThC.XTBN.Y.n98 XThC.XTBN.Y.t46 212.081
R17793 XThC.XTBN.Y.n93 XThC.XTBN.Y.t12 212.081
R17794 XThC.XTBN.Y.n92 XThC.XTBN.Y.t6 212.081
R17795 XThC.XTBN.Y.n122 XThC.XTBN.Y.t34 212.081
R17796 XThC.XTBN.Y.n121 XThC.XTBN.Y.t30 212.081
R17797 XThC.XTBN.Y.n116 XThC.XTBN.Y.t103 212.081
R17798 XThC.XTBN.Y.n115 XThC.XTBN.Y.t98 212.081
R17799 XThC.XTBN.Y.n146 XThC.XTBN.Y.t91 212.081
R17800 XThC.XTBN.Y.n145 XThC.XTBN.Y.t88 212.081
R17801 XThC.XTBN.Y.n140 XThC.XTBN.Y.t40 212.081
R17802 XThC.XTBN.Y.n139 XThC.XTBN.Y.t37 212.081
R17803 XThC.XTBN.Y.n170 XThC.XTBN.Y.t28 212.081
R17804 XThC.XTBN.Y.n169 XThC.XTBN.Y.t23 212.081
R17805 XThC.XTBN.Y.n164 XThC.XTBN.Y.t97 212.081
R17806 XThC.XTBN.Y.n163 XThC.XTBN.Y.t95 212.081
R17807 XThC.XTBN.Y.n110 XThC.XTBN.Y.t42 212.081
R17808 XThC.XTBN.Y.n109 XThC.XTBN.Y.t38 212.081
R17809 XThC.XTBN.Y.n104 XThC.XTBN.Y.t119 212.081
R17810 XThC.XTBN.Y.n103 XThC.XTBN.Y.t113 212.081
R17811 XThC.XTBN.Y.n134 XThC.XTBN.Y.t99 212.081
R17812 XThC.XTBN.Y.n133 XThC.XTBN.Y.t96 212.081
R17813 XThC.XTBN.Y.n128 XThC.XTBN.Y.t58 212.081
R17814 XThC.XTBN.Y.n127 XThC.XTBN.Y.t51 212.081
R17815 XThC.XTBN.Y.n158 XThC.XTBN.Y.t13 212.081
R17816 XThC.XTBN.Y.n157 XThC.XTBN.Y.t7 212.081
R17817 XThC.XTBN.Y.n152 XThC.XTBN.Y.t86 212.081
R17818 XThC.XTBN.Y.n151 XThC.XTBN.Y.t81 212.081
R17819 XThC.XTBN.Y.n189 XThC.XTBN.Y.n188 208.965
R17820 XThC.XTBN.Y.n176 XThC.XTBN.Y.n0 188.516
R17821 XThC.XTBN.Y.n88 XThC.XTBN.Y.n87 180.482
R17822 XThC.XTBN.Y.n62 XThC.XTBN.Y.n61 180.482
R17823 XThC.XTBN.Y.n36 XThC.XTBN.Y.n35 180.482
R17824 XThC.XTBN.Y.n11 XThC.XTBN.Y.n10 180.482
R17825 XThC.XTBN.Y.n75 XThC.XTBN.Y.n74 180.482
R17826 XThC.XTBN.Y.n49 XThC.XTBN.Y.n48 180.482
R17827 XThC.XTBN.Y.n23 XThC.XTBN.Y.n22 180.482
R17828 XThC.XTBN.Y.n95 XThC.XTBN.Y.n94 173.761
R17829 XThC.XTBN.Y.n118 XThC.XTBN.Y.n117 173.761
R17830 XThC.XTBN.Y.n142 XThC.XTBN.Y.n141 173.761
R17831 XThC.XTBN.Y.n166 XThC.XTBN.Y.n165 173.761
R17832 XThC.XTBN.Y.n106 XThC.XTBN.Y.n105 173.761
R17833 XThC.XTBN.Y.n130 XThC.XTBN.Y.n129 173.761
R17834 XThC.XTBN.Y.n154 XThC.XTBN.Y.n153 173.761
R17835 XThC.XTBN.Y.n81 XThC.XTBN.Y.n79 152
R17836 XThC.XTBN.Y.n84 XThC.XTBN.Y.n83 152
R17837 XThC.XTBN.Y.n86 XThC.XTBN.Y.n85 152
R17838 XThC.XTBN.Y.n55 XThC.XTBN.Y.n53 152
R17839 XThC.XTBN.Y.n58 XThC.XTBN.Y.n57 152
R17840 XThC.XTBN.Y.n60 XThC.XTBN.Y.n59 152
R17841 XThC.XTBN.Y.n29 XThC.XTBN.Y.n27 152
R17842 XThC.XTBN.Y.n32 XThC.XTBN.Y.n31 152
R17843 XThC.XTBN.Y.n34 XThC.XTBN.Y.n33 152
R17844 XThC.XTBN.Y.n4 XThC.XTBN.Y.n2 152
R17845 XThC.XTBN.Y.n7 XThC.XTBN.Y.n6 152
R17846 XThC.XTBN.Y.n9 XThC.XTBN.Y.n8 152
R17847 XThC.XTBN.Y.n68 XThC.XTBN.Y.n66 152
R17848 XThC.XTBN.Y.n71 XThC.XTBN.Y.n70 152
R17849 XThC.XTBN.Y.n73 XThC.XTBN.Y.n72 152
R17850 XThC.XTBN.Y.n42 XThC.XTBN.Y.n40 152
R17851 XThC.XTBN.Y.n45 XThC.XTBN.Y.n44 152
R17852 XThC.XTBN.Y.n47 XThC.XTBN.Y.n46 152
R17853 XThC.XTBN.Y.n16 XThC.XTBN.Y.n14 152
R17854 XThC.XTBN.Y.n19 XThC.XTBN.Y.n18 152
R17855 XThC.XTBN.Y.n21 XThC.XTBN.Y.n20 152
R17856 XThC.XTBN.Y.n95 XThC.XTBN.Y.n91 152
R17857 XThC.XTBN.Y.n97 XThC.XTBN.Y.n96 152
R17858 XThC.XTBN.Y.n101 XThC.XTBN.Y.n100 152
R17859 XThC.XTBN.Y.n118 XThC.XTBN.Y.n114 152
R17860 XThC.XTBN.Y.n120 XThC.XTBN.Y.n119 152
R17861 XThC.XTBN.Y.n124 XThC.XTBN.Y.n123 152
R17862 XThC.XTBN.Y.n142 XThC.XTBN.Y.n138 152
R17863 XThC.XTBN.Y.n144 XThC.XTBN.Y.n143 152
R17864 XThC.XTBN.Y.n148 XThC.XTBN.Y.n147 152
R17865 XThC.XTBN.Y.n166 XThC.XTBN.Y.n162 152
R17866 XThC.XTBN.Y.n168 XThC.XTBN.Y.n167 152
R17867 XThC.XTBN.Y.n172 XThC.XTBN.Y.n171 152
R17868 XThC.XTBN.Y.n106 XThC.XTBN.Y.n102 152
R17869 XThC.XTBN.Y.n108 XThC.XTBN.Y.n107 152
R17870 XThC.XTBN.Y.n112 XThC.XTBN.Y.n111 152
R17871 XThC.XTBN.Y.n130 XThC.XTBN.Y.n126 152
R17872 XThC.XTBN.Y.n132 XThC.XTBN.Y.n131 152
R17873 XThC.XTBN.Y.n136 XThC.XTBN.Y.n135 152
R17874 XThC.XTBN.Y.n154 XThC.XTBN.Y.n150 152
R17875 XThC.XTBN.Y.n156 XThC.XTBN.Y.n155 152
R17876 XThC.XTBN.Y.n160 XThC.XTBN.Y.n159 152
R17877 XThC.XTBN.Y.n178 XThC.XTBN.Y.n177 152
R17878 XThC.XTBN.Y.n180 XThC.XTBN.Y.n179 152
R17879 XThC.XTBN.Y.n184 XThC.XTBN.Y.n183 152
R17880 XThC.XTBN.Y.n182 XThC.XTBN.Y.t14 139.78
R17881 XThC.XTBN.Y.n181 XThC.XTBN.Y.t105 139.78
R17882 XThC.XTBN.Y.n175 XThC.XTBN.Y.t69 139.78
R17883 XThC.XTBN.Y.n176 XThC.XTBN.Y.t61 139.78
R17884 XThC.XTBN.Y.n87 XThC.XTBN.Y.t123 139.78
R17885 XThC.XTBN.Y.n78 XThC.XTBN.Y.t85 139.78
R17886 XThC.XTBN.Y.n82 XThC.XTBN.Y.t74 139.78
R17887 XThC.XTBN.Y.n80 XThC.XTBN.Y.t65 139.78
R17888 XThC.XTBN.Y.n61 XThC.XTBN.Y.t31 139.78
R17889 XThC.XTBN.Y.n52 XThC.XTBN.Y.t104 139.78
R17890 XThC.XTBN.Y.n56 XThC.XTBN.Y.t94 139.78
R17891 XThC.XTBN.Y.n54 XThC.XTBN.Y.t92 139.78
R17892 XThC.XTBN.Y.n35 XThC.XTBN.Y.t89 139.78
R17893 XThC.XTBN.Y.n26 XThC.XTBN.Y.t41 139.78
R17894 XThC.XTBN.Y.n30 XThC.XTBN.Y.t35 139.78
R17895 XThC.XTBN.Y.n28 XThC.XTBN.Y.t32 139.78
R17896 XThC.XTBN.Y.n10 XThC.XTBN.Y.t118 139.78
R17897 XThC.XTBN.Y.n1 XThC.XTBN.Y.t83 139.78
R17898 XThC.XTBN.Y.n5 XThC.XTBN.Y.t71 139.78
R17899 XThC.XTBN.Y.n3 XThC.XTBN.Y.t62 139.78
R17900 XThC.XTBN.Y.n74 XThC.XTBN.Y.t107 139.78
R17901 XThC.XTBN.Y.n65 XThC.XTBN.Y.t72 139.78
R17902 XThC.XTBN.Y.n69 XThC.XTBN.Y.t57 139.78
R17903 XThC.XTBN.Y.n67 XThC.XTBN.Y.t49 139.78
R17904 XThC.XTBN.Y.n48 XThC.XTBN.Y.t43 139.78
R17905 XThC.XTBN.Y.n39 XThC.XTBN.Y.t10 139.78
R17906 XThC.XTBN.Y.n43 XThC.XTBN.Y.t112 139.78
R17907 XThC.XTBN.Y.n41 XThC.XTBN.Y.t108 139.78
R17908 XThC.XTBN.Y.n22 XThC.XTBN.Y.t121 139.78
R17909 XThC.XTBN.Y.n13 XThC.XTBN.Y.t84 139.78
R17910 XThC.XTBN.Y.n17 XThC.XTBN.Y.t73 139.78
R17911 XThC.XTBN.Y.n15 XThC.XTBN.Y.t64 139.78
R17912 XThC.XTBN.Y.n99 XThC.XTBN.Y.t76 139.78
R17913 XThC.XTBN.Y.n98 XThC.XTBN.Y.t67 139.78
R17914 XThC.XTBN.Y.n93 XThC.XTBN.Y.t29 139.78
R17915 XThC.XTBN.Y.n92 XThC.XTBN.Y.t24 139.78
R17916 XThC.XTBN.Y.n122 XThC.XTBN.Y.t15 139.78
R17917 XThC.XTBN.Y.n121 XThC.XTBN.Y.t8 139.78
R17918 XThC.XTBN.Y.n116 XThC.XTBN.Y.t87 139.78
R17919 XThC.XTBN.Y.n115 XThC.XTBN.Y.t82 139.78
R17920 XThC.XTBN.Y.n146 XThC.XTBN.Y.t66 139.78
R17921 XThC.XTBN.Y.n145 XThC.XTBN.Y.t60 139.78
R17922 XThC.XTBN.Y.n140 XThC.XTBN.Y.t22 139.78
R17923 XThC.XTBN.Y.n139 XThC.XTBN.Y.t20 139.78
R17924 XThC.XTBN.Y.n170 XThC.XTBN.Y.t4 139.78
R17925 XThC.XTBN.Y.n169 XThC.XTBN.Y.t117 139.78
R17926 XThC.XTBN.Y.n164 XThC.XTBN.Y.t80 139.78
R17927 XThC.XTBN.Y.n163 XThC.XTBN.Y.t78 139.78
R17928 XThC.XTBN.Y.n110 XThC.XTBN.Y.t59 139.78
R17929 XThC.XTBN.Y.n109 XThC.XTBN.Y.t55 139.78
R17930 XThC.XTBN.Y.n104 XThC.XTBN.Y.t19 139.78
R17931 XThC.XTBN.Y.n103 XThC.XTBN.Y.t16 139.78
R17932 XThC.XTBN.Y.n134 XThC.XTBN.Y.t115 139.78
R17933 XThC.XTBN.Y.n133 XThC.XTBN.Y.t110 139.78
R17934 XThC.XTBN.Y.n128 XThC.XTBN.Y.t77 139.78
R17935 XThC.XTBN.Y.n127 XThC.XTBN.Y.t68 139.78
R17936 XThC.XTBN.Y.n158 XThC.XTBN.Y.t53 139.78
R17937 XThC.XTBN.Y.n157 XThC.XTBN.Y.t45 139.78
R17938 XThC.XTBN.Y.n152 XThC.XTBN.Y.t11 139.78
R17939 XThC.XTBN.Y.n151 XThC.XTBN.Y.t5 139.78
R17940 XThC.XTBN.Y XThC.XTBN.Y.n192 96.8352
R17941 XThC.XTBN.Y.n187 XThC.XTBN.Y.n0 64.6909
R17942 XThC.XTBN.Y.n97 XThC.XTBN.Y.n91 49.6611
R17943 XThC.XTBN.Y.n120 XThC.XTBN.Y.n114 49.6611
R17944 XThC.XTBN.Y.n144 XThC.XTBN.Y.n138 49.6611
R17945 XThC.XTBN.Y.n168 XThC.XTBN.Y.n162 49.6611
R17946 XThC.XTBN.Y.n108 XThC.XTBN.Y.n102 49.6611
R17947 XThC.XTBN.Y.n132 XThC.XTBN.Y.n126 49.6611
R17948 XThC.XTBN.Y.n156 XThC.XTBN.Y.n150 49.6611
R17949 XThC.XTBN.Y.n100 XThC.XTBN.Y.n98 44.549
R17950 XThC.XTBN.Y.n123 XThC.XTBN.Y.n121 44.549
R17951 XThC.XTBN.Y.n147 XThC.XTBN.Y.n145 44.549
R17952 XThC.XTBN.Y.n171 XThC.XTBN.Y.n169 44.549
R17953 XThC.XTBN.Y.n111 XThC.XTBN.Y.n109 44.549
R17954 XThC.XTBN.Y.n135 XThC.XTBN.Y.n133 44.549
R17955 XThC.XTBN.Y.n159 XThC.XTBN.Y.n157 44.549
R17956 XThC.XTBN.Y.n94 XThC.XTBN.Y.n93 43.0884
R17957 XThC.XTBN.Y.n117 XThC.XTBN.Y.n116 43.0884
R17958 XThC.XTBN.Y.n141 XThC.XTBN.Y.n140 43.0884
R17959 XThC.XTBN.Y.n165 XThC.XTBN.Y.n164 43.0884
R17960 XThC.XTBN.Y.n105 XThC.XTBN.Y.n104 43.0884
R17961 XThC.XTBN.Y.n129 XThC.XTBN.Y.n128 43.0884
R17962 XThC.XTBN.Y.n153 XThC.XTBN.Y.n152 43.0884
R17963 XThC.XTBN.Y.n177 XThC.XTBN.Y.n176 30.6732
R17964 XThC.XTBN.Y.n177 XThC.XTBN.Y.n175 30.6732
R17965 XThC.XTBN.Y.n180 XThC.XTBN.Y.n175 30.6732
R17966 XThC.XTBN.Y.n181 XThC.XTBN.Y.n180 30.6732
R17967 XThC.XTBN.Y.n183 XThC.XTBN.Y.n181 30.6732
R17968 XThC.XTBN.Y.n183 XThC.XTBN.Y.n182 30.6732
R17969 XThC.XTBN.Y.n81 XThC.XTBN.Y.n80 30.6732
R17970 XThC.XTBN.Y.n82 XThC.XTBN.Y.n81 30.6732
R17971 XThC.XTBN.Y.n83 XThC.XTBN.Y.n82 30.6732
R17972 XThC.XTBN.Y.n83 XThC.XTBN.Y.n78 30.6732
R17973 XThC.XTBN.Y.n86 XThC.XTBN.Y.n78 30.6732
R17974 XThC.XTBN.Y.n87 XThC.XTBN.Y.n86 30.6732
R17975 XThC.XTBN.Y.n55 XThC.XTBN.Y.n54 30.6732
R17976 XThC.XTBN.Y.n56 XThC.XTBN.Y.n55 30.6732
R17977 XThC.XTBN.Y.n57 XThC.XTBN.Y.n56 30.6732
R17978 XThC.XTBN.Y.n57 XThC.XTBN.Y.n52 30.6732
R17979 XThC.XTBN.Y.n60 XThC.XTBN.Y.n52 30.6732
R17980 XThC.XTBN.Y.n61 XThC.XTBN.Y.n60 30.6732
R17981 XThC.XTBN.Y.n29 XThC.XTBN.Y.n28 30.6732
R17982 XThC.XTBN.Y.n30 XThC.XTBN.Y.n29 30.6732
R17983 XThC.XTBN.Y.n31 XThC.XTBN.Y.n30 30.6732
R17984 XThC.XTBN.Y.n31 XThC.XTBN.Y.n26 30.6732
R17985 XThC.XTBN.Y.n34 XThC.XTBN.Y.n26 30.6732
R17986 XThC.XTBN.Y.n35 XThC.XTBN.Y.n34 30.6732
R17987 XThC.XTBN.Y.n4 XThC.XTBN.Y.n3 30.6732
R17988 XThC.XTBN.Y.n5 XThC.XTBN.Y.n4 30.6732
R17989 XThC.XTBN.Y.n6 XThC.XTBN.Y.n5 30.6732
R17990 XThC.XTBN.Y.n6 XThC.XTBN.Y.n1 30.6732
R17991 XThC.XTBN.Y.n9 XThC.XTBN.Y.n1 30.6732
R17992 XThC.XTBN.Y.n10 XThC.XTBN.Y.n9 30.6732
R17993 XThC.XTBN.Y.n68 XThC.XTBN.Y.n67 30.6732
R17994 XThC.XTBN.Y.n69 XThC.XTBN.Y.n68 30.6732
R17995 XThC.XTBN.Y.n70 XThC.XTBN.Y.n69 30.6732
R17996 XThC.XTBN.Y.n70 XThC.XTBN.Y.n65 30.6732
R17997 XThC.XTBN.Y.n73 XThC.XTBN.Y.n65 30.6732
R17998 XThC.XTBN.Y.n74 XThC.XTBN.Y.n73 30.6732
R17999 XThC.XTBN.Y.n42 XThC.XTBN.Y.n41 30.6732
R18000 XThC.XTBN.Y.n43 XThC.XTBN.Y.n42 30.6732
R18001 XThC.XTBN.Y.n44 XThC.XTBN.Y.n43 30.6732
R18002 XThC.XTBN.Y.n44 XThC.XTBN.Y.n39 30.6732
R18003 XThC.XTBN.Y.n47 XThC.XTBN.Y.n39 30.6732
R18004 XThC.XTBN.Y.n48 XThC.XTBN.Y.n47 30.6732
R18005 XThC.XTBN.Y.n16 XThC.XTBN.Y.n15 30.6732
R18006 XThC.XTBN.Y.n17 XThC.XTBN.Y.n16 30.6732
R18007 XThC.XTBN.Y.n18 XThC.XTBN.Y.n17 30.6732
R18008 XThC.XTBN.Y.n18 XThC.XTBN.Y.n13 30.6732
R18009 XThC.XTBN.Y.n21 XThC.XTBN.Y.n13 30.6732
R18010 XThC.XTBN.Y.n22 XThC.XTBN.Y.n21 30.6732
R18011 XThC.XTBN.Y.n188 XThC.XTBN.Y.t2 26.5955
R18012 XThC.XTBN.Y.n188 XThC.XTBN.Y.t3 26.5955
R18013 XThC.XTBN.Y.n192 XThC.XTBN.Y.t1 24.9236
R18014 XThC.XTBN.Y.n192 XThC.XTBN.Y.t0 24.9236
R18015 XThC.XTBN.Y.n96 XThC.XTBN.Y.n95 21.7605
R18016 XThC.XTBN.Y.n119 XThC.XTBN.Y.n118 21.7605
R18017 XThC.XTBN.Y.n143 XThC.XTBN.Y.n142 21.7605
R18018 XThC.XTBN.Y.n167 XThC.XTBN.Y.n166 21.7605
R18019 XThC.XTBN.Y.n107 XThC.XTBN.Y.n106 21.7605
R18020 XThC.XTBN.Y.n131 XThC.XTBN.Y.n130 21.7605
R18021 XThC.XTBN.Y.n155 XThC.XTBN.Y.n154 21.7605
R18022 XThC.XTBN.Y.n84 XThC.XTBN.Y.n79 21.5045
R18023 XThC.XTBN.Y.n58 XThC.XTBN.Y.n53 21.5045
R18024 XThC.XTBN.Y.n32 XThC.XTBN.Y.n27 21.5045
R18025 XThC.XTBN.Y.n7 XThC.XTBN.Y.n2 21.5045
R18026 XThC.XTBN.Y.n71 XThC.XTBN.Y.n66 21.5045
R18027 XThC.XTBN.Y.n45 XThC.XTBN.Y.n40 21.5045
R18028 XThC.XTBN.Y.n19 XThC.XTBN.Y.n14 21.5045
R18029 XThC.XTBN.Y.n178 XThC.XTBN.Y 21.2485
R18030 XThC.XTBN.Y.n85 XThC.XTBN.Y 19.9685
R18031 XThC.XTBN.Y.n59 XThC.XTBN.Y 19.9685
R18032 XThC.XTBN.Y.n33 XThC.XTBN.Y 19.9685
R18033 XThC.XTBN.Y.n8 XThC.XTBN.Y 19.9685
R18034 XThC.XTBN.Y.n72 XThC.XTBN.Y 19.9685
R18035 XThC.XTBN.Y.n46 XThC.XTBN.Y 19.9685
R18036 XThC.XTBN.Y.n20 XThC.XTBN.Y 19.9685
R18037 XThC.XTBN.Y.n179 XThC.XTBN.Y 19.2005
R18038 XThC.XTBN.Y.n94 XThC.XTBN.Y.n92 18.2581
R18039 XThC.XTBN.Y.n117 XThC.XTBN.Y.n115 18.2581
R18040 XThC.XTBN.Y.n141 XThC.XTBN.Y.n139 18.2581
R18041 XThC.XTBN.Y.n165 XThC.XTBN.Y.n163 18.2581
R18042 XThC.XTBN.Y.n105 XThC.XTBN.Y.n103 18.2581
R18043 XThC.XTBN.Y.n129 XThC.XTBN.Y.n127 18.2581
R18044 XThC.XTBN.Y.n153 XThC.XTBN.Y.n151 18.2581
R18045 XThC.XTBN.Y.n113 XThC.XTBN.Y.n101 17.1655
R18046 XThC.XTBN.Y.n88 XThC.XTBN.Y 17.1525
R18047 XThC.XTBN.Y.n62 XThC.XTBN.Y 17.1525
R18048 XThC.XTBN.Y.n36 XThC.XTBN.Y 17.1525
R18049 XThC.XTBN.Y.n11 XThC.XTBN.Y 17.1525
R18050 XThC.XTBN.Y.n75 XThC.XTBN.Y 17.1525
R18051 XThC.XTBN.Y.n49 XThC.XTBN.Y 17.1525
R18052 XThC.XTBN.Y.n23 XThC.XTBN.Y 17.1525
R18053 XThC.XTBN.Y.n100 XThC.XTBN.Y.n99 16.7975
R18054 XThC.XTBN.Y.n123 XThC.XTBN.Y.n122 16.7975
R18055 XThC.XTBN.Y.n147 XThC.XTBN.Y.n146 16.7975
R18056 XThC.XTBN.Y.n171 XThC.XTBN.Y.n170 16.7975
R18057 XThC.XTBN.Y.n111 XThC.XTBN.Y.n110 16.7975
R18058 XThC.XTBN.Y.n135 XThC.XTBN.Y.n134 16.7975
R18059 XThC.XTBN.Y.n159 XThC.XTBN.Y.n158 16.7975
R18060 XThC.XTBN.Y.n125 XThC.XTBN.Y.n124 16.0405
R18061 XThC.XTBN.Y.n149 XThC.XTBN.Y.n148 16.0405
R18062 XThC.XTBN.Y.n173 XThC.XTBN.Y.n172 16.0405
R18063 XThC.XTBN.Y.n113 XThC.XTBN.Y.n112 16.0405
R18064 XThC.XTBN.Y.n137 XThC.XTBN.Y.n136 16.0405
R18065 XThC.XTBN.Y.n161 XThC.XTBN.Y.n160 16.0405
R18066 XThC.XTBN.Y.n25 XThC.XTBN.Y.n12 15.262
R18067 XThC.XTBN.Y.n101 XThC.XTBN.Y 15.0405
R18068 XThC.XTBN.Y.n124 XThC.XTBN.Y 15.0405
R18069 XThC.XTBN.Y.n148 XThC.XTBN.Y 15.0405
R18070 XThC.XTBN.Y.n172 XThC.XTBN.Y 15.0405
R18071 XThC.XTBN.Y.n112 XThC.XTBN.Y 15.0405
R18072 XThC.XTBN.Y.n136 XThC.XTBN.Y 15.0405
R18073 XThC.XTBN.Y.n160 XThC.XTBN.Y 15.0405
R18074 XThC.XTBN.Y.n90 XThC.XTBN.Y.n89 13.8005
R18075 XThC.XTBN.Y.n64 XThC.XTBN.Y.n63 13.8005
R18076 XThC.XTBN.Y.n38 XThC.XTBN.Y.n37 13.8005
R18077 XThC.XTBN.Y.n77 XThC.XTBN.Y.n76 13.8005
R18078 XThC.XTBN.Y.n51 XThC.XTBN.Y.n50 13.8005
R18079 XThC.XTBN.Y.n25 XThC.XTBN.Y.n24 13.8005
R18080 XThC.XTBN.Y.n190 XThC.XTBN.Y 12.5445
R18081 XThC.XTBN.Y.n191 XThC.XTBN.Y 11.2645
R18082 XThC.XTBN.Y.n185 XThC.XTBN.Y.n184 9.2165
R18083 XThC.XTBN.Y.n185 XThC.XTBN.Y 7.9365
R18084 XThC.XTBN.Y.n96 XThC.XTBN.Y 6.7205
R18085 XThC.XTBN.Y.n119 XThC.XTBN.Y 6.7205
R18086 XThC.XTBN.Y.n143 XThC.XTBN.Y 6.7205
R18087 XThC.XTBN.Y.n167 XThC.XTBN.Y 6.7205
R18088 XThC.XTBN.Y.n107 XThC.XTBN.Y 6.7205
R18089 XThC.XTBN.Y.n131 XThC.XTBN.Y 6.7205
R18090 XThC.XTBN.Y.n155 XThC.XTBN.Y 6.7205
R18091 XThC.XTBN.Y.n93 XThC.XTBN.Y.n91 6.57323
R18092 XThC.XTBN.Y.n116 XThC.XTBN.Y.n114 6.57323
R18093 XThC.XTBN.Y.n140 XThC.XTBN.Y.n138 6.57323
R18094 XThC.XTBN.Y.n164 XThC.XTBN.Y.n162 6.57323
R18095 XThC.XTBN.Y.n104 XThC.XTBN.Y.n102 6.57323
R18096 XThC.XTBN.Y.n128 XThC.XTBN.Y.n126 6.57323
R18097 XThC.XTBN.Y.n152 XThC.XTBN.Y.n150 6.57323
R18098 XThC.XTBN.Y.n184 XThC.XTBN.Y 6.4005
R18099 XThC.XTBN.Y.n191 XThC.XTBN.Y 6.1445
R18100 XThC.XTBN.Y.n187 XThC.XTBN.Y.n186 5.74665
R18101 XThC.XTBN.Y.n186 XThC.XTBN.Y.n174 5.68319
R18102 XThC.XTBN.Y.n98 XThC.XTBN.Y.n97 5.11262
R18103 XThC.XTBN.Y.n121 XThC.XTBN.Y.n120 5.11262
R18104 XThC.XTBN.Y.n145 XThC.XTBN.Y.n144 5.11262
R18105 XThC.XTBN.Y.n169 XThC.XTBN.Y.n168 5.11262
R18106 XThC.XTBN.Y.n109 XThC.XTBN.Y.n108 5.11262
R18107 XThC.XTBN.Y.n133 XThC.XTBN.Y.n132 5.11262
R18108 XThC.XTBN.Y.n157 XThC.XTBN.Y.n156 5.11262
R18109 XThC.XTBN.Y.n190 XThC.XTBN.Y.n187 5.06717
R18110 XThC.XTBN.Y XThC.XTBN.Y.n190 4.8645
R18111 XThC.XTBN.Y XThC.XTBN.Y.n191 4.65505
R18112 XThC.XTBN.Y.n186 XThC.XTBN.Y.n185 4.6505
R18113 XThC.XTBN.Y.n89 XThC.XTBN.Y 4.6085
R18114 XThC.XTBN.Y.n63 XThC.XTBN.Y 4.6085
R18115 XThC.XTBN.Y.n37 XThC.XTBN.Y 4.6085
R18116 XThC.XTBN.Y.n12 XThC.XTBN.Y 4.6085
R18117 XThC.XTBN.Y.n76 XThC.XTBN.Y 4.6085
R18118 XThC.XTBN.Y.n50 XThC.XTBN.Y 4.6085
R18119 XThC.XTBN.Y.n24 XThC.XTBN.Y 4.6085
R18120 XThC.XTBN.Y.n179 XThC.XTBN.Y 4.3525
R18121 XThC.XTBN.Y.n85 XThC.XTBN.Y 3.5845
R18122 XThC.XTBN.Y.n59 XThC.XTBN.Y 3.5845
R18123 XThC.XTBN.Y.n33 XThC.XTBN.Y 3.5845
R18124 XThC.XTBN.Y.n8 XThC.XTBN.Y 3.5845
R18125 XThC.XTBN.Y.n72 XThC.XTBN.Y 3.5845
R18126 XThC.XTBN.Y.n46 XThC.XTBN.Y 3.5845
R18127 XThC.XTBN.Y.n20 XThC.XTBN.Y 3.5845
R18128 XThC.XTBN.Y XThC.XTBN.Y.n0 2.3045
R18129 XThC.XTBN.Y XThC.XTBN.Y.n178 2.3045
R18130 XThC.XTBN.Y XThC.XTBN.Y.n189 2.0485
R18131 XThC.XTBN.Y.n89 XThC.XTBN.Y.n88 1.7925
R18132 XThC.XTBN.Y.n63 XThC.XTBN.Y.n62 1.7925
R18133 XThC.XTBN.Y.n37 XThC.XTBN.Y.n36 1.7925
R18134 XThC.XTBN.Y.n12 XThC.XTBN.Y.n11 1.7925
R18135 XThC.XTBN.Y.n76 XThC.XTBN.Y.n75 1.7925
R18136 XThC.XTBN.Y.n50 XThC.XTBN.Y.n49 1.7925
R18137 XThC.XTBN.Y.n24 XThC.XTBN.Y.n23 1.7925
R18138 XThC.XTBN.Y.n174 XThC.XTBN.Y.n173 1.59665
R18139 XThC.XTBN.Y.n189 XThC.XTBN.Y 1.55202
R18140 XThC.XTBN.Y XThC.XTBN.Y.n84 1.5365
R18141 XThC.XTBN.Y XThC.XTBN.Y.n58 1.5365
R18142 XThC.XTBN.Y XThC.XTBN.Y.n32 1.5365
R18143 XThC.XTBN.Y XThC.XTBN.Y.n7 1.5365
R18144 XThC.XTBN.Y XThC.XTBN.Y.n71 1.5365
R18145 XThC.XTBN.Y XThC.XTBN.Y.n45 1.5365
R18146 XThC.XTBN.Y XThC.XTBN.Y.n19 1.5365
R18147 XThC.XTBN.Y.n149 XThC.XTBN.Y.n137 1.49088
R18148 XThC.XTBN.Y.n125 XThC.XTBN.Y.n113 1.49088
R18149 XThC.XTBN.Y.n173 XThC.XTBN.Y.n161 1.48608
R18150 XThC.XTBN.Y.n51 XThC.XTBN.Y.n38 1.46204
R18151 XThC.XTBN.Y.n77 XThC.XTBN.Y.n64 1.46204
R18152 XThC.XTBN.Y.n38 XThC.XTBN.Y.n25 1.15435
R18153 XThC.XTBN.Y.n64 XThC.XTBN.Y.n51 1.15435
R18154 XThC.XTBN.Y.n90 XThC.XTBN.Y.n77 1.15435
R18155 XThC.XTBN.Y.n174 XThC.XTBN.Y.n90 1.14473
R18156 XThC.XTBN.Y.n161 XThC.XTBN.Y.n149 1.13031
R18157 XThC.XTBN.Y.n137 XThC.XTBN.Y.n125 1.1255
R18158 XThC.XTBN.Y.n79 XThC.XTBN.Y 0.5125
R18159 XThC.XTBN.Y.n53 XThC.XTBN.Y 0.5125
R18160 XThC.XTBN.Y.n27 XThC.XTBN.Y 0.5125
R18161 XThC.XTBN.Y.n2 XThC.XTBN.Y 0.5125
R18162 XThC.XTBN.Y.n66 XThC.XTBN.Y 0.5125
R18163 XThC.XTBN.Y.n40 XThC.XTBN.Y 0.5125
R18164 XThC.XTBN.Y.n14 XThC.XTBN.Y 0.5125
R18165 XThC.Tn[6].n2 XThC.Tn[6].n1 332.332
R18166 XThC.Tn[6].n2 XThC.Tn[6].n0 296.493
R18167 XThC.Tn[6].n12 XThC.Tn[6].n10 161.406
R18168 XThC.Tn[6].n15 XThC.Tn[6].n13 161.406
R18169 XThC.Tn[6].n18 XThC.Tn[6].n16 161.406
R18170 XThC.Tn[6].n21 XThC.Tn[6].n19 161.406
R18171 XThC.Tn[6].n24 XThC.Tn[6].n22 161.406
R18172 XThC.Tn[6].n27 XThC.Tn[6].n25 161.406
R18173 XThC.Tn[6].n30 XThC.Tn[6].n28 161.406
R18174 XThC.Tn[6].n33 XThC.Tn[6].n31 161.406
R18175 XThC.Tn[6].n36 XThC.Tn[6].n34 161.406
R18176 XThC.Tn[6].n39 XThC.Tn[6].n37 161.406
R18177 XThC.Tn[6].n42 XThC.Tn[6].n40 161.406
R18178 XThC.Tn[6].n45 XThC.Tn[6].n43 161.406
R18179 XThC.Tn[6].n48 XThC.Tn[6].n46 161.406
R18180 XThC.Tn[6].n51 XThC.Tn[6].n49 161.406
R18181 XThC.Tn[6].n54 XThC.Tn[6].n52 161.406
R18182 XThC.Tn[6].n57 XThC.Tn[6].n55 161.406
R18183 XThC.Tn[6].n10 XThC.Tn[6].t26 161.202
R18184 XThC.Tn[6].n13 XThC.Tn[6].t13 161.202
R18185 XThC.Tn[6].n16 XThC.Tn[6].t17 161.202
R18186 XThC.Tn[6].n19 XThC.Tn[6].t18 161.202
R18187 XThC.Tn[6].n22 XThC.Tn[6].t37 161.202
R18188 XThC.Tn[6].n25 XThC.Tn[6].t38 161.202
R18189 XThC.Tn[6].n28 XThC.Tn[6].t22 161.202
R18190 XThC.Tn[6].n31 XThC.Tn[6].t29 161.202
R18191 XThC.Tn[6].n34 XThC.Tn[6].t31 161.202
R18192 XThC.Tn[6].n37 XThC.Tn[6].t19 161.202
R18193 XThC.Tn[6].n40 XThC.Tn[6].t21 161.202
R18194 XThC.Tn[6].n43 XThC.Tn[6].t32 161.202
R18195 XThC.Tn[6].n46 XThC.Tn[6].t41 161.202
R18196 XThC.Tn[6].n49 XThC.Tn[6].t43 161.202
R18197 XThC.Tn[6].n52 XThC.Tn[6].t24 161.202
R18198 XThC.Tn[6].n55 XThC.Tn[6].t34 161.202
R18199 XThC.Tn[6].n10 XThC.Tn[6].t23 145.137
R18200 XThC.Tn[6].n13 XThC.Tn[6].t40 145.137
R18201 XThC.Tn[6].n16 XThC.Tn[6].t42 145.137
R18202 XThC.Tn[6].n19 XThC.Tn[6].t12 145.137
R18203 XThC.Tn[6].n22 XThC.Tn[6].t33 145.137
R18204 XThC.Tn[6].n25 XThC.Tn[6].t35 145.137
R18205 XThC.Tn[6].n28 XThC.Tn[6].t16 145.137
R18206 XThC.Tn[6].n31 XThC.Tn[6].t25 145.137
R18207 XThC.Tn[6].n34 XThC.Tn[6].t27 145.137
R18208 XThC.Tn[6].n37 XThC.Tn[6].t14 145.137
R18209 XThC.Tn[6].n40 XThC.Tn[6].t15 145.137
R18210 XThC.Tn[6].n43 XThC.Tn[6].t28 145.137
R18211 XThC.Tn[6].n46 XThC.Tn[6].t36 145.137
R18212 XThC.Tn[6].n49 XThC.Tn[6].t39 145.137
R18213 XThC.Tn[6].n52 XThC.Tn[6].t20 145.137
R18214 XThC.Tn[6].n55 XThC.Tn[6].t30 145.137
R18215 XThC.Tn[6].n7 XThC.Tn[6].n6 135.248
R18216 XThC.Tn[6].n9 XThC.Tn[6].n3 98.982
R18217 XThC.Tn[6].n8 XThC.Tn[6].n4 98.982
R18218 XThC.Tn[6].n7 XThC.Tn[6].n5 98.982
R18219 XThC.Tn[6].n9 XThC.Tn[6].n8 36.2672
R18220 XThC.Tn[6].n8 XThC.Tn[6].n7 36.2672
R18221 XThC.Tn[6].n59 XThC.Tn[6].n9 32.6405
R18222 XThC.Tn[6].n1 XThC.Tn[6].t5 26.5955
R18223 XThC.Tn[6].n1 XThC.Tn[6].t4 26.5955
R18224 XThC.Tn[6].n0 XThC.Tn[6].t7 26.5955
R18225 XThC.Tn[6].n0 XThC.Tn[6].t6 26.5955
R18226 XThC.Tn[6].n3 XThC.Tn[6].t8 24.9236
R18227 XThC.Tn[6].n3 XThC.Tn[6].t11 24.9236
R18228 XThC.Tn[6].n4 XThC.Tn[6].t10 24.9236
R18229 XThC.Tn[6].n4 XThC.Tn[6].t9 24.9236
R18230 XThC.Tn[6].n5 XThC.Tn[6].t1 24.9236
R18231 XThC.Tn[6].n5 XThC.Tn[6].t0 24.9236
R18232 XThC.Tn[6].n6 XThC.Tn[6].t3 24.9236
R18233 XThC.Tn[6].n6 XThC.Tn[6].t2 24.9236
R18234 XThC.Tn[6].n60 XThC.Tn[6].n2 18.5605
R18235 XThC.Tn[6].n60 XThC.Tn[6].n59 11.5205
R18236 XThC.Tn[6].n59 XThC.Tn[6].n58 3.18344
R18237 XThC.Tn[6].n58 XThC.Tn[6] 3.09179
R18238 XThC.Tn[6].n15 XThC.Tn[6] 0.931056
R18239 XThC.Tn[6].n18 XThC.Tn[6] 0.931056
R18240 XThC.Tn[6].n21 XThC.Tn[6] 0.931056
R18241 XThC.Tn[6].n24 XThC.Tn[6] 0.931056
R18242 XThC.Tn[6].n27 XThC.Tn[6] 0.931056
R18243 XThC.Tn[6].n30 XThC.Tn[6] 0.931056
R18244 XThC.Tn[6].n33 XThC.Tn[6] 0.931056
R18245 XThC.Tn[6].n36 XThC.Tn[6] 0.931056
R18246 XThC.Tn[6].n39 XThC.Tn[6] 0.931056
R18247 XThC.Tn[6].n42 XThC.Tn[6] 0.931056
R18248 XThC.Tn[6].n45 XThC.Tn[6] 0.931056
R18249 XThC.Tn[6].n48 XThC.Tn[6] 0.931056
R18250 XThC.Tn[6].n51 XThC.Tn[6] 0.931056
R18251 XThC.Tn[6].n54 XThC.Tn[6] 0.931056
R18252 XThC.Tn[6].n57 XThC.Tn[6] 0.931056
R18253 XThC.Tn[6] XThC.Tn[6].n60 0.6405
R18254 XThC.Tn[6] XThC.Tn[6].n12 0.396333
R18255 XThC.Tn[6] XThC.Tn[6].n15 0.396333
R18256 XThC.Tn[6] XThC.Tn[6].n18 0.396333
R18257 XThC.Tn[6] XThC.Tn[6].n21 0.396333
R18258 XThC.Tn[6] XThC.Tn[6].n24 0.396333
R18259 XThC.Tn[6] XThC.Tn[6].n27 0.396333
R18260 XThC.Tn[6] XThC.Tn[6].n30 0.396333
R18261 XThC.Tn[6] XThC.Tn[6].n33 0.396333
R18262 XThC.Tn[6] XThC.Tn[6].n36 0.396333
R18263 XThC.Tn[6] XThC.Tn[6].n39 0.396333
R18264 XThC.Tn[6] XThC.Tn[6].n42 0.396333
R18265 XThC.Tn[6] XThC.Tn[6].n45 0.396333
R18266 XThC.Tn[6] XThC.Tn[6].n48 0.396333
R18267 XThC.Tn[6] XThC.Tn[6].n51 0.396333
R18268 XThC.Tn[6] XThC.Tn[6].n54 0.396333
R18269 XThC.Tn[6] XThC.Tn[6].n57 0.396333
R18270 XThC.Tn[6].n11 XThC.Tn[6] 0.104667
R18271 XThC.Tn[6].n14 XThC.Tn[6] 0.104667
R18272 XThC.Tn[6].n17 XThC.Tn[6] 0.104667
R18273 XThC.Tn[6].n20 XThC.Tn[6] 0.104667
R18274 XThC.Tn[6].n23 XThC.Tn[6] 0.104667
R18275 XThC.Tn[6].n26 XThC.Tn[6] 0.104667
R18276 XThC.Tn[6].n29 XThC.Tn[6] 0.104667
R18277 XThC.Tn[6].n32 XThC.Tn[6] 0.104667
R18278 XThC.Tn[6].n35 XThC.Tn[6] 0.104667
R18279 XThC.Tn[6].n38 XThC.Tn[6] 0.104667
R18280 XThC.Tn[6].n41 XThC.Tn[6] 0.104667
R18281 XThC.Tn[6].n44 XThC.Tn[6] 0.104667
R18282 XThC.Tn[6].n47 XThC.Tn[6] 0.104667
R18283 XThC.Tn[6].n50 XThC.Tn[6] 0.104667
R18284 XThC.Tn[6].n53 XThC.Tn[6] 0.104667
R18285 XThC.Tn[6].n56 XThC.Tn[6] 0.104667
R18286 XThC.Tn[6].n11 XThC.Tn[6] 0.0309878
R18287 XThC.Tn[6].n14 XThC.Tn[6] 0.0309878
R18288 XThC.Tn[6].n17 XThC.Tn[6] 0.0309878
R18289 XThC.Tn[6].n20 XThC.Tn[6] 0.0309878
R18290 XThC.Tn[6].n23 XThC.Tn[6] 0.0309878
R18291 XThC.Tn[6].n26 XThC.Tn[6] 0.0309878
R18292 XThC.Tn[6].n29 XThC.Tn[6] 0.0309878
R18293 XThC.Tn[6].n32 XThC.Tn[6] 0.0309878
R18294 XThC.Tn[6].n35 XThC.Tn[6] 0.0309878
R18295 XThC.Tn[6].n38 XThC.Tn[6] 0.0309878
R18296 XThC.Tn[6].n41 XThC.Tn[6] 0.0309878
R18297 XThC.Tn[6].n44 XThC.Tn[6] 0.0309878
R18298 XThC.Tn[6].n47 XThC.Tn[6] 0.0309878
R18299 XThC.Tn[6].n50 XThC.Tn[6] 0.0309878
R18300 XThC.Tn[6].n53 XThC.Tn[6] 0.0309878
R18301 XThC.Tn[6].n56 XThC.Tn[6] 0.0309878
R18302 XThC.Tn[6].n12 XThC.Tn[6].n11 0.027939
R18303 XThC.Tn[6].n15 XThC.Tn[6].n14 0.027939
R18304 XThC.Tn[6].n18 XThC.Tn[6].n17 0.027939
R18305 XThC.Tn[6].n21 XThC.Tn[6].n20 0.027939
R18306 XThC.Tn[6].n24 XThC.Tn[6].n23 0.027939
R18307 XThC.Tn[6].n27 XThC.Tn[6].n26 0.027939
R18308 XThC.Tn[6].n30 XThC.Tn[6].n29 0.027939
R18309 XThC.Tn[6].n33 XThC.Tn[6].n32 0.027939
R18310 XThC.Tn[6].n36 XThC.Tn[6].n35 0.027939
R18311 XThC.Tn[6].n39 XThC.Tn[6].n38 0.027939
R18312 XThC.Tn[6].n42 XThC.Tn[6].n41 0.027939
R18313 XThC.Tn[6].n45 XThC.Tn[6].n44 0.027939
R18314 XThC.Tn[6].n48 XThC.Tn[6].n47 0.027939
R18315 XThC.Tn[6].n51 XThC.Tn[6].n50 0.027939
R18316 XThC.Tn[6].n54 XThC.Tn[6].n53 0.027939
R18317 XThC.Tn[6].n57 XThC.Tn[6].n56 0.027939
R18318 XThC.Tn[6].n58 XThC.Tn[6] 0.0140108
R18319 XThR.Tn[9].n87 XThR.Tn[9].n86 256.104
R18320 XThR.Tn[9].n2 XThR.Tn[9].n0 243.68
R18321 XThR.Tn[9].n5 XThR.Tn[9].n3 241.847
R18322 XThR.Tn[9].n2 XThR.Tn[9].n1 205.28
R18323 XThR.Tn[9].n87 XThR.Tn[9].n85 202.094
R18324 XThR.Tn[9].n5 XThR.Tn[9].n4 185
R18325 XThR.Tn[9] XThR.Tn[9].n78 161.363
R18326 XThR.Tn[9] XThR.Tn[9].n73 161.363
R18327 XThR.Tn[9] XThR.Tn[9].n68 161.363
R18328 XThR.Tn[9] XThR.Tn[9].n63 161.363
R18329 XThR.Tn[9] XThR.Tn[9].n58 161.363
R18330 XThR.Tn[9] XThR.Tn[9].n53 161.363
R18331 XThR.Tn[9] XThR.Tn[9].n48 161.363
R18332 XThR.Tn[9] XThR.Tn[9].n43 161.363
R18333 XThR.Tn[9] XThR.Tn[9].n38 161.363
R18334 XThR.Tn[9] XThR.Tn[9].n33 161.363
R18335 XThR.Tn[9] XThR.Tn[9].n28 161.363
R18336 XThR.Tn[9] XThR.Tn[9].n23 161.363
R18337 XThR.Tn[9] XThR.Tn[9].n18 161.363
R18338 XThR.Tn[9] XThR.Tn[9].n13 161.363
R18339 XThR.Tn[9] XThR.Tn[9].n8 161.363
R18340 XThR.Tn[9] XThR.Tn[9].n6 161.363
R18341 XThR.Tn[9].n80 XThR.Tn[9].n79 161.3
R18342 XThR.Tn[9].n75 XThR.Tn[9].n74 161.3
R18343 XThR.Tn[9].n70 XThR.Tn[9].n69 161.3
R18344 XThR.Tn[9].n65 XThR.Tn[9].n64 161.3
R18345 XThR.Tn[9].n60 XThR.Tn[9].n59 161.3
R18346 XThR.Tn[9].n55 XThR.Tn[9].n54 161.3
R18347 XThR.Tn[9].n50 XThR.Tn[9].n49 161.3
R18348 XThR.Tn[9].n45 XThR.Tn[9].n44 161.3
R18349 XThR.Tn[9].n40 XThR.Tn[9].n39 161.3
R18350 XThR.Tn[9].n35 XThR.Tn[9].n34 161.3
R18351 XThR.Tn[9].n30 XThR.Tn[9].n29 161.3
R18352 XThR.Tn[9].n25 XThR.Tn[9].n24 161.3
R18353 XThR.Tn[9].n20 XThR.Tn[9].n19 161.3
R18354 XThR.Tn[9].n15 XThR.Tn[9].n14 161.3
R18355 XThR.Tn[9].n10 XThR.Tn[9].n9 161.3
R18356 XThR.Tn[9].n78 XThR.Tn[9].t63 161.106
R18357 XThR.Tn[9].n73 XThR.Tn[9].t69 161.106
R18358 XThR.Tn[9].n68 XThR.Tn[9].t47 161.106
R18359 XThR.Tn[9].n63 XThR.Tn[9].t34 161.106
R18360 XThR.Tn[9].n58 XThR.Tn[9].t62 161.106
R18361 XThR.Tn[9].n53 XThR.Tn[9].t24 161.106
R18362 XThR.Tn[9].n48 XThR.Tn[9].t66 161.106
R18363 XThR.Tn[9].n43 XThR.Tn[9].t45 161.106
R18364 XThR.Tn[9].n38 XThR.Tn[9].t32 161.106
R18365 XThR.Tn[9].n33 XThR.Tn[9].t37 161.106
R18366 XThR.Tn[9].n28 XThR.Tn[9].t23 161.106
R18367 XThR.Tn[9].n23 XThR.Tn[9].t46 161.106
R18368 XThR.Tn[9].n18 XThR.Tn[9].t21 161.106
R18369 XThR.Tn[9].n13 XThR.Tn[9].t64 161.106
R18370 XThR.Tn[9].n8 XThR.Tn[9].t28 161.106
R18371 XThR.Tn[9].n6 XThR.Tn[9].t71 161.106
R18372 XThR.Tn[9].n79 XThR.Tn[9].t54 159.978
R18373 XThR.Tn[9].n74 XThR.Tn[9].t61 159.978
R18374 XThR.Tn[9].n69 XThR.Tn[9].t43 159.978
R18375 XThR.Tn[9].n64 XThR.Tn[9].t27 159.978
R18376 XThR.Tn[9].n59 XThR.Tn[9].t52 159.978
R18377 XThR.Tn[9].n54 XThR.Tn[9].t18 159.978
R18378 XThR.Tn[9].n49 XThR.Tn[9].t60 159.978
R18379 XThR.Tn[9].n44 XThR.Tn[9].t40 159.978
R18380 XThR.Tn[9].n39 XThR.Tn[9].t25 159.978
R18381 XThR.Tn[9].n34 XThR.Tn[9].t33 159.978
R18382 XThR.Tn[9].n29 XThR.Tn[9].t16 159.978
R18383 XThR.Tn[9].n24 XThR.Tn[9].t42 159.978
R18384 XThR.Tn[9].n19 XThR.Tn[9].t15 159.978
R18385 XThR.Tn[9].n14 XThR.Tn[9].t59 159.978
R18386 XThR.Tn[9].n9 XThR.Tn[9].t19 159.978
R18387 XThR.Tn[9].n78 XThR.Tn[9].t49 145.038
R18388 XThR.Tn[9].n73 XThR.Tn[9].t14 145.038
R18389 XThR.Tn[9].n68 XThR.Tn[9].t57 145.038
R18390 XThR.Tn[9].n63 XThR.Tn[9].t38 145.038
R18391 XThR.Tn[9].n58 XThR.Tn[9].t70 145.038
R18392 XThR.Tn[9].n53 XThR.Tn[9].t48 145.038
R18393 XThR.Tn[9].n48 XThR.Tn[9].t58 145.038
R18394 XThR.Tn[9].n43 XThR.Tn[9].t39 145.038
R18395 XThR.Tn[9].n38 XThR.Tn[9].t36 145.038
R18396 XThR.Tn[9].n33 XThR.Tn[9].t67 145.038
R18397 XThR.Tn[9].n28 XThR.Tn[9].t31 145.038
R18398 XThR.Tn[9].n23 XThR.Tn[9].t56 145.038
R18399 XThR.Tn[9].n18 XThR.Tn[9].t29 145.038
R18400 XThR.Tn[9].n13 XThR.Tn[9].t72 145.038
R18401 XThR.Tn[9].n8 XThR.Tn[9].t35 145.038
R18402 XThR.Tn[9].n6 XThR.Tn[9].t17 145.038
R18403 XThR.Tn[9].n79 XThR.Tn[9].t68 143.911
R18404 XThR.Tn[9].n74 XThR.Tn[9].t30 143.911
R18405 XThR.Tn[9].n69 XThR.Tn[9].t12 143.911
R18406 XThR.Tn[9].n64 XThR.Tn[9].t53 143.911
R18407 XThR.Tn[9].n59 XThR.Tn[9].t22 143.911
R18408 XThR.Tn[9].n54 XThR.Tn[9].t65 143.911
R18409 XThR.Tn[9].n49 XThR.Tn[9].t13 143.911
R18410 XThR.Tn[9].n44 XThR.Tn[9].t55 143.911
R18411 XThR.Tn[9].n39 XThR.Tn[9].t51 143.911
R18412 XThR.Tn[9].n34 XThR.Tn[9].t20 143.911
R18413 XThR.Tn[9].n29 XThR.Tn[9].t44 143.911
R18414 XThR.Tn[9].n24 XThR.Tn[9].t73 143.911
R18415 XThR.Tn[9].n19 XThR.Tn[9].t41 143.911
R18416 XThR.Tn[9].n14 XThR.Tn[9].t26 143.911
R18417 XThR.Tn[9].n9 XThR.Tn[9].t50 143.911
R18418 XThR.Tn[9] XThR.Tn[9].n2 35.7652
R18419 XThR.Tn[9].n0 XThR.Tn[9].t2 26.5955
R18420 XThR.Tn[9].n0 XThR.Tn[9].t0 26.5955
R18421 XThR.Tn[9].n85 XThR.Tn[9].t10 26.5955
R18422 XThR.Tn[9].n85 XThR.Tn[9].t8 26.5955
R18423 XThR.Tn[9].n86 XThR.Tn[9].t11 26.5955
R18424 XThR.Tn[9].n86 XThR.Tn[9].t9 26.5955
R18425 XThR.Tn[9].n1 XThR.Tn[9].t3 26.5955
R18426 XThR.Tn[9].n1 XThR.Tn[9].t1 26.5955
R18427 XThR.Tn[9].n4 XThR.Tn[9].t4 24.9236
R18428 XThR.Tn[9].n4 XThR.Tn[9].t6 24.9236
R18429 XThR.Tn[9].n3 XThR.Tn[9].t5 24.9236
R18430 XThR.Tn[9].n3 XThR.Tn[9].t7 24.9236
R18431 XThR.Tn[9] XThR.Tn[9].n5 22.9615
R18432 XThR.Tn[9].n88 XThR.Tn[9].n87 13.5534
R18433 XThR.Tn[9].n84 XThR.Tn[9] 7.97984
R18434 XThR.Tn[9] XThR.Tn[9].n7 5.34038
R18435 XThR.Tn[9].n12 XThR.Tn[9].n11 4.5005
R18436 XThR.Tn[9].n17 XThR.Tn[9].n16 4.5005
R18437 XThR.Tn[9].n22 XThR.Tn[9].n21 4.5005
R18438 XThR.Tn[9].n27 XThR.Tn[9].n26 4.5005
R18439 XThR.Tn[9].n32 XThR.Tn[9].n31 4.5005
R18440 XThR.Tn[9].n37 XThR.Tn[9].n36 4.5005
R18441 XThR.Tn[9].n42 XThR.Tn[9].n41 4.5005
R18442 XThR.Tn[9].n47 XThR.Tn[9].n46 4.5005
R18443 XThR.Tn[9].n52 XThR.Tn[9].n51 4.5005
R18444 XThR.Tn[9].n57 XThR.Tn[9].n56 4.5005
R18445 XThR.Tn[9].n62 XThR.Tn[9].n61 4.5005
R18446 XThR.Tn[9].n67 XThR.Tn[9].n66 4.5005
R18447 XThR.Tn[9].n72 XThR.Tn[9].n71 4.5005
R18448 XThR.Tn[9].n77 XThR.Tn[9].n76 4.5005
R18449 XThR.Tn[9].n82 XThR.Tn[9].n81 4.5005
R18450 XThR.Tn[9].n83 XThR.Tn[9] 3.70586
R18451 XThR.Tn[9].n88 XThR.Tn[9].n84 2.99115
R18452 XThR.Tn[9].n88 XThR.Tn[9] 2.87153
R18453 XThR.Tn[9].n12 XThR.Tn[9] 2.52282
R18454 XThR.Tn[9].n17 XThR.Tn[9] 2.52282
R18455 XThR.Tn[9].n22 XThR.Tn[9] 2.52282
R18456 XThR.Tn[9].n27 XThR.Tn[9] 2.52282
R18457 XThR.Tn[9].n32 XThR.Tn[9] 2.52282
R18458 XThR.Tn[9].n37 XThR.Tn[9] 2.52282
R18459 XThR.Tn[9].n42 XThR.Tn[9] 2.52282
R18460 XThR.Tn[9].n47 XThR.Tn[9] 2.52282
R18461 XThR.Tn[9].n52 XThR.Tn[9] 2.52282
R18462 XThR.Tn[9].n57 XThR.Tn[9] 2.52282
R18463 XThR.Tn[9].n62 XThR.Tn[9] 2.52282
R18464 XThR.Tn[9].n67 XThR.Tn[9] 2.52282
R18465 XThR.Tn[9].n72 XThR.Tn[9] 2.52282
R18466 XThR.Tn[9].n77 XThR.Tn[9] 2.52282
R18467 XThR.Tn[9].n82 XThR.Tn[9] 2.52282
R18468 XThR.Tn[9].n84 XThR.Tn[9] 2.2734
R18469 XThR.Tn[9] XThR.Tn[9].n88 1.50638
R18470 XThR.Tn[9].n80 XThR.Tn[9] 1.08677
R18471 XThR.Tn[9].n75 XThR.Tn[9] 1.08677
R18472 XThR.Tn[9].n70 XThR.Tn[9] 1.08677
R18473 XThR.Tn[9].n65 XThR.Tn[9] 1.08677
R18474 XThR.Tn[9].n60 XThR.Tn[9] 1.08677
R18475 XThR.Tn[9].n55 XThR.Tn[9] 1.08677
R18476 XThR.Tn[9].n50 XThR.Tn[9] 1.08677
R18477 XThR.Tn[9].n45 XThR.Tn[9] 1.08677
R18478 XThR.Tn[9].n40 XThR.Tn[9] 1.08677
R18479 XThR.Tn[9].n35 XThR.Tn[9] 1.08677
R18480 XThR.Tn[9].n30 XThR.Tn[9] 1.08677
R18481 XThR.Tn[9].n25 XThR.Tn[9] 1.08677
R18482 XThR.Tn[9].n20 XThR.Tn[9] 1.08677
R18483 XThR.Tn[9].n15 XThR.Tn[9] 1.08677
R18484 XThR.Tn[9].n10 XThR.Tn[9] 1.08677
R18485 XThR.Tn[9] XThR.Tn[9].n12 0.839786
R18486 XThR.Tn[9] XThR.Tn[9].n17 0.839786
R18487 XThR.Tn[9] XThR.Tn[9].n22 0.839786
R18488 XThR.Tn[9] XThR.Tn[9].n27 0.839786
R18489 XThR.Tn[9] XThR.Tn[9].n32 0.839786
R18490 XThR.Tn[9] XThR.Tn[9].n37 0.839786
R18491 XThR.Tn[9] XThR.Tn[9].n42 0.839786
R18492 XThR.Tn[9] XThR.Tn[9].n47 0.839786
R18493 XThR.Tn[9] XThR.Tn[9].n52 0.839786
R18494 XThR.Tn[9] XThR.Tn[9].n57 0.839786
R18495 XThR.Tn[9] XThR.Tn[9].n62 0.839786
R18496 XThR.Tn[9] XThR.Tn[9].n67 0.839786
R18497 XThR.Tn[9] XThR.Tn[9].n72 0.839786
R18498 XThR.Tn[9] XThR.Tn[9].n77 0.839786
R18499 XThR.Tn[9] XThR.Tn[9].n82 0.839786
R18500 XThR.Tn[9].n7 XThR.Tn[9] 0.499542
R18501 XThR.Tn[9].n81 XThR.Tn[9] 0.063
R18502 XThR.Tn[9].n76 XThR.Tn[9] 0.063
R18503 XThR.Tn[9].n71 XThR.Tn[9] 0.063
R18504 XThR.Tn[9].n66 XThR.Tn[9] 0.063
R18505 XThR.Tn[9].n61 XThR.Tn[9] 0.063
R18506 XThR.Tn[9].n56 XThR.Tn[9] 0.063
R18507 XThR.Tn[9].n51 XThR.Tn[9] 0.063
R18508 XThR.Tn[9].n46 XThR.Tn[9] 0.063
R18509 XThR.Tn[9].n41 XThR.Tn[9] 0.063
R18510 XThR.Tn[9].n36 XThR.Tn[9] 0.063
R18511 XThR.Tn[9].n31 XThR.Tn[9] 0.063
R18512 XThR.Tn[9].n26 XThR.Tn[9] 0.063
R18513 XThR.Tn[9].n21 XThR.Tn[9] 0.063
R18514 XThR.Tn[9].n16 XThR.Tn[9] 0.063
R18515 XThR.Tn[9].n11 XThR.Tn[9] 0.063
R18516 XThR.Tn[9].n83 XThR.Tn[9] 0.0540714
R18517 XThR.Tn[9] XThR.Tn[9].n83 0.038
R18518 XThR.Tn[9].n7 XThR.Tn[9] 0.0143889
R18519 XThR.Tn[9].n81 XThR.Tn[9].n80 0.00771154
R18520 XThR.Tn[9].n76 XThR.Tn[9].n75 0.00771154
R18521 XThR.Tn[9].n71 XThR.Tn[9].n70 0.00771154
R18522 XThR.Tn[9].n66 XThR.Tn[9].n65 0.00771154
R18523 XThR.Tn[9].n61 XThR.Tn[9].n60 0.00771154
R18524 XThR.Tn[9].n56 XThR.Tn[9].n55 0.00771154
R18525 XThR.Tn[9].n51 XThR.Tn[9].n50 0.00771154
R18526 XThR.Tn[9].n46 XThR.Tn[9].n45 0.00771154
R18527 XThR.Tn[9].n41 XThR.Tn[9].n40 0.00771154
R18528 XThR.Tn[9].n36 XThR.Tn[9].n35 0.00771154
R18529 XThR.Tn[9].n31 XThR.Tn[9].n30 0.00771154
R18530 XThR.Tn[9].n26 XThR.Tn[9].n25 0.00771154
R18531 XThR.Tn[9].n21 XThR.Tn[9].n20 0.00771154
R18532 XThR.Tn[9].n16 XThR.Tn[9].n15 0.00771154
R18533 XThR.Tn[9].n11 XThR.Tn[9].n10 0.00771154
R18534 XThC.Tn[5].n2 XThC.Tn[5].n1 332.332
R18535 XThC.Tn[5].n2 XThC.Tn[5].n0 296.493
R18536 XThC.Tn[5].n12 XThC.Tn[5].n10 161.406
R18537 XThC.Tn[5].n15 XThC.Tn[5].n13 161.406
R18538 XThC.Tn[5].n18 XThC.Tn[5].n16 161.406
R18539 XThC.Tn[5].n21 XThC.Tn[5].n19 161.406
R18540 XThC.Tn[5].n24 XThC.Tn[5].n22 161.406
R18541 XThC.Tn[5].n27 XThC.Tn[5].n25 161.406
R18542 XThC.Tn[5].n30 XThC.Tn[5].n28 161.406
R18543 XThC.Tn[5].n33 XThC.Tn[5].n31 161.406
R18544 XThC.Tn[5].n36 XThC.Tn[5].n34 161.406
R18545 XThC.Tn[5].n39 XThC.Tn[5].n37 161.406
R18546 XThC.Tn[5].n42 XThC.Tn[5].n40 161.406
R18547 XThC.Tn[5].n45 XThC.Tn[5].n43 161.406
R18548 XThC.Tn[5].n48 XThC.Tn[5].n46 161.406
R18549 XThC.Tn[5].n51 XThC.Tn[5].n49 161.406
R18550 XThC.Tn[5].n54 XThC.Tn[5].n52 161.406
R18551 XThC.Tn[5].n57 XThC.Tn[5].n55 161.406
R18552 XThC.Tn[5].n10 XThC.Tn[5].t33 161.202
R18553 XThC.Tn[5].n13 XThC.Tn[5].t19 161.202
R18554 XThC.Tn[5].n16 XThC.Tn[5].t23 161.202
R18555 XThC.Tn[5].n19 XThC.Tn[5].t24 161.202
R18556 XThC.Tn[5].n22 XThC.Tn[5].t13 161.202
R18557 XThC.Tn[5].n25 XThC.Tn[5].t14 161.202
R18558 XThC.Tn[5].n28 XThC.Tn[5].t27 161.202
R18559 XThC.Tn[5].n31 XThC.Tn[5].t35 161.202
R18560 XThC.Tn[5].n34 XThC.Tn[5].t37 161.202
R18561 XThC.Tn[5].n37 XThC.Tn[5].t25 161.202
R18562 XThC.Tn[5].n40 XThC.Tn[5].t26 161.202
R18563 XThC.Tn[5].n43 XThC.Tn[5].t39 161.202
R18564 XThC.Tn[5].n46 XThC.Tn[5].t16 161.202
R18565 XThC.Tn[5].n49 XThC.Tn[5].t18 161.202
R18566 XThC.Tn[5].n52 XThC.Tn[5].t30 161.202
R18567 XThC.Tn[5].n55 XThC.Tn[5].t41 161.202
R18568 XThC.Tn[5].n10 XThC.Tn[5].t15 145.137
R18569 XThC.Tn[5].n13 XThC.Tn[5].t34 145.137
R18570 XThC.Tn[5].n16 XThC.Tn[5].t36 145.137
R18571 XThC.Tn[5].n19 XThC.Tn[5].t38 145.137
R18572 XThC.Tn[5].n22 XThC.Tn[5].t28 145.137
R18573 XThC.Tn[5].n25 XThC.Tn[5].t29 145.137
R18574 XThC.Tn[5].n28 XThC.Tn[5].t43 145.137
R18575 XThC.Tn[5].n31 XThC.Tn[5].t17 145.137
R18576 XThC.Tn[5].n34 XThC.Tn[5].t20 145.137
R18577 XThC.Tn[5].n37 XThC.Tn[5].t40 145.137
R18578 XThC.Tn[5].n40 XThC.Tn[5].t42 145.137
R18579 XThC.Tn[5].n43 XThC.Tn[5].t21 145.137
R18580 XThC.Tn[5].n46 XThC.Tn[5].t31 145.137
R18581 XThC.Tn[5].n49 XThC.Tn[5].t32 145.137
R18582 XThC.Tn[5].n52 XThC.Tn[5].t12 145.137
R18583 XThC.Tn[5].n55 XThC.Tn[5].t22 145.137
R18584 XThC.Tn[5].n7 XThC.Tn[5].n6 135.249
R18585 XThC.Tn[5].n9 XThC.Tn[5].n3 98.981
R18586 XThC.Tn[5].n8 XThC.Tn[5].n4 98.981
R18587 XThC.Tn[5].n7 XThC.Tn[5].n5 98.981
R18588 XThC.Tn[5].n9 XThC.Tn[5].n8 36.2672
R18589 XThC.Tn[5].n8 XThC.Tn[5].n7 36.2672
R18590 XThC.Tn[5].n59 XThC.Tn[5].n9 32.6405
R18591 XThC.Tn[5].n1 XThC.Tn[5].t9 26.5955
R18592 XThC.Tn[5].n1 XThC.Tn[5].t8 26.5955
R18593 XThC.Tn[5].n0 XThC.Tn[5].t11 26.5955
R18594 XThC.Tn[5].n0 XThC.Tn[5].t10 26.5955
R18595 XThC.Tn[5].n3 XThC.Tn[5].t5 24.9236
R18596 XThC.Tn[5].n3 XThC.Tn[5].t4 24.9236
R18597 XThC.Tn[5].n4 XThC.Tn[5].t7 24.9236
R18598 XThC.Tn[5].n4 XThC.Tn[5].t6 24.9236
R18599 XThC.Tn[5].n5 XThC.Tn[5].t2 24.9236
R18600 XThC.Tn[5].n5 XThC.Tn[5].t1 24.9236
R18601 XThC.Tn[5].n6 XThC.Tn[5].t0 24.9236
R18602 XThC.Tn[5].n6 XThC.Tn[5].t3 24.9236
R18603 XThC.Tn[5] XThC.Tn[5].n2 23.3605
R18604 XThC.Tn[5] XThC.Tn[5].n59 6.7205
R18605 XThC.Tn[5].n58 XThC.Tn[5] 3.62266
R18606 XThC.Tn[5].n59 XThC.Tn[5].n58 3.18437
R18607 XThC.Tn[5].n15 XThC.Tn[5] 0.931056
R18608 XThC.Tn[5].n18 XThC.Tn[5] 0.931056
R18609 XThC.Tn[5].n21 XThC.Tn[5] 0.931056
R18610 XThC.Tn[5].n24 XThC.Tn[5] 0.931056
R18611 XThC.Tn[5].n27 XThC.Tn[5] 0.931056
R18612 XThC.Tn[5].n30 XThC.Tn[5] 0.931056
R18613 XThC.Tn[5].n33 XThC.Tn[5] 0.931056
R18614 XThC.Tn[5].n36 XThC.Tn[5] 0.931056
R18615 XThC.Tn[5].n39 XThC.Tn[5] 0.931056
R18616 XThC.Tn[5].n42 XThC.Tn[5] 0.931056
R18617 XThC.Tn[5].n45 XThC.Tn[5] 0.931056
R18618 XThC.Tn[5].n48 XThC.Tn[5] 0.931056
R18619 XThC.Tn[5].n51 XThC.Tn[5] 0.931056
R18620 XThC.Tn[5].n54 XThC.Tn[5] 0.931056
R18621 XThC.Tn[5].n57 XThC.Tn[5] 0.931056
R18622 XThC.Tn[5] XThC.Tn[5].n12 0.396333
R18623 XThC.Tn[5] XThC.Tn[5].n15 0.396333
R18624 XThC.Tn[5] XThC.Tn[5].n18 0.396333
R18625 XThC.Tn[5] XThC.Tn[5].n21 0.396333
R18626 XThC.Tn[5] XThC.Tn[5].n24 0.396333
R18627 XThC.Tn[5] XThC.Tn[5].n27 0.396333
R18628 XThC.Tn[5] XThC.Tn[5].n30 0.396333
R18629 XThC.Tn[5] XThC.Tn[5].n33 0.396333
R18630 XThC.Tn[5] XThC.Tn[5].n36 0.396333
R18631 XThC.Tn[5] XThC.Tn[5].n39 0.396333
R18632 XThC.Tn[5] XThC.Tn[5].n42 0.396333
R18633 XThC.Tn[5] XThC.Tn[5].n45 0.396333
R18634 XThC.Tn[5] XThC.Tn[5].n48 0.396333
R18635 XThC.Tn[5] XThC.Tn[5].n51 0.396333
R18636 XThC.Tn[5] XThC.Tn[5].n54 0.396333
R18637 XThC.Tn[5] XThC.Tn[5].n57 0.396333
R18638 XThC.Tn[5].n11 XThC.Tn[5] 0.104667
R18639 XThC.Tn[5].n14 XThC.Tn[5] 0.104667
R18640 XThC.Tn[5].n17 XThC.Tn[5] 0.104667
R18641 XThC.Tn[5].n20 XThC.Tn[5] 0.104667
R18642 XThC.Tn[5].n23 XThC.Tn[5] 0.104667
R18643 XThC.Tn[5].n26 XThC.Tn[5] 0.104667
R18644 XThC.Tn[5].n29 XThC.Tn[5] 0.104667
R18645 XThC.Tn[5].n32 XThC.Tn[5] 0.104667
R18646 XThC.Tn[5].n35 XThC.Tn[5] 0.104667
R18647 XThC.Tn[5].n38 XThC.Tn[5] 0.104667
R18648 XThC.Tn[5].n41 XThC.Tn[5] 0.104667
R18649 XThC.Tn[5].n44 XThC.Tn[5] 0.104667
R18650 XThC.Tn[5].n47 XThC.Tn[5] 0.104667
R18651 XThC.Tn[5].n50 XThC.Tn[5] 0.104667
R18652 XThC.Tn[5].n53 XThC.Tn[5] 0.104667
R18653 XThC.Tn[5].n56 XThC.Tn[5] 0.104667
R18654 XThC.Tn[5].n11 XThC.Tn[5] 0.0309878
R18655 XThC.Tn[5].n14 XThC.Tn[5] 0.0309878
R18656 XThC.Tn[5].n17 XThC.Tn[5] 0.0309878
R18657 XThC.Tn[5].n20 XThC.Tn[5] 0.0309878
R18658 XThC.Tn[5].n23 XThC.Tn[5] 0.0309878
R18659 XThC.Tn[5].n26 XThC.Tn[5] 0.0309878
R18660 XThC.Tn[5].n29 XThC.Tn[5] 0.0309878
R18661 XThC.Tn[5].n32 XThC.Tn[5] 0.0309878
R18662 XThC.Tn[5].n35 XThC.Tn[5] 0.0309878
R18663 XThC.Tn[5].n38 XThC.Tn[5] 0.0309878
R18664 XThC.Tn[5].n41 XThC.Tn[5] 0.0309878
R18665 XThC.Tn[5].n44 XThC.Tn[5] 0.0309878
R18666 XThC.Tn[5].n47 XThC.Tn[5] 0.0309878
R18667 XThC.Tn[5].n50 XThC.Tn[5] 0.0309878
R18668 XThC.Tn[5].n53 XThC.Tn[5] 0.0309878
R18669 XThC.Tn[5].n56 XThC.Tn[5] 0.0309878
R18670 XThC.Tn[5].n12 XThC.Tn[5].n11 0.027939
R18671 XThC.Tn[5].n15 XThC.Tn[5].n14 0.027939
R18672 XThC.Tn[5].n18 XThC.Tn[5].n17 0.027939
R18673 XThC.Tn[5].n21 XThC.Tn[5].n20 0.027939
R18674 XThC.Tn[5].n24 XThC.Tn[5].n23 0.027939
R18675 XThC.Tn[5].n27 XThC.Tn[5].n26 0.027939
R18676 XThC.Tn[5].n30 XThC.Tn[5].n29 0.027939
R18677 XThC.Tn[5].n33 XThC.Tn[5].n32 0.027939
R18678 XThC.Tn[5].n36 XThC.Tn[5].n35 0.027939
R18679 XThC.Tn[5].n39 XThC.Tn[5].n38 0.027939
R18680 XThC.Tn[5].n42 XThC.Tn[5].n41 0.027939
R18681 XThC.Tn[5].n45 XThC.Tn[5].n44 0.027939
R18682 XThC.Tn[5].n48 XThC.Tn[5].n47 0.027939
R18683 XThC.Tn[5].n51 XThC.Tn[5].n50 0.027939
R18684 XThC.Tn[5].n54 XThC.Tn[5].n53 0.027939
R18685 XThC.Tn[5].n57 XThC.Tn[5].n56 0.027939
R18686 XThC.Tn[5].n58 XThC.Tn[5] 0.0129681
R18687 XThC.Tn[9].n54 XThC.Tn[9].n53 265.341
R18688 XThC.Tn[9].n58 XThC.Tn[9].n56 243.68
R18689 XThC.Tn[9].n2 XThC.Tn[9].n0 241.847
R18690 XThC.Tn[9].n58 XThC.Tn[9].n57 205.28
R18691 XThC.Tn[9].n54 XThC.Tn[9].n52 202.094
R18692 XThC.Tn[9].n2 XThC.Tn[9].n1 185
R18693 XThC.Tn[9].n5 XThC.Tn[9].n3 161.406
R18694 XThC.Tn[9].n8 XThC.Tn[9].n6 161.406
R18695 XThC.Tn[9].n11 XThC.Tn[9].n9 161.406
R18696 XThC.Tn[9].n14 XThC.Tn[9].n12 161.406
R18697 XThC.Tn[9].n17 XThC.Tn[9].n15 161.406
R18698 XThC.Tn[9].n20 XThC.Tn[9].n18 161.406
R18699 XThC.Tn[9].n23 XThC.Tn[9].n21 161.406
R18700 XThC.Tn[9].n26 XThC.Tn[9].n24 161.406
R18701 XThC.Tn[9].n29 XThC.Tn[9].n27 161.406
R18702 XThC.Tn[9].n32 XThC.Tn[9].n30 161.406
R18703 XThC.Tn[9].n35 XThC.Tn[9].n33 161.406
R18704 XThC.Tn[9].n38 XThC.Tn[9].n36 161.406
R18705 XThC.Tn[9].n41 XThC.Tn[9].n39 161.406
R18706 XThC.Tn[9].n44 XThC.Tn[9].n42 161.406
R18707 XThC.Tn[9].n47 XThC.Tn[9].n45 161.406
R18708 XThC.Tn[9].n50 XThC.Tn[9].n48 161.406
R18709 XThC.Tn[9].n3 XThC.Tn[9].t12 161.202
R18710 XThC.Tn[9].n6 XThC.Tn[9].t30 161.202
R18711 XThC.Tn[9].n9 XThC.Tn[9].t34 161.202
R18712 XThC.Tn[9].n12 XThC.Tn[9].t35 161.202
R18713 XThC.Tn[9].n15 XThC.Tn[9].t24 161.202
R18714 XThC.Tn[9].n18 XThC.Tn[9].t25 161.202
R18715 XThC.Tn[9].n21 XThC.Tn[9].t38 161.202
R18716 XThC.Tn[9].n24 XThC.Tn[9].t14 161.202
R18717 XThC.Tn[9].n27 XThC.Tn[9].t16 161.202
R18718 XThC.Tn[9].n30 XThC.Tn[9].t36 161.202
R18719 XThC.Tn[9].n33 XThC.Tn[9].t37 161.202
R18720 XThC.Tn[9].n36 XThC.Tn[9].t18 161.202
R18721 XThC.Tn[9].n39 XThC.Tn[9].t27 161.202
R18722 XThC.Tn[9].n42 XThC.Tn[9].t29 161.202
R18723 XThC.Tn[9].n45 XThC.Tn[9].t41 161.202
R18724 XThC.Tn[9].n48 XThC.Tn[9].t20 161.202
R18725 XThC.Tn[9].n3 XThC.Tn[9].t26 145.137
R18726 XThC.Tn[9].n6 XThC.Tn[9].t13 145.137
R18727 XThC.Tn[9].n9 XThC.Tn[9].t15 145.137
R18728 XThC.Tn[9].n12 XThC.Tn[9].t17 145.137
R18729 XThC.Tn[9].n15 XThC.Tn[9].t39 145.137
R18730 XThC.Tn[9].n18 XThC.Tn[9].t40 145.137
R18731 XThC.Tn[9].n21 XThC.Tn[9].t22 145.137
R18732 XThC.Tn[9].n24 XThC.Tn[9].t28 145.137
R18733 XThC.Tn[9].n27 XThC.Tn[9].t31 145.137
R18734 XThC.Tn[9].n30 XThC.Tn[9].t19 145.137
R18735 XThC.Tn[9].n33 XThC.Tn[9].t21 145.137
R18736 XThC.Tn[9].n36 XThC.Tn[9].t32 145.137
R18737 XThC.Tn[9].n39 XThC.Tn[9].t42 145.137
R18738 XThC.Tn[9].n42 XThC.Tn[9].t43 145.137
R18739 XThC.Tn[9].n45 XThC.Tn[9].t23 145.137
R18740 XThC.Tn[9].n48 XThC.Tn[9].t33 145.137
R18741 XThC.Tn[9].n53 XThC.Tn[9].t2 26.5955
R18742 XThC.Tn[9].n53 XThC.Tn[9].t1 26.5955
R18743 XThC.Tn[9].n56 XThC.Tn[9].t9 26.5955
R18744 XThC.Tn[9].n56 XThC.Tn[9].t8 26.5955
R18745 XThC.Tn[9].n57 XThC.Tn[9].t11 26.5955
R18746 XThC.Tn[9].n57 XThC.Tn[9].t10 26.5955
R18747 XThC.Tn[9].n52 XThC.Tn[9].t0 26.5955
R18748 XThC.Tn[9].n52 XThC.Tn[9].t3 26.5955
R18749 XThC.Tn[9].n1 XThC.Tn[9].t6 24.9236
R18750 XThC.Tn[9].n1 XThC.Tn[9].t7 24.9236
R18751 XThC.Tn[9].n0 XThC.Tn[9].t5 24.9236
R18752 XThC.Tn[9].n0 XThC.Tn[9].t4 24.9236
R18753 XThC.Tn[9] XThC.Tn[9].n58 22.9652
R18754 XThC.Tn[9] XThC.Tn[9].n2 18.8943
R18755 XThC.Tn[9].n55 XThC.Tn[9].n54 13.9299
R18756 XThC.Tn[9] XThC.Tn[9].n55 13.9299
R18757 XThC.Tn[9].n51 XThC.Tn[9] 6.34069
R18758 XThC.Tn[9].n51 XThC.Tn[9] 5.13485
R18759 XThC.Tn[9] XThC.Tn[9].n51 1.79489
R18760 XThC.Tn[9].n55 XThC.Tn[9] 1.19676
R18761 XThC.Tn[9].n8 XThC.Tn[9] 0.931056
R18762 XThC.Tn[9].n11 XThC.Tn[9] 0.931056
R18763 XThC.Tn[9].n14 XThC.Tn[9] 0.931056
R18764 XThC.Tn[9].n17 XThC.Tn[9] 0.931056
R18765 XThC.Tn[9].n20 XThC.Tn[9] 0.931056
R18766 XThC.Tn[9].n23 XThC.Tn[9] 0.931056
R18767 XThC.Tn[9].n26 XThC.Tn[9] 0.931056
R18768 XThC.Tn[9].n29 XThC.Tn[9] 0.931056
R18769 XThC.Tn[9].n32 XThC.Tn[9] 0.931056
R18770 XThC.Tn[9].n35 XThC.Tn[9] 0.931056
R18771 XThC.Tn[9].n38 XThC.Tn[9] 0.931056
R18772 XThC.Tn[9].n41 XThC.Tn[9] 0.931056
R18773 XThC.Tn[9].n44 XThC.Tn[9] 0.931056
R18774 XThC.Tn[9].n47 XThC.Tn[9] 0.931056
R18775 XThC.Tn[9].n50 XThC.Tn[9] 0.931056
R18776 XThC.Tn[9] XThC.Tn[9].n5 0.396333
R18777 XThC.Tn[9] XThC.Tn[9].n8 0.396333
R18778 XThC.Tn[9] XThC.Tn[9].n11 0.396333
R18779 XThC.Tn[9] XThC.Tn[9].n14 0.396333
R18780 XThC.Tn[9] XThC.Tn[9].n17 0.396333
R18781 XThC.Tn[9] XThC.Tn[9].n20 0.396333
R18782 XThC.Tn[9] XThC.Tn[9].n23 0.396333
R18783 XThC.Tn[9] XThC.Tn[9].n26 0.396333
R18784 XThC.Tn[9] XThC.Tn[9].n29 0.396333
R18785 XThC.Tn[9] XThC.Tn[9].n32 0.396333
R18786 XThC.Tn[9] XThC.Tn[9].n35 0.396333
R18787 XThC.Tn[9] XThC.Tn[9].n38 0.396333
R18788 XThC.Tn[9] XThC.Tn[9].n41 0.396333
R18789 XThC.Tn[9] XThC.Tn[9].n44 0.396333
R18790 XThC.Tn[9] XThC.Tn[9].n47 0.396333
R18791 XThC.Tn[9] XThC.Tn[9].n50 0.396333
R18792 XThC.Tn[9].n4 XThC.Tn[9] 0.104667
R18793 XThC.Tn[9].n7 XThC.Tn[9] 0.104667
R18794 XThC.Tn[9].n10 XThC.Tn[9] 0.104667
R18795 XThC.Tn[9].n13 XThC.Tn[9] 0.104667
R18796 XThC.Tn[9].n16 XThC.Tn[9] 0.104667
R18797 XThC.Tn[9].n19 XThC.Tn[9] 0.104667
R18798 XThC.Tn[9].n22 XThC.Tn[9] 0.104667
R18799 XThC.Tn[9].n25 XThC.Tn[9] 0.104667
R18800 XThC.Tn[9].n28 XThC.Tn[9] 0.104667
R18801 XThC.Tn[9].n31 XThC.Tn[9] 0.104667
R18802 XThC.Tn[9].n34 XThC.Tn[9] 0.104667
R18803 XThC.Tn[9].n37 XThC.Tn[9] 0.104667
R18804 XThC.Tn[9].n40 XThC.Tn[9] 0.104667
R18805 XThC.Tn[9].n43 XThC.Tn[9] 0.104667
R18806 XThC.Tn[9].n46 XThC.Tn[9] 0.104667
R18807 XThC.Tn[9].n49 XThC.Tn[9] 0.104667
R18808 XThC.Tn[9].n4 XThC.Tn[9] 0.0309878
R18809 XThC.Tn[9].n7 XThC.Tn[9] 0.0309878
R18810 XThC.Tn[9].n10 XThC.Tn[9] 0.0309878
R18811 XThC.Tn[9].n13 XThC.Tn[9] 0.0309878
R18812 XThC.Tn[9].n16 XThC.Tn[9] 0.0309878
R18813 XThC.Tn[9].n19 XThC.Tn[9] 0.0309878
R18814 XThC.Tn[9].n22 XThC.Tn[9] 0.0309878
R18815 XThC.Tn[9].n25 XThC.Tn[9] 0.0309878
R18816 XThC.Tn[9].n28 XThC.Tn[9] 0.0309878
R18817 XThC.Tn[9].n31 XThC.Tn[9] 0.0309878
R18818 XThC.Tn[9].n34 XThC.Tn[9] 0.0309878
R18819 XThC.Tn[9].n37 XThC.Tn[9] 0.0309878
R18820 XThC.Tn[9].n40 XThC.Tn[9] 0.0309878
R18821 XThC.Tn[9].n43 XThC.Tn[9] 0.0309878
R18822 XThC.Tn[9].n46 XThC.Tn[9] 0.0309878
R18823 XThC.Tn[9].n49 XThC.Tn[9] 0.0309878
R18824 XThC.Tn[9].n5 XThC.Tn[9].n4 0.027939
R18825 XThC.Tn[9].n8 XThC.Tn[9].n7 0.027939
R18826 XThC.Tn[9].n11 XThC.Tn[9].n10 0.027939
R18827 XThC.Tn[9].n14 XThC.Tn[9].n13 0.027939
R18828 XThC.Tn[9].n17 XThC.Tn[9].n16 0.027939
R18829 XThC.Tn[9].n20 XThC.Tn[9].n19 0.027939
R18830 XThC.Tn[9].n23 XThC.Tn[9].n22 0.027939
R18831 XThC.Tn[9].n26 XThC.Tn[9].n25 0.027939
R18832 XThC.Tn[9].n29 XThC.Tn[9].n28 0.027939
R18833 XThC.Tn[9].n32 XThC.Tn[9].n31 0.027939
R18834 XThC.Tn[9].n35 XThC.Tn[9].n34 0.027939
R18835 XThC.Tn[9].n38 XThC.Tn[9].n37 0.027939
R18836 XThC.Tn[9].n41 XThC.Tn[9].n40 0.027939
R18837 XThC.Tn[9].n44 XThC.Tn[9].n43 0.027939
R18838 XThC.Tn[9].n47 XThC.Tn[9].n46 0.027939
R18839 XThC.Tn[9].n50 XThC.Tn[9].n49 0.027939
R18840 XThC.Tn[11].n2 XThC.Tn[11].n1 265.341
R18841 XThC.Tn[11].n5 XThC.Tn[11].n3 243.68
R18842 XThC.Tn[11].n58 XThC.Tn[11].n57 241.847
R18843 XThC.Tn[11].n5 XThC.Tn[11].n4 205.28
R18844 XThC.Tn[11].n2 XThC.Tn[11].n0 202.094
R18845 XThC.Tn[11].n58 XThC.Tn[11].n56 185
R18846 XThC.Tn[11].n9 XThC.Tn[11].n7 161.406
R18847 XThC.Tn[11].n12 XThC.Tn[11].n10 161.406
R18848 XThC.Tn[11].n15 XThC.Tn[11].n13 161.406
R18849 XThC.Tn[11].n18 XThC.Tn[11].n16 161.406
R18850 XThC.Tn[11].n21 XThC.Tn[11].n19 161.406
R18851 XThC.Tn[11].n24 XThC.Tn[11].n22 161.406
R18852 XThC.Tn[11].n27 XThC.Tn[11].n25 161.406
R18853 XThC.Tn[11].n30 XThC.Tn[11].n28 161.406
R18854 XThC.Tn[11].n33 XThC.Tn[11].n31 161.406
R18855 XThC.Tn[11].n36 XThC.Tn[11].n34 161.406
R18856 XThC.Tn[11].n39 XThC.Tn[11].n37 161.406
R18857 XThC.Tn[11].n42 XThC.Tn[11].n40 161.406
R18858 XThC.Tn[11].n45 XThC.Tn[11].n43 161.406
R18859 XThC.Tn[11].n48 XThC.Tn[11].n46 161.406
R18860 XThC.Tn[11].n51 XThC.Tn[11].n49 161.406
R18861 XThC.Tn[11].n54 XThC.Tn[11].n52 161.406
R18862 XThC.Tn[11].n7 XThC.Tn[11].t18 161.202
R18863 XThC.Tn[11].n10 XThC.Tn[11].t35 161.202
R18864 XThC.Tn[11].n13 XThC.Tn[11].t37 161.202
R18865 XThC.Tn[11].n16 XThC.Tn[11].t39 161.202
R18866 XThC.Tn[11].n19 XThC.Tn[11].t28 161.202
R18867 XThC.Tn[11].n22 XThC.Tn[11].t29 161.202
R18868 XThC.Tn[11].n25 XThC.Tn[11].t42 161.202
R18869 XThC.Tn[11].n28 XThC.Tn[11].t19 161.202
R18870 XThC.Tn[11].n31 XThC.Tn[11].t21 161.202
R18871 XThC.Tn[11].n34 XThC.Tn[11].t40 161.202
R18872 XThC.Tn[11].n37 XThC.Tn[11].t41 161.202
R18873 XThC.Tn[11].n40 XThC.Tn[11].t22 161.202
R18874 XThC.Tn[11].n43 XThC.Tn[11].t30 161.202
R18875 XThC.Tn[11].n46 XThC.Tn[11].t33 161.202
R18876 XThC.Tn[11].n49 XThC.Tn[11].t14 161.202
R18877 XThC.Tn[11].n52 XThC.Tn[11].t24 161.202
R18878 XThC.Tn[11].n7 XThC.Tn[11].t20 145.137
R18879 XThC.Tn[11].n10 XThC.Tn[11].t38 145.137
R18880 XThC.Tn[11].n13 XThC.Tn[11].t43 145.137
R18881 XThC.Tn[11].n16 XThC.Tn[11].t12 145.137
R18882 XThC.Tn[11].n19 XThC.Tn[11].t31 145.137
R18883 XThC.Tn[11].n22 XThC.Tn[11].t32 145.137
R18884 XThC.Tn[11].n25 XThC.Tn[11].t16 145.137
R18885 XThC.Tn[11].n28 XThC.Tn[11].t23 145.137
R18886 XThC.Tn[11].n31 XThC.Tn[11].t25 145.137
R18887 XThC.Tn[11].n34 XThC.Tn[11].t13 145.137
R18888 XThC.Tn[11].n37 XThC.Tn[11].t15 145.137
R18889 XThC.Tn[11].n40 XThC.Tn[11].t26 145.137
R18890 XThC.Tn[11].n43 XThC.Tn[11].t34 145.137
R18891 XThC.Tn[11].n46 XThC.Tn[11].t36 145.137
R18892 XThC.Tn[11].n49 XThC.Tn[11].t17 145.137
R18893 XThC.Tn[11].n52 XThC.Tn[11].t27 145.137
R18894 XThC.Tn[11].n1 XThC.Tn[11].t3 26.5955
R18895 XThC.Tn[11].n1 XThC.Tn[11].t1 26.5955
R18896 XThC.Tn[11].n0 XThC.Tn[11].t11 26.5955
R18897 XThC.Tn[11].n0 XThC.Tn[11].t8 26.5955
R18898 XThC.Tn[11].n3 XThC.Tn[11].t4 26.5955
R18899 XThC.Tn[11].n3 XThC.Tn[11].t7 26.5955
R18900 XThC.Tn[11].n4 XThC.Tn[11].t6 26.5955
R18901 XThC.Tn[11].n4 XThC.Tn[11].t5 26.5955
R18902 XThC.Tn[11].n56 XThC.Tn[11].t2 24.9236
R18903 XThC.Tn[11].n56 XThC.Tn[11].t10 24.9236
R18904 XThC.Tn[11].n57 XThC.Tn[11].t0 24.9236
R18905 XThC.Tn[11].n57 XThC.Tn[11].t9 24.9236
R18906 XThC.Tn[11] XThC.Tn[11].n5 22.9652
R18907 XThC.Tn[11] XThC.Tn[11].n58 18.8943
R18908 XThC.Tn[11].n6 XThC.Tn[11].n2 13.9299
R18909 XThC.Tn[11].n6 XThC.Tn[11] 13.9299
R18910 XThC.Tn[11] XThC.Tn[11].n55 6.34069
R18911 XThC.Tn[11].n55 XThC.Tn[11] 5.13485
R18912 XThC.Tn[11].n55 XThC.Tn[11] 1.79489
R18913 XThC.Tn[11] XThC.Tn[11].n6 1.19676
R18914 XThC.Tn[11].n12 XThC.Tn[11] 0.931056
R18915 XThC.Tn[11].n15 XThC.Tn[11] 0.931056
R18916 XThC.Tn[11].n18 XThC.Tn[11] 0.931056
R18917 XThC.Tn[11].n21 XThC.Tn[11] 0.931056
R18918 XThC.Tn[11].n24 XThC.Tn[11] 0.931056
R18919 XThC.Tn[11].n27 XThC.Tn[11] 0.931056
R18920 XThC.Tn[11].n30 XThC.Tn[11] 0.931056
R18921 XThC.Tn[11].n33 XThC.Tn[11] 0.931056
R18922 XThC.Tn[11].n36 XThC.Tn[11] 0.931056
R18923 XThC.Tn[11].n39 XThC.Tn[11] 0.931056
R18924 XThC.Tn[11].n42 XThC.Tn[11] 0.931056
R18925 XThC.Tn[11].n45 XThC.Tn[11] 0.931056
R18926 XThC.Tn[11].n48 XThC.Tn[11] 0.931056
R18927 XThC.Tn[11].n51 XThC.Tn[11] 0.931056
R18928 XThC.Tn[11].n54 XThC.Tn[11] 0.931056
R18929 XThC.Tn[11] XThC.Tn[11].n9 0.396333
R18930 XThC.Tn[11] XThC.Tn[11].n12 0.396333
R18931 XThC.Tn[11] XThC.Tn[11].n15 0.396333
R18932 XThC.Tn[11] XThC.Tn[11].n18 0.396333
R18933 XThC.Tn[11] XThC.Tn[11].n21 0.396333
R18934 XThC.Tn[11] XThC.Tn[11].n24 0.396333
R18935 XThC.Tn[11] XThC.Tn[11].n27 0.396333
R18936 XThC.Tn[11] XThC.Tn[11].n30 0.396333
R18937 XThC.Tn[11] XThC.Tn[11].n33 0.396333
R18938 XThC.Tn[11] XThC.Tn[11].n36 0.396333
R18939 XThC.Tn[11] XThC.Tn[11].n39 0.396333
R18940 XThC.Tn[11] XThC.Tn[11].n42 0.396333
R18941 XThC.Tn[11] XThC.Tn[11].n45 0.396333
R18942 XThC.Tn[11] XThC.Tn[11].n48 0.396333
R18943 XThC.Tn[11] XThC.Tn[11].n51 0.396333
R18944 XThC.Tn[11] XThC.Tn[11].n54 0.396333
R18945 XThC.Tn[11].n8 XThC.Tn[11] 0.104667
R18946 XThC.Tn[11].n11 XThC.Tn[11] 0.104667
R18947 XThC.Tn[11].n14 XThC.Tn[11] 0.104667
R18948 XThC.Tn[11].n17 XThC.Tn[11] 0.104667
R18949 XThC.Tn[11].n20 XThC.Tn[11] 0.104667
R18950 XThC.Tn[11].n23 XThC.Tn[11] 0.104667
R18951 XThC.Tn[11].n26 XThC.Tn[11] 0.104667
R18952 XThC.Tn[11].n29 XThC.Tn[11] 0.104667
R18953 XThC.Tn[11].n32 XThC.Tn[11] 0.104667
R18954 XThC.Tn[11].n35 XThC.Tn[11] 0.104667
R18955 XThC.Tn[11].n38 XThC.Tn[11] 0.104667
R18956 XThC.Tn[11].n41 XThC.Tn[11] 0.104667
R18957 XThC.Tn[11].n44 XThC.Tn[11] 0.104667
R18958 XThC.Tn[11].n47 XThC.Tn[11] 0.104667
R18959 XThC.Tn[11].n50 XThC.Tn[11] 0.104667
R18960 XThC.Tn[11].n53 XThC.Tn[11] 0.104667
R18961 XThC.Tn[11].n8 XThC.Tn[11] 0.0309878
R18962 XThC.Tn[11].n11 XThC.Tn[11] 0.0309878
R18963 XThC.Tn[11].n14 XThC.Tn[11] 0.0309878
R18964 XThC.Tn[11].n17 XThC.Tn[11] 0.0309878
R18965 XThC.Tn[11].n20 XThC.Tn[11] 0.0309878
R18966 XThC.Tn[11].n23 XThC.Tn[11] 0.0309878
R18967 XThC.Tn[11].n26 XThC.Tn[11] 0.0309878
R18968 XThC.Tn[11].n29 XThC.Tn[11] 0.0309878
R18969 XThC.Tn[11].n32 XThC.Tn[11] 0.0309878
R18970 XThC.Tn[11].n35 XThC.Tn[11] 0.0309878
R18971 XThC.Tn[11].n38 XThC.Tn[11] 0.0309878
R18972 XThC.Tn[11].n41 XThC.Tn[11] 0.0309878
R18973 XThC.Tn[11].n44 XThC.Tn[11] 0.0309878
R18974 XThC.Tn[11].n47 XThC.Tn[11] 0.0309878
R18975 XThC.Tn[11].n50 XThC.Tn[11] 0.0309878
R18976 XThC.Tn[11].n53 XThC.Tn[11] 0.0309878
R18977 XThC.Tn[11].n9 XThC.Tn[11].n8 0.027939
R18978 XThC.Tn[11].n12 XThC.Tn[11].n11 0.027939
R18979 XThC.Tn[11].n15 XThC.Tn[11].n14 0.027939
R18980 XThC.Tn[11].n18 XThC.Tn[11].n17 0.027939
R18981 XThC.Tn[11].n21 XThC.Tn[11].n20 0.027939
R18982 XThC.Tn[11].n24 XThC.Tn[11].n23 0.027939
R18983 XThC.Tn[11].n27 XThC.Tn[11].n26 0.027939
R18984 XThC.Tn[11].n30 XThC.Tn[11].n29 0.027939
R18985 XThC.Tn[11].n33 XThC.Tn[11].n32 0.027939
R18986 XThC.Tn[11].n36 XThC.Tn[11].n35 0.027939
R18987 XThC.Tn[11].n39 XThC.Tn[11].n38 0.027939
R18988 XThC.Tn[11].n42 XThC.Tn[11].n41 0.027939
R18989 XThC.Tn[11].n45 XThC.Tn[11].n44 0.027939
R18990 XThC.Tn[11].n48 XThC.Tn[11].n47 0.027939
R18991 XThC.Tn[11].n51 XThC.Tn[11].n50 0.027939
R18992 XThC.Tn[11].n54 XThC.Tn[11].n53 0.027939
R18993 XThC.Tn[12].n5 XThC.Tn[12].n4 256.104
R18994 XThC.Tn[12].n8 XThC.Tn[12].n6 243.68
R18995 XThC.Tn[12].n2 XThC.Tn[12].n1 241.847
R18996 XThC.Tn[12].n8 XThC.Tn[12].n7 205.28
R18997 XThC.Tn[12].n5 XThC.Tn[12].n3 202.095
R18998 XThC.Tn[12].n2 XThC.Tn[12].n0 185
R18999 XThC.Tn[12].n12 XThC.Tn[12].n10 161.406
R19000 XThC.Tn[12].n15 XThC.Tn[12].n13 161.406
R19001 XThC.Tn[12].n18 XThC.Tn[12].n16 161.406
R19002 XThC.Tn[12].n21 XThC.Tn[12].n19 161.406
R19003 XThC.Tn[12].n24 XThC.Tn[12].n22 161.406
R19004 XThC.Tn[12].n27 XThC.Tn[12].n25 161.406
R19005 XThC.Tn[12].n30 XThC.Tn[12].n28 161.406
R19006 XThC.Tn[12].n33 XThC.Tn[12].n31 161.406
R19007 XThC.Tn[12].n36 XThC.Tn[12].n34 161.406
R19008 XThC.Tn[12].n39 XThC.Tn[12].n37 161.406
R19009 XThC.Tn[12].n42 XThC.Tn[12].n40 161.406
R19010 XThC.Tn[12].n45 XThC.Tn[12].n43 161.406
R19011 XThC.Tn[12].n48 XThC.Tn[12].n46 161.406
R19012 XThC.Tn[12].n51 XThC.Tn[12].n49 161.406
R19013 XThC.Tn[12].n54 XThC.Tn[12].n52 161.406
R19014 XThC.Tn[12].n57 XThC.Tn[12].n55 161.406
R19015 XThC.Tn[12].n10 XThC.Tn[12].t35 161.202
R19016 XThC.Tn[12].n13 XThC.Tn[12].t20 161.202
R19017 XThC.Tn[12].n16 XThC.Tn[12].t22 161.202
R19018 XThC.Tn[12].n19 XThC.Tn[12].t24 161.202
R19019 XThC.Tn[12].n22 XThC.Tn[12].t13 161.202
R19020 XThC.Tn[12].n25 XThC.Tn[12].t14 161.202
R19021 XThC.Tn[12].n28 XThC.Tn[12].t27 161.202
R19022 XThC.Tn[12].n31 XThC.Tn[12].t36 161.202
R19023 XThC.Tn[12].n34 XThC.Tn[12].t38 161.202
R19024 XThC.Tn[12].n37 XThC.Tn[12].t25 161.202
R19025 XThC.Tn[12].n40 XThC.Tn[12].t26 161.202
R19026 XThC.Tn[12].n43 XThC.Tn[12].t39 161.202
R19027 XThC.Tn[12].n46 XThC.Tn[12].t15 161.202
R19028 XThC.Tn[12].n49 XThC.Tn[12].t18 161.202
R19029 XThC.Tn[12].n52 XThC.Tn[12].t31 161.202
R19030 XThC.Tn[12].n55 XThC.Tn[12].t41 161.202
R19031 XThC.Tn[12].n10 XThC.Tn[12].t37 145.137
R19032 XThC.Tn[12].n13 XThC.Tn[12].t23 145.137
R19033 XThC.Tn[12].n16 XThC.Tn[12].t28 145.137
R19034 XThC.Tn[12].n19 XThC.Tn[12].t29 145.137
R19035 XThC.Tn[12].n22 XThC.Tn[12].t16 145.137
R19036 XThC.Tn[12].n25 XThC.Tn[12].t17 145.137
R19037 XThC.Tn[12].n28 XThC.Tn[12].t33 145.137
R19038 XThC.Tn[12].n31 XThC.Tn[12].t40 145.137
R19039 XThC.Tn[12].n34 XThC.Tn[12].t42 145.137
R19040 XThC.Tn[12].n37 XThC.Tn[12].t30 145.137
R19041 XThC.Tn[12].n40 XThC.Tn[12].t32 145.137
R19042 XThC.Tn[12].n43 XThC.Tn[12].t43 145.137
R19043 XThC.Tn[12].n46 XThC.Tn[12].t19 145.137
R19044 XThC.Tn[12].n49 XThC.Tn[12].t21 145.137
R19045 XThC.Tn[12].n52 XThC.Tn[12].t34 145.137
R19046 XThC.Tn[12].n55 XThC.Tn[12].t12 145.137
R19047 XThC.Tn[12].n3 XThC.Tn[12].t5 26.5955
R19048 XThC.Tn[12].n3 XThC.Tn[12].t6 26.5955
R19049 XThC.Tn[12].n4 XThC.Tn[12].t4 26.5955
R19050 XThC.Tn[12].n4 XThC.Tn[12].t7 26.5955
R19051 XThC.Tn[12].n6 XThC.Tn[12].t9 26.5955
R19052 XThC.Tn[12].n6 XThC.Tn[12].t8 26.5955
R19053 XThC.Tn[12].n7 XThC.Tn[12].t11 26.5955
R19054 XThC.Tn[12].n7 XThC.Tn[12].t10 26.5955
R19055 XThC.Tn[12].n0 XThC.Tn[12].t1 24.9236
R19056 XThC.Tn[12].n0 XThC.Tn[12].t0 24.9236
R19057 XThC.Tn[12].n1 XThC.Tn[12].t3 24.9236
R19058 XThC.Tn[12].n1 XThC.Tn[12].t2 24.9236
R19059 XThC.Tn[12] XThC.Tn[12].n8 22.9652
R19060 XThC.Tn[12] XThC.Tn[12].n2 22.9615
R19061 XThC.Tn[12].n9 XThC.Tn[12].n5 13.9299
R19062 XThC.Tn[12].n9 XThC.Tn[12] 13.9299
R19063 XThC.Tn[12].n59 XThC.Tn[12].n58 5.13244
R19064 XThC.Tn[12].n58 XThC.Tn[12] 3.8444
R19065 XThC.Tn[12].n59 XThC.Tn[12].n9 2.99115
R19066 XThC.Tn[12].n9 XThC.Tn[12] 2.87153
R19067 XThC.Tn[12] XThC.Tn[12].n59 2.2734
R19068 XThC.Tn[12].n15 XThC.Tn[12] 0.931056
R19069 XThC.Tn[12].n18 XThC.Tn[12] 0.931056
R19070 XThC.Tn[12].n21 XThC.Tn[12] 0.931056
R19071 XThC.Tn[12].n24 XThC.Tn[12] 0.931056
R19072 XThC.Tn[12].n27 XThC.Tn[12] 0.931056
R19073 XThC.Tn[12].n30 XThC.Tn[12] 0.931056
R19074 XThC.Tn[12].n33 XThC.Tn[12] 0.931056
R19075 XThC.Tn[12].n36 XThC.Tn[12] 0.931056
R19076 XThC.Tn[12].n39 XThC.Tn[12] 0.931056
R19077 XThC.Tn[12].n42 XThC.Tn[12] 0.931056
R19078 XThC.Tn[12].n45 XThC.Tn[12] 0.931056
R19079 XThC.Tn[12].n48 XThC.Tn[12] 0.931056
R19080 XThC.Tn[12].n51 XThC.Tn[12] 0.931056
R19081 XThC.Tn[12].n54 XThC.Tn[12] 0.931056
R19082 XThC.Tn[12].n57 XThC.Tn[12] 0.931056
R19083 XThC.Tn[12] XThC.Tn[12].n12 0.396333
R19084 XThC.Tn[12] XThC.Tn[12].n15 0.396333
R19085 XThC.Tn[12] XThC.Tn[12].n18 0.396333
R19086 XThC.Tn[12] XThC.Tn[12].n21 0.396333
R19087 XThC.Tn[12] XThC.Tn[12].n24 0.396333
R19088 XThC.Tn[12] XThC.Tn[12].n27 0.396333
R19089 XThC.Tn[12] XThC.Tn[12].n30 0.396333
R19090 XThC.Tn[12] XThC.Tn[12].n33 0.396333
R19091 XThC.Tn[12] XThC.Tn[12].n36 0.396333
R19092 XThC.Tn[12] XThC.Tn[12].n39 0.396333
R19093 XThC.Tn[12] XThC.Tn[12].n42 0.396333
R19094 XThC.Tn[12] XThC.Tn[12].n45 0.396333
R19095 XThC.Tn[12] XThC.Tn[12].n48 0.396333
R19096 XThC.Tn[12] XThC.Tn[12].n51 0.396333
R19097 XThC.Tn[12] XThC.Tn[12].n54 0.396333
R19098 XThC.Tn[12] XThC.Tn[12].n57 0.396333
R19099 XThC.Tn[12].n11 XThC.Tn[12] 0.104667
R19100 XThC.Tn[12].n14 XThC.Tn[12] 0.104667
R19101 XThC.Tn[12].n17 XThC.Tn[12] 0.104667
R19102 XThC.Tn[12].n20 XThC.Tn[12] 0.104667
R19103 XThC.Tn[12].n23 XThC.Tn[12] 0.104667
R19104 XThC.Tn[12].n26 XThC.Tn[12] 0.104667
R19105 XThC.Tn[12].n29 XThC.Tn[12] 0.104667
R19106 XThC.Tn[12].n32 XThC.Tn[12] 0.104667
R19107 XThC.Tn[12].n35 XThC.Tn[12] 0.104667
R19108 XThC.Tn[12].n38 XThC.Tn[12] 0.104667
R19109 XThC.Tn[12].n41 XThC.Tn[12] 0.104667
R19110 XThC.Tn[12].n44 XThC.Tn[12] 0.104667
R19111 XThC.Tn[12].n47 XThC.Tn[12] 0.104667
R19112 XThC.Tn[12].n50 XThC.Tn[12] 0.104667
R19113 XThC.Tn[12].n53 XThC.Tn[12] 0.104667
R19114 XThC.Tn[12].n56 XThC.Tn[12] 0.104667
R19115 XThC.Tn[12].n11 XThC.Tn[12] 0.0309878
R19116 XThC.Tn[12].n14 XThC.Tn[12] 0.0309878
R19117 XThC.Tn[12].n17 XThC.Tn[12] 0.0309878
R19118 XThC.Tn[12].n20 XThC.Tn[12] 0.0309878
R19119 XThC.Tn[12].n23 XThC.Tn[12] 0.0309878
R19120 XThC.Tn[12].n26 XThC.Tn[12] 0.0309878
R19121 XThC.Tn[12].n29 XThC.Tn[12] 0.0309878
R19122 XThC.Tn[12].n32 XThC.Tn[12] 0.0309878
R19123 XThC.Tn[12].n35 XThC.Tn[12] 0.0309878
R19124 XThC.Tn[12].n38 XThC.Tn[12] 0.0309878
R19125 XThC.Tn[12].n41 XThC.Tn[12] 0.0309878
R19126 XThC.Tn[12].n44 XThC.Tn[12] 0.0309878
R19127 XThC.Tn[12].n47 XThC.Tn[12] 0.0309878
R19128 XThC.Tn[12].n50 XThC.Tn[12] 0.0309878
R19129 XThC.Tn[12].n53 XThC.Tn[12] 0.0309878
R19130 XThC.Tn[12].n56 XThC.Tn[12] 0.0309878
R19131 XThC.Tn[12].n12 XThC.Tn[12].n11 0.027939
R19132 XThC.Tn[12].n15 XThC.Tn[12].n14 0.027939
R19133 XThC.Tn[12].n18 XThC.Tn[12].n17 0.027939
R19134 XThC.Tn[12].n21 XThC.Tn[12].n20 0.027939
R19135 XThC.Tn[12].n24 XThC.Tn[12].n23 0.027939
R19136 XThC.Tn[12].n27 XThC.Tn[12].n26 0.027939
R19137 XThC.Tn[12].n30 XThC.Tn[12].n29 0.027939
R19138 XThC.Tn[12].n33 XThC.Tn[12].n32 0.027939
R19139 XThC.Tn[12].n36 XThC.Tn[12].n35 0.027939
R19140 XThC.Tn[12].n39 XThC.Tn[12].n38 0.027939
R19141 XThC.Tn[12].n42 XThC.Tn[12].n41 0.027939
R19142 XThC.Tn[12].n45 XThC.Tn[12].n44 0.027939
R19143 XThC.Tn[12].n48 XThC.Tn[12].n47 0.027939
R19144 XThC.Tn[12].n51 XThC.Tn[12].n50 0.027939
R19145 XThC.Tn[12].n54 XThC.Tn[12].n53 0.027939
R19146 XThC.Tn[12].n57 XThC.Tn[12].n56 0.027939
R19147 XThC.Tn[12].n58 XThC.Tn[12] 0.00316553
R19148 XThC.Tn[13].n2 XThC.Tn[13].n1 265.341
R19149 XThC.Tn[13].n5 XThC.Tn[13].n3 243.68
R19150 XThC.Tn[13].n59 XThC.Tn[13].n58 241.847
R19151 XThC.Tn[13].n5 XThC.Tn[13].n4 205.28
R19152 XThC.Tn[13].n2 XThC.Tn[13].n0 202.094
R19153 XThC.Tn[13].n59 XThC.Tn[13].n57 185
R19154 XThC.Tn[13].n9 XThC.Tn[13].n7 161.406
R19155 XThC.Tn[13].n12 XThC.Tn[13].n10 161.406
R19156 XThC.Tn[13].n15 XThC.Tn[13].n13 161.406
R19157 XThC.Tn[13].n18 XThC.Tn[13].n16 161.406
R19158 XThC.Tn[13].n21 XThC.Tn[13].n19 161.406
R19159 XThC.Tn[13].n24 XThC.Tn[13].n22 161.406
R19160 XThC.Tn[13].n27 XThC.Tn[13].n25 161.406
R19161 XThC.Tn[13].n30 XThC.Tn[13].n28 161.406
R19162 XThC.Tn[13].n33 XThC.Tn[13].n31 161.406
R19163 XThC.Tn[13].n36 XThC.Tn[13].n34 161.406
R19164 XThC.Tn[13].n39 XThC.Tn[13].n37 161.406
R19165 XThC.Tn[13].n42 XThC.Tn[13].n40 161.406
R19166 XThC.Tn[13].n45 XThC.Tn[13].n43 161.406
R19167 XThC.Tn[13].n48 XThC.Tn[13].n46 161.406
R19168 XThC.Tn[13].n51 XThC.Tn[13].n49 161.406
R19169 XThC.Tn[13].n54 XThC.Tn[13].n52 161.406
R19170 XThC.Tn[13].n7 XThC.Tn[13].t27 161.202
R19171 XThC.Tn[13].n10 XThC.Tn[13].t12 161.202
R19172 XThC.Tn[13].n13 XThC.Tn[13].t14 161.202
R19173 XThC.Tn[13].n16 XThC.Tn[13].t16 161.202
R19174 XThC.Tn[13].n19 XThC.Tn[13].t37 161.202
R19175 XThC.Tn[13].n22 XThC.Tn[13].t38 161.202
R19176 XThC.Tn[13].n25 XThC.Tn[13].t19 161.202
R19177 XThC.Tn[13].n28 XThC.Tn[13].t28 161.202
R19178 XThC.Tn[13].n31 XThC.Tn[13].t30 161.202
R19179 XThC.Tn[13].n34 XThC.Tn[13].t17 161.202
R19180 XThC.Tn[13].n37 XThC.Tn[13].t18 161.202
R19181 XThC.Tn[13].n40 XThC.Tn[13].t31 161.202
R19182 XThC.Tn[13].n43 XThC.Tn[13].t39 161.202
R19183 XThC.Tn[13].n46 XThC.Tn[13].t42 161.202
R19184 XThC.Tn[13].n49 XThC.Tn[13].t23 161.202
R19185 XThC.Tn[13].n52 XThC.Tn[13].t33 161.202
R19186 XThC.Tn[13].n7 XThC.Tn[13].t29 145.137
R19187 XThC.Tn[13].n10 XThC.Tn[13].t15 145.137
R19188 XThC.Tn[13].n13 XThC.Tn[13].t20 145.137
R19189 XThC.Tn[13].n16 XThC.Tn[13].t21 145.137
R19190 XThC.Tn[13].n19 XThC.Tn[13].t40 145.137
R19191 XThC.Tn[13].n22 XThC.Tn[13].t41 145.137
R19192 XThC.Tn[13].n25 XThC.Tn[13].t25 145.137
R19193 XThC.Tn[13].n28 XThC.Tn[13].t32 145.137
R19194 XThC.Tn[13].n31 XThC.Tn[13].t34 145.137
R19195 XThC.Tn[13].n34 XThC.Tn[13].t22 145.137
R19196 XThC.Tn[13].n37 XThC.Tn[13].t24 145.137
R19197 XThC.Tn[13].n40 XThC.Tn[13].t35 145.137
R19198 XThC.Tn[13].n43 XThC.Tn[13].t43 145.137
R19199 XThC.Tn[13].n46 XThC.Tn[13].t13 145.137
R19200 XThC.Tn[13].n49 XThC.Tn[13].t26 145.137
R19201 XThC.Tn[13].n52 XThC.Tn[13].t36 145.137
R19202 XThC.Tn[13].n1 XThC.Tn[13].t4 26.5955
R19203 XThC.Tn[13].n1 XThC.Tn[13].t7 26.5955
R19204 XThC.Tn[13].n0 XThC.Tn[13].t6 26.5955
R19205 XThC.Tn[13].n0 XThC.Tn[13].t5 26.5955
R19206 XThC.Tn[13].n3 XThC.Tn[13].t9 26.5955
R19207 XThC.Tn[13].n3 XThC.Tn[13].t8 26.5955
R19208 XThC.Tn[13].n4 XThC.Tn[13].t11 26.5955
R19209 XThC.Tn[13].n4 XThC.Tn[13].t10 26.5955
R19210 XThC.Tn[13].n57 XThC.Tn[13].t0 24.9236
R19211 XThC.Tn[13].n57 XThC.Tn[13].t2 24.9236
R19212 XThC.Tn[13].n58 XThC.Tn[13].t3 24.9236
R19213 XThC.Tn[13].n58 XThC.Tn[13].t1 24.9236
R19214 XThC.Tn[13] XThC.Tn[13].n5 22.9652
R19215 XThC.Tn[13] XThC.Tn[13].n59 18.8943
R19216 XThC.Tn[13].n6 XThC.Tn[13].n2 13.9299
R19217 XThC.Tn[13].n6 XThC.Tn[13] 13.9299
R19218 XThC.Tn[13] XThC.Tn[13].n56 6.34069
R19219 XThC.Tn[13].n56 XThC.Tn[13].n55 5.13021
R19220 XThC.Tn[13].n55 XThC.Tn[13] 4.03795
R19221 XThC.Tn[13].n56 XThC.Tn[13] 1.79489
R19222 XThC.Tn[13] XThC.Tn[13].n6 1.19676
R19223 XThC.Tn[13].n12 XThC.Tn[13] 0.931056
R19224 XThC.Tn[13].n15 XThC.Tn[13] 0.931056
R19225 XThC.Tn[13].n18 XThC.Tn[13] 0.931056
R19226 XThC.Tn[13].n21 XThC.Tn[13] 0.931056
R19227 XThC.Tn[13].n24 XThC.Tn[13] 0.931056
R19228 XThC.Tn[13].n27 XThC.Tn[13] 0.931056
R19229 XThC.Tn[13].n30 XThC.Tn[13] 0.931056
R19230 XThC.Tn[13].n33 XThC.Tn[13] 0.931056
R19231 XThC.Tn[13].n36 XThC.Tn[13] 0.931056
R19232 XThC.Tn[13].n39 XThC.Tn[13] 0.931056
R19233 XThC.Tn[13].n42 XThC.Tn[13] 0.931056
R19234 XThC.Tn[13].n45 XThC.Tn[13] 0.931056
R19235 XThC.Tn[13].n48 XThC.Tn[13] 0.931056
R19236 XThC.Tn[13].n51 XThC.Tn[13] 0.931056
R19237 XThC.Tn[13].n54 XThC.Tn[13] 0.931056
R19238 XThC.Tn[13] XThC.Tn[13].n9 0.396333
R19239 XThC.Tn[13] XThC.Tn[13].n12 0.396333
R19240 XThC.Tn[13] XThC.Tn[13].n15 0.396333
R19241 XThC.Tn[13] XThC.Tn[13].n18 0.396333
R19242 XThC.Tn[13] XThC.Tn[13].n21 0.396333
R19243 XThC.Tn[13] XThC.Tn[13].n24 0.396333
R19244 XThC.Tn[13] XThC.Tn[13].n27 0.396333
R19245 XThC.Tn[13] XThC.Tn[13].n30 0.396333
R19246 XThC.Tn[13] XThC.Tn[13].n33 0.396333
R19247 XThC.Tn[13] XThC.Tn[13].n36 0.396333
R19248 XThC.Tn[13] XThC.Tn[13].n39 0.396333
R19249 XThC.Tn[13] XThC.Tn[13].n42 0.396333
R19250 XThC.Tn[13] XThC.Tn[13].n45 0.396333
R19251 XThC.Tn[13] XThC.Tn[13].n48 0.396333
R19252 XThC.Tn[13] XThC.Tn[13].n51 0.396333
R19253 XThC.Tn[13] XThC.Tn[13].n54 0.396333
R19254 XThC.Tn[13].n8 XThC.Tn[13] 0.104667
R19255 XThC.Tn[13].n11 XThC.Tn[13] 0.104667
R19256 XThC.Tn[13].n14 XThC.Tn[13] 0.104667
R19257 XThC.Tn[13].n17 XThC.Tn[13] 0.104667
R19258 XThC.Tn[13].n20 XThC.Tn[13] 0.104667
R19259 XThC.Tn[13].n23 XThC.Tn[13] 0.104667
R19260 XThC.Tn[13].n26 XThC.Tn[13] 0.104667
R19261 XThC.Tn[13].n29 XThC.Tn[13] 0.104667
R19262 XThC.Tn[13].n32 XThC.Tn[13] 0.104667
R19263 XThC.Tn[13].n35 XThC.Tn[13] 0.104667
R19264 XThC.Tn[13].n38 XThC.Tn[13] 0.104667
R19265 XThC.Tn[13].n41 XThC.Tn[13] 0.104667
R19266 XThC.Tn[13].n44 XThC.Tn[13] 0.104667
R19267 XThC.Tn[13].n47 XThC.Tn[13] 0.104667
R19268 XThC.Tn[13].n50 XThC.Tn[13] 0.104667
R19269 XThC.Tn[13].n53 XThC.Tn[13] 0.104667
R19270 XThC.Tn[13].n8 XThC.Tn[13] 0.0309878
R19271 XThC.Tn[13].n11 XThC.Tn[13] 0.0309878
R19272 XThC.Tn[13].n14 XThC.Tn[13] 0.0309878
R19273 XThC.Tn[13].n17 XThC.Tn[13] 0.0309878
R19274 XThC.Tn[13].n20 XThC.Tn[13] 0.0309878
R19275 XThC.Tn[13].n23 XThC.Tn[13] 0.0309878
R19276 XThC.Tn[13].n26 XThC.Tn[13] 0.0309878
R19277 XThC.Tn[13].n29 XThC.Tn[13] 0.0309878
R19278 XThC.Tn[13].n32 XThC.Tn[13] 0.0309878
R19279 XThC.Tn[13].n35 XThC.Tn[13] 0.0309878
R19280 XThC.Tn[13].n38 XThC.Tn[13] 0.0309878
R19281 XThC.Tn[13].n41 XThC.Tn[13] 0.0309878
R19282 XThC.Tn[13].n44 XThC.Tn[13] 0.0309878
R19283 XThC.Tn[13].n47 XThC.Tn[13] 0.0309878
R19284 XThC.Tn[13].n50 XThC.Tn[13] 0.0309878
R19285 XThC.Tn[13].n53 XThC.Tn[13] 0.0309878
R19286 XThC.Tn[13].n9 XThC.Tn[13].n8 0.027939
R19287 XThC.Tn[13].n12 XThC.Tn[13].n11 0.027939
R19288 XThC.Tn[13].n15 XThC.Tn[13].n14 0.027939
R19289 XThC.Tn[13].n18 XThC.Tn[13].n17 0.027939
R19290 XThC.Tn[13].n21 XThC.Tn[13].n20 0.027939
R19291 XThC.Tn[13].n24 XThC.Tn[13].n23 0.027939
R19292 XThC.Tn[13].n27 XThC.Tn[13].n26 0.027939
R19293 XThC.Tn[13].n30 XThC.Tn[13].n29 0.027939
R19294 XThC.Tn[13].n33 XThC.Tn[13].n32 0.027939
R19295 XThC.Tn[13].n36 XThC.Tn[13].n35 0.027939
R19296 XThC.Tn[13].n39 XThC.Tn[13].n38 0.027939
R19297 XThC.Tn[13].n42 XThC.Tn[13].n41 0.027939
R19298 XThC.Tn[13].n45 XThC.Tn[13].n44 0.027939
R19299 XThC.Tn[13].n48 XThC.Tn[13].n47 0.027939
R19300 XThC.Tn[13].n51 XThC.Tn[13].n50 0.027939
R19301 XThC.Tn[13].n54 XThC.Tn[13].n53 0.027939
R19302 XThC.Tn[13].n55 XThC.Tn[13] 0.00548355
R19303 XThC.Tn[0].n2 XThC.Tn[0].n1 332.332
R19304 XThC.Tn[0].n2 XThC.Tn[0].n0 296.493
R19305 XThC.Tn[0].n12 XThC.Tn[0].n10 161.406
R19306 XThC.Tn[0].n15 XThC.Tn[0].n13 161.406
R19307 XThC.Tn[0].n18 XThC.Tn[0].n16 161.406
R19308 XThC.Tn[0].n21 XThC.Tn[0].n19 161.406
R19309 XThC.Tn[0].n24 XThC.Tn[0].n22 161.406
R19310 XThC.Tn[0].n27 XThC.Tn[0].n25 161.406
R19311 XThC.Tn[0].n30 XThC.Tn[0].n28 161.406
R19312 XThC.Tn[0].n33 XThC.Tn[0].n31 161.406
R19313 XThC.Tn[0].n36 XThC.Tn[0].n34 161.406
R19314 XThC.Tn[0].n39 XThC.Tn[0].n37 161.406
R19315 XThC.Tn[0].n42 XThC.Tn[0].n40 161.406
R19316 XThC.Tn[0].n45 XThC.Tn[0].n43 161.406
R19317 XThC.Tn[0].n48 XThC.Tn[0].n46 161.406
R19318 XThC.Tn[0].n51 XThC.Tn[0].n49 161.406
R19319 XThC.Tn[0].n54 XThC.Tn[0].n52 161.406
R19320 XThC.Tn[0].n57 XThC.Tn[0].n55 161.406
R19321 XThC.Tn[0].n10 XThC.Tn[0].t22 161.202
R19322 XThC.Tn[0].n13 XThC.Tn[0].t41 161.202
R19323 XThC.Tn[0].n16 XThC.Tn[0].t12 161.202
R19324 XThC.Tn[0].n19 XThC.Tn[0].t13 161.202
R19325 XThC.Tn[0].n22 XThC.Tn[0].t32 161.202
R19326 XThC.Tn[0].n25 XThC.Tn[0].t34 161.202
R19327 XThC.Tn[0].n28 XThC.Tn[0].t17 161.202
R19328 XThC.Tn[0].n31 XThC.Tn[0].t25 161.202
R19329 XThC.Tn[0].n34 XThC.Tn[0].t26 161.202
R19330 XThC.Tn[0].n37 XThC.Tn[0].t15 161.202
R19331 XThC.Tn[0].n40 XThC.Tn[0].t16 161.202
R19332 XThC.Tn[0].n43 XThC.Tn[0].t27 161.202
R19333 XThC.Tn[0].n46 XThC.Tn[0].t36 161.202
R19334 XThC.Tn[0].n49 XThC.Tn[0].t38 161.202
R19335 XThC.Tn[0].n52 XThC.Tn[0].t19 161.202
R19336 XThC.Tn[0].n55 XThC.Tn[0].t29 161.202
R19337 XThC.Tn[0].n10 XThC.Tn[0].t18 145.137
R19338 XThC.Tn[0].n13 XThC.Tn[0].t35 145.137
R19339 XThC.Tn[0].n16 XThC.Tn[0].t37 145.137
R19340 XThC.Tn[0].n19 XThC.Tn[0].t39 145.137
R19341 XThC.Tn[0].n22 XThC.Tn[0].t28 145.137
R19342 XThC.Tn[0].n25 XThC.Tn[0].t30 145.137
R19343 XThC.Tn[0].n28 XThC.Tn[0].t43 145.137
R19344 XThC.Tn[0].n31 XThC.Tn[0].t20 145.137
R19345 XThC.Tn[0].n34 XThC.Tn[0].t21 145.137
R19346 XThC.Tn[0].n37 XThC.Tn[0].t40 145.137
R19347 XThC.Tn[0].n40 XThC.Tn[0].t42 145.137
R19348 XThC.Tn[0].n43 XThC.Tn[0].t23 145.137
R19349 XThC.Tn[0].n46 XThC.Tn[0].t31 145.137
R19350 XThC.Tn[0].n49 XThC.Tn[0].t33 145.137
R19351 XThC.Tn[0].n52 XThC.Tn[0].t14 145.137
R19352 XThC.Tn[0].n55 XThC.Tn[0].t24 145.137
R19353 XThC.Tn[0].n7 XThC.Tn[0].n6 135.248
R19354 XThC.Tn[0].n9 XThC.Tn[0].n3 98.982
R19355 XThC.Tn[0].n8 XThC.Tn[0].n4 98.982
R19356 XThC.Tn[0].n7 XThC.Tn[0].n5 98.982
R19357 XThC.Tn[0].n9 XThC.Tn[0].n8 36.2672
R19358 XThC.Tn[0].n8 XThC.Tn[0].n7 36.2672
R19359 XThC.Tn[0].n59 XThC.Tn[0].n9 32.6405
R19360 XThC.Tn[0].n1 XThC.Tn[0].t6 26.5955
R19361 XThC.Tn[0].n1 XThC.Tn[0].t5 26.5955
R19362 XThC.Tn[0].n0 XThC.Tn[0].t4 26.5955
R19363 XThC.Tn[0].n0 XThC.Tn[0].t3 26.5955
R19364 XThC.Tn[0].n3 XThC.Tn[0].t8 24.9236
R19365 XThC.Tn[0].n3 XThC.Tn[0].t7 24.9236
R19366 XThC.Tn[0].n4 XThC.Tn[0].t10 24.9236
R19367 XThC.Tn[0].n4 XThC.Tn[0].t9 24.9236
R19368 XThC.Tn[0].n5 XThC.Tn[0].t1 24.9236
R19369 XThC.Tn[0].n5 XThC.Tn[0].t2 24.9236
R19370 XThC.Tn[0].n6 XThC.Tn[0].t11 24.9236
R19371 XThC.Tn[0].n6 XThC.Tn[0].t0 24.9236
R19372 XThC.Tn[0].n60 XThC.Tn[0].n2 18.5605
R19373 XThC.Tn[0].n60 XThC.Tn[0].n59 11.5205
R19374 XThC.Tn[0].n59 XThC.Tn[0].n58 3.16389
R19375 XThC.Tn[0].n15 XThC.Tn[0] 0.931056
R19376 XThC.Tn[0].n18 XThC.Tn[0] 0.931056
R19377 XThC.Tn[0].n21 XThC.Tn[0] 0.931056
R19378 XThC.Tn[0].n24 XThC.Tn[0] 0.931056
R19379 XThC.Tn[0].n27 XThC.Tn[0] 0.931056
R19380 XThC.Tn[0].n30 XThC.Tn[0] 0.931056
R19381 XThC.Tn[0].n33 XThC.Tn[0] 0.931056
R19382 XThC.Tn[0].n36 XThC.Tn[0] 0.931056
R19383 XThC.Tn[0].n39 XThC.Tn[0] 0.931056
R19384 XThC.Tn[0].n42 XThC.Tn[0] 0.931056
R19385 XThC.Tn[0].n45 XThC.Tn[0] 0.931056
R19386 XThC.Tn[0].n48 XThC.Tn[0] 0.931056
R19387 XThC.Tn[0].n51 XThC.Tn[0] 0.931056
R19388 XThC.Tn[0].n54 XThC.Tn[0] 0.931056
R19389 XThC.Tn[0].n57 XThC.Tn[0] 0.931056
R19390 XThC.Tn[0] XThC.Tn[0].n60 0.6405
R19391 XThC.Tn[0] XThC.Tn[0].n12 0.396333
R19392 XThC.Tn[0] XThC.Tn[0].n15 0.396333
R19393 XThC.Tn[0] XThC.Tn[0].n18 0.396333
R19394 XThC.Tn[0] XThC.Tn[0].n21 0.396333
R19395 XThC.Tn[0] XThC.Tn[0].n24 0.396333
R19396 XThC.Tn[0] XThC.Tn[0].n27 0.396333
R19397 XThC.Tn[0] XThC.Tn[0].n30 0.396333
R19398 XThC.Tn[0] XThC.Tn[0].n33 0.396333
R19399 XThC.Tn[0] XThC.Tn[0].n36 0.396333
R19400 XThC.Tn[0] XThC.Tn[0].n39 0.396333
R19401 XThC.Tn[0] XThC.Tn[0].n42 0.396333
R19402 XThC.Tn[0] XThC.Tn[0].n45 0.396333
R19403 XThC.Tn[0] XThC.Tn[0].n48 0.396333
R19404 XThC.Tn[0] XThC.Tn[0].n51 0.396333
R19405 XThC.Tn[0] XThC.Tn[0].n54 0.396333
R19406 XThC.Tn[0] XThC.Tn[0].n57 0.396333
R19407 XThC.Tn[0].n58 XThC.Tn[0] 0.243556
R19408 XThC.Tn[0].n11 XThC.Tn[0] 0.104667
R19409 XThC.Tn[0].n14 XThC.Tn[0] 0.104667
R19410 XThC.Tn[0].n17 XThC.Tn[0] 0.104667
R19411 XThC.Tn[0].n20 XThC.Tn[0] 0.104667
R19412 XThC.Tn[0].n23 XThC.Tn[0] 0.104667
R19413 XThC.Tn[0].n26 XThC.Tn[0] 0.104667
R19414 XThC.Tn[0].n29 XThC.Tn[0] 0.104667
R19415 XThC.Tn[0].n32 XThC.Tn[0] 0.104667
R19416 XThC.Tn[0].n35 XThC.Tn[0] 0.104667
R19417 XThC.Tn[0].n38 XThC.Tn[0] 0.104667
R19418 XThC.Tn[0].n41 XThC.Tn[0] 0.104667
R19419 XThC.Tn[0].n44 XThC.Tn[0] 0.104667
R19420 XThC.Tn[0].n47 XThC.Tn[0] 0.104667
R19421 XThC.Tn[0].n50 XThC.Tn[0] 0.104667
R19422 XThC.Tn[0].n53 XThC.Tn[0] 0.104667
R19423 XThC.Tn[0].n56 XThC.Tn[0] 0.104667
R19424 XThC.Tn[0].n58 XThC.Tn[0] 0.0326429
R19425 XThC.Tn[0].n11 XThC.Tn[0] 0.0309878
R19426 XThC.Tn[0].n14 XThC.Tn[0] 0.0309878
R19427 XThC.Tn[0].n17 XThC.Tn[0] 0.0309878
R19428 XThC.Tn[0].n20 XThC.Tn[0] 0.0309878
R19429 XThC.Tn[0].n23 XThC.Tn[0] 0.0309878
R19430 XThC.Tn[0].n26 XThC.Tn[0] 0.0309878
R19431 XThC.Tn[0].n29 XThC.Tn[0] 0.0309878
R19432 XThC.Tn[0].n32 XThC.Tn[0] 0.0309878
R19433 XThC.Tn[0].n35 XThC.Tn[0] 0.0309878
R19434 XThC.Tn[0].n38 XThC.Tn[0] 0.0309878
R19435 XThC.Tn[0].n41 XThC.Tn[0] 0.0309878
R19436 XThC.Tn[0].n44 XThC.Tn[0] 0.0309878
R19437 XThC.Tn[0].n47 XThC.Tn[0] 0.0309878
R19438 XThC.Tn[0].n50 XThC.Tn[0] 0.0309878
R19439 XThC.Tn[0].n53 XThC.Tn[0] 0.0309878
R19440 XThC.Tn[0].n56 XThC.Tn[0] 0.0309878
R19441 XThC.Tn[0].n12 XThC.Tn[0].n11 0.027939
R19442 XThC.Tn[0].n15 XThC.Tn[0].n14 0.027939
R19443 XThC.Tn[0].n18 XThC.Tn[0].n17 0.027939
R19444 XThC.Tn[0].n21 XThC.Tn[0].n20 0.027939
R19445 XThC.Tn[0].n24 XThC.Tn[0].n23 0.027939
R19446 XThC.Tn[0].n27 XThC.Tn[0].n26 0.027939
R19447 XThC.Tn[0].n30 XThC.Tn[0].n29 0.027939
R19448 XThC.Tn[0].n33 XThC.Tn[0].n32 0.027939
R19449 XThC.Tn[0].n36 XThC.Tn[0].n35 0.027939
R19450 XThC.Tn[0].n39 XThC.Tn[0].n38 0.027939
R19451 XThC.Tn[0].n42 XThC.Tn[0].n41 0.027939
R19452 XThC.Tn[0].n45 XThC.Tn[0].n44 0.027939
R19453 XThC.Tn[0].n48 XThC.Tn[0].n47 0.027939
R19454 XThC.Tn[0].n51 XThC.Tn[0].n50 0.027939
R19455 XThC.Tn[0].n54 XThC.Tn[0].n53 0.027939
R19456 XThC.Tn[0].n57 XThC.Tn[0].n56 0.027939
R19457 XThC.XTB4.Y.t0 XThC.XTB4.Y.n21 268.738
R19458 XThC.XTB4.Y.n22 XThC.XTB4.Y.t0 268.077
R19459 XThC.XTB4.Y.n0 XThC.XTB4.Y.t1 235.56
R19460 XThC.XTB4.Y.n4 XThC.XTB4.Y.t3 212.081
R19461 XThC.XTB4.Y.n3 XThC.XTB4.Y.t2 212.081
R19462 XThC.XTB4.Y.n9 XThC.XTB4.Y.t17 212.081
R19463 XThC.XTB4.Y.n1 XThC.XTB4.Y.t13 212.081
R19464 XThC.XTB4.Y.n13 XThC.XTB4.Y.t8 212.081
R19465 XThC.XTB4.Y.n14 XThC.XTB4.Y.t12 212.081
R19466 XThC.XTB4.Y.n16 XThC.XTB4.Y.t6 212.081
R19467 XThC.XTB4.Y.n12 XThC.XTB4.Y.t16 212.081
R19468 XThC.XTB4.Y.n6 XThC.XTB4.Y.n5 173.761
R19469 XThC.XTB4.Y.n15 XThC.XTB4.Y 158.656
R19470 XThC.XTB4.Y.n8 XThC.XTB4.Y.n7 152
R19471 XThC.XTB4.Y.n6 XThC.XTB4.Y.n2 152
R19472 XThC.XTB4.Y.n11 XThC.XTB4.Y.n10 152
R19473 XThC.XTB4.Y.n18 XThC.XTB4.Y.n17 152
R19474 XThC.XTB4.Y.n4 XThC.XTB4.Y.t14 139.78
R19475 XThC.XTB4.Y.n3 XThC.XTB4.Y.t10 139.78
R19476 XThC.XTB4.Y.n9 XThC.XTB4.Y.t7 139.78
R19477 XThC.XTB4.Y.n1 XThC.XTB4.Y.t4 139.78
R19478 XThC.XTB4.Y.n13 XThC.XTB4.Y.t11 139.78
R19479 XThC.XTB4.Y.n14 XThC.XTB4.Y.t15 139.78
R19480 XThC.XTB4.Y.n16 XThC.XTB4.Y.t9 139.78
R19481 XThC.XTB4.Y.n12 XThC.XTB4.Y.t5 139.78
R19482 XThC.XTB4.Y.n20 XThC.XTB4.Y.n11 72.9296
R19483 XThC.XTB4.Y.n14 XThC.XTB4.Y.n13 61.346
R19484 XThC.XTB4.Y.n8 XThC.XTB4.Y.n2 49.6611
R19485 XThC.XTB4.Y.n10 XThC.XTB4.Y.n9 45.2793
R19486 XThC.XTB4.Y.n5 XThC.XTB4.Y.n3 42.3581
R19487 XThC.XTB4.Y.n20 XThC.XTB4.Y.n19 38.1854
R19488 XThC.XTB4.Y.n17 XThC.XTB4.Y.n12 30.6732
R19489 XThC.XTB4.Y.n17 XThC.XTB4.Y.n16 30.6732
R19490 XThC.XTB4.Y.n16 XThC.XTB4.Y.n15 30.6732
R19491 XThC.XTB4.Y.n15 XThC.XTB4.Y.n14 30.6732
R19492 XThC.XTB4.Y.n7 XThC.XTB4.Y.n6 21.7605
R19493 XThC.XTB4.Y.n5 XThC.XTB4.Y.n4 18.9884
R19494 XThC.XTB4.Y XThC.XTB4.Y.n22 17.8682
R19495 XThC.XTB4.Y.n10 XThC.XTB4.Y.n1 16.0672
R19496 XThC.XTB4.Y.n18 XThC.XTB4.Y 14.7905
R19497 XThC.XTB4.Y.n11 XThC.XTB4.Y 11.5205
R19498 XThC.XTB4.Y.n21 XThC.XTB4.Y.n20 10.353
R19499 XThC.XTB4.Y.n7 XThC.XTB4.Y 10.2405
R19500 XThC.XTB4.Y.n3 XThC.XTB4.Y.n2 7.30353
R19501 XThC.XTB4.Y.n19 XThC.XTB4.Y.n18 7.24578
R19502 XThC.XTB4.Y.n9 XThC.XTB4.Y.n8 4.38232
R19503 XThC.XTB4.Y.n22 XThC.XTB4.Y.n21 3.29747
R19504 XThC.XTB4.Y XThC.XTB4.Y.n0 2.22659
R19505 XThC.XTB4.Y.n0 XThC.XTB4.Y 1.55202
R19506 XThC.XTB4.Y.n19 XThC.XTB4.Y 0.966538
R19507 XThR.Tn[3].n2 XThR.Tn[3].n1 332.332
R19508 XThR.Tn[3].n2 XThR.Tn[3].n0 296.493
R19509 XThR.Tn[3] XThR.Tn[3].n82 161.363
R19510 XThR.Tn[3] XThR.Tn[3].n77 161.363
R19511 XThR.Tn[3] XThR.Tn[3].n72 161.363
R19512 XThR.Tn[3] XThR.Tn[3].n67 161.363
R19513 XThR.Tn[3] XThR.Tn[3].n62 161.363
R19514 XThR.Tn[3] XThR.Tn[3].n57 161.363
R19515 XThR.Tn[3] XThR.Tn[3].n52 161.363
R19516 XThR.Tn[3] XThR.Tn[3].n47 161.363
R19517 XThR.Tn[3] XThR.Tn[3].n42 161.363
R19518 XThR.Tn[3] XThR.Tn[3].n37 161.363
R19519 XThR.Tn[3] XThR.Tn[3].n32 161.363
R19520 XThR.Tn[3] XThR.Tn[3].n27 161.363
R19521 XThR.Tn[3] XThR.Tn[3].n22 161.363
R19522 XThR.Tn[3] XThR.Tn[3].n17 161.363
R19523 XThR.Tn[3] XThR.Tn[3].n12 161.363
R19524 XThR.Tn[3] XThR.Tn[3].n10 161.363
R19525 XThR.Tn[3].n84 XThR.Tn[3].n83 161.3
R19526 XThR.Tn[3].n79 XThR.Tn[3].n78 161.3
R19527 XThR.Tn[3].n74 XThR.Tn[3].n73 161.3
R19528 XThR.Tn[3].n69 XThR.Tn[3].n68 161.3
R19529 XThR.Tn[3].n64 XThR.Tn[3].n63 161.3
R19530 XThR.Tn[3].n59 XThR.Tn[3].n58 161.3
R19531 XThR.Tn[3].n54 XThR.Tn[3].n53 161.3
R19532 XThR.Tn[3].n49 XThR.Tn[3].n48 161.3
R19533 XThR.Tn[3].n44 XThR.Tn[3].n43 161.3
R19534 XThR.Tn[3].n39 XThR.Tn[3].n38 161.3
R19535 XThR.Tn[3].n34 XThR.Tn[3].n33 161.3
R19536 XThR.Tn[3].n29 XThR.Tn[3].n28 161.3
R19537 XThR.Tn[3].n24 XThR.Tn[3].n23 161.3
R19538 XThR.Tn[3].n19 XThR.Tn[3].n18 161.3
R19539 XThR.Tn[3].n14 XThR.Tn[3].n13 161.3
R19540 XThR.Tn[3].n82 XThR.Tn[3].t46 161.106
R19541 XThR.Tn[3].n77 XThR.Tn[3].t53 161.106
R19542 XThR.Tn[3].n72 XThR.Tn[3].t34 161.106
R19543 XThR.Tn[3].n67 XThR.Tn[3].t17 161.106
R19544 XThR.Tn[3].n62 XThR.Tn[3].t44 161.106
R19545 XThR.Tn[3].n57 XThR.Tn[3].t69 161.106
R19546 XThR.Tn[3].n52 XThR.Tn[3].t51 161.106
R19547 XThR.Tn[3].n47 XThR.Tn[3].t31 161.106
R19548 XThR.Tn[3].n42 XThR.Tn[3].t14 161.106
R19549 XThR.Tn[3].n37 XThR.Tn[3].t20 161.106
R19550 XThR.Tn[3].n32 XThR.Tn[3].t68 161.106
R19551 XThR.Tn[3].n27 XThR.Tn[3].t33 161.106
R19552 XThR.Tn[3].n22 XThR.Tn[3].t67 161.106
R19553 XThR.Tn[3].n17 XThR.Tn[3].t49 161.106
R19554 XThR.Tn[3].n12 XThR.Tn[3].t70 161.106
R19555 XThR.Tn[3].n10 XThR.Tn[3].t57 161.106
R19556 XThR.Tn[3].n83 XThR.Tn[3].t27 159.978
R19557 XThR.Tn[3].n78 XThR.Tn[3].t32 159.978
R19558 XThR.Tn[3].n73 XThR.Tn[3].t15 159.978
R19559 XThR.Tn[3].n68 XThR.Tn[3].t63 159.978
R19560 XThR.Tn[3].n63 XThR.Tn[3].t25 159.978
R19561 XThR.Tn[3].n58 XThR.Tn[3].t50 159.978
R19562 XThR.Tn[3].n53 XThR.Tn[3].t30 159.978
R19563 XThR.Tn[3].n48 XThR.Tn[3].t73 159.978
R19564 XThR.Tn[3].n43 XThR.Tn[3].t61 159.978
R19565 XThR.Tn[3].n38 XThR.Tn[3].t66 159.978
R19566 XThR.Tn[3].n33 XThR.Tn[3].t48 159.978
R19567 XThR.Tn[3].n28 XThR.Tn[3].t13 159.978
R19568 XThR.Tn[3].n23 XThR.Tn[3].t47 159.978
R19569 XThR.Tn[3].n18 XThR.Tn[3].t29 159.978
R19570 XThR.Tn[3].n13 XThR.Tn[3].t55 159.978
R19571 XThR.Tn[3].n82 XThR.Tn[3].t36 145.038
R19572 XThR.Tn[3].n77 XThR.Tn[3].t60 145.038
R19573 XThR.Tn[3].n72 XThR.Tn[3].t40 145.038
R19574 XThR.Tn[3].n67 XThR.Tn[3].t21 145.038
R19575 XThR.Tn[3].n62 XThR.Tn[3].t54 145.038
R19576 XThR.Tn[3].n57 XThR.Tn[3].t35 145.038
R19577 XThR.Tn[3].n52 XThR.Tn[3].t41 145.038
R19578 XThR.Tn[3].n47 XThR.Tn[3].t22 145.038
R19579 XThR.Tn[3].n42 XThR.Tn[3].t19 145.038
R19580 XThR.Tn[3].n37 XThR.Tn[3].t52 145.038
R19581 XThR.Tn[3].n32 XThR.Tn[3].t72 145.038
R19582 XThR.Tn[3].n27 XThR.Tn[3].t39 145.038
R19583 XThR.Tn[3].n22 XThR.Tn[3].t71 145.038
R19584 XThR.Tn[3].n17 XThR.Tn[3].t59 145.038
R19585 XThR.Tn[3].n12 XThR.Tn[3].t18 145.038
R19586 XThR.Tn[3].n10 XThR.Tn[3].t64 145.038
R19587 XThR.Tn[3].n83 XThR.Tn[3].t38 143.911
R19588 XThR.Tn[3].n78 XThR.Tn[3].t65 143.911
R19589 XThR.Tn[3].n73 XThR.Tn[3].t43 143.911
R19590 XThR.Tn[3].n68 XThR.Tn[3].t26 143.911
R19591 XThR.Tn[3].n63 XThR.Tn[3].t58 143.911
R19592 XThR.Tn[3].n58 XThR.Tn[3].t37 143.911
R19593 XThR.Tn[3].n53 XThR.Tn[3].t45 143.911
R19594 XThR.Tn[3].n48 XThR.Tn[3].t28 143.911
R19595 XThR.Tn[3].n43 XThR.Tn[3].t23 143.911
R19596 XThR.Tn[3].n38 XThR.Tn[3].t56 143.911
R19597 XThR.Tn[3].n33 XThR.Tn[3].t16 143.911
R19598 XThR.Tn[3].n28 XThR.Tn[3].t42 143.911
R19599 XThR.Tn[3].n23 XThR.Tn[3].t12 143.911
R19600 XThR.Tn[3].n18 XThR.Tn[3].t62 143.911
R19601 XThR.Tn[3].n13 XThR.Tn[3].t24 143.911
R19602 XThR.Tn[3].n7 XThR.Tn[3].n5 135.249
R19603 XThR.Tn[3].n9 XThR.Tn[3].n3 98.981
R19604 XThR.Tn[3].n8 XThR.Tn[3].n4 98.981
R19605 XThR.Tn[3].n7 XThR.Tn[3].n6 98.981
R19606 XThR.Tn[3].n9 XThR.Tn[3].n8 36.2672
R19607 XThR.Tn[3].n8 XThR.Tn[3].n7 36.2672
R19608 XThR.Tn[3].n88 XThR.Tn[3].n9 32.6405
R19609 XThR.Tn[3].n1 XThR.Tn[3].t8 26.5955
R19610 XThR.Tn[3].n1 XThR.Tn[3].t11 26.5955
R19611 XThR.Tn[3].n0 XThR.Tn[3].t9 26.5955
R19612 XThR.Tn[3].n0 XThR.Tn[3].t10 26.5955
R19613 XThR.Tn[3].n3 XThR.Tn[3].t7 24.9236
R19614 XThR.Tn[3].n3 XThR.Tn[3].t4 24.9236
R19615 XThR.Tn[3].n4 XThR.Tn[3].t6 24.9236
R19616 XThR.Tn[3].n4 XThR.Tn[3].t5 24.9236
R19617 XThR.Tn[3].n5 XThR.Tn[3].t0 24.9236
R19618 XThR.Tn[3].n5 XThR.Tn[3].t1 24.9236
R19619 XThR.Tn[3].n6 XThR.Tn[3].t3 24.9236
R19620 XThR.Tn[3].n6 XThR.Tn[3].t2 24.9236
R19621 XThR.Tn[3].n89 XThR.Tn[3].n2 18.5605
R19622 XThR.Tn[3].n89 XThR.Tn[3].n88 11.5205
R19623 XThR.Tn[3].n88 XThR.Tn[3] 6.21508
R19624 XThR.Tn[3] XThR.Tn[3].n11 5.34038
R19625 XThR.Tn[3].n16 XThR.Tn[3].n15 4.5005
R19626 XThR.Tn[3].n21 XThR.Tn[3].n20 4.5005
R19627 XThR.Tn[3].n26 XThR.Tn[3].n25 4.5005
R19628 XThR.Tn[3].n31 XThR.Tn[3].n30 4.5005
R19629 XThR.Tn[3].n36 XThR.Tn[3].n35 4.5005
R19630 XThR.Tn[3].n41 XThR.Tn[3].n40 4.5005
R19631 XThR.Tn[3].n46 XThR.Tn[3].n45 4.5005
R19632 XThR.Tn[3].n51 XThR.Tn[3].n50 4.5005
R19633 XThR.Tn[3].n56 XThR.Tn[3].n55 4.5005
R19634 XThR.Tn[3].n61 XThR.Tn[3].n60 4.5005
R19635 XThR.Tn[3].n66 XThR.Tn[3].n65 4.5005
R19636 XThR.Tn[3].n71 XThR.Tn[3].n70 4.5005
R19637 XThR.Tn[3].n76 XThR.Tn[3].n75 4.5005
R19638 XThR.Tn[3].n81 XThR.Tn[3].n80 4.5005
R19639 XThR.Tn[3].n86 XThR.Tn[3].n85 4.5005
R19640 XThR.Tn[3].n87 XThR.Tn[3] 3.70586
R19641 XThR.Tn[3].n16 XThR.Tn[3] 2.52282
R19642 XThR.Tn[3].n21 XThR.Tn[3] 2.52282
R19643 XThR.Tn[3].n26 XThR.Tn[3] 2.52282
R19644 XThR.Tn[3].n31 XThR.Tn[3] 2.52282
R19645 XThR.Tn[3].n36 XThR.Tn[3] 2.52282
R19646 XThR.Tn[3].n41 XThR.Tn[3] 2.52282
R19647 XThR.Tn[3].n46 XThR.Tn[3] 2.52282
R19648 XThR.Tn[3].n51 XThR.Tn[3] 2.52282
R19649 XThR.Tn[3].n56 XThR.Tn[3] 2.52282
R19650 XThR.Tn[3].n61 XThR.Tn[3] 2.52282
R19651 XThR.Tn[3].n66 XThR.Tn[3] 2.52282
R19652 XThR.Tn[3].n71 XThR.Tn[3] 2.52282
R19653 XThR.Tn[3].n76 XThR.Tn[3] 2.52282
R19654 XThR.Tn[3].n81 XThR.Tn[3] 2.52282
R19655 XThR.Tn[3].n86 XThR.Tn[3] 2.52282
R19656 XThR.Tn[3].n84 XThR.Tn[3] 1.08677
R19657 XThR.Tn[3].n79 XThR.Tn[3] 1.08677
R19658 XThR.Tn[3].n74 XThR.Tn[3] 1.08677
R19659 XThR.Tn[3].n69 XThR.Tn[3] 1.08677
R19660 XThR.Tn[3].n64 XThR.Tn[3] 1.08677
R19661 XThR.Tn[3].n59 XThR.Tn[3] 1.08677
R19662 XThR.Tn[3].n54 XThR.Tn[3] 1.08677
R19663 XThR.Tn[3].n49 XThR.Tn[3] 1.08677
R19664 XThR.Tn[3].n44 XThR.Tn[3] 1.08677
R19665 XThR.Tn[3].n39 XThR.Tn[3] 1.08677
R19666 XThR.Tn[3].n34 XThR.Tn[3] 1.08677
R19667 XThR.Tn[3].n29 XThR.Tn[3] 1.08677
R19668 XThR.Tn[3].n24 XThR.Tn[3] 1.08677
R19669 XThR.Tn[3].n19 XThR.Tn[3] 1.08677
R19670 XThR.Tn[3].n14 XThR.Tn[3] 1.08677
R19671 XThR.Tn[3] XThR.Tn[3].n16 0.839786
R19672 XThR.Tn[3] XThR.Tn[3].n21 0.839786
R19673 XThR.Tn[3] XThR.Tn[3].n26 0.839786
R19674 XThR.Tn[3] XThR.Tn[3].n31 0.839786
R19675 XThR.Tn[3] XThR.Tn[3].n36 0.839786
R19676 XThR.Tn[3] XThR.Tn[3].n41 0.839786
R19677 XThR.Tn[3] XThR.Tn[3].n46 0.839786
R19678 XThR.Tn[3] XThR.Tn[3].n51 0.839786
R19679 XThR.Tn[3] XThR.Tn[3].n56 0.839786
R19680 XThR.Tn[3] XThR.Tn[3].n61 0.839786
R19681 XThR.Tn[3] XThR.Tn[3].n66 0.839786
R19682 XThR.Tn[3] XThR.Tn[3].n71 0.839786
R19683 XThR.Tn[3] XThR.Tn[3].n76 0.839786
R19684 XThR.Tn[3] XThR.Tn[3].n81 0.839786
R19685 XThR.Tn[3] XThR.Tn[3].n86 0.839786
R19686 XThR.Tn[3] XThR.Tn[3].n89 0.6405
R19687 XThR.Tn[3].n11 XThR.Tn[3] 0.499542
R19688 XThR.Tn[3].n85 XThR.Tn[3] 0.063
R19689 XThR.Tn[3].n80 XThR.Tn[3] 0.063
R19690 XThR.Tn[3].n75 XThR.Tn[3] 0.063
R19691 XThR.Tn[3].n70 XThR.Tn[3] 0.063
R19692 XThR.Tn[3].n65 XThR.Tn[3] 0.063
R19693 XThR.Tn[3].n60 XThR.Tn[3] 0.063
R19694 XThR.Tn[3].n55 XThR.Tn[3] 0.063
R19695 XThR.Tn[3].n50 XThR.Tn[3] 0.063
R19696 XThR.Tn[3].n45 XThR.Tn[3] 0.063
R19697 XThR.Tn[3].n40 XThR.Tn[3] 0.063
R19698 XThR.Tn[3].n35 XThR.Tn[3] 0.063
R19699 XThR.Tn[3].n30 XThR.Tn[3] 0.063
R19700 XThR.Tn[3].n25 XThR.Tn[3] 0.063
R19701 XThR.Tn[3].n20 XThR.Tn[3] 0.063
R19702 XThR.Tn[3].n15 XThR.Tn[3] 0.063
R19703 XThR.Tn[3].n87 XThR.Tn[3] 0.0540714
R19704 XThR.Tn[3] XThR.Tn[3].n87 0.038
R19705 XThR.Tn[3].n11 XThR.Tn[3] 0.0143889
R19706 XThR.Tn[3].n85 XThR.Tn[3].n84 0.00771154
R19707 XThR.Tn[3].n80 XThR.Tn[3].n79 0.00771154
R19708 XThR.Tn[3].n75 XThR.Tn[3].n74 0.00771154
R19709 XThR.Tn[3].n70 XThR.Tn[3].n69 0.00771154
R19710 XThR.Tn[3].n65 XThR.Tn[3].n64 0.00771154
R19711 XThR.Tn[3].n60 XThR.Tn[3].n59 0.00771154
R19712 XThR.Tn[3].n55 XThR.Tn[3].n54 0.00771154
R19713 XThR.Tn[3].n50 XThR.Tn[3].n49 0.00771154
R19714 XThR.Tn[3].n45 XThR.Tn[3].n44 0.00771154
R19715 XThR.Tn[3].n40 XThR.Tn[3].n39 0.00771154
R19716 XThR.Tn[3].n35 XThR.Tn[3].n34 0.00771154
R19717 XThR.Tn[3].n30 XThR.Tn[3].n29 0.00771154
R19718 XThR.Tn[3].n25 XThR.Tn[3].n24 0.00771154
R19719 XThR.Tn[3].n20 XThR.Tn[3].n19 0.00771154
R19720 XThR.Tn[3].n15 XThR.Tn[3].n14 0.00771154
R19721 XThR.Tn[5].n2 XThR.Tn[5].n1 332.332
R19722 XThR.Tn[5].n2 XThR.Tn[5].n0 296.493
R19723 XThR.Tn[5] XThR.Tn[5].n82 161.363
R19724 XThR.Tn[5] XThR.Tn[5].n77 161.363
R19725 XThR.Tn[5] XThR.Tn[5].n72 161.363
R19726 XThR.Tn[5] XThR.Tn[5].n67 161.363
R19727 XThR.Tn[5] XThR.Tn[5].n62 161.363
R19728 XThR.Tn[5] XThR.Tn[5].n57 161.363
R19729 XThR.Tn[5] XThR.Tn[5].n52 161.363
R19730 XThR.Tn[5] XThR.Tn[5].n47 161.363
R19731 XThR.Tn[5] XThR.Tn[5].n42 161.363
R19732 XThR.Tn[5] XThR.Tn[5].n37 161.363
R19733 XThR.Tn[5] XThR.Tn[5].n32 161.363
R19734 XThR.Tn[5] XThR.Tn[5].n27 161.363
R19735 XThR.Tn[5] XThR.Tn[5].n22 161.363
R19736 XThR.Tn[5] XThR.Tn[5].n17 161.363
R19737 XThR.Tn[5] XThR.Tn[5].n12 161.363
R19738 XThR.Tn[5] XThR.Tn[5].n10 161.363
R19739 XThR.Tn[5].n84 XThR.Tn[5].n83 161.3
R19740 XThR.Tn[5].n79 XThR.Tn[5].n78 161.3
R19741 XThR.Tn[5].n74 XThR.Tn[5].n73 161.3
R19742 XThR.Tn[5].n69 XThR.Tn[5].n68 161.3
R19743 XThR.Tn[5].n64 XThR.Tn[5].n63 161.3
R19744 XThR.Tn[5].n59 XThR.Tn[5].n58 161.3
R19745 XThR.Tn[5].n54 XThR.Tn[5].n53 161.3
R19746 XThR.Tn[5].n49 XThR.Tn[5].n48 161.3
R19747 XThR.Tn[5].n44 XThR.Tn[5].n43 161.3
R19748 XThR.Tn[5].n39 XThR.Tn[5].n38 161.3
R19749 XThR.Tn[5].n34 XThR.Tn[5].n33 161.3
R19750 XThR.Tn[5].n29 XThR.Tn[5].n28 161.3
R19751 XThR.Tn[5].n24 XThR.Tn[5].n23 161.3
R19752 XThR.Tn[5].n19 XThR.Tn[5].n18 161.3
R19753 XThR.Tn[5].n14 XThR.Tn[5].n13 161.3
R19754 XThR.Tn[5].n82 XThR.Tn[5].t62 161.106
R19755 XThR.Tn[5].n77 XThR.Tn[5].t70 161.106
R19756 XThR.Tn[5].n72 XThR.Tn[5].t52 161.106
R19757 XThR.Tn[5].n67 XThR.Tn[5].t35 161.106
R19758 XThR.Tn[5].n62 XThR.Tn[5].t60 161.106
R19759 XThR.Tn[5].n57 XThR.Tn[5].t24 161.106
R19760 XThR.Tn[5].n52 XThR.Tn[5].t68 161.106
R19761 XThR.Tn[5].n47 XThR.Tn[5].t49 161.106
R19762 XThR.Tn[5].n42 XThR.Tn[5].t32 161.106
R19763 XThR.Tn[5].n37 XThR.Tn[5].t40 161.106
R19764 XThR.Tn[5].n32 XThR.Tn[5].t22 161.106
R19765 XThR.Tn[5].n27 XThR.Tn[5].t51 161.106
R19766 XThR.Tn[5].n22 XThR.Tn[5].t21 161.106
R19767 XThR.Tn[5].n17 XThR.Tn[5].t66 161.106
R19768 XThR.Tn[5].n12 XThR.Tn[5].t26 161.106
R19769 XThR.Tn[5].n10 XThR.Tn[5].t72 161.106
R19770 XThR.Tn[5].n83 XThR.Tn[5].t59 159.978
R19771 XThR.Tn[5].n78 XThR.Tn[5].t64 159.978
R19772 XThR.Tn[5].n73 XThR.Tn[5].t47 159.978
R19773 XThR.Tn[5].n68 XThR.Tn[5].t31 159.978
R19774 XThR.Tn[5].n63 XThR.Tn[5].t57 159.978
R19775 XThR.Tn[5].n58 XThR.Tn[5].t20 159.978
R19776 XThR.Tn[5].n53 XThR.Tn[5].t63 159.978
R19777 XThR.Tn[5].n48 XThR.Tn[5].t45 159.978
R19778 XThR.Tn[5].n43 XThR.Tn[5].t29 159.978
R19779 XThR.Tn[5].n38 XThR.Tn[5].t37 159.978
R19780 XThR.Tn[5].n33 XThR.Tn[5].t19 159.978
R19781 XThR.Tn[5].n28 XThR.Tn[5].t46 159.978
R19782 XThR.Tn[5].n23 XThR.Tn[5].t18 159.978
R19783 XThR.Tn[5].n18 XThR.Tn[5].t61 159.978
R19784 XThR.Tn[5].n13 XThR.Tn[5].t23 159.978
R19785 XThR.Tn[5].n82 XThR.Tn[5].t54 145.038
R19786 XThR.Tn[5].n77 XThR.Tn[5].t12 145.038
R19787 XThR.Tn[5].n72 XThR.Tn[5].t56 145.038
R19788 XThR.Tn[5].n67 XThR.Tn[5].t41 145.038
R19789 XThR.Tn[5].n62 XThR.Tn[5].t71 145.038
R19790 XThR.Tn[5].n57 XThR.Tn[5].t53 145.038
R19791 XThR.Tn[5].n52 XThR.Tn[5].t58 145.038
R19792 XThR.Tn[5].n47 XThR.Tn[5].t42 145.038
R19793 XThR.Tn[5].n42 XThR.Tn[5].t38 145.038
R19794 XThR.Tn[5].n37 XThR.Tn[5].t69 145.038
R19795 XThR.Tn[5].n32 XThR.Tn[5].t30 145.038
R19796 XThR.Tn[5].n27 XThR.Tn[5].t55 145.038
R19797 XThR.Tn[5].n22 XThR.Tn[5].t28 145.038
R19798 XThR.Tn[5].n17 XThR.Tn[5].t73 145.038
R19799 XThR.Tn[5].n12 XThR.Tn[5].t39 145.038
R19800 XThR.Tn[5].n10 XThR.Tn[5].t17 145.038
R19801 XThR.Tn[5].n83 XThR.Tn[5].t27 143.911
R19802 XThR.Tn[5].n78 XThR.Tn[5].t50 143.911
R19803 XThR.Tn[5].n73 XThR.Tn[5].t34 143.911
R19804 XThR.Tn[5].n68 XThR.Tn[5].t15 143.911
R19805 XThR.Tn[5].n63 XThR.Tn[5].t44 143.911
R19806 XThR.Tn[5].n58 XThR.Tn[5].t25 143.911
R19807 XThR.Tn[5].n53 XThR.Tn[5].t36 143.911
R19808 XThR.Tn[5].n48 XThR.Tn[5].t16 143.911
R19809 XThR.Tn[5].n43 XThR.Tn[5].t14 143.911
R19810 XThR.Tn[5].n38 XThR.Tn[5].t43 143.911
R19811 XThR.Tn[5].n33 XThR.Tn[5].t67 143.911
R19812 XThR.Tn[5].n28 XThR.Tn[5].t33 143.911
R19813 XThR.Tn[5].n23 XThR.Tn[5].t65 143.911
R19814 XThR.Tn[5].n18 XThR.Tn[5].t48 143.911
R19815 XThR.Tn[5].n13 XThR.Tn[5].t13 143.911
R19816 XThR.Tn[5].n7 XThR.Tn[5].n5 135.249
R19817 XThR.Tn[5].n9 XThR.Tn[5].n3 98.981
R19818 XThR.Tn[5].n8 XThR.Tn[5].n4 98.981
R19819 XThR.Tn[5].n7 XThR.Tn[5].n6 98.981
R19820 XThR.Tn[5].n9 XThR.Tn[5].n8 36.2672
R19821 XThR.Tn[5].n8 XThR.Tn[5].n7 36.2672
R19822 XThR.Tn[5].n88 XThR.Tn[5].n9 32.6405
R19823 XThR.Tn[5].n1 XThR.Tn[5].t5 26.5955
R19824 XThR.Tn[5].n1 XThR.Tn[5].t4 26.5955
R19825 XThR.Tn[5].n0 XThR.Tn[5].t6 26.5955
R19826 XThR.Tn[5].n0 XThR.Tn[5].t7 26.5955
R19827 XThR.Tn[5].n3 XThR.Tn[5].t11 24.9236
R19828 XThR.Tn[5].n3 XThR.Tn[5].t8 24.9236
R19829 XThR.Tn[5].n4 XThR.Tn[5].t10 24.9236
R19830 XThR.Tn[5].n4 XThR.Tn[5].t9 24.9236
R19831 XThR.Tn[5].n5 XThR.Tn[5].t0 24.9236
R19832 XThR.Tn[5].n5 XThR.Tn[5].t1 24.9236
R19833 XThR.Tn[5].n6 XThR.Tn[5].t3 24.9236
R19834 XThR.Tn[5].n6 XThR.Tn[5].t2 24.9236
R19835 XThR.Tn[5].n89 XThR.Tn[5].n2 18.5605
R19836 XThR.Tn[5].n89 XThR.Tn[5].n88 11.5205
R19837 XThR.Tn[5].n88 XThR.Tn[5] 5.71508
R19838 XThR.Tn[5] XThR.Tn[5].n11 5.34038
R19839 XThR.Tn[5].n16 XThR.Tn[5].n15 4.5005
R19840 XThR.Tn[5].n21 XThR.Tn[5].n20 4.5005
R19841 XThR.Tn[5].n26 XThR.Tn[5].n25 4.5005
R19842 XThR.Tn[5].n31 XThR.Tn[5].n30 4.5005
R19843 XThR.Tn[5].n36 XThR.Tn[5].n35 4.5005
R19844 XThR.Tn[5].n41 XThR.Tn[5].n40 4.5005
R19845 XThR.Tn[5].n46 XThR.Tn[5].n45 4.5005
R19846 XThR.Tn[5].n51 XThR.Tn[5].n50 4.5005
R19847 XThR.Tn[5].n56 XThR.Tn[5].n55 4.5005
R19848 XThR.Tn[5].n61 XThR.Tn[5].n60 4.5005
R19849 XThR.Tn[5].n66 XThR.Tn[5].n65 4.5005
R19850 XThR.Tn[5].n71 XThR.Tn[5].n70 4.5005
R19851 XThR.Tn[5].n76 XThR.Tn[5].n75 4.5005
R19852 XThR.Tn[5].n81 XThR.Tn[5].n80 4.5005
R19853 XThR.Tn[5].n86 XThR.Tn[5].n85 4.5005
R19854 XThR.Tn[5].n87 XThR.Tn[5] 3.70586
R19855 XThR.Tn[5].n16 XThR.Tn[5] 2.52282
R19856 XThR.Tn[5].n21 XThR.Tn[5] 2.52282
R19857 XThR.Tn[5].n26 XThR.Tn[5] 2.52282
R19858 XThR.Tn[5].n31 XThR.Tn[5] 2.52282
R19859 XThR.Tn[5].n36 XThR.Tn[5] 2.52282
R19860 XThR.Tn[5].n41 XThR.Tn[5] 2.52282
R19861 XThR.Tn[5].n46 XThR.Tn[5] 2.52282
R19862 XThR.Tn[5].n51 XThR.Tn[5] 2.52282
R19863 XThR.Tn[5].n56 XThR.Tn[5] 2.52282
R19864 XThR.Tn[5].n61 XThR.Tn[5] 2.52282
R19865 XThR.Tn[5].n66 XThR.Tn[5] 2.52282
R19866 XThR.Tn[5].n71 XThR.Tn[5] 2.52282
R19867 XThR.Tn[5].n76 XThR.Tn[5] 2.52282
R19868 XThR.Tn[5].n81 XThR.Tn[5] 2.52282
R19869 XThR.Tn[5].n86 XThR.Tn[5] 2.52282
R19870 XThR.Tn[5].n84 XThR.Tn[5] 1.08677
R19871 XThR.Tn[5].n79 XThR.Tn[5] 1.08677
R19872 XThR.Tn[5].n74 XThR.Tn[5] 1.08677
R19873 XThR.Tn[5].n69 XThR.Tn[5] 1.08677
R19874 XThR.Tn[5].n64 XThR.Tn[5] 1.08677
R19875 XThR.Tn[5].n59 XThR.Tn[5] 1.08677
R19876 XThR.Tn[5].n54 XThR.Tn[5] 1.08677
R19877 XThR.Tn[5].n49 XThR.Tn[5] 1.08677
R19878 XThR.Tn[5].n44 XThR.Tn[5] 1.08677
R19879 XThR.Tn[5].n39 XThR.Tn[5] 1.08677
R19880 XThR.Tn[5].n34 XThR.Tn[5] 1.08677
R19881 XThR.Tn[5].n29 XThR.Tn[5] 1.08677
R19882 XThR.Tn[5].n24 XThR.Tn[5] 1.08677
R19883 XThR.Tn[5].n19 XThR.Tn[5] 1.08677
R19884 XThR.Tn[5].n14 XThR.Tn[5] 1.08677
R19885 XThR.Tn[5] XThR.Tn[5].n16 0.839786
R19886 XThR.Tn[5] XThR.Tn[5].n21 0.839786
R19887 XThR.Tn[5] XThR.Tn[5].n26 0.839786
R19888 XThR.Tn[5] XThR.Tn[5].n31 0.839786
R19889 XThR.Tn[5] XThR.Tn[5].n36 0.839786
R19890 XThR.Tn[5] XThR.Tn[5].n41 0.839786
R19891 XThR.Tn[5] XThR.Tn[5].n46 0.839786
R19892 XThR.Tn[5] XThR.Tn[5].n51 0.839786
R19893 XThR.Tn[5] XThR.Tn[5].n56 0.839786
R19894 XThR.Tn[5] XThR.Tn[5].n61 0.839786
R19895 XThR.Tn[5] XThR.Tn[5].n66 0.839786
R19896 XThR.Tn[5] XThR.Tn[5].n71 0.839786
R19897 XThR.Tn[5] XThR.Tn[5].n76 0.839786
R19898 XThR.Tn[5] XThR.Tn[5].n81 0.839786
R19899 XThR.Tn[5] XThR.Tn[5].n86 0.839786
R19900 XThR.Tn[5] XThR.Tn[5].n89 0.6405
R19901 XThR.Tn[5].n11 XThR.Tn[5] 0.499542
R19902 XThR.Tn[5].n85 XThR.Tn[5] 0.063
R19903 XThR.Tn[5].n80 XThR.Tn[5] 0.063
R19904 XThR.Tn[5].n75 XThR.Tn[5] 0.063
R19905 XThR.Tn[5].n70 XThR.Tn[5] 0.063
R19906 XThR.Tn[5].n65 XThR.Tn[5] 0.063
R19907 XThR.Tn[5].n60 XThR.Tn[5] 0.063
R19908 XThR.Tn[5].n55 XThR.Tn[5] 0.063
R19909 XThR.Tn[5].n50 XThR.Tn[5] 0.063
R19910 XThR.Tn[5].n45 XThR.Tn[5] 0.063
R19911 XThR.Tn[5].n40 XThR.Tn[5] 0.063
R19912 XThR.Tn[5].n35 XThR.Tn[5] 0.063
R19913 XThR.Tn[5].n30 XThR.Tn[5] 0.063
R19914 XThR.Tn[5].n25 XThR.Tn[5] 0.063
R19915 XThR.Tn[5].n20 XThR.Tn[5] 0.063
R19916 XThR.Tn[5].n15 XThR.Tn[5] 0.063
R19917 XThR.Tn[5].n87 XThR.Tn[5] 0.0540714
R19918 XThR.Tn[5] XThR.Tn[5].n87 0.038
R19919 XThR.Tn[5].n11 XThR.Tn[5] 0.0143889
R19920 XThR.Tn[5].n85 XThR.Tn[5].n84 0.00771154
R19921 XThR.Tn[5].n80 XThR.Tn[5].n79 0.00771154
R19922 XThR.Tn[5].n75 XThR.Tn[5].n74 0.00771154
R19923 XThR.Tn[5].n70 XThR.Tn[5].n69 0.00771154
R19924 XThR.Tn[5].n65 XThR.Tn[5].n64 0.00771154
R19925 XThR.Tn[5].n60 XThR.Tn[5].n59 0.00771154
R19926 XThR.Tn[5].n55 XThR.Tn[5].n54 0.00771154
R19927 XThR.Tn[5].n50 XThR.Tn[5].n49 0.00771154
R19928 XThR.Tn[5].n45 XThR.Tn[5].n44 0.00771154
R19929 XThR.Tn[5].n40 XThR.Tn[5].n39 0.00771154
R19930 XThR.Tn[5].n35 XThR.Tn[5].n34 0.00771154
R19931 XThR.Tn[5].n30 XThR.Tn[5].n29 0.00771154
R19932 XThR.Tn[5].n25 XThR.Tn[5].n24 0.00771154
R19933 XThR.Tn[5].n20 XThR.Tn[5].n19 0.00771154
R19934 XThR.Tn[5].n15 XThR.Tn[5].n14 0.00771154
R19935 XThC.Tn[4].n2 XThC.Tn[4].n1 332.332
R19936 XThC.Tn[4].n2 XThC.Tn[4].n0 296.493
R19937 XThC.Tn[4].n12 XThC.Tn[4].n10 161.406
R19938 XThC.Tn[4].n15 XThC.Tn[4].n13 161.406
R19939 XThC.Tn[4].n18 XThC.Tn[4].n16 161.406
R19940 XThC.Tn[4].n21 XThC.Tn[4].n19 161.406
R19941 XThC.Tn[4].n24 XThC.Tn[4].n22 161.406
R19942 XThC.Tn[4].n27 XThC.Tn[4].n25 161.406
R19943 XThC.Tn[4].n30 XThC.Tn[4].n28 161.406
R19944 XThC.Tn[4].n33 XThC.Tn[4].n31 161.406
R19945 XThC.Tn[4].n36 XThC.Tn[4].n34 161.406
R19946 XThC.Tn[4].n39 XThC.Tn[4].n37 161.406
R19947 XThC.Tn[4].n42 XThC.Tn[4].n40 161.406
R19948 XThC.Tn[4].n45 XThC.Tn[4].n43 161.406
R19949 XThC.Tn[4].n48 XThC.Tn[4].n46 161.406
R19950 XThC.Tn[4].n51 XThC.Tn[4].n49 161.406
R19951 XThC.Tn[4].n54 XThC.Tn[4].n52 161.406
R19952 XThC.Tn[4].n57 XThC.Tn[4].n55 161.406
R19953 XThC.Tn[4].n10 XThC.Tn[4].t26 161.202
R19954 XThC.Tn[4].n13 XThC.Tn[4].t43 161.202
R19955 XThC.Tn[4].n16 XThC.Tn[4].t13 161.202
R19956 XThC.Tn[4].n19 XThC.Tn[4].t15 161.202
R19957 XThC.Tn[4].n22 XThC.Tn[4].t36 161.202
R19958 XThC.Tn[4].n25 XThC.Tn[4].t37 161.202
R19959 XThC.Tn[4].n28 XThC.Tn[4].t18 161.202
R19960 XThC.Tn[4].n31 XThC.Tn[4].t27 161.202
R19961 XThC.Tn[4].n34 XThC.Tn[4].t29 161.202
R19962 XThC.Tn[4].n37 XThC.Tn[4].t16 161.202
R19963 XThC.Tn[4].n40 XThC.Tn[4].t17 161.202
R19964 XThC.Tn[4].n43 XThC.Tn[4].t30 161.202
R19965 XThC.Tn[4].n46 XThC.Tn[4].t38 161.202
R19966 XThC.Tn[4].n49 XThC.Tn[4].t41 161.202
R19967 XThC.Tn[4].n52 XThC.Tn[4].t22 161.202
R19968 XThC.Tn[4].n55 XThC.Tn[4].t32 161.202
R19969 XThC.Tn[4].n10 XThC.Tn[4].t28 145.137
R19970 XThC.Tn[4].n13 XThC.Tn[4].t14 145.137
R19971 XThC.Tn[4].n16 XThC.Tn[4].t19 145.137
R19972 XThC.Tn[4].n19 XThC.Tn[4].t20 145.137
R19973 XThC.Tn[4].n22 XThC.Tn[4].t39 145.137
R19974 XThC.Tn[4].n25 XThC.Tn[4].t40 145.137
R19975 XThC.Tn[4].n28 XThC.Tn[4].t24 145.137
R19976 XThC.Tn[4].n31 XThC.Tn[4].t31 145.137
R19977 XThC.Tn[4].n34 XThC.Tn[4].t33 145.137
R19978 XThC.Tn[4].n37 XThC.Tn[4].t21 145.137
R19979 XThC.Tn[4].n40 XThC.Tn[4].t23 145.137
R19980 XThC.Tn[4].n43 XThC.Tn[4].t34 145.137
R19981 XThC.Tn[4].n46 XThC.Tn[4].t42 145.137
R19982 XThC.Tn[4].n49 XThC.Tn[4].t12 145.137
R19983 XThC.Tn[4].n52 XThC.Tn[4].t25 145.137
R19984 XThC.Tn[4].n55 XThC.Tn[4].t35 145.137
R19985 XThC.Tn[4].n7 XThC.Tn[4].n6 135.248
R19986 XThC.Tn[4].n9 XThC.Tn[4].n3 98.982
R19987 XThC.Tn[4].n8 XThC.Tn[4].n4 98.982
R19988 XThC.Tn[4].n7 XThC.Tn[4].n5 98.982
R19989 XThC.Tn[4].n9 XThC.Tn[4].n8 36.2672
R19990 XThC.Tn[4].n8 XThC.Tn[4].n7 36.2672
R19991 XThC.Tn[4].n59 XThC.Tn[4].n9 32.6405
R19992 XThC.Tn[4].n1 XThC.Tn[4].t11 26.5955
R19993 XThC.Tn[4].n1 XThC.Tn[4].t10 26.5955
R19994 XThC.Tn[4].n0 XThC.Tn[4].t9 26.5955
R19995 XThC.Tn[4].n0 XThC.Tn[4].t8 26.5955
R19996 XThC.Tn[4].n3 XThC.Tn[4].t5 24.9236
R19997 XThC.Tn[4].n3 XThC.Tn[4].t4 24.9236
R19998 XThC.Tn[4].n4 XThC.Tn[4].t7 24.9236
R19999 XThC.Tn[4].n4 XThC.Tn[4].t6 24.9236
R20000 XThC.Tn[4].n5 XThC.Tn[4].t2 24.9236
R20001 XThC.Tn[4].n5 XThC.Tn[4].t1 24.9236
R20002 XThC.Tn[4].n6 XThC.Tn[4].t0 24.9236
R20003 XThC.Tn[4].n6 XThC.Tn[4].t3 24.9236
R20004 XThC.Tn[4].n60 XThC.Tn[4].n2 18.5605
R20005 XThC.Tn[4].n60 XThC.Tn[4].n59 11.5205
R20006 XThC.Tn[4].n58 XThC.Tn[4] 4.63701
R20007 XThC.Tn[4].n59 XThC.Tn[4].n58 3.1844
R20008 XThC.Tn[4].n15 XThC.Tn[4] 0.931056
R20009 XThC.Tn[4].n18 XThC.Tn[4] 0.931056
R20010 XThC.Tn[4].n21 XThC.Tn[4] 0.931056
R20011 XThC.Tn[4].n24 XThC.Tn[4] 0.931056
R20012 XThC.Tn[4].n27 XThC.Tn[4] 0.931056
R20013 XThC.Tn[4].n30 XThC.Tn[4] 0.931056
R20014 XThC.Tn[4].n33 XThC.Tn[4] 0.931056
R20015 XThC.Tn[4].n36 XThC.Tn[4] 0.931056
R20016 XThC.Tn[4].n39 XThC.Tn[4] 0.931056
R20017 XThC.Tn[4].n42 XThC.Tn[4] 0.931056
R20018 XThC.Tn[4].n45 XThC.Tn[4] 0.931056
R20019 XThC.Tn[4].n48 XThC.Tn[4] 0.931056
R20020 XThC.Tn[4].n51 XThC.Tn[4] 0.931056
R20021 XThC.Tn[4].n54 XThC.Tn[4] 0.931056
R20022 XThC.Tn[4].n57 XThC.Tn[4] 0.931056
R20023 XThC.Tn[4] XThC.Tn[4].n60 0.6405
R20024 XThC.Tn[4] XThC.Tn[4].n12 0.396333
R20025 XThC.Tn[4] XThC.Tn[4].n15 0.396333
R20026 XThC.Tn[4] XThC.Tn[4].n18 0.396333
R20027 XThC.Tn[4] XThC.Tn[4].n21 0.396333
R20028 XThC.Tn[4] XThC.Tn[4].n24 0.396333
R20029 XThC.Tn[4] XThC.Tn[4].n27 0.396333
R20030 XThC.Tn[4] XThC.Tn[4].n30 0.396333
R20031 XThC.Tn[4] XThC.Tn[4].n33 0.396333
R20032 XThC.Tn[4] XThC.Tn[4].n36 0.396333
R20033 XThC.Tn[4] XThC.Tn[4].n39 0.396333
R20034 XThC.Tn[4] XThC.Tn[4].n42 0.396333
R20035 XThC.Tn[4] XThC.Tn[4].n45 0.396333
R20036 XThC.Tn[4] XThC.Tn[4].n48 0.396333
R20037 XThC.Tn[4] XThC.Tn[4].n51 0.396333
R20038 XThC.Tn[4] XThC.Tn[4].n54 0.396333
R20039 XThC.Tn[4] XThC.Tn[4].n57 0.396333
R20040 XThC.Tn[4].n11 XThC.Tn[4] 0.104667
R20041 XThC.Tn[4].n14 XThC.Tn[4] 0.104667
R20042 XThC.Tn[4].n17 XThC.Tn[4] 0.104667
R20043 XThC.Tn[4].n20 XThC.Tn[4] 0.104667
R20044 XThC.Tn[4].n23 XThC.Tn[4] 0.104667
R20045 XThC.Tn[4].n26 XThC.Tn[4] 0.104667
R20046 XThC.Tn[4].n29 XThC.Tn[4] 0.104667
R20047 XThC.Tn[4].n32 XThC.Tn[4] 0.104667
R20048 XThC.Tn[4].n35 XThC.Tn[4] 0.104667
R20049 XThC.Tn[4].n38 XThC.Tn[4] 0.104667
R20050 XThC.Tn[4].n41 XThC.Tn[4] 0.104667
R20051 XThC.Tn[4].n44 XThC.Tn[4] 0.104667
R20052 XThC.Tn[4].n47 XThC.Tn[4] 0.104667
R20053 XThC.Tn[4].n50 XThC.Tn[4] 0.104667
R20054 XThC.Tn[4].n53 XThC.Tn[4] 0.104667
R20055 XThC.Tn[4].n56 XThC.Tn[4] 0.104667
R20056 XThC.Tn[4].n11 XThC.Tn[4] 0.0309878
R20057 XThC.Tn[4].n14 XThC.Tn[4] 0.0309878
R20058 XThC.Tn[4].n17 XThC.Tn[4] 0.0309878
R20059 XThC.Tn[4].n20 XThC.Tn[4] 0.0309878
R20060 XThC.Tn[4].n23 XThC.Tn[4] 0.0309878
R20061 XThC.Tn[4].n26 XThC.Tn[4] 0.0309878
R20062 XThC.Tn[4].n29 XThC.Tn[4] 0.0309878
R20063 XThC.Tn[4].n32 XThC.Tn[4] 0.0309878
R20064 XThC.Tn[4].n35 XThC.Tn[4] 0.0309878
R20065 XThC.Tn[4].n38 XThC.Tn[4] 0.0309878
R20066 XThC.Tn[4].n41 XThC.Tn[4] 0.0309878
R20067 XThC.Tn[4].n44 XThC.Tn[4] 0.0309878
R20068 XThC.Tn[4].n47 XThC.Tn[4] 0.0309878
R20069 XThC.Tn[4].n50 XThC.Tn[4] 0.0309878
R20070 XThC.Tn[4].n53 XThC.Tn[4] 0.0309878
R20071 XThC.Tn[4].n56 XThC.Tn[4] 0.0309878
R20072 XThC.Tn[4].n12 XThC.Tn[4].n11 0.027939
R20073 XThC.Tn[4].n15 XThC.Tn[4].n14 0.027939
R20074 XThC.Tn[4].n18 XThC.Tn[4].n17 0.027939
R20075 XThC.Tn[4].n21 XThC.Tn[4].n20 0.027939
R20076 XThC.Tn[4].n24 XThC.Tn[4].n23 0.027939
R20077 XThC.Tn[4].n27 XThC.Tn[4].n26 0.027939
R20078 XThC.Tn[4].n30 XThC.Tn[4].n29 0.027939
R20079 XThC.Tn[4].n33 XThC.Tn[4].n32 0.027939
R20080 XThC.Tn[4].n36 XThC.Tn[4].n35 0.027939
R20081 XThC.Tn[4].n39 XThC.Tn[4].n38 0.027939
R20082 XThC.Tn[4].n42 XThC.Tn[4].n41 0.027939
R20083 XThC.Tn[4].n45 XThC.Tn[4].n44 0.027939
R20084 XThC.Tn[4].n48 XThC.Tn[4].n47 0.027939
R20085 XThC.Tn[4].n51 XThC.Tn[4].n50 0.027939
R20086 XThC.Tn[4].n54 XThC.Tn[4].n53 0.027939
R20087 XThC.Tn[4].n57 XThC.Tn[4].n56 0.027939
R20088 XThC.Tn[4].n58 XThC.Tn[4] 0.0129465
R20089 XThC.Tn[2].n2 XThC.Tn[2].n1 332.332
R20090 XThC.Tn[2].n2 XThC.Tn[2].n0 296.493
R20091 XThC.Tn[2].n12 XThC.Tn[2].n10 161.406
R20092 XThC.Tn[2].n15 XThC.Tn[2].n13 161.406
R20093 XThC.Tn[2].n18 XThC.Tn[2].n16 161.406
R20094 XThC.Tn[2].n21 XThC.Tn[2].n19 161.406
R20095 XThC.Tn[2].n24 XThC.Tn[2].n22 161.406
R20096 XThC.Tn[2].n27 XThC.Tn[2].n25 161.406
R20097 XThC.Tn[2].n30 XThC.Tn[2].n28 161.406
R20098 XThC.Tn[2].n33 XThC.Tn[2].n31 161.406
R20099 XThC.Tn[2].n36 XThC.Tn[2].n34 161.406
R20100 XThC.Tn[2].n39 XThC.Tn[2].n37 161.406
R20101 XThC.Tn[2].n42 XThC.Tn[2].n40 161.406
R20102 XThC.Tn[2].n45 XThC.Tn[2].n43 161.406
R20103 XThC.Tn[2].n48 XThC.Tn[2].n46 161.406
R20104 XThC.Tn[2].n51 XThC.Tn[2].n49 161.406
R20105 XThC.Tn[2].n54 XThC.Tn[2].n52 161.406
R20106 XThC.Tn[2].n57 XThC.Tn[2].n55 161.406
R20107 XThC.Tn[2].n10 XThC.Tn[2].t18 161.202
R20108 XThC.Tn[2].n13 XThC.Tn[2].t35 161.202
R20109 XThC.Tn[2].n16 XThC.Tn[2].t37 161.202
R20110 XThC.Tn[2].n19 XThC.Tn[2].t39 161.202
R20111 XThC.Tn[2].n22 XThC.Tn[2].t28 161.202
R20112 XThC.Tn[2].n25 XThC.Tn[2].t29 161.202
R20113 XThC.Tn[2].n28 XThC.Tn[2].t42 161.202
R20114 XThC.Tn[2].n31 XThC.Tn[2].t19 161.202
R20115 XThC.Tn[2].n34 XThC.Tn[2].t21 161.202
R20116 XThC.Tn[2].n37 XThC.Tn[2].t40 161.202
R20117 XThC.Tn[2].n40 XThC.Tn[2].t41 161.202
R20118 XThC.Tn[2].n43 XThC.Tn[2].t22 161.202
R20119 XThC.Tn[2].n46 XThC.Tn[2].t30 161.202
R20120 XThC.Tn[2].n49 XThC.Tn[2].t33 161.202
R20121 XThC.Tn[2].n52 XThC.Tn[2].t14 161.202
R20122 XThC.Tn[2].n55 XThC.Tn[2].t24 161.202
R20123 XThC.Tn[2].n10 XThC.Tn[2].t20 145.137
R20124 XThC.Tn[2].n13 XThC.Tn[2].t38 145.137
R20125 XThC.Tn[2].n16 XThC.Tn[2].t43 145.137
R20126 XThC.Tn[2].n19 XThC.Tn[2].t12 145.137
R20127 XThC.Tn[2].n22 XThC.Tn[2].t31 145.137
R20128 XThC.Tn[2].n25 XThC.Tn[2].t32 145.137
R20129 XThC.Tn[2].n28 XThC.Tn[2].t16 145.137
R20130 XThC.Tn[2].n31 XThC.Tn[2].t23 145.137
R20131 XThC.Tn[2].n34 XThC.Tn[2].t25 145.137
R20132 XThC.Tn[2].n37 XThC.Tn[2].t13 145.137
R20133 XThC.Tn[2].n40 XThC.Tn[2].t15 145.137
R20134 XThC.Tn[2].n43 XThC.Tn[2].t26 145.137
R20135 XThC.Tn[2].n46 XThC.Tn[2].t34 145.137
R20136 XThC.Tn[2].n49 XThC.Tn[2].t36 145.137
R20137 XThC.Tn[2].n52 XThC.Tn[2].t17 145.137
R20138 XThC.Tn[2].n55 XThC.Tn[2].t27 145.137
R20139 XThC.Tn[2].n7 XThC.Tn[2].n6 135.248
R20140 XThC.Tn[2].n9 XThC.Tn[2].n3 98.982
R20141 XThC.Tn[2].n8 XThC.Tn[2].n4 98.982
R20142 XThC.Tn[2].n7 XThC.Tn[2].n5 98.982
R20143 XThC.Tn[2].n9 XThC.Tn[2].n8 36.2672
R20144 XThC.Tn[2].n8 XThC.Tn[2].n7 36.2672
R20145 XThC.Tn[2].n59 XThC.Tn[2].n9 32.6405
R20146 XThC.Tn[2].n1 XThC.Tn[2].t5 26.5955
R20147 XThC.Tn[2].n1 XThC.Tn[2].t4 26.5955
R20148 XThC.Tn[2].n0 XThC.Tn[2].t7 26.5955
R20149 XThC.Tn[2].n0 XThC.Tn[2].t6 26.5955
R20150 XThC.Tn[2].n3 XThC.Tn[2].t11 24.9236
R20151 XThC.Tn[2].n3 XThC.Tn[2].t10 24.9236
R20152 XThC.Tn[2].n4 XThC.Tn[2].t9 24.9236
R20153 XThC.Tn[2].n4 XThC.Tn[2].t8 24.9236
R20154 XThC.Tn[2].n5 XThC.Tn[2].t1 24.9236
R20155 XThC.Tn[2].n5 XThC.Tn[2].t2 24.9236
R20156 XThC.Tn[2].n6 XThC.Tn[2].t3 24.9236
R20157 XThC.Tn[2].n6 XThC.Tn[2].t0 24.9236
R20158 XThC.Tn[2].n60 XThC.Tn[2].n2 18.5605
R20159 XThC.Tn[2].n60 XThC.Tn[2].n59 11.5205
R20160 XThC.Tn[2].n58 XThC.Tn[2] 6.32799
R20161 XThC.Tn[2].n59 XThC.Tn[2].n58 3.18175
R20162 XThC.Tn[2].n15 XThC.Tn[2] 0.931056
R20163 XThC.Tn[2].n18 XThC.Tn[2] 0.931056
R20164 XThC.Tn[2].n21 XThC.Tn[2] 0.931056
R20165 XThC.Tn[2].n24 XThC.Tn[2] 0.931056
R20166 XThC.Tn[2].n27 XThC.Tn[2] 0.931056
R20167 XThC.Tn[2].n30 XThC.Tn[2] 0.931056
R20168 XThC.Tn[2].n33 XThC.Tn[2] 0.931056
R20169 XThC.Tn[2].n36 XThC.Tn[2] 0.931056
R20170 XThC.Tn[2].n39 XThC.Tn[2] 0.931056
R20171 XThC.Tn[2].n42 XThC.Tn[2] 0.931056
R20172 XThC.Tn[2].n45 XThC.Tn[2] 0.931056
R20173 XThC.Tn[2].n48 XThC.Tn[2] 0.931056
R20174 XThC.Tn[2].n51 XThC.Tn[2] 0.931056
R20175 XThC.Tn[2].n54 XThC.Tn[2] 0.931056
R20176 XThC.Tn[2].n57 XThC.Tn[2] 0.931056
R20177 XThC.Tn[2] XThC.Tn[2].n60 0.6405
R20178 XThC.Tn[2] XThC.Tn[2].n12 0.396333
R20179 XThC.Tn[2] XThC.Tn[2].n15 0.396333
R20180 XThC.Tn[2] XThC.Tn[2].n18 0.396333
R20181 XThC.Tn[2] XThC.Tn[2].n21 0.396333
R20182 XThC.Tn[2] XThC.Tn[2].n24 0.396333
R20183 XThC.Tn[2] XThC.Tn[2].n27 0.396333
R20184 XThC.Tn[2] XThC.Tn[2].n30 0.396333
R20185 XThC.Tn[2] XThC.Tn[2].n33 0.396333
R20186 XThC.Tn[2] XThC.Tn[2].n36 0.396333
R20187 XThC.Tn[2] XThC.Tn[2].n39 0.396333
R20188 XThC.Tn[2] XThC.Tn[2].n42 0.396333
R20189 XThC.Tn[2] XThC.Tn[2].n45 0.396333
R20190 XThC.Tn[2] XThC.Tn[2].n48 0.396333
R20191 XThC.Tn[2] XThC.Tn[2].n51 0.396333
R20192 XThC.Tn[2] XThC.Tn[2].n54 0.396333
R20193 XThC.Tn[2] XThC.Tn[2].n57 0.396333
R20194 XThC.Tn[2].n11 XThC.Tn[2] 0.104667
R20195 XThC.Tn[2].n14 XThC.Tn[2] 0.104667
R20196 XThC.Tn[2].n17 XThC.Tn[2] 0.104667
R20197 XThC.Tn[2].n20 XThC.Tn[2] 0.104667
R20198 XThC.Tn[2].n23 XThC.Tn[2] 0.104667
R20199 XThC.Tn[2].n26 XThC.Tn[2] 0.104667
R20200 XThC.Tn[2].n29 XThC.Tn[2] 0.104667
R20201 XThC.Tn[2].n32 XThC.Tn[2] 0.104667
R20202 XThC.Tn[2].n35 XThC.Tn[2] 0.104667
R20203 XThC.Tn[2].n38 XThC.Tn[2] 0.104667
R20204 XThC.Tn[2].n41 XThC.Tn[2] 0.104667
R20205 XThC.Tn[2].n44 XThC.Tn[2] 0.104667
R20206 XThC.Tn[2].n47 XThC.Tn[2] 0.104667
R20207 XThC.Tn[2].n50 XThC.Tn[2] 0.104667
R20208 XThC.Tn[2].n53 XThC.Tn[2] 0.104667
R20209 XThC.Tn[2].n56 XThC.Tn[2] 0.104667
R20210 XThC.Tn[2].n11 XThC.Tn[2] 0.0309878
R20211 XThC.Tn[2].n14 XThC.Tn[2] 0.0309878
R20212 XThC.Tn[2].n17 XThC.Tn[2] 0.0309878
R20213 XThC.Tn[2].n20 XThC.Tn[2] 0.0309878
R20214 XThC.Tn[2].n23 XThC.Tn[2] 0.0309878
R20215 XThC.Tn[2].n26 XThC.Tn[2] 0.0309878
R20216 XThC.Tn[2].n29 XThC.Tn[2] 0.0309878
R20217 XThC.Tn[2].n32 XThC.Tn[2] 0.0309878
R20218 XThC.Tn[2].n35 XThC.Tn[2] 0.0309878
R20219 XThC.Tn[2].n38 XThC.Tn[2] 0.0309878
R20220 XThC.Tn[2].n41 XThC.Tn[2] 0.0309878
R20221 XThC.Tn[2].n44 XThC.Tn[2] 0.0309878
R20222 XThC.Tn[2].n47 XThC.Tn[2] 0.0309878
R20223 XThC.Tn[2].n50 XThC.Tn[2] 0.0309878
R20224 XThC.Tn[2].n53 XThC.Tn[2] 0.0309878
R20225 XThC.Tn[2].n56 XThC.Tn[2] 0.0309878
R20226 XThC.Tn[2].n12 XThC.Tn[2].n11 0.027939
R20227 XThC.Tn[2].n15 XThC.Tn[2].n14 0.027939
R20228 XThC.Tn[2].n18 XThC.Tn[2].n17 0.027939
R20229 XThC.Tn[2].n21 XThC.Tn[2].n20 0.027939
R20230 XThC.Tn[2].n24 XThC.Tn[2].n23 0.027939
R20231 XThC.Tn[2].n27 XThC.Tn[2].n26 0.027939
R20232 XThC.Tn[2].n30 XThC.Tn[2].n29 0.027939
R20233 XThC.Tn[2].n33 XThC.Tn[2].n32 0.027939
R20234 XThC.Tn[2].n36 XThC.Tn[2].n35 0.027939
R20235 XThC.Tn[2].n39 XThC.Tn[2].n38 0.027939
R20236 XThC.Tn[2].n42 XThC.Tn[2].n41 0.027939
R20237 XThC.Tn[2].n45 XThC.Tn[2].n44 0.027939
R20238 XThC.Tn[2].n48 XThC.Tn[2].n47 0.027939
R20239 XThC.Tn[2].n51 XThC.Tn[2].n50 0.027939
R20240 XThC.Tn[2].n54 XThC.Tn[2].n53 0.027939
R20241 XThC.Tn[2].n57 XThC.Tn[2].n56 0.027939
R20242 XThC.Tn[2].n58 XThC.Tn[2] 0.0156819
R20243 Vbias.t4 Vbias.n512 313.474
R20244 Vbias.t6 Vbias.n518 313.464
R20245 Vbias.n516 Vbias.t4 313.13
R20246 Vbias.n522 Vbias.t6 313.13
R20247 Vbias.n515 Vbias.n514 299.471
R20248 Vbias.n521 Vbias.n520 299.471
R20249 Vbias.n515 Vbias.n513 299.144
R20250 Vbias.n521 Vbias.n519 299.144
R20251 Vbias.n509 Vbias.t187 119.309
R20252 Vbias.n507 Vbias.t30 119.309
R20253 Vbias.n505 Vbias.t18 119.309
R20254 Vbias.n503 Vbias.t254 119.309
R20255 Vbias.n501 Vbias.t101 119.309
R20256 Vbias.n499 Vbias.t81 119.309
R20257 Vbias.n497 Vbias.t252 119.309
R20258 Vbias.n495 Vbias.t175 119.309
R20259 Vbias.n493 Vbias.t153 119.309
R20260 Vbias.n491 Vbias.t66 119.309
R20261 Vbias.n489 Vbias.t233 119.309
R20262 Vbias.n487 Vbias.t147 119.309
R20263 Vbias.n485 Vbias.t62 119.309
R20264 Vbias.n483 Vbias.t47 119.309
R20265 Vbias.n481 Vbias.t207 119.309
R20266 Vbias.n480 Vbias.t135 119.309
R20267 Vbias.n477 Vbias.t116 119.309
R20268 Vbias.n475 Vbias.t216 119.309
R20269 Vbias.n473 Vbias.t199 119.309
R20270 Vbias.n471 Vbias.t179 119.309
R20271 Vbias.n469 Vbias.t31 119.309
R20272 Vbias.n467 Vbias.t264 119.309
R20273 Vbias.n465 Vbias.t177 119.309
R20274 Vbias.n463 Vbias.t102 119.309
R20275 Vbias.n461 Vbias.t82 119.309
R20276 Vbias.n459 Vbias.t253 119.309
R20277 Vbias.n457 Vbias.t162 119.309
R20278 Vbias.n455 Vbias.t75 119.309
R20279 Vbias.n453 Vbias.t248 119.309
R20280 Vbias.n451 Vbias.t235 119.309
R20281 Vbias.n449 Vbias.t136 119.309
R20282 Vbias.n448 Vbias.t63 119.309
R20283 Vbias.n445 Vbias.t152 119.309
R20284 Vbias.n443 Vbias.t244 119.309
R20285 Vbias.n441 Vbias.t231 119.309
R20286 Vbias.n439 Vbias.t211 119.309
R20287 Vbias.n437 Vbias.t58 119.309
R20288 Vbias.n435 Vbias.t38 119.309
R20289 Vbias.n433 Vbias.t205 119.309
R20290 Vbias.n431 Vbias.t131 119.309
R20291 Vbias.n429 Vbias.t108 119.309
R20292 Vbias.n427 Vbias.t24 119.309
R20293 Vbias.n425 Vbias.t189 119.309
R20294 Vbias.n423 Vbias.t105 119.309
R20295 Vbias.n421 Vbias.t20 119.309
R20296 Vbias.n419 Vbias.t267 119.309
R20297 Vbias.n417 Vbias.t166 119.309
R20298 Vbias.n416 Vbias.t93 119.309
R20299 Vbias.n413 Vbias.t79 119.309
R20300 Vbias.n411 Vbias.t171 119.309
R20301 Vbias.n409 Vbias.t159 119.309
R20302 Vbias.n407 Vbias.t139 119.309
R20303 Vbias.n405 Vbias.t245 119.309
R20304 Vbias.n403 Vbias.t223 119.309
R20305 Vbias.n401 Vbias.t132 119.309
R20306 Vbias.n399 Vbias.t59 119.309
R20307 Vbias.n397 Vbias.t39 119.309
R20308 Vbias.n395 Vbias.t206 119.309
R20309 Vbias.n393 Vbias.t118 119.309
R20310 Vbias.n391 Vbias.t35 119.309
R20311 Vbias.n389 Vbias.t202 119.309
R20312 Vbias.n387 Vbias.t191 119.309
R20313 Vbias.n385 Vbias.t94 119.309
R20314 Vbias.n384 Vbias.t22 119.309
R20315 Vbias.n381 Vbias.t261 119.309
R20316 Vbias.n379 Vbias.t98 119.309
R20317 Vbias.n377 Vbias.t87 119.309
R20318 Vbias.n375 Vbias.t68 119.309
R20319 Vbias.n373 Vbias.t172 119.309
R20320 Vbias.n371 Vbias.t150 119.309
R20321 Vbias.n369 Vbias.t60 119.309
R20322 Vbias.n367 Vbias.t246 119.309
R20323 Vbias.n365 Vbias.t225 119.309
R20324 Vbias.n363 Vbias.t133 119.309
R20325 Vbias.n361 Vbias.t46 119.309
R20326 Vbias.n359 Vbias.t219 119.309
R20327 Vbias.n357 Vbias.t130 119.309
R20328 Vbias.n355 Vbias.t119 119.309
R20329 Vbias.n353 Vbias.t23 119.309
R20330 Vbias.n352 Vbias.t204 119.309
R20331 Vbias.n349 Vbias.t182 119.309
R20332 Vbias.n347 Vbias.t26 119.309
R20333 Vbias.n345 Vbias.t13 119.309
R20334 Vbias.n343 Vbias.t249 119.309
R20335 Vbias.n341 Vbias.t96 119.309
R20336 Vbias.n339 Vbias.t71 119.309
R20337 Vbias.n337 Vbias.t242 119.309
R20338 Vbias.n335 Vbias.t169 119.309
R20339 Vbias.n333 Vbias.t144 119.309
R20340 Vbias.n331 Vbias.t56 119.309
R20341 Vbias.n329 Vbias.t227 119.309
R20342 Vbias.n327 Vbias.t141 119.309
R20343 Vbias.n325 Vbias.t54 119.309
R20344 Vbias.n323 Vbias.t43 119.309
R20345 Vbias.n321 Vbias.t201 119.309
R20346 Vbias.n320 Vbias.t127 119.309
R20347 Vbias.n317 Vbias.t111 119.309
R20348 Vbias.n315 Vbias.t210 119.309
R20349 Vbias.n313 Vbias.t193 119.309
R20350 Vbias.n311 Vbias.t174 119.309
R20351 Vbias.n309 Vbias.t27 119.309
R20352 Vbias.n307 Vbias.t257 119.309
R20353 Vbias.n305 Vbias.t170 119.309
R20354 Vbias.n303 Vbias.t97 119.309
R20355 Vbias.n301 Vbias.t74 119.309
R20356 Vbias.n299 Vbias.t243 119.309
R20357 Vbias.n297 Vbias.t156 119.309
R20358 Vbias.n295 Vbias.t69 119.309
R20359 Vbias.n293 Vbias.t241 119.309
R20360 Vbias.n291 Vbias.t228 119.309
R20361 Vbias.n289 Vbias.t128 119.309
R20362 Vbias.n288 Vbias.t55 119.309
R20363 Vbias.n285 Vbias.t143 119.309
R20364 Vbias.n283 Vbias.t238 119.309
R20365 Vbias.n281 Vbias.t226 119.309
R20366 Vbias.n279 Vbias.t203 119.309
R20367 Vbias.n277 Vbias.t50 119.309
R20368 Vbias.n275 Vbias.t33 119.309
R20369 Vbias.n273 Vbias.t196 119.309
R20370 Vbias.n271 Vbias.t124 119.309
R20371 Vbias.n269 Vbias.t104 119.309
R20372 Vbias.n267 Vbias.t17 119.309
R20373 Vbias.n265 Vbias.t185 119.309
R20374 Vbias.n263 Vbias.t99 119.309
R20375 Vbias.n261 Vbias.t14 119.309
R20376 Vbias.n259 Vbias.t263 119.309
R20377 Vbias.n257 Vbias.t160 119.309
R20378 Vbias.n256 Vbias.t88 119.309
R20379 Vbias.n253 Vbias.t70 119.309
R20380 Vbias.n251 Vbias.t167 119.309
R20381 Vbias.n249 Vbias.t155 119.309
R20382 Vbias.n247 Vbias.t129 119.309
R20383 Vbias.n245 Vbias.t239 119.309
R20384 Vbias.n243 Vbias.t217 119.309
R20385 Vbias.n241 Vbias.t125 119.309
R20386 Vbias.n239 Vbias.t51 119.309
R20387 Vbias.n237 Vbias.t34 119.309
R20388 Vbias.n235 Vbias.t198 119.309
R20389 Vbias.n233 Vbias.t113 119.309
R20390 Vbias.n231 Vbias.t29 119.309
R20391 Vbias.n229 Vbias.t194 119.309
R20392 Vbias.n227 Vbias.t186 119.309
R20393 Vbias.n225 Vbias.t89 119.309
R20394 Vbias.n224 Vbias.t15 119.309
R20395 Vbias.n221 Vbias.t256 119.309
R20396 Vbias.n219 Vbias.t95 119.309
R20397 Vbias.n217 Vbias.t86 119.309
R20398 Vbias.n215 Vbias.t57 119.309
R20399 Vbias.n213 Vbias.t168 119.309
R20400 Vbias.n211 Vbias.t142 119.309
R20401 Vbias.n209 Vbias.t52 119.309
R20402 Vbias.n207 Vbias.t240 119.309
R20403 Vbias.n205 Vbias.t218 119.309
R20404 Vbias.n203 Vbias.t126 119.309
R20405 Vbias.n201 Vbias.t42 119.309
R20406 Vbias.n199 Vbias.t214 119.309
R20407 Vbias.n197 Vbias.t123 119.309
R20408 Vbias.n195 Vbias.t114 119.309
R20409 Vbias.n193 Vbias.t16 119.309
R20410 Vbias.n192 Vbias.t195 119.309
R20411 Vbias.n189 Vbias.t115 119.309
R20412 Vbias.n187 Vbias.t213 119.309
R20413 Vbias.n185 Vbias.t197 119.309
R20414 Vbias.n183 Vbias.t178 119.309
R20415 Vbias.n181 Vbias.t28 119.309
R20416 Vbias.n179 Vbias.t262 119.309
R20417 Vbias.n177 Vbias.t173 119.309
R20418 Vbias.n175 Vbias.t100 119.309
R20419 Vbias.n173 Vbias.t80 119.309
R20420 Vbias.n171 Vbias.t250 119.309
R20421 Vbias.n169 Vbias.t161 119.309
R20422 Vbias.n167 Vbias.t72 119.309
R20423 Vbias.n165 Vbias.t247 119.309
R20424 Vbias.n163 Vbias.t232 119.309
R20425 Vbias.n161 Vbias.t134 119.309
R20426 Vbias.n160 Vbias.t61 119.309
R20427 Vbias.n157 Vbias.t255 119.309
R20428 Vbias.n155 Vbias.t91 119.309
R20429 Vbias.n153 Vbias.t84 119.309
R20430 Vbias.n151 Vbias.t53 119.309
R20431 Vbias.n149 Vbias.t165 119.309
R20432 Vbias.n147 Vbias.t140 119.309
R20433 Vbias.n145 Vbias.t49 119.309
R20434 Vbias.n143 Vbias.t237 119.309
R20435 Vbias.n141 Vbias.t215 119.309
R20436 Vbias.n139 Vbias.t122 119.309
R20437 Vbias.n137 Vbias.t40 119.309
R20438 Vbias.n135 Vbias.t212 119.309
R20439 Vbias.n133 Vbias.t121 119.309
R20440 Vbias.n131 Vbias.t109 119.309
R20441 Vbias.n129 Vbias.t12 119.309
R20442 Vbias.n128 Vbias.t192 119.309
R20443 Vbias.n125 Vbias.t92 119.309
R20444 Vbias.n123 Vbias.t181 119.309
R20445 Vbias.n121 Vbias.t176 119.309
R20446 Vbias.n119 Vbias.t154 119.309
R20447 Vbias.n117 Vbias.t258 119.309
R20448 Vbias.n115 Vbias.t234 119.309
R20449 Vbias.n113 Vbias.t149 119.309
R20450 Vbias.n111 Vbias.t76 119.309
R20451 Vbias.n109 Vbias.t48 119.309
R20452 Vbias.n107 Vbias.t224 119.309
R20453 Vbias.n105 Vbias.t137 119.309
R20454 Vbias.n103 Vbias.t44 119.309
R20455 Vbias.n101 Vbias.t220 119.309
R20456 Vbias.n99 Vbias.t209 119.309
R20457 Vbias.n97 Vbias.t106 119.309
R20458 Vbias.n96 Vbias.t36 119.309
R20459 Vbias.n93 Vbias.t19 119.309
R20460 Vbias.n91 Vbias.t110 119.309
R20461 Vbias.n89 Vbias.t103 119.309
R20462 Vbias.n87 Vbias.t83 119.309
R20463 Vbias.n85 Vbias.t183 119.309
R20464 Vbias.n83 Vbias.t163 119.309
R20465 Vbias.n81 Vbias.t77 119.309
R20466 Vbias.n79 Vbias.t259 119.309
R20467 Vbias.n77 Vbias.t236 119.309
R20468 Vbias.n75 Vbias.t151 119.309
R20469 Vbias.n73 Vbias.t64 119.309
R20470 Vbias.n71 Vbias.t230 119.309
R20471 Vbias.n69 Vbias.t145 119.309
R20472 Vbias.n67 Vbias.t138 119.309
R20473 Vbias.n65 Vbias.t37 119.309
R20474 Vbias.n64 Vbias.t221 119.309
R20475 Vbias.n61 Vbias.t200 119.309
R20476 Vbias.n59 Vbias.t41 119.309
R20477 Vbias.n57 Vbias.t32 119.309
R20478 Vbias.n55 Vbias.t265 119.309
R20479 Vbias.n53 Vbias.t112 119.309
R20480 Vbias.n51 Vbias.t90 119.309
R20481 Vbias.n49 Vbias.t260 119.309
R20482 Vbias.n47 Vbias.t184 119.309
R20483 Vbias.n45 Vbias.t164 119.309
R20484 Vbias.n43 Vbias.t78 119.309
R20485 Vbias.n41 Vbias.t251 119.309
R20486 Vbias.n39 Vbias.t158 119.309
R20487 Vbias.n37 Vbias.t73 119.309
R20488 Vbias.n35 Vbias.t65 119.309
R20489 Vbias.n33 Vbias.t222 119.309
R20490 Vbias.n32 Vbias.t146 119.309
R20491 Vbias.n29 Vbias.t67 119.309
R20492 Vbias.n27 Vbias.t157 119.309
R20493 Vbias.n25 Vbias.t148 119.309
R20494 Vbias.n23 Vbias.t120 119.309
R20495 Vbias.n21 Vbias.t229 119.309
R20496 Vbias.n19 Vbias.t208 119.309
R20497 Vbias.n17 Vbias.t117 119.309
R20498 Vbias.n15 Vbias.t45 119.309
R20499 Vbias.n13 Vbias.t25 119.309
R20500 Vbias.n11 Vbias.t190 119.309
R20501 Vbias.n9 Vbias.t107 119.309
R20502 Vbias.n7 Vbias.t21 119.309
R20503 Vbias.n5 Vbias.t188 119.309
R20504 Vbias.n3 Vbias.t180 119.309
R20505 Vbias.n1 Vbias.t85 119.309
R20506 Vbias.n0 Vbias.t266 119.309
R20507 Vbias.n513 Vbias.t9 53.3064
R20508 Vbias.n513 Vbias.t0 53.3064
R20509 Vbias.n519 Vbias.t3 53.3064
R20510 Vbias.n519 Vbias.t11 53.3064
R20511 Vbias.n512 Vbias.t5 34.1153
R20512 Vbias.n518 Vbias.t7 34.1153
R20513 Vbias.n514 Vbias.t2 33.6064
R20514 Vbias.n514 Vbias.t8 33.6064
R20515 Vbias.n520 Vbias.t1 33.6064
R20516 Vbias.n520 Vbias.t10 33.6064
R20517 Vbias Vbias.n480 8.00727
R20518 Vbias Vbias.n448 8.00727
R20519 Vbias Vbias.n416 8.00727
R20520 Vbias Vbias.n384 8.00727
R20521 Vbias Vbias.n352 8.00727
R20522 Vbias Vbias.n320 8.00727
R20523 Vbias Vbias.n288 8.00727
R20524 Vbias Vbias.n256 8.00727
R20525 Vbias Vbias.n224 8.00727
R20526 Vbias Vbias.n192 8.00727
R20527 Vbias Vbias.n160 8.00727
R20528 Vbias Vbias.n128 8.00727
R20529 Vbias Vbias.n96 8.00727
R20530 Vbias Vbias.n64 8.00727
R20531 Vbias Vbias.n32 8.00727
R20532 Vbias Vbias.n0 8.00727
R20533 Vbias.n510 Vbias.n509 7.9105
R20534 Vbias.n508 Vbias.n507 7.9105
R20535 Vbias.n506 Vbias.n505 7.9105
R20536 Vbias.n504 Vbias.n503 7.9105
R20537 Vbias.n502 Vbias.n501 7.9105
R20538 Vbias.n500 Vbias.n499 7.9105
R20539 Vbias.n498 Vbias.n497 7.9105
R20540 Vbias.n496 Vbias.n495 7.9105
R20541 Vbias.n494 Vbias.n493 7.9105
R20542 Vbias.n492 Vbias.n491 7.9105
R20543 Vbias.n490 Vbias.n489 7.9105
R20544 Vbias.n488 Vbias.n487 7.9105
R20545 Vbias.n486 Vbias.n485 7.9105
R20546 Vbias.n484 Vbias.n483 7.9105
R20547 Vbias.n482 Vbias.n481 7.9105
R20548 Vbias.n478 Vbias.n477 7.9105
R20549 Vbias.n476 Vbias.n475 7.9105
R20550 Vbias.n474 Vbias.n473 7.9105
R20551 Vbias.n472 Vbias.n471 7.9105
R20552 Vbias.n470 Vbias.n469 7.9105
R20553 Vbias.n468 Vbias.n467 7.9105
R20554 Vbias.n466 Vbias.n465 7.9105
R20555 Vbias.n464 Vbias.n463 7.9105
R20556 Vbias.n462 Vbias.n461 7.9105
R20557 Vbias.n460 Vbias.n459 7.9105
R20558 Vbias.n458 Vbias.n457 7.9105
R20559 Vbias.n456 Vbias.n455 7.9105
R20560 Vbias.n454 Vbias.n453 7.9105
R20561 Vbias.n452 Vbias.n451 7.9105
R20562 Vbias.n450 Vbias.n449 7.9105
R20563 Vbias.n446 Vbias.n445 7.9105
R20564 Vbias.n444 Vbias.n443 7.9105
R20565 Vbias.n442 Vbias.n441 7.9105
R20566 Vbias.n440 Vbias.n439 7.9105
R20567 Vbias.n438 Vbias.n437 7.9105
R20568 Vbias.n436 Vbias.n435 7.9105
R20569 Vbias.n434 Vbias.n433 7.9105
R20570 Vbias.n432 Vbias.n431 7.9105
R20571 Vbias.n430 Vbias.n429 7.9105
R20572 Vbias.n428 Vbias.n427 7.9105
R20573 Vbias.n426 Vbias.n425 7.9105
R20574 Vbias.n424 Vbias.n423 7.9105
R20575 Vbias.n422 Vbias.n421 7.9105
R20576 Vbias.n420 Vbias.n419 7.9105
R20577 Vbias.n418 Vbias.n417 7.9105
R20578 Vbias.n414 Vbias.n413 7.9105
R20579 Vbias.n412 Vbias.n411 7.9105
R20580 Vbias.n410 Vbias.n409 7.9105
R20581 Vbias.n408 Vbias.n407 7.9105
R20582 Vbias.n406 Vbias.n405 7.9105
R20583 Vbias.n404 Vbias.n403 7.9105
R20584 Vbias.n402 Vbias.n401 7.9105
R20585 Vbias.n400 Vbias.n399 7.9105
R20586 Vbias.n398 Vbias.n397 7.9105
R20587 Vbias.n396 Vbias.n395 7.9105
R20588 Vbias.n394 Vbias.n393 7.9105
R20589 Vbias.n392 Vbias.n391 7.9105
R20590 Vbias.n390 Vbias.n389 7.9105
R20591 Vbias.n388 Vbias.n387 7.9105
R20592 Vbias.n386 Vbias.n385 7.9105
R20593 Vbias.n382 Vbias.n381 7.9105
R20594 Vbias.n380 Vbias.n379 7.9105
R20595 Vbias.n378 Vbias.n377 7.9105
R20596 Vbias.n376 Vbias.n375 7.9105
R20597 Vbias.n374 Vbias.n373 7.9105
R20598 Vbias.n372 Vbias.n371 7.9105
R20599 Vbias.n370 Vbias.n369 7.9105
R20600 Vbias.n368 Vbias.n367 7.9105
R20601 Vbias.n366 Vbias.n365 7.9105
R20602 Vbias.n364 Vbias.n363 7.9105
R20603 Vbias.n362 Vbias.n361 7.9105
R20604 Vbias.n360 Vbias.n359 7.9105
R20605 Vbias.n358 Vbias.n357 7.9105
R20606 Vbias.n356 Vbias.n355 7.9105
R20607 Vbias.n354 Vbias.n353 7.9105
R20608 Vbias.n350 Vbias.n349 7.9105
R20609 Vbias.n348 Vbias.n347 7.9105
R20610 Vbias.n346 Vbias.n345 7.9105
R20611 Vbias.n344 Vbias.n343 7.9105
R20612 Vbias.n342 Vbias.n341 7.9105
R20613 Vbias.n340 Vbias.n339 7.9105
R20614 Vbias.n338 Vbias.n337 7.9105
R20615 Vbias.n336 Vbias.n335 7.9105
R20616 Vbias.n334 Vbias.n333 7.9105
R20617 Vbias.n332 Vbias.n331 7.9105
R20618 Vbias.n330 Vbias.n329 7.9105
R20619 Vbias.n328 Vbias.n327 7.9105
R20620 Vbias.n326 Vbias.n325 7.9105
R20621 Vbias.n324 Vbias.n323 7.9105
R20622 Vbias.n322 Vbias.n321 7.9105
R20623 Vbias.n318 Vbias.n317 7.9105
R20624 Vbias.n316 Vbias.n315 7.9105
R20625 Vbias.n314 Vbias.n313 7.9105
R20626 Vbias.n312 Vbias.n311 7.9105
R20627 Vbias.n310 Vbias.n309 7.9105
R20628 Vbias.n308 Vbias.n307 7.9105
R20629 Vbias.n306 Vbias.n305 7.9105
R20630 Vbias.n304 Vbias.n303 7.9105
R20631 Vbias.n302 Vbias.n301 7.9105
R20632 Vbias.n300 Vbias.n299 7.9105
R20633 Vbias.n298 Vbias.n297 7.9105
R20634 Vbias.n296 Vbias.n295 7.9105
R20635 Vbias.n294 Vbias.n293 7.9105
R20636 Vbias.n292 Vbias.n291 7.9105
R20637 Vbias.n290 Vbias.n289 7.9105
R20638 Vbias.n286 Vbias.n285 7.9105
R20639 Vbias.n284 Vbias.n283 7.9105
R20640 Vbias.n282 Vbias.n281 7.9105
R20641 Vbias.n280 Vbias.n279 7.9105
R20642 Vbias.n278 Vbias.n277 7.9105
R20643 Vbias.n276 Vbias.n275 7.9105
R20644 Vbias.n274 Vbias.n273 7.9105
R20645 Vbias.n272 Vbias.n271 7.9105
R20646 Vbias.n270 Vbias.n269 7.9105
R20647 Vbias.n268 Vbias.n267 7.9105
R20648 Vbias.n266 Vbias.n265 7.9105
R20649 Vbias.n264 Vbias.n263 7.9105
R20650 Vbias.n262 Vbias.n261 7.9105
R20651 Vbias.n260 Vbias.n259 7.9105
R20652 Vbias.n258 Vbias.n257 7.9105
R20653 Vbias.n254 Vbias.n253 7.9105
R20654 Vbias.n252 Vbias.n251 7.9105
R20655 Vbias.n250 Vbias.n249 7.9105
R20656 Vbias.n248 Vbias.n247 7.9105
R20657 Vbias.n246 Vbias.n245 7.9105
R20658 Vbias.n244 Vbias.n243 7.9105
R20659 Vbias.n242 Vbias.n241 7.9105
R20660 Vbias.n240 Vbias.n239 7.9105
R20661 Vbias.n238 Vbias.n237 7.9105
R20662 Vbias.n236 Vbias.n235 7.9105
R20663 Vbias.n234 Vbias.n233 7.9105
R20664 Vbias.n232 Vbias.n231 7.9105
R20665 Vbias.n230 Vbias.n229 7.9105
R20666 Vbias.n228 Vbias.n227 7.9105
R20667 Vbias.n226 Vbias.n225 7.9105
R20668 Vbias.n222 Vbias.n221 7.9105
R20669 Vbias.n220 Vbias.n219 7.9105
R20670 Vbias.n218 Vbias.n217 7.9105
R20671 Vbias.n216 Vbias.n215 7.9105
R20672 Vbias.n214 Vbias.n213 7.9105
R20673 Vbias.n212 Vbias.n211 7.9105
R20674 Vbias.n210 Vbias.n209 7.9105
R20675 Vbias.n208 Vbias.n207 7.9105
R20676 Vbias.n206 Vbias.n205 7.9105
R20677 Vbias.n204 Vbias.n203 7.9105
R20678 Vbias.n202 Vbias.n201 7.9105
R20679 Vbias.n200 Vbias.n199 7.9105
R20680 Vbias.n198 Vbias.n197 7.9105
R20681 Vbias.n196 Vbias.n195 7.9105
R20682 Vbias.n194 Vbias.n193 7.9105
R20683 Vbias.n190 Vbias.n189 7.9105
R20684 Vbias.n188 Vbias.n187 7.9105
R20685 Vbias.n186 Vbias.n185 7.9105
R20686 Vbias.n184 Vbias.n183 7.9105
R20687 Vbias.n182 Vbias.n181 7.9105
R20688 Vbias.n180 Vbias.n179 7.9105
R20689 Vbias.n178 Vbias.n177 7.9105
R20690 Vbias.n176 Vbias.n175 7.9105
R20691 Vbias.n174 Vbias.n173 7.9105
R20692 Vbias.n172 Vbias.n171 7.9105
R20693 Vbias.n170 Vbias.n169 7.9105
R20694 Vbias.n168 Vbias.n167 7.9105
R20695 Vbias.n166 Vbias.n165 7.9105
R20696 Vbias.n164 Vbias.n163 7.9105
R20697 Vbias.n162 Vbias.n161 7.9105
R20698 Vbias.n158 Vbias.n157 7.9105
R20699 Vbias.n156 Vbias.n155 7.9105
R20700 Vbias.n154 Vbias.n153 7.9105
R20701 Vbias.n152 Vbias.n151 7.9105
R20702 Vbias.n150 Vbias.n149 7.9105
R20703 Vbias.n148 Vbias.n147 7.9105
R20704 Vbias.n146 Vbias.n145 7.9105
R20705 Vbias.n144 Vbias.n143 7.9105
R20706 Vbias.n142 Vbias.n141 7.9105
R20707 Vbias.n140 Vbias.n139 7.9105
R20708 Vbias.n138 Vbias.n137 7.9105
R20709 Vbias.n136 Vbias.n135 7.9105
R20710 Vbias.n134 Vbias.n133 7.9105
R20711 Vbias.n132 Vbias.n131 7.9105
R20712 Vbias.n130 Vbias.n129 7.9105
R20713 Vbias.n126 Vbias.n125 7.9105
R20714 Vbias.n124 Vbias.n123 7.9105
R20715 Vbias.n122 Vbias.n121 7.9105
R20716 Vbias.n120 Vbias.n119 7.9105
R20717 Vbias.n118 Vbias.n117 7.9105
R20718 Vbias.n116 Vbias.n115 7.9105
R20719 Vbias.n114 Vbias.n113 7.9105
R20720 Vbias.n112 Vbias.n111 7.9105
R20721 Vbias.n110 Vbias.n109 7.9105
R20722 Vbias.n108 Vbias.n107 7.9105
R20723 Vbias.n106 Vbias.n105 7.9105
R20724 Vbias.n104 Vbias.n103 7.9105
R20725 Vbias.n102 Vbias.n101 7.9105
R20726 Vbias.n100 Vbias.n99 7.9105
R20727 Vbias.n98 Vbias.n97 7.9105
R20728 Vbias.n94 Vbias.n93 7.9105
R20729 Vbias.n92 Vbias.n91 7.9105
R20730 Vbias.n90 Vbias.n89 7.9105
R20731 Vbias.n88 Vbias.n87 7.9105
R20732 Vbias.n86 Vbias.n85 7.9105
R20733 Vbias.n84 Vbias.n83 7.9105
R20734 Vbias.n82 Vbias.n81 7.9105
R20735 Vbias.n80 Vbias.n79 7.9105
R20736 Vbias.n78 Vbias.n77 7.9105
R20737 Vbias.n76 Vbias.n75 7.9105
R20738 Vbias.n74 Vbias.n73 7.9105
R20739 Vbias.n72 Vbias.n71 7.9105
R20740 Vbias.n70 Vbias.n69 7.9105
R20741 Vbias.n68 Vbias.n67 7.9105
R20742 Vbias.n66 Vbias.n65 7.9105
R20743 Vbias.n62 Vbias.n61 7.9105
R20744 Vbias.n60 Vbias.n59 7.9105
R20745 Vbias.n58 Vbias.n57 7.9105
R20746 Vbias.n56 Vbias.n55 7.9105
R20747 Vbias.n54 Vbias.n53 7.9105
R20748 Vbias.n52 Vbias.n51 7.9105
R20749 Vbias.n50 Vbias.n49 7.9105
R20750 Vbias.n48 Vbias.n47 7.9105
R20751 Vbias.n46 Vbias.n45 7.9105
R20752 Vbias.n44 Vbias.n43 7.9105
R20753 Vbias.n42 Vbias.n41 7.9105
R20754 Vbias.n40 Vbias.n39 7.9105
R20755 Vbias.n38 Vbias.n37 7.9105
R20756 Vbias.n36 Vbias.n35 7.9105
R20757 Vbias.n34 Vbias.n33 7.9105
R20758 Vbias.n30 Vbias.n29 7.9105
R20759 Vbias.n28 Vbias.n27 7.9105
R20760 Vbias.n26 Vbias.n25 7.9105
R20761 Vbias.n24 Vbias.n23 7.9105
R20762 Vbias.n22 Vbias.n21 7.9105
R20763 Vbias.n20 Vbias.n19 7.9105
R20764 Vbias.n18 Vbias.n17 7.9105
R20765 Vbias.n16 Vbias.n15 7.9105
R20766 Vbias.n14 Vbias.n13 7.9105
R20767 Vbias.n12 Vbias.n11 7.9105
R20768 Vbias.n10 Vbias.n9 7.9105
R20769 Vbias.n8 Vbias.n7 7.9105
R20770 Vbias.n6 Vbias.n5 7.9105
R20771 Vbias.n4 Vbias.n3 7.9105
R20772 Vbias.n2 Vbias.n1 7.9105
R20773 Vbias.n524 Vbias 6.41494
R20774 Vbias.n516 Vbias.n515 2.87046
R20775 Vbias.n522 Vbias.n521 2.87046
R20776 Vbias.n511 Vbias 1.6647
R20777 Vbias.n479 Vbias 1.6647
R20778 Vbias.n447 Vbias 1.6647
R20779 Vbias.n415 Vbias 1.6647
R20780 Vbias.n383 Vbias 1.6647
R20781 Vbias.n351 Vbias 1.6647
R20782 Vbias.n319 Vbias 1.6647
R20783 Vbias.n287 Vbias 1.6647
R20784 Vbias.n255 Vbias 1.6647
R20785 Vbias.n223 Vbias 1.6647
R20786 Vbias.n191 Vbias 1.6647
R20787 Vbias.n159 Vbias 1.6647
R20788 Vbias.n127 Vbias 1.6647
R20789 Vbias.n95 Vbias 1.6647
R20790 Vbias.n63 Vbias 1.6647
R20791 Vbias.n31 Vbias 1.6647
R20792 Vbias.n524 Vbias.n511 0.5692
R20793 Vbias.n63 Vbias.n31 0.410967
R20794 Vbias.n95 Vbias.n63 0.410967
R20795 Vbias.n127 Vbias.n95 0.410967
R20796 Vbias.n159 Vbias.n127 0.410967
R20797 Vbias.n191 Vbias.n159 0.410967
R20798 Vbias.n223 Vbias.n191 0.410967
R20799 Vbias.n255 Vbias.n223 0.410967
R20800 Vbias.n287 Vbias.n255 0.410967
R20801 Vbias.n319 Vbias.n287 0.410967
R20802 Vbias.n351 Vbias.n319 0.410967
R20803 Vbias.n383 Vbias.n351 0.410967
R20804 Vbias.n415 Vbias.n383 0.410967
R20805 Vbias.n447 Vbias.n415 0.410967
R20806 Vbias.n479 Vbias.n447 0.410967
R20807 Vbias.n511 Vbias.n479 0.410967
R20808 Vbias.n31 Vbias 0.383811
R20809 Vbias.n482 Vbias 0.252372
R20810 Vbias.n484 Vbias 0.252372
R20811 Vbias.n486 Vbias 0.252372
R20812 Vbias.n488 Vbias 0.252372
R20813 Vbias.n490 Vbias 0.252372
R20814 Vbias.n492 Vbias 0.252372
R20815 Vbias.n494 Vbias 0.252372
R20816 Vbias.n496 Vbias 0.252372
R20817 Vbias.n498 Vbias 0.252372
R20818 Vbias.n500 Vbias 0.252372
R20819 Vbias.n502 Vbias 0.252372
R20820 Vbias.n504 Vbias 0.252372
R20821 Vbias.n506 Vbias 0.252372
R20822 Vbias.n508 Vbias 0.252372
R20823 Vbias.n510 Vbias 0.252372
R20824 Vbias.n450 Vbias 0.252372
R20825 Vbias.n452 Vbias 0.252372
R20826 Vbias.n454 Vbias 0.252372
R20827 Vbias.n456 Vbias 0.252372
R20828 Vbias.n458 Vbias 0.252372
R20829 Vbias.n460 Vbias 0.252372
R20830 Vbias.n462 Vbias 0.252372
R20831 Vbias.n464 Vbias 0.252372
R20832 Vbias.n466 Vbias 0.252372
R20833 Vbias.n468 Vbias 0.252372
R20834 Vbias.n470 Vbias 0.252372
R20835 Vbias.n472 Vbias 0.252372
R20836 Vbias.n474 Vbias 0.252372
R20837 Vbias.n476 Vbias 0.252372
R20838 Vbias.n478 Vbias 0.252372
R20839 Vbias.n418 Vbias 0.252372
R20840 Vbias.n420 Vbias 0.252372
R20841 Vbias.n422 Vbias 0.252372
R20842 Vbias.n424 Vbias 0.252372
R20843 Vbias.n426 Vbias 0.252372
R20844 Vbias.n428 Vbias 0.252372
R20845 Vbias.n430 Vbias 0.252372
R20846 Vbias.n432 Vbias 0.252372
R20847 Vbias.n434 Vbias 0.252372
R20848 Vbias.n436 Vbias 0.252372
R20849 Vbias.n438 Vbias 0.252372
R20850 Vbias.n440 Vbias 0.252372
R20851 Vbias.n442 Vbias 0.252372
R20852 Vbias.n444 Vbias 0.252372
R20853 Vbias.n446 Vbias 0.252372
R20854 Vbias.n386 Vbias 0.252372
R20855 Vbias.n388 Vbias 0.252372
R20856 Vbias.n390 Vbias 0.252372
R20857 Vbias.n392 Vbias 0.252372
R20858 Vbias.n394 Vbias 0.252372
R20859 Vbias.n396 Vbias 0.252372
R20860 Vbias.n398 Vbias 0.252372
R20861 Vbias.n400 Vbias 0.252372
R20862 Vbias.n402 Vbias 0.252372
R20863 Vbias.n404 Vbias 0.252372
R20864 Vbias.n406 Vbias 0.252372
R20865 Vbias.n408 Vbias 0.252372
R20866 Vbias.n410 Vbias 0.252372
R20867 Vbias.n412 Vbias 0.252372
R20868 Vbias.n414 Vbias 0.252372
R20869 Vbias.n354 Vbias 0.252372
R20870 Vbias.n356 Vbias 0.252372
R20871 Vbias.n358 Vbias 0.252372
R20872 Vbias.n360 Vbias 0.252372
R20873 Vbias.n362 Vbias 0.252372
R20874 Vbias.n364 Vbias 0.252372
R20875 Vbias.n366 Vbias 0.252372
R20876 Vbias.n368 Vbias 0.252372
R20877 Vbias.n370 Vbias 0.252372
R20878 Vbias.n372 Vbias 0.252372
R20879 Vbias.n374 Vbias 0.252372
R20880 Vbias.n376 Vbias 0.252372
R20881 Vbias.n378 Vbias 0.252372
R20882 Vbias.n380 Vbias 0.252372
R20883 Vbias.n382 Vbias 0.252372
R20884 Vbias.n322 Vbias 0.252372
R20885 Vbias.n324 Vbias 0.252372
R20886 Vbias.n326 Vbias 0.252372
R20887 Vbias.n328 Vbias 0.252372
R20888 Vbias.n330 Vbias 0.252372
R20889 Vbias.n332 Vbias 0.252372
R20890 Vbias.n334 Vbias 0.252372
R20891 Vbias.n336 Vbias 0.252372
R20892 Vbias.n338 Vbias 0.252372
R20893 Vbias.n340 Vbias 0.252372
R20894 Vbias.n342 Vbias 0.252372
R20895 Vbias.n344 Vbias 0.252372
R20896 Vbias.n346 Vbias 0.252372
R20897 Vbias.n348 Vbias 0.252372
R20898 Vbias.n350 Vbias 0.252372
R20899 Vbias.n290 Vbias 0.252372
R20900 Vbias.n292 Vbias 0.252372
R20901 Vbias.n294 Vbias 0.252372
R20902 Vbias.n296 Vbias 0.252372
R20903 Vbias.n298 Vbias 0.252372
R20904 Vbias.n300 Vbias 0.252372
R20905 Vbias.n302 Vbias 0.252372
R20906 Vbias.n304 Vbias 0.252372
R20907 Vbias.n306 Vbias 0.252372
R20908 Vbias.n308 Vbias 0.252372
R20909 Vbias.n310 Vbias 0.252372
R20910 Vbias.n312 Vbias 0.252372
R20911 Vbias.n314 Vbias 0.252372
R20912 Vbias.n316 Vbias 0.252372
R20913 Vbias.n318 Vbias 0.252372
R20914 Vbias.n258 Vbias 0.252372
R20915 Vbias.n260 Vbias 0.252372
R20916 Vbias.n262 Vbias 0.252372
R20917 Vbias.n264 Vbias 0.252372
R20918 Vbias.n266 Vbias 0.252372
R20919 Vbias.n268 Vbias 0.252372
R20920 Vbias.n270 Vbias 0.252372
R20921 Vbias.n272 Vbias 0.252372
R20922 Vbias.n274 Vbias 0.252372
R20923 Vbias.n276 Vbias 0.252372
R20924 Vbias.n278 Vbias 0.252372
R20925 Vbias.n280 Vbias 0.252372
R20926 Vbias.n282 Vbias 0.252372
R20927 Vbias.n284 Vbias 0.252372
R20928 Vbias.n286 Vbias 0.252372
R20929 Vbias.n226 Vbias 0.252372
R20930 Vbias.n228 Vbias 0.252372
R20931 Vbias.n230 Vbias 0.252372
R20932 Vbias.n232 Vbias 0.252372
R20933 Vbias.n234 Vbias 0.252372
R20934 Vbias.n236 Vbias 0.252372
R20935 Vbias.n238 Vbias 0.252372
R20936 Vbias.n240 Vbias 0.252372
R20937 Vbias.n242 Vbias 0.252372
R20938 Vbias.n244 Vbias 0.252372
R20939 Vbias.n246 Vbias 0.252372
R20940 Vbias.n248 Vbias 0.252372
R20941 Vbias.n250 Vbias 0.252372
R20942 Vbias.n252 Vbias 0.252372
R20943 Vbias.n254 Vbias 0.252372
R20944 Vbias.n194 Vbias 0.252372
R20945 Vbias.n196 Vbias 0.252372
R20946 Vbias.n198 Vbias 0.252372
R20947 Vbias.n200 Vbias 0.252372
R20948 Vbias.n202 Vbias 0.252372
R20949 Vbias.n204 Vbias 0.252372
R20950 Vbias.n206 Vbias 0.252372
R20951 Vbias.n208 Vbias 0.252372
R20952 Vbias.n210 Vbias 0.252372
R20953 Vbias.n212 Vbias 0.252372
R20954 Vbias.n214 Vbias 0.252372
R20955 Vbias.n216 Vbias 0.252372
R20956 Vbias.n218 Vbias 0.252372
R20957 Vbias.n220 Vbias 0.252372
R20958 Vbias.n222 Vbias 0.252372
R20959 Vbias.n162 Vbias 0.252372
R20960 Vbias.n164 Vbias 0.252372
R20961 Vbias.n166 Vbias 0.252372
R20962 Vbias.n168 Vbias 0.252372
R20963 Vbias.n170 Vbias 0.252372
R20964 Vbias.n172 Vbias 0.252372
R20965 Vbias.n174 Vbias 0.252372
R20966 Vbias.n176 Vbias 0.252372
R20967 Vbias.n178 Vbias 0.252372
R20968 Vbias.n180 Vbias 0.252372
R20969 Vbias.n182 Vbias 0.252372
R20970 Vbias.n184 Vbias 0.252372
R20971 Vbias.n186 Vbias 0.252372
R20972 Vbias.n188 Vbias 0.252372
R20973 Vbias.n190 Vbias 0.252372
R20974 Vbias.n130 Vbias 0.252372
R20975 Vbias.n132 Vbias 0.252372
R20976 Vbias.n134 Vbias 0.252372
R20977 Vbias.n136 Vbias 0.252372
R20978 Vbias.n138 Vbias 0.252372
R20979 Vbias.n140 Vbias 0.252372
R20980 Vbias.n142 Vbias 0.252372
R20981 Vbias.n144 Vbias 0.252372
R20982 Vbias.n146 Vbias 0.252372
R20983 Vbias.n148 Vbias 0.252372
R20984 Vbias.n150 Vbias 0.252372
R20985 Vbias.n152 Vbias 0.252372
R20986 Vbias.n154 Vbias 0.252372
R20987 Vbias.n156 Vbias 0.252372
R20988 Vbias.n158 Vbias 0.252372
R20989 Vbias.n98 Vbias 0.252372
R20990 Vbias.n100 Vbias 0.252372
R20991 Vbias.n102 Vbias 0.252372
R20992 Vbias.n104 Vbias 0.252372
R20993 Vbias.n106 Vbias 0.252372
R20994 Vbias.n108 Vbias 0.252372
R20995 Vbias.n110 Vbias 0.252372
R20996 Vbias.n112 Vbias 0.252372
R20997 Vbias.n114 Vbias 0.252372
R20998 Vbias.n116 Vbias 0.252372
R20999 Vbias.n118 Vbias 0.252372
R21000 Vbias.n120 Vbias 0.252372
R21001 Vbias.n122 Vbias 0.252372
R21002 Vbias.n124 Vbias 0.252372
R21003 Vbias.n126 Vbias 0.252372
R21004 Vbias.n66 Vbias 0.252372
R21005 Vbias.n68 Vbias 0.252372
R21006 Vbias.n70 Vbias 0.252372
R21007 Vbias.n72 Vbias 0.252372
R21008 Vbias.n74 Vbias 0.252372
R21009 Vbias.n76 Vbias 0.252372
R21010 Vbias.n78 Vbias 0.252372
R21011 Vbias.n80 Vbias 0.252372
R21012 Vbias.n82 Vbias 0.252372
R21013 Vbias.n84 Vbias 0.252372
R21014 Vbias.n86 Vbias 0.252372
R21015 Vbias.n88 Vbias 0.252372
R21016 Vbias.n90 Vbias 0.252372
R21017 Vbias.n92 Vbias 0.252372
R21018 Vbias.n94 Vbias 0.252372
R21019 Vbias.n34 Vbias 0.252372
R21020 Vbias.n36 Vbias 0.252372
R21021 Vbias.n38 Vbias 0.252372
R21022 Vbias.n40 Vbias 0.252372
R21023 Vbias.n42 Vbias 0.252372
R21024 Vbias.n44 Vbias 0.252372
R21025 Vbias.n46 Vbias 0.252372
R21026 Vbias.n48 Vbias 0.252372
R21027 Vbias.n50 Vbias 0.252372
R21028 Vbias.n52 Vbias 0.252372
R21029 Vbias.n54 Vbias 0.252372
R21030 Vbias.n56 Vbias 0.252372
R21031 Vbias.n58 Vbias 0.252372
R21032 Vbias.n60 Vbias 0.252372
R21033 Vbias.n62 Vbias 0.252372
R21034 Vbias.n2 Vbias 0.252372
R21035 Vbias.n4 Vbias 0.252372
R21036 Vbias.n6 Vbias 0.252372
R21037 Vbias.n8 Vbias 0.252372
R21038 Vbias.n10 Vbias 0.252372
R21039 Vbias.n12 Vbias 0.252372
R21040 Vbias.n14 Vbias 0.252372
R21041 Vbias.n16 Vbias 0.252372
R21042 Vbias.n18 Vbias 0.252372
R21043 Vbias.n20 Vbias 0.252372
R21044 Vbias.n22 Vbias 0.252372
R21045 Vbias.n24 Vbias 0.252372
R21046 Vbias.n26 Vbias 0.252372
R21047 Vbias.n28 Vbias 0.252372
R21048 Vbias.n30 Vbias 0.252372
R21049 Vbias Vbias.n524 0.237067
R21050 Vbias.n517 Vbias.n512 0.215542
R21051 Vbias.n523 Vbias.n518 0.215542
R21052 Vbias Vbias.n517 0.175939
R21053 Vbias.n517 Vbias.n516 0.150018
R21054 Vbias.n523 Vbias.n522 0.150018
R21055 Vbias Vbias.n523 0.127693
R21056 Vbias Vbias.n482 0.0972718
R21057 Vbias Vbias.n484 0.0972718
R21058 Vbias Vbias.n486 0.0972718
R21059 Vbias Vbias.n488 0.0972718
R21060 Vbias Vbias.n490 0.0972718
R21061 Vbias Vbias.n492 0.0972718
R21062 Vbias Vbias.n494 0.0972718
R21063 Vbias Vbias.n496 0.0972718
R21064 Vbias Vbias.n498 0.0972718
R21065 Vbias Vbias.n500 0.0972718
R21066 Vbias Vbias.n502 0.0972718
R21067 Vbias Vbias.n504 0.0972718
R21068 Vbias Vbias.n506 0.0972718
R21069 Vbias Vbias.n508 0.0972718
R21070 Vbias Vbias.n510 0.0972718
R21071 Vbias Vbias.n450 0.0972718
R21072 Vbias Vbias.n452 0.0972718
R21073 Vbias Vbias.n454 0.0972718
R21074 Vbias Vbias.n456 0.0972718
R21075 Vbias Vbias.n458 0.0972718
R21076 Vbias Vbias.n460 0.0972718
R21077 Vbias Vbias.n462 0.0972718
R21078 Vbias Vbias.n464 0.0972718
R21079 Vbias Vbias.n466 0.0972718
R21080 Vbias Vbias.n468 0.0972718
R21081 Vbias Vbias.n470 0.0972718
R21082 Vbias Vbias.n472 0.0972718
R21083 Vbias Vbias.n474 0.0972718
R21084 Vbias Vbias.n476 0.0972718
R21085 Vbias Vbias.n478 0.0972718
R21086 Vbias Vbias.n418 0.0972718
R21087 Vbias Vbias.n420 0.0972718
R21088 Vbias Vbias.n422 0.0972718
R21089 Vbias Vbias.n424 0.0972718
R21090 Vbias Vbias.n426 0.0972718
R21091 Vbias Vbias.n428 0.0972718
R21092 Vbias Vbias.n430 0.0972718
R21093 Vbias Vbias.n432 0.0972718
R21094 Vbias Vbias.n434 0.0972718
R21095 Vbias Vbias.n436 0.0972718
R21096 Vbias Vbias.n438 0.0972718
R21097 Vbias Vbias.n440 0.0972718
R21098 Vbias Vbias.n442 0.0972718
R21099 Vbias Vbias.n444 0.0972718
R21100 Vbias Vbias.n446 0.0972718
R21101 Vbias Vbias.n386 0.0972718
R21102 Vbias Vbias.n388 0.0972718
R21103 Vbias Vbias.n390 0.0972718
R21104 Vbias Vbias.n392 0.0972718
R21105 Vbias Vbias.n394 0.0972718
R21106 Vbias Vbias.n396 0.0972718
R21107 Vbias Vbias.n398 0.0972718
R21108 Vbias Vbias.n400 0.0972718
R21109 Vbias Vbias.n402 0.0972718
R21110 Vbias Vbias.n404 0.0972718
R21111 Vbias Vbias.n406 0.0972718
R21112 Vbias Vbias.n408 0.0972718
R21113 Vbias Vbias.n410 0.0972718
R21114 Vbias Vbias.n412 0.0972718
R21115 Vbias Vbias.n414 0.0972718
R21116 Vbias Vbias.n354 0.0972718
R21117 Vbias Vbias.n356 0.0972718
R21118 Vbias Vbias.n358 0.0972718
R21119 Vbias Vbias.n360 0.0972718
R21120 Vbias Vbias.n362 0.0972718
R21121 Vbias Vbias.n364 0.0972718
R21122 Vbias Vbias.n366 0.0972718
R21123 Vbias Vbias.n368 0.0972718
R21124 Vbias Vbias.n370 0.0972718
R21125 Vbias Vbias.n372 0.0972718
R21126 Vbias Vbias.n374 0.0972718
R21127 Vbias Vbias.n376 0.0972718
R21128 Vbias Vbias.n378 0.0972718
R21129 Vbias Vbias.n380 0.0972718
R21130 Vbias Vbias.n382 0.0972718
R21131 Vbias Vbias.n322 0.0972718
R21132 Vbias Vbias.n324 0.0972718
R21133 Vbias Vbias.n326 0.0972718
R21134 Vbias Vbias.n328 0.0972718
R21135 Vbias Vbias.n330 0.0972718
R21136 Vbias Vbias.n332 0.0972718
R21137 Vbias Vbias.n334 0.0972718
R21138 Vbias Vbias.n336 0.0972718
R21139 Vbias Vbias.n338 0.0972718
R21140 Vbias Vbias.n340 0.0972718
R21141 Vbias Vbias.n342 0.0972718
R21142 Vbias Vbias.n344 0.0972718
R21143 Vbias Vbias.n346 0.0972718
R21144 Vbias Vbias.n348 0.0972718
R21145 Vbias Vbias.n350 0.0972718
R21146 Vbias Vbias.n290 0.0972718
R21147 Vbias Vbias.n292 0.0972718
R21148 Vbias Vbias.n294 0.0972718
R21149 Vbias Vbias.n296 0.0972718
R21150 Vbias Vbias.n298 0.0972718
R21151 Vbias Vbias.n300 0.0972718
R21152 Vbias Vbias.n302 0.0972718
R21153 Vbias Vbias.n304 0.0972718
R21154 Vbias Vbias.n306 0.0972718
R21155 Vbias Vbias.n308 0.0972718
R21156 Vbias Vbias.n310 0.0972718
R21157 Vbias Vbias.n312 0.0972718
R21158 Vbias Vbias.n314 0.0972718
R21159 Vbias Vbias.n316 0.0972718
R21160 Vbias Vbias.n318 0.0972718
R21161 Vbias Vbias.n258 0.0972718
R21162 Vbias Vbias.n260 0.0972718
R21163 Vbias Vbias.n262 0.0972718
R21164 Vbias Vbias.n264 0.0972718
R21165 Vbias Vbias.n266 0.0972718
R21166 Vbias Vbias.n268 0.0972718
R21167 Vbias Vbias.n270 0.0972718
R21168 Vbias Vbias.n272 0.0972718
R21169 Vbias Vbias.n274 0.0972718
R21170 Vbias Vbias.n276 0.0972718
R21171 Vbias Vbias.n278 0.0972718
R21172 Vbias Vbias.n280 0.0972718
R21173 Vbias Vbias.n282 0.0972718
R21174 Vbias Vbias.n284 0.0972718
R21175 Vbias Vbias.n286 0.0972718
R21176 Vbias Vbias.n226 0.0972718
R21177 Vbias Vbias.n228 0.0972718
R21178 Vbias Vbias.n230 0.0972718
R21179 Vbias Vbias.n232 0.0972718
R21180 Vbias Vbias.n234 0.0972718
R21181 Vbias Vbias.n236 0.0972718
R21182 Vbias Vbias.n238 0.0972718
R21183 Vbias Vbias.n240 0.0972718
R21184 Vbias Vbias.n242 0.0972718
R21185 Vbias Vbias.n244 0.0972718
R21186 Vbias Vbias.n246 0.0972718
R21187 Vbias Vbias.n248 0.0972718
R21188 Vbias Vbias.n250 0.0972718
R21189 Vbias Vbias.n252 0.0972718
R21190 Vbias Vbias.n254 0.0972718
R21191 Vbias Vbias.n194 0.0972718
R21192 Vbias Vbias.n196 0.0972718
R21193 Vbias Vbias.n198 0.0972718
R21194 Vbias Vbias.n200 0.0972718
R21195 Vbias Vbias.n202 0.0972718
R21196 Vbias Vbias.n204 0.0972718
R21197 Vbias Vbias.n206 0.0972718
R21198 Vbias Vbias.n208 0.0972718
R21199 Vbias Vbias.n210 0.0972718
R21200 Vbias Vbias.n212 0.0972718
R21201 Vbias Vbias.n214 0.0972718
R21202 Vbias Vbias.n216 0.0972718
R21203 Vbias Vbias.n218 0.0972718
R21204 Vbias Vbias.n220 0.0972718
R21205 Vbias Vbias.n222 0.0972718
R21206 Vbias Vbias.n162 0.0972718
R21207 Vbias Vbias.n164 0.0972718
R21208 Vbias Vbias.n166 0.0972718
R21209 Vbias Vbias.n168 0.0972718
R21210 Vbias Vbias.n170 0.0972718
R21211 Vbias Vbias.n172 0.0972718
R21212 Vbias Vbias.n174 0.0972718
R21213 Vbias Vbias.n176 0.0972718
R21214 Vbias Vbias.n178 0.0972718
R21215 Vbias Vbias.n180 0.0972718
R21216 Vbias Vbias.n182 0.0972718
R21217 Vbias Vbias.n184 0.0972718
R21218 Vbias Vbias.n186 0.0972718
R21219 Vbias Vbias.n188 0.0972718
R21220 Vbias Vbias.n190 0.0972718
R21221 Vbias Vbias.n130 0.0972718
R21222 Vbias Vbias.n132 0.0972718
R21223 Vbias Vbias.n134 0.0972718
R21224 Vbias Vbias.n136 0.0972718
R21225 Vbias Vbias.n138 0.0972718
R21226 Vbias Vbias.n140 0.0972718
R21227 Vbias Vbias.n142 0.0972718
R21228 Vbias Vbias.n144 0.0972718
R21229 Vbias Vbias.n146 0.0972718
R21230 Vbias Vbias.n148 0.0972718
R21231 Vbias Vbias.n150 0.0972718
R21232 Vbias Vbias.n152 0.0972718
R21233 Vbias Vbias.n154 0.0972718
R21234 Vbias Vbias.n156 0.0972718
R21235 Vbias Vbias.n158 0.0972718
R21236 Vbias Vbias.n98 0.0972718
R21237 Vbias Vbias.n100 0.0972718
R21238 Vbias Vbias.n102 0.0972718
R21239 Vbias Vbias.n104 0.0972718
R21240 Vbias Vbias.n106 0.0972718
R21241 Vbias Vbias.n108 0.0972718
R21242 Vbias Vbias.n110 0.0972718
R21243 Vbias Vbias.n112 0.0972718
R21244 Vbias Vbias.n114 0.0972718
R21245 Vbias Vbias.n116 0.0972718
R21246 Vbias Vbias.n118 0.0972718
R21247 Vbias Vbias.n120 0.0972718
R21248 Vbias Vbias.n122 0.0972718
R21249 Vbias Vbias.n124 0.0972718
R21250 Vbias Vbias.n126 0.0972718
R21251 Vbias Vbias.n66 0.0972718
R21252 Vbias Vbias.n68 0.0972718
R21253 Vbias Vbias.n70 0.0972718
R21254 Vbias Vbias.n72 0.0972718
R21255 Vbias Vbias.n74 0.0972718
R21256 Vbias Vbias.n76 0.0972718
R21257 Vbias Vbias.n78 0.0972718
R21258 Vbias Vbias.n80 0.0972718
R21259 Vbias Vbias.n82 0.0972718
R21260 Vbias Vbias.n84 0.0972718
R21261 Vbias Vbias.n86 0.0972718
R21262 Vbias Vbias.n88 0.0972718
R21263 Vbias Vbias.n90 0.0972718
R21264 Vbias Vbias.n92 0.0972718
R21265 Vbias Vbias.n94 0.0972718
R21266 Vbias Vbias.n34 0.0972718
R21267 Vbias Vbias.n36 0.0972718
R21268 Vbias Vbias.n38 0.0972718
R21269 Vbias Vbias.n40 0.0972718
R21270 Vbias Vbias.n42 0.0972718
R21271 Vbias Vbias.n44 0.0972718
R21272 Vbias Vbias.n46 0.0972718
R21273 Vbias Vbias.n48 0.0972718
R21274 Vbias Vbias.n50 0.0972718
R21275 Vbias Vbias.n52 0.0972718
R21276 Vbias Vbias.n54 0.0972718
R21277 Vbias Vbias.n56 0.0972718
R21278 Vbias Vbias.n58 0.0972718
R21279 Vbias Vbias.n60 0.0972718
R21280 Vbias Vbias.n62 0.0972718
R21281 Vbias Vbias.n2 0.0972718
R21282 Vbias Vbias.n4 0.0972718
R21283 Vbias Vbias.n6 0.0972718
R21284 Vbias Vbias.n8 0.0972718
R21285 Vbias Vbias.n10 0.0972718
R21286 Vbias Vbias.n12 0.0972718
R21287 Vbias Vbias.n14 0.0972718
R21288 Vbias Vbias.n16 0.0972718
R21289 Vbias Vbias.n18 0.0972718
R21290 Vbias Vbias.n20 0.0972718
R21291 Vbias Vbias.n22 0.0972718
R21292 Vbias Vbias.n24 0.0972718
R21293 Vbias Vbias.n26 0.0972718
R21294 Vbias Vbias.n28 0.0972718
R21295 Vbias Vbias.n30 0.0972718
R21296 Vbias.n509 Vbias 0.0489375
R21297 Vbias.n507 Vbias 0.0489375
R21298 Vbias.n505 Vbias 0.0489375
R21299 Vbias.n503 Vbias 0.0489375
R21300 Vbias.n501 Vbias 0.0489375
R21301 Vbias.n499 Vbias 0.0489375
R21302 Vbias.n497 Vbias 0.0489375
R21303 Vbias.n495 Vbias 0.0489375
R21304 Vbias.n493 Vbias 0.0489375
R21305 Vbias.n491 Vbias 0.0489375
R21306 Vbias.n489 Vbias 0.0489375
R21307 Vbias.n487 Vbias 0.0489375
R21308 Vbias.n485 Vbias 0.0489375
R21309 Vbias.n483 Vbias 0.0489375
R21310 Vbias.n481 Vbias 0.0489375
R21311 Vbias.n480 Vbias 0.0489375
R21312 Vbias.n477 Vbias 0.0489375
R21313 Vbias.n475 Vbias 0.0489375
R21314 Vbias.n473 Vbias 0.0489375
R21315 Vbias.n471 Vbias 0.0489375
R21316 Vbias.n469 Vbias 0.0489375
R21317 Vbias.n467 Vbias 0.0489375
R21318 Vbias.n465 Vbias 0.0489375
R21319 Vbias.n463 Vbias 0.0489375
R21320 Vbias.n461 Vbias 0.0489375
R21321 Vbias.n459 Vbias 0.0489375
R21322 Vbias.n457 Vbias 0.0489375
R21323 Vbias.n455 Vbias 0.0489375
R21324 Vbias.n453 Vbias 0.0489375
R21325 Vbias.n451 Vbias 0.0489375
R21326 Vbias.n449 Vbias 0.0489375
R21327 Vbias.n448 Vbias 0.0489375
R21328 Vbias.n445 Vbias 0.0489375
R21329 Vbias.n443 Vbias 0.0489375
R21330 Vbias.n441 Vbias 0.0489375
R21331 Vbias.n439 Vbias 0.0489375
R21332 Vbias.n437 Vbias 0.0489375
R21333 Vbias.n435 Vbias 0.0489375
R21334 Vbias.n433 Vbias 0.0489375
R21335 Vbias.n431 Vbias 0.0489375
R21336 Vbias.n429 Vbias 0.0489375
R21337 Vbias.n427 Vbias 0.0489375
R21338 Vbias.n425 Vbias 0.0489375
R21339 Vbias.n423 Vbias 0.0489375
R21340 Vbias.n421 Vbias 0.0489375
R21341 Vbias.n419 Vbias 0.0489375
R21342 Vbias.n417 Vbias 0.0489375
R21343 Vbias.n416 Vbias 0.0489375
R21344 Vbias.n413 Vbias 0.0489375
R21345 Vbias.n411 Vbias 0.0489375
R21346 Vbias.n409 Vbias 0.0489375
R21347 Vbias.n407 Vbias 0.0489375
R21348 Vbias.n405 Vbias 0.0489375
R21349 Vbias.n403 Vbias 0.0489375
R21350 Vbias.n401 Vbias 0.0489375
R21351 Vbias.n399 Vbias 0.0489375
R21352 Vbias.n397 Vbias 0.0489375
R21353 Vbias.n395 Vbias 0.0489375
R21354 Vbias.n393 Vbias 0.0489375
R21355 Vbias.n391 Vbias 0.0489375
R21356 Vbias.n389 Vbias 0.0489375
R21357 Vbias.n387 Vbias 0.0489375
R21358 Vbias.n385 Vbias 0.0489375
R21359 Vbias.n384 Vbias 0.0489375
R21360 Vbias.n381 Vbias 0.0489375
R21361 Vbias.n379 Vbias 0.0489375
R21362 Vbias.n377 Vbias 0.0489375
R21363 Vbias.n375 Vbias 0.0489375
R21364 Vbias.n373 Vbias 0.0489375
R21365 Vbias.n371 Vbias 0.0489375
R21366 Vbias.n369 Vbias 0.0489375
R21367 Vbias.n367 Vbias 0.0489375
R21368 Vbias.n365 Vbias 0.0489375
R21369 Vbias.n363 Vbias 0.0489375
R21370 Vbias.n361 Vbias 0.0489375
R21371 Vbias.n359 Vbias 0.0489375
R21372 Vbias.n357 Vbias 0.0489375
R21373 Vbias.n355 Vbias 0.0489375
R21374 Vbias.n353 Vbias 0.0489375
R21375 Vbias.n352 Vbias 0.0489375
R21376 Vbias.n349 Vbias 0.0489375
R21377 Vbias.n347 Vbias 0.0489375
R21378 Vbias.n345 Vbias 0.0489375
R21379 Vbias.n343 Vbias 0.0489375
R21380 Vbias.n341 Vbias 0.0489375
R21381 Vbias.n339 Vbias 0.0489375
R21382 Vbias.n337 Vbias 0.0489375
R21383 Vbias.n335 Vbias 0.0489375
R21384 Vbias.n333 Vbias 0.0489375
R21385 Vbias.n331 Vbias 0.0489375
R21386 Vbias.n329 Vbias 0.0489375
R21387 Vbias.n327 Vbias 0.0489375
R21388 Vbias.n325 Vbias 0.0489375
R21389 Vbias.n323 Vbias 0.0489375
R21390 Vbias.n321 Vbias 0.0489375
R21391 Vbias.n320 Vbias 0.0489375
R21392 Vbias.n317 Vbias 0.0489375
R21393 Vbias.n315 Vbias 0.0489375
R21394 Vbias.n313 Vbias 0.0489375
R21395 Vbias.n311 Vbias 0.0489375
R21396 Vbias.n309 Vbias 0.0489375
R21397 Vbias.n307 Vbias 0.0489375
R21398 Vbias.n305 Vbias 0.0489375
R21399 Vbias.n303 Vbias 0.0489375
R21400 Vbias.n301 Vbias 0.0489375
R21401 Vbias.n299 Vbias 0.0489375
R21402 Vbias.n297 Vbias 0.0489375
R21403 Vbias.n295 Vbias 0.0489375
R21404 Vbias.n293 Vbias 0.0489375
R21405 Vbias.n291 Vbias 0.0489375
R21406 Vbias.n289 Vbias 0.0489375
R21407 Vbias.n288 Vbias 0.0489375
R21408 Vbias.n285 Vbias 0.0489375
R21409 Vbias.n283 Vbias 0.0489375
R21410 Vbias.n281 Vbias 0.0489375
R21411 Vbias.n279 Vbias 0.0489375
R21412 Vbias.n277 Vbias 0.0489375
R21413 Vbias.n275 Vbias 0.0489375
R21414 Vbias.n273 Vbias 0.0489375
R21415 Vbias.n271 Vbias 0.0489375
R21416 Vbias.n269 Vbias 0.0489375
R21417 Vbias.n267 Vbias 0.0489375
R21418 Vbias.n265 Vbias 0.0489375
R21419 Vbias.n263 Vbias 0.0489375
R21420 Vbias.n261 Vbias 0.0489375
R21421 Vbias.n259 Vbias 0.0489375
R21422 Vbias.n257 Vbias 0.0489375
R21423 Vbias.n256 Vbias 0.0489375
R21424 Vbias.n253 Vbias 0.0489375
R21425 Vbias.n251 Vbias 0.0489375
R21426 Vbias.n249 Vbias 0.0489375
R21427 Vbias.n247 Vbias 0.0489375
R21428 Vbias.n245 Vbias 0.0489375
R21429 Vbias.n243 Vbias 0.0489375
R21430 Vbias.n241 Vbias 0.0489375
R21431 Vbias.n239 Vbias 0.0489375
R21432 Vbias.n237 Vbias 0.0489375
R21433 Vbias.n235 Vbias 0.0489375
R21434 Vbias.n233 Vbias 0.0489375
R21435 Vbias.n231 Vbias 0.0489375
R21436 Vbias.n229 Vbias 0.0489375
R21437 Vbias.n227 Vbias 0.0489375
R21438 Vbias.n225 Vbias 0.0489375
R21439 Vbias.n224 Vbias 0.0489375
R21440 Vbias.n221 Vbias 0.0489375
R21441 Vbias.n219 Vbias 0.0489375
R21442 Vbias.n217 Vbias 0.0489375
R21443 Vbias.n215 Vbias 0.0489375
R21444 Vbias.n213 Vbias 0.0489375
R21445 Vbias.n211 Vbias 0.0489375
R21446 Vbias.n209 Vbias 0.0489375
R21447 Vbias.n207 Vbias 0.0489375
R21448 Vbias.n205 Vbias 0.0489375
R21449 Vbias.n203 Vbias 0.0489375
R21450 Vbias.n201 Vbias 0.0489375
R21451 Vbias.n199 Vbias 0.0489375
R21452 Vbias.n197 Vbias 0.0489375
R21453 Vbias.n195 Vbias 0.0489375
R21454 Vbias.n193 Vbias 0.0489375
R21455 Vbias.n192 Vbias 0.0489375
R21456 Vbias.n189 Vbias 0.0489375
R21457 Vbias.n187 Vbias 0.0489375
R21458 Vbias.n185 Vbias 0.0489375
R21459 Vbias.n183 Vbias 0.0489375
R21460 Vbias.n181 Vbias 0.0489375
R21461 Vbias.n179 Vbias 0.0489375
R21462 Vbias.n177 Vbias 0.0489375
R21463 Vbias.n175 Vbias 0.0489375
R21464 Vbias.n173 Vbias 0.0489375
R21465 Vbias.n171 Vbias 0.0489375
R21466 Vbias.n169 Vbias 0.0489375
R21467 Vbias.n167 Vbias 0.0489375
R21468 Vbias.n165 Vbias 0.0489375
R21469 Vbias.n163 Vbias 0.0489375
R21470 Vbias.n161 Vbias 0.0489375
R21471 Vbias.n160 Vbias 0.0489375
R21472 Vbias.n157 Vbias 0.0489375
R21473 Vbias.n155 Vbias 0.0489375
R21474 Vbias.n153 Vbias 0.0489375
R21475 Vbias.n151 Vbias 0.0489375
R21476 Vbias.n149 Vbias 0.0489375
R21477 Vbias.n147 Vbias 0.0489375
R21478 Vbias.n145 Vbias 0.0489375
R21479 Vbias.n143 Vbias 0.0489375
R21480 Vbias.n141 Vbias 0.0489375
R21481 Vbias.n139 Vbias 0.0489375
R21482 Vbias.n137 Vbias 0.0489375
R21483 Vbias.n135 Vbias 0.0489375
R21484 Vbias.n133 Vbias 0.0489375
R21485 Vbias.n131 Vbias 0.0489375
R21486 Vbias.n129 Vbias 0.0489375
R21487 Vbias.n128 Vbias 0.0489375
R21488 Vbias.n125 Vbias 0.0489375
R21489 Vbias.n123 Vbias 0.0489375
R21490 Vbias.n121 Vbias 0.0489375
R21491 Vbias.n119 Vbias 0.0489375
R21492 Vbias.n117 Vbias 0.0489375
R21493 Vbias.n115 Vbias 0.0489375
R21494 Vbias.n113 Vbias 0.0489375
R21495 Vbias.n111 Vbias 0.0489375
R21496 Vbias.n109 Vbias 0.0489375
R21497 Vbias.n107 Vbias 0.0489375
R21498 Vbias.n105 Vbias 0.0489375
R21499 Vbias.n103 Vbias 0.0489375
R21500 Vbias.n101 Vbias 0.0489375
R21501 Vbias.n99 Vbias 0.0489375
R21502 Vbias.n97 Vbias 0.0489375
R21503 Vbias.n96 Vbias 0.0489375
R21504 Vbias.n93 Vbias 0.0489375
R21505 Vbias.n91 Vbias 0.0489375
R21506 Vbias.n89 Vbias 0.0489375
R21507 Vbias.n87 Vbias 0.0489375
R21508 Vbias.n85 Vbias 0.0489375
R21509 Vbias.n83 Vbias 0.0489375
R21510 Vbias.n81 Vbias 0.0489375
R21511 Vbias.n79 Vbias 0.0489375
R21512 Vbias.n77 Vbias 0.0489375
R21513 Vbias.n75 Vbias 0.0489375
R21514 Vbias.n73 Vbias 0.0489375
R21515 Vbias.n71 Vbias 0.0489375
R21516 Vbias.n69 Vbias 0.0489375
R21517 Vbias.n67 Vbias 0.0489375
R21518 Vbias.n65 Vbias 0.0489375
R21519 Vbias.n64 Vbias 0.0489375
R21520 Vbias.n61 Vbias 0.0489375
R21521 Vbias.n59 Vbias 0.0489375
R21522 Vbias.n57 Vbias 0.0489375
R21523 Vbias.n55 Vbias 0.0489375
R21524 Vbias.n53 Vbias 0.0489375
R21525 Vbias.n51 Vbias 0.0489375
R21526 Vbias.n49 Vbias 0.0489375
R21527 Vbias.n47 Vbias 0.0489375
R21528 Vbias.n45 Vbias 0.0489375
R21529 Vbias.n43 Vbias 0.0489375
R21530 Vbias.n41 Vbias 0.0489375
R21531 Vbias.n39 Vbias 0.0489375
R21532 Vbias.n37 Vbias 0.0489375
R21533 Vbias.n35 Vbias 0.0489375
R21534 Vbias.n33 Vbias 0.0489375
R21535 Vbias.n32 Vbias 0.0489375
R21536 Vbias.n29 Vbias 0.0489375
R21537 Vbias.n27 Vbias 0.0489375
R21538 Vbias.n25 Vbias 0.0489375
R21539 Vbias.n23 Vbias 0.0489375
R21540 Vbias.n21 Vbias 0.0489375
R21541 Vbias.n19 Vbias 0.0489375
R21542 Vbias.n17 Vbias 0.0489375
R21543 Vbias.n15 Vbias 0.0489375
R21544 Vbias.n13 Vbias 0.0489375
R21545 Vbias.n11 Vbias 0.0489375
R21546 Vbias.n9 Vbias 0.0489375
R21547 Vbias.n7 Vbias 0.0489375
R21548 Vbias.n5 Vbias 0.0489375
R21549 Vbias.n3 Vbias 0.0489375
R21550 Vbias.n1 Vbias 0.0489375
R21551 Vbias.n0 Vbias 0.0489375
R21552 XThC.Tn[1].n2 XThC.Tn[1].n1 332.332
R21553 XThC.Tn[1].n2 XThC.Tn[1].n0 296.493
R21554 XThC.Tn[1].n12 XThC.Tn[1].n10 161.406
R21555 XThC.Tn[1].n15 XThC.Tn[1].n13 161.406
R21556 XThC.Tn[1].n18 XThC.Tn[1].n16 161.406
R21557 XThC.Tn[1].n21 XThC.Tn[1].n19 161.406
R21558 XThC.Tn[1].n24 XThC.Tn[1].n22 161.406
R21559 XThC.Tn[1].n27 XThC.Tn[1].n25 161.406
R21560 XThC.Tn[1].n30 XThC.Tn[1].n28 161.406
R21561 XThC.Tn[1].n33 XThC.Tn[1].n31 161.406
R21562 XThC.Tn[1].n36 XThC.Tn[1].n34 161.406
R21563 XThC.Tn[1].n39 XThC.Tn[1].n37 161.406
R21564 XThC.Tn[1].n42 XThC.Tn[1].n40 161.406
R21565 XThC.Tn[1].n45 XThC.Tn[1].n43 161.406
R21566 XThC.Tn[1].n48 XThC.Tn[1].n46 161.406
R21567 XThC.Tn[1].n51 XThC.Tn[1].n49 161.406
R21568 XThC.Tn[1].n54 XThC.Tn[1].n52 161.406
R21569 XThC.Tn[1].n57 XThC.Tn[1].n55 161.406
R21570 XThC.Tn[1].n10 XThC.Tn[1].t29 161.202
R21571 XThC.Tn[1].n13 XThC.Tn[1].t14 161.202
R21572 XThC.Tn[1].n16 XThC.Tn[1].t16 161.202
R21573 XThC.Tn[1].n19 XThC.Tn[1].t18 161.202
R21574 XThC.Tn[1].n22 XThC.Tn[1].t39 161.202
R21575 XThC.Tn[1].n25 XThC.Tn[1].t40 161.202
R21576 XThC.Tn[1].n28 XThC.Tn[1].t21 161.202
R21577 XThC.Tn[1].n31 XThC.Tn[1].t30 161.202
R21578 XThC.Tn[1].n34 XThC.Tn[1].t32 161.202
R21579 XThC.Tn[1].n37 XThC.Tn[1].t19 161.202
R21580 XThC.Tn[1].n40 XThC.Tn[1].t20 161.202
R21581 XThC.Tn[1].n43 XThC.Tn[1].t33 161.202
R21582 XThC.Tn[1].n46 XThC.Tn[1].t41 161.202
R21583 XThC.Tn[1].n49 XThC.Tn[1].t12 161.202
R21584 XThC.Tn[1].n52 XThC.Tn[1].t25 161.202
R21585 XThC.Tn[1].n55 XThC.Tn[1].t35 161.202
R21586 XThC.Tn[1].n10 XThC.Tn[1].t31 145.137
R21587 XThC.Tn[1].n13 XThC.Tn[1].t17 145.137
R21588 XThC.Tn[1].n16 XThC.Tn[1].t22 145.137
R21589 XThC.Tn[1].n19 XThC.Tn[1].t23 145.137
R21590 XThC.Tn[1].n22 XThC.Tn[1].t42 145.137
R21591 XThC.Tn[1].n25 XThC.Tn[1].t43 145.137
R21592 XThC.Tn[1].n28 XThC.Tn[1].t27 145.137
R21593 XThC.Tn[1].n31 XThC.Tn[1].t34 145.137
R21594 XThC.Tn[1].n34 XThC.Tn[1].t36 145.137
R21595 XThC.Tn[1].n37 XThC.Tn[1].t24 145.137
R21596 XThC.Tn[1].n40 XThC.Tn[1].t26 145.137
R21597 XThC.Tn[1].n43 XThC.Tn[1].t37 145.137
R21598 XThC.Tn[1].n46 XThC.Tn[1].t13 145.137
R21599 XThC.Tn[1].n49 XThC.Tn[1].t15 145.137
R21600 XThC.Tn[1].n52 XThC.Tn[1].t28 145.137
R21601 XThC.Tn[1].n55 XThC.Tn[1].t38 145.137
R21602 XThC.Tn[1].n7 XThC.Tn[1].n6 135.249
R21603 XThC.Tn[1].n9 XThC.Tn[1].n3 98.981
R21604 XThC.Tn[1].n8 XThC.Tn[1].n4 98.981
R21605 XThC.Tn[1].n7 XThC.Tn[1].n5 98.981
R21606 XThC.Tn[1].n9 XThC.Tn[1].n8 36.2672
R21607 XThC.Tn[1].n8 XThC.Tn[1].n7 36.2672
R21608 XThC.Tn[1].n59 XThC.Tn[1].n9 32.6405
R21609 XThC.Tn[1].n1 XThC.Tn[1].t9 26.5955
R21610 XThC.Tn[1].n1 XThC.Tn[1].t8 26.5955
R21611 XThC.Tn[1].n0 XThC.Tn[1].t11 26.5955
R21612 XThC.Tn[1].n0 XThC.Tn[1].t10 26.5955
R21613 XThC.Tn[1].n3 XThC.Tn[1].t5 24.9236
R21614 XThC.Tn[1].n3 XThC.Tn[1].t4 24.9236
R21615 XThC.Tn[1].n4 XThC.Tn[1].t7 24.9236
R21616 XThC.Tn[1].n4 XThC.Tn[1].t6 24.9236
R21617 XThC.Tn[1].n5 XThC.Tn[1].t1 24.9236
R21618 XThC.Tn[1].n5 XThC.Tn[1].t0 24.9236
R21619 XThC.Tn[1].n6 XThC.Tn[1].t3 24.9236
R21620 XThC.Tn[1].n6 XThC.Tn[1].t2 24.9236
R21621 XThC.Tn[1] XThC.Tn[1].n2 23.3605
R21622 XThC.Tn[1].n58 XThC.Tn[1] 7.29217
R21623 XThC.Tn[1] XThC.Tn[1].n59 6.7205
R21624 XThC.Tn[1].n59 XThC.Tn[1].n58 3.13711
R21625 XThC.Tn[1].n15 XThC.Tn[1] 0.931056
R21626 XThC.Tn[1].n18 XThC.Tn[1] 0.931056
R21627 XThC.Tn[1].n21 XThC.Tn[1] 0.931056
R21628 XThC.Tn[1].n24 XThC.Tn[1] 0.931056
R21629 XThC.Tn[1].n27 XThC.Tn[1] 0.931056
R21630 XThC.Tn[1].n30 XThC.Tn[1] 0.931056
R21631 XThC.Tn[1].n33 XThC.Tn[1] 0.931056
R21632 XThC.Tn[1].n36 XThC.Tn[1] 0.931056
R21633 XThC.Tn[1].n39 XThC.Tn[1] 0.931056
R21634 XThC.Tn[1].n42 XThC.Tn[1] 0.931056
R21635 XThC.Tn[1].n45 XThC.Tn[1] 0.931056
R21636 XThC.Tn[1].n48 XThC.Tn[1] 0.931056
R21637 XThC.Tn[1].n51 XThC.Tn[1] 0.931056
R21638 XThC.Tn[1].n54 XThC.Tn[1] 0.931056
R21639 XThC.Tn[1].n57 XThC.Tn[1] 0.931056
R21640 XThC.Tn[1] XThC.Tn[1].n12 0.396333
R21641 XThC.Tn[1] XThC.Tn[1].n15 0.396333
R21642 XThC.Tn[1] XThC.Tn[1].n18 0.396333
R21643 XThC.Tn[1] XThC.Tn[1].n21 0.396333
R21644 XThC.Tn[1] XThC.Tn[1].n24 0.396333
R21645 XThC.Tn[1] XThC.Tn[1].n27 0.396333
R21646 XThC.Tn[1] XThC.Tn[1].n30 0.396333
R21647 XThC.Tn[1] XThC.Tn[1].n33 0.396333
R21648 XThC.Tn[1] XThC.Tn[1].n36 0.396333
R21649 XThC.Tn[1] XThC.Tn[1].n39 0.396333
R21650 XThC.Tn[1] XThC.Tn[1].n42 0.396333
R21651 XThC.Tn[1] XThC.Tn[1].n45 0.396333
R21652 XThC.Tn[1] XThC.Tn[1].n48 0.396333
R21653 XThC.Tn[1] XThC.Tn[1].n51 0.396333
R21654 XThC.Tn[1] XThC.Tn[1].n54 0.396333
R21655 XThC.Tn[1] XThC.Tn[1].n57 0.396333
R21656 XThC.Tn[1].n11 XThC.Tn[1] 0.104667
R21657 XThC.Tn[1].n14 XThC.Tn[1] 0.104667
R21658 XThC.Tn[1].n17 XThC.Tn[1] 0.104667
R21659 XThC.Tn[1].n20 XThC.Tn[1] 0.104667
R21660 XThC.Tn[1].n23 XThC.Tn[1] 0.104667
R21661 XThC.Tn[1].n26 XThC.Tn[1] 0.104667
R21662 XThC.Tn[1].n29 XThC.Tn[1] 0.104667
R21663 XThC.Tn[1].n32 XThC.Tn[1] 0.104667
R21664 XThC.Tn[1].n35 XThC.Tn[1] 0.104667
R21665 XThC.Tn[1].n38 XThC.Tn[1] 0.104667
R21666 XThC.Tn[1].n41 XThC.Tn[1] 0.104667
R21667 XThC.Tn[1].n44 XThC.Tn[1] 0.104667
R21668 XThC.Tn[1].n47 XThC.Tn[1] 0.104667
R21669 XThC.Tn[1].n50 XThC.Tn[1] 0.104667
R21670 XThC.Tn[1].n53 XThC.Tn[1] 0.104667
R21671 XThC.Tn[1].n56 XThC.Tn[1] 0.104667
R21672 XThC.Tn[1].n58 XThC.Tn[1] 0.0594286
R21673 XThC.Tn[1].n11 XThC.Tn[1] 0.0309878
R21674 XThC.Tn[1].n14 XThC.Tn[1] 0.0309878
R21675 XThC.Tn[1].n17 XThC.Tn[1] 0.0309878
R21676 XThC.Tn[1].n20 XThC.Tn[1] 0.0309878
R21677 XThC.Tn[1].n23 XThC.Tn[1] 0.0309878
R21678 XThC.Tn[1].n26 XThC.Tn[1] 0.0309878
R21679 XThC.Tn[1].n29 XThC.Tn[1] 0.0309878
R21680 XThC.Tn[1].n32 XThC.Tn[1] 0.0309878
R21681 XThC.Tn[1].n35 XThC.Tn[1] 0.0309878
R21682 XThC.Tn[1].n38 XThC.Tn[1] 0.0309878
R21683 XThC.Tn[1].n41 XThC.Tn[1] 0.0309878
R21684 XThC.Tn[1].n44 XThC.Tn[1] 0.0309878
R21685 XThC.Tn[1].n47 XThC.Tn[1] 0.0309878
R21686 XThC.Tn[1].n50 XThC.Tn[1] 0.0309878
R21687 XThC.Tn[1].n53 XThC.Tn[1] 0.0309878
R21688 XThC.Tn[1].n56 XThC.Tn[1] 0.0309878
R21689 XThC.Tn[1].n12 XThC.Tn[1].n11 0.027939
R21690 XThC.Tn[1].n15 XThC.Tn[1].n14 0.027939
R21691 XThC.Tn[1].n18 XThC.Tn[1].n17 0.027939
R21692 XThC.Tn[1].n21 XThC.Tn[1].n20 0.027939
R21693 XThC.Tn[1].n24 XThC.Tn[1].n23 0.027939
R21694 XThC.Tn[1].n27 XThC.Tn[1].n26 0.027939
R21695 XThC.Tn[1].n30 XThC.Tn[1].n29 0.027939
R21696 XThC.Tn[1].n33 XThC.Tn[1].n32 0.027939
R21697 XThC.Tn[1].n36 XThC.Tn[1].n35 0.027939
R21698 XThC.Tn[1].n39 XThC.Tn[1].n38 0.027939
R21699 XThC.Tn[1].n42 XThC.Tn[1].n41 0.027939
R21700 XThC.Tn[1].n45 XThC.Tn[1].n44 0.027939
R21701 XThC.Tn[1].n48 XThC.Tn[1].n47 0.027939
R21702 XThC.Tn[1].n51 XThC.Tn[1].n50 0.027939
R21703 XThC.Tn[1].n54 XThC.Tn[1].n53 0.027939
R21704 XThC.Tn[1].n57 XThC.Tn[1].n56 0.027939
R21705 XThC.Tn[3].n2 XThC.Tn[3].n1 332.332
R21706 XThC.Tn[3].n2 XThC.Tn[3].n0 296.493
R21707 XThC.Tn[3].n12 XThC.Tn[3].n10 161.406
R21708 XThC.Tn[3].n15 XThC.Tn[3].n13 161.406
R21709 XThC.Tn[3].n18 XThC.Tn[3].n16 161.406
R21710 XThC.Tn[3].n21 XThC.Tn[3].n19 161.406
R21711 XThC.Tn[3].n24 XThC.Tn[3].n22 161.406
R21712 XThC.Tn[3].n27 XThC.Tn[3].n25 161.406
R21713 XThC.Tn[3].n30 XThC.Tn[3].n28 161.406
R21714 XThC.Tn[3].n33 XThC.Tn[3].n31 161.406
R21715 XThC.Tn[3].n36 XThC.Tn[3].n34 161.406
R21716 XThC.Tn[3].n39 XThC.Tn[3].n37 161.406
R21717 XThC.Tn[3].n42 XThC.Tn[3].n40 161.406
R21718 XThC.Tn[3].n45 XThC.Tn[3].n43 161.406
R21719 XThC.Tn[3].n48 XThC.Tn[3].n46 161.406
R21720 XThC.Tn[3].n51 XThC.Tn[3].n49 161.406
R21721 XThC.Tn[3].n54 XThC.Tn[3].n52 161.406
R21722 XThC.Tn[3].n57 XThC.Tn[3].n55 161.406
R21723 XThC.Tn[3].n10 XThC.Tn[3].t42 161.202
R21724 XThC.Tn[3].n13 XThC.Tn[3].t27 161.202
R21725 XThC.Tn[3].n16 XThC.Tn[3].t29 161.202
R21726 XThC.Tn[3].n19 XThC.Tn[3].t31 161.202
R21727 XThC.Tn[3].n22 XThC.Tn[3].t20 161.202
R21728 XThC.Tn[3].n25 XThC.Tn[3].t21 161.202
R21729 XThC.Tn[3].n28 XThC.Tn[3].t34 161.202
R21730 XThC.Tn[3].n31 XThC.Tn[3].t43 161.202
R21731 XThC.Tn[3].n34 XThC.Tn[3].t13 161.202
R21732 XThC.Tn[3].n37 XThC.Tn[3].t32 161.202
R21733 XThC.Tn[3].n40 XThC.Tn[3].t33 161.202
R21734 XThC.Tn[3].n43 XThC.Tn[3].t14 161.202
R21735 XThC.Tn[3].n46 XThC.Tn[3].t22 161.202
R21736 XThC.Tn[3].n49 XThC.Tn[3].t25 161.202
R21737 XThC.Tn[3].n52 XThC.Tn[3].t38 161.202
R21738 XThC.Tn[3].n55 XThC.Tn[3].t16 161.202
R21739 XThC.Tn[3].n10 XThC.Tn[3].t12 145.137
R21740 XThC.Tn[3].n13 XThC.Tn[3].t30 145.137
R21741 XThC.Tn[3].n16 XThC.Tn[3].t35 145.137
R21742 XThC.Tn[3].n19 XThC.Tn[3].t36 145.137
R21743 XThC.Tn[3].n22 XThC.Tn[3].t23 145.137
R21744 XThC.Tn[3].n25 XThC.Tn[3].t24 145.137
R21745 XThC.Tn[3].n28 XThC.Tn[3].t40 145.137
R21746 XThC.Tn[3].n31 XThC.Tn[3].t15 145.137
R21747 XThC.Tn[3].n34 XThC.Tn[3].t17 145.137
R21748 XThC.Tn[3].n37 XThC.Tn[3].t37 145.137
R21749 XThC.Tn[3].n40 XThC.Tn[3].t39 145.137
R21750 XThC.Tn[3].n43 XThC.Tn[3].t18 145.137
R21751 XThC.Tn[3].n46 XThC.Tn[3].t26 145.137
R21752 XThC.Tn[3].n49 XThC.Tn[3].t28 145.137
R21753 XThC.Tn[3].n52 XThC.Tn[3].t41 145.137
R21754 XThC.Tn[3].n55 XThC.Tn[3].t19 145.137
R21755 XThC.Tn[3].n6 XThC.Tn[3].n4 135.249
R21756 XThC.Tn[3].n9 XThC.Tn[3].n3 98.981
R21757 XThC.Tn[3].n6 XThC.Tn[3].n5 98.981
R21758 XThC.Tn[3].n8 XThC.Tn[3].n7 98.981
R21759 XThC.Tn[3].n8 XThC.Tn[3].n6 36.2672
R21760 XThC.Tn[3].n9 XThC.Tn[3].n8 36.2672
R21761 XThC.Tn[3].n58 XThC.Tn[3].n9 32.6405
R21762 XThC.Tn[3].n1 XThC.Tn[3].t7 26.5955
R21763 XThC.Tn[3].n1 XThC.Tn[3].t6 26.5955
R21764 XThC.Tn[3].n0 XThC.Tn[3].t5 26.5955
R21765 XThC.Tn[3].n0 XThC.Tn[3].t4 26.5955
R21766 XThC.Tn[3].n3 XThC.Tn[3].t1 24.9236
R21767 XThC.Tn[3].n3 XThC.Tn[3].t0 24.9236
R21768 XThC.Tn[3].n4 XThC.Tn[3].t11 24.9236
R21769 XThC.Tn[3].n4 XThC.Tn[3].t10 24.9236
R21770 XThC.Tn[3].n5 XThC.Tn[3].t9 24.9236
R21771 XThC.Tn[3].n5 XThC.Tn[3].t8 24.9236
R21772 XThC.Tn[3].n7 XThC.Tn[3].t3 24.9236
R21773 XThC.Tn[3].n7 XThC.Tn[3].t2 24.9236
R21774 XThC.Tn[3] XThC.Tn[3].n2 23.3605
R21775 XThC.Tn[3] XThC.Tn[3].n58 6.7205
R21776 XThC.Tn[3].n58 XThC.Tn[3] 3.19574
R21777 XThC.Tn[3].n15 XThC.Tn[3] 0.931056
R21778 XThC.Tn[3].n18 XThC.Tn[3] 0.931056
R21779 XThC.Tn[3].n21 XThC.Tn[3] 0.931056
R21780 XThC.Tn[3].n24 XThC.Tn[3] 0.931056
R21781 XThC.Tn[3].n27 XThC.Tn[3] 0.931056
R21782 XThC.Tn[3].n30 XThC.Tn[3] 0.931056
R21783 XThC.Tn[3].n33 XThC.Tn[3] 0.931056
R21784 XThC.Tn[3].n36 XThC.Tn[3] 0.931056
R21785 XThC.Tn[3].n39 XThC.Tn[3] 0.931056
R21786 XThC.Tn[3].n42 XThC.Tn[3] 0.931056
R21787 XThC.Tn[3].n45 XThC.Tn[3] 0.931056
R21788 XThC.Tn[3].n48 XThC.Tn[3] 0.931056
R21789 XThC.Tn[3].n51 XThC.Tn[3] 0.931056
R21790 XThC.Tn[3].n54 XThC.Tn[3] 0.931056
R21791 XThC.Tn[3].n57 XThC.Tn[3] 0.931056
R21792 XThC.Tn[3] XThC.Tn[3].n12 0.396333
R21793 XThC.Tn[3] XThC.Tn[3].n15 0.396333
R21794 XThC.Tn[3] XThC.Tn[3].n18 0.396333
R21795 XThC.Tn[3] XThC.Tn[3].n21 0.396333
R21796 XThC.Tn[3] XThC.Tn[3].n24 0.396333
R21797 XThC.Tn[3] XThC.Tn[3].n27 0.396333
R21798 XThC.Tn[3] XThC.Tn[3].n30 0.396333
R21799 XThC.Tn[3] XThC.Tn[3].n33 0.396333
R21800 XThC.Tn[3] XThC.Tn[3].n36 0.396333
R21801 XThC.Tn[3] XThC.Tn[3].n39 0.396333
R21802 XThC.Tn[3] XThC.Tn[3].n42 0.396333
R21803 XThC.Tn[3] XThC.Tn[3].n45 0.396333
R21804 XThC.Tn[3] XThC.Tn[3].n48 0.396333
R21805 XThC.Tn[3] XThC.Tn[3].n51 0.396333
R21806 XThC.Tn[3] XThC.Tn[3].n54 0.396333
R21807 XThC.Tn[3] XThC.Tn[3].n57 0.396333
R21808 XThC.Tn[3].n11 XThC.Tn[3] 0.104667
R21809 XThC.Tn[3].n14 XThC.Tn[3] 0.104667
R21810 XThC.Tn[3].n17 XThC.Tn[3] 0.104667
R21811 XThC.Tn[3].n20 XThC.Tn[3] 0.104667
R21812 XThC.Tn[3].n23 XThC.Tn[3] 0.104667
R21813 XThC.Tn[3].n26 XThC.Tn[3] 0.104667
R21814 XThC.Tn[3].n29 XThC.Tn[3] 0.104667
R21815 XThC.Tn[3].n32 XThC.Tn[3] 0.104667
R21816 XThC.Tn[3].n35 XThC.Tn[3] 0.104667
R21817 XThC.Tn[3].n38 XThC.Tn[3] 0.104667
R21818 XThC.Tn[3].n41 XThC.Tn[3] 0.104667
R21819 XThC.Tn[3].n44 XThC.Tn[3] 0.104667
R21820 XThC.Tn[3].n47 XThC.Tn[3] 0.104667
R21821 XThC.Tn[3].n50 XThC.Tn[3] 0.104667
R21822 XThC.Tn[3].n53 XThC.Tn[3] 0.104667
R21823 XThC.Tn[3].n56 XThC.Tn[3] 0.104667
R21824 XThC.Tn[3].n11 XThC.Tn[3] 0.0309878
R21825 XThC.Tn[3].n14 XThC.Tn[3] 0.0309878
R21826 XThC.Tn[3].n17 XThC.Tn[3] 0.0309878
R21827 XThC.Tn[3].n20 XThC.Tn[3] 0.0309878
R21828 XThC.Tn[3].n23 XThC.Tn[3] 0.0309878
R21829 XThC.Tn[3].n26 XThC.Tn[3] 0.0309878
R21830 XThC.Tn[3].n29 XThC.Tn[3] 0.0309878
R21831 XThC.Tn[3].n32 XThC.Tn[3] 0.0309878
R21832 XThC.Tn[3].n35 XThC.Tn[3] 0.0309878
R21833 XThC.Tn[3].n38 XThC.Tn[3] 0.0309878
R21834 XThC.Tn[3].n41 XThC.Tn[3] 0.0309878
R21835 XThC.Tn[3].n44 XThC.Tn[3] 0.0309878
R21836 XThC.Tn[3].n47 XThC.Tn[3] 0.0309878
R21837 XThC.Tn[3].n50 XThC.Tn[3] 0.0309878
R21838 XThC.Tn[3].n53 XThC.Tn[3] 0.0309878
R21839 XThC.Tn[3].n56 XThC.Tn[3] 0.0309878
R21840 XThC.Tn[3].n12 XThC.Tn[3].n11 0.027939
R21841 XThC.Tn[3].n15 XThC.Tn[3].n14 0.027939
R21842 XThC.Tn[3].n18 XThC.Tn[3].n17 0.027939
R21843 XThC.Tn[3].n21 XThC.Tn[3].n20 0.027939
R21844 XThC.Tn[3].n24 XThC.Tn[3].n23 0.027939
R21845 XThC.Tn[3].n27 XThC.Tn[3].n26 0.027939
R21846 XThC.Tn[3].n30 XThC.Tn[3].n29 0.027939
R21847 XThC.Tn[3].n33 XThC.Tn[3].n32 0.027939
R21848 XThC.Tn[3].n36 XThC.Tn[3].n35 0.027939
R21849 XThC.Tn[3].n39 XThC.Tn[3].n38 0.027939
R21850 XThC.Tn[3].n42 XThC.Tn[3].n41 0.027939
R21851 XThC.Tn[3].n45 XThC.Tn[3].n44 0.027939
R21852 XThC.Tn[3].n48 XThC.Tn[3].n47 0.027939
R21853 XThC.Tn[3].n51 XThC.Tn[3].n50 0.027939
R21854 XThC.Tn[3].n54 XThC.Tn[3].n53 0.027939
R21855 XThC.Tn[3].n57 XThC.Tn[3].n56 0.027939
R21856 XThR.Tn[10].n5 XThR.Tn[10].n4 256.103
R21857 XThR.Tn[10].n2 XThR.Tn[10].n0 243.68
R21858 XThR.Tn[10].n88 XThR.Tn[10].n86 241.847
R21859 XThR.Tn[10].n2 XThR.Tn[10].n1 205.28
R21860 XThR.Tn[10].n5 XThR.Tn[10].n3 202.095
R21861 XThR.Tn[10].n88 XThR.Tn[10].n87 185
R21862 XThR.Tn[10] XThR.Tn[10].n79 161.363
R21863 XThR.Tn[10] XThR.Tn[10].n74 161.363
R21864 XThR.Tn[10] XThR.Tn[10].n69 161.363
R21865 XThR.Tn[10] XThR.Tn[10].n64 161.363
R21866 XThR.Tn[10] XThR.Tn[10].n59 161.363
R21867 XThR.Tn[10] XThR.Tn[10].n54 161.363
R21868 XThR.Tn[10] XThR.Tn[10].n49 161.363
R21869 XThR.Tn[10] XThR.Tn[10].n44 161.363
R21870 XThR.Tn[10] XThR.Tn[10].n39 161.363
R21871 XThR.Tn[10] XThR.Tn[10].n34 161.363
R21872 XThR.Tn[10] XThR.Tn[10].n29 161.363
R21873 XThR.Tn[10] XThR.Tn[10].n24 161.363
R21874 XThR.Tn[10] XThR.Tn[10].n19 161.363
R21875 XThR.Tn[10] XThR.Tn[10].n14 161.363
R21876 XThR.Tn[10] XThR.Tn[10].n9 161.363
R21877 XThR.Tn[10] XThR.Tn[10].n7 161.363
R21878 XThR.Tn[10].n81 XThR.Tn[10].n80 161.3
R21879 XThR.Tn[10].n76 XThR.Tn[10].n75 161.3
R21880 XThR.Tn[10].n71 XThR.Tn[10].n70 161.3
R21881 XThR.Tn[10].n66 XThR.Tn[10].n65 161.3
R21882 XThR.Tn[10].n61 XThR.Tn[10].n60 161.3
R21883 XThR.Tn[10].n56 XThR.Tn[10].n55 161.3
R21884 XThR.Tn[10].n51 XThR.Tn[10].n50 161.3
R21885 XThR.Tn[10].n46 XThR.Tn[10].n45 161.3
R21886 XThR.Tn[10].n41 XThR.Tn[10].n40 161.3
R21887 XThR.Tn[10].n36 XThR.Tn[10].n35 161.3
R21888 XThR.Tn[10].n31 XThR.Tn[10].n30 161.3
R21889 XThR.Tn[10].n26 XThR.Tn[10].n25 161.3
R21890 XThR.Tn[10].n21 XThR.Tn[10].n20 161.3
R21891 XThR.Tn[10].n16 XThR.Tn[10].n15 161.3
R21892 XThR.Tn[10].n11 XThR.Tn[10].n10 161.3
R21893 XThR.Tn[10].n79 XThR.Tn[10].t37 161.106
R21894 XThR.Tn[10].n74 XThR.Tn[10].t45 161.106
R21895 XThR.Tn[10].n69 XThR.Tn[10].t27 161.106
R21896 XThR.Tn[10].n64 XThR.Tn[10].t72 161.106
R21897 XThR.Tn[10].n59 XThR.Tn[10].t35 161.106
R21898 XThR.Tn[10].n54 XThR.Tn[10].t61 161.106
R21899 XThR.Tn[10].n49 XThR.Tn[10].t43 161.106
R21900 XThR.Tn[10].n44 XThR.Tn[10].t24 161.106
R21901 XThR.Tn[10].n39 XThR.Tn[10].t69 161.106
R21902 XThR.Tn[10].n34 XThR.Tn[10].t15 161.106
R21903 XThR.Tn[10].n29 XThR.Tn[10].t59 161.106
R21904 XThR.Tn[10].n24 XThR.Tn[10].t26 161.106
R21905 XThR.Tn[10].n19 XThR.Tn[10].t58 161.106
R21906 XThR.Tn[10].n14 XThR.Tn[10].t41 161.106
R21907 XThR.Tn[10].n9 XThR.Tn[10].t63 161.106
R21908 XThR.Tn[10].n7 XThR.Tn[10].t47 161.106
R21909 XThR.Tn[10].n80 XThR.Tn[10].t34 159.978
R21910 XThR.Tn[10].n75 XThR.Tn[10].t39 159.978
R21911 XThR.Tn[10].n70 XThR.Tn[10].t22 159.978
R21912 XThR.Tn[10].n65 XThR.Tn[10].t68 159.978
R21913 XThR.Tn[10].n60 XThR.Tn[10].t32 159.978
R21914 XThR.Tn[10].n55 XThR.Tn[10].t57 159.978
R21915 XThR.Tn[10].n50 XThR.Tn[10].t38 159.978
R21916 XThR.Tn[10].n45 XThR.Tn[10].t20 159.978
R21917 XThR.Tn[10].n40 XThR.Tn[10].t66 159.978
R21918 XThR.Tn[10].n35 XThR.Tn[10].t12 159.978
R21919 XThR.Tn[10].n30 XThR.Tn[10].t56 159.978
R21920 XThR.Tn[10].n25 XThR.Tn[10].t21 159.978
R21921 XThR.Tn[10].n20 XThR.Tn[10].t55 159.978
R21922 XThR.Tn[10].n15 XThR.Tn[10].t36 159.978
R21923 XThR.Tn[10].n10 XThR.Tn[10].t60 159.978
R21924 XThR.Tn[10].n79 XThR.Tn[10].t29 145.038
R21925 XThR.Tn[10].n74 XThR.Tn[10].t49 145.038
R21926 XThR.Tn[10].n69 XThR.Tn[10].t31 145.038
R21927 XThR.Tn[10].n64 XThR.Tn[10].t16 145.038
R21928 XThR.Tn[10].n59 XThR.Tn[10].t46 145.038
R21929 XThR.Tn[10].n54 XThR.Tn[10].t28 145.038
R21930 XThR.Tn[10].n49 XThR.Tn[10].t33 145.038
R21931 XThR.Tn[10].n44 XThR.Tn[10].t17 145.038
R21932 XThR.Tn[10].n39 XThR.Tn[10].t14 145.038
R21933 XThR.Tn[10].n34 XThR.Tn[10].t44 145.038
R21934 XThR.Tn[10].n29 XThR.Tn[10].t67 145.038
R21935 XThR.Tn[10].n24 XThR.Tn[10].t30 145.038
R21936 XThR.Tn[10].n19 XThR.Tn[10].t65 145.038
R21937 XThR.Tn[10].n14 XThR.Tn[10].t48 145.038
R21938 XThR.Tn[10].n9 XThR.Tn[10].t13 145.038
R21939 XThR.Tn[10].n7 XThR.Tn[10].t54 145.038
R21940 XThR.Tn[10].n80 XThR.Tn[10].t64 143.911
R21941 XThR.Tn[10].n75 XThR.Tn[10].t25 143.911
R21942 XThR.Tn[10].n70 XThR.Tn[10].t71 143.911
R21943 XThR.Tn[10].n65 XThR.Tn[10].t52 143.911
R21944 XThR.Tn[10].n60 XThR.Tn[10].t19 143.911
R21945 XThR.Tn[10].n55 XThR.Tn[10].t62 143.911
R21946 XThR.Tn[10].n50 XThR.Tn[10].t73 143.911
R21947 XThR.Tn[10].n45 XThR.Tn[10].t53 143.911
R21948 XThR.Tn[10].n40 XThR.Tn[10].t51 143.911
R21949 XThR.Tn[10].n35 XThR.Tn[10].t18 143.911
R21950 XThR.Tn[10].n30 XThR.Tn[10].t42 143.911
R21951 XThR.Tn[10].n25 XThR.Tn[10].t70 143.911
R21952 XThR.Tn[10].n20 XThR.Tn[10].t40 143.911
R21953 XThR.Tn[10].n15 XThR.Tn[10].t23 143.911
R21954 XThR.Tn[10].n10 XThR.Tn[10].t50 143.911
R21955 XThR.Tn[10] XThR.Tn[10].n2 35.7652
R21956 XThR.Tn[10].n3 XThR.Tn[10].t6 26.5955
R21957 XThR.Tn[10].n3 XThR.Tn[10].t10 26.5955
R21958 XThR.Tn[10].n4 XThR.Tn[10].t7 26.5955
R21959 XThR.Tn[10].n4 XThR.Tn[10].t9 26.5955
R21960 XThR.Tn[10].n0 XThR.Tn[10].t4 26.5955
R21961 XThR.Tn[10].n0 XThR.Tn[10].t2 26.5955
R21962 XThR.Tn[10].n1 XThR.Tn[10].t5 26.5955
R21963 XThR.Tn[10].n1 XThR.Tn[10].t3 26.5955
R21964 XThR.Tn[10].n86 XThR.Tn[10].t11 24.9236
R21965 XThR.Tn[10].n86 XThR.Tn[10].t1 24.9236
R21966 XThR.Tn[10].n87 XThR.Tn[10].t0 24.9236
R21967 XThR.Tn[10].n87 XThR.Tn[10].t8 24.9236
R21968 XThR.Tn[10] XThR.Tn[10].n88 18.8943
R21969 XThR.Tn[10].n6 XThR.Tn[10].n5 13.5534
R21970 XThR.Tn[10].n85 XThR.Tn[10] 7.84567
R21971 XThR.Tn[10] XThR.Tn[10].n85 6.34069
R21972 XThR.Tn[10] XThR.Tn[10].n8 5.34038
R21973 XThR.Tn[10].n13 XThR.Tn[10].n12 4.5005
R21974 XThR.Tn[10].n18 XThR.Tn[10].n17 4.5005
R21975 XThR.Tn[10].n23 XThR.Tn[10].n22 4.5005
R21976 XThR.Tn[10].n28 XThR.Tn[10].n27 4.5005
R21977 XThR.Tn[10].n33 XThR.Tn[10].n32 4.5005
R21978 XThR.Tn[10].n38 XThR.Tn[10].n37 4.5005
R21979 XThR.Tn[10].n43 XThR.Tn[10].n42 4.5005
R21980 XThR.Tn[10].n48 XThR.Tn[10].n47 4.5005
R21981 XThR.Tn[10].n53 XThR.Tn[10].n52 4.5005
R21982 XThR.Tn[10].n58 XThR.Tn[10].n57 4.5005
R21983 XThR.Tn[10].n63 XThR.Tn[10].n62 4.5005
R21984 XThR.Tn[10].n68 XThR.Tn[10].n67 4.5005
R21985 XThR.Tn[10].n73 XThR.Tn[10].n72 4.5005
R21986 XThR.Tn[10].n78 XThR.Tn[10].n77 4.5005
R21987 XThR.Tn[10].n83 XThR.Tn[10].n82 4.5005
R21988 XThR.Tn[10].n84 XThR.Tn[10] 3.70586
R21989 XThR.Tn[10].n13 XThR.Tn[10] 2.52282
R21990 XThR.Tn[10].n18 XThR.Tn[10] 2.52282
R21991 XThR.Tn[10].n23 XThR.Tn[10] 2.52282
R21992 XThR.Tn[10].n28 XThR.Tn[10] 2.52282
R21993 XThR.Tn[10].n33 XThR.Tn[10] 2.52282
R21994 XThR.Tn[10].n38 XThR.Tn[10] 2.52282
R21995 XThR.Tn[10].n43 XThR.Tn[10] 2.52282
R21996 XThR.Tn[10].n48 XThR.Tn[10] 2.52282
R21997 XThR.Tn[10].n53 XThR.Tn[10] 2.52282
R21998 XThR.Tn[10].n58 XThR.Tn[10] 2.52282
R21999 XThR.Tn[10].n63 XThR.Tn[10] 2.52282
R22000 XThR.Tn[10].n68 XThR.Tn[10] 2.52282
R22001 XThR.Tn[10].n73 XThR.Tn[10] 2.52282
R22002 XThR.Tn[10].n78 XThR.Tn[10] 2.52282
R22003 XThR.Tn[10].n83 XThR.Tn[10] 2.52282
R22004 XThR.Tn[10].n85 XThR.Tn[10] 1.79489
R22005 XThR.Tn[10].n6 XThR.Tn[10] 1.50638
R22006 XThR.Tn[10] XThR.Tn[10].n6 1.19676
R22007 XThR.Tn[10].n81 XThR.Tn[10] 1.08677
R22008 XThR.Tn[10].n76 XThR.Tn[10] 1.08677
R22009 XThR.Tn[10].n71 XThR.Tn[10] 1.08677
R22010 XThR.Tn[10].n66 XThR.Tn[10] 1.08677
R22011 XThR.Tn[10].n61 XThR.Tn[10] 1.08677
R22012 XThR.Tn[10].n56 XThR.Tn[10] 1.08677
R22013 XThR.Tn[10].n51 XThR.Tn[10] 1.08677
R22014 XThR.Tn[10].n46 XThR.Tn[10] 1.08677
R22015 XThR.Tn[10].n41 XThR.Tn[10] 1.08677
R22016 XThR.Tn[10].n36 XThR.Tn[10] 1.08677
R22017 XThR.Tn[10].n31 XThR.Tn[10] 1.08677
R22018 XThR.Tn[10].n26 XThR.Tn[10] 1.08677
R22019 XThR.Tn[10].n21 XThR.Tn[10] 1.08677
R22020 XThR.Tn[10].n16 XThR.Tn[10] 1.08677
R22021 XThR.Tn[10].n11 XThR.Tn[10] 1.08677
R22022 XThR.Tn[10] XThR.Tn[10].n13 0.839786
R22023 XThR.Tn[10] XThR.Tn[10].n18 0.839786
R22024 XThR.Tn[10] XThR.Tn[10].n23 0.839786
R22025 XThR.Tn[10] XThR.Tn[10].n28 0.839786
R22026 XThR.Tn[10] XThR.Tn[10].n33 0.839786
R22027 XThR.Tn[10] XThR.Tn[10].n38 0.839786
R22028 XThR.Tn[10] XThR.Tn[10].n43 0.839786
R22029 XThR.Tn[10] XThR.Tn[10].n48 0.839786
R22030 XThR.Tn[10] XThR.Tn[10].n53 0.839786
R22031 XThR.Tn[10] XThR.Tn[10].n58 0.839786
R22032 XThR.Tn[10] XThR.Tn[10].n63 0.839786
R22033 XThR.Tn[10] XThR.Tn[10].n68 0.839786
R22034 XThR.Tn[10] XThR.Tn[10].n73 0.839786
R22035 XThR.Tn[10] XThR.Tn[10].n78 0.839786
R22036 XThR.Tn[10] XThR.Tn[10].n83 0.839786
R22037 XThR.Tn[10].n8 XThR.Tn[10] 0.499542
R22038 XThR.Tn[10].n82 XThR.Tn[10] 0.063
R22039 XThR.Tn[10].n77 XThR.Tn[10] 0.063
R22040 XThR.Tn[10].n72 XThR.Tn[10] 0.063
R22041 XThR.Tn[10].n67 XThR.Tn[10] 0.063
R22042 XThR.Tn[10].n62 XThR.Tn[10] 0.063
R22043 XThR.Tn[10].n57 XThR.Tn[10] 0.063
R22044 XThR.Tn[10].n52 XThR.Tn[10] 0.063
R22045 XThR.Tn[10].n47 XThR.Tn[10] 0.063
R22046 XThR.Tn[10].n42 XThR.Tn[10] 0.063
R22047 XThR.Tn[10].n37 XThR.Tn[10] 0.063
R22048 XThR.Tn[10].n32 XThR.Tn[10] 0.063
R22049 XThR.Tn[10].n27 XThR.Tn[10] 0.063
R22050 XThR.Tn[10].n22 XThR.Tn[10] 0.063
R22051 XThR.Tn[10].n17 XThR.Tn[10] 0.063
R22052 XThR.Tn[10].n12 XThR.Tn[10] 0.063
R22053 XThR.Tn[10].n84 XThR.Tn[10] 0.0540714
R22054 XThR.Tn[10] XThR.Tn[10].n84 0.038
R22055 XThR.Tn[10].n8 XThR.Tn[10] 0.0143889
R22056 XThR.Tn[10].n82 XThR.Tn[10].n81 0.00771154
R22057 XThR.Tn[10].n77 XThR.Tn[10].n76 0.00771154
R22058 XThR.Tn[10].n72 XThR.Tn[10].n71 0.00771154
R22059 XThR.Tn[10].n67 XThR.Tn[10].n66 0.00771154
R22060 XThR.Tn[10].n62 XThR.Tn[10].n61 0.00771154
R22061 XThR.Tn[10].n57 XThR.Tn[10].n56 0.00771154
R22062 XThR.Tn[10].n52 XThR.Tn[10].n51 0.00771154
R22063 XThR.Tn[10].n47 XThR.Tn[10].n46 0.00771154
R22064 XThR.Tn[10].n42 XThR.Tn[10].n41 0.00771154
R22065 XThR.Tn[10].n37 XThR.Tn[10].n36 0.00771154
R22066 XThR.Tn[10].n32 XThR.Tn[10].n31 0.00771154
R22067 XThR.Tn[10].n27 XThR.Tn[10].n26 0.00771154
R22068 XThR.Tn[10].n22 XThR.Tn[10].n21 0.00771154
R22069 XThR.Tn[10].n17 XThR.Tn[10].n16 0.00771154
R22070 XThR.Tn[10].n12 XThR.Tn[10].n11 0.00771154
R22071 XThC.Tn[14].n5 XThC.Tn[14].n4 256.104
R22072 XThC.Tn[14].n8 XThC.Tn[14].n6 243.68
R22073 XThC.Tn[14].n2 XThC.Tn[14].n0 241.847
R22074 XThC.Tn[14].n8 XThC.Tn[14].n7 205.28
R22075 XThC.Tn[14].n5 XThC.Tn[14].n3 202.095
R22076 XThC.Tn[14].n2 XThC.Tn[14].n1 185
R22077 XThC.Tn[14].n12 XThC.Tn[14].n10 161.406
R22078 XThC.Tn[14].n15 XThC.Tn[14].n13 161.406
R22079 XThC.Tn[14].n18 XThC.Tn[14].n16 161.406
R22080 XThC.Tn[14].n21 XThC.Tn[14].n19 161.406
R22081 XThC.Tn[14].n24 XThC.Tn[14].n22 161.406
R22082 XThC.Tn[14].n27 XThC.Tn[14].n25 161.406
R22083 XThC.Tn[14].n30 XThC.Tn[14].n28 161.406
R22084 XThC.Tn[14].n33 XThC.Tn[14].n31 161.406
R22085 XThC.Tn[14].n36 XThC.Tn[14].n34 161.406
R22086 XThC.Tn[14].n39 XThC.Tn[14].n37 161.406
R22087 XThC.Tn[14].n42 XThC.Tn[14].n40 161.406
R22088 XThC.Tn[14].n45 XThC.Tn[14].n43 161.406
R22089 XThC.Tn[14].n48 XThC.Tn[14].n46 161.406
R22090 XThC.Tn[14].n51 XThC.Tn[14].n49 161.406
R22091 XThC.Tn[14].n54 XThC.Tn[14].n52 161.406
R22092 XThC.Tn[14].n57 XThC.Tn[14].n55 161.406
R22093 XThC.Tn[14].n10 XThC.Tn[14].t38 161.202
R22094 XThC.Tn[14].n13 XThC.Tn[14].t22 161.202
R22095 XThC.Tn[14].n16 XThC.Tn[14].t25 161.202
R22096 XThC.Tn[14].n19 XThC.Tn[14].t26 161.202
R22097 XThC.Tn[14].n22 XThC.Tn[14].t14 161.202
R22098 XThC.Tn[14].n25 XThC.Tn[14].t17 161.202
R22099 XThC.Tn[14].n28 XThC.Tn[14].t31 161.202
R22100 XThC.Tn[14].n31 XThC.Tn[14].t39 161.202
R22101 XThC.Tn[14].n34 XThC.Tn[14].t41 161.202
R22102 XThC.Tn[14].n37 XThC.Tn[14].t27 161.202
R22103 XThC.Tn[14].n40 XThC.Tn[14].t30 161.202
R22104 XThC.Tn[14].n43 XThC.Tn[14].t42 161.202
R22105 XThC.Tn[14].n46 XThC.Tn[14].t19 161.202
R22106 XThC.Tn[14].n49 XThC.Tn[14].t21 161.202
R22107 XThC.Tn[14].n52 XThC.Tn[14].t33 161.202
R22108 XThC.Tn[14].n55 XThC.Tn[14].t12 161.202
R22109 XThC.Tn[14].n10 XThC.Tn[14].t43 145.137
R22110 XThC.Tn[14].n13 XThC.Tn[14].t29 145.137
R22111 XThC.Tn[14].n16 XThC.Tn[14].t32 145.137
R22112 XThC.Tn[14].n19 XThC.Tn[14].t34 145.137
R22113 XThC.Tn[14].n22 XThC.Tn[14].t20 145.137
R22114 XThC.Tn[14].n25 XThC.Tn[14].t23 145.137
R22115 XThC.Tn[14].n28 XThC.Tn[14].t37 145.137
R22116 XThC.Tn[14].n31 XThC.Tn[14].t13 145.137
R22117 XThC.Tn[14].n34 XThC.Tn[14].t15 145.137
R22118 XThC.Tn[14].n37 XThC.Tn[14].t35 145.137
R22119 XThC.Tn[14].n40 XThC.Tn[14].t36 145.137
R22120 XThC.Tn[14].n43 XThC.Tn[14].t16 145.137
R22121 XThC.Tn[14].n46 XThC.Tn[14].t24 145.137
R22122 XThC.Tn[14].n49 XThC.Tn[14].t28 145.137
R22123 XThC.Tn[14].n52 XThC.Tn[14].t40 145.137
R22124 XThC.Tn[14].n55 XThC.Tn[14].t18 145.137
R22125 XThC.Tn[14].n3 XThC.Tn[14].t4 26.5955
R22126 XThC.Tn[14].n3 XThC.Tn[14].t5 26.5955
R22127 XThC.Tn[14].n4 XThC.Tn[14].t7 26.5955
R22128 XThC.Tn[14].n4 XThC.Tn[14].t6 26.5955
R22129 XThC.Tn[14].n6 XThC.Tn[14].t11 26.5955
R22130 XThC.Tn[14].n6 XThC.Tn[14].t10 26.5955
R22131 XThC.Tn[14].n7 XThC.Tn[14].t9 26.5955
R22132 XThC.Tn[14].n7 XThC.Tn[14].t8 26.5955
R22133 XThC.Tn[14].n0 XThC.Tn[14].t0 24.9236
R22134 XThC.Tn[14].n0 XThC.Tn[14].t2 24.9236
R22135 XThC.Tn[14].n1 XThC.Tn[14].t1 24.9236
R22136 XThC.Tn[14].n1 XThC.Tn[14].t3 24.9236
R22137 XThC.Tn[14] XThC.Tn[14].n8 22.9652
R22138 XThC.Tn[14] XThC.Tn[14].n2 22.9615
R22139 XThC.Tn[14].n9 XThC.Tn[14].n5 13.9299
R22140 XThC.Tn[14].n9 XThC.Tn[14] 13.9299
R22141 XThC.Tn[14].n58 XThC.Tn[14] 5.65386
R22142 XThC.Tn[14].n59 XThC.Tn[14].n58 5.13312
R22143 XThC.Tn[14].n59 XThC.Tn[14].n9 2.99115
R22144 XThC.Tn[14].n9 XThC.Tn[14] 2.87153
R22145 XThC.Tn[14] XThC.Tn[14].n59 2.2734
R22146 XThC.Tn[14].n15 XThC.Tn[14] 0.931056
R22147 XThC.Tn[14].n18 XThC.Tn[14] 0.931056
R22148 XThC.Tn[14].n21 XThC.Tn[14] 0.931056
R22149 XThC.Tn[14].n24 XThC.Tn[14] 0.931056
R22150 XThC.Tn[14].n27 XThC.Tn[14] 0.931056
R22151 XThC.Tn[14].n30 XThC.Tn[14] 0.931056
R22152 XThC.Tn[14].n33 XThC.Tn[14] 0.931056
R22153 XThC.Tn[14].n36 XThC.Tn[14] 0.931056
R22154 XThC.Tn[14].n39 XThC.Tn[14] 0.931056
R22155 XThC.Tn[14].n42 XThC.Tn[14] 0.931056
R22156 XThC.Tn[14].n45 XThC.Tn[14] 0.931056
R22157 XThC.Tn[14].n48 XThC.Tn[14] 0.931056
R22158 XThC.Tn[14].n51 XThC.Tn[14] 0.931056
R22159 XThC.Tn[14].n54 XThC.Tn[14] 0.931056
R22160 XThC.Tn[14].n57 XThC.Tn[14] 0.931056
R22161 XThC.Tn[14] XThC.Tn[14].n12 0.396333
R22162 XThC.Tn[14] XThC.Tn[14].n15 0.396333
R22163 XThC.Tn[14] XThC.Tn[14].n18 0.396333
R22164 XThC.Tn[14] XThC.Tn[14].n21 0.396333
R22165 XThC.Tn[14] XThC.Tn[14].n24 0.396333
R22166 XThC.Tn[14] XThC.Tn[14].n27 0.396333
R22167 XThC.Tn[14] XThC.Tn[14].n30 0.396333
R22168 XThC.Tn[14] XThC.Tn[14].n33 0.396333
R22169 XThC.Tn[14] XThC.Tn[14].n36 0.396333
R22170 XThC.Tn[14] XThC.Tn[14].n39 0.396333
R22171 XThC.Tn[14] XThC.Tn[14].n42 0.396333
R22172 XThC.Tn[14] XThC.Tn[14].n45 0.396333
R22173 XThC.Tn[14] XThC.Tn[14].n48 0.396333
R22174 XThC.Tn[14] XThC.Tn[14].n51 0.396333
R22175 XThC.Tn[14] XThC.Tn[14].n54 0.396333
R22176 XThC.Tn[14] XThC.Tn[14].n57 0.396333
R22177 XThC.Tn[14].n11 XThC.Tn[14] 0.104667
R22178 XThC.Tn[14].n14 XThC.Tn[14] 0.104667
R22179 XThC.Tn[14].n17 XThC.Tn[14] 0.104667
R22180 XThC.Tn[14].n20 XThC.Tn[14] 0.104667
R22181 XThC.Tn[14].n23 XThC.Tn[14] 0.104667
R22182 XThC.Tn[14].n26 XThC.Tn[14] 0.104667
R22183 XThC.Tn[14].n29 XThC.Tn[14] 0.104667
R22184 XThC.Tn[14].n32 XThC.Tn[14] 0.104667
R22185 XThC.Tn[14].n35 XThC.Tn[14] 0.104667
R22186 XThC.Tn[14].n38 XThC.Tn[14] 0.104667
R22187 XThC.Tn[14].n41 XThC.Tn[14] 0.104667
R22188 XThC.Tn[14].n44 XThC.Tn[14] 0.104667
R22189 XThC.Tn[14].n47 XThC.Tn[14] 0.104667
R22190 XThC.Tn[14].n50 XThC.Tn[14] 0.104667
R22191 XThC.Tn[14].n53 XThC.Tn[14] 0.104667
R22192 XThC.Tn[14].n56 XThC.Tn[14] 0.104667
R22193 XThC.Tn[14].n11 XThC.Tn[14] 0.0309878
R22194 XThC.Tn[14].n14 XThC.Tn[14] 0.0309878
R22195 XThC.Tn[14].n17 XThC.Tn[14] 0.0309878
R22196 XThC.Tn[14].n20 XThC.Tn[14] 0.0309878
R22197 XThC.Tn[14].n23 XThC.Tn[14] 0.0309878
R22198 XThC.Tn[14].n26 XThC.Tn[14] 0.0309878
R22199 XThC.Tn[14].n29 XThC.Tn[14] 0.0309878
R22200 XThC.Tn[14].n32 XThC.Tn[14] 0.0309878
R22201 XThC.Tn[14].n35 XThC.Tn[14] 0.0309878
R22202 XThC.Tn[14].n38 XThC.Tn[14] 0.0309878
R22203 XThC.Tn[14].n41 XThC.Tn[14] 0.0309878
R22204 XThC.Tn[14].n44 XThC.Tn[14] 0.0309878
R22205 XThC.Tn[14].n47 XThC.Tn[14] 0.0309878
R22206 XThC.Tn[14].n50 XThC.Tn[14] 0.0309878
R22207 XThC.Tn[14].n53 XThC.Tn[14] 0.0309878
R22208 XThC.Tn[14].n56 XThC.Tn[14] 0.0309878
R22209 XThC.Tn[14].n12 XThC.Tn[14].n11 0.027939
R22210 XThC.Tn[14].n15 XThC.Tn[14].n14 0.027939
R22211 XThC.Tn[14].n18 XThC.Tn[14].n17 0.027939
R22212 XThC.Tn[14].n21 XThC.Tn[14].n20 0.027939
R22213 XThC.Tn[14].n24 XThC.Tn[14].n23 0.027939
R22214 XThC.Tn[14].n27 XThC.Tn[14].n26 0.027939
R22215 XThC.Tn[14].n30 XThC.Tn[14].n29 0.027939
R22216 XThC.Tn[14].n33 XThC.Tn[14].n32 0.027939
R22217 XThC.Tn[14].n36 XThC.Tn[14].n35 0.027939
R22218 XThC.Tn[14].n39 XThC.Tn[14].n38 0.027939
R22219 XThC.Tn[14].n42 XThC.Tn[14].n41 0.027939
R22220 XThC.Tn[14].n45 XThC.Tn[14].n44 0.027939
R22221 XThC.Tn[14].n48 XThC.Tn[14].n47 0.027939
R22222 XThC.Tn[14].n51 XThC.Tn[14].n50 0.027939
R22223 XThC.Tn[14].n54 XThC.Tn[14].n53 0.027939
R22224 XThC.Tn[14].n57 XThC.Tn[14].n56 0.027939
R22225 XThC.Tn[14].n58 XThC.Tn[14] 0.00250754
R22226 XThC.XTB1.Y.n6 XThC.XTB1.Y.t11 212.081
R22227 XThC.XTB1.Y.n5 XThC.XTB1.Y.t8 212.081
R22228 XThC.XTB1.Y.n11 XThC.XTB1.Y.t6 212.081
R22229 XThC.XTB1.Y.n3 XThC.XTB1.Y.t17 212.081
R22230 XThC.XTB1.Y.n15 XThC.XTB1.Y.t10 212.081
R22231 XThC.XTB1.Y.n16 XThC.XTB1.Y.t14 212.081
R22232 XThC.XTB1.Y.n18 XThC.XTB1.Y.t7 212.081
R22233 XThC.XTB1.Y.n14 XThC.XTB1.Y.t18 212.081
R22234 XThC.XTB1.Y.n22 XThC.XTB1.Y.n2 201.288
R22235 XThC.XTB1.Y.n8 XThC.XTB1.Y.n7 173.761
R22236 XThC.XTB1.Y.n17 XThC.XTB1.Y 158.656
R22237 XThC.XTB1.Y.n10 XThC.XTB1.Y.n9 152
R22238 XThC.XTB1.Y.n8 XThC.XTB1.Y.n4 152
R22239 XThC.XTB1.Y.n13 XThC.XTB1.Y.n12 152
R22240 XThC.XTB1.Y.n20 XThC.XTB1.Y.n19 152
R22241 XThC.XTB1.Y.n6 XThC.XTB1.Y.t16 139.78
R22242 XThC.XTB1.Y.n5 XThC.XTB1.Y.t13 139.78
R22243 XThC.XTB1.Y.n11 XThC.XTB1.Y.t12 139.78
R22244 XThC.XTB1.Y.n3 XThC.XTB1.Y.t5 139.78
R22245 XThC.XTB1.Y.n15 XThC.XTB1.Y.t4 139.78
R22246 XThC.XTB1.Y.n16 XThC.XTB1.Y.t3 139.78
R22247 XThC.XTB1.Y.n18 XThC.XTB1.Y.t15 139.78
R22248 XThC.XTB1.Y.n14 XThC.XTB1.Y.t9 139.78
R22249 XThC.XTB1.Y.n0 XThC.XTB1.Y.t1 132.067
R22250 XThC.XTB1.Y.n21 XThC.XTB1.Y 83.4676
R22251 XThC.XTB1.Y.n21 XThC.XTB1.Y.n13 61.4091
R22252 XThC.XTB1.Y.n16 XThC.XTB1.Y.n15 61.346
R22253 XThC.XTB1.Y.n10 XThC.XTB1.Y.n4 49.6611
R22254 XThC.XTB1.Y.n12 XThC.XTB1.Y.n11 45.2793
R22255 XThC.XTB1.Y.n7 XThC.XTB1.Y.n5 42.3581
R22256 XThC.XTB1.Y.n19 XThC.XTB1.Y.n14 30.6732
R22257 XThC.XTB1.Y.n19 XThC.XTB1.Y.n18 30.6732
R22258 XThC.XTB1.Y.n18 XThC.XTB1.Y.n17 30.6732
R22259 XThC.XTB1.Y.n17 XThC.XTB1.Y.n16 30.6732
R22260 XThC.XTB1.Y.n2 XThC.XTB1.Y.t2 26.5955
R22261 XThC.XTB1.Y.n2 XThC.XTB1.Y.t0 26.5955
R22262 XThC.XTB1.Y XThC.XTB1.Y.n22 23.489
R22263 XThC.XTB1.Y.n9 XThC.XTB1.Y.n8 21.7605
R22264 XThC.XTB1.Y.n7 XThC.XTB1.Y.n6 18.9884
R22265 XThC.XTB1.Y.n12 XThC.XTB1.Y.n3 16.0672
R22266 XThC.XTB1.Y.n20 XThC.XTB1.Y 14.8485
R22267 XThC.XTB1.Y.n13 XThC.XTB1.Y 11.5205
R22268 XThC.XTB1.Y.n22 XThC.XTB1.Y.n21 10.7939
R22269 XThC.XTB1.Y.n9 XThC.XTB1.Y 10.2405
R22270 XThC.XTB1.Y XThC.XTB1.Y.n20 8.7045
R22271 XThC.XTB1.Y.n5 XThC.XTB1.Y.n4 7.30353
R22272 XThC.XTB1.Y.n11 XThC.XTB1.Y.n10 4.38232
R22273 XThC.XTB1.Y.n1 XThC.XTB1.Y.n0 4.15748
R22274 XThC.XTB1.Y XThC.XTB1.Y.n1 3.76521
R22275 XThC.XTB1.Y.n0 XThC.XTB1.Y 1.17559
R22276 XThC.XTB1.Y.n1 XThC.XTB1.Y 0.921363
R22277 XThC.Tn[8].n5 XThC.Tn[8].n4 256.104
R22278 XThC.Tn[8].n8 XThC.Tn[8].n6 243.68
R22279 XThC.Tn[8].n2 XThC.Tn[8].n0 241.847
R22280 XThC.Tn[8].n8 XThC.Tn[8].n7 205.28
R22281 XThC.Tn[8].n5 XThC.Tn[8].n3 202.095
R22282 XThC.Tn[8].n2 XThC.Tn[8].n1 185
R22283 XThC.Tn[8].n12 XThC.Tn[8].n10 161.406
R22284 XThC.Tn[8].n15 XThC.Tn[8].n13 161.406
R22285 XThC.Tn[8].n18 XThC.Tn[8].n16 161.406
R22286 XThC.Tn[8].n21 XThC.Tn[8].n19 161.406
R22287 XThC.Tn[8].n24 XThC.Tn[8].n22 161.406
R22288 XThC.Tn[8].n27 XThC.Tn[8].n25 161.406
R22289 XThC.Tn[8].n30 XThC.Tn[8].n28 161.406
R22290 XThC.Tn[8].n33 XThC.Tn[8].n31 161.406
R22291 XThC.Tn[8].n36 XThC.Tn[8].n34 161.406
R22292 XThC.Tn[8].n39 XThC.Tn[8].n37 161.406
R22293 XThC.Tn[8].n42 XThC.Tn[8].n40 161.406
R22294 XThC.Tn[8].n45 XThC.Tn[8].n43 161.406
R22295 XThC.Tn[8].n48 XThC.Tn[8].n46 161.406
R22296 XThC.Tn[8].n51 XThC.Tn[8].n49 161.406
R22297 XThC.Tn[8].n54 XThC.Tn[8].n52 161.406
R22298 XThC.Tn[8].n57 XThC.Tn[8].n55 161.406
R22299 XThC.Tn[8].n10 XThC.Tn[8].t41 161.202
R22300 XThC.Tn[8].n13 XThC.Tn[8].t26 161.202
R22301 XThC.Tn[8].n16 XThC.Tn[8].t28 161.202
R22302 XThC.Tn[8].n19 XThC.Tn[8].t30 161.202
R22303 XThC.Tn[8].n22 XThC.Tn[8].t19 161.202
R22304 XThC.Tn[8].n25 XThC.Tn[8].t20 161.202
R22305 XThC.Tn[8].n28 XThC.Tn[8].t33 161.202
R22306 XThC.Tn[8].n31 XThC.Tn[8].t42 161.202
R22307 XThC.Tn[8].n34 XThC.Tn[8].t12 161.202
R22308 XThC.Tn[8].n37 XThC.Tn[8].t31 161.202
R22309 XThC.Tn[8].n40 XThC.Tn[8].t32 161.202
R22310 XThC.Tn[8].n43 XThC.Tn[8].t13 161.202
R22311 XThC.Tn[8].n46 XThC.Tn[8].t21 161.202
R22312 XThC.Tn[8].n49 XThC.Tn[8].t24 161.202
R22313 XThC.Tn[8].n52 XThC.Tn[8].t37 161.202
R22314 XThC.Tn[8].n55 XThC.Tn[8].t15 161.202
R22315 XThC.Tn[8].n10 XThC.Tn[8].t43 145.137
R22316 XThC.Tn[8].n13 XThC.Tn[8].t29 145.137
R22317 XThC.Tn[8].n16 XThC.Tn[8].t34 145.137
R22318 XThC.Tn[8].n19 XThC.Tn[8].t35 145.137
R22319 XThC.Tn[8].n22 XThC.Tn[8].t22 145.137
R22320 XThC.Tn[8].n25 XThC.Tn[8].t23 145.137
R22321 XThC.Tn[8].n28 XThC.Tn[8].t39 145.137
R22322 XThC.Tn[8].n31 XThC.Tn[8].t14 145.137
R22323 XThC.Tn[8].n34 XThC.Tn[8].t16 145.137
R22324 XThC.Tn[8].n37 XThC.Tn[8].t36 145.137
R22325 XThC.Tn[8].n40 XThC.Tn[8].t38 145.137
R22326 XThC.Tn[8].n43 XThC.Tn[8].t17 145.137
R22327 XThC.Tn[8].n46 XThC.Tn[8].t25 145.137
R22328 XThC.Tn[8].n49 XThC.Tn[8].t27 145.137
R22329 XThC.Tn[8].n52 XThC.Tn[8].t40 145.137
R22330 XThC.Tn[8].n55 XThC.Tn[8].t18 145.137
R22331 XThC.Tn[8].n3 XThC.Tn[8].t5 26.5955
R22332 XThC.Tn[8].n3 XThC.Tn[8].t6 26.5955
R22333 XThC.Tn[8].n4 XThC.Tn[8].t4 26.5955
R22334 XThC.Tn[8].n4 XThC.Tn[8].t7 26.5955
R22335 XThC.Tn[8].n6 XThC.Tn[8].t8 26.5955
R22336 XThC.Tn[8].n6 XThC.Tn[8].t11 26.5955
R22337 XThC.Tn[8].n7 XThC.Tn[8].t10 26.5955
R22338 XThC.Tn[8].n7 XThC.Tn[8].t9 26.5955
R22339 XThC.Tn[8].n0 XThC.Tn[8].t1 24.9236
R22340 XThC.Tn[8].n0 XThC.Tn[8].t0 24.9236
R22341 XThC.Tn[8].n1 XThC.Tn[8].t3 24.9236
R22342 XThC.Tn[8].n1 XThC.Tn[8].t2 24.9236
R22343 XThC.Tn[8] XThC.Tn[8].n8 22.9652
R22344 XThC.Tn[8] XThC.Tn[8].n2 22.9615
R22345 XThC.Tn[8].n9 XThC.Tn[8].n5 13.9299
R22346 XThC.Tn[8].n9 XThC.Tn[8] 13.9299
R22347 XThC.Tn[8].n60 XThC.Tn[8].n59 5.09639
R22348 XThC.Tn[8].n60 XThC.Tn[8].n9 2.99115
R22349 XThC.Tn[8].n9 XThC.Tn[8] 2.87153
R22350 XThC.Tn[8] XThC.Tn[8].n60 2.2734
R22351 XThC.Tn[8].n58 XThC.Tn[8] 1.14336
R22352 XThC.Tn[8].n15 XThC.Tn[8] 0.931056
R22353 XThC.Tn[8].n18 XThC.Tn[8] 0.931056
R22354 XThC.Tn[8].n21 XThC.Tn[8] 0.931056
R22355 XThC.Tn[8].n24 XThC.Tn[8] 0.931056
R22356 XThC.Tn[8].n27 XThC.Tn[8] 0.931056
R22357 XThC.Tn[8].n30 XThC.Tn[8] 0.931056
R22358 XThC.Tn[8].n33 XThC.Tn[8] 0.931056
R22359 XThC.Tn[8].n36 XThC.Tn[8] 0.931056
R22360 XThC.Tn[8].n39 XThC.Tn[8] 0.931056
R22361 XThC.Tn[8].n42 XThC.Tn[8] 0.931056
R22362 XThC.Tn[8].n45 XThC.Tn[8] 0.931056
R22363 XThC.Tn[8].n48 XThC.Tn[8] 0.931056
R22364 XThC.Tn[8].n51 XThC.Tn[8] 0.931056
R22365 XThC.Tn[8].n54 XThC.Tn[8] 0.931056
R22366 XThC.Tn[8].n57 XThC.Tn[8] 0.931056
R22367 XThC.Tn[8] XThC.Tn[8].n12 0.396333
R22368 XThC.Tn[8] XThC.Tn[8].n15 0.396333
R22369 XThC.Tn[8] XThC.Tn[8].n18 0.396333
R22370 XThC.Tn[8] XThC.Tn[8].n21 0.396333
R22371 XThC.Tn[8] XThC.Tn[8].n24 0.396333
R22372 XThC.Tn[8] XThC.Tn[8].n27 0.396333
R22373 XThC.Tn[8] XThC.Tn[8].n30 0.396333
R22374 XThC.Tn[8] XThC.Tn[8].n33 0.396333
R22375 XThC.Tn[8] XThC.Tn[8].n36 0.396333
R22376 XThC.Tn[8] XThC.Tn[8].n39 0.396333
R22377 XThC.Tn[8] XThC.Tn[8].n42 0.396333
R22378 XThC.Tn[8] XThC.Tn[8].n45 0.396333
R22379 XThC.Tn[8] XThC.Tn[8].n48 0.396333
R22380 XThC.Tn[8] XThC.Tn[8].n51 0.396333
R22381 XThC.Tn[8] XThC.Tn[8].n54 0.396333
R22382 XThC.Tn[8] XThC.Tn[8].n57 0.396333
R22383 XThC.Tn[8].n59 XThC.Tn[8].n58 0.166125
R22384 XThC.Tn[8].n11 XThC.Tn[8] 0.104667
R22385 XThC.Tn[8].n14 XThC.Tn[8] 0.104667
R22386 XThC.Tn[8].n17 XThC.Tn[8] 0.104667
R22387 XThC.Tn[8].n20 XThC.Tn[8] 0.104667
R22388 XThC.Tn[8].n23 XThC.Tn[8] 0.104667
R22389 XThC.Tn[8].n26 XThC.Tn[8] 0.104667
R22390 XThC.Tn[8].n29 XThC.Tn[8] 0.104667
R22391 XThC.Tn[8].n32 XThC.Tn[8] 0.104667
R22392 XThC.Tn[8].n35 XThC.Tn[8] 0.104667
R22393 XThC.Tn[8].n38 XThC.Tn[8] 0.104667
R22394 XThC.Tn[8].n41 XThC.Tn[8] 0.104667
R22395 XThC.Tn[8].n44 XThC.Tn[8] 0.104667
R22396 XThC.Tn[8].n47 XThC.Tn[8] 0.104667
R22397 XThC.Tn[8].n50 XThC.Tn[8] 0.104667
R22398 XThC.Tn[8].n53 XThC.Tn[8] 0.104667
R22399 XThC.Tn[8].n56 XThC.Tn[8] 0.104667
R22400 XThC.Tn[8].n59 XThC.Tn[8] 0.0389615
R22401 XThC.Tn[8].n58 XThC.Tn[8] 0.038
R22402 XThC.Tn[8].n11 XThC.Tn[8] 0.0309878
R22403 XThC.Tn[8].n14 XThC.Tn[8] 0.0309878
R22404 XThC.Tn[8].n17 XThC.Tn[8] 0.0309878
R22405 XThC.Tn[8].n20 XThC.Tn[8] 0.0309878
R22406 XThC.Tn[8].n23 XThC.Tn[8] 0.0309878
R22407 XThC.Tn[8].n26 XThC.Tn[8] 0.0309878
R22408 XThC.Tn[8].n29 XThC.Tn[8] 0.0309878
R22409 XThC.Tn[8].n32 XThC.Tn[8] 0.0309878
R22410 XThC.Tn[8].n35 XThC.Tn[8] 0.0309878
R22411 XThC.Tn[8].n38 XThC.Tn[8] 0.0309878
R22412 XThC.Tn[8].n41 XThC.Tn[8] 0.0309878
R22413 XThC.Tn[8].n44 XThC.Tn[8] 0.0309878
R22414 XThC.Tn[8].n47 XThC.Tn[8] 0.0309878
R22415 XThC.Tn[8].n50 XThC.Tn[8] 0.0309878
R22416 XThC.Tn[8].n53 XThC.Tn[8] 0.0309878
R22417 XThC.Tn[8].n56 XThC.Tn[8] 0.0309878
R22418 XThC.Tn[8].n12 XThC.Tn[8].n11 0.027939
R22419 XThC.Tn[8].n15 XThC.Tn[8].n14 0.027939
R22420 XThC.Tn[8].n18 XThC.Tn[8].n17 0.027939
R22421 XThC.Tn[8].n21 XThC.Tn[8].n20 0.027939
R22422 XThC.Tn[8].n24 XThC.Tn[8].n23 0.027939
R22423 XThC.Tn[8].n27 XThC.Tn[8].n26 0.027939
R22424 XThC.Tn[8].n30 XThC.Tn[8].n29 0.027939
R22425 XThC.Tn[8].n33 XThC.Tn[8].n32 0.027939
R22426 XThC.Tn[8].n36 XThC.Tn[8].n35 0.027939
R22427 XThC.Tn[8].n39 XThC.Tn[8].n38 0.027939
R22428 XThC.Tn[8].n42 XThC.Tn[8].n41 0.027939
R22429 XThC.Tn[8].n45 XThC.Tn[8].n44 0.027939
R22430 XThC.Tn[8].n48 XThC.Tn[8].n47 0.027939
R22431 XThC.Tn[8].n51 XThC.Tn[8].n50 0.027939
R22432 XThC.Tn[8].n54 XThC.Tn[8].n53 0.027939
R22433 XThC.Tn[8].n57 XThC.Tn[8].n56 0.027939
R22434 XThR.Tn[1].n88 XThR.Tn[1].n87 332.334
R22435 XThR.Tn[1].n88 XThR.Tn[1].n86 296.493
R22436 XThR.Tn[1] XThR.Tn[1].n79 161.363
R22437 XThR.Tn[1] XThR.Tn[1].n74 161.363
R22438 XThR.Tn[1] XThR.Tn[1].n69 161.363
R22439 XThR.Tn[1] XThR.Tn[1].n64 161.363
R22440 XThR.Tn[1] XThR.Tn[1].n59 161.363
R22441 XThR.Tn[1] XThR.Tn[1].n54 161.363
R22442 XThR.Tn[1] XThR.Tn[1].n49 161.363
R22443 XThR.Tn[1] XThR.Tn[1].n44 161.363
R22444 XThR.Tn[1] XThR.Tn[1].n39 161.363
R22445 XThR.Tn[1] XThR.Tn[1].n34 161.363
R22446 XThR.Tn[1] XThR.Tn[1].n29 161.363
R22447 XThR.Tn[1] XThR.Tn[1].n24 161.363
R22448 XThR.Tn[1] XThR.Tn[1].n19 161.363
R22449 XThR.Tn[1] XThR.Tn[1].n14 161.363
R22450 XThR.Tn[1] XThR.Tn[1].n9 161.363
R22451 XThR.Tn[1] XThR.Tn[1].n7 161.363
R22452 XThR.Tn[1].n81 XThR.Tn[1].n80 161.3
R22453 XThR.Tn[1].n76 XThR.Tn[1].n75 161.3
R22454 XThR.Tn[1].n71 XThR.Tn[1].n70 161.3
R22455 XThR.Tn[1].n66 XThR.Tn[1].n65 161.3
R22456 XThR.Tn[1].n61 XThR.Tn[1].n60 161.3
R22457 XThR.Tn[1].n56 XThR.Tn[1].n55 161.3
R22458 XThR.Tn[1].n51 XThR.Tn[1].n50 161.3
R22459 XThR.Tn[1].n46 XThR.Tn[1].n45 161.3
R22460 XThR.Tn[1].n41 XThR.Tn[1].n40 161.3
R22461 XThR.Tn[1].n36 XThR.Tn[1].n35 161.3
R22462 XThR.Tn[1].n31 XThR.Tn[1].n30 161.3
R22463 XThR.Tn[1].n26 XThR.Tn[1].n25 161.3
R22464 XThR.Tn[1].n21 XThR.Tn[1].n20 161.3
R22465 XThR.Tn[1].n16 XThR.Tn[1].n15 161.3
R22466 XThR.Tn[1].n11 XThR.Tn[1].n10 161.3
R22467 XThR.Tn[1].n79 XThR.Tn[1].t70 161.106
R22468 XThR.Tn[1].n74 XThR.Tn[1].t14 161.106
R22469 XThR.Tn[1].n69 XThR.Tn[1].t56 161.106
R22470 XThR.Tn[1].n64 XThR.Tn[1].t42 161.106
R22471 XThR.Tn[1].n59 XThR.Tn[1].t68 161.106
R22472 XThR.Tn[1].n54 XThR.Tn[1].t31 161.106
R22473 XThR.Tn[1].n49 XThR.Tn[1].t12 161.106
R22474 XThR.Tn[1].n44 XThR.Tn[1].t54 161.106
R22475 XThR.Tn[1].n39 XThR.Tn[1].t41 161.106
R22476 XThR.Tn[1].n34 XThR.Tn[1].t46 161.106
R22477 XThR.Tn[1].n29 XThR.Tn[1].t29 161.106
R22478 XThR.Tn[1].n24 XThR.Tn[1].t55 161.106
R22479 XThR.Tn[1].n19 XThR.Tn[1].t28 161.106
R22480 XThR.Tn[1].n14 XThR.Tn[1].t73 161.106
R22481 XThR.Tn[1].n9 XThR.Tn[1].t34 161.106
R22482 XThR.Tn[1].n7 XThR.Tn[1].t18 161.106
R22483 XThR.Tn[1].n80 XThR.Tn[1].t66 159.978
R22484 XThR.Tn[1].n75 XThR.Tn[1].t72 159.978
R22485 XThR.Tn[1].n70 XThR.Tn[1].t52 159.978
R22486 XThR.Tn[1].n65 XThR.Tn[1].t39 159.978
R22487 XThR.Tn[1].n60 XThR.Tn[1].t63 159.978
R22488 XThR.Tn[1].n55 XThR.Tn[1].t27 159.978
R22489 XThR.Tn[1].n50 XThR.Tn[1].t71 159.978
R22490 XThR.Tn[1].n45 XThR.Tn[1].t49 159.978
R22491 XThR.Tn[1].n40 XThR.Tn[1].t36 159.978
R22492 XThR.Tn[1].n35 XThR.Tn[1].t43 159.978
R22493 XThR.Tn[1].n30 XThR.Tn[1].t26 159.978
R22494 XThR.Tn[1].n25 XThR.Tn[1].t51 159.978
R22495 XThR.Tn[1].n20 XThR.Tn[1].t25 159.978
R22496 XThR.Tn[1].n15 XThR.Tn[1].t69 159.978
R22497 XThR.Tn[1].n10 XThR.Tn[1].t30 159.978
R22498 XThR.Tn[1].n79 XThR.Tn[1].t58 145.038
R22499 XThR.Tn[1].n74 XThR.Tn[1].t20 145.038
R22500 XThR.Tn[1].n69 XThR.Tn[1].t62 145.038
R22501 XThR.Tn[1].n64 XThR.Tn[1].t47 145.038
R22502 XThR.Tn[1].n59 XThR.Tn[1].t15 145.038
R22503 XThR.Tn[1].n54 XThR.Tn[1].t57 145.038
R22504 XThR.Tn[1].n49 XThR.Tn[1].t64 145.038
R22505 XThR.Tn[1].n44 XThR.Tn[1].t48 145.038
R22506 XThR.Tn[1].n39 XThR.Tn[1].t45 145.038
R22507 XThR.Tn[1].n34 XThR.Tn[1].t13 145.038
R22508 XThR.Tn[1].n29 XThR.Tn[1].t37 145.038
R22509 XThR.Tn[1].n24 XThR.Tn[1].t59 145.038
R22510 XThR.Tn[1].n19 XThR.Tn[1].t35 145.038
R22511 XThR.Tn[1].n14 XThR.Tn[1].t19 145.038
R22512 XThR.Tn[1].n9 XThR.Tn[1].t44 145.038
R22513 XThR.Tn[1].n7 XThR.Tn[1].t24 145.038
R22514 XThR.Tn[1].n80 XThR.Tn[1].t17 143.911
R22515 XThR.Tn[1].n75 XThR.Tn[1].t40 143.911
R22516 XThR.Tn[1].n70 XThR.Tn[1].t22 143.911
R22517 XThR.Tn[1].n65 XThR.Tn[1].t65 143.911
R22518 XThR.Tn[1].n60 XThR.Tn[1].t33 143.911
R22519 XThR.Tn[1].n55 XThR.Tn[1].t16 143.911
R22520 XThR.Tn[1].n50 XThR.Tn[1].t23 143.911
R22521 XThR.Tn[1].n45 XThR.Tn[1].t67 143.911
R22522 XThR.Tn[1].n40 XThR.Tn[1].t60 143.911
R22523 XThR.Tn[1].n35 XThR.Tn[1].t32 143.911
R22524 XThR.Tn[1].n30 XThR.Tn[1].t53 143.911
R22525 XThR.Tn[1].n25 XThR.Tn[1].t21 143.911
R22526 XThR.Tn[1].n20 XThR.Tn[1].t50 143.911
R22527 XThR.Tn[1].n15 XThR.Tn[1].t38 143.911
R22528 XThR.Tn[1].n10 XThR.Tn[1].t61 143.911
R22529 XThR.Tn[1].n2 XThR.Tn[1].n0 135.249
R22530 XThR.Tn[1].n2 XThR.Tn[1].n1 98.981
R22531 XThR.Tn[1].n4 XThR.Tn[1].n3 98.981
R22532 XThR.Tn[1].n6 XThR.Tn[1].n5 98.981
R22533 XThR.Tn[1].n4 XThR.Tn[1].n2 36.2672
R22534 XThR.Tn[1].n6 XThR.Tn[1].n4 36.2672
R22535 XThR.Tn[1].n85 XThR.Tn[1].n6 32.6405
R22536 XThR.Tn[1].n86 XThR.Tn[1].t0 26.5955
R22537 XThR.Tn[1].n86 XThR.Tn[1].t1 26.5955
R22538 XThR.Tn[1].n87 XThR.Tn[1].t3 26.5955
R22539 XThR.Tn[1].n87 XThR.Tn[1].t2 26.5955
R22540 XThR.Tn[1].n0 XThR.Tn[1].t11 24.9236
R22541 XThR.Tn[1].n0 XThR.Tn[1].t8 24.9236
R22542 XThR.Tn[1].n1 XThR.Tn[1].t10 24.9236
R22543 XThR.Tn[1].n1 XThR.Tn[1].t9 24.9236
R22544 XThR.Tn[1].n3 XThR.Tn[1].t6 24.9236
R22545 XThR.Tn[1].n3 XThR.Tn[1].t5 24.9236
R22546 XThR.Tn[1].n5 XThR.Tn[1].t7 24.9236
R22547 XThR.Tn[1].n5 XThR.Tn[1].t4 24.9236
R22548 XThR.Tn[1].n89 XThR.Tn[1].n88 18.5605
R22549 XThR.Tn[1].n89 XThR.Tn[1].n85 11.5205
R22550 XThR.Tn[1].n85 XThR.Tn[1] 6.42118
R22551 XThR.Tn[1] XThR.Tn[1].n8 5.34038
R22552 XThR.Tn[1].n13 XThR.Tn[1].n12 4.5005
R22553 XThR.Tn[1].n18 XThR.Tn[1].n17 4.5005
R22554 XThR.Tn[1].n23 XThR.Tn[1].n22 4.5005
R22555 XThR.Tn[1].n28 XThR.Tn[1].n27 4.5005
R22556 XThR.Tn[1].n33 XThR.Tn[1].n32 4.5005
R22557 XThR.Tn[1].n38 XThR.Tn[1].n37 4.5005
R22558 XThR.Tn[1].n43 XThR.Tn[1].n42 4.5005
R22559 XThR.Tn[1].n48 XThR.Tn[1].n47 4.5005
R22560 XThR.Tn[1].n53 XThR.Tn[1].n52 4.5005
R22561 XThR.Tn[1].n58 XThR.Tn[1].n57 4.5005
R22562 XThR.Tn[1].n63 XThR.Tn[1].n62 4.5005
R22563 XThR.Tn[1].n68 XThR.Tn[1].n67 4.5005
R22564 XThR.Tn[1].n73 XThR.Tn[1].n72 4.5005
R22565 XThR.Tn[1].n78 XThR.Tn[1].n77 4.5005
R22566 XThR.Tn[1].n83 XThR.Tn[1].n82 4.5005
R22567 XThR.Tn[1].n84 XThR.Tn[1] 3.70586
R22568 XThR.Tn[1].n13 XThR.Tn[1] 2.52282
R22569 XThR.Tn[1].n18 XThR.Tn[1] 2.52282
R22570 XThR.Tn[1].n23 XThR.Tn[1] 2.52282
R22571 XThR.Tn[1].n28 XThR.Tn[1] 2.52282
R22572 XThR.Tn[1].n33 XThR.Tn[1] 2.52282
R22573 XThR.Tn[1].n38 XThR.Tn[1] 2.52282
R22574 XThR.Tn[1].n43 XThR.Tn[1] 2.52282
R22575 XThR.Tn[1].n48 XThR.Tn[1] 2.52282
R22576 XThR.Tn[1].n53 XThR.Tn[1] 2.52282
R22577 XThR.Tn[1].n58 XThR.Tn[1] 2.52282
R22578 XThR.Tn[1].n63 XThR.Tn[1] 2.52282
R22579 XThR.Tn[1].n68 XThR.Tn[1] 2.52282
R22580 XThR.Tn[1].n73 XThR.Tn[1] 2.52282
R22581 XThR.Tn[1].n78 XThR.Tn[1] 2.52282
R22582 XThR.Tn[1].n83 XThR.Tn[1] 2.52282
R22583 XThR.Tn[1].n81 XThR.Tn[1] 1.08677
R22584 XThR.Tn[1].n76 XThR.Tn[1] 1.08677
R22585 XThR.Tn[1].n71 XThR.Tn[1] 1.08677
R22586 XThR.Tn[1].n66 XThR.Tn[1] 1.08677
R22587 XThR.Tn[1].n61 XThR.Tn[1] 1.08677
R22588 XThR.Tn[1].n56 XThR.Tn[1] 1.08677
R22589 XThR.Tn[1].n51 XThR.Tn[1] 1.08677
R22590 XThR.Tn[1].n46 XThR.Tn[1] 1.08677
R22591 XThR.Tn[1].n41 XThR.Tn[1] 1.08677
R22592 XThR.Tn[1].n36 XThR.Tn[1] 1.08677
R22593 XThR.Tn[1].n31 XThR.Tn[1] 1.08677
R22594 XThR.Tn[1].n26 XThR.Tn[1] 1.08677
R22595 XThR.Tn[1].n21 XThR.Tn[1] 1.08677
R22596 XThR.Tn[1].n16 XThR.Tn[1] 1.08677
R22597 XThR.Tn[1].n11 XThR.Tn[1] 1.08677
R22598 XThR.Tn[1] XThR.Tn[1].n13 0.839786
R22599 XThR.Tn[1] XThR.Tn[1].n18 0.839786
R22600 XThR.Tn[1] XThR.Tn[1].n23 0.839786
R22601 XThR.Tn[1] XThR.Tn[1].n28 0.839786
R22602 XThR.Tn[1] XThR.Tn[1].n33 0.839786
R22603 XThR.Tn[1] XThR.Tn[1].n38 0.839786
R22604 XThR.Tn[1] XThR.Tn[1].n43 0.839786
R22605 XThR.Tn[1] XThR.Tn[1].n48 0.839786
R22606 XThR.Tn[1] XThR.Tn[1].n53 0.839786
R22607 XThR.Tn[1] XThR.Tn[1].n58 0.839786
R22608 XThR.Tn[1] XThR.Tn[1].n63 0.839786
R22609 XThR.Tn[1] XThR.Tn[1].n68 0.839786
R22610 XThR.Tn[1] XThR.Tn[1].n73 0.839786
R22611 XThR.Tn[1] XThR.Tn[1].n78 0.839786
R22612 XThR.Tn[1] XThR.Tn[1].n83 0.839786
R22613 XThR.Tn[1] XThR.Tn[1].n89 0.6405
R22614 XThR.Tn[1].n8 XThR.Tn[1] 0.499542
R22615 XThR.Tn[1].n82 XThR.Tn[1] 0.063
R22616 XThR.Tn[1].n77 XThR.Tn[1] 0.063
R22617 XThR.Tn[1].n72 XThR.Tn[1] 0.063
R22618 XThR.Tn[1].n67 XThR.Tn[1] 0.063
R22619 XThR.Tn[1].n62 XThR.Tn[1] 0.063
R22620 XThR.Tn[1].n57 XThR.Tn[1] 0.063
R22621 XThR.Tn[1].n52 XThR.Tn[1] 0.063
R22622 XThR.Tn[1].n47 XThR.Tn[1] 0.063
R22623 XThR.Tn[1].n42 XThR.Tn[1] 0.063
R22624 XThR.Tn[1].n37 XThR.Tn[1] 0.063
R22625 XThR.Tn[1].n32 XThR.Tn[1] 0.063
R22626 XThR.Tn[1].n27 XThR.Tn[1] 0.063
R22627 XThR.Tn[1].n22 XThR.Tn[1] 0.063
R22628 XThR.Tn[1].n17 XThR.Tn[1] 0.063
R22629 XThR.Tn[1].n12 XThR.Tn[1] 0.063
R22630 XThR.Tn[1].n84 XThR.Tn[1] 0.0540714
R22631 XThR.Tn[1] XThR.Tn[1].n84 0.038
R22632 XThR.Tn[1].n8 XThR.Tn[1] 0.0143889
R22633 XThR.Tn[1].n82 XThR.Tn[1].n81 0.00771154
R22634 XThR.Tn[1].n77 XThR.Tn[1].n76 0.00771154
R22635 XThR.Tn[1].n72 XThR.Tn[1].n71 0.00771154
R22636 XThR.Tn[1].n67 XThR.Tn[1].n66 0.00771154
R22637 XThR.Tn[1].n62 XThR.Tn[1].n61 0.00771154
R22638 XThR.Tn[1].n57 XThR.Tn[1].n56 0.00771154
R22639 XThR.Tn[1].n52 XThR.Tn[1].n51 0.00771154
R22640 XThR.Tn[1].n47 XThR.Tn[1].n46 0.00771154
R22641 XThR.Tn[1].n42 XThR.Tn[1].n41 0.00771154
R22642 XThR.Tn[1].n37 XThR.Tn[1].n36 0.00771154
R22643 XThR.Tn[1].n32 XThR.Tn[1].n31 0.00771154
R22644 XThR.Tn[1].n27 XThR.Tn[1].n26 0.00771154
R22645 XThR.Tn[1].n22 XThR.Tn[1].n21 0.00771154
R22646 XThR.Tn[1].n17 XThR.Tn[1].n16 0.00771154
R22647 XThR.Tn[1].n12 XThR.Tn[1].n11 0.00771154
R22648 XThC.Tn[7].n2 XThC.Tn[7].n1 255.096
R22649 XThC.Tn[7].n55 XThC.Tn[7].n53 236.589
R22650 XThC.Tn[7].n2 XThC.Tn[7].n0 201.845
R22651 XThC.Tn[7].n55 XThC.Tn[7].n54 200.321
R22652 XThC.Tn[7].n5 XThC.Tn[7].n3 161.406
R22653 XThC.Tn[7].n8 XThC.Tn[7].n6 161.406
R22654 XThC.Tn[7].n11 XThC.Tn[7].n9 161.406
R22655 XThC.Tn[7].n14 XThC.Tn[7].n12 161.406
R22656 XThC.Tn[7].n17 XThC.Tn[7].n15 161.406
R22657 XThC.Tn[7].n20 XThC.Tn[7].n18 161.406
R22658 XThC.Tn[7].n23 XThC.Tn[7].n21 161.406
R22659 XThC.Tn[7].n26 XThC.Tn[7].n24 161.406
R22660 XThC.Tn[7].n29 XThC.Tn[7].n27 161.406
R22661 XThC.Tn[7].n32 XThC.Tn[7].n30 161.406
R22662 XThC.Tn[7].n35 XThC.Tn[7].n33 161.406
R22663 XThC.Tn[7].n38 XThC.Tn[7].n36 161.406
R22664 XThC.Tn[7].n41 XThC.Tn[7].n39 161.406
R22665 XThC.Tn[7].n44 XThC.Tn[7].n42 161.406
R22666 XThC.Tn[7].n47 XThC.Tn[7].n45 161.406
R22667 XThC.Tn[7].n50 XThC.Tn[7].n48 161.406
R22668 XThC.Tn[7].n3 XThC.Tn[7].t11 161.202
R22669 XThC.Tn[7].n6 XThC.Tn[7].t30 161.202
R22670 XThC.Tn[7].n9 XThC.Tn[7].t34 161.202
R22671 XThC.Tn[7].n12 XThC.Tn[7].t35 161.202
R22672 XThC.Tn[7].n15 XThC.Tn[7].t22 161.202
R22673 XThC.Tn[7].n18 XThC.Tn[7].t23 161.202
R22674 XThC.Tn[7].n21 XThC.Tn[7].t39 161.202
R22675 XThC.Tn[7].n24 XThC.Tn[7].t14 161.202
R22676 XThC.Tn[7].n27 XThC.Tn[7].t16 161.202
R22677 XThC.Tn[7].n30 XThC.Tn[7].t36 161.202
R22678 XThC.Tn[7].n33 XThC.Tn[7].t38 161.202
R22679 XThC.Tn[7].n36 XThC.Tn[7].t17 161.202
R22680 XThC.Tn[7].n39 XThC.Tn[7].t26 161.202
R22681 XThC.Tn[7].n42 XThC.Tn[7].t28 161.202
R22682 XThC.Tn[7].n45 XThC.Tn[7].t9 161.202
R22683 XThC.Tn[7].n48 XThC.Tn[7].t19 161.202
R22684 XThC.Tn[7].n3 XThC.Tn[7].t8 145.137
R22685 XThC.Tn[7].n6 XThC.Tn[7].t25 145.137
R22686 XThC.Tn[7].n9 XThC.Tn[7].t27 145.137
R22687 XThC.Tn[7].n12 XThC.Tn[7].t29 145.137
R22688 XThC.Tn[7].n15 XThC.Tn[7].t18 145.137
R22689 XThC.Tn[7].n18 XThC.Tn[7].t20 145.137
R22690 XThC.Tn[7].n21 XThC.Tn[7].t33 145.137
R22691 XThC.Tn[7].n24 XThC.Tn[7].t10 145.137
R22692 XThC.Tn[7].n27 XThC.Tn[7].t12 145.137
R22693 XThC.Tn[7].n30 XThC.Tn[7].t31 145.137
R22694 XThC.Tn[7].n33 XThC.Tn[7].t32 145.137
R22695 XThC.Tn[7].n36 XThC.Tn[7].t13 145.137
R22696 XThC.Tn[7].n39 XThC.Tn[7].t21 145.137
R22697 XThC.Tn[7].n42 XThC.Tn[7].t24 145.137
R22698 XThC.Tn[7].n45 XThC.Tn[7].t37 145.137
R22699 XThC.Tn[7].n48 XThC.Tn[7].t15 145.137
R22700 XThC.Tn[7].n0 XThC.Tn[7].t4 26.5955
R22701 XThC.Tn[7].n0 XThC.Tn[7].t7 26.5955
R22702 XThC.Tn[7].n1 XThC.Tn[7].t6 26.5955
R22703 XThC.Tn[7].n1 XThC.Tn[7].t5 26.5955
R22704 XThC.Tn[7] XThC.Tn[7].n2 26.5002
R22705 XThC.Tn[7].n53 XThC.Tn[7].t2 24.9236
R22706 XThC.Tn[7].n53 XThC.Tn[7].t1 24.9236
R22707 XThC.Tn[7].n54 XThC.Tn[7].t0 24.9236
R22708 XThC.Tn[7].n54 XThC.Tn[7].t3 24.9236
R22709 XThC.Tn[7].n56 XThC.Tn[7].n55 12.0894
R22710 XThC.Tn[7].n56 XThC.Tn[7] 9.64206
R22711 XThC.Tn[7].n52 XThC.Tn[7] 8.14595
R22712 XThC.Tn[7].n52 XThC.Tn[7].n51 3.36239
R22713 XThC.Tn[7] XThC.Tn[7].n52 3.15894
R22714 XThC.Tn[7].n51 XThC.Tn[7] 2.07622
R22715 XThC.Tn[7] XThC.Tn[7].n56 1.66284
R22716 XThC.Tn[7].n8 XThC.Tn[7] 0.931056
R22717 XThC.Tn[7].n11 XThC.Tn[7] 0.931056
R22718 XThC.Tn[7].n14 XThC.Tn[7] 0.931056
R22719 XThC.Tn[7].n17 XThC.Tn[7] 0.931056
R22720 XThC.Tn[7].n20 XThC.Tn[7] 0.931056
R22721 XThC.Tn[7].n23 XThC.Tn[7] 0.931056
R22722 XThC.Tn[7].n26 XThC.Tn[7] 0.931056
R22723 XThC.Tn[7].n29 XThC.Tn[7] 0.931056
R22724 XThC.Tn[7].n32 XThC.Tn[7] 0.931056
R22725 XThC.Tn[7].n35 XThC.Tn[7] 0.931056
R22726 XThC.Tn[7].n38 XThC.Tn[7] 0.931056
R22727 XThC.Tn[7].n41 XThC.Tn[7] 0.931056
R22728 XThC.Tn[7].n44 XThC.Tn[7] 0.931056
R22729 XThC.Tn[7].n47 XThC.Tn[7] 0.931056
R22730 XThC.Tn[7].n50 XThC.Tn[7] 0.931056
R22731 XThC.Tn[7] XThC.Tn[7].n5 0.396333
R22732 XThC.Tn[7] XThC.Tn[7].n8 0.396333
R22733 XThC.Tn[7] XThC.Tn[7].n11 0.396333
R22734 XThC.Tn[7] XThC.Tn[7].n14 0.396333
R22735 XThC.Tn[7] XThC.Tn[7].n17 0.396333
R22736 XThC.Tn[7] XThC.Tn[7].n20 0.396333
R22737 XThC.Tn[7] XThC.Tn[7].n23 0.396333
R22738 XThC.Tn[7] XThC.Tn[7].n26 0.396333
R22739 XThC.Tn[7] XThC.Tn[7].n29 0.396333
R22740 XThC.Tn[7] XThC.Tn[7].n32 0.396333
R22741 XThC.Tn[7] XThC.Tn[7].n35 0.396333
R22742 XThC.Tn[7] XThC.Tn[7].n38 0.396333
R22743 XThC.Tn[7] XThC.Tn[7].n41 0.396333
R22744 XThC.Tn[7] XThC.Tn[7].n44 0.396333
R22745 XThC.Tn[7] XThC.Tn[7].n47 0.396333
R22746 XThC.Tn[7] XThC.Tn[7].n50 0.396333
R22747 XThC.Tn[7].n4 XThC.Tn[7] 0.104667
R22748 XThC.Tn[7].n7 XThC.Tn[7] 0.104667
R22749 XThC.Tn[7].n10 XThC.Tn[7] 0.104667
R22750 XThC.Tn[7].n13 XThC.Tn[7] 0.104667
R22751 XThC.Tn[7].n16 XThC.Tn[7] 0.104667
R22752 XThC.Tn[7].n19 XThC.Tn[7] 0.104667
R22753 XThC.Tn[7].n22 XThC.Tn[7] 0.104667
R22754 XThC.Tn[7].n25 XThC.Tn[7] 0.104667
R22755 XThC.Tn[7].n28 XThC.Tn[7] 0.104667
R22756 XThC.Tn[7].n31 XThC.Tn[7] 0.104667
R22757 XThC.Tn[7].n34 XThC.Tn[7] 0.104667
R22758 XThC.Tn[7].n37 XThC.Tn[7] 0.104667
R22759 XThC.Tn[7].n40 XThC.Tn[7] 0.104667
R22760 XThC.Tn[7].n43 XThC.Tn[7] 0.104667
R22761 XThC.Tn[7].n46 XThC.Tn[7] 0.104667
R22762 XThC.Tn[7].n49 XThC.Tn[7] 0.104667
R22763 XThC.Tn[7].n4 XThC.Tn[7] 0.0309878
R22764 XThC.Tn[7].n7 XThC.Tn[7] 0.0309878
R22765 XThC.Tn[7].n10 XThC.Tn[7] 0.0309878
R22766 XThC.Tn[7].n13 XThC.Tn[7] 0.0309878
R22767 XThC.Tn[7].n16 XThC.Tn[7] 0.0309878
R22768 XThC.Tn[7].n19 XThC.Tn[7] 0.0309878
R22769 XThC.Tn[7].n22 XThC.Tn[7] 0.0309878
R22770 XThC.Tn[7].n25 XThC.Tn[7] 0.0309878
R22771 XThC.Tn[7].n28 XThC.Tn[7] 0.0309878
R22772 XThC.Tn[7].n31 XThC.Tn[7] 0.0309878
R22773 XThC.Tn[7].n34 XThC.Tn[7] 0.0309878
R22774 XThC.Tn[7].n37 XThC.Tn[7] 0.0309878
R22775 XThC.Tn[7].n40 XThC.Tn[7] 0.0309878
R22776 XThC.Tn[7].n43 XThC.Tn[7] 0.0309878
R22777 XThC.Tn[7].n46 XThC.Tn[7] 0.0309878
R22778 XThC.Tn[7].n49 XThC.Tn[7] 0.0309878
R22779 XThC.Tn[7].n5 XThC.Tn[7].n4 0.027939
R22780 XThC.Tn[7].n8 XThC.Tn[7].n7 0.027939
R22781 XThC.Tn[7].n11 XThC.Tn[7].n10 0.027939
R22782 XThC.Tn[7].n14 XThC.Tn[7].n13 0.027939
R22783 XThC.Tn[7].n17 XThC.Tn[7].n16 0.027939
R22784 XThC.Tn[7].n20 XThC.Tn[7].n19 0.027939
R22785 XThC.Tn[7].n23 XThC.Tn[7].n22 0.027939
R22786 XThC.Tn[7].n26 XThC.Tn[7].n25 0.027939
R22787 XThC.Tn[7].n29 XThC.Tn[7].n28 0.027939
R22788 XThC.Tn[7].n32 XThC.Tn[7].n31 0.027939
R22789 XThC.Tn[7].n35 XThC.Tn[7].n34 0.027939
R22790 XThC.Tn[7].n38 XThC.Tn[7].n37 0.027939
R22791 XThC.Tn[7].n41 XThC.Tn[7].n40 0.027939
R22792 XThC.Tn[7].n44 XThC.Tn[7].n43 0.027939
R22793 XThC.Tn[7].n47 XThC.Tn[7].n46 0.027939
R22794 XThC.Tn[7].n50 XThC.Tn[7].n49 0.027939
R22795 XThC.Tn[7].n51 XThC.Tn[7] 0.00240908
R22796 XThR.Tn[4].n2 XThR.Tn[4].n1 332.334
R22797 XThR.Tn[4].n2 XThR.Tn[4].n0 296.493
R22798 XThR.Tn[4] XThR.Tn[4].n82 161.363
R22799 XThR.Tn[4] XThR.Tn[4].n77 161.363
R22800 XThR.Tn[4] XThR.Tn[4].n72 161.363
R22801 XThR.Tn[4] XThR.Tn[4].n67 161.363
R22802 XThR.Tn[4] XThR.Tn[4].n62 161.363
R22803 XThR.Tn[4] XThR.Tn[4].n57 161.363
R22804 XThR.Tn[4] XThR.Tn[4].n52 161.363
R22805 XThR.Tn[4] XThR.Tn[4].n47 161.363
R22806 XThR.Tn[4] XThR.Tn[4].n42 161.363
R22807 XThR.Tn[4] XThR.Tn[4].n37 161.363
R22808 XThR.Tn[4] XThR.Tn[4].n32 161.363
R22809 XThR.Tn[4] XThR.Tn[4].n27 161.363
R22810 XThR.Tn[4] XThR.Tn[4].n22 161.363
R22811 XThR.Tn[4] XThR.Tn[4].n17 161.363
R22812 XThR.Tn[4] XThR.Tn[4].n12 161.363
R22813 XThR.Tn[4] XThR.Tn[4].n10 161.363
R22814 XThR.Tn[4].n84 XThR.Tn[4].n83 161.3
R22815 XThR.Tn[4].n79 XThR.Tn[4].n78 161.3
R22816 XThR.Tn[4].n74 XThR.Tn[4].n73 161.3
R22817 XThR.Tn[4].n69 XThR.Tn[4].n68 161.3
R22818 XThR.Tn[4].n64 XThR.Tn[4].n63 161.3
R22819 XThR.Tn[4].n59 XThR.Tn[4].n58 161.3
R22820 XThR.Tn[4].n54 XThR.Tn[4].n53 161.3
R22821 XThR.Tn[4].n49 XThR.Tn[4].n48 161.3
R22822 XThR.Tn[4].n44 XThR.Tn[4].n43 161.3
R22823 XThR.Tn[4].n39 XThR.Tn[4].n38 161.3
R22824 XThR.Tn[4].n34 XThR.Tn[4].n33 161.3
R22825 XThR.Tn[4].n29 XThR.Tn[4].n28 161.3
R22826 XThR.Tn[4].n24 XThR.Tn[4].n23 161.3
R22827 XThR.Tn[4].n19 XThR.Tn[4].n18 161.3
R22828 XThR.Tn[4].n14 XThR.Tn[4].n13 161.3
R22829 XThR.Tn[4].n82 XThR.Tn[4].t28 161.106
R22830 XThR.Tn[4].n77 XThR.Tn[4].t34 161.106
R22831 XThR.Tn[4].n72 XThR.Tn[4].t14 161.106
R22832 XThR.Tn[4].n67 XThR.Tn[4].t62 161.106
R22833 XThR.Tn[4].n62 XThR.Tn[4].t26 161.106
R22834 XThR.Tn[4].n57 XThR.Tn[4].t51 161.106
R22835 XThR.Tn[4].n52 XThR.Tn[4].t32 161.106
R22836 XThR.Tn[4].n47 XThR.Tn[4].t12 161.106
R22837 XThR.Tn[4].n42 XThR.Tn[4].t61 161.106
R22838 XThR.Tn[4].n37 XThR.Tn[4].t66 161.106
R22839 XThR.Tn[4].n32 XThR.Tn[4].t49 161.106
R22840 XThR.Tn[4].n27 XThR.Tn[4].t13 161.106
R22841 XThR.Tn[4].n22 XThR.Tn[4].t48 161.106
R22842 XThR.Tn[4].n17 XThR.Tn[4].t31 161.106
R22843 XThR.Tn[4].n12 XThR.Tn[4].t54 161.106
R22844 XThR.Tn[4].n10 XThR.Tn[4].t38 161.106
R22845 XThR.Tn[4].n83 XThR.Tn[4].t24 159.978
R22846 XThR.Tn[4].n78 XThR.Tn[4].t30 159.978
R22847 XThR.Tn[4].n73 XThR.Tn[4].t72 159.978
R22848 XThR.Tn[4].n68 XThR.Tn[4].t59 159.978
R22849 XThR.Tn[4].n63 XThR.Tn[4].t21 159.978
R22850 XThR.Tn[4].n58 XThR.Tn[4].t47 159.978
R22851 XThR.Tn[4].n53 XThR.Tn[4].t29 159.978
R22852 XThR.Tn[4].n48 XThR.Tn[4].t69 159.978
R22853 XThR.Tn[4].n43 XThR.Tn[4].t56 159.978
R22854 XThR.Tn[4].n38 XThR.Tn[4].t63 159.978
R22855 XThR.Tn[4].n33 XThR.Tn[4].t46 159.978
R22856 XThR.Tn[4].n28 XThR.Tn[4].t71 159.978
R22857 XThR.Tn[4].n23 XThR.Tn[4].t45 159.978
R22858 XThR.Tn[4].n18 XThR.Tn[4].t27 159.978
R22859 XThR.Tn[4].n13 XThR.Tn[4].t50 159.978
R22860 XThR.Tn[4].n82 XThR.Tn[4].t16 145.038
R22861 XThR.Tn[4].n77 XThR.Tn[4].t40 145.038
R22862 XThR.Tn[4].n72 XThR.Tn[4].t20 145.038
R22863 XThR.Tn[4].n67 XThR.Tn[4].t67 145.038
R22864 XThR.Tn[4].n62 XThR.Tn[4].t35 145.038
R22865 XThR.Tn[4].n57 XThR.Tn[4].t15 145.038
R22866 XThR.Tn[4].n52 XThR.Tn[4].t22 145.038
R22867 XThR.Tn[4].n47 XThR.Tn[4].t68 145.038
R22868 XThR.Tn[4].n42 XThR.Tn[4].t64 145.038
R22869 XThR.Tn[4].n37 XThR.Tn[4].t33 145.038
R22870 XThR.Tn[4].n32 XThR.Tn[4].t57 145.038
R22871 XThR.Tn[4].n27 XThR.Tn[4].t17 145.038
R22872 XThR.Tn[4].n22 XThR.Tn[4].t55 145.038
R22873 XThR.Tn[4].n17 XThR.Tn[4].t39 145.038
R22874 XThR.Tn[4].n12 XThR.Tn[4].t65 145.038
R22875 XThR.Tn[4].n10 XThR.Tn[4].t44 145.038
R22876 XThR.Tn[4].n83 XThR.Tn[4].t37 143.911
R22877 XThR.Tn[4].n78 XThR.Tn[4].t60 143.911
R22878 XThR.Tn[4].n73 XThR.Tn[4].t42 143.911
R22879 XThR.Tn[4].n68 XThR.Tn[4].t23 143.911
R22880 XThR.Tn[4].n63 XThR.Tn[4].t53 143.911
R22881 XThR.Tn[4].n58 XThR.Tn[4].t36 143.911
R22882 XThR.Tn[4].n53 XThR.Tn[4].t43 143.911
R22883 XThR.Tn[4].n48 XThR.Tn[4].t25 143.911
R22884 XThR.Tn[4].n43 XThR.Tn[4].t18 143.911
R22885 XThR.Tn[4].n38 XThR.Tn[4].t52 143.911
R22886 XThR.Tn[4].n33 XThR.Tn[4].t73 143.911
R22887 XThR.Tn[4].n28 XThR.Tn[4].t41 143.911
R22888 XThR.Tn[4].n23 XThR.Tn[4].t70 143.911
R22889 XThR.Tn[4].n18 XThR.Tn[4].t58 143.911
R22890 XThR.Tn[4].n13 XThR.Tn[4].t19 143.911
R22891 XThR.Tn[4].n5 XThR.Tn[4].n3 135.249
R22892 XThR.Tn[4].n5 XThR.Tn[4].n4 98.982
R22893 XThR.Tn[4].n7 XThR.Tn[4].n6 98.982
R22894 XThR.Tn[4].n9 XThR.Tn[4].n8 98.982
R22895 XThR.Tn[4].n7 XThR.Tn[4].n5 36.2672
R22896 XThR.Tn[4].n9 XThR.Tn[4].n7 36.2672
R22897 XThR.Tn[4].n88 XThR.Tn[4].n9 32.6405
R22898 XThR.Tn[4].n0 XThR.Tn[4].t1 26.5955
R22899 XThR.Tn[4].n0 XThR.Tn[4].t2 26.5955
R22900 XThR.Tn[4].n1 XThR.Tn[4].t0 26.5955
R22901 XThR.Tn[4].n1 XThR.Tn[4].t3 26.5955
R22902 XThR.Tn[4].n3 XThR.Tn[4].t8 24.9236
R22903 XThR.Tn[4].n3 XThR.Tn[4].t9 24.9236
R22904 XThR.Tn[4].n4 XThR.Tn[4].t11 24.9236
R22905 XThR.Tn[4].n4 XThR.Tn[4].t10 24.9236
R22906 XThR.Tn[4].n6 XThR.Tn[4].t6 24.9236
R22907 XThR.Tn[4].n6 XThR.Tn[4].t5 24.9236
R22908 XThR.Tn[4].n8 XThR.Tn[4].t7 24.9236
R22909 XThR.Tn[4].n8 XThR.Tn[4].t4 24.9236
R22910 XThR.Tn[4] XThR.Tn[4].n2 23.3605
R22911 XThR.Tn[4] XThR.Tn[4].n88 6.7205
R22912 XThR.Tn[4].n88 XThR.Tn[4] 5.80883
R22913 XThR.Tn[4] XThR.Tn[4].n11 5.34038
R22914 XThR.Tn[4].n16 XThR.Tn[4].n15 4.5005
R22915 XThR.Tn[4].n21 XThR.Tn[4].n20 4.5005
R22916 XThR.Tn[4].n26 XThR.Tn[4].n25 4.5005
R22917 XThR.Tn[4].n31 XThR.Tn[4].n30 4.5005
R22918 XThR.Tn[4].n36 XThR.Tn[4].n35 4.5005
R22919 XThR.Tn[4].n41 XThR.Tn[4].n40 4.5005
R22920 XThR.Tn[4].n46 XThR.Tn[4].n45 4.5005
R22921 XThR.Tn[4].n51 XThR.Tn[4].n50 4.5005
R22922 XThR.Tn[4].n56 XThR.Tn[4].n55 4.5005
R22923 XThR.Tn[4].n61 XThR.Tn[4].n60 4.5005
R22924 XThR.Tn[4].n66 XThR.Tn[4].n65 4.5005
R22925 XThR.Tn[4].n71 XThR.Tn[4].n70 4.5005
R22926 XThR.Tn[4].n76 XThR.Tn[4].n75 4.5005
R22927 XThR.Tn[4].n81 XThR.Tn[4].n80 4.5005
R22928 XThR.Tn[4].n86 XThR.Tn[4].n85 4.5005
R22929 XThR.Tn[4].n87 XThR.Tn[4] 3.70586
R22930 XThR.Tn[4].n16 XThR.Tn[4] 2.52282
R22931 XThR.Tn[4].n21 XThR.Tn[4] 2.52282
R22932 XThR.Tn[4].n26 XThR.Tn[4] 2.52282
R22933 XThR.Tn[4].n31 XThR.Tn[4] 2.52282
R22934 XThR.Tn[4].n36 XThR.Tn[4] 2.52282
R22935 XThR.Tn[4].n41 XThR.Tn[4] 2.52282
R22936 XThR.Tn[4].n46 XThR.Tn[4] 2.52282
R22937 XThR.Tn[4].n51 XThR.Tn[4] 2.52282
R22938 XThR.Tn[4].n56 XThR.Tn[4] 2.52282
R22939 XThR.Tn[4].n61 XThR.Tn[4] 2.52282
R22940 XThR.Tn[4].n66 XThR.Tn[4] 2.52282
R22941 XThR.Tn[4].n71 XThR.Tn[4] 2.52282
R22942 XThR.Tn[4].n76 XThR.Tn[4] 2.52282
R22943 XThR.Tn[4].n81 XThR.Tn[4] 2.52282
R22944 XThR.Tn[4].n86 XThR.Tn[4] 2.52282
R22945 XThR.Tn[4].n84 XThR.Tn[4] 1.08677
R22946 XThR.Tn[4].n79 XThR.Tn[4] 1.08677
R22947 XThR.Tn[4].n74 XThR.Tn[4] 1.08677
R22948 XThR.Tn[4].n69 XThR.Tn[4] 1.08677
R22949 XThR.Tn[4].n64 XThR.Tn[4] 1.08677
R22950 XThR.Tn[4].n59 XThR.Tn[4] 1.08677
R22951 XThR.Tn[4].n54 XThR.Tn[4] 1.08677
R22952 XThR.Tn[4].n49 XThR.Tn[4] 1.08677
R22953 XThR.Tn[4].n44 XThR.Tn[4] 1.08677
R22954 XThR.Tn[4].n39 XThR.Tn[4] 1.08677
R22955 XThR.Tn[4].n34 XThR.Tn[4] 1.08677
R22956 XThR.Tn[4].n29 XThR.Tn[4] 1.08677
R22957 XThR.Tn[4].n24 XThR.Tn[4] 1.08677
R22958 XThR.Tn[4].n19 XThR.Tn[4] 1.08677
R22959 XThR.Tn[4].n14 XThR.Tn[4] 1.08677
R22960 XThR.Tn[4] XThR.Tn[4].n16 0.839786
R22961 XThR.Tn[4] XThR.Tn[4].n21 0.839786
R22962 XThR.Tn[4] XThR.Tn[4].n26 0.839786
R22963 XThR.Tn[4] XThR.Tn[4].n31 0.839786
R22964 XThR.Tn[4] XThR.Tn[4].n36 0.839786
R22965 XThR.Tn[4] XThR.Tn[4].n41 0.839786
R22966 XThR.Tn[4] XThR.Tn[4].n46 0.839786
R22967 XThR.Tn[4] XThR.Tn[4].n51 0.839786
R22968 XThR.Tn[4] XThR.Tn[4].n56 0.839786
R22969 XThR.Tn[4] XThR.Tn[4].n61 0.839786
R22970 XThR.Tn[4] XThR.Tn[4].n66 0.839786
R22971 XThR.Tn[4] XThR.Tn[4].n71 0.839786
R22972 XThR.Tn[4] XThR.Tn[4].n76 0.839786
R22973 XThR.Tn[4] XThR.Tn[4].n81 0.839786
R22974 XThR.Tn[4] XThR.Tn[4].n86 0.839786
R22975 XThR.Tn[4].n11 XThR.Tn[4] 0.499542
R22976 XThR.Tn[4].n85 XThR.Tn[4] 0.063
R22977 XThR.Tn[4].n80 XThR.Tn[4] 0.063
R22978 XThR.Tn[4].n75 XThR.Tn[4] 0.063
R22979 XThR.Tn[4].n70 XThR.Tn[4] 0.063
R22980 XThR.Tn[4].n65 XThR.Tn[4] 0.063
R22981 XThR.Tn[4].n60 XThR.Tn[4] 0.063
R22982 XThR.Tn[4].n55 XThR.Tn[4] 0.063
R22983 XThR.Tn[4].n50 XThR.Tn[4] 0.063
R22984 XThR.Tn[4].n45 XThR.Tn[4] 0.063
R22985 XThR.Tn[4].n40 XThR.Tn[4] 0.063
R22986 XThR.Tn[4].n35 XThR.Tn[4] 0.063
R22987 XThR.Tn[4].n30 XThR.Tn[4] 0.063
R22988 XThR.Tn[4].n25 XThR.Tn[4] 0.063
R22989 XThR.Tn[4].n20 XThR.Tn[4] 0.063
R22990 XThR.Tn[4].n15 XThR.Tn[4] 0.063
R22991 XThR.Tn[4].n87 XThR.Tn[4] 0.0540714
R22992 XThR.Tn[4] XThR.Tn[4].n87 0.038
R22993 XThR.Tn[4].n11 XThR.Tn[4] 0.0143889
R22994 XThR.Tn[4].n85 XThR.Tn[4].n84 0.00771154
R22995 XThR.Tn[4].n80 XThR.Tn[4].n79 0.00771154
R22996 XThR.Tn[4].n75 XThR.Tn[4].n74 0.00771154
R22997 XThR.Tn[4].n70 XThR.Tn[4].n69 0.00771154
R22998 XThR.Tn[4].n65 XThR.Tn[4].n64 0.00771154
R22999 XThR.Tn[4].n60 XThR.Tn[4].n59 0.00771154
R23000 XThR.Tn[4].n55 XThR.Tn[4].n54 0.00771154
R23001 XThR.Tn[4].n50 XThR.Tn[4].n49 0.00771154
R23002 XThR.Tn[4].n45 XThR.Tn[4].n44 0.00771154
R23003 XThR.Tn[4].n40 XThR.Tn[4].n39 0.00771154
R23004 XThR.Tn[4].n35 XThR.Tn[4].n34 0.00771154
R23005 XThR.Tn[4].n30 XThR.Tn[4].n29 0.00771154
R23006 XThR.Tn[4].n25 XThR.Tn[4].n24 0.00771154
R23007 XThR.Tn[4].n20 XThR.Tn[4].n19 0.00771154
R23008 XThR.Tn[4].n15 XThR.Tn[4].n14 0.00771154
R23009 XThR.Tn[11].n8 XThR.Tn[11].n7 256.104
R23010 XThR.Tn[11].n5 XThR.Tn[11].n3 243.68
R23011 XThR.Tn[11].n2 XThR.Tn[11].n1 241.847
R23012 XThR.Tn[11].n5 XThR.Tn[11].n4 205.28
R23013 XThR.Tn[11].n8 XThR.Tn[11].n6 202.094
R23014 XThR.Tn[11].n2 XThR.Tn[11].n0 185
R23015 XThR.Tn[11] XThR.Tn[11].n82 161.363
R23016 XThR.Tn[11] XThR.Tn[11].n77 161.363
R23017 XThR.Tn[11] XThR.Tn[11].n72 161.363
R23018 XThR.Tn[11] XThR.Tn[11].n67 161.363
R23019 XThR.Tn[11] XThR.Tn[11].n62 161.363
R23020 XThR.Tn[11] XThR.Tn[11].n57 161.363
R23021 XThR.Tn[11] XThR.Tn[11].n52 161.363
R23022 XThR.Tn[11] XThR.Tn[11].n47 161.363
R23023 XThR.Tn[11] XThR.Tn[11].n42 161.363
R23024 XThR.Tn[11] XThR.Tn[11].n37 161.363
R23025 XThR.Tn[11] XThR.Tn[11].n32 161.363
R23026 XThR.Tn[11] XThR.Tn[11].n27 161.363
R23027 XThR.Tn[11] XThR.Tn[11].n22 161.363
R23028 XThR.Tn[11] XThR.Tn[11].n17 161.363
R23029 XThR.Tn[11] XThR.Tn[11].n12 161.363
R23030 XThR.Tn[11] XThR.Tn[11].n10 161.363
R23031 XThR.Tn[11].n84 XThR.Tn[11].n83 161.3
R23032 XThR.Tn[11].n79 XThR.Tn[11].n78 161.3
R23033 XThR.Tn[11].n74 XThR.Tn[11].n73 161.3
R23034 XThR.Tn[11].n69 XThR.Tn[11].n68 161.3
R23035 XThR.Tn[11].n64 XThR.Tn[11].n63 161.3
R23036 XThR.Tn[11].n59 XThR.Tn[11].n58 161.3
R23037 XThR.Tn[11].n54 XThR.Tn[11].n53 161.3
R23038 XThR.Tn[11].n49 XThR.Tn[11].n48 161.3
R23039 XThR.Tn[11].n44 XThR.Tn[11].n43 161.3
R23040 XThR.Tn[11].n39 XThR.Tn[11].n38 161.3
R23041 XThR.Tn[11].n34 XThR.Tn[11].n33 161.3
R23042 XThR.Tn[11].n29 XThR.Tn[11].n28 161.3
R23043 XThR.Tn[11].n24 XThR.Tn[11].n23 161.3
R23044 XThR.Tn[11].n19 XThR.Tn[11].n18 161.3
R23045 XThR.Tn[11].n14 XThR.Tn[11].n13 161.3
R23046 XThR.Tn[11].n82 XThR.Tn[11].t40 161.106
R23047 XThR.Tn[11].n77 XThR.Tn[11].t46 161.106
R23048 XThR.Tn[11].n72 XThR.Tn[11].t24 161.106
R23049 XThR.Tn[11].n67 XThR.Tn[11].t73 161.106
R23050 XThR.Tn[11].n62 XThR.Tn[11].t39 161.106
R23051 XThR.Tn[11].n57 XThR.Tn[11].t63 161.106
R23052 XThR.Tn[11].n52 XThR.Tn[11].t43 161.106
R23053 XThR.Tn[11].n47 XThR.Tn[11].t22 161.106
R23054 XThR.Tn[11].n42 XThR.Tn[11].t71 161.106
R23055 XThR.Tn[11].n37 XThR.Tn[11].t14 161.106
R23056 XThR.Tn[11].n32 XThR.Tn[11].t62 161.106
R23057 XThR.Tn[11].n27 XThR.Tn[11].t23 161.106
R23058 XThR.Tn[11].n22 XThR.Tn[11].t60 161.106
R23059 XThR.Tn[11].n17 XThR.Tn[11].t41 161.106
R23060 XThR.Tn[11].n12 XThR.Tn[11].t67 161.106
R23061 XThR.Tn[11].n10 XThR.Tn[11].t48 161.106
R23062 XThR.Tn[11].n83 XThR.Tn[11].t31 159.978
R23063 XThR.Tn[11].n78 XThR.Tn[11].t38 159.978
R23064 XThR.Tn[11].n73 XThR.Tn[11].t20 159.978
R23065 XThR.Tn[11].n68 XThR.Tn[11].t66 159.978
R23066 XThR.Tn[11].n63 XThR.Tn[11].t29 159.978
R23067 XThR.Tn[11].n58 XThR.Tn[11].t57 159.978
R23068 XThR.Tn[11].n53 XThR.Tn[11].t37 159.978
R23069 XThR.Tn[11].n48 XThR.Tn[11].t17 159.978
R23070 XThR.Tn[11].n43 XThR.Tn[11].t64 159.978
R23071 XThR.Tn[11].n38 XThR.Tn[11].t72 159.978
R23072 XThR.Tn[11].n33 XThR.Tn[11].t55 159.978
R23073 XThR.Tn[11].n28 XThR.Tn[11].t19 159.978
R23074 XThR.Tn[11].n23 XThR.Tn[11].t54 159.978
R23075 XThR.Tn[11].n18 XThR.Tn[11].t36 159.978
R23076 XThR.Tn[11].n13 XThR.Tn[11].t58 159.978
R23077 XThR.Tn[11].n82 XThR.Tn[11].t26 145.038
R23078 XThR.Tn[11].n77 XThR.Tn[11].t53 145.038
R23079 XThR.Tn[11].n72 XThR.Tn[11].t34 145.038
R23080 XThR.Tn[11].n67 XThR.Tn[11].t15 145.038
R23081 XThR.Tn[11].n62 XThR.Tn[11].t47 145.038
R23082 XThR.Tn[11].n57 XThR.Tn[11].t25 145.038
R23083 XThR.Tn[11].n52 XThR.Tn[11].t35 145.038
R23084 XThR.Tn[11].n47 XThR.Tn[11].t16 145.038
R23085 XThR.Tn[11].n42 XThR.Tn[11].t13 145.038
R23086 XThR.Tn[11].n37 XThR.Tn[11].t44 145.038
R23087 XThR.Tn[11].n32 XThR.Tn[11].t70 145.038
R23088 XThR.Tn[11].n27 XThR.Tn[11].t33 145.038
R23089 XThR.Tn[11].n22 XThR.Tn[11].t68 145.038
R23090 XThR.Tn[11].n17 XThR.Tn[11].t49 145.038
R23091 XThR.Tn[11].n12 XThR.Tn[11].t12 145.038
R23092 XThR.Tn[11].n10 XThR.Tn[11].t56 145.038
R23093 XThR.Tn[11].n83 XThR.Tn[11].t45 143.911
R23094 XThR.Tn[11].n78 XThR.Tn[11].t69 143.911
R23095 XThR.Tn[11].n73 XThR.Tn[11].t51 143.911
R23096 XThR.Tn[11].n68 XThR.Tn[11].t30 143.911
R23097 XThR.Tn[11].n63 XThR.Tn[11].t61 143.911
R23098 XThR.Tn[11].n58 XThR.Tn[11].t42 143.911
R23099 XThR.Tn[11].n53 XThR.Tn[11].t52 143.911
R23100 XThR.Tn[11].n48 XThR.Tn[11].t32 143.911
R23101 XThR.Tn[11].n43 XThR.Tn[11].t28 143.911
R23102 XThR.Tn[11].n38 XThR.Tn[11].t59 143.911
R23103 XThR.Tn[11].n33 XThR.Tn[11].t21 143.911
R23104 XThR.Tn[11].n28 XThR.Tn[11].t50 143.911
R23105 XThR.Tn[11].n23 XThR.Tn[11].t18 143.911
R23106 XThR.Tn[11].n18 XThR.Tn[11].t65 143.911
R23107 XThR.Tn[11].n13 XThR.Tn[11].t27 143.911
R23108 XThR.Tn[11] XThR.Tn[11].n5 35.7652
R23109 XThR.Tn[11].n6 XThR.Tn[11].t4 26.5955
R23110 XThR.Tn[11].n6 XThR.Tn[11].t6 26.5955
R23111 XThR.Tn[11].n7 XThR.Tn[11].t5 26.5955
R23112 XThR.Tn[11].n7 XThR.Tn[11].t7 26.5955
R23113 XThR.Tn[11].n3 XThR.Tn[11].t8 26.5955
R23114 XThR.Tn[11].n3 XThR.Tn[11].t10 26.5955
R23115 XThR.Tn[11].n4 XThR.Tn[11].t9 26.5955
R23116 XThR.Tn[11].n4 XThR.Tn[11].t11 26.5955
R23117 XThR.Tn[11].n0 XThR.Tn[11].t2 24.9236
R23118 XThR.Tn[11].n0 XThR.Tn[11].t0 24.9236
R23119 XThR.Tn[11].n1 XThR.Tn[11].t3 24.9236
R23120 XThR.Tn[11].n1 XThR.Tn[11].t1 24.9236
R23121 XThR.Tn[11] XThR.Tn[11].n2 22.9615
R23122 XThR.Tn[11].n9 XThR.Tn[11].n8 13.5534
R23123 XThR.Tn[11].n88 XThR.Tn[11] 8.41462
R23124 XThR.Tn[11] XThR.Tn[11].n11 5.34038
R23125 XThR.Tn[11].n16 XThR.Tn[11].n15 4.5005
R23126 XThR.Tn[11].n21 XThR.Tn[11].n20 4.5005
R23127 XThR.Tn[11].n26 XThR.Tn[11].n25 4.5005
R23128 XThR.Tn[11].n31 XThR.Tn[11].n30 4.5005
R23129 XThR.Tn[11].n36 XThR.Tn[11].n35 4.5005
R23130 XThR.Tn[11].n41 XThR.Tn[11].n40 4.5005
R23131 XThR.Tn[11].n46 XThR.Tn[11].n45 4.5005
R23132 XThR.Tn[11].n51 XThR.Tn[11].n50 4.5005
R23133 XThR.Tn[11].n56 XThR.Tn[11].n55 4.5005
R23134 XThR.Tn[11].n61 XThR.Tn[11].n60 4.5005
R23135 XThR.Tn[11].n66 XThR.Tn[11].n65 4.5005
R23136 XThR.Tn[11].n71 XThR.Tn[11].n70 4.5005
R23137 XThR.Tn[11].n76 XThR.Tn[11].n75 4.5005
R23138 XThR.Tn[11].n81 XThR.Tn[11].n80 4.5005
R23139 XThR.Tn[11].n86 XThR.Tn[11].n85 4.5005
R23140 XThR.Tn[11].n87 XThR.Tn[11] 3.70586
R23141 XThR.Tn[11].n88 XThR.Tn[11].n9 2.99115
R23142 XThR.Tn[11].n9 XThR.Tn[11] 2.87153
R23143 XThR.Tn[11].n16 XThR.Tn[11] 2.52282
R23144 XThR.Tn[11].n21 XThR.Tn[11] 2.52282
R23145 XThR.Tn[11].n26 XThR.Tn[11] 2.52282
R23146 XThR.Tn[11].n31 XThR.Tn[11] 2.52282
R23147 XThR.Tn[11].n36 XThR.Tn[11] 2.52282
R23148 XThR.Tn[11].n41 XThR.Tn[11] 2.52282
R23149 XThR.Tn[11].n46 XThR.Tn[11] 2.52282
R23150 XThR.Tn[11].n51 XThR.Tn[11] 2.52282
R23151 XThR.Tn[11].n56 XThR.Tn[11] 2.52282
R23152 XThR.Tn[11].n61 XThR.Tn[11] 2.52282
R23153 XThR.Tn[11].n66 XThR.Tn[11] 2.52282
R23154 XThR.Tn[11].n71 XThR.Tn[11] 2.52282
R23155 XThR.Tn[11].n76 XThR.Tn[11] 2.52282
R23156 XThR.Tn[11].n81 XThR.Tn[11] 2.52282
R23157 XThR.Tn[11].n86 XThR.Tn[11] 2.52282
R23158 XThR.Tn[11] XThR.Tn[11].n88 2.2734
R23159 XThR.Tn[11].n9 XThR.Tn[11] 1.50638
R23160 XThR.Tn[11].n84 XThR.Tn[11] 1.08677
R23161 XThR.Tn[11].n79 XThR.Tn[11] 1.08677
R23162 XThR.Tn[11].n74 XThR.Tn[11] 1.08677
R23163 XThR.Tn[11].n69 XThR.Tn[11] 1.08677
R23164 XThR.Tn[11].n64 XThR.Tn[11] 1.08677
R23165 XThR.Tn[11].n59 XThR.Tn[11] 1.08677
R23166 XThR.Tn[11].n54 XThR.Tn[11] 1.08677
R23167 XThR.Tn[11].n49 XThR.Tn[11] 1.08677
R23168 XThR.Tn[11].n44 XThR.Tn[11] 1.08677
R23169 XThR.Tn[11].n39 XThR.Tn[11] 1.08677
R23170 XThR.Tn[11].n34 XThR.Tn[11] 1.08677
R23171 XThR.Tn[11].n29 XThR.Tn[11] 1.08677
R23172 XThR.Tn[11].n24 XThR.Tn[11] 1.08677
R23173 XThR.Tn[11].n19 XThR.Tn[11] 1.08677
R23174 XThR.Tn[11].n14 XThR.Tn[11] 1.08677
R23175 XThR.Tn[11] XThR.Tn[11].n16 0.839786
R23176 XThR.Tn[11] XThR.Tn[11].n21 0.839786
R23177 XThR.Tn[11] XThR.Tn[11].n26 0.839786
R23178 XThR.Tn[11] XThR.Tn[11].n31 0.839786
R23179 XThR.Tn[11] XThR.Tn[11].n36 0.839786
R23180 XThR.Tn[11] XThR.Tn[11].n41 0.839786
R23181 XThR.Tn[11] XThR.Tn[11].n46 0.839786
R23182 XThR.Tn[11] XThR.Tn[11].n51 0.839786
R23183 XThR.Tn[11] XThR.Tn[11].n56 0.839786
R23184 XThR.Tn[11] XThR.Tn[11].n61 0.839786
R23185 XThR.Tn[11] XThR.Tn[11].n66 0.839786
R23186 XThR.Tn[11] XThR.Tn[11].n71 0.839786
R23187 XThR.Tn[11] XThR.Tn[11].n76 0.839786
R23188 XThR.Tn[11] XThR.Tn[11].n81 0.839786
R23189 XThR.Tn[11] XThR.Tn[11].n86 0.839786
R23190 XThR.Tn[11].n11 XThR.Tn[11] 0.499542
R23191 XThR.Tn[11].n85 XThR.Tn[11] 0.063
R23192 XThR.Tn[11].n80 XThR.Tn[11] 0.063
R23193 XThR.Tn[11].n75 XThR.Tn[11] 0.063
R23194 XThR.Tn[11].n70 XThR.Tn[11] 0.063
R23195 XThR.Tn[11].n65 XThR.Tn[11] 0.063
R23196 XThR.Tn[11].n60 XThR.Tn[11] 0.063
R23197 XThR.Tn[11].n55 XThR.Tn[11] 0.063
R23198 XThR.Tn[11].n50 XThR.Tn[11] 0.063
R23199 XThR.Tn[11].n45 XThR.Tn[11] 0.063
R23200 XThR.Tn[11].n40 XThR.Tn[11] 0.063
R23201 XThR.Tn[11].n35 XThR.Tn[11] 0.063
R23202 XThR.Tn[11].n30 XThR.Tn[11] 0.063
R23203 XThR.Tn[11].n25 XThR.Tn[11] 0.063
R23204 XThR.Tn[11].n20 XThR.Tn[11] 0.063
R23205 XThR.Tn[11].n15 XThR.Tn[11] 0.063
R23206 XThR.Tn[11].n87 XThR.Tn[11] 0.0540714
R23207 XThR.Tn[11] XThR.Tn[11].n87 0.038
R23208 XThR.Tn[11].n11 XThR.Tn[11] 0.0143889
R23209 XThR.Tn[11].n85 XThR.Tn[11].n84 0.00771154
R23210 XThR.Tn[11].n80 XThR.Tn[11].n79 0.00771154
R23211 XThR.Tn[11].n75 XThR.Tn[11].n74 0.00771154
R23212 XThR.Tn[11].n70 XThR.Tn[11].n69 0.00771154
R23213 XThR.Tn[11].n65 XThR.Tn[11].n64 0.00771154
R23214 XThR.Tn[11].n60 XThR.Tn[11].n59 0.00771154
R23215 XThR.Tn[11].n55 XThR.Tn[11].n54 0.00771154
R23216 XThR.Tn[11].n50 XThR.Tn[11].n49 0.00771154
R23217 XThR.Tn[11].n45 XThR.Tn[11].n44 0.00771154
R23218 XThR.Tn[11].n40 XThR.Tn[11].n39 0.00771154
R23219 XThR.Tn[11].n35 XThR.Tn[11].n34 0.00771154
R23220 XThR.Tn[11].n30 XThR.Tn[11].n29 0.00771154
R23221 XThR.Tn[11].n25 XThR.Tn[11].n24 0.00771154
R23222 XThR.Tn[11].n20 XThR.Tn[11].n19 0.00771154
R23223 XThR.Tn[11].n15 XThR.Tn[11].n14 0.00771154
R23224 XThR.Tn[7].n5 XThR.Tn[7].n3 244.069
R23225 XThR.Tn[7].n2 XThR.Tn[7].n1 236.589
R23226 XThR.Tn[7].n5 XThR.Tn[7].n4 204.893
R23227 XThR.Tn[7].n2 XThR.Tn[7].n0 200.321
R23228 XThR.Tn[7] XThR.Tn[7].n79 161.363
R23229 XThR.Tn[7] XThR.Tn[7].n74 161.363
R23230 XThR.Tn[7] XThR.Tn[7].n69 161.363
R23231 XThR.Tn[7] XThR.Tn[7].n64 161.363
R23232 XThR.Tn[7] XThR.Tn[7].n59 161.363
R23233 XThR.Tn[7] XThR.Tn[7].n54 161.363
R23234 XThR.Tn[7] XThR.Tn[7].n49 161.363
R23235 XThR.Tn[7] XThR.Tn[7].n44 161.363
R23236 XThR.Tn[7] XThR.Tn[7].n39 161.363
R23237 XThR.Tn[7] XThR.Tn[7].n34 161.363
R23238 XThR.Tn[7] XThR.Tn[7].n29 161.363
R23239 XThR.Tn[7] XThR.Tn[7].n24 161.363
R23240 XThR.Tn[7] XThR.Tn[7].n19 161.363
R23241 XThR.Tn[7] XThR.Tn[7].n14 161.363
R23242 XThR.Tn[7] XThR.Tn[7].n9 161.363
R23243 XThR.Tn[7] XThR.Tn[7].n7 161.363
R23244 XThR.Tn[7].n81 XThR.Tn[7].n80 161.3
R23245 XThR.Tn[7].n76 XThR.Tn[7].n75 161.3
R23246 XThR.Tn[7].n71 XThR.Tn[7].n70 161.3
R23247 XThR.Tn[7].n66 XThR.Tn[7].n65 161.3
R23248 XThR.Tn[7].n61 XThR.Tn[7].n60 161.3
R23249 XThR.Tn[7].n56 XThR.Tn[7].n55 161.3
R23250 XThR.Tn[7].n51 XThR.Tn[7].n50 161.3
R23251 XThR.Tn[7].n46 XThR.Tn[7].n45 161.3
R23252 XThR.Tn[7].n41 XThR.Tn[7].n40 161.3
R23253 XThR.Tn[7].n36 XThR.Tn[7].n35 161.3
R23254 XThR.Tn[7].n31 XThR.Tn[7].n30 161.3
R23255 XThR.Tn[7].n26 XThR.Tn[7].n25 161.3
R23256 XThR.Tn[7].n21 XThR.Tn[7].n20 161.3
R23257 XThR.Tn[7].n16 XThR.Tn[7].n15 161.3
R23258 XThR.Tn[7].n11 XThR.Tn[7].n10 161.3
R23259 XThR.Tn[7].n79 XThR.Tn[7].t35 161.106
R23260 XThR.Tn[7].n74 XThR.Tn[7].t41 161.106
R23261 XThR.Tn[7].n69 XThR.Tn[7].t22 161.106
R23262 XThR.Tn[7].n64 XThR.Tn[7].t69 161.106
R23263 XThR.Tn[7].n59 XThR.Tn[7].t33 161.106
R23264 XThR.Tn[7].n54 XThR.Tn[7].t57 161.106
R23265 XThR.Tn[7].n49 XThR.Tn[7].t39 161.106
R23266 XThR.Tn[7].n44 XThR.Tn[7].t20 161.106
R23267 XThR.Tn[7].n39 XThR.Tn[7].t68 161.106
R23268 XThR.Tn[7].n34 XThR.Tn[7].t11 161.106
R23269 XThR.Tn[7].n29 XThR.Tn[7].t56 161.106
R23270 XThR.Tn[7].n24 XThR.Tn[7].t21 161.106
R23271 XThR.Tn[7].n19 XThR.Tn[7].t55 161.106
R23272 XThR.Tn[7].n14 XThR.Tn[7].t37 161.106
R23273 XThR.Tn[7].n9 XThR.Tn[7].t60 161.106
R23274 XThR.Tn[7].n7 XThR.Tn[7].t45 161.106
R23275 XThR.Tn[7].n80 XThR.Tn[7].t13 159.978
R23276 XThR.Tn[7].n75 XThR.Tn[7].t17 159.978
R23277 XThR.Tn[7].n70 XThR.Tn[7].t64 159.978
R23278 XThR.Tn[7].n65 XThR.Tn[7].t48 159.978
R23279 XThR.Tn[7].n60 XThR.Tn[7].t10 159.978
R23280 XThR.Tn[7].n55 XThR.Tn[7].t36 159.978
R23281 XThR.Tn[7].n50 XThR.Tn[7].t16 159.978
R23282 XThR.Tn[7].n45 XThR.Tn[7].t61 159.978
R23283 XThR.Tn[7].n40 XThR.Tn[7].t46 159.978
R23284 XThR.Tn[7].n35 XThR.Tn[7].t54 159.978
R23285 XThR.Tn[7].n30 XThR.Tn[7].t34 159.978
R23286 XThR.Tn[7].n25 XThR.Tn[7].t63 159.978
R23287 XThR.Tn[7].n20 XThR.Tn[7].t32 159.978
R23288 XThR.Tn[7].n15 XThR.Tn[7].t15 159.978
R23289 XThR.Tn[7].n10 XThR.Tn[7].t38 159.978
R23290 XThR.Tn[7].n79 XThR.Tn[7].t24 145.038
R23291 XThR.Tn[7].n74 XThR.Tn[7].t49 145.038
R23292 XThR.Tn[7].n69 XThR.Tn[7].t28 145.038
R23293 XThR.Tn[7].n64 XThR.Tn[7].t12 145.038
R23294 XThR.Tn[7].n59 XThR.Tn[7].t42 145.038
R23295 XThR.Tn[7].n54 XThR.Tn[7].t23 145.038
R23296 XThR.Tn[7].n49 XThR.Tn[7].t29 145.038
R23297 XThR.Tn[7].n44 XThR.Tn[7].t14 145.038
R23298 XThR.Tn[7].n39 XThR.Tn[7].t9 145.038
R23299 XThR.Tn[7].n34 XThR.Tn[7].t40 145.038
R23300 XThR.Tn[7].n29 XThR.Tn[7].t65 145.038
R23301 XThR.Tn[7].n24 XThR.Tn[7].t25 145.038
R23302 XThR.Tn[7].n19 XThR.Tn[7].t62 145.038
R23303 XThR.Tn[7].n14 XThR.Tn[7].t47 145.038
R23304 XThR.Tn[7].n9 XThR.Tn[7].t8 145.038
R23305 XThR.Tn[7].n7 XThR.Tn[7].t53 145.038
R23306 XThR.Tn[7].n80 XThR.Tn[7].t44 143.911
R23307 XThR.Tn[7].n75 XThR.Tn[7].t67 143.911
R23308 XThR.Tn[7].n70 XThR.Tn[7].t51 143.911
R23309 XThR.Tn[7].n65 XThR.Tn[7].t30 143.911
R23310 XThR.Tn[7].n60 XThR.Tn[7].t59 143.911
R23311 XThR.Tn[7].n55 XThR.Tn[7].t43 143.911
R23312 XThR.Tn[7].n50 XThR.Tn[7].t52 143.911
R23313 XThR.Tn[7].n45 XThR.Tn[7].t31 143.911
R23314 XThR.Tn[7].n40 XThR.Tn[7].t27 143.911
R23315 XThR.Tn[7].n35 XThR.Tn[7].t58 143.911
R23316 XThR.Tn[7].n30 XThR.Tn[7].t19 143.911
R23317 XThR.Tn[7].n25 XThR.Tn[7].t50 143.911
R23318 XThR.Tn[7].n20 XThR.Tn[7].t18 143.911
R23319 XThR.Tn[7].n15 XThR.Tn[7].t66 143.911
R23320 XThR.Tn[7].n10 XThR.Tn[7].t26 143.911
R23321 XThR.Tn[7].n4 XThR.Tn[7].t5 26.5955
R23322 XThR.Tn[7].n4 XThR.Tn[7].t4 26.5955
R23323 XThR.Tn[7].n3 XThR.Tn[7].t6 26.5955
R23324 XThR.Tn[7].n3 XThR.Tn[7].t7 26.5955
R23325 XThR.Tn[7].n0 XThR.Tn[7].t2 24.9236
R23326 XThR.Tn[7].n0 XThR.Tn[7].t1 24.9236
R23327 XThR.Tn[7].n1 XThR.Tn[7].t3 24.9236
R23328 XThR.Tn[7].n1 XThR.Tn[7].t0 24.9236
R23329 XThR.Tn[7] XThR.Tn[7].n2 16.079
R23330 XThR.Tn[7].n6 XThR.Tn[7].n5 11.4531
R23331 XThR.Tn[7] XThR.Tn[7].n6 10.4732
R23332 XThR.Tn[7] XThR.Tn[7].n85 8.81089
R23333 XThR.Tn[7] XThR.Tn[7].n8 5.34038
R23334 XThR.Tn[7].n85 XThR.Tn[7] 5.25732
R23335 XThR.Tn[7].n13 XThR.Tn[7].n12 4.5005
R23336 XThR.Tn[7].n18 XThR.Tn[7].n17 4.5005
R23337 XThR.Tn[7].n23 XThR.Tn[7].n22 4.5005
R23338 XThR.Tn[7].n28 XThR.Tn[7].n27 4.5005
R23339 XThR.Tn[7].n33 XThR.Tn[7].n32 4.5005
R23340 XThR.Tn[7].n38 XThR.Tn[7].n37 4.5005
R23341 XThR.Tn[7].n43 XThR.Tn[7].n42 4.5005
R23342 XThR.Tn[7].n48 XThR.Tn[7].n47 4.5005
R23343 XThR.Tn[7].n53 XThR.Tn[7].n52 4.5005
R23344 XThR.Tn[7].n58 XThR.Tn[7].n57 4.5005
R23345 XThR.Tn[7].n63 XThR.Tn[7].n62 4.5005
R23346 XThR.Tn[7].n68 XThR.Tn[7].n67 4.5005
R23347 XThR.Tn[7].n73 XThR.Tn[7].n72 4.5005
R23348 XThR.Tn[7].n78 XThR.Tn[7].n77 4.5005
R23349 XThR.Tn[7].n83 XThR.Tn[7].n82 4.5005
R23350 XThR.Tn[7].n84 XThR.Tn[7] 3.70586
R23351 XThR.Tn[7].n13 XThR.Tn[7] 2.52282
R23352 XThR.Tn[7].n18 XThR.Tn[7] 2.52282
R23353 XThR.Tn[7].n23 XThR.Tn[7] 2.52282
R23354 XThR.Tn[7].n28 XThR.Tn[7] 2.52282
R23355 XThR.Tn[7].n33 XThR.Tn[7] 2.52282
R23356 XThR.Tn[7].n38 XThR.Tn[7] 2.52282
R23357 XThR.Tn[7].n43 XThR.Tn[7] 2.52282
R23358 XThR.Tn[7].n48 XThR.Tn[7] 2.52282
R23359 XThR.Tn[7].n53 XThR.Tn[7] 2.52282
R23360 XThR.Tn[7].n58 XThR.Tn[7] 2.52282
R23361 XThR.Tn[7].n63 XThR.Tn[7] 2.52282
R23362 XThR.Tn[7].n68 XThR.Tn[7] 2.52282
R23363 XThR.Tn[7].n73 XThR.Tn[7] 2.52282
R23364 XThR.Tn[7].n78 XThR.Tn[7] 2.52282
R23365 XThR.Tn[7].n83 XThR.Tn[7] 2.52282
R23366 XThR.Tn[7].n85 XThR.Tn[7] 2.49401
R23367 XThR.Tn[7].n81 XThR.Tn[7] 1.08677
R23368 XThR.Tn[7].n76 XThR.Tn[7] 1.08677
R23369 XThR.Tn[7].n71 XThR.Tn[7] 1.08677
R23370 XThR.Tn[7].n66 XThR.Tn[7] 1.08677
R23371 XThR.Tn[7].n61 XThR.Tn[7] 1.08677
R23372 XThR.Tn[7].n56 XThR.Tn[7] 1.08677
R23373 XThR.Tn[7].n51 XThR.Tn[7] 1.08677
R23374 XThR.Tn[7].n46 XThR.Tn[7] 1.08677
R23375 XThR.Tn[7].n41 XThR.Tn[7] 1.08677
R23376 XThR.Tn[7].n36 XThR.Tn[7] 1.08677
R23377 XThR.Tn[7].n31 XThR.Tn[7] 1.08677
R23378 XThR.Tn[7].n26 XThR.Tn[7] 1.08677
R23379 XThR.Tn[7].n21 XThR.Tn[7] 1.08677
R23380 XThR.Tn[7].n16 XThR.Tn[7] 1.08677
R23381 XThR.Tn[7].n11 XThR.Tn[7] 1.08677
R23382 XThR.Tn[7] XThR.Tn[7].n13 0.839786
R23383 XThR.Tn[7] XThR.Tn[7].n18 0.839786
R23384 XThR.Tn[7] XThR.Tn[7].n23 0.839786
R23385 XThR.Tn[7] XThR.Tn[7].n28 0.839786
R23386 XThR.Tn[7] XThR.Tn[7].n33 0.839786
R23387 XThR.Tn[7] XThR.Tn[7].n38 0.839786
R23388 XThR.Tn[7] XThR.Tn[7].n43 0.839786
R23389 XThR.Tn[7] XThR.Tn[7].n48 0.839786
R23390 XThR.Tn[7] XThR.Tn[7].n53 0.839786
R23391 XThR.Tn[7] XThR.Tn[7].n58 0.839786
R23392 XThR.Tn[7] XThR.Tn[7].n63 0.839786
R23393 XThR.Tn[7] XThR.Tn[7].n68 0.839786
R23394 XThR.Tn[7] XThR.Tn[7].n73 0.839786
R23395 XThR.Tn[7] XThR.Tn[7].n78 0.839786
R23396 XThR.Tn[7] XThR.Tn[7].n83 0.839786
R23397 XThR.Tn[7].n6 XThR.Tn[7] 0.829611
R23398 XThR.Tn[7].n8 XThR.Tn[7] 0.499542
R23399 XThR.Tn[7].n82 XThR.Tn[7] 0.063
R23400 XThR.Tn[7].n77 XThR.Tn[7] 0.063
R23401 XThR.Tn[7].n72 XThR.Tn[7] 0.063
R23402 XThR.Tn[7].n67 XThR.Tn[7] 0.063
R23403 XThR.Tn[7].n62 XThR.Tn[7] 0.063
R23404 XThR.Tn[7].n57 XThR.Tn[7] 0.063
R23405 XThR.Tn[7].n52 XThR.Tn[7] 0.063
R23406 XThR.Tn[7].n47 XThR.Tn[7] 0.063
R23407 XThR.Tn[7].n42 XThR.Tn[7] 0.063
R23408 XThR.Tn[7].n37 XThR.Tn[7] 0.063
R23409 XThR.Tn[7].n32 XThR.Tn[7] 0.063
R23410 XThR.Tn[7].n27 XThR.Tn[7] 0.063
R23411 XThR.Tn[7].n22 XThR.Tn[7] 0.063
R23412 XThR.Tn[7].n17 XThR.Tn[7] 0.063
R23413 XThR.Tn[7].n12 XThR.Tn[7] 0.063
R23414 XThR.Tn[7].n84 XThR.Tn[7] 0.0540714
R23415 XThR.Tn[7] XThR.Tn[7].n84 0.038
R23416 XThR.Tn[7].n8 XThR.Tn[7] 0.0143889
R23417 XThR.Tn[7].n82 XThR.Tn[7].n81 0.00771154
R23418 XThR.Tn[7].n77 XThR.Tn[7].n76 0.00771154
R23419 XThR.Tn[7].n72 XThR.Tn[7].n71 0.00771154
R23420 XThR.Tn[7].n67 XThR.Tn[7].n66 0.00771154
R23421 XThR.Tn[7].n62 XThR.Tn[7].n61 0.00771154
R23422 XThR.Tn[7].n57 XThR.Tn[7].n56 0.00771154
R23423 XThR.Tn[7].n52 XThR.Tn[7].n51 0.00771154
R23424 XThR.Tn[7].n47 XThR.Tn[7].n46 0.00771154
R23425 XThR.Tn[7].n42 XThR.Tn[7].n41 0.00771154
R23426 XThR.Tn[7].n37 XThR.Tn[7].n36 0.00771154
R23427 XThR.Tn[7].n32 XThR.Tn[7].n31 0.00771154
R23428 XThR.Tn[7].n27 XThR.Tn[7].n26 0.00771154
R23429 XThR.Tn[7].n22 XThR.Tn[7].n21 0.00771154
R23430 XThR.Tn[7].n17 XThR.Tn[7].n16 0.00771154
R23431 XThR.Tn[7].n12 XThR.Tn[7].n11 0.00771154
R23432 XThR.Tn[0].n2 XThR.Tn[0].n1 332.332
R23433 XThR.Tn[0].n2 XThR.Tn[0].n0 296.493
R23434 XThR.Tn[0] XThR.Tn[0].n82 161.363
R23435 XThR.Tn[0] XThR.Tn[0].n77 161.363
R23436 XThR.Tn[0] XThR.Tn[0].n72 161.363
R23437 XThR.Tn[0] XThR.Tn[0].n67 161.363
R23438 XThR.Tn[0] XThR.Tn[0].n62 161.363
R23439 XThR.Tn[0] XThR.Tn[0].n57 161.363
R23440 XThR.Tn[0] XThR.Tn[0].n52 161.363
R23441 XThR.Tn[0] XThR.Tn[0].n47 161.363
R23442 XThR.Tn[0] XThR.Tn[0].n42 161.363
R23443 XThR.Tn[0] XThR.Tn[0].n37 161.363
R23444 XThR.Tn[0] XThR.Tn[0].n32 161.363
R23445 XThR.Tn[0] XThR.Tn[0].n27 161.363
R23446 XThR.Tn[0] XThR.Tn[0].n22 161.363
R23447 XThR.Tn[0] XThR.Tn[0].n17 161.363
R23448 XThR.Tn[0] XThR.Tn[0].n12 161.363
R23449 XThR.Tn[0] XThR.Tn[0].n10 161.363
R23450 XThR.Tn[0].n84 XThR.Tn[0].n83 161.3
R23451 XThR.Tn[0].n79 XThR.Tn[0].n78 161.3
R23452 XThR.Tn[0].n74 XThR.Tn[0].n73 161.3
R23453 XThR.Tn[0].n69 XThR.Tn[0].n68 161.3
R23454 XThR.Tn[0].n64 XThR.Tn[0].n63 161.3
R23455 XThR.Tn[0].n59 XThR.Tn[0].n58 161.3
R23456 XThR.Tn[0].n54 XThR.Tn[0].n53 161.3
R23457 XThR.Tn[0].n49 XThR.Tn[0].n48 161.3
R23458 XThR.Tn[0].n44 XThR.Tn[0].n43 161.3
R23459 XThR.Tn[0].n39 XThR.Tn[0].n38 161.3
R23460 XThR.Tn[0].n34 XThR.Tn[0].n33 161.3
R23461 XThR.Tn[0].n29 XThR.Tn[0].n28 161.3
R23462 XThR.Tn[0].n24 XThR.Tn[0].n23 161.3
R23463 XThR.Tn[0].n19 XThR.Tn[0].n18 161.3
R23464 XThR.Tn[0].n14 XThR.Tn[0].n13 161.3
R23465 XThR.Tn[0].n82 XThR.Tn[0].t32 161.106
R23466 XThR.Tn[0].n77 XThR.Tn[0].t36 161.106
R23467 XThR.Tn[0].n72 XThR.Tn[0].t16 161.106
R23468 XThR.Tn[0].n67 XThR.Tn[0].t65 161.106
R23469 XThR.Tn[0].n62 XThR.Tn[0].t31 161.106
R23470 XThR.Tn[0].n57 XThR.Tn[0].t53 161.106
R23471 XThR.Tn[0].n52 XThR.Tn[0].t34 161.106
R23472 XThR.Tn[0].n47 XThR.Tn[0].t14 161.106
R23473 XThR.Tn[0].n42 XThR.Tn[0].t63 161.106
R23474 XThR.Tn[0].n37 XThR.Tn[0].t68 161.106
R23475 XThR.Tn[0].n32 XThR.Tn[0].t52 161.106
R23476 XThR.Tn[0].n27 XThR.Tn[0].t15 161.106
R23477 XThR.Tn[0].n22 XThR.Tn[0].t51 161.106
R23478 XThR.Tn[0].n17 XThR.Tn[0].t33 161.106
R23479 XThR.Tn[0].n12 XThR.Tn[0].t58 161.106
R23480 XThR.Tn[0].n10 XThR.Tn[0].t40 161.106
R23481 XThR.Tn[0].n83 XThR.Tn[0].t20 159.978
R23482 XThR.Tn[0].n78 XThR.Tn[0].t30 159.978
R23483 XThR.Tn[0].n73 XThR.Tn[0].t73 159.978
R23484 XThR.Tn[0].n68 XThR.Tn[0].t57 159.978
R23485 XThR.Tn[0].n63 XThR.Tn[0].t19 159.978
R23486 XThR.Tn[0].n58 XThR.Tn[0].t49 159.978
R23487 XThR.Tn[0].n53 XThR.Tn[0].t29 159.978
R23488 XThR.Tn[0].n48 XThR.Tn[0].t71 159.978
R23489 XThR.Tn[0].n43 XThR.Tn[0].t55 159.978
R23490 XThR.Tn[0].n38 XThR.Tn[0].t64 159.978
R23491 XThR.Tn[0].n33 XThR.Tn[0].t46 159.978
R23492 XThR.Tn[0].n28 XThR.Tn[0].t72 159.978
R23493 XThR.Tn[0].n23 XThR.Tn[0].t44 159.978
R23494 XThR.Tn[0].n18 XThR.Tn[0].t26 159.978
R23495 XThR.Tn[0].n13 XThR.Tn[0].t50 159.978
R23496 XThR.Tn[0].n82 XThR.Tn[0].t18 145.038
R23497 XThR.Tn[0].n77 XThR.Tn[0].t42 145.038
R23498 XThR.Tn[0].n72 XThR.Tn[0].t22 145.038
R23499 XThR.Tn[0].n67 XThR.Tn[0].t69 145.038
R23500 XThR.Tn[0].n62 XThR.Tn[0].t37 145.038
R23501 XThR.Tn[0].n57 XThR.Tn[0].t17 145.038
R23502 XThR.Tn[0].n52 XThR.Tn[0].t25 145.038
R23503 XThR.Tn[0].n47 XThR.Tn[0].t70 145.038
R23504 XThR.Tn[0].n42 XThR.Tn[0].t66 145.038
R23505 XThR.Tn[0].n37 XThR.Tn[0].t35 145.038
R23506 XThR.Tn[0].n32 XThR.Tn[0].t60 145.038
R23507 XThR.Tn[0].n27 XThR.Tn[0].t21 145.038
R23508 XThR.Tn[0].n22 XThR.Tn[0].t59 145.038
R23509 XThR.Tn[0].n17 XThR.Tn[0].t41 145.038
R23510 XThR.Tn[0].n12 XThR.Tn[0].t67 145.038
R23511 XThR.Tn[0].n10 XThR.Tn[0].t48 145.038
R23512 XThR.Tn[0].n83 XThR.Tn[0].t39 143.911
R23513 XThR.Tn[0].n78 XThR.Tn[0].t62 143.911
R23514 XThR.Tn[0].n73 XThR.Tn[0].t45 143.911
R23515 XThR.Tn[0].n68 XThR.Tn[0].t27 143.911
R23516 XThR.Tn[0].n63 XThR.Tn[0].t56 143.911
R23517 XThR.Tn[0].n58 XThR.Tn[0].t38 143.911
R23518 XThR.Tn[0].n53 XThR.Tn[0].t47 143.911
R23519 XThR.Tn[0].n48 XThR.Tn[0].t28 143.911
R23520 XThR.Tn[0].n43 XThR.Tn[0].t23 143.911
R23521 XThR.Tn[0].n38 XThR.Tn[0].t54 143.911
R23522 XThR.Tn[0].n33 XThR.Tn[0].t13 143.911
R23523 XThR.Tn[0].n28 XThR.Tn[0].t43 143.911
R23524 XThR.Tn[0].n23 XThR.Tn[0].t12 143.911
R23525 XThR.Tn[0].n18 XThR.Tn[0].t61 143.911
R23526 XThR.Tn[0].n13 XThR.Tn[0].t24 143.911
R23527 XThR.Tn[0].n7 XThR.Tn[0].n6 135.249
R23528 XThR.Tn[0].n9 XThR.Tn[0].n3 98.982
R23529 XThR.Tn[0].n8 XThR.Tn[0].n4 98.982
R23530 XThR.Tn[0].n7 XThR.Tn[0].n5 98.982
R23531 XThR.Tn[0].n9 XThR.Tn[0].n8 36.2672
R23532 XThR.Tn[0].n8 XThR.Tn[0].n7 36.2672
R23533 XThR.Tn[0].n88 XThR.Tn[0].n9 32.6405
R23534 XThR.Tn[0].n1 XThR.Tn[0].t2 26.5955
R23535 XThR.Tn[0].n1 XThR.Tn[0].t1 26.5955
R23536 XThR.Tn[0].n0 XThR.Tn[0].t3 26.5955
R23537 XThR.Tn[0].n0 XThR.Tn[0].t4 26.5955
R23538 XThR.Tn[0].n3 XThR.Tn[0].t6 24.9236
R23539 XThR.Tn[0].n3 XThR.Tn[0].t7 24.9236
R23540 XThR.Tn[0].n4 XThR.Tn[0].t5 24.9236
R23541 XThR.Tn[0].n4 XThR.Tn[0].t8 24.9236
R23542 XThR.Tn[0].n5 XThR.Tn[0].t11 24.9236
R23543 XThR.Tn[0].n5 XThR.Tn[0].t9 24.9236
R23544 XThR.Tn[0].n6 XThR.Tn[0].t0 24.9236
R23545 XThR.Tn[0].n6 XThR.Tn[0].t10 24.9236
R23546 XThR.Tn[0] XThR.Tn[0].n2 23.3605
R23547 XThR.Tn[0] XThR.Tn[0].n88 6.7205
R23548 XThR.Tn[0].n88 XThR.Tn[0] 6.36522
R23549 XThR.Tn[0] XThR.Tn[0].n11 5.34038
R23550 XThR.Tn[0].n16 XThR.Tn[0].n15 4.5005
R23551 XThR.Tn[0].n21 XThR.Tn[0].n20 4.5005
R23552 XThR.Tn[0].n26 XThR.Tn[0].n25 4.5005
R23553 XThR.Tn[0].n31 XThR.Tn[0].n30 4.5005
R23554 XThR.Tn[0].n36 XThR.Tn[0].n35 4.5005
R23555 XThR.Tn[0].n41 XThR.Tn[0].n40 4.5005
R23556 XThR.Tn[0].n46 XThR.Tn[0].n45 4.5005
R23557 XThR.Tn[0].n51 XThR.Tn[0].n50 4.5005
R23558 XThR.Tn[0].n56 XThR.Tn[0].n55 4.5005
R23559 XThR.Tn[0].n61 XThR.Tn[0].n60 4.5005
R23560 XThR.Tn[0].n66 XThR.Tn[0].n65 4.5005
R23561 XThR.Tn[0].n71 XThR.Tn[0].n70 4.5005
R23562 XThR.Tn[0].n76 XThR.Tn[0].n75 4.5005
R23563 XThR.Tn[0].n81 XThR.Tn[0].n80 4.5005
R23564 XThR.Tn[0].n86 XThR.Tn[0].n85 4.5005
R23565 XThR.Tn[0].n87 XThR.Tn[0] 3.70586
R23566 XThR.Tn[0].n16 XThR.Tn[0] 2.52282
R23567 XThR.Tn[0].n21 XThR.Tn[0] 2.52282
R23568 XThR.Tn[0].n26 XThR.Tn[0] 2.52282
R23569 XThR.Tn[0].n31 XThR.Tn[0] 2.52282
R23570 XThR.Tn[0].n36 XThR.Tn[0] 2.52282
R23571 XThR.Tn[0].n41 XThR.Tn[0] 2.52282
R23572 XThR.Tn[0].n46 XThR.Tn[0] 2.52282
R23573 XThR.Tn[0].n51 XThR.Tn[0] 2.52282
R23574 XThR.Tn[0].n56 XThR.Tn[0] 2.52282
R23575 XThR.Tn[0].n61 XThR.Tn[0] 2.52282
R23576 XThR.Tn[0].n66 XThR.Tn[0] 2.52282
R23577 XThR.Tn[0].n71 XThR.Tn[0] 2.52282
R23578 XThR.Tn[0].n76 XThR.Tn[0] 2.52282
R23579 XThR.Tn[0].n81 XThR.Tn[0] 2.52282
R23580 XThR.Tn[0].n86 XThR.Tn[0] 2.52282
R23581 XThR.Tn[0].n84 XThR.Tn[0] 1.08677
R23582 XThR.Tn[0].n79 XThR.Tn[0] 1.08677
R23583 XThR.Tn[0].n74 XThR.Tn[0] 1.08677
R23584 XThR.Tn[0].n69 XThR.Tn[0] 1.08677
R23585 XThR.Tn[0].n64 XThR.Tn[0] 1.08677
R23586 XThR.Tn[0].n59 XThR.Tn[0] 1.08677
R23587 XThR.Tn[0].n54 XThR.Tn[0] 1.08677
R23588 XThR.Tn[0].n49 XThR.Tn[0] 1.08677
R23589 XThR.Tn[0].n44 XThR.Tn[0] 1.08677
R23590 XThR.Tn[0].n39 XThR.Tn[0] 1.08677
R23591 XThR.Tn[0].n34 XThR.Tn[0] 1.08677
R23592 XThR.Tn[0].n29 XThR.Tn[0] 1.08677
R23593 XThR.Tn[0].n24 XThR.Tn[0] 1.08677
R23594 XThR.Tn[0].n19 XThR.Tn[0] 1.08677
R23595 XThR.Tn[0].n14 XThR.Tn[0] 1.08677
R23596 XThR.Tn[0] XThR.Tn[0].n16 0.839786
R23597 XThR.Tn[0] XThR.Tn[0].n21 0.839786
R23598 XThR.Tn[0] XThR.Tn[0].n26 0.839786
R23599 XThR.Tn[0] XThR.Tn[0].n31 0.839786
R23600 XThR.Tn[0] XThR.Tn[0].n36 0.839786
R23601 XThR.Tn[0] XThR.Tn[0].n41 0.839786
R23602 XThR.Tn[0] XThR.Tn[0].n46 0.839786
R23603 XThR.Tn[0] XThR.Tn[0].n51 0.839786
R23604 XThR.Tn[0] XThR.Tn[0].n56 0.839786
R23605 XThR.Tn[0] XThR.Tn[0].n61 0.839786
R23606 XThR.Tn[0] XThR.Tn[0].n66 0.839786
R23607 XThR.Tn[0] XThR.Tn[0].n71 0.839786
R23608 XThR.Tn[0] XThR.Tn[0].n76 0.839786
R23609 XThR.Tn[0] XThR.Tn[0].n81 0.839786
R23610 XThR.Tn[0] XThR.Tn[0].n86 0.839786
R23611 XThR.Tn[0].n11 XThR.Tn[0] 0.499542
R23612 XThR.Tn[0].n85 XThR.Tn[0] 0.063
R23613 XThR.Tn[0].n80 XThR.Tn[0] 0.063
R23614 XThR.Tn[0].n75 XThR.Tn[0] 0.063
R23615 XThR.Tn[0].n70 XThR.Tn[0] 0.063
R23616 XThR.Tn[0].n65 XThR.Tn[0] 0.063
R23617 XThR.Tn[0].n60 XThR.Tn[0] 0.063
R23618 XThR.Tn[0].n55 XThR.Tn[0] 0.063
R23619 XThR.Tn[0].n50 XThR.Tn[0] 0.063
R23620 XThR.Tn[0].n45 XThR.Tn[0] 0.063
R23621 XThR.Tn[0].n40 XThR.Tn[0] 0.063
R23622 XThR.Tn[0].n35 XThR.Tn[0] 0.063
R23623 XThR.Tn[0].n30 XThR.Tn[0] 0.063
R23624 XThR.Tn[0].n25 XThR.Tn[0] 0.063
R23625 XThR.Tn[0].n20 XThR.Tn[0] 0.063
R23626 XThR.Tn[0].n15 XThR.Tn[0] 0.063
R23627 XThR.Tn[0].n87 XThR.Tn[0] 0.0540714
R23628 XThR.Tn[0] XThR.Tn[0].n87 0.038
R23629 XThR.Tn[0].n11 XThR.Tn[0] 0.0143889
R23630 XThR.Tn[0].n85 XThR.Tn[0].n84 0.00771154
R23631 XThR.Tn[0].n80 XThR.Tn[0].n79 0.00771154
R23632 XThR.Tn[0].n75 XThR.Tn[0].n74 0.00771154
R23633 XThR.Tn[0].n70 XThR.Tn[0].n69 0.00771154
R23634 XThR.Tn[0].n65 XThR.Tn[0].n64 0.00771154
R23635 XThR.Tn[0].n60 XThR.Tn[0].n59 0.00771154
R23636 XThR.Tn[0].n55 XThR.Tn[0].n54 0.00771154
R23637 XThR.Tn[0].n50 XThR.Tn[0].n49 0.00771154
R23638 XThR.Tn[0].n45 XThR.Tn[0].n44 0.00771154
R23639 XThR.Tn[0].n40 XThR.Tn[0].n39 0.00771154
R23640 XThR.Tn[0].n35 XThR.Tn[0].n34 0.00771154
R23641 XThR.Tn[0].n30 XThR.Tn[0].n29 0.00771154
R23642 XThR.Tn[0].n25 XThR.Tn[0].n24 0.00771154
R23643 XThR.Tn[0].n20 XThR.Tn[0].n19 0.00771154
R23644 XThR.Tn[0].n15 XThR.Tn[0].n14 0.00771154
R23645 XThR.Tn[8].n87 XThR.Tn[8].n86 256.103
R23646 XThR.Tn[8].n2 XThR.Tn[8].n0 243.68
R23647 XThR.Tn[8].n5 XThR.Tn[8].n3 241.847
R23648 XThR.Tn[8].n2 XThR.Tn[8].n1 205.28
R23649 XThR.Tn[8].n87 XThR.Tn[8].n85 202.094
R23650 XThR.Tn[8].n5 XThR.Tn[8].n4 185
R23651 XThR.Tn[8] XThR.Tn[8].n78 161.363
R23652 XThR.Tn[8] XThR.Tn[8].n73 161.363
R23653 XThR.Tn[8] XThR.Tn[8].n68 161.363
R23654 XThR.Tn[8] XThR.Tn[8].n63 161.363
R23655 XThR.Tn[8] XThR.Tn[8].n58 161.363
R23656 XThR.Tn[8] XThR.Tn[8].n53 161.363
R23657 XThR.Tn[8] XThR.Tn[8].n48 161.363
R23658 XThR.Tn[8] XThR.Tn[8].n43 161.363
R23659 XThR.Tn[8] XThR.Tn[8].n38 161.363
R23660 XThR.Tn[8] XThR.Tn[8].n33 161.363
R23661 XThR.Tn[8] XThR.Tn[8].n28 161.363
R23662 XThR.Tn[8] XThR.Tn[8].n23 161.363
R23663 XThR.Tn[8] XThR.Tn[8].n18 161.363
R23664 XThR.Tn[8] XThR.Tn[8].n13 161.363
R23665 XThR.Tn[8] XThR.Tn[8].n8 161.363
R23666 XThR.Tn[8] XThR.Tn[8].n6 161.363
R23667 XThR.Tn[8].n80 XThR.Tn[8].n79 161.3
R23668 XThR.Tn[8].n75 XThR.Tn[8].n74 161.3
R23669 XThR.Tn[8].n70 XThR.Tn[8].n69 161.3
R23670 XThR.Tn[8].n65 XThR.Tn[8].n64 161.3
R23671 XThR.Tn[8].n60 XThR.Tn[8].n59 161.3
R23672 XThR.Tn[8].n55 XThR.Tn[8].n54 161.3
R23673 XThR.Tn[8].n50 XThR.Tn[8].n49 161.3
R23674 XThR.Tn[8].n45 XThR.Tn[8].n44 161.3
R23675 XThR.Tn[8].n40 XThR.Tn[8].n39 161.3
R23676 XThR.Tn[8].n35 XThR.Tn[8].n34 161.3
R23677 XThR.Tn[8].n30 XThR.Tn[8].n29 161.3
R23678 XThR.Tn[8].n25 XThR.Tn[8].n24 161.3
R23679 XThR.Tn[8].n20 XThR.Tn[8].n19 161.3
R23680 XThR.Tn[8].n15 XThR.Tn[8].n14 161.3
R23681 XThR.Tn[8].n10 XThR.Tn[8].n9 161.3
R23682 XThR.Tn[8].n78 XThR.Tn[8].t23 161.106
R23683 XThR.Tn[8].n73 XThR.Tn[8].t29 161.106
R23684 XThR.Tn[8].n68 XThR.Tn[8].t71 161.106
R23685 XThR.Tn[8].n63 XThR.Tn[8].t57 161.106
R23686 XThR.Tn[8].n58 XThR.Tn[8].t21 161.106
R23687 XThR.Tn[8].n53 XThR.Tn[8].t46 161.106
R23688 XThR.Tn[8].n48 XThR.Tn[8].t27 161.106
R23689 XThR.Tn[8].n43 XThR.Tn[8].t69 161.106
R23690 XThR.Tn[8].n38 XThR.Tn[8].t56 161.106
R23691 XThR.Tn[8].n33 XThR.Tn[8].t61 161.106
R23692 XThR.Tn[8].n28 XThR.Tn[8].t44 161.106
R23693 XThR.Tn[8].n23 XThR.Tn[8].t70 161.106
R23694 XThR.Tn[8].n18 XThR.Tn[8].t43 161.106
R23695 XThR.Tn[8].n13 XThR.Tn[8].t26 161.106
R23696 XThR.Tn[8].n8 XThR.Tn[8].t49 161.106
R23697 XThR.Tn[8].n6 XThR.Tn[8].t33 161.106
R23698 XThR.Tn[8].n79 XThR.Tn[8].t19 159.978
R23699 XThR.Tn[8].n74 XThR.Tn[8].t25 159.978
R23700 XThR.Tn[8].n69 XThR.Tn[8].t67 159.978
R23701 XThR.Tn[8].n64 XThR.Tn[8].t54 159.978
R23702 XThR.Tn[8].n59 XThR.Tn[8].t16 159.978
R23703 XThR.Tn[8].n54 XThR.Tn[8].t42 159.978
R23704 XThR.Tn[8].n49 XThR.Tn[8].t24 159.978
R23705 XThR.Tn[8].n44 XThR.Tn[8].t64 159.978
R23706 XThR.Tn[8].n39 XThR.Tn[8].t51 159.978
R23707 XThR.Tn[8].n34 XThR.Tn[8].t58 159.978
R23708 XThR.Tn[8].n29 XThR.Tn[8].t41 159.978
R23709 XThR.Tn[8].n24 XThR.Tn[8].t66 159.978
R23710 XThR.Tn[8].n19 XThR.Tn[8].t40 159.978
R23711 XThR.Tn[8].n14 XThR.Tn[8].t22 159.978
R23712 XThR.Tn[8].n9 XThR.Tn[8].t45 159.978
R23713 XThR.Tn[8].n78 XThR.Tn[8].t73 145.038
R23714 XThR.Tn[8].n73 XThR.Tn[8].t35 145.038
R23715 XThR.Tn[8].n68 XThR.Tn[8].t15 145.038
R23716 XThR.Tn[8].n63 XThR.Tn[8].t62 145.038
R23717 XThR.Tn[8].n58 XThR.Tn[8].t30 145.038
R23718 XThR.Tn[8].n53 XThR.Tn[8].t72 145.038
R23719 XThR.Tn[8].n48 XThR.Tn[8].t17 145.038
R23720 XThR.Tn[8].n43 XThR.Tn[8].t63 145.038
R23721 XThR.Tn[8].n38 XThR.Tn[8].t60 145.038
R23722 XThR.Tn[8].n33 XThR.Tn[8].t28 145.038
R23723 XThR.Tn[8].n28 XThR.Tn[8].t52 145.038
R23724 XThR.Tn[8].n23 XThR.Tn[8].t12 145.038
R23725 XThR.Tn[8].n18 XThR.Tn[8].t50 145.038
R23726 XThR.Tn[8].n13 XThR.Tn[8].t34 145.038
R23727 XThR.Tn[8].n8 XThR.Tn[8].t59 145.038
R23728 XThR.Tn[8].n6 XThR.Tn[8].t39 145.038
R23729 XThR.Tn[8].n79 XThR.Tn[8].t32 143.911
R23730 XThR.Tn[8].n74 XThR.Tn[8].t55 143.911
R23731 XThR.Tn[8].n69 XThR.Tn[8].t37 143.911
R23732 XThR.Tn[8].n64 XThR.Tn[8].t18 143.911
R23733 XThR.Tn[8].n59 XThR.Tn[8].t48 143.911
R23734 XThR.Tn[8].n54 XThR.Tn[8].t31 143.911
R23735 XThR.Tn[8].n49 XThR.Tn[8].t38 143.911
R23736 XThR.Tn[8].n44 XThR.Tn[8].t20 143.911
R23737 XThR.Tn[8].n39 XThR.Tn[8].t14 143.911
R23738 XThR.Tn[8].n34 XThR.Tn[8].t47 143.911
R23739 XThR.Tn[8].n29 XThR.Tn[8].t68 143.911
R23740 XThR.Tn[8].n24 XThR.Tn[8].t36 143.911
R23741 XThR.Tn[8].n19 XThR.Tn[8].t65 143.911
R23742 XThR.Tn[8].n14 XThR.Tn[8].t53 143.911
R23743 XThR.Tn[8].n9 XThR.Tn[8].t13 143.911
R23744 XThR.Tn[8] XThR.Tn[8].n2 35.7652
R23745 XThR.Tn[8].n86 XThR.Tn[8].t10 26.5955
R23746 XThR.Tn[8].n86 XThR.Tn[8].t1 26.5955
R23747 XThR.Tn[8].n0 XThR.Tn[8].t6 26.5955
R23748 XThR.Tn[8].n0 XThR.Tn[8].t4 26.5955
R23749 XThR.Tn[8].n1 XThR.Tn[8].t7 26.5955
R23750 XThR.Tn[8].n1 XThR.Tn[8].t5 26.5955
R23751 XThR.Tn[8].n85 XThR.Tn[8].t0 26.5955
R23752 XThR.Tn[8].n85 XThR.Tn[8].t2 26.5955
R23753 XThR.Tn[8].n4 XThR.Tn[8].t11 24.9236
R23754 XThR.Tn[8].n4 XThR.Tn[8].t9 24.9236
R23755 XThR.Tn[8].n3 XThR.Tn[8].t3 24.9236
R23756 XThR.Tn[8].n3 XThR.Tn[8].t8 24.9236
R23757 XThR.Tn[8] XThR.Tn[8].n5 18.8943
R23758 XThR.Tn[8].n88 XThR.Tn[8].n87 13.5534
R23759 XThR.Tn[8].n84 XThR.Tn[8] 7.82692
R23760 XThR.Tn[8].n84 XThR.Tn[8] 6.34069
R23761 XThR.Tn[8] XThR.Tn[8].n7 5.34038
R23762 XThR.Tn[8].n12 XThR.Tn[8].n11 4.5005
R23763 XThR.Tn[8].n17 XThR.Tn[8].n16 4.5005
R23764 XThR.Tn[8].n22 XThR.Tn[8].n21 4.5005
R23765 XThR.Tn[8].n27 XThR.Tn[8].n26 4.5005
R23766 XThR.Tn[8].n32 XThR.Tn[8].n31 4.5005
R23767 XThR.Tn[8].n37 XThR.Tn[8].n36 4.5005
R23768 XThR.Tn[8].n42 XThR.Tn[8].n41 4.5005
R23769 XThR.Tn[8].n47 XThR.Tn[8].n46 4.5005
R23770 XThR.Tn[8].n52 XThR.Tn[8].n51 4.5005
R23771 XThR.Tn[8].n57 XThR.Tn[8].n56 4.5005
R23772 XThR.Tn[8].n62 XThR.Tn[8].n61 4.5005
R23773 XThR.Tn[8].n67 XThR.Tn[8].n66 4.5005
R23774 XThR.Tn[8].n72 XThR.Tn[8].n71 4.5005
R23775 XThR.Tn[8].n77 XThR.Tn[8].n76 4.5005
R23776 XThR.Tn[8].n82 XThR.Tn[8].n81 4.5005
R23777 XThR.Tn[8].n83 XThR.Tn[8] 3.70586
R23778 XThR.Tn[8].n12 XThR.Tn[8] 2.52282
R23779 XThR.Tn[8].n17 XThR.Tn[8] 2.52282
R23780 XThR.Tn[8].n22 XThR.Tn[8] 2.52282
R23781 XThR.Tn[8].n27 XThR.Tn[8] 2.52282
R23782 XThR.Tn[8].n32 XThR.Tn[8] 2.52282
R23783 XThR.Tn[8].n37 XThR.Tn[8] 2.52282
R23784 XThR.Tn[8].n42 XThR.Tn[8] 2.52282
R23785 XThR.Tn[8].n47 XThR.Tn[8] 2.52282
R23786 XThR.Tn[8].n52 XThR.Tn[8] 2.52282
R23787 XThR.Tn[8].n57 XThR.Tn[8] 2.52282
R23788 XThR.Tn[8].n62 XThR.Tn[8] 2.52282
R23789 XThR.Tn[8].n67 XThR.Tn[8] 2.52282
R23790 XThR.Tn[8].n72 XThR.Tn[8] 2.52282
R23791 XThR.Tn[8].n77 XThR.Tn[8] 2.52282
R23792 XThR.Tn[8].n82 XThR.Tn[8] 2.52282
R23793 XThR.Tn[8] XThR.Tn[8].n84 1.79489
R23794 XThR.Tn[8] XThR.Tn[8].n88 1.50638
R23795 XThR.Tn[8].n88 XThR.Tn[8] 1.19676
R23796 XThR.Tn[8].n80 XThR.Tn[8] 1.08677
R23797 XThR.Tn[8].n75 XThR.Tn[8] 1.08677
R23798 XThR.Tn[8].n70 XThR.Tn[8] 1.08677
R23799 XThR.Tn[8].n65 XThR.Tn[8] 1.08677
R23800 XThR.Tn[8].n60 XThR.Tn[8] 1.08677
R23801 XThR.Tn[8].n55 XThR.Tn[8] 1.08677
R23802 XThR.Tn[8].n50 XThR.Tn[8] 1.08677
R23803 XThR.Tn[8].n45 XThR.Tn[8] 1.08677
R23804 XThR.Tn[8].n40 XThR.Tn[8] 1.08677
R23805 XThR.Tn[8].n35 XThR.Tn[8] 1.08677
R23806 XThR.Tn[8].n30 XThR.Tn[8] 1.08677
R23807 XThR.Tn[8].n25 XThR.Tn[8] 1.08677
R23808 XThR.Tn[8].n20 XThR.Tn[8] 1.08677
R23809 XThR.Tn[8].n15 XThR.Tn[8] 1.08677
R23810 XThR.Tn[8].n10 XThR.Tn[8] 1.08677
R23811 XThR.Tn[8] XThR.Tn[8].n12 0.839786
R23812 XThR.Tn[8] XThR.Tn[8].n17 0.839786
R23813 XThR.Tn[8] XThR.Tn[8].n22 0.839786
R23814 XThR.Tn[8] XThR.Tn[8].n27 0.839786
R23815 XThR.Tn[8] XThR.Tn[8].n32 0.839786
R23816 XThR.Tn[8] XThR.Tn[8].n37 0.839786
R23817 XThR.Tn[8] XThR.Tn[8].n42 0.839786
R23818 XThR.Tn[8] XThR.Tn[8].n47 0.839786
R23819 XThR.Tn[8] XThR.Tn[8].n52 0.839786
R23820 XThR.Tn[8] XThR.Tn[8].n57 0.839786
R23821 XThR.Tn[8] XThR.Tn[8].n62 0.839786
R23822 XThR.Tn[8] XThR.Tn[8].n67 0.839786
R23823 XThR.Tn[8] XThR.Tn[8].n72 0.839786
R23824 XThR.Tn[8] XThR.Tn[8].n77 0.839786
R23825 XThR.Tn[8] XThR.Tn[8].n82 0.839786
R23826 XThR.Tn[8].n7 XThR.Tn[8] 0.499542
R23827 XThR.Tn[8].n81 XThR.Tn[8] 0.063
R23828 XThR.Tn[8].n76 XThR.Tn[8] 0.063
R23829 XThR.Tn[8].n71 XThR.Tn[8] 0.063
R23830 XThR.Tn[8].n66 XThR.Tn[8] 0.063
R23831 XThR.Tn[8].n61 XThR.Tn[8] 0.063
R23832 XThR.Tn[8].n56 XThR.Tn[8] 0.063
R23833 XThR.Tn[8].n51 XThR.Tn[8] 0.063
R23834 XThR.Tn[8].n46 XThR.Tn[8] 0.063
R23835 XThR.Tn[8].n41 XThR.Tn[8] 0.063
R23836 XThR.Tn[8].n36 XThR.Tn[8] 0.063
R23837 XThR.Tn[8].n31 XThR.Tn[8] 0.063
R23838 XThR.Tn[8].n26 XThR.Tn[8] 0.063
R23839 XThR.Tn[8].n21 XThR.Tn[8] 0.063
R23840 XThR.Tn[8].n16 XThR.Tn[8] 0.063
R23841 XThR.Tn[8].n11 XThR.Tn[8] 0.063
R23842 XThR.Tn[8].n83 XThR.Tn[8] 0.0540714
R23843 XThR.Tn[8] XThR.Tn[8].n83 0.038
R23844 XThR.Tn[8].n7 XThR.Tn[8] 0.0143889
R23845 XThR.Tn[8].n81 XThR.Tn[8].n80 0.00771154
R23846 XThR.Tn[8].n76 XThR.Tn[8].n75 0.00771154
R23847 XThR.Tn[8].n71 XThR.Tn[8].n70 0.00771154
R23848 XThR.Tn[8].n66 XThR.Tn[8].n65 0.00771154
R23849 XThR.Tn[8].n61 XThR.Tn[8].n60 0.00771154
R23850 XThR.Tn[8].n56 XThR.Tn[8].n55 0.00771154
R23851 XThR.Tn[8].n51 XThR.Tn[8].n50 0.00771154
R23852 XThR.Tn[8].n46 XThR.Tn[8].n45 0.00771154
R23853 XThR.Tn[8].n41 XThR.Tn[8].n40 0.00771154
R23854 XThR.Tn[8].n36 XThR.Tn[8].n35 0.00771154
R23855 XThR.Tn[8].n31 XThR.Tn[8].n30 0.00771154
R23856 XThR.Tn[8].n26 XThR.Tn[8].n25 0.00771154
R23857 XThR.Tn[8].n21 XThR.Tn[8].n20 0.00771154
R23858 XThR.Tn[8].n16 XThR.Tn[8].n15 0.00771154
R23859 XThR.Tn[8].n11 XThR.Tn[8].n10 0.00771154
R23860 XThC.XTB3.Y.n6 XThC.XTB3.Y.t3 212.081
R23861 XThC.XTB3.Y.n5 XThC.XTB3.Y.t15 212.081
R23862 XThC.XTB3.Y.n11 XThC.XTB3.Y.t14 212.081
R23863 XThC.XTB3.Y.n3 XThC.XTB3.Y.t10 212.081
R23864 XThC.XTB3.Y.n15 XThC.XTB3.Y.t11 212.081
R23865 XThC.XTB3.Y.n16 XThC.XTB3.Y.t12 212.081
R23866 XThC.XTB3.Y.n18 XThC.XTB3.Y.t4 212.081
R23867 XThC.XTB3.Y.n14 XThC.XTB3.Y.t16 212.081
R23868 XThC.XTB3.Y.n22 XThC.XTB3.Y.n2 201.288
R23869 XThC.XTB3.Y.n8 XThC.XTB3.Y.n7 173.761
R23870 XThC.XTB3.Y.n17 XThC.XTB3.Y 158.656
R23871 XThC.XTB3.Y.n10 XThC.XTB3.Y.n9 152
R23872 XThC.XTB3.Y.n8 XThC.XTB3.Y.n4 152
R23873 XThC.XTB3.Y.n13 XThC.XTB3.Y.n12 152
R23874 XThC.XTB3.Y.n20 XThC.XTB3.Y.n19 152
R23875 XThC.XTB3.Y.n6 XThC.XTB3.Y.t9 139.78
R23876 XThC.XTB3.Y.n5 XThC.XTB3.Y.t6 139.78
R23877 XThC.XTB3.Y.n11 XThC.XTB3.Y.t5 139.78
R23878 XThC.XTB3.Y.n3 XThC.XTB3.Y.t17 139.78
R23879 XThC.XTB3.Y.n15 XThC.XTB3.Y.t8 139.78
R23880 XThC.XTB3.Y.n16 XThC.XTB3.Y.t18 139.78
R23881 XThC.XTB3.Y.n18 XThC.XTB3.Y.t13 139.78
R23882 XThC.XTB3.Y.n14 XThC.XTB3.Y.t7 139.78
R23883 XThC.XTB3.Y.n0 XThC.XTB3.Y.t1 132.067
R23884 XThC.XTB3.Y.n21 XThC.XTB3.Y.n13 61.4096
R23885 XThC.XTB3.Y.n16 XThC.XTB3.Y.n15 61.346
R23886 XThC.XTB3.Y.n21 XThC.XTB3.Y 54.2785
R23887 XThC.XTB3.Y.n10 XThC.XTB3.Y.n4 49.6611
R23888 XThC.XTB3.Y.n12 XThC.XTB3.Y.n11 45.2793
R23889 XThC.XTB3.Y.n7 XThC.XTB3.Y.n5 42.3581
R23890 XThC.XTB3.Y.n19 XThC.XTB3.Y.n14 30.6732
R23891 XThC.XTB3.Y.n19 XThC.XTB3.Y.n18 30.6732
R23892 XThC.XTB3.Y.n18 XThC.XTB3.Y.n17 30.6732
R23893 XThC.XTB3.Y.n17 XThC.XTB3.Y.n16 30.6732
R23894 XThC.XTB3.Y.n2 XThC.XTB3.Y.t2 26.5955
R23895 XThC.XTB3.Y.n2 XThC.XTB3.Y.t0 26.5955
R23896 XThC.XTB3.Y XThC.XTB3.Y.n22 23.489
R23897 XThC.XTB3.Y.n9 XThC.XTB3.Y.n8 21.7605
R23898 XThC.XTB3.Y.n7 XThC.XTB3.Y.n6 18.9884
R23899 XThC.XTB3.Y.n12 XThC.XTB3.Y.n3 16.0672
R23900 XThC.XTB3.Y.n20 XThC.XTB3.Y 14.8485
R23901 XThC.XTB3.Y.n13 XThC.XTB3.Y 11.5205
R23902 XThC.XTB3.Y.n22 XThC.XTB3.Y.n21 10.8207
R23903 XThC.XTB3.Y.n9 XThC.XTB3.Y 10.2405
R23904 XThC.XTB3.Y XThC.XTB3.Y.n20 8.7045
R23905 XThC.XTB3.Y.n5 XThC.XTB3.Y.n4 7.30353
R23906 XThC.XTB3.Y.n11 XThC.XTB3.Y.n10 4.38232
R23907 XThC.XTB3.Y.n1 XThC.XTB3.Y.n0 4.15748
R23908 XThC.XTB3.Y XThC.XTB3.Y.n1 3.76521
R23909 XThC.XTB3.Y.n0 XThC.XTB3.Y 1.17559
R23910 XThC.XTB3.Y.n1 XThC.XTB3.Y 0.921363
R23911 data[4].n3 data[4].t0 231.835
R23912 data[4].n0 data[4].t3 230.155
R23913 data[4].n0 data[4].t1 157.856
R23914 data[4].n3 data[4].t2 157.07
R23915 data[4].n1 data[4].n0 152
R23916 data[4].n4 data[4].n3 152
R23917 data[4].n2 data[4].n1 25.6681
R23918 data[4].n4 data[4].n2 10.7642
R23919 data[4].n2 data[4] 2.763
R23920 data[4].n1 data[4] 2.10199
R23921 data[4] data[4].n4 2.01193
R23922 XThR.Tn[13].n8 XThR.Tn[13].n7 256.104
R23923 XThR.Tn[13].n5 XThR.Tn[13].n3 243.68
R23924 XThR.Tn[13].n2 XThR.Tn[13].n1 241.847
R23925 XThR.Tn[13].n5 XThR.Tn[13].n4 205.28
R23926 XThR.Tn[13].n8 XThR.Tn[13].n6 202.094
R23927 XThR.Tn[13].n2 XThR.Tn[13].n0 185
R23928 XThR.Tn[13] XThR.Tn[13].n82 161.363
R23929 XThR.Tn[13] XThR.Tn[13].n77 161.363
R23930 XThR.Tn[13] XThR.Tn[13].n72 161.363
R23931 XThR.Tn[13] XThR.Tn[13].n67 161.363
R23932 XThR.Tn[13] XThR.Tn[13].n62 161.363
R23933 XThR.Tn[13] XThR.Tn[13].n57 161.363
R23934 XThR.Tn[13] XThR.Tn[13].n52 161.363
R23935 XThR.Tn[13] XThR.Tn[13].n47 161.363
R23936 XThR.Tn[13] XThR.Tn[13].n42 161.363
R23937 XThR.Tn[13] XThR.Tn[13].n37 161.363
R23938 XThR.Tn[13] XThR.Tn[13].n32 161.363
R23939 XThR.Tn[13] XThR.Tn[13].n27 161.363
R23940 XThR.Tn[13] XThR.Tn[13].n22 161.363
R23941 XThR.Tn[13] XThR.Tn[13].n17 161.363
R23942 XThR.Tn[13] XThR.Tn[13].n12 161.363
R23943 XThR.Tn[13] XThR.Tn[13].n10 161.363
R23944 XThR.Tn[13].n84 XThR.Tn[13].n83 161.3
R23945 XThR.Tn[13].n79 XThR.Tn[13].n78 161.3
R23946 XThR.Tn[13].n74 XThR.Tn[13].n73 161.3
R23947 XThR.Tn[13].n69 XThR.Tn[13].n68 161.3
R23948 XThR.Tn[13].n64 XThR.Tn[13].n63 161.3
R23949 XThR.Tn[13].n59 XThR.Tn[13].n58 161.3
R23950 XThR.Tn[13].n54 XThR.Tn[13].n53 161.3
R23951 XThR.Tn[13].n49 XThR.Tn[13].n48 161.3
R23952 XThR.Tn[13].n44 XThR.Tn[13].n43 161.3
R23953 XThR.Tn[13].n39 XThR.Tn[13].n38 161.3
R23954 XThR.Tn[13].n34 XThR.Tn[13].n33 161.3
R23955 XThR.Tn[13].n29 XThR.Tn[13].n28 161.3
R23956 XThR.Tn[13].n24 XThR.Tn[13].n23 161.3
R23957 XThR.Tn[13].n19 XThR.Tn[13].n18 161.3
R23958 XThR.Tn[13].n14 XThR.Tn[13].n13 161.3
R23959 XThR.Tn[13].n82 XThR.Tn[13].t56 161.106
R23960 XThR.Tn[13].n77 XThR.Tn[13].t62 161.106
R23961 XThR.Tn[13].n72 XThR.Tn[13].t40 161.106
R23962 XThR.Tn[13].n67 XThR.Tn[13].t27 161.106
R23963 XThR.Tn[13].n62 XThR.Tn[13].t55 161.106
R23964 XThR.Tn[13].n57 XThR.Tn[13].t17 161.106
R23965 XThR.Tn[13].n52 XThR.Tn[13].t59 161.106
R23966 XThR.Tn[13].n47 XThR.Tn[13].t38 161.106
R23967 XThR.Tn[13].n42 XThR.Tn[13].t25 161.106
R23968 XThR.Tn[13].n37 XThR.Tn[13].t30 161.106
R23969 XThR.Tn[13].n32 XThR.Tn[13].t16 161.106
R23970 XThR.Tn[13].n27 XThR.Tn[13].t39 161.106
R23971 XThR.Tn[13].n22 XThR.Tn[13].t14 161.106
R23972 XThR.Tn[13].n17 XThR.Tn[13].t57 161.106
R23973 XThR.Tn[13].n12 XThR.Tn[13].t21 161.106
R23974 XThR.Tn[13].n10 XThR.Tn[13].t64 161.106
R23975 XThR.Tn[13].n83 XThR.Tn[13].t47 159.978
R23976 XThR.Tn[13].n78 XThR.Tn[13].t54 159.978
R23977 XThR.Tn[13].n73 XThR.Tn[13].t36 159.978
R23978 XThR.Tn[13].n68 XThR.Tn[13].t20 159.978
R23979 XThR.Tn[13].n63 XThR.Tn[13].t45 159.978
R23980 XThR.Tn[13].n58 XThR.Tn[13].t73 159.978
R23981 XThR.Tn[13].n53 XThR.Tn[13].t53 159.978
R23982 XThR.Tn[13].n48 XThR.Tn[13].t33 159.978
R23983 XThR.Tn[13].n43 XThR.Tn[13].t18 159.978
R23984 XThR.Tn[13].n38 XThR.Tn[13].t26 159.978
R23985 XThR.Tn[13].n33 XThR.Tn[13].t71 159.978
R23986 XThR.Tn[13].n28 XThR.Tn[13].t35 159.978
R23987 XThR.Tn[13].n23 XThR.Tn[13].t70 159.978
R23988 XThR.Tn[13].n18 XThR.Tn[13].t52 159.978
R23989 XThR.Tn[13].n13 XThR.Tn[13].t12 159.978
R23990 XThR.Tn[13].n82 XThR.Tn[13].t42 145.038
R23991 XThR.Tn[13].n77 XThR.Tn[13].t69 145.038
R23992 XThR.Tn[13].n72 XThR.Tn[13].t50 145.038
R23993 XThR.Tn[13].n67 XThR.Tn[13].t31 145.038
R23994 XThR.Tn[13].n62 XThR.Tn[13].t63 145.038
R23995 XThR.Tn[13].n57 XThR.Tn[13].t41 145.038
R23996 XThR.Tn[13].n52 XThR.Tn[13].t51 145.038
R23997 XThR.Tn[13].n47 XThR.Tn[13].t32 145.038
R23998 XThR.Tn[13].n42 XThR.Tn[13].t29 145.038
R23999 XThR.Tn[13].n37 XThR.Tn[13].t60 145.038
R24000 XThR.Tn[13].n32 XThR.Tn[13].t24 145.038
R24001 XThR.Tn[13].n27 XThR.Tn[13].t49 145.038
R24002 XThR.Tn[13].n22 XThR.Tn[13].t22 145.038
R24003 XThR.Tn[13].n17 XThR.Tn[13].t65 145.038
R24004 XThR.Tn[13].n12 XThR.Tn[13].t28 145.038
R24005 XThR.Tn[13].n10 XThR.Tn[13].t72 145.038
R24006 XThR.Tn[13].n83 XThR.Tn[13].t61 143.911
R24007 XThR.Tn[13].n78 XThR.Tn[13].t23 143.911
R24008 XThR.Tn[13].n73 XThR.Tn[13].t67 143.911
R24009 XThR.Tn[13].n68 XThR.Tn[13].t46 143.911
R24010 XThR.Tn[13].n63 XThR.Tn[13].t15 143.911
R24011 XThR.Tn[13].n58 XThR.Tn[13].t58 143.911
R24012 XThR.Tn[13].n53 XThR.Tn[13].t68 143.911
R24013 XThR.Tn[13].n48 XThR.Tn[13].t48 143.911
R24014 XThR.Tn[13].n43 XThR.Tn[13].t43 143.911
R24015 XThR.Tn[13].n38 XThR.Tn[13].t13 143.911
R24016 XThR.Tn[13].n33 XThR.Tn[13].t37 143.911
R24017 XThR.Tn[13].n28 XThR.Tn[13].t66 143.911
R24018 XThR.Tn[13].n23 XThR.Tn[13].t34 143.911
R24019 XThR.Tn[13].n18 XThR.Tn[13].t19 143.911
R24020 XThR.Tn[13].n13 XThR.Tn[13].t44 143.911
R24021 XThR.Tn[13] XThR.Tn[13].n5 35.7652
R24022 XThR.Tn[13].n6 XThR.Tn[13].t6 26.5955
R24023 XThR.Tn[13].n6 XThR.Tn[13].t4 26.5955
R24024 XThR.Tn[13].n7 XThR.Tn[13].t7 26.5955
R24025 XThR.Tn[13].n7 XThR.Tn[13].t5 26.5955
R24026 XThR.Tn[13].n3 XThR.Tn[13].t9 26.5955
R24027 XThR.Tn[13].n3 XThR.Tn[13].t11 26.5955
R24028 XThR.Tn[13].n4 XThR.Tn[13].t10 26.5955
R24029 XThR.Tn[13].n4 XThR.Tn[13].t8 26.5955
R24030 XThR.Tn[13].n0 XThR.Tn[13].t2 24.9236
R24031 XThR.Tn[13].n0 XThR.Tn[13].t0 24.9236
R24032 XThR.Tn[13].n1 XThR.Tn[13].t3 24.9236
R24033 XThR.Tn[13].n1 XThR.Tn[13].t1 24.9236
R24034 XThR.Tn[13] XThR.Tn[13].n2 22.9615
R24035 XThR.Tn[13].n9 XThR.Tn[13].n8 13.5534
R24036 XThR.Tn[13].n88 XThR.Tn[13] 8.8494
R24037 XThR.Tn[13] XThR.Tn[13].n11 5.34038
R24038 XThR.Tn[13].n16 XThR.Tn[13].n15 4.5005
R24039 XThR.Tn[13].n21 XThR.Tn[13].n20 4.5005
R24040 XThR.Tn[13].n26 XThR.Tn[13].n25 4.5005
R24041 XThR.Tn[13].n31 XThR.Tn[13].n30 4.5005
R24042 XThR.Tn[13].n36 XThR.Tn[13].n35 4.5005
R24043 XThR.Tn[13].n41 XThR.Tn[13].n40 4.5005
R24044 XThR.Tn[13].n46 XThR.Tn[13].n45 4.5005
R24045 XThR.Tn[13].n51 XThR.Tn[13].n50 4.5005
R24046 XThR.Tn[13].n56 XThR.Tn[13].n55 4.5005
R24047 XThR.Tn[13].n61 XThR.Tn[13].n60 4.5005
R24048 XThR.Tn[13].n66 XThR.Tn[13].n65 4.5005
R24049 XThR.Tn[13].n71 XThR.Tn[13].n70 4.5005
R24050 XThR.Tn[13].n76 XThR.Tn[13].n75 4.5005
R24051 XThR.Tn[13].n81 XThR.Tn[13].n80 4.5005
R24052 XThR.Tn[13].n86 XThR.Tn[13].n85 4.5005
R24053 XThR.Tn[13].n87 XThR.Tn[13] 3.70586
R24054 XThR.Tn[13].n88 XThR.Tn[13].n9 2.99115
R24055 XThR.Tn[13].n9 XThR.Tn[13] 2.87153
R24056 XThR.Tn[13].n16 XThR.Tn[13] 2.52282
R24057 XThR.Tn[13].n21 XThR.Tn[13] 2.52282
R24058 XThR.Tn[13].n26 XThR.Tn[13] 2.52282
R24059 XThR.Tn[13].n31 XThR.Tn[13] 2.52282
R24060 XThR.Tn[13].n36 XThR.Tn[13] 2.52282
R24061 XThR.Tn[13].n41 XThR.Tn[13] 2.52282
R24062 XThR.Tn[13].n46 XThR.Tn[13] 2.52282
R24063 XThR.Tn[13].n51 XThR.Tn[13] 2.52282
R24064 XThR.Tn[13].n56 XThR.Tn[13] 2.52282
R24065 XThR.Tn[13].n61 XThR.Tn[13] 2.52282
R24066 XThR.Tn[13].n66 XThR.Tn[13] 2.52282
R24067 XThR.Tn[13].n71 XThR.Tn[13] 2.52282
R24068 XThR.Tn[13].n76 XThR.Tn[13] 2.52282
R24069 XThR.Tn[13].n81 XThR.Tn[13] 2.52282
R24070 XThR.Tn[13].n86 XThR.Tn[13] 2.52282
R24071 XThR.Tn[13] XThR.Tn[13].n88 2.2734
R24072 XThR.Tn[13].n9 XThR.Tn[13] 1.50638
R24073 XThR.Tn[13].n84 XThR.Tn[13] 1.08677
R24074 XThR.Tn[13].n79 XThR.Tn[13] 1.08677
R24075 XThR.Tn[13].n74 XThR.Tn[13] 1.08677
R24076 XThR.Tn[13].n69 XThR.Tn[13] 1.08677
R24077 XThR.Tn[13].n64 XThR.Tn[13] 1.08677
R24078 XThR.Tn[13].n59 XThR.Tn[13] 1.08677
R24079 XThR.Tn[13].n54 XThR.Tn[13] 1.08677
R24080 XThR.Tn[13].n49 XThR.Tn[13] 1.08677
R24081 XThR.Tn[13].n44 XThR.Tn[13] 1.08677
R24082 XThR.Tn[13].n39 XThR.Tn[13] 1.08677
R24083 XThR.Tn[13].n34 XThR.Tn[13] 1.08677
R24084 XThR.Tn[13].n29 XThR.Tn[13] 1.08677
R24085 XThR.Tn[13].n24 XThR.Tn[13] 1.08677
R24086 XThR.Tn[13].n19 XThR.Tn[13] 1.08677
R24087 XThR.Tn[13].n14 XThR.Tn[13] 1.08677
R24088 XThR.Tn[13] XThR.Tn[13].n16 0.839786
R24089 XThR.Tn[13] XThR.Tn[13].n21 0.839786
R24090 XThR.Tn[13] XThR.Tn[13].n26 0.839786
R24091 XThR.Tn[13] XThR.Tn[13].n31 0.839786
R24092 XThR.Tn[13] XThR.Tn[13].n36 0.839786
R24093 XThR.Tn[13] XThR.Tn[13].n41 0.839786
R24094 XThR.Tn[13] XThR.Tn[13].n46 0.839786
R24095 XThR.Tn[13] XThR.Tn[13].n51 0.839786
R24096 XThR.Tn[13] XThR.Tn[13].n56 0.839786
R24097 XThR.Tn[13] XThR.Tn[13].n61 0.839786
R24098 XThR.Tn[13] XThR.Tn[13].n66 0.839786
R24099 XThR.Tn[13] XThR.Tn[13].n71 0.839786
R24100 XThR.Tn[13] XThR.Tn[13].n76 0.839786
R24101 XThR.Tn[13] XThR.Tn[13].n81 0.839786
R24102 XThR.Tn[13] XThR.Tn[13].n86 0.839786
R24103 XThR.Tn[13].n11 XThR.Tn[13] 0.499542
R24104 XThR.Tn[13].n85 XThR.Tn[13] 0.063
R24105 XThR.Tn[13].n80 XThR.Tn[13] 0.063
R24106 XThR.Tn[13].n75 XThR.Tn[13] 0.063
R24107 XThR.Tn[13].n70 XThR.Tn[13] 0.063
R24108 XThR.Tn[13].n65 XThR.Tn[13] 0.063
R24109 XThR.Tn[13].n60 XThR.Tn[13] 0.063
R24110 XThR.Tn[13].n55 XThR.Tn[13] 0.063
R24111 XThR.Tn[13].n50 XThR.Tn[13] 0.063
R24112 XThR.Tn[13].n45 XThR.Tn[13] 0.063
R24113 XThR.Tn[13].n40 XThR.Tn[13] 0.063
R24114 XThR.Tn[13].n35 XThR.Tn[13] 0.063
R24115 XThR.Tn[13].n30 XThR.Tn[13] 0.063
R24116 XThR.Tn[13].n25 XThR.Tn[13] 0.063
R24117 XThR.Tn[13].n20 XThR.Tn[13] 0.063
R24118 XThR.Tn[13].n15 XThR.Tn[13] 0.063
R24119 XThR.Tn[13].n87 XThR.Tn[13] 0.0540714
R24120 XThR.Tn[13] XThR.Tn[13].n87 0.038
R24121 XThR.Tn[13].n11 XThR.Tn[13] 0.0143889
R24122 XThR.Tn[13].n85 XThR.Tn[13].n84 0.00771154
R24123 XThR.Tn[13].n80 XThR.Tn[13].n79 0.00771154
R24124 XThR.Tn[13].n75 XThR.Tn[13].n74 0.00771154
R24125 XThR.Tn[13].n70 XThR.Tn[13].n69 0.00771154
R24126 XThR.Tn[13].n65 XThR.Tn[13].n64 0.00771154
R24127 XThR.Tn[13].n60 XThR.Tn[13].n59 0.00771154
R24128 XThR.Tn[13].n55 XThR.Tn[13].n54 0.00771154
R24129 XThR.Tn[13].n50 XThR.Tn[13].n49 0.00771154
R24130 XThR.Tn[13].n45 XThR.Tn[13].n44 0.00771154
R24131 XThR.Tn[13].n40 XThR.Tn[13].n39 0.00771154
R24132 XThR.Tn[13].n35 XThR.Tn[13].n34 0.00771154
R24133 XThR.Tn[13].n30 XThR.Tn[13].n29 0.00771154
R24134 XThR.Tn[13].n25 XThR.Tn[13].n24 0.00771154
R24135 XThR.Tn[13].n20 XThR.Tn[13].n19 0.00771154
R24136 XThR.Tn[13].n15 XThR.Tn[13].n14 0.00771154
R24137 data[0].n1 data[0].t0 230.155
R24138 data[0].n0 data[0].t2 228.463
R24139 data[0].n1 data[0].t1 157.856
R24140 data[0].n0 data[0].t3 157.07
R24141 data[0].n2 data[0].n1 152.768
R24142 data[0].n4 data[0].n0 152.256
R24143 data[0].n3 data[0].n2 24.1398
R24144 data[0].n4 data[0].n3 9.48418
R24145 data[0] data[0].n4 6.1445
R24146 data[0].n2 data[0] 5.6325
R24147 data[0].n3 data[0] 2.638
R24148 XThR.XTB1.Y.n9 XThR.XTB1.Y.t12 212.081
R24149 XThR.XTB1.Y.n10 XThR.XTB1.Y.t17 212.081
R24150 XThR.XTB1.Y.n15 XThR.XTB1.Y.t6 212.081
R24151 XThR.XTB1.Y.n16 XThR.XTB1.Y.t3 212.081
R24152 XThR.XTB1.Y.n1 XThR.XTB1.Y.t10 212.081
R24153 XThR.XTB1.Y.n2 XThR.XTB1.Y.t14 212.081
R24154 XThR.XTB1.Y.n4 XThR.XTB1.Y.t8 212.081
R24155 XThR.XTB1.Y.n5 XThR.XTB1.Y.t13 212.081
R24156 XThR.XTB1.Y.n21 XThR.XTB1.Y.n20 201.288
R24157 XThR.XTB1.Y.n12 XThR.XTB1.Y.n11 173.761
R24158 XThR.XTB1.Y.n3 XThR.XTB1.Y 167.361
R24159 XThR.XTB1.Y.n18 XThR.XTB1.Y.n17 152
R24160 XThR.XTB1.Y.n14 XThR.XTB1.Y.n13 152
R24161 XThR.XTB1.Y.n12 XThR.XTB1.Y.n8 152
R24162 XThR.XTB1.Y.n7 XThR.XTB1.Y.n6 152
R24163 XThR.XTB1.Y.n9 XThR.XTB1.Y.t16 139.78
R24164 XThR.XTB1.Y.n10 XThR.XTB1.Y.t5 139.78
R24165 XThR.XTB1.Y.n15 XThR.XTB1.Y.t11 139.78
R24166 XThR.XTB1.Y.n16 XThR.XTB1.Y.t9 139.78
R24167 XThR.XTB1.Y.n1 XThR.XTB1.Y.t18 139.78
R24168 XThR.XTB1.Y.n2 XThR.XTB1.Y.t7 139.78
R24169 XThR.XTB1.Y.n4 XThR.XTB1.Y.t15 139.78
R24170 XThR.XTB1.Y.n5 XThR.XTB1.Y.t4 139.78
R24171 XThR.XTB1.Y.n0 XThR.XTB1.Y.t1 130.548
R24172 XThR.XTB1.Y.n19 XThR.XTB1.Y 74.7655
R24173 XThR.XTB1.Y.n19 XThR.XTB1.Y.n18 61.4072
R24174 XThR.XTB1.Y.n2 XThR.XTB1.Y.n1 61.346
R24175 XThR.XTB1.Y.n14 XThR.XTB1.Y.n8 49.6611
R24176 XThR.XTB1.Y.n17 XThR.XTB1.Y.n15 45.2793
R24177 XThR.XTB1.Y.n11 XThR.XTB1.Y.n10 42.3581
R24178 XThR.XTB1.Y XThR.XTB1.Y.n21 36.289
R24179 XThR.XTB1.Y.n3 XThR.XTB1.Y.n2 30.6732
R24180 XThR.XTB1.Y.n4 XThR.XTB1.Y.n3 30.6732
R24181 XThR.XTB1.Y.n6 XThR.XTB1.Y.n4 30.6732
R24182 XThR.XTB1.Y.n6 XThR.XTB1.Y.n5 30.6732
R24183 XThR.XTB1.Y.n20 XThR.XTB1.Y.t0 26.5955
R24184 XThR.XTB1.Y.n20 XThR.XTB1.Y.t2 26.5955
R24185 XThR.XTB1.Y.n13 XThR.XTB1.Y.n12 21.7605
R24186 XThR.XTB1.Y.n13 XThR.XTB1.Y 21.1205
R24187 XThR.XTB1.Y.n11 XThR.XTB1.Y.n9 18.9884
R24188 XThR.XTB1.Y XThR.XTB1.Y.n7 17.4085
R24189 XThR.XTB1.Y.n22 XThR.XTB1.Y 16.5652
R24190 XThR.XTB1.Y.n17 XThR.XTB1.Y.n16 16.0672
R24191 XThR.XTB1.Y.n21 XThR.XTB1.Y.n19 10.8571
R24192 XThR.XTB1.Y XThR.XTB1.Y.n22 9.03579
R24193 XThR.XTB1.Y.n10 XThR.XTB1.Y.n8 7.30353
R24194 XThR.XTB1.Y.n7 XThR.XTB1.Y 6.1445
R24195 XThR.XTB1.Y.n15 XThR.XTB1.Y.n14 4.38232
R24196 XThR.XTB1.Y XThR.XTB1.Y.n0 3.46739
R24197 XThR.XTB1.Y.n0 XThR.XTB1.Y 2.74112
R24198 XThR.XTB1.Y.n22 XThR.XTB1.Y 2.21057
R24199 XThR.XTB1.Y.n18 XThR.XTB1.Y 0.6405
R24200 XThR.XTB3.Y.n9 XThR.XTB3.Y.t7 212.081
R24201 XThR.XTB3.Y.n10 XThR.XTB3.Y.t11 212.081
R24202 XThR.XTB3.Y.n15 XThR.XTB3.Y.t18 212.081
R24203 XThR.XTB3.Y.n16 XThR.XTB3.Y.t14 212.081
R24204 XThR.XTB3.Y.n1 XThR.XTB3.Y.t9 212.081
R24205 XThR.XTB3.Y.n2 XThR.XTB3.Y.t13 212.081
R24206 XThR.XTB3.Y.n4 XThR.XTB3.Y.t8 212.081
R24207 XThR.XTB3.Y.n5 XThR.XTB3.Y.t12 212.081
R24208 XThR.XTB3.Y.n21 XThR.XTB3.Y.n20 201.288
R24209 XThR.XTB3.Y.n12 XThR.XTB3.Y.n11 173.761
R24210 XThR.XTB3.Y.n3 XThR.XTB3.Y 167.361
R24211 XThR.XTB3.Y.n18 XThR.XTB3.Y.n17 152
R24212 XThR.XTB3.Y.n14 XThR.XTB3.Y.n13 152
R24213 XThR.XTB3.Y.n12 XThR.XTB3.Y.n8 152
R24214 XThR.XTB3.Y.n7 XThR.XTB3.Y.n6 152
R24215 XThR.XTB3.Y.n9 XThR.XTB3.Y.t10 139.78
R24216 XThR.XTB3.Y.n10 XThR.XTB3.Y.t16 139.78
R24217 XThR.XTB3.Y.n15 XThR.XTB3.Y.t5 139.78
R24218 XThR.XTB3.Y.n16 XThR.XTB3.Y.t3 139.78
R24219 XThR.XTB3.Y.n1 XThR.XTB3.Y.t17 139.78
R24220 XThR.XTB3.Y.n2 XThR.XTB3.Y.t6 139.78
R24221 XThR.XTB3.Y.n4 XThR.XTB3.Y.t15 139.78
R24222 XThR.XTB3.Y.n5 XThR.XTB3.Y.t4 139.78
R24223 XThR.XTB3.Y.n0 XThR.XTB3.Y.t1 130.548
R24224 XThR.XTB3.Y.n19 XThR.XTB3.Y.n18 61.4096
R24225 XThR.XTB3.Y.n2 XThR.XTB3.Y.n1 61.346
R24226 XThR.XTB3.Y.n14 XThR.XTB3.Y.n8 49.6611
R24227 XThR.XTB3.Y.n19 XThR.XTB3.Y 45.5863
R24228 XThR.XTB3.Y.n17 XThR.XTB3.Y.n15 45.2793
R24229 XThR.XTB3.Y.n11 XThR.XTB3.Y.n10 42.3581
R24230 XThR.XTB3.Y XThR.XTB3.Y.n21 36.289
R24231 XThR.XTB3.Y.n3 XThR.XTB3.Y.n2 30.6732
R24232 XThR.XTB3.Y.n4 XThR.XTB3.Y.n3 30.6732
R24233 XThR.XTB3.Y.n6 XThR.XTB3.Y.n4 30.6732
R24234 XThR.XTB3.Y.n6 XThR.XTB3.Y.n5 30.6732
R24235 XThR.XTB3.Y.n20 XThR.XTB3.Y.t0 26.5955
R24236 XThR.XTB3.Y.n20 XThR.XTB3.Y.t2 26.5955
R24237 XThR.XTB3.Y.n13 XThR.XTB3.Y.n12 21.7605
R24238 XThR.XTB3.Y.n13 XThR.XTB3.Y 21.1205
R24239 XThR.XTB3.Y.n11 XThR.XTB3.Y.n9 18.9884
R24240 XThR.XTB3.Y XThR.XTB3.Y.n7 17.4085
R24241 XThR.XTB3.Y.n22 XThR.XTB3.Y 16.5652
R24242 XThR.XTB3.Y.n17 XThR.XTB3.Y.n16 16.0672
R24243 XThR.XTB3.Y.n21 XThR.XTB3.Y.n19 10.8207
R24244 XThR.XTB3.Y XThR.XTB3.Y.n22 9.03579
R24245 XThR.XTB3.Y.n10 XThR.XTB3.Y.n8 7.30353
R24246 XThR.XTB3.Y.n7 XThR.XTB3.Y 6.1445
R24247 XThR.XTB3.Y.n15 XThR.XTB3.Y.n14 4.38232
R24248 XThR.XTB3.Y XThR.XTB3.Y.n0 3.46739
R24249 XThR.XTB3.Y.n0 XThR.XTB3.Y 2.74112
R24250 XThR.XTB3.Y.n22 XThR.XTB3.Y 2.21057
R24251 XThR.XTB3.Y.n18 XThR.XTB3.Y 0.6405
R24252 data[6].n0 data[6].t0 230.576
R24253 data[6].n0 data[6].t1 158.275
R24254 data[6].n1 data[6].n0 152
R24255 data[6].n1 data[6] 11.9995
R24256 data[6] data[6].n1 6.66717
R24257 data[1].n4 data[1].t2 230.576
R24258 data[1].n1 data[1].t0 230.363
R24259 data[1].n0 data[1].t4 229.369
R24260 data[1].n4 data[1].t5 158.275
R24261 data[1].n1 data[1].t3 158.064
R24262 data[1].n0 data[1].t1 157.07
R24263 data[1].n2 data[1].n1 153.28
R24264 data[1].n7 data[1].n0 153.147
R24265 data[1].n5 data[1].n4 152
R24266 data[1].n7 data[1].n6 16.3874
R24267 data[1].n6 data[1].n5 14.9641
R24268 data[1].n3 data[1].n2 9.3005
R24269 data[1].n6 data[1].n3 6.49639
R24270 data[1] data[1].n7 3.24826
R24271 data[1].n2 data[1] 2.92621
R24272 data[1].n3 data[1] 2.15819
R24273 data[1].n5 data[1] 2.13383
R24274 data[2].n0 data[2].t0 230.576
R24275 data[2].n0 data[2].t1 158.275
R24276 data[2].n1 data[2].n0 152
R24277 data[2].n1 data[2] 12.7714
R24278 data[2] data[2].n1 2.13383
R24279 data[5].n4 data[5].t2 230.576
R24280 data[5].n1 data[5].t0 230.363
R24281 data[5].n0 data[5].t1 229.369
R24282 data[5].n4 data[5].t5 158.275
R24283 data[5].n1 data[5].t3 158.064
R24284 data[5].n0 data[5].t4 157.07
R24285 data[5].n2 data[5].n1 152.256
R24286 data[5].n7 data[5].n0 152.238
R24287 data[5].n5 data[5].n4 152
R24288 data[5].n7 data[5].n6 16.3874
R24289 data[5].n6 data[5].n5 14.6005
R24290 data[5].n3 data[5].n2 9.3005
R24291 data[5].n5 data[5] 6.66717
R24292 data[5].n6 data[5].n3 6.49639
R24293 data[5].n2 data[5] 6.1445
R24294 data[5] data[5].n7 5.68939
R24295 data[5].n3 data[5] 2.28319
R24296 bias[1].n0 bias[1].t1 81.1889
R24297 bias[1].n2 bias[1].t0 81.1889
R24298 bias[1].n1 bias[1] 9.32819
R24299 bias[1].n1 bias[1].n0 1.06523
R24300 bias[1].n2 bias[1].n1 0.895589
R24301 bias[1] bias[1].n2 0.301839
R24302 bias[1].n0 bias[1] 0.221482
R24303 data[3].n0 data[3].t1 230.576
R24304 data[3].n0 data[3].t0 158.275
R24305 data[3].n1 data[3].n0 153.553
R24306 data[3].n1 data[3] 11.6078
R24307 data[3] data[3].n1 2.90959
R24308 data[7].n0 data[7].t0 230.576
R24309 data[7].n0 data[7].t1 158.275
R24310 data[7].n1 data[7].n0 152
R24311 data[7].n1 data[7] 11.9995
R24312 data[7] data[7].n1 6.66717
R24313 bias[2].n0 bias[2].t1 136.779
R24314 bias[2].n2 bias[2].t0 136.779
R24315 bias[2].n1 bias[2] 7.84903
R24316 bias[2].n1 bias[2].n0 1.2438
R24317 bias[2].n2 bias[2].n1 0.717018
R24318 bias[2] bias[2].n2 0.301839
R24319 bias[2].n0 bias[2] 0.221482
R24320 bias[0].n0 bias[0].t0 57.5124
R24321 bias[0].n2 bias[0].t1 57.5124
R24322 bias[0].n1 bias[0] 11.1563
R24323 bias[0].n2 bias[0].n1 1.10095
R24324 bias[0].n1 bias[0].n0 0.859875
R24325 bias[0] bias[0].n2 0.301839
R24326 bias[0].n0 bias[0] 0.221482
C0 XA.XIR[2].XIC[14].icell.Ien XA.XIR[3].XIC[14].icell.PDM 0.02104f
C1 XThR.XTBN.Y a_n1049_6699# 0.07601f
C2 XThR.Tn[5] XA.XIR[6].XIC[9].icell.PDM 0.04035f
C3 XA.XIR[7].XIC_15.icell.Ien XA.XIR[8].XIC_15.icell.PDM 0.02104f
C4 XThC.Tn[7] XThR.Tn[7] 0.40738f
C5 XA.XIR[11].XIC[2].icell.PDM Vbias 0.03928f
C6 XThC.Tn[13] Iout 0.22423f
C7 XThR.Tn[2] XA.XIR[3].XIC[1].icell.PDM 0.04035f
C8 XThC.XTB5.Y XThC.Tn[9] 0.01732f
C9 XA.XIR[10].XIC[6].icell.PDM Vbias 0.03928f
C10 XA.XIR[5].XIC[8].icell.Ien Iout 0.06801f
C11 XThC.XTB6.Y XThC.Tn[13] 0.32317f
C12 XThR.Tn[6] XA.XIR[7].XIC[8].icell.PDM 0.04035f
C13 XA.XIR[10].XIC_dummy_left.icell.Iout Iout 0.03553f
C14 XThR.XTB7.A data[4] 0.8689f
C15 XThC.Tn[4] XA.XIR[14].XIC[4].icell.Ien 0.04604f
C16 XThC.Tn[11] XThR.Tn[1] 0.40744f
C17 XA.XIR[11].XIC[5].icell.Ien XA.XIR[12].XIC[5].icell.PDM 0.02104f
C18 XA.XIR[15].XIC[6].icell.Ien Vbias 0.15966f
C19 XThR.Tn[8] XA.XIR[8].XIC[14].icell.Ien 0.144f
C20 XThR.XTB4.Y a_n1049_6699# 0.23756f
C21 XA.XIR[6].XIC_15.icell.PDM XA.XIR[6].XIC_15.icell.Ien 0.04854f
C22 XA.XIR[10].XIC_dummy_left.icell.Iout XA.XIR[11].XIC_dummy_left.icell.Iout 0.03665f
C23 XThR.XTB6.A XThR.XTB3.Y 0.03869f
C24 XThR.XTB2.Y XThR.XTB7.A 0.2319f
C25 XA.XIR[11].XIC[3].icell.PDM VPWR 0.01171f
C26 XThC.Tn[11] XThR.Tn[12] 0.40738f
C27 XA.XIR[4].XIC[9].icell.Ien Vbias 0.19161f
C28 XA.XIR[12].XIC[3].icell.Ien Iout 0.06801f
C29 XThC.Tn[1] XA.XIR[3].XIC[1].icell.Ien 0.04604f
C30 XA.XIR[0].XIC[0].icell.Ien Vbias 0.19201f
C31 XA.XIR[10].XIC[7].icell.PDM VPWR 0.01171f
C32 XA.XIR[10].XIC[13].icell.PDM XA.XIR[10].XIC[13].icell.Ien 0.04854f
C33 XA.XIR[14].XIC[14].icell.Ien Iout 0.06801f
C34 XA.XIR[10].XIC[8].icell.Ien XA.XIR[11].XIC[8].icell.PDM 0.02104f
C35 XThR.XTB7.B XThR.Tn[8] 0.05091f
C36 XA.XIR[8].XIC[3].icell.Ien Vbias 0.19161f
C37 XThC.XTBN.Y XThC.Tn[9] 0.39932f
C38 XThC.Tn[6] XThR.Tn[3] 0.40738f
C39 XThC.Tn[12] XA.XIR[15].XIC[12].icell.PDM 0.02601f
C40 XA.XIR[10].XIC[9].icell.PDM XA.XIR[10].XIC[9].icell.Ien 0.04854f
C41 XThR.Tn[5] XA.XIR[5].XIC[13].icell.Ien 0.14211f
C42 XA.XIR[0].XIC_dummy_left.icell.PDM VPWR 0.08179f
C43 XA.XIR[0].XIC[14].icell.PDM Vbias 0.03945f
C44 XA.XIR[5].XIC[7].icell.Ien VPWR 0.18829f
C45 XThR.XTB7.A a_n1049_5611# 0.01824f
C46 XA.XIR[9].XIC[12].icell.Ien Vbias 0.19161f
C47 XThC.Tn[10] XThR.Tn[10] 0.40738f
C48 XThC.Tn[0] XThR.Tn[0] 0.41303f
C49 XThC.Tn[2] XThR.Tn[5] 0.40738f
C50 XThC.Tn[10] XA.XIR[6].XIC[10].icell.PDM 0.02601f
C51 XA.XIR[0].XIC[5].icell.Ien Vbias 0.19213f
C52 XThC.Tn[9] XThC.Tn[10] 0.0671f
C53 XA.XIR[11].XIC[10].icell.Ien Iout 0.06801f
C54 XThR.Tn[13] a_n997_1579# 0.19413f
C55 XA.XIR[12].XIC[2].icell.Ien VPWR 0.18829f
C56 XThR.Tn[9] XA.XIR[10].XIC[11].icell.PDM 0.04035f
C57 XA.XIR[0].XIC_15.icell.PDM VPWR 0.07389f
C58 XThC.XTB7.Y VPWR 1.07721f
C59 XA.XIR[11].XIC[1].icell.Ien XA.XIR[12].XIC[1].icell.PDM 0.02104f
C60 XA.XIR[7].XIC[8].icell.Ien Vbias 0.19161f
C61 XA.XIR[2].XIC[7].icell.Ien XA.XIR[3].XIC[7].icell.PDM 0.02104f
C62 XA.XIR[7].XIC[8].icell.Ien XA.XIR[8].XIC[8].icell.PDM 0.02104f
C63 XThR.Tn[4] XA.XIR[4].XIC[3].icell.Ien 0.14211f
C64 XThC.XTBN.A XThC.XTB6.Y 0.06405f
C65 XThR.XTBN.A XThR.Tn[9] 0.12398f
C66 XA.XIR[11].XIC[0].icell.Ien Iout 0.06795f
C67 XA.XIR[1].XIC[10].icell.Ien XA.XIR[2].XIC[10].icell.PDM 0.02104f
C68 XA.XIR[8].XIC_15.icell.PDM XA.XIR[8].XIC_15.icell.Ien 0.04854f
C69 XA.XIR[10].XIC_dummy_left.icell.PUM VPWR 0.01604f
C70 XThC.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.02602f
C71 XA.XIR[0].XIC[14].icell.Ien XA.XIR[1].XIC[14].icell.PDM 0.02104f
C72 XThR.XTB6.A VPWR 0.68801f
C73 XThC.Tn[8] XThR.Tn[14] 0.40738f
C74 XThR.Tn[7] XA.XIR[8].XIC[1].icell.PDM 0.04035f
C75 XA.XIR[10].XIC[0].icell.Ien Vbias 0.19149f
C76 XA.XIR[6].XIC[8].icell.PDM XA.XIR[6].XIC[8].icell.Ien 0.04854f
C77 XA.XIR[14].XIC[12].icell.Ien Iout 0.06801f
C78 XThR.Tn[1] XA.XIR[2].XIC_dummy_left.icell.Iout 0.01728f
C79 XA.XIR[13].XIC_dummy_left.icell.Ien VPWR 0.39002f
C80 XThC.Tn[0] XA.XIR[4].XIC[0].icell.PDM 0.02601f
C81 XA.XIR[15].XIC[7].icell.PDM XA.XIR[15].XIC[7].icell.Ien 0.04854f
C82 XA.XIR[6].XIC[5].icell.PDM Vbias 0.03928f
C83 XThC.Tn[9] XA.XIR[15].XIC[9].icell.Ien 0.04292f
C84 XThR.XTB1.Y a_n1049_8581# 0.21263f
C85 XA.XIR[5].XIC[12].icell.PDM Vbias 0.03928f
C86 XA.XIR[14].XIC[2].icell.PDM Vbias 0.03928f
C87 XThR.Tn[3] XA.XIR[3].XIC[6].icell.Ien 0.14211f
C88 XThC.Tn[5] XA.XIR[0].XIC[5].icell.Ien 0.04659f
C89 XA.XIR[9].XIC[7].icell.Ien XA.XIR[10].XIC[7].icell.PDM 0.02104f
C90 XThR.XTB7.B data[4] 0.01382f
C91 XA.XIR[10].XIC[2].icell.PDM XA.XIR[10].XIC[2].icell.Ien 0.04854f
C92 XA.XIR[13].XIC[6].icell.PDM Vbias 0.03928f
C93 XA.XIR[9].XIC[4].icell.Ien Iout 0.06801f
C94 XThR.Tn[0] VPWR 8.10551f
C95 XThC.XTB4.Y XThC.XTBN.A 0.03415f
C96 XThR.Tn[3] XA.XIR[4].XIC[2].icell.PDM 0.04035f
C97 XA.XIR[13].XIC_dummy_left.icell.Iout Iout 0.03553f
C98 XThR.XTB7.B XThR.XTB2.Y 0.22599f
C99 XThR.XTB7.B a_n997_3755# 0.01174f
C100 XThC.Tn[4] XThR.Tn[6] 0.40738f
C101 XA.XIR[5].XIC_dummy_right.icell.Iout XA.XIR[6].XIC_dummy_right.icell.Iout 0.04047f
C102 XThR.XTBN.Y XThR.Tn[8] 0.4783f
C103 XA.XIR[6].XIC[6].icell.PDM VPWR 0.01171f
C104 XA.XIR[0].XIC[0].icell.PDM XA.XIR[0].XIC[0].icell.Ien 0.04854f
C105 XA.XIR[5].XIC[13].icell.PDM VPWR 0.01171f
C106 XA.XIR[14].XIC[3].icell.PDM VPWR 0.01171f
C107 XA.XIR[5].XIC[13].icell.Ien Iout 0.06801f
C108 XThC.Tn[7] XA.XIR[4].XIC[7].icell.Ien 0.04604f
C109 XThC.Tn[6] XThR.Tn[11] 0.40738f
C110 XA.XIR[3].XIC[5].icell.Ien Vbias 0.19161f
C111 XA.XIR[13].XIC[7].icell.PDM VPWR 0.01171f
C112 XA.XIR[9].XIC[11].icell.Ien XA.XIR[10].XIC[11].icell.PDM 0.02104f
C113 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.PDM 0.02104f
C114 XThC.Tn[2] Iout 0.22439f
C115 XA.XIR[9].XIC[11].icell.PDM XA.XIR[9].XIC[11].icell.Ien 0.04854f
C116 XThC.XTB3.Y XThC.XTB6.Y 0.04428f
C117 XA.XIR[7].XIC[9].icell.PDM XA.XIR[7].XIC[9].icell.Ien 0.04854f
C118 XA.XIR[9].XIC[3].icell.Ien VPWR 0.18829f
C119 XThC.Tn[1] XA.XIR[11].XIC[1].icell.PDM 0.02601f
C120 XThC.Tn[12] Vbias 0.8219f
C121 XA.XIR[3].XIC[7].icell.PDM Vbias 0.03928f
C122 XA.XIR[4].XIC[14].icell.Ien Vbias 0.19161f
C123 XA.XIR[8].XIC[9].icell.PDM Vbias 0.03928f
C124 XA.XIR[11].XIC_15.icell.Ien Iout 0.0694f
C125 VPWR data[7] 0.212f
C126 XA.XIR[4].XIC[10].icell.PDM XA.XIR[4].XIC[10].icell.Ien 0.04854f
C127 XA.XIR[12].XIC[8].icell.Ien Iout 0.06801f
C128 XThR.XTB4.Y XThR.Tn[8] 0.01306f
C129 XThC.Tn[0] XA.XIR[1].XIC[0].icell.Ien 0.04606f
C130 XThC.Tn[10] XThR.Tn[13] 0.40738f
C131 XA.XIR[2].XIC[13].icell.PDM Vbias 0.03928f
C132 XThC.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.02601f
C133 XThC.Tn[0] XThR.Tn[1] 0.40748f
C134 XThC.Tn[0] XA.XIR[4].XIC[0].icell.Ien 0.04604f
C135 XA.XIR[8].XIC[8].icell.Ien Vbias 0.19161f
C136 XThC.Tn[12] XA.XIR[2].XIC[12].icell.PDM 0.02602f
C137 XThR.Tn[9] XA.XIR[10].XIC[10].icell.PDM 0.04035f
C138 XA.XIR[1].XIC[0].icell.PDM VPWR 0.01171f
C139 XThC.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.02601f
C140 XA.XIR[1].XIC[3].icell.Ien XA.XIR[2].XIC[3].icell.PDM 0.02104f
C141 XThR.XTB6.Y XThR.Tn[9] 0.0246f
C142 XA.XIR[8].XIC[8].icell.PDM XA.XIR[8].XIC[8].icell.Ien 0.04854f
C143 XA.XIR[10].XIC_15.icell.PDM Vbias 0.03927f
C144 XThR.XTB7.A XThR.Tn[3] 0.0306f
C145 XA.XIR[14].XIC[10].icell.Ien Iout 0.06801f
C146 XA.XIR[11].XIC[14].icell.Ien XA.XIR[12].XIC[14].icell.PDM 0.02104f
C147 XThC.Tn[13] XThR.Tn[9] 0.40739f
C148 XA.XIR[4].XIC[0].icell.PDM VPWR 0.01171f
C149 XThC.Tn[0] XThR.Tn[12] 0.40738f
C150 XThC.Tn[9] XThR.Tn[8] 0.40738f
C151 XA.XIR[5].XIC[12].icell.Ien VPWR 0.18829f
C152 XA.XIR[0].XIC[7].icell.Ien XA.XIR[1].XIC[7].icell.PDM 0.02104f
C153 XA.XIR[3].XIC[8].icell.PDM VPWR 0.01171f
C154 XThC.XTB6.A VPWR 0.68179f
C155 XA.XIR[4].XIC_15.icell.PUM VPWR 0.01655f
C156 XA.XIR[8].XIC[10].icell.PDM VPWR 0.01171f
C157 XThC.XTB7.B XThC.XTB7.Y 0.33493f
C158 XThR.Tn[9] XA.XIR[10].XIC_dummy_left.icell.Iout 0.01779f
C159 XThC.XTBN.A a_7875_9569# 0.01939f
C160 XA.XIR[8].XIC_15.icell.Ien XA.XIR[9].XIC_15.icell.PDM 0.02104f
C161 XThR.XTB7.A XThR.XTB7.Y 0.37429f
C162 XA.XIR[2].XIC[14].icell.PDM VPWR 0.0118f
C163 XA.XIR[0].XIC[10].icell.Ien Vbias 0.19213f
C164 XThC.XTBN.Y XThC.Tn[7] 0.85979f
C165 XA.XIR[11].XIC_dummy_right.icell.Iout Iout 0.01732f
C166 XThR.Tn[12] XA.XIR[13].XIC[4].icell.PDM 0.04035f
C167 XThC.Tn[4] XThR.Tn[4] 0.40738f
C168 XThC.XTB2.Y XThC.XTBN.A 0.04716f
C169 XThC.XTB3.Y XThC.XTB4.Y 2.13136f
C170 XA.XIR[3].XIC[14].icell.Ien XA.XIR[4].XIC[14].icell.PDM 0.02104f
C171 XA.XIR[12].XIC[7].icell.Ien VPWR 0.18829f
C172 XA.XIR[10].XIC_dummy_right.icell.PDM VPWR 0.08209f
C173 XA.XIR[4].XIC[1].icell.Ien Iout 0.06801f
C174 XThC.Tn[5] XA.XIR[3].XIC[5].icell.Ien 0.04604f
C175 XA.XIR[7].XIC_dummy_right.icell.Iout XA.XIR[8].XIC_dummy_right.icell.Iout 0.04047f
C176 XA.XIR[7].XIC[13].icell.Ien Vbias 0.19161f
C177 XThC.Tn[12] XA.XIR[2].XIC[12].icell.Ien 0.04605f
C178 XA.XIR[13].XIC_dummy_left.icell.PUM VPWR 0.01669f
C179 XThR.Tn[4] XA.XIR[4].XIC[8].icell.Ien 0.14211f
C180 XThR.Tn[11] XA.XIR[11].XIC[13].icell.Ien 0.14211f
C181 XThC.XTBN.A data[1] 0.01444f
C182 XA.XIR[13].XIC[0].icell.Ien Vbias 0.19149f
C183 XA.XIR[3].XIC[1].icell.Ien XA.XIR[4].XIC[1].icell.PDM 0.02104f
C184 XA.XIR[15].XIC[3].icell.Ien Iout 0.07192f
C185 XA.XIR[6].XIC_dummy_left.icell.Ien VPWR 0.38995f
C186 XThR.Tn[0] XA.XIR[1].XIC[12].icell.PDM 0.04035f
C187 XThR.Tn[1] XA.XIR[2].XIC[11].icell.PDM 0.04035f
C188 XThC.XTB1.Y XThC.XTB6.Y 0.05752f
C189 XA.XIR[4].XIC[6].icell.Ien Iout 0.06801f
C190 XA.XIR[6].XIC[10].icell.Ien XA.XIR[7].XIC[10].icell.PDM 0.02104f
C191 XA.XIR[1].XIC[0].icell.Ien VPWR 0.18829f
C192 XThR.XTBN.Y XThR.XTB2.Y 0.2075f
C193 XThR.XTBN.Y a_n997_3755# 0.229f
C194 XThR.Tn[2] XA.XIR[2].XIC[1].icell.Ien 0.14211f
C195 XA.XIR[7].XIC[13].icell.PDM Vbias 0.03928f
C196 XA.XIR[9].XIC[4].icell.PDM XA.XIR[9].XIC[4].icell.Ien 0.04854f
C197 XA.XIR[7].XIC[2].icell.PDM XA.XIR[7].XIC[2].icell.Ien 0.04854f
C198 XA.XIR[4].XIC[0].icell.Ien VPWR 0.18829f
C199 XThR.Tn[1] VPWR 8.09427f
C200 XThC.Tn[12] XA.XIR[7].XIC[12].icell.PDM 0.02601f
C201 XA.XIR[4].XIC[3].icell.PDM XA.XIR[4].XIC[3].icell.Ien 0.04854f
C202 XThR.Tn[12] XA.XIR[12].XIC[6].icell.Ien 0.14211f
C203 XThC.XTBN.Y a_3773_9615# 0.08456f
C204 XA.XIR[7].XIC[0].icell.Ien Iout 0.06795f
C205 XThR.Tn[3] XA.XIR[3].XIC[11].icell.Ien 0.14211f
C206 XThR.Tn[12] VPWR 8.99609f
C207 XA.XIR[14].XIC[5].icell.Ien XA.XIR[15].XIC[5].icell.PDM 0.02104f
C208 XA.XIR[13].XIC_dummy_left.icell.Iout XA.XIR[14].XIC_dummy_left.icell.Iout 0.03665f
C209 XA.XIR[9].XIC[9].icell.Ien Iout 0.06801f
C210 XThR.XTBN.Y a_n1049_5611# 0.0768f
C211 XA.XIR[9].XIC_dummy_left.icell.PDM XA.XIR[9].XIC_dummy_left.icell.Ien 0.04854f
C212 a_10915_9569# Vbias 0.01451f
C213 XA.XIR[9].XIC[9].icell.PDM Vbias 0.03928f
C214 XThR.XTB2.Y XThR.XTB4.Y 0.04006f
C215 XThC.Tn[6] XThR.Tn[14] 0.40738f
C216 XA.XIR[0].XIC[1].icell.PDM Vbias 0.03945f
C217 XA.XIR[15].XIC[2].icell.Ien VPWR 0.31713f
C218 XA.XIR[13].XIC[13].icell.PDM XA.XIR[13].XIC[13].icell.Ien 0.04854f
C219 XA.XIR[7].XIC[14].icell.PDM VPWR 0.0118f
C220 XA.XIR[0].XIC[2].icell.Ien Iout 0.0675f
C221 XA.XIR[13].XIC[8].icell.Ien XA.XIR[14].XIC[8].icell.PDM 0.02104f
C222 XThR.Tn[2] XA.XIR[2].XIC[6].icell.Ien 0.14211f
C223 XA.XIR[7].XIC[1].icell.Ien XA.XIR[8].XIC[1].icell.PDM 0.02104f
C224 XThC.Tn[3] XA.XIR[10].XIC[3].icell.Ien 0.04604f
C225 XThC.XTB2.Y XThC.XTB3.Y 2.04808f
C226 XThC.XTB1.Y XThC.XTB4.Y 0.05121f
C227 XA.XIR[13].XIC[9].icell.PDM XA.XIR[13].XIC[9].icell.Ien 0.04854f
C228 XA.XIR[4].XIC[5].icell.Ien VPWR 0.18829f
C229 XA.XIR[8].XIC[8].icell.Ien XA.XIR[9].XIC[8].icell.PDM 0.02104f
C230 XThC.Tn[1] XA.XIR[14].XIC[1].icell.PDM 0.02601f
C231 XA.XIR[7].XIC[5].icell.Ien Iout 0.06801f
C232 XA.XIR[14].XIC_15.icell.Ien Iout 0.0694f
C233 XA.XIR[1].XIC_dummy_left.icell.PDM VPWR 0.08221f
C234 XA.XIR[3].XIC[10].icell.Ien Vbias 0.19161f
C235 XA.XIR[3].XIC[7].icell.Ien XA.XIR[4].XIC[7].icell.PDM 0.02104f
C236 XA.XIR[1].XIC[14].icell.PDM Vbias 0.03928f
C237 XA.XIR[10].XIC[14].icell.PDM Vbias 0.03928f
C238 XA.XIR[9].XIC[10].icell.PDM VPWR 0.01171f
C239 XThC.Tn[6] XA.XIR[5].XIC[6].icell.Ien 0.04604f
C240 XThC.Tn[7] XA.XIR[2].XIC[7].icell.PDM 0.02602f
C241 XThC.Tn[8] VPWR 4.5473f
C242 XA.XIR[4].XIC_dummy_left.icell.PDM VPWR 0.08221f
C243 XA.XIR[0].XIC[2].icell.PDM VPWR 0.01132f
C244 XA.XIR[3].XIC[9].icell.PDM XA.XIR[3].XIC[9].icell.Ien 0.04854f
C245 XThC.Tn[0] XA.XIR[5].XIC[0].icell.PDM 0.02601f
C246 XA.XIR[4].XIC[14].icell.PDM Vbias 0.03928f
C247 XA.XIR[2].XIC[3].icell.Ien Vbias 0.19161f
C248 XThR.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.14211f
C249 XA.XIR[9].XIC[8].icell.Ien VPWR 0.18829f
C250 XA.XIR[6].XIC[1].icell.PDM XA.XIR[6].XIC[1].icell.Ien 0.04854f
C251 XA.XIR[13].XIC_15.icell.PDM Vbias 0.03927f
C252 XA.XIR[1].XIC[5].icell.Ien Vbias 0.19173f
C253 XThR.XTB7.B XThR.XTB7.Y 0.33493f
C254 XA.XIR[15].XIC[0].icell.PDM XA.XIR[15].XIC[0].icell.Ien 0.04854f
C255 XThR.Tn[9] XA.XIR[9].XIC[4].icell.Ien 0.14211f
C256 XThC.XTB6.A XThC.XTB7.B 1.47641f
C257 XThC.Tn[2] XA.XIR[7].XIC[2].icell.Ien 0.04604f
C258 XThR.XTB5.Y a_n1319_6405# 0.01188f
C259 XThR.Tn[4] XA.XIR[5].XIC[9].icell.PDM 0.04035f
C260 XA.XIR[8].XIC[13].icell.Ien Vbias 0.19161f
C261 XA.XIR[14].XIC[1].icell.Ien XA.XIR[15].XIC[1].icell.PDM 0.02104f
C262 a_n1049_5317# VPWR 0.72036f
C263 XA.XIR[1].XIC_15.icell.PDM VPWR 0.07527f
C264 XA.XIR[14].XIC_dummy_right.icell.Iout Iout 0.01732f
C265 XThC.Tn[1] Vbias 0.8372f
C266 XA.XIR[4].XIC_15.icell.PDM VPWR 0.07527f
C267 XA.XIR[7].XIC[4].icell.Ien VPWR 0.18829f
C268 XA.XIR[10].XIC[11].icell.PDM XA.XIR[10].XIC[11].icell.Ien 0.04854f
C269 XA.XIR[6].XIC[3].icell.Ien XA.XIR[7].XIC[3].icell.PDM 0.02104f
C270 XThR.Tn[2] XThR.Tn[3] 0.15335f
C271 XA.XIR[13].XIC_dummy_right.icell.PDM VPWR 0.08209f
C272 XA.XIR[11].XIC_15.icell.Ien XA.XIR[12].XIC_15.icell.PDM 0.02104f
C273 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.Iout 0.06446f
C274 XThR.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.14251f
C275 XA.XIR[0].XIC_15.icell.Ien Vbias 0.19241f
C276 XThR.Tn[8] XA.XIR[9].XIC[14].icell.PDM 0.04056f
C277 XThC.Tn[2] XThR.Tn[9] 0.40738f
C278 XThR.XTBN.Y a_n997_715# 0.21503f
C279 XThC.Tn[4] XA.XIR[9].XIC[4].icell.Ien 0.04604f
C280 XThR.Tn[7] XA.XIR[7].XIC[1].icell.Ien 0.14211f
C281 XA.XIR[6].XIC[0].icell.Ien Vbias 0.19149f
C282 XThC.Tn[7] XThR.Tn[8] 0.40738f
C283 XA.XIR[1].XIC[14].icell.PDM XA.XIR[1].XIC[14].icell.Ien 0.04854f
C284 XA.XIR[4].XIC[10].icell.Ien XA.XIR[5].XIC[10].icell.PDM 0.02104f
C285 XThC.XTB1.Y XThC.XTB2.Y 2.14864f
C286 XThC.Tn[11] XA.XIR[0].XIC[11].icell.Ien 0.04662f
C287 XThR.Tn[4] XA.XIR[4].XIC[13].icell.Ien 0.14211f
C288 XThR.Tn[5] XA.XIR[6].XIC[11].icell.PDM 0.04035f
C289 XA.XIR[11].XIC[4].icell.PDM Vbias 0.03928f
C290 XA.XIR[0].XIC_dummy_right.icell.PUM VPWR 0.01499f
C291 XA.XIR[3].XIC[2].icell.Ien Iout 0.06801f
C292 XA.XIR[13].XIC[2].icell.PDM XA.XIR[13].XIC[2].icell.Ien 0.04854f
C293 XThR.Tn[0] XA.XIR[0].XIC[5].icell.Ien 0.14211f
C294 XThR.Tn[2] XA.XIR[3].XIC[3].icell.PDM 0.04035f
C295 XThR.XTB7.B a_n997_2667# 0.02071f
C296 XThC.Tn[5] XA.XIR[1].XIC[5].icell.Ien 0.04606f
C297 XThR.Tn[10] XA.XIR[10].XIC[4].icell.Ien 0.14211f
C298 XThC.Tn[7] XA.XIR[7].XIC[7].icell.PDM 0.02601f
C299 XA.XIR[10].XIC[8].icell.PDM Vbias 0.03928f
C300 XThC.Tn[13] XA.XIR[10].XIC[13].icell.Ien 0.04604f
C301 XA.XIR[5].XIC[0].icell.PDM VPWR 0.01171f
C302 XA.XIR[12].XIC[3].icell.Ien XA.XIR[13].XIC[3].icell.PDM 0.02104f
C303 XA.XIR[15].XIC[8].icell.Ien Iout 0.07192f
C304 XThR.Tn[6] XA.XIR[7].XIC[10].icell.PDM 0.04035f
C305 XThC.Tn[11] XA.XIR[11].XIC[11].icell.Ien 0.04604f
C306 XA.XIR[4].XIC[11].icell.Ien Iout 0.06801f
C307 XA.XIR[6].XIC[5].icell.Ien Vbias 0.19161f
C308 a_n1049_6405# VPWR 0.72095f
C309 XThR.Tn[7] XA.XIR[7].XIC[6].icell.Ien 0.14211f
C310 XA.XIR[8].XIC[1].icell.PDM XA.XIR[8].XIC[1].icell.Ien 0.04854f
C311 XA.XIR[8].XIC_dummy_left.icell.Ien XThR.Tn[8] 0.0125f
C312 XA.XIR[3].XIC[2].icell.PDM XA.XIR[3].XIC[2].icell.Ien 0.04854f
C313 XThC.Tn[13] XA.XIR[4].XIC[13].icell.Ien 0.04604f
C314 XThC.Tn[13] XA.XIR[12].XIC[13].icell.PDM 0.02601f
C315 XA.XIR[0].XIC[0].icell.Ien XA.XIR[1].XIC[0].icell.PDM 0.02104f
C316 XA.XIR[8].XIC[5].icell.Ien Iout 0.06801f
C317 XA.XIR[11].XIC[5].icell.PDM VPWR 0.01171f
C318 XA.XIR[11].XIC[7].icell.PDM XA.XIR[11].XIC[7].icell.Ien 0.04854f
C319 XA.XIR[10].XIC[9].icell.PDM VPWR 0.01171f
C320 VPWR data[3] 0.20846f
C321 XThC.Tn[1] XA.XIR[12].XIC[1].icell.Ien 0.04604f
C322 XA.XIR[12].XIC_dummy_left.icell.PDM XA.XIR[12].XIC_dummy_left.icell.Ien 0.04854f
C323 XA.XIR[2].XIC[0].icell.PDM Vbias 0.03915f
C324 XThC.Tn[3] XA.XIR[13].XIC[3].icell.Ien 0.04604f
C325 XA.XIR[9].XIC[0].icell.Ien XA.XIR[10].XIC[0].icell.PDM 0.02104f
C326 XThR.XTBN.Y XThR.Tn[3] 0.62501f
C327 XA.XIR[10].XIC[13].icell.PDM Vbias 0.03928f
C328 XA.XIR[11].XIC_dummy_left.icell.Ien XThR.Tn[11] 0.01244f
C329 XA.XIR[9].XIC[14].icell.Ien Iout 0.06801f
C330 a_n1049_8581# XThR.Tn[0] 0.2685f
C331 XThR.XTB7.B XThR.Tn[11] 0.03888f
C332 XThC.Tn[10] XThR.Tn[7] 0.40738f
C333 XA.XIR[15].XIC[7].icell.Ien VPWR 0.31713f
C334 XA.XIR[11].XIC[4].icell.Ien Vbias 0.19161f
C335 XA.XIR[0].XIC[7].icell.Ien Iout 0.0675f
C336 XThC.Tn[0] XA.XIR[2].XIC[0].icell.Ien 0.04605f
C337 XA.XIR[0].XIC_dummy_left.icell.PDM XA.XIR[0].XIC_dummy_left.icell.Ien 0.04854f
C338 XThC.Tn[2] XA.XIR[8].XIC[2].icell.Ien 0.04604f
C339 XThC.XTB7.B XThC.Tn[8] 0.05151f
C340 XThR.Tn[2] XA.XIR[2].XIC[11].icell.Ien 0.14211f
C341 XA.XIR[13].XIC[14].icell.PDM Vbias 0.03928f
C342 XThR.XTBN.Y XThR.XTB7.Y 0.50018f
C343 XA.XIR[7].XIC_dummy_left.icell.Ien VPWR 0.38902f
C344 XA.XIR[10].XIC[6].icell.Ien Vbias 0.19161f
C345 XThC.XTB7.Y XThC.Tn[12] 0.07091f
C346 XA.XIR[4].XIC[10].icell.Ien VPWR 0.18829f
C347 XA.XIR[0].XIC[1].icell.Ien VPWR 0.18776f
C348 XA.XIR[2].XIC[1].icell.PDM VPWR 0.01171f
C349 XA.XIR[7].XIC[10].icell.Ien Iout 0.06801f
C350 XA.XIR[14].XIC[14].icell.Ien XA.XIR[15].XIC[14].icell.PDM 0.02104f
C351 XA.XIR[8].XIC[4].icell.Ien VPWR 0.18829f
C352 XA.XIR[3].XIC_15.icell.Ien Vbias 0.19195f
C353 XThR.XTB4.Y XThR.Tn[3] 0.1895f
C354 XA.XIR[1].XIC[7].icell.PDM XA.XIR[1].XIC[7].icell.Ien 0.04854f
C355 XA.XIR[4].XIC[3].icell.Ien XA.XIR[5].XIC[3].icell.PDM 0.02104f
C356 XA.XIR[2].XIC[8].icell.Ien Vbias 0.19161f
C357 XThR.Tn[11] XA.XIR[12].XIC[1].icell.PDM 0.04035f
C358 XThC.Tn[5] XA.XIR[6].XIC[5].icell.Ien 0.04604f
C359 XA.XIR[8].XIC[0].icell.Ien Iout 0.06795f
C360 XA.XIR[9].XIC[13].icell.Ien VPWR 0.18829f
C361 XA.XIR[1].XIC[10].icell.Ien Vbias 0.19173f
C362 XThR.XTB4.Y XThR.XTB7.Y 0.03475f
C363 XThC.Tn[11] XA.XIR[3].XIC[11].icell.Ien 0.04604f
C364 XThR.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.14211f
C365 XA.XIR[0].XIC[6].icell.Ien VPWR 0.1878f
C366 XThC.Tn[9] XThR.Tn[3] 0.40738f
C367 XA.XIR[2].XIC[9].icell.PDM XA.XIR[2].XIC[9].icell.Ien 0.04854f
C368 XA.XIR[2].XIC_dummy_left.icell.PUM VPWR 0.01604f
C369 XThC.Tn[6] XA.XIR[12].XIC[6].icell.Ien 0.04604f
C370 XThR.XTB7.Y XThR.Tn[10] 0.07406f
C371 XA.XIR[3].XIC_dummy_right.icell.PUM VPWR 0.01691f
C372 XThC.Tn[6] VPWR 3.63495f
C373 XA.XIR[10].XIC_dummy_right.icell.PDM XA.XIR[10].XIC_dummy_right.icell.Ien 0.04854f
C374 XThR.Tn[5] XA.XIR[5].XIC[0].icell.Ien 0.1423f
C375 XA.XIR[7].XIC[9].icell.Ien VPWR 0.18829f
C376 XThR.Tn[14] XA.XIR[14].XIC[13].icell.Ien 0.14211f
C377 XThC.Tn[12] XThR.Tn[0] 0.40763f
C378 XA.XIR[7].XIC[0].icell.PDM Vbias 0.03915f
C379 XThC.Tn[14] XThR.Tn[5] 0.40742f
C380 XThR.Tn[7] XA.XIR[8].XIC[3].icell.PDM 0.04035f
C381 XThR.XTBN.Y a_n997_2667# 0.22784f
C382 XA.XIR[9].XIC_dummy_left.icell.Iout XA.XIR[10].XIC_dummy_left.icell.Iout 0.03665f
C383 XA.XIR[6].XIC[7].icell.PDM Vbias 0.03928f
C384 XA.XIR[5].XIC_dummy_left.icell.PDM VPWR 0.08221f
C385 XA.XIR[8].XIC[1].icell.Ien XA.XIR[9].XIC[1].icell.PDM 0.02104f
C386 XA.XIR[11].XIC[12].icell.Ien XA.XIR[12].XIC[12].icell.PDM 0.02104f
C387 XThR.Tn[8] a_n997_3979# 0.1927f
C388 XA.XIR[14].XIC[4].icell.PDM Vbias 0.03928f
C389 XA.XIR[5].XIC[14].icell.PDM Vbias 0.03928f
C390 XA.XIR[5].XIC[12].icell.PDM XA.XIR[5].XIC[12].icell.Ien 0.04854f
C391 XA.XIR[2].XIC[0].icell.Ien VPWR 0.18829f
C392 XThC.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.04604f
C393 XA.XIR[13].XIC[8].icell.PDM Vbias 0.03928f
C394 XThC.Tn[2] XA.XIR[6].XIC[2].icell.PDM 0.02601f
C395 XThR.Tn[3] XA.XIR[4].XIC[4].icell.PDM 0.04035f
C396 XThR.Tn[11] XA.XIR[11].XIC[5].icell.Ien 0.14211f
C397 XThC.Tn[9] XA.XIR[2].XIC[9].icell.PDM 0.02602f
C398 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Ien 0.01557f
C399 XA.XIR[10].XIC[1].icell.Ien VPWR 0.18829f
C400 XThC.Tn[11] XA.XIR[14].XIC[11].icell.Ien 0.04604f
C401 XA.XIR[7].XIC[1].icell.PDM VPWR 0.01171f
C402 XThR.XTB4.Y a_n997_2667# 0.07199f
C403 XA.XIR[3].XIC[7].icell.Ien Iout 0.06801f
C404 XThR.Tn[10] XA.XIR[10].XIC[9].icell.Ien 0.14211f
C405 XA.XIR[6].XIC[8].icell.PDM VPWR 0.01171f
C406 XThR.Tn[0] XA.XIR[0].XIC[10].icell.Ien 0.14211f
C407 XThC.Tn[13] XA.XIR[15].XIC[13].icell.PDM 0.02601f
C408 XA.XIR[5].XIC_15.icell.PDM VPWR 0.07527f
C409 XThR.Tn[6] XA.XIR[6].XIC[4].icell.Ien 0.14211f
C410 XA.XIR[14].XIC[5].icell.PDM VPWR 0.01171f
C411 XThC.Tn[9] XA.XIR[10].XIC[9].icell.Ien 0.04604f
C412 XThR.XTBN.Y XThR.Tn[11] 0.52268f
C413 XA.XIR[5].XIC_dummy_right.icell.PDM XA.XIR[5].XIC_dummy_right.icell.Ien 0.04854f
C414 XA.XIR[10].XIC[12].icell.PDM Vbias 0.03928f
C415 XThC.Tn[11] XThR.Tn[2] 0.40741f
C416 XA.XIR[13].XIC[9].icell.PDM VPWR 0.01171f
C417 XA.XIR[1].XIC[1].icell.PDM Vbias 0.03928f
C418 XA.XIR[12].XIC[8].icell.PDM XA.XIR[12].XIC[8].icell.Ien 0.04854f
C419 XA.XIR[6].XIC[10].icell.Ien Vbias 0.19161f
C420 XThR.Tn[7] XA.XIR[7].XIC[11].icell.Ien 0.14211f
C421 XA.XIR[1].XIC[2].icell.Ien Iout 0.06801f
C422 XThC.XTB7.Y a_10915_9569# 0.06874f
C423 XA.XIR[13].XIC[13].icell.PDM Vbias 0.03928f
C424 XThR.XTB7.A XThR.XTB3.Y 0.57441f
C425 XA.XIR[4].XIC[1].icell.PDM Vbias 0.03928f
C426 XA.XIR[7].XIC_dummy_left.icell.PUM VPWR 0.01604f
C427 XA.XIR[8].XIC[10].icell.Ien Iout 0.06801f
C428 data[5] data[6] 0.01513f
C429 XThC.Tn[12] XA.XIR[5].XIC[12].icell.Ien 0.04604f
C430 XA.XIR[3].XIC[9].icell.PDM Vbias 0.03928f
C431 XA.XIR[8].XIC[11].icell.PDM Vbias 0.03928f
C432 XA.XIR[14].XIC[4].icell.Ien Vbias 0.19161f
C433 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.Iout 0.06446f
C434 XThR.Tn[7] XThR.Tn[8] 0.12208f
C435 XA.XIR[11].XIC[13].icell.Ien VPWR 0.18829f
C436 XA.XIR[2].XIC_15.icell.PDM Vbias 0.03927f
C437 XA.XIR[5].XIC[0].icell.Ien XA.XIR[6].XIC[0].icell.PDM 0.02104f
C438 XA.XIR[13].XIC[6].icell.Ien Vbias 0.19161f
C439 XA.XIR[2].XIC[2].icell.PDM XA.XIR[2].XIC[2].icell.Ien 0.04854f
C440 XA.XIR[3].XIC[6].icell.Ien VPWR 0.18829f
C441 XThR.Tn[14] XA.XIR[14].XIC[11].icell.Ien 0.14211f
C442 XA.XIR[1].XIC[2].icell.PDM VPWR 0.01171f
C443 XThR.XTB4.Y XThR.Tn[11] 0.3042f
C444 XThC.Tn[8] XA.XIR[7].XIC[8].icell.Ien 0.04604f
C445 XA.XIR[11].XIC[9].icell.Ien Vbias 0.19161f
C446 XA.XIR[0].XIC[12].icell.Ien Iout 0.0675f
C447 XA.XIR[4].XIC[2].icell.PDM VPWR 0.01171f
C448 XThR.Tn[10] XThR.Tn[11] 0.10691f
C449 XA.XIR[3].XIC[10].icell.PDM VPWR 0.01171f
C450 XA.XIR[4].XIC_15.icell.Ien VPWR 0.26829f
C451 XA.XIR[8].XIC[12].icell.PDM VPWR 0.01171f
C452 XThC.XTB5.Y XThC.XTBN.Y 0.162f
C453 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[14].XIC_dummy_left.icell.Iout 0.06446f
C454 XThC.Tn[9] XThR.Tn[11] 0.40738f
C455 XA.XIR[2].XIC_dummy_right.icell.PDM VPWR 0.08209f
C456 XThC.XTBN.A a_8963_9569# 0.01679f
C457 XThR.Tn[8] XA.XIR[9].XIC[1].icell.PDM 0.04035f
C458 XThR.Tn[12] XA.XIR[13].XIC[6].icell.PDM 0.04035f
C459 XA.XIR[7].XIC_15.icell.Ien Iout 0.0694f
C460 XA.XIR[8].XIC[9].icell.Ien VPWR 0.18829f
C461 XThC.Tn[9] XA.XIR[7].XIC[9].icell.PDM 0.02601f
C462 XA.XIR[13].XIC[11].icell.PDM XA.XIR[13].XIC[11].icell.Ien 0.04854f
C463 XA.XIR[5].XIC[0].icell.Ien Iout 0.06795f
C464 XA.XIR[14].XIC_15.icell.Ien XA.XIR[15].XIC_15.icell.PDM 0.02104f
C465 XA.XIR[5].XIC[5].icell.PDM XA.XIR[5].XIC[5].icell.Ien 0.04854f
C466 XThR.XTB7.Y XThR.Tn[13] 0.10781f
C467 XA.XIR[4].XIC_dummy_left.icell.Iout Iout 0.03553f
C468 XA.XIR[2].XIC[13].icell.Ien Vbias 0.19161f
C469 XThC.Tn[14] Iout 0.22441f
C470 XThC.XTB7.B XThC.Tn[6] 0.04318f
C471 XThC.XTB5.Y XThC.Tn[10] 0.01755f
C472 XA.XIR[1].XIC_15.icell.Ien Vbias 0.19206f
C473 XThC.Tn[10] XA.XIR[9].XIC[10].icell.Ien 0.04604f
C474 XThR.Tn[9] XA.XIR[9].XIC[14].icell.Ien 0.144f
C475 XA.XIR[0].XIC_15.icell.PDM XA.XIR[0].XIC_15.icell.Ien 0.04854f
C476 XA.XIR[0].XIC[11].icell.Ien VPWR 0.18882f
C477 XThR.Tn[12] XA.XIR[12].XIC_dummy_left.icell.Iout 0.03385f
C478 XA.XIR[4].XIC_dummy_right.icell.Iout VPWR 0.11567f
C479 XA.XIR[6].XIC[2].icell.Ien Iout 0.06801f
C480 XThC.Tn[12] XThR.Tn[1] 0.40744f
C481 XThR.Tn[0] XA.XIR[1].XIC[14].icell.PDM 0.04056f
C482 XA.XIR[7].XIC_dummy_right.icell.Iout Iout 0.01732f
C483 bias[1] Vbias 0.68866f
C484 XA.XIR[6].XIC_dummy_left.icell.Iout XA.XIR[7].XIC_dummy_left.icell.Iout 0.03665f
C485 XThC.Tn[11] XA.XIR[1].XIC[11].icell.Ien 0.04606f
C486 XThR.Tn[1] XA.XIR[2].XIC[13].icell.PDM 0.0404f
C487 XThC.Tn[12] XThR.Tn[12] 0.40738f
C488 XA.XIR[7].XIC[14].icell.Ien VPWR 0.18835f
C489 XThR.XTB5.Y XThR.XTBN.A 0.10854f
C490 XThR.XTB7.A VPWR 0.88595f
C491 XThR.Tn[10] XA.XIR[10].XIC[14].icell.Ien 0.144f
C492 XThR.Tn[13] XA.XIR[13].XIC[4].icell.Ien 0.14211f
C493 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Iout 0.03842f
C494 XThC.Tn[4] XA.XIR[2].XIC[4].icell.PDM 0.02602f
C495 XA.XIR[1].XIC_dummy_right.icell.PUM VPWR 0.01691f
C496 XA.XIR[5].XIC[3].icell.Ien Vbias 0.19161f
C497 XA.XIR[11].XIC[11].icell.Ien VPWR 0.18829f
C498 XA.XIR[7].XIC_15.icell.PDM Vbias 0.03927f
C499 XThC.Tn[7] XThR.Tn[3] 0.40738f
C500 XThC.XTBN.Y XThC.Tn[10] 0.4511f
C501 XThC.Tn[7] XA.XIR[12].XIC[7].icell.PDM 0.02601f
C502 XA.XIR[5].XIC[14].icell.Ien XA.XIR[6].XIC[14].icell.PDM 0.02104f
C503 XA.XIR[13].XIC[1].icell.Ien VPWR 0.18829f
C504 XThC.XTBN.Y a_4861_9615# 0.07601f
C505 XA.XIR[10].XIC[11].icell.PDM Vbias 0.03928f
C506 XThC.Tn[13] XA.XIR[0].XIC[13].icell.PDM 0.0279f
C507 XThC.Tn[1] XThR.Tn[0] 0.40762f
C508 XThC.Tn[11] XThR.Tn[10] 0.40738f
C509 XA.XIR[10].XIC[3].icell.Ien Iout 0.06801f
C510 XA.XIR[14].XIC[7].icell.PDM XA.XIR[14].XIC[7].icell.Ien 0.04854f
C511 XThC.Tn[3] XThR.Tn[5] 0.40738f
C512 XThR.XTB7.B XThR.XTB3.Y 0.23315f
C513 XA.XIR[9].XIC[11].icell.PDM Vbias 0.03928f
C514 XA.XIR[13].XIC[12].icell.PDM Vbias 0.03928f
C515 XThC.XTB5.Y a_5155_10571# 0.01188f
C516 XA.XIR[11].XIC_dummy_left.icell.PDM XA.XIR[11].XIC_dummy_left.icell.Ien 0.04854f
C517 XThC.Tn[9] XA.XIR[13].XIC[9].icell.Ien 0.04604f
C518 XA.XIR[0].XIC[3].icell.PDM Vbias 0.03945f
C519 XThR.XTBN.Y XThR.Tn[14] 0.47807f
C520 XA.XIR[7].XIC_dummy_right.icell.PDM VPWR 0.08209f
C521 XThR.Tn[0] XA.XIR[0].XIC_15.icell.Ien 0.13564f
C522 XA.XIR[3].XIC[12].icell.Ien Iout 0.06801f
C523 XThC.Tn[6] XA.XIR[10].XIC[6].icell.PDM 0.02601f
C524 XThR.Tn[6] XA.XIR[6].XIC[9].icell.Ien 0.14211f
C525 XThC.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.04604f
C526 XA.XIR[2].XIC[5].icell.Ien Iout 0.06801f
C527 XA.XIR[11].XIC[14].icell.Ien Vbias 0.19161f
C528 XThR.Tn[6] Vbias 1.39526f
C529 XA.XIR[14].XIC[13].icell.Ien VPWR 0.18883f
C530 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.PDM 0.02104f
C531 XA.XIR[1].XIC[7].icell.Ien Iout 0.06801f
C532 XThC.Tn[6] XA.XIR[15].XIC[6].icell.Ien 0.04292f
C533 XA.XIR[6].XIC_15.icell.Ien Vbias 0.19195f
C534 XA.XIR[9].XIC[12].icell.PDM VPWR 0.01171f
C535 XThR.XTB1.Y XThR.XTBN.A 0.12307f
C536 XA.XIR[0].XIC[4].icell.PDM VPWR 0.01136f
C537 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.Iout 0.06446f
C538 XA.XIR[1].XIC[1].icell.Ien VPWR 0.18829f
C539 XA.XIR[8].XIC_15.icell.Ien Iout 0.0694f
C540 XThR.XTB3.Y XThR.Tn[2] 0.18254f
C541 XA.XIR[10].XIC[2].icell.Ien VPWR 0.18829f
C542 XA.XIR[14].XIC[9].icell.Ien Vbias 0.19161f
C543 XThC.Tn[7] XA.XIR[11].XIC[7].icell.Ien 0.04604f
C544 XA.XIR[0].XIC[8].icell.PDM XA.XIR[0].XIC[8].icell.Ien 0.04854f
C545 XThC.Tn[0] XThR.Tn[2] 0.40744f
C546 XThR.Tn[10] XA.XIR[11].XIC[0].icell.PDM 0.04035f
C547 XThC.Tn[11] XA.XIR[6].XIC[11].icell.Ien 0.04604f
C548 XThC.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.04605f
C549 XThR.Tn[4] XA.XIR[5].XIC[11].icell.PDM 0.04035f
C550 XThR.XTB5.Y XThR.Tn[4] 0.19957f
C551 XThR.Tn[14] XA.XIR[15].XIC[1].icell.PDM 0.04035f
C552 XA.XIR[3].XIC[11].icell.Ien VPWR 0.18829f
C553 XA.XIR[6].XIC_dummy_right.icell.PUM VPWR 0.01691f
C554 XThR.Tn[10] XA.XIR[10].XIC[12].icell.Ien 0.14211f
C555 XThC.Tn[9] XThR.Tn[14] 0.40738f
C556 XThC.Tn[4] XA.XIR[7].XIC[4].icell.PDM 0.02601f
C557 XA.XIR[2].XIC[4].icell.Ien VPWR 0.18829f
C558 XThR.Tn[1] a_n1049_7787# 0.26879f
C559 XA.XIR[1].XIC[6].icell.Ien VPWR 0.18829f
C560 XThR.XTB5.Y XThR.XTB6.Y 2.12831f
C561 XA.XIR[8].XIC_dummy_right.icell.Iout Iout 0.01732f
C562 XA.XIR[5].XIC[7].icell.Ien XA.XIR[6].XIC[7].icell.PDM 0.02104f
C563 XA.XIR[13].XIC_dummy_right.icell.PDM XA.XIR[13].XIC_dummy_right.icell.Ien 0.04854f
C564 XA.XIR[8].XIC[14].icell.Ien VPWR 0.18835f
C565 XA.XIR[5].XIC[1].icell.PDM Vbias 0.03928f
C566 XA.XIR[11].XIC_dummy_left.icell.Ien VPWR 0.38914f
C567 XThC.Tn[5] XThR.Tn[6] 0.40738f
C568 XThR.Tn[7] XA.XIR[7].XIC_dummy_left.icell.Iout 0.0402f
C569 XThR.XTB7.B VPWR 1.67716f
C570 XThR.Tn[4] Vbias 1.39526f
C571 XA.XIR[12].XIC[0].icell.PDM Vbias 0.03915f
C572 XA.XIR[14].XIC[12].icell.Ien XA.XIR[15].XIC[12].icell.PDM 0.02104f
C573 XThR.Tn[5] XA.XIR[6].XIC[13].icell.PDM 0.0404f
C574 XA.XIR[2].XIC_15.icell.Ien XA.XIR[3].XIC_15.icell.PDM 0.02104f
C575 XThC.Tn[7] XThR.Tn[11] 0.40738f
C576 XA.XIR[11].XIC[6].icell.PDM Vbias 0.03928f
C577 XA.XIR[11].XIC[12].icell.Ien Vbias 0.19161f
C578 XThR.Tn[2] XA.XIR[3].XIC[5].icell.PDM 0.04035f
C579 XA.XIR[6].XIC[7].icell.Ien Iout 0.06801f
C580 XA.XIR[14].XIC[11].icell.Ien VPWR 0.18883f
C581 XThR.Tn[1] XA.XIR[1].XIC[5].icell.Ien 0.14211f
C582 XThR.Tn[14] XA.XIR[14].XIC[5].icell.Ien 0.14211f
C583 XA.XIR[10].XIC[10].icell.PDM Vbias 0.03928f
C584 XA.XIR[5].XIC[2].icell.PDM VPWR 0.01171f
C585 XThC.Tn[3] Iout 0.22443f
C586 XThC.Tn[7] XA.XIR[15].XIC[7].icell.PDM 0.02601f
C587 XThR.XTBN.Y XThR.XTB3.Y 0.17246f
C588 XA.XIR[6].XIC[1].icell.Ien VPWR 0.18829f
C589 XThR.Tn[6] XA.XIR[7].XIC[12].icell.PDM 0.04035f
C590 XThC.Tn[13] Vbias 0.82511f
C591 XThC.Tn[10] XA.XIR[12].XIC[10].icell.Ien 0.04604f
C592 XA.XIR[13].XIC[11].icell.PDM Vbias 0.03928f
C593 XThR.Tn[13] XA.XIR[13].XIC[9].icell.Ien 0.14211f
C594 XA.XIR[12].XIC[1].icell.PDM VPWR 0.01171f
C595 XA.XIR[11].XIC[6].icell.Ien XA.XIR[12].XIC[6].icell.PDM 0.02104f
C596 XThC.Tn[11] XThR.Tn[13] 0.40738f
C597 XThR.Tn[2] VPWR 8.04926f
C598 XA.XIR[13].XIC[3].icell.Ien Iout 0.06801f
C599 XA.XIR[5].XIC[8].icell.Ien Vbias 0.19161f
C600 XThC.Tn[1] XThR.Tn[1] 0.40744f
C601 XA.XIR[10].XIC[13].icell.Ien XA.XIR[11].XIC[13].icell.PDM 0.02104f
C602 XA.XIR[11].XIC[7].icell.PDM VPWR 0.01171f
C603 XThR.XTB1.Y XThR.XTB6.Y 0.05751f
C604 XThR.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.14211f
C605 XA.XIR[10].XIC[9].icell.Ien XA.XIR[11].XIC[9].icell.PDM 0.02104f
C606 XA.XIR[2].XIC[2].icell.PDM Vbias 0.03928f
C607 XThC.Tn[14] XThR.Tn[9] 0.40742f
C608 XA.XIR[11].XIC[6].icell.Ien Iout 0.06801f
C609 XThC.Tn[1] XThR.Tn[12] 0.40738f
C610 XThC.Tn[6] XA.XIR[13].XIC[6].icell.PDM 0.02601f
C611 XThC.Tn[10] XThR.Tn[8] 0.40738f
C612 XThR.XTB3.Y XThR.XTB4.Y 2.13136f
C613 XA.XIR[12].XIC[3].icell.Ien Vbias 0.19161f
C614 XA.XIR[6].XIC[6].icell.Ien VPWR 0.18829f
C615 XA.XIR[10].XIC[8].icell.Ien Iout 0.06801f
C616 XA.XIR[14].XIC[14].icell.Ien Vbias 0.19161f
C617 XA.XIR[11].XIC[10].icell.Ien XA.XIR[12].XIC[10].icell.PDM 0.02104f
C618 XThC.Tn[5] XThR.Tn[4] 0.40738f
C619 XThC.XTBN.Y a_7651_9569# 0.23021f
C620 XThR.XTB3.Y XThR.Tn[10] 0.29462f
C621 XA.XIR[0].XIC_dummy_left.icell.Iout VPWR 0.1175f
C622 XThC.XTB4.Y XThC.Tn[3] 0.1917f
C623 XThR.Tn[6] XA.XIR[6].XIC[14].icell.Ien 0.144f
C624 XThC.Tn[0] XThR.Tn[10] 0.40734f
C625 XA.XIR[14].XIC[0].icell.Ien XThR.Tn[14] 0.14211f
C626 XA.XIR[2].XIC[3].icell.PDM VPWR 0.01171f
C627 XA.XIR[2].XIC[10].icell.Ien Iout 0.06801f
C628 XA.XIR[13].XIC[2].icell.Ien VPWR 0.18829f
C629 XThC.Tn[7] XA.XIR[14].XIC[7].icell.Ien 0.04604f
C630 XA.XIR[3].XIC_dummy_left.icell.PDM XA.XIR[3].XIC_dummy_left.icell.Ien 0.04854f
C631 XThR.Tn[13] XThR.Tn[14] 0.20347f
C632 XA.XIR[1].XIC[12].icell.Ien Iout 0.06801f
C633 XThR.Tn[11] XA.XIR[12].XIC[3].icell.PDM 0.04035f
C634 XA.XIR[11].XIC[5].icell.Ien VPWR 0.18829f
C635 XA.XIR[11].XIC[10].icell.Ien Vbias 0.19161f
C636 XThR.Tn[8] XA.XIR[8].XIC[1].icell.Ien 0.14211f
C637 XA.XIR[10].XIC[7].icell.Ien VPWR 0.18829f
C638 XA.XIR[2].XIC[8].icell.Ien XA.XIR[3].XIC[8].icell.PDM 0.02104f
C639 XA.XIR[4].XIC_dummy_right.icell.Ien VPWR 0.35722f
C640 XThR.XTB7.Y XThR.Tn[7] 0.0835f
C641 XA.XIR[7].XIC[9].icell.Ien XA.XIR[8].XIC[9].icell.PDM 0.02104f
C642 XThC.XTB2.Y a_4067_9615# 0.02133f
C643 XThR.Tn[7] XA.XIR[8].XIC_dummy_left.icell.Iout 0.01728f
C644 XThC.Tn[9] XA.XIR[12].XIC[9].icell.PDM 0.02601f
C645 XA.XIR[1].XIC[0].icell.Ien XA.XIR[2].XIC[0].icell.PDM 0.02104f
C646 XThC.XTBN.A Vbias 0.01693f
C647 XThR.Tn[0] XA.XIR[1].XIC[1].icell.PDM 0.04035f
C648 XA.XIR[1].XIC[11].icell.Ien XA.XIR[2].XIC[11].icell.PDM 0.02104f
C649 XA.XIR[11].XIC_dummy_left.icell.PUM VPWR 0.01604f
C650 XThR.XTBN.Y VPWR 4.54558f
C651 XThR.Tn[1] XA.XIR[2].XIC[0].icell.PDM 0.0404f
C652 XA.XIR[2].XIC[9].icell.Ien VPWR 0.18829f
C653 XA.XIR[11].XIC[0].icell.Ien Vbias 0.19149f
C654 XA.XIR[0].XIC_15.icell.Ien XA.XIR[1].XIC_15.icell.PDM 0.02104f
C655 XA.XIR[1].XIC[11].icell.Ien VPWR 0.18829f
C656 XA.XIR[6].XIC[9].icell.PDM XA.XIR[6].XIC[9].icell.Ien 0.04854f
C657 XThR.Tn[8] XA.XIR[8].XIC[6].icell.Ien 0.14211f
C658 XThR.Tn[7] XA.XIR[8].XIC[5].icell.PDM 0.04035f
C659 XA.XIR[7].XIC[2].icell.PDM Vbias 0.03928f
C660 XA.XIR[15].XIC[0].icell.PDM Vbias 0.03915f
C661 XA.XIR[15].XIC[8].icell.PDM XA.XIR[15].XIC[8].icell.Ien 0.04854f
C662 XThC.Tn[3] XA.XIR[4].XIC[3].icell.Ien 0.04604f
C663 XA.XIR[6].XIC[9].icell.PDM Vbias 0.03928f
C664 XThC.Tn[8] XA.XIR[10].XIC[8].icell.PDM 0.02601f
C665 XThC.Tn[7] XThR.Tn[14] 0.40738f
C666 XA.XIR[10].XIC[2].icell.Ien XA.XIR[11].XIC[2].icell.PDM 0.02104f
C667 XA.XIR[14].XIC[6].icell.PDM Vbias 0.03928f
C668 XA.XIR[14].XIC[12].icell.Ien Vbias 0.19161f
C669 XThR.Tn[13] XA.XIR[13].XIC[14].icell.Ien 0.144f
C670 XThC.Tn[14] XA.XIR[12].XIC[14].icell.PDM 0.02601f
C671 a_10051_9569# XThC.Tn[13] 0.1927f
C672 XA.XIR[9].XIC[8].icell.Ien XA.XIR[10].XIC[8].icell.PDM 0.02104f
C673 XThR.XTB4.Y VPWR 0.92827f
C674 XA.XIR[10].XIC[3].icell.PDM XA.XIR[10].XIC[3].icell.Ien 0.04854f
C675 XThR.Tn[12] XA.XIR[13].XIC[14].icell.PDM 0.04056f
C676 XA.XIR[13].XIC[10].icell.PDM Vbias 0.03928f
C677 XA.XIR[12].XIC[13].icell.Ien Iout 0.06801f
C678 XThR.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.14211f
C679 XThR.Tn[3] XA.XIR[4].XIC[6].icell.PDM 0.04035f
C680 XA.XIR[7].XIC[3].icell.PDM VPWR 0.01171f
C681 XThR.Tn[10] XA.XIR[10].XIC_15.icell.Ien 0.13564f
C682 XThR.Tn[10] VPWR 8.95184f
C683 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Ien 0.01557f
C684 XA.XIR[9].XIC[4].icell.Ien Vbias 0.19161f
C685 XA.XIR[15].XIC[1].icell.PDM VPWR 0.01512f
C686 XA.XIR[6].XIC[10].icell.PDM VPWR 0.01171f
C687 XA.XIR[0].XIC[1].icell.PDM XA.XIR[0].XIC[1].icell.Ien 0.04854f
C688 XA.XIR[6].XIC[12].icell.Ien Iout 0.06801f
C689 XThC.Tn[9] VPWR 4.54443f
C690 XThC.Tn[13] XA.XIR[1].XIC[13].icell.PDM 0.02602f
C691 XThR.Tn[1] XA.XIR[1].XIC[10].icell.Ien 0.14211f
C692 XThR.XTB5.A a_n1335_4229# 0.01243f
C693 XA.XIR[14].XIC[7].icell.PDM VPWR 0.01171f
C694 XA.XIR[1].XIC[3].icell.PDM Vbias 0.03928f
C695 XThC.Tn[13] XA.XIR[4].XIC[13].icell.PDM 0.02601f
C696 XA.XIR[14].XIC[6].icell.Ien Iout 0.06801f
C697 XA.XIR[4].XIC[3].icell.PDM Vbias 0.03928f
C698 XA.XIR[5].XIC[13].icell.Ien Vbias 0.19161f
C699 XA.XIR[13].XIC[8].icell.Ien Iout 0.06801f
C700 XA.XIR[9].XIC[12].icell.PDM XA.XIR[9].XIC[12].icell.Ien 0.04854f
C701 XA.XIR[7].XIC[10].icell.PDM XA.XIR[7].XIC[10].icell.Ien 0.04854f
C702 XA.XIR[1].XIC_dummy_left.icell.Iout XA.XIR[2].XIC_dummy_left.icell.Iout 0.03665f
C703 XThC.XTB3.Y Vbias 0.01224f
C704 XA.XIR[3].XIC[11].icell.PDM Vbias 0.03928f
C705 XA.XIR[4].XIC[11].icell.PDM XA.XIR[4].XIC[11].icell.Ien 0.04854f
C706 XThC.XTB7.A XThC.XTB5.Y 0.11935f
C707 XA.XIR[8].XIC[13].icell.PDM Vbias 0.03928f
C708 XA.XIR[7].XIC[2].icell.Ien XA.XIR[8].XIC[2].icell.PDM 0.02104f
C709 XThC.Tn[12] XA.XIR[8].XIC[12].icell.PDM 0.02601f
C710 XThC.Tn[2] Vbias 0.83223f
C711 XA.XIR[1].XIC_dummy_left.icell.PDM XA.XIR[1].XIC_dummy_left.icell.Ien 0.04854f
C712 XThC.Tn[0] XA.XIR[14].XIC[0].icell.Ien 0.04604f
C713 XA.XIR[11].XIC_15.icell.PDM Vbias 0.03927f
C714 XA.XIR[11].XIC_15.icell.Ien Vbias 0.19195f
C715 XA.XIR[1].XIC[4].icell.PDM VPWR 0.01171f
C716 XA.XIR[12].XIC[8].icell.Ien Vbias 0.19161f
C717 XThC.Tn[0] XThR.Tn[13] 0.40741f
C718 XA.XIR[1].XIC[4].icell.Ien XA.XIR[2].XIC[4].icell.PDM 0.02104f
C719 XA.XIR[6].XIC[11].icell.Ien VPWR 0.18829f
C720 XA.XIR[14].XIC[0].icell.PDM XA.XIR[14].XIC[0].icell.Ien 0.04854f
C721 XThC.Tn[8] XA.XIR[2].XIC[8].icell.Ien 0.04605f
C722 XA.XIR[8].XIC[9].icell.PDM XA.XIR[8].XIC[9].icell.Ien 0.04854f
C723 XA.XIR[4].XIC[4].icell.PDM VPWR 0.01171f
C724 XThR.Tn[13] XA.XIR[14].XIC[0].icell.PDM 0.04042f
C725 XA.XIR[9].XIC_dummy_right.icell.PDM XA.XIR[9].XIC_dummy_right.icell.Ien 0.04854f
C726 XA.XIR[4].XIC_dummy_left.icell.PDM XA.XIR[4].XIC_dummy_left.icell.Ien 0.04854f
C727 XA.XIR[0].XIC[8].icell.Ien XA.XIR[1].XIC[8].icell.PDM 0.02104f
C728 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.Iout 0.06446f
C729 XA.XIR[3].XIC[12].icell.PDM VPWR 0.01171f
C730 XThC.Tn[3] XThR.Tn[9] 0.40738f
C731 XA.XIR[8].XIC[14].icell.PDM VPWR 0.0118f
C732 XA.XIR[6].XIC[2].icell.PDM XA.XIR[6].XIC[2].icell.Ien 0.04854f
C733 XA.XIR[14].XIC[5].icell.Ien VPWR 0.18883f
C734 XThC.Tn[1] XA.XIR[0].XIC[1].icell.Ien 0.04659f
C735 XA.XIR[14].XIC[10].icell.Ien Vbias 0.19161f
C736 XThR.Tn[13] XA.XIR[13].XIC[12].icell.Ien 0.14211f
C737 XThC.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.02602f
C738 XThC.XTB7.A XThC.XTBN.Y 0.59539f
C739 XA.XIR[13].XIC[7].icell.Ien VPWR 0.18829f
C740 XA.XIR[2].XIC_15.icell.Ien Iout 0.0694f
C741 XThR.Tn[8] XA.XIR[9].XIC[3].icell.PDM 0.04035f
C742 XThR.Tn[12] XA.XIR[13].XIC[8].icell.PDM 0.04035f
C743 XA.XIR[12].XIC[11].icell.Ien Iout 0.06801f
C744 XThR.XTB6.A XThR.XTBN.A 0.0512f
C745 XA.XIR[11].XIC_dummy_right.icell.PDM VPWR 0.08209f
C746 XThR.XTB7.Y a_n997_1579# 0.013f
C747 XA.XIR[11].XIC_dummy_right.icell.PUM VPWR 0.01691f
C748 XA.XIR[3].XIC_15.icell.Ien XA.XIR[4].XIC_15.icell.PDM 0.02104f
C749 XThC.Tn[4] XA.XIR[12].XIC[4].icell.PDM 0.02601f
C750 XThC.Tn[9] XA.XIR[15].XIC[9].icell.PDM 0.02601f
C751 a_n997_1803# VPWR 0.01991f
C752 XThC.Tn[10] XA.XIR[0].XIC[10].icell.PDM 0.02792f
C753 XThC.Tn[10] XA.XIR[15].XIC[10].icell.Ien 0.04292f
C754 XThR.Tn[5] XA.XIR[6].XIC[0].icell.PDM 0.0404f
C755 XA.XIR[9].XIC_dummy_left.icell.Ien XThR.Tn[9] 0.01244f
C756 XA.XIR[4].XIC[1].icell.Ien Vbias 0.19161f
C757 XThC.XTB7.A a_4861_9615# 0.02294f
C758 XThC.Tn[3] XA.XIR[10].XIC[3].icell.PDM 0.02601f
C759 XThC.Tn[3] XThC.Tn[4] 0.45992f
C760 XThR.Tn[12] XA.XIR[13].XIC[13].icell.PDM 0.0404f
C761 XA.XIR[2].XIC_dummy_right.icell.Iout Iout 0.01732f
C762 XA.XIR[5].XIC[5].icell.Ien Iout 0.06801f
C763 XThC.Tn[8] XA.XIR[13].XIC[8].icell.PDM 0.02601f
C764 XA.XIR[2].XIC[14].icell.Ien VPWR 0.18835f
C765 XA.XIR[6].XIC[11].icell.Ien XA.XIR[7].XIC[11].icell.PDM 0.02104f
C766 XThC.XTB1.Y Vbias 0.01576f
C767 XThC.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.02601f
C768 XThC.XTB5.A XThC.XTB5.Y 0.0538f
C769 XA.XIR[15].XIC[3].icell.Ien Vbias 0.15966f
C770 XA.XIR[9].XIC[5].icell.PDM XA.XIR[9].XIC[5].icell.Ien 0.04854f
C771 XThR.Tn[8] XA.XIR[8].XIC[11].icell.Ien 0.14211f
C772 XA.XIR[7].XIC[3].icell.PDM XA.XIR[7].XIC[3].icell.Ien 0.04854f
C773 XA.XIR[14].XIC[0].icell.Ien VPWR 0.18883f
C774 XA.XIR[4].XIC[6].icell.Ien Vbias 0.19161f
C775 XA.XIR[4].XIC[4].icell.PDM XA.XIR[4].XIC[4].icell.Ien 0.04854f
C776 XThR.Tn[8] data[4] 0.01643f
C777 XThR.Tn[5] Iout 1.12761f
C778 XThR.Tn[13] VPWR 9.0331f
C779 data[1] data[2] 0.01393f
C780 XThC.XTBN.Y a_5949_9615# 0.07703f
C781 XThC.Tn[11] XThR.Tn[7] 0.40738f
C782 XThC.Tn[2] XA.XIR[5].XIC[2].icell.Ien 0.04604f
C783 XA.XIR[14].XIC[6].icell.Ien XA.XIR[15].XIC[6].icell.PDM 0.02104f
C784 XThC.XTB7.B XThC.Tn[9] 0.05542f
C785 XThR.XTBN.A data[7] 0.07741f
C786 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.PDM 0.02104f
C787 XA.XIR[13].XIC[13].icell.Ien XA.XIR[14].XIC[13].icell.PDM 0.02104f
C788 XThC.XTB7.Y XThC.Tn[13] 0.10846f
C789 XThR.Tn[5] XA.XIR[5].XIC[10].icell.Ien 0.14211f
C790 XA.XIR[9].XIC[13].icell.PDM Vbias 0.03928f
C791 XA.XIR[8].XIC[2].icell.PDM XA.XIR[8].XIC[2].icell.Ien 0.04854f
C792 XThC.Tn[1] XA.XIR[7].XIC[1].icell.PDM 0.02601f
C793 XA.XIR[7].XIC[0].icell.Ien Vbias 0.19149f
C794 XA.XIR[0].XIC[5].icell.PDM Vbias 0.03945f
C795 XA.XIR[5].XIC[4].icell.Ien VPWR 0.18829f
C796 XThC.Tn[1] XA.XIR[10].XIC[1].icell.Ien 0.04604f
C797 XThR.Tn[13] XA.XIR[13].XIC[10].icell.Ien 0.14211f
C798 XA.XIR[13].XIC[9].icell.Ien XA.XIR[14].XIC[9].icell.PDM 0.02104f
C799 XThC.Tn[12] XA.XIR[9].XIC[12].icell.PDM 0.02601f
C800 XA.XIR[9].XIC[9].icell.Ien Vbias 0.19161f
C801 XA.XIR[2].XIC[1].icell.Ien XA.XIR[3].XIC[1].icell.PDM 0.02104f
C802 XThR.Tn[3] a_n1049_6699# 0.27008f
C803 XThR.Tn[1] XA.XIR[1].XIC_15.icell.Ien 0.13564f
C804 XA.XIR[0].XIC[2].icell.Ien Vbias 0.19213f
C805 XA.XIR[8].XIC[9].icell.Ien XA.XIR[9].XIC[9].icell.PDM 0.02104f
C806 XA.XIR[11].XIC[14].icell.PDM Vbias 0.03928f
C807 XThC.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.02601f
C808 XA.XIR[14].XIC[10].icell.Ien XA.XIR[15].XIC[10].icell.PDM 0.02104f
C809 XA.XIR[3].XIC[8].icell.Ien XA.XIR[4].XIC[8].icell.PDM 0.02104f
C810 XA.XIR[9].XIC[14].icell.PDM VPWR 0.0118f
C811 XThR.XTB6.A XThR.XTB6.Y 0.10153f
C812 XA.XIR[9].XIC[13].icell.Ien XA.XIR[10].XIC[13].icell.PDM 0.02104f
C813 XA.XIR[0].XIC[6].icell.PDM VPWR 0.01138f
C814 XA.XIR[14].XIC_15.icell.PDM Vbias 0.03927f
C815 XA.XIR[3].XIC[10].icell.PDM XA.XIR[3].XIC[10].icell.Ien 0.04854f
C816 XThC.Tn[10] XThR.Tn[3] 0.40738f
C817 XA.XIR[14].XIC_15.icell.Ien Vbias 0.19195f
C818 XA.XIR[7].XIC[5].icell.Ien Vbias 0.19161f
C819 XA.XIR[1].XIC_dummy_left.icell.Iout VPWR 0.11048f
C820 XThC.Tn[7] VPWR 3.9785f
C821 XA.XIR[15].XIC[1].icell.PDM XA.XIR[15].XIC[1].icell.Ien 0.04854f
C822 XThR.Tn[10] XA.XIR[11].XIC[2].icell.PDM 0.04035f
C823 XThR.Tn[4] XA.XIR[5].XIC[13].icell.PDM 0.0404f
C824 XThR.Tn[14] XA.XIR[15].XIC[3].icell.PDM 0.04035f
C825 XThC.Tn[13] XThR.Tn[0] 0.40764f
C826 XA.XIR[9].XIC[1].icell.Ien XA.XIR[10].XIC[1].icell.PDM 0.02104f
C827 XA.XIR[10].XIC[11].icell.Ien XA.XIR[11].XIC[11].icell.PDM 0.02104f
C828 XA.XIR[14].XIC_dummy_right.icell.PDM VPWR 0.08209f
C829 XThC.Tn[4] XA.XIR[15].XIC[4].icell.PDM 0.02601f
C830 XA.XIR[14].XIC_dummy_right.icell.PUM VPWR 0.01691f
C831 XA.XIR[6].XIC[4].icell.Ien XA.XIR[7].XIC[4].icell.PDM 0.02104f
C832 XThC.Tn[6] XA.XIR[10].XIC[6].icell.Ien 0.04604f
C833 XA.XIR[15].XIC[13].icell.Ien Iout 0.07192f
C834 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.Iout 0.06446f
C835 XThC.Tn[5] XA.XIR[0].XIC[5].icell.PDM 0.02803f
C836 XA.XIR[2].XIC[0].icell.PDM XA.XIR[2].XIC[0].icell.Ien 0.04854f
C837 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Ien 0.01263f
C838 XA.XIR[8].XIC_dummy_left.icell.Ien VPWR 0.38999f
C839 a_2979_9615# Vbias 0.01381f
C840 XThC.Tn[13] XA.XIR[5].XIC[13].icell.PDM 0.02601f
C841 XThC.XTBN.A XThC.XTB7.Y 1.11562f
C842 XThR.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.04035f
C843 XA.XIR[5].XIC[3].icell.PDM Vbias 0.03928f
C844 XThR.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.14211f
C845 XThR.XTB5.A data[5] 0.11096f
C846 XThC.Tn[9] XA.XIR[4].XIC[9].icell.Ien 0.04604f
C847 XA.XIR[1].XIC_15.icell.PDM XA.XIR[1].XIC_15.icell.Ien 0.04854f
C848 XThC.Tn[3] XA.XIR[13].XIC[3].icell.PDM 0.02601f
C849 XA.XIR[4].XIC[11].icell.Ien XA.XIR[5].XIC[11].icell.PDM 0.02104f
C850 XThR.XTBN.A XThR.Tn[12] 0.22096f
C851 XA.XIR[12].XIC[2].icell.PDM Vbias 0.03928f
C852 XA.XIR[13].XIC[2].icell.Ien XA.XIR[14].XIC[2].icell.PDM 0.02104f
C853 XThC.Tn[5] XA.XIR[7].XIC[5].icell.Ien 0.04604f
C854 a_3773_9615# VPWR 0.70508f
C855 XA.XIR[11].XIC[8].icell.PDM Vbias 0.03928f
C856 XA.XIR[13].XIC[3].icell.PDM XA.XIR[13].XIC[3].icell.Ien 0.04854f
C857 XThC.Tn[12] XThR.Tn[2] 0.40741f
C858 XThR.XTB2.Y a_n997_3755# 0.06476f
C859 XThR.Tn[2] XA.XIR[3].XIC[7].icell.PDM 0.04035f
C860 XA.XIR[11].XIC_dummy_left.icell.Iout Iout 0.03553f
C861 XA.XIR[5].XIC[4].icell.PDM VPWR 0.01171f
C862 XA.XIR[12].XIC[4].icell.Ien XA.XIR[13].XIC[4].icell.PDM 0.02104f
C863 XA.XIR[8].XIC[2].icell.Ien XA.XIR[9].XIC[2].icell.PDM 0.02104f
C864 XA.XIR[5].XIC[10].icell.Ien Iout 0.06801f
C865 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.Iout 0.06446f
C866 XThC.XTB4.Y a_5155_9615# 0.01546f
C867 XThR.XTBN.Y a_n1049_8581# 0.0607f
C868 XThR.Tn[13] XA.XIR[13].XIC_15.icell.Ien 0.13564f
C869 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.PDM 0.02104f
C870 XThR.Tn[6] XA.XIR[7].XIC[14].icell.PDM 0.04056f
C871 XA.XIR[3].XIC[2].icell.Ien Vbias 0.19161f
C872 XA.XIR[6].XIC_dummy_left.icell.Iout VPWR 0.11008f
C873 XA.XIR[15].XIC[8].icell.Ien Vbias 0.15966f
C874 XA.XIR[3].XIC[3].icell.PDM XA.XIR[3].XIC[3].icell.Ien 0.04854f
C875 XA.XIR[12].XIC[3].icell.PDM VPWR 0.01171f
C876 XA.XIR[0].XIC[1].icell.Ien XA.XIR[1].XIC[1].icell.PDM 0.02104f
C877 XThC.Tn[7] XA.XIR[9].XIC[7].icell.PDM 0.02601f
C878 XA.XIR[11].XIC[9].icell.PDM VPWR 0.01171f
C879 XA.XIR[11].XIC[8].icell.PDM XA.XIR[11].XIC[8].icell.Ien 0.04854f
C880 XA.XIR[8].XIC[0].icell.PDM Vbias 0.03915f
C881 XA.XIR[4].XIC[11].icell.Ien Vbias 0.19161f
C882 XThC.Tn[1] XA.XIR[13].XIC[1].icell.Ien 0.04604f
C883 XA.XIR[12].XIC[5].icell.Ien Iout 0.06801f
C884 XA.XIR[11].XIC[13].icell.PDM Vbias 0.03928f
C885 XA.XIR[2].XIC[4].icell.PDM Vbias 0.03928f
C886 XThC.Tn[8] XThR.Tn[6] 0.40738f
C887 XThC.Tn[7] XA.XIR[9].XIC[7].icell.Ien 0.04604f
C888 XA.XIR[8].XIC[5].icell.Ien Vbias 0.19161f
C889 XThR.Tn[9] XA.XIR[10].XIC[1].icell.PDM 0.04035f
C890 XThC.Tn[14] XA.XIR[0].XIC[14].icell.Ien 0.04662f
C891 XA.XIR[15].XIC[11].icell.Ien Iout 0.07192f
C892 XThR.Tn[5] XA.XIR[5].XIC_15.icell.Ien 0.13564f
C893 XA.XIR[14].XIC[14].icell.PDM Vbias 0.03928f
C894 XThR.XTB3.Y a_n997_2891# 0.07285f
C895 XThC.Tn[10] XThR.Tn[11] 0.40738f
C896 XA.XIR[5].XIC[9].icell.Ien VPWR 0.18829f
C897 XThC.XTBN.Y a_8739_9569# 0.22804f
C898 XThC.Tn[0] XThR.Tn[7] 0.40736f
C899 XA.XIR[9].XIC[14].icell.Ien Vbias 0.19161f
C900 XThC.XTB3.Y XThC.XTB7.Y 0.03772f
C901 XThC.XTB4.Y XThC.XTB6.Y 0.04273f
C902 XA.XIR[8].XIC[1].icell.PDM VPWR 0.01171f
C903 XThC.Tn[2] XA.XIR[12].XIC[2].icell.Ien 0.04604f
C904 XThR.Tn[4] XA.XIR[4].XIC[0].icell.Ien 0.1423f
C905 a_n1049_5317# XThR.Tn[6] 0.26047f
C906 XA.XIR[10].XIC[0].icell.Ien XThR.Tn[10] 0.14211f
C907 XA.XIR[2].XIC[5].icell.PDM VPWR 0.01171f
C908 XA.XIR[0].XIC[7].icell.Ien Vbias 0.19213f
C909 XThR.Tn[3] XA.XIR[3].XIC[0].icell.Ien 0.14251f
C910 XA.XIR[12].XIC[0].icell.Ien XA.XIR[13].XIC[0].icell.PDM 0.02104f
C911 XA.XIR[0].XIC_dummy_left.icell.Ien XA.XIR[0].XIC_dummy_left.icell.Iout 0.06446f
C912 XThC.XTB7.B XThC.Tn[7] 0.07854f
C913 XThC.XTB5.Y XThC.Tn[11] 0.02112f
C914 XA.XIR[12].XIC[4].icell.Ien VPWR 0.18829f
C915 XA.XIR[13].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.Iout 0.06446f
C916 XA.XIR[1].XIC[8].icell.PDM XA.XIR[1].XIC[8].icell.Ien 0.04854f
C917 XA.XIR[4].XIC[4].icell.Ien XA.XIR[5].XIC[4].icell.PDM 0.02104f
C918 a_8739_9569# XThC.Tn[10] 0.21014f
C919 XThR.XTB7.Y XThR.Tn[8] 0.07806f
C920 a_n997_3979# VPWR 0.01662f
C921 XThR.Tn[11] XA.XIR[12].XIC[5].icell.PDM 0.04035f
C922 XA.XIR[7].XIC[10].icell.Ien Vbias 0.19161f
C923 XThC.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.04606f
C924 XThC.Tn[13] XThR.Tn[1] 0.40745f
C925 XA.XIR[9].XIC_15.icell.PUM VPWR 0.01655f
C926 XThR.Tn[8] XA.XIR[8].XIC_dummy_left.icell.Iout 0.03962f
C927 XA.XIR[8].XIC_dummy_left.icell.PUM VPWR 0.01604f
C928 XThR.Tn[4] XA.XIR[4].XIC[5].icell.Ien 0.14211f
C929 XThC.Tn[6] XA.XIR[13].XIC[6].icell.Ien 0.04604f
C930 XA.XIR[7].XIC_dummy_left.icell.PDM XA.XIR[7].XIC_dummy_left.icell.Ien 0.04854f
C931 XThR.XTB6.Y XThR.Tn[12] 0.02431f
C932 XA.XIR[2].XIC[10].icell.PDM XA.XIR[2].XIC[10].icell.Ien 0.04854f
C933 XThC.Tn[13] XThR.Tn[12] 0.40739f
C934 XThR.Tn[12] XA.XIR[13].XIC[11].icell.PDM 0.04035f
C935 XA.XIR[8].XIC[0].icell.Ien Vbias 0.19149f
C936 XThR.Tn[0] XA.XIR[1].XIC[3].icell.PDM 0.04035f
C937 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.PDM 0.02104f
C938 XThC.XTB6.A XThC.XTBN.A 0.0513f
C939 XA.XIR[9].XIC[1].icell.Ien Iout 0.06801f
C940 XThC.Tn[10] XA.XIR[1].XIC[10].icell.PDM 0.02602f
C941 XThC.XTBN.Y XThC.Tn[11] 0.40412f
C942 XThC.Tn[8] XThR.Tn[4] 0.40738f
C943 XThC.Tn[5] XA.XIR[8].XIC[5].icell.Ien 0.04604f
C944 XThR.Tn[1] XA.XIR[2].XIC[2].icell.PDM 0.04035f
C945 XA.XIR[5].XIC_dummy_left.icell.Ien VPWR 0.38939f
C946 XA.XIR[4].XIC[3].icell.Ien Iout 0.06801f
C947 XThC.Tn[10] XA.XIR[4].XIC[10].icell.PDM 0.02601f
C948 XA.XIR[7].XIC[4].icell.PDM Vbias 0.03928f
C949 XThR.Tn[7] XA.XIR[8].XIC[7].icell.PDM 0.04035f
C950 XA.XIR[6].XIC[11].icell.PDM Vbias 0.03928f
C951 XA.XIR[15].XIC[2].icell.PDM Vbias 0.03928f
C952 XThC.Tn[2] XThR.Tn[0] 0.40765f
C953 XThC.Tn[12] XThR.Tn[10] 0.40738f
C954 XThC.Tn[4] XThR.Tn[5] 0.40738f
C955 XThR.Tn[12] XA.XIR[12].XIC[3].icell.Ien 0.14211f
C956 XA.XIR[14].XIC[8].icell.PDM Vbias 0.03928f
C957 XThR.Tn[3] XA.XIR[3].XIC[8].icell.Ien 0.14211f
C958 XA.XIR[5].XIC[13].icell.PDM XA.XIR[5].XIC[13].icell.Ien 0.04854f
C959 XThC.Tn[10] XThC.Tn[11] 0.07237f
C960 XThC.Tn[9] XA.XIR[8].XIC[9].icell.PDM 0.02601f
C961 XA.XIR[9].XIC[6].icell.Ien Iout 0.06801f
C962 XA.XIR[14].XIC_dummy_left.icell.Iout Iout 0.03553f
C963 XThR.Tn[7] VPWR 8.3986f
C964 a_n997_2891# VPWR 0.01347f
C965 XA.XIR[9].XIC[0].icell.PDM Vbias 0.03915f
C966 XThR.Tn[3] XA.XIR[4].XIC[8].icell.PDM 0.04035f
C967 XThC.XTB1.Y XThC.XTB7.Y 0.05222f
C968 XThC.Tn[8] XA.XIR[5].XIC[8].icell.Ien 0.04604f
C969 XThC.XTB2.Y XThC.XTB6.Y 0.04959f
C970 XThC.Tn[14] XA.XIR[3].XIC[14].icell.Ien 0.04604f
C971 XA.XIR[7].XIC[5].icell.PDM VPWR 0.01171f
C972 XThR.Tn[2] XA.XIR[2].XIC[3].icell.Ien 0.14211f
C973 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.Iout 0.06446f
C974 XA.XIR[15].XIC[3].icell.PDM VPWR 0.01512f
C975 XA.XIR[4].XIC[2].icell.Ien VPWR 0.18829f
C976 XA.XIR[6].XIC[12].icell.PDM VPWR 0.01171f
C977 XThR.XTB6.Y a_n1049_5317# 0.01199f
C978 XA.XIR[3].XIC_dummy_right.icell.Iout XA.XIR[4].XIC_dummy_right.icell.Iout 0.04047f
C979 XA.XIR[11].XIC[12].icell.PDM Vbias 0.03928f
C980 XThC.Tn[0] XA.XIR[9].XIC[0].icell.Ien 0.04604f
C981 XA.XIR[12].XIC[13].icell.PDM XA.XIR[12].XIC[13].icell.Ien 0.04854f
C982 XA.XIR[14].XIC[9].icell.PDM VPWR 0.01171f
C983 XA.XIR[5].XIC_15.icell.Ien Iout 0.0694f
C984 XA.XIR[7].XIC[2].icell.Ien Iout 0.06801f
C985 XThC.Tn[1] XA.XIR[6].XIC[1].icell.Ien 0.04604f
C986 XA.XIR[3].XIC[7].icell.Ien Vbias 0.19161f
C987 XA.XIR[1].XIC[5].icell.PDM Vbias 0.03928f
C988 XA.XIR[12].XIC[9].icell.PDM XA.XIR[12].XIC[9].icell.Ien 0.04854f
C989 XA.XIR[14].XIC[13].icell.PDM Vbias 0.03928f
C990 XA.XIR[9].XIC[1].icell.PDM VPWR 0.01171f
C991 XThC.Tn[1] XA.XIR[12].XIC[1].icell.PDM 0.02601f
C992 XThC.Tn[1] XThR.Tn[2] 0.40741f
C993 XA.XIR[4].XIC[5].icell.PDM Vbias 0.03928f
C994 XA.XIR[9].XIC[5].icell.Ien VPWR 0.18829f
C995 XA.XIR[1].XIC[2].icell.Ien Vbias 0.19173f
C996 XA.XIR[8].XIC_15.icell.PDM Vbias 0.03927f
C997 XA.XIR[3].XIC[13].icell.PDM Vbias 0.03928f
C998 XThC.Tn[10] XThR.Tn[14] 0.40738f
C999 XThR.XTBN.Y a_n1049_7787# 0.08456f
C1000 XThC.Tn[12] XA.XIR[3].XIC[12].icell.PDM 0.02601f
C1001 XThC.XTB2.Y XThC.XTB4.Y 0.04006f
C1002 XThC.XTB6.A XThC.XTB3.Y 0.03869f
C1003 XA.XIR[2].XIC[3].icell.PDM XA.XIR[2].XIC[3].icell.Ien 0.04854f
C1004 XThR.Tn[4] XA.XIR[5].XIC[0].icell.PDM 0.0404f
C1005 XA.XIR[8].XIC[10].icell.Ien Vbias 0.19161f
C1006 XThR.XTB2.Y XThR.XTB7.Y 0.0437f
C1007 XA.XIR[1].XIC[6].icell.PDM VPWR 0.01171f
C1008 XThR.Tn[9] Iout 1.12762f
C1009 XA.XIR[5].XIC_dummy_right.icell.Iout Iout 0.01732f
C1010 XThC.Tn[0] XA.XIR[10].XIC[0].icell.PDM 0.02601f
C1011 XA.XIR[5].XIC_dummy_left.icell.Iout XA.XIR[6].XIC_dummy_left.icell.Iout 0.03665f
C1012 XA.XIR[11].XIC[1].icell.Ien XThR.Tn[11] 0.14211f
C1013 XA.XIR[9].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1014 a_n1049_6405# XThR.Tn[4] 0.26564f
C1015 a_5155_9615# XThC.Tn[4] 0.27224f
C1016 XA.XIR[4].XIC[6].icell.PDM VPWR 0.01171f
C1017 XA.XIR[5].XIC[14].icell.Ien VPWR 0.18835f
C1018 XThR.Tn[13] XA.XIR[14].XIC[2].icell.PDM 0.04035f
C1019 XA.XIR[3].XIC[14].icell.PDM VPWR 0.0118f
C1020 XA.XIR[8].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1021 XA.XIR[13].XIC[11].icell.Ien XA.XIR[14].XIC[11].icell.PDM 0.02104f
C1022 XThC.XTBN.A XThC.Tn[8] 0.13691f
C1023 XThC.Tn[6] XThR.Tn[6] 0.40738f
C1024 XA.XIR[12].XIC_15.icell.PUM VPWR 0.01655f
C1025 XThR.Tn[8] XA.XIR[9].XIC[5].icell.PDM 0.04035f
C1026 XA.XIR[0].XIC[12].icell.Ien Vbias 0.19213f
C1027 XThR.Tn[12] XA.XIR[13].XIC[10].icell.PDM 0.04035f
C1028 XA.XIR[15].XIC[0].icell.Ien Iout 0.07185f
C1029 XA.XIR[5].XIC[6].icell.PDM XA.XIR[5].XIC[6].icell.Ien 0.04854f
C1030 XA.XIR[12].XIC[9].icell.Ien VPWR 0.18829f
C1031 XA.XIR[5].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1032 XA.XIR[7].XIC_15.icell.Ien Vbias 0.19195f
C1033 XThC.Tn[5] XA.XIR[1].XIC[5].icell.PDM 0.02602f
C1034 XA.XIR[5].XIC[0].icell.Ien Vbias 0.19149f
C1035 XA.XIR[9].XIC[0].icell.Ien VPWR 0.18829f
C1036 XThR.Tn[12] XA.XIR[13].XIC_dummy_left.icell.Iout 0.01828f
C1037 XThR.Tn[5] XA.XIR[6].XIC[2].icell.PDM 0.04035f
C1038 XThC.Tn[5] XA.XIR[4].XIC[5].icell.PDM 0.02601f
C1039 XThC.Tn[4] Iout 0.22518f
C1040 XThR.Tn[4] XA.XIR[4].XIC[10].icell.Ien 0.14211f
C1041 XThC.Tn[9] XA.XIR[9].XIC[9].icell.PDM 0.02601f
C1042 XThC.Tn[14] Vbias 0.8291f
C1043 XThR.Tn[0] XA.XIR[0].XIC[2].icell.Ien 0.14211f
C1044 XThC.XTB7.A a_5949_9615# 0.01824f
C1045 XThC.Tn[11] XA.XIR[7].XIC[11].icell.Ien 0.04604f
C1046 XA.XIR[15].XIC[5].icell.Ien Iout 0.07192f
C1047 XThC.Tn[12] XThR.Tn[13] 0.40738f
C1048 XThC.Tn[2] XThR.Tn[1] 0.40744f
C1049 XThR.Tn[6] XA.XIR[7].XIC[1].icell.PDM 0.04035f
C1050 XA.XIR[12].XIC[2].icell.PDM XA.XIR[12].XIC[2].icell.Ien 0.04854f
C1051 XA.XIR[6].XIC[2].icell.Ien Vbias 0.19161f
C1052 XA.XIR[4].XIC[8].icell.Ien Iout 0.06801f
C1053 XA.XIR[7].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1054 XThR.Tn[7] XA.XIR[7].XIC[3].icell.Ien 0.14211f
C1055 XThC.Tn[4] XA.XIR[8].XIC[4].icell.PDM 0.02601f
C1056 XThC.XTB2.Y a_7875_9569# 0.06476f
C1057 XThC.Tn[2] XThR.Tn[12] 0.40738f
C1058 XThC.XTB1.Y XThC.XTB6.A 0.01609f
C1059 XThC.XTB5.A XThC.XTB7.A 0.07824f
C1060 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.Iout 0.06446f
C1061 XThC.Tn[11] XThR.Tn[8] 0.40738f
C1062 a_n997_1579# VPWR 0.02417f
C1063 XA.XIR[8].XIC[2].icell.Ien Iout 0.06801f
C1064 XThC.Tn[10] XA.XIR[10].XIC[10].icell.Ien 0.04604f
C1065 XA.XIR[11].XIC[11].icell.PDM Vbias 0.03928f
C1066 XA.XIR[5].XIC_15.icell.Ien XA.XIR[6].XIC_15.icell.PDM 0.02104f
C1067 XThR.Tn[12] XA.XIR[12].XIC[8].icell.Ien 0.14211f
C1068 XA.XIR[10].XIC[0].icell.PDM VPWR 0.01171f
C1069 XThC.XTBN.Y XThC.Tn[0] 0.45269f
C1070 XA.XIR[7].XIC_dummy_left.icell.Iout XA.XIR[8].XIC_dummy_left.icell.Iout 0.03665f
C1071 XThC.Tn[2] XA.XIR[15].XIC[2].icell.Ien 0.04292f
C1072 XThR.Tn[3] XA.XIR[3].XIC[13].icell.Ien 0.14211f
C1073 XThC.Tn[6] XThR.Tn[4] 0.40738f
C1074 XA.XIR[14].XIC[12].icell.PDM Vbias 0.03928f
C1075 XA.XIR[9].XIC[11].icell.Ien Iout 0.06801f
C1076 XA.XIR[14].XIC[8].icell.PDM XA.XIR[14].XIC[8].icell.Ien 0.04854f
C1077 XA.XIR[9].XIC_15.icell.PDM Vbias 0.03927f
C1078 XA.XIR[1].XIC[1].icell.PDM XA.XIR[1].XIC[1].icell.Ien 0.04854f
C1079 XThC.Tn[13] XA.XIR[9].XIC[13].icell.Ien 0.04604f
C1080 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[5].XIC_dummy_left.icell.Iout 0.06446f
C1081 XThC.XTB2.Y data[1] 0.017f
C1082 XA.XIR[0].XIC[7].icell.PDM Vbias 0.03945f
C1083 XA.XIR[15].XIC[4].icell.Ien VPWR 0.31713f
C1084 XThC.Tn[1] XThR.Tn[10] 0.40738f
C1085 XA.XIR[0].XIC[4].icell.Ien Iout 0.0675f
C1086 XThC.Tn[6] XA.XIR[11].XIC[6].icell.PDM 0.02601f
C1087 XThC.Tn[3] XA.XIR[11].XIC[3].icell.Ien 0.04604f
C1088 XThR.Tn[2] XA.XIR[2].XIC[8].icell.Ien 0.14211f
C1089 XThC.Tn[1] XA.XIR[15].XIC[1].icell.PDM 0.02601f
C1090 XA.XIR[10].XIC[3].icell.Ien Vbias 0.19161f
C1091 XA.XIR[4].XIC[7].icell.Ien VPWR 0.18829f
C1092 XThR.Tn[9] XA.XIR[9].XIC[1].icell.Ien 0.14211f
C1093 XThC.Tn[2] XA.XIR[0].XIC[2].icell.PDM 0.02803f
C1094 XThR.XTB7.Y a_n997_715# 0.06874f
C1095 XThC.Tn[14] XA.XIR[1].XIC[14].icell.Ien 0.04606f
C1096 XA.XIR[7].XIC[7].icell.Ien Iout 0.06801f
C1097 XThC.Tn[7] XA.XIR[3].XIC[7].icell.PDM 0.02601f
C1098 XThC.Tn[10] XA.XIR[5].XIC[10].icell.PDM 0.02601f
C1099 XThC.Tn[8] XA.XIR[12].XIC[8].icell.Ien 0.04604f
C1100 XA.XIR[3].XIC[12].icell.Ien Vbias 0.19161f
C1101 XA.XIR[3].XIC_dummy_left.icell.Iout XA.XIR[4].XIC_dummy_left.icell.Iout 0.03665f
C1102 XA.XIR[9].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1103 XA.XIR[7].XIC[1].icell.Ien VPWR 0.18829f
C1104 XA.XIR[13].XIC[0].icell.Ien XThR.Tn[13] 0.14211f
C1105 XA.XIR[0].XIC[8].icell.PDM VPWR 0.01451f
C1106 XThC.XTBN.A data[3] 0.07741f
C1107 XThC.XTB5.Y VPWR 1.01219f
C1108 XA.XIR[2].XIC[5].icell.Ien Vbias 0.19161f
C1109 XA.XIR[9].XIC[10].icell.Ien VPWR 0.18829f
C1110 XThC.Tn[0] XA.XIR[13].XIC[0].icell.PDM 0.02601f
C1111 XThC.XTB7.A data[0] 0.86893f
C1112 XA.XIR[1].XIC[7].icell.Ien Vbias 0.19173f
C1113 XA.XIR[12].XIC[14].icell.Ien VPWR 0.18835f
C1114 XA.XIR[0].XIC[9].icell.PDM XA.XIR[0].XIC[9].icell.Ien 0.04854f
C1115 XThR.Tn[9] XA.XIR[9].XIC[6].icell.Ien 0.14211f
C1116 XA.XIR[0].XIC[3].icell.Ien VPWR 0.18776f
C1117 XThR.Tn[10] XA.XIR[11].XIC[4].icell.PDM 0.04035f
C1118 XA.XIR[8].XIC_15.icell.Ien Vbias 0.19195f
C1119 XThR.Tn[14] XA.XIR[15].XIC[5].icell.PDM 0.04035f
C1120 XA.XIR[7].XIC[6].icell.Ien VPWR 0.18829f
C1121 XThC.XTBN.Y VPWR 4.12335f
C1122 XThC.Tn[11] XA.XIR[8].XIC[11].icell.Ien 0.04604f
C1123 XThC.XTB6.Y a_6243_9615# 0.01199f
C1124 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.PDM 0.02104f
C1125 a_n1049_6699# VPWR 0.72162f
C1126 XThR.XTB7.A XThR.XTBN.A 0.19736f
C1127 XA.XIR[5].XIC[8].icell.Ien XA.XIR[6].XIC[8].icell.PDM 0.02104f
C1128 XA.XIR[8].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1129 XThC.Tn[4] XA.XIR[9].XIC[4].icell.PDM 0.02601f
C1130 XThR.XTB7.A XThR.Tn[6] 0.1056f
C1131 XA.XIR[5].XIC[5].icell.PDM Vbias 0.03928f
C1132 XThC.XTB1.Y XThC.Tn[8] 0.29214f
C1133 XThR.Tn[11] XA.XIR[11].XIC[2].icell.Ien 0.14211f
C1134 XThC.Tn[10] VPWR 4.54895f
C1135 XA.XIR[12].XIC[4].icell.PDM Vbias 0.03928f
C1136 XThC.Tn[14] XA.XIR[6].XIC[14].icell.Ien 0.04604f
C1137 XThC.Tn[5] XA.XIR[2].XIC[5].icell.Ien 0.04605f
C1138 XThR.Tn[4] XA.XIR[4].XIC_15.icell.Ien 0.13564f
C1139 a_4861_9615# VPWR 0.70519f
C1140 XThC.Tn[13] XA.XIR[11].XIC[13].icell.Ien 0.04604f
C1141 XA.XIR[11].XIC[10].icell.PDM Vbias 0.03928f
C1142 XA.XIR[3].XIC[4].icell.Ien Iout 0.06801f
C1143 XA.XIR[10].XIC[13].icell.Ien Iout 0.06801f
C1144 XThR.Tn[0] XA.XIR[0].XIC[7].icell.Ien 0.14211f
C1145 XA.XIR[10].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1146 XThR.Tn[10] XA.XIR[10].XIC[6].icell.Ien 0.14211f
C1147 XThR.Tn[2] XA.XIR[3].XIC[9].icell.PDM 0.04035f
C1148 XA.XIR[5].XIC[6].icell.PDM VPWR 0.01171f
C1149 XThC.Tn[10] XA.XIR[13].XIC[10].icell.Ien 0.04604f
C1150 XA.XIR[14].XIC[11].icell.PDM Vbias 0.03928f
C1151 XA.XIR[13].XIC[0].icell.PDM VPWR 0.01171f
C1152 XThR.Tn[7] XA.XIR[7].XIC[8].icell.Ien 0.14211f
C1153 XA.XIR[4].XIC[13].icell.Ien Iout 0.06801f
C1154 XA.XIR[6].XIC[7].icell.Ien Vbias 0.19161f
C1155 XThC.XTB5.A data[0] 0.14415f
C1156 XThC.XTB5.Y a_9827_9569# 0.06458f
C1157 XA.XIR[12].XIC[5].icell.PDM VPWR 0.01171f
C1158 XA.XIR[11].XIC[7].icell.Ien XA.XIR[12].XIC[7].icell.PDM 0.02104f
C1159 XA.XIR[12].XIC[12].icell.Ien VPWR 0.18829f
C1160 XThC.Tn[3] Vbias 0.84088f
C1161 XA.XIR[8].XIC[7].icell.Ien Iout 0.06801f
C1162 XA.XIR[8].XIC[2].icell.PDM Vbias 0.03928f
C1163 XA.XIR[3].XIC[0].icell.PDM Vbias 0.03915f
C1164 XThC.Tn[6] XA.XIR[14].XIC[6].icell.PDM 0.02601f
C1165 XThC.Tn[3] XA.XIR[14].XIC[3].icell.Ien 0.04604f
C1166 XThC.Tn[1] XThR.Tn[13] 0.40738f
C1167 XA.XIR[0].XIC[2].icell.PDM XA.XIR[0].XIC[2].icell.Ien 0.04854f
C1168 XA.XIR[8].XIC[1].icell.Ien VPWR 0.18829f
C1169 XA.XIR[2].XIC[6].icell.PDM Vbias 0.03928f
C1170 XA.XIR[13].XIC[3].icell.Ien Vbias 0.19161f
C1171 XA.XIR[3].XIC[3].icell.Ien VPWR 0.18829f
C1172 XThR.Tn[9] XA.XIR[10].XIC[3].icell.PDM 0.04035f
C1173 XA.XIR[15].XIC_15.icell.PUM VPWR 0.01655f
C1174 XThC.Tn[4] XThR.Tn[9] 0.40738f
C1175 XThC.Tn[5] XA.XIR[5].XIC[5].icell.PDM 0.02601f
C1176 XThC.Tn[0] XThR.Tn[8] 0.40736f
C1177 XThC.Tn[0] XA.XIR[3].XIC[0].icell.Ien 0.04604f
C1178 XThR.XTB7.A XThR.Tn[4] 0.02736f
C1179 XA.XIR[15].XIC[9].icell.Ien VPWR 0.31713f
C1180 XA.XIR[11].XIC[6].icell.Ien Vbias 0.19161f
C1181 XA.XIR[0].XIC[9].icell.Ien Iout 0.0675f
C1182 XThC.XTBN.Y a_9827_9569# 0.22873f
C1183 XThR.Tn[2] XA.XIR[2].XIC[13].icell.Ien 0.14211f
C1184 XThR.XTB7.A a_n1049_7493# 0.0127f
C1185 XA.XIR[3].XIC[1].icell.PDM VPWR 0.01171f
C1186 XA.XIR[10].XIC[8].icell.Ien Vbias 0.19161f
C1187 XThC.XTB5.Y XThC.XTB7.B 0.30234f
C1188 XA.XIR[8].XIC[3].icell.PDM VPWR 0.01171f
C1189 XA.XIR[4].XIC[12].icell.Ien VPWR 0.18829f
C1190 XA.XIR[2].XIC[7].icell.PDM VPWR 0.01171f
C1191 XA.XIR[14].XIC[1].icell.Ien XThR.Tn[14] 0.14211f
C1192 XA.XIR[7].XIC[12].icell.Ien Iout 0.06801f
C1193 XA.XIR[8].XIC[6].icell.Ien VPWR 0.18829f
C1194 XThR.XTB7.A XThR.XTB6.Y 0.19112f
C1195 XA.XIR[2].XIC[10].icell.Ien Vbias 0.19161f
C1196 XThR.Tn[11] XA.XIR[12].XIC[7].icell.PDM 0.04035f
C1197 XA.XIR[10].XIC[11].icell.Ien Iout 0.06801f
C1198 XA.XIR[12].XIC[11].icell.PDM XA.XIR[12].XIC[11].icell.Ien 0.04854f
C1199 XA.XIR[9].XIC_15.icell.Ien VPWR 0.26829f
C1200 XA.XIR[3].XIC[1].icell.Ien Iout 0.06801f
C1201 XA.XIR[2].XIC[9].icell.Ien XA.XIR[3].XIC[9].icell.PDM 0.02104f
C1202 XA.XIR[1].XIC[12].icell.Ien Vbias 0.19173f
C1203 XA.XIR[3].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1204 XThR.XTB7.B XThR.XTBN.A 0.35142f
C1205 XA.XIR[7].XIC[10].icell.Ien XA.XIR[8].XIC[10].icell.PDM 0.02104f
C1206 XThR.Tn[9] XA.XIR[9].XIC[11].icell.Ien 0.14211f
C1207 XThR.XTB7.Y XThR.Tn[11] 0.07412f
C1208 XA.XIR[0].XIC[8].icell.Ien VPWR 0.18959f
C1209 XThC.XTB7.B XThC.XTBN.Y 0.38751f
C1210 XThR.XTB7.B XThR.Tn[6] 0.04822f
C1211 XA.XIR[1].XIC[12].icell.Ien XA.XIR[2].XIC[12].icell.PDM 0.02104f
C1212 XThR.Tn[0] XA.XIR[1].XIC[5].icell.PDM 0.04035f
C1213 XA.XIR[12].XIC[10].icell.Ien VPWR 0.18829f
C1214 XA.XIR[9].XIC_dummy_left.icell.Iout Iout 0.03553f
C1215 XThR.Tn[1] XA.XIR[2].XIC[4].icell.PDM 0.04035f
C1216 XA.XIR[7].XIC[11].icell.Ien VPWR 0.18829f
C1217 XThC.Tn[12] XThR.Tn[7] 0.40738f
C1218 XA.XIR[15].XIC[13].icell.PDM XA.XIR[15].XIC[13].icell.Ien 0.04854f
C1219 XA.XIR[7].XIC[6].icell.PDM Vbias 0.03928f
C1220 XThR.Tn[7] XA.XIR[8].XIC[9].icell.PDM 0.04035f
C1221 XThC.Tn[8] XA.XIR[11].XIC[8].icell.PDM 0.02601f
C1222 XA.XIR[6].XIC[10].icell.PDM XA.XIR[6].XIC[10].icell.Ien 0.04854f
C1223 XThC.XTB7.B XThC.Tn[10] 0.0672f
C1224 XA.XIR[9].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1225 XThC.XTB7.Y XThC.Tn[14] 0.4237f
C1226 XA.XIR[6].XIC[13].icell.PDM Vbias 0.03928f
C1227 XA.XIR[15].XIC[9].icell.PDM XA.XIR[15].XIC[9].icell.Ien 0.04854f
C1228 XA.XIR[15].XIC[4].icell.PDM Vbias 0.03928f
C1229 XA.XIR[3].XIC[0].icell.Ien VPWR 0.18829f
C1230 XThR.Tn[6] XA.XIR[6].XIC[1].icell.Ien 0.14211f
C1231 XThR.Tn[8] VPWR 8.93422f
C1232 XThC.Tn[12] XA.XIR[6].XIC[12].icell.PDM 0.02601f
C1233 XThC.Tn[13] XA.XIR[14].XIC[13].icell.Ien 0.04604f
C1234 XA.XIR[10].XIC[3].icell.Ien XA.XIR[11].XIC[3].icell.PDM 0.02104f
C1235 XA.XIR[13].XIC[13].icell.Ien Iout 0.06801f
C1236 XA.XIR[14].XIC[10].icell.PDM Vbias 0.03928f
C1237 XA.XIR[9].XIC[9].icell.Ien XA.XIR[10].XIC[9].icell.PDM 0.02104f
C1238 XA.XIR[13].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1239 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[2].XIC_dummy_right.icell.PDM 0.02104f
C1240 XThC.Tn[9] XA.XIR[3].XIC[9].icell.PDM 0.02601f
C1241 XA.XIR[10].XIC[4].icell.PDM XA.XIR[10].XIC[4].icell.Ien 0.04854f
C1242 bias[0] Vbias 0.82324f
C1243 XA.XIR[11].XIC[1].icell.Ien VPWR 0.18829f
C1244 XThR.XTB3.Y data[4] 0.03253f
C1245 XThR.Tn[11] XA.XIR[11].XIC[7].icell.Ien 0.14211f
C1246 XThC.Tn[8] XA.XIR[15].XIC[8].icell.Ien 0.04292f
C1247 XA.XIR[9].XIC[2].icell.PDM Vbias 0.03928f
C1248 XThR.Tn[3] XA.XIR[4].XIC[10].icell.PDM 0.04035f
C1249 XThC.Tn[4] XA.XIR[0].XIC[4].icell.Ien 0.04658f
C1250 XA.XIR[7].XIC[7].icell.PDM VPWR 0.01171f
C1251 XThR.XTB2.Y XThR.XTB3.Y 2.04808f
C1252 a_3773_9615# XThC.Tn[1] 0.26251f
C1253 XThR.Tn[14] a_n997_715# 0.1927f
C1254 XA.XIR[12].XIC[13].icell.Ien Vbias 0.19161f
C1255 XA.XIR[3].XIC[9].icell.Ien Iout 0.06801f
C1256 XA.XIR[6].XIC[14].icell.PDM VPWR 0.0118f
C1257 XThR.Tn[0] XA.XIR[0].XIC[12].icell.Ien 0.14211f
C1258 XA.XIR[15].XIC[5].icell.PDM VPWR 0.01512f
C1259 XThR.Tn[11] a_n997_2667# 0.19413f
C1260 XThC.Tn[9] XA.XIR[11].XIC[9].icell.Ien 0.04604f
C1261 XThR.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.14211f
C1262 XA.XIR[9].XIC_dummy_right.icell.Iout XA.XIR[10].XIC_dummy_right.icell.Iout 0.04047f
C1263 XThC.Tn[11] XThR.Tn[3] 0.40738f
C1264 XA.XIR[2].XIC[2].icell.Ien Iout 0.06801f
C1265 XA.XIR[15].XIC[14].icell.Ien VPWR 0.31908f
C1266 XA.XIR[1].XIC[7].icell.PDM Vbias 0.03928f
C1267 XThR.Tn[2] XA.XIR[2].XIC_dummy_left.icell.Ien 0.01569f
C1268 XA.XIR[1].XIC[4].icell.Ien Iout 0.06801f
C1269 XA.XIR[6].XIC[12].icell.Ien Vbias 0.19161f
C1270 XThR.Tn[7] XA.XIR[7].XIC[13].icell.Ien 0.14211f
C1271 XA.XIR[9].XIC[3].icell.PDM VPWR 0.01171f
C1272 XA.XIR[9].XIC[13].icell.PDM XA.XIR[9].XIC[13].icell.Ien 0.04854f
C1273 XA.XIR[4].XIC[7].icell.PDM Vbias 0.03928f
C1274 XA.XIR[7].XIC[11].icell.PDM XA.XIR[7].XIC[11].icell.Ien 0.04854f
C1275 XThC.Tn[6] XA.XIR[4].XIC[6].icell.Ien 0.04604f
C1276 XA.XIR[8].XIC[12].icell.Ien Iout 0.06801f
C1277 XThC.Tn[2] XA.XIR[1].XIC[2].icell.PDM 0.02602f
C1278 XA.XIR[4].XIC[12].icell.PDM XA.XIR[4].XIC[12].icell.Ien 0.04854f
C1279 XA.XIR[2].XIC[2].icell.Ien XA.XIR[3].XIC[2].icell.PDM 0.02104f
C1280 XThC.XTB4.Y a_8963_9569# 0.07199f
C1281 XA.XIR[3].XIC_15.icell.PDM Vbias 0.03927f
C1282 XThC.Tn[14] XThR.Tn[0] 0.40766f
C1283 XA.XIR[14].XIC[6].icell.Ien Vbias 0.19161f
C1284 XA.XIR[7].XIC[3].icell.Ien XA.XIR[8].XIC[3].icell.PDM 0.02104f
C1285 XA.XIR[5].XIC[1].icell.Ien XA.XIR[6].XIC[1].icell.PDM 0.02104f
C1286 XThC.Tn[2] XA.XIR[4].XIC[2].icell.PDM 0.02601f
C1287 XThR.Tn[4] XA.XIR[5].XIC[2].icell.PDM 0.04035f
C1288 XA.XIR[13].XIC[8].icell.Ien Vbias 0.19161f
C1289 XThR.XTB7.B XThR.XTB6.Y 0.30244f
C1290 XA.XIR[3].XIC[8].icell.Ien VPWR 0.18829f
C1291 XA.XIR[10].XIC[0].icell.PDM XA.XIR[10].XIC[0].icell.Ien 0.04854f
C1292 XA.XIR[1].XIC[8].icell.PDM VPWR 0.01171f
C1293 XA.XIR[1].XIC[5].icell.Ien XA.XIR[2].XIC[5].icell.PDM 0.02104f
C1294 XA.XIR[8].XIC[10].icell.PDM XA.XIR[8].XIC[10].icell.Ien 0.04854f
C1295 XA.XIR[4].XIC[8].icell.PDM VPWR 0.01171f
C1296 XA.XIR[0].XIC[14].icell.Ien Iout 0.0675f
C1297 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[1].XIC_dummy_left.icell.Iout 0.06446f
C1298 XThR.Tn[13] XA.XIR[14].XIC[4].icell.PDM 0.04035f
C1299 XThR.XTBN.Y XThR.XTBN.A 0.77119f
C1300 XA.XIR[0].XIC[9].icell.Ien XA.XIR[1].XIC[9].icell.PDM 0.02104f
C1301 XA.XIR[1].XIC[3].icell.Ien VPWR 0.18829f
C1302 XA.XIR[3].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1303 XThC.Tn[1] XA.XIR[8].XIC[1].icell.PDM 0.02601f
C1304 XThC.XTB7.Y a_6243_10571# 0.01283f
C1305 XA.XIR[6].XIC[3].icell.PDM XA.XIR[6].XIC[3].icell.Ien 0.04854f
C1306 XA.XIR[13].XIC[11].icell.Ien Iout 0.06801f
C1307 XA.XIR[4].XIC_dummy_right.icell.PDM XA.XIR[4].XIC_dummy_right.icell.Ien 0.04854f
C1308 a_n1049_7493# XThR.Tn[2] 0.26564f
C1309 XA.XIR[15].XIC[2].icell.PDM XA.XIR[15].XIC[2].icell.Ien 0.04854f
C1310 XA.XIR[12].XIC_15.icell.Ien VPWR 0.26829f
C1311 XThR.XTBN.Y XThR.Tn[6] 0.59897f
C1312 XThR.Tn[8] XA.XIR[9].XIC[7].icell.PDM 0.04035f
C1313 XA.XIR[8].XIC[11].icell.Ien VPWR 0.18829f
C1314 XThR.XTB7.Y XThR.Tn[14] 0.4222f
C1315 XA.XIR[9].XIC[2].icell.Ien XA.XIR[10].XIC[2].icell.PDM 0.02104f
C1316 VPWR data[4] 0.5303f
C1317 XA.XIR[12].XIC_dummy_right.icell.PDM XA.XIR[12].XIC_dummy_right.icell.Ien 0.04854f
C1318 XThC.Tn[13] XThR.Tn[2] 0.40742f
C1319 XA.XIR[2].XIC_15.icell.Ien Vbias 0.19195f
C1320 XA.XIR[12].XIC[11].icell.Ien Vbias 0.19161f
C1321 XThR.XTB4.Y XThR.XTBN.A 0.03415f
C1322 XThR.XTB2.Y VPWR 0.99055f
C1323 a_n997_3755# VPWR 0.0133f
C1324 XThR.Tn[5] XA.XIR[6].XIC[4].icell.PDM 0.04035f
C1325 XA.XIR[15].XIC[12].icell.Ien VPWR 0.31713f
C1326 XThC.Tn[3] XA.XIR[11].XIC[3].icell.PDM 0.02601f
C1327 XA.XIR[0].XIC[13].icell.Ien VPWR 0.18776f
C1328 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.Iout 0.06446f
C1329 XThC.Tn[4] XA.XIR[3].XIC[4].icell.Ien 0.04604f
C1330 XThR.XTB5.Y XThR.Tn[5] 0.01094f
C1331 XA.XIR[6].XIC[4].icell.Ien Iout 0.06801f
C1332 XThR.XTBN.A XThR.Tn[10] 0.12147f
C1333 XThC.Tn[8] XA.XIR[14].XIC[8].icell.PDM 0.02601f
C1334 XA.XIR[10].XIC[1].icell.PDM Vbias 0.03928f
C1335 XThR.Tn[14] XA.XIR[14].XIC[2].icell.Ien 0.14211f
C1336 XThC.Tn[11] XA.XIR[2].XIC[11].icell.Ien 0.04605f
C1337 XThR.Tn[1] XA.XIR[1].XIC[2].icell.Ien 0.14211f
C1338 XA.XIR[12].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1339 XThC.Tn[7] XA.XIR[6].XIC[7].icell.PDM 0.02601f
C1340 data[6] data[7] 0.04128f
C1341 XThR.Tn[6] XA.XIR[7].XIC[3].icell.PDM 0.04035f
C1342 XA.XIR[2].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1343 XThC.Tn[14] XA.XIR[2].XIC[14].icell.PDM 0.02602f
C1344 XThC.Tn[4] XA.XIR[3].XIC[4].icell.PDM 0.02601f
C1345 XA.XIR[6].XIC[12].icell.Ien XA.XIR[7].XIC[12].icell.PDM 0.02104f
C1346 XThR.Tn[13] XA.XIR[13].XIC[6].icell.Ien 0.14211f
C1347 a_n1049_5611# VPWR 0.71817f
C1348 XA.XIR[5].XIC[5].icell.Ien Vbias 0.19161f
C1349 XThC.Tn[9] XThR.Tn[6] 0.40738f
C1350 XA.XIR[9].XIC[6].icell.PDM XA.XIR[9].XIC[6].icell.Ien 0.04854f
C1351 XA.XIR[7].XIC[4].icell.PDM XA.XIR[7].XIC[4].icell.Ien 0.04854f
C1352 XA.XIR[14].XIC[1].icell.Ien VPWR 0.18883f
C1353 XA.XIR[4].XIC[5].icell.PDM XA.XIR[4].XIC[5].icell.Ien 0.04854f
C1354 XA.XIR[10].XIC[2].icell.PDM VPWR 0.01171f
C1355 XThC.Tn[11] XThR.Tn[11] 0.40738f
C1356 XA.XIR[11].XIC[3].icell.Ien Iout 0.06801f
C1357 XA.XIR[14].XIC[7].icell.Ien XA.XIR[15].XIC[7].icell.PDM 0.02104f
C1358 XThR.XTBN.Y XThR.Tn[4] 0.6035f
C1359 XThC.Tn[9] XA.XIR[14].XIC[9].icell.Ien 0.04604f
C1360 XThC.Tn[1] XThR.Tn[7] 0.40738f
C1361 XA.XIR[10].XIC[5].icell.Ien Iout 0.06801f
C1362 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.PDM 0.02104f
C1363 XA.XIR[6].XIC[3].icell.Ien VPWR 0.18829f
C1364 XThR.Tn[5] Vbias 1.39526f
C1365 XA.XIR[8].XIC[3].icell.PDM XA.XIR[8].XIC[3].icell.Ien 0.04854f
C1366 XThR.XTBN.Y a_n1049_7493# 0.08456f
C1367 XA.XIR[0].XIC[9].icell.PDM Vbias 0.03945f
C1368 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[7].XIC_dummy_right.icell.PDM 0.02104f
C1369 XThC.XTB7.B a_7651_9569# 0.01152f
C1370 XA.XIR[0].XIC[2].icell.Ien XA.XIR[1].XIC[2].icell.PDM 0.02104f
C1371 XA.XIR[3].XIC[14].icell.Ien Iout 0.06801f
C1372 XThC.XTB5.Y XThC.Tn[12] 0.32158f
C1373 XThR.Tn[9] XA.XIR[9].XIC_dummy_left.icell.Iout 0.03386f
C1374 XThR.XTBN.Y XThR.XTB6.Y 0.1894f
C1375 XA.XIR[8].XIC[10].icell.Ien XA.XIR[9].XIC[10].icell.PDM 0.02104f
C1376 XThR.Tn[6] XA.XIR[6].XIC[11].icell.Ien 0.14211f
C1377 XA.XIR[2].XIC[7].icell.Ien Iout 0.06801f
C1378 XThC.Tn[14] XThR.Tn[1] 0.40747f
C1379 XThC.Tn[2] XA.XIR[10].XIC[2].icell.Ien 0.04604f
C1380 XA.XIR[3].XIC[9].icell.Ien XA.XIR[4].XIC[9].icell.PDM 0.02104f
C1381 XA.XIR[15].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.Iout 0.06446f
C1382 XThC.Tn[1] XA.XIR[9].XIC[1].icell.PDM 0.02601f
C1383 XA.XIR[1].XIC[9].icell.Ien Iout 0.06801f
C1384 XA.XIR[2].XIC[1].icell.Ien VPWR 0.18829f
C1385 XThR.XTB3.Y XThR.Tn[3] 0.01287f
C1386 XA.XIR[0].XIC[10].icell.PDM VPWR 0.01132f
C1387 XA.XIR[7].XIC_dummy_left.icell.Iout VPWR 0.10954f
C1388 XA.XIR[3].XIC[11].icell.PDM XA.XIR[3].XIC[11].icell.Ien 0.04854f
C1389 XA.XIR[11].XIC[2].icell.Ien VPWR 0.18829f
C1390 XA.XIR[15].XIC[10].icell.Ien VPWR 0.31713f
C1391 XThC.Tn[14] XThR.Tn[12] 0.40742f
C1392 XA.XIR[10].XIC[4].icell.Ien VPWR 0.18829f
C1393 XThC.XTB7.A VPWR 0.87269f
C1394 XThC.Tn[0] XThR.Tn[3] 0.40742f
C1395 XThC.Tn[5] XA.XIR[5].XIC[5].icell.Ien 0.04604f
C1396 XThR.XTBN.A a_n997_1803# 0.09118f
C1397 XThC.XTBN.Y XThC.Tn[12] 0.46758f
C1398 XThR.Tn[10] XA.XIR[11].XIC[6].icell.PDM 0.04035f
C1399 XThC.Tn[9] XThR.Tn[4] 0.40738f
C1400 XThR.XTB3.Y XThR.XTB7.Y 0.03772f
C1401 XThR.XTB4.Y XThR.XTB6.Y 0.04273f
C1402 XThC.Tn[14] XA.XIR[7].XIC[14].icell.PDM 0.02601f
C1403 XThR.Tn[14] XA.XIR[15].XIC[7].icell.PDM 0.04035f
C1404 XA.XIR[3].XIC[13].icell.Ien VPWR 0.18829f
C1405 XThR.XTB6.Y XThR.Tn[10] 0.02461f
C1406 XThC.Tn[13] XThR.Tn[10] 0.40739f
C1407 XA.XIR[2].XIC[6].icell.Ien VPWR 0.18829f
C1408 XThC.Tn[3] XThR.Tn[0] 0.40763f
C1409 a_n997_715# VPWR 0.02818f
C1410 XThC.Tn[5] XThR.Tn[5] 0.40738f
C1411 XA.XIR[6].XIC[5].icell.Ien XA.XIR[7].XIC[5].icell.PDM 0.02104f
C1412 XA.XIR[1].XIC[8].icell.Ien VPWR 0.18829f
C1413 XThR.Tn[8] XA.XIR[8].XIC[3].icell.Ien 0.14211f
C1414 XA.XIR[9].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1415 XThR.Tn[10] XA.XIR[10].XIC_dummy_left.icell.Iout 0.03385f
C1416 XA.XIR[6].XIC[0].icell.PDM Vbias 0.03915f
C1417 XA.XIR[15].XIC[13].icell.Ien Vbias 0.15966f
C1418 XThC.Tn[3] XA.XIR[14].XIC[3].icell.PDM 0.02601f
C1419 XA.XIR[5].XIC[7].icell.PDM Vbias 0.03928f
C1420 XA.XIR[13].XIC[1].icell.PDM Vbias 0.03928f
C1421 XA.XIR[4].XIC[12].icell.Ien XA.XIR[5].XIC[12].icell.PDM 0.02104f
C1422 XThR.Tn[5] XA.XIR[5].XIC[2].icell.Ien 0.14211f
C1423 XA.XIR[12].XIC[6].icell.PDM Vbias 0.03928f
C1424 XThC.Tn[2] XA.XIR[5].XIC[2].icell.PDM 0.02601f
C1425 XA.XIR[13].XIC[3].icell.Ien XA.XIR[14].XIC[3].icell.PDM 0.02104f
C1426 a_5949_9615# VPWR 0.7053f
C1427 XThC.Tn[3] XA.XIR[9].XIC[3].icell.Ien 0.04604f
C1428 XThC.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.04604f
C1429 XA.XIR[6].XIC[1].icell.PDM VPWR 0.01171f
C1430 XA.XIR[13].XIC[4].icell.PDM XA.XIR[13].XIC[4].icell.Ien 0.04854f
C1431 XThR.Tn[2] XA.XIR[3].XIC[11].icell.PDM 0.04035f
C1432 XA.XIR[6].XIC[9].icell.Ien Iout 0.06801f
C1433 XThC.Tn[10] XA.XIR[0].XIC[10].icell.Ien 0.04662f
C1434 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[8].XIC_dummy_left.icell.PDM 0.02104f
C1435 XThR.Tn[14] XA.XIR[14].XIC[7].icell.Ien 0.14211f
C1436 XA.XIR[5].XIC[8].icell.PDM VPWR 0.01171f
C1437 XThR.Tn[1] XA.XIR[1].XIC[7].icell.Ien 0.14211f
C1438 XA.XIR[8].XIC[3].icell.Ien XA.XIR[9].XIC[3].icell.PDM 0.02104f
C1439 XA.XIR[12].XIC[5].icell.Ien XA.XIR[13].XIC[5].icell.PDM 0.02104f
C1440 XThC.Tn[2] XThR.Tn[2] 0.40741f
C1441 Vbias Iout 74.00211f
C1442 XA.XIR[13].XIC[2].icell.PDM VPWR 0.01171f
C1443 XA.XIR[3].XIC[2].icell.Ien XA.XIR[4].XIC[2].icell.PDM 0.02104f
C1444 XThC.Tn[4] XA.XIR[1].XIC[4].icell.Ien 0.04607f
C1445 XThR.Tn[3] VPWR 8.06517f
C1446 XThC.Tn[11] XThR.Tn[14] 0.40738f
C1447 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.Iout 0.06446f
C1448 XThC.XTB6.Y Vbias 0.01779f
C1449 XA.XIR[14].XIC[3].icell.Ien Iout 0.06801f
C1450 XThC.XTB5.A VPWR 0.82807f
C1451 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[5].XIC_dummy_right.icell.PDM 0.02104f
C1452 XA.XIR[3].XIC[4].icell.PDM XA.XIR[3].XIC[4].icell.Ien 0.04854f
C1453 XA.XIR[11].XIC[13].icell.PDM XA.XIR[11].XIC[13].icell.Ien 0.04854f
C1454 XA.XIR[12].XIC[7].icell.PDM VPWR 0.01171f
C1455 XA.XIR[5].XIC[10].icell.Ien Vbias 0.19161f
C1456 XA.XIR[12].XIC_dummy_right.icell.Iout XA.XIR[13].XIC_dummy_right.icell.Iout 0.04047f
C1457 XA.XIR[13].XIC[5].icell.Ien Iout 0.06801f
C1458 XA.XIR[3].XIC[2].icell.PDM Vbias 0.03928f
C1459 XA.XIR[11].XIC[9].icell.PDM XA.XIR[11].XIC[9].icell.Ien 0.04854f
C1460 XA.XIR[8].XIC[4].icell.PDM Vbias 0.03928f
C1461 XThR.XTB7.Y VPWR 1.14768f
C1462 XThC.Tn[12] XA.XIR[4].XIC[12].icell.Ien 0.04604f
C1463 XA.XIR[2].XIC[8].icell.PDM Vbias 0.03928f
C1464 XThR.XTB5.A XThR.XTB5.Y 0.0538f
C1465 XA.XIR[8].XIC_dummy_left.icell.Iout VPWR 0.11f
C1466 XA.XIR[11].XIC[8].icell.Ien Iout 0.06801f
C1467 XA.XIR[15].XIC[11].icell.PDM XA.XIR[15].XIC[11].icell.Ien 0.04854f
C1468 XA.XIR[15].XIC_15.icell.Ien VPWR 0.37868f
C1469 XA.XIR[5].XIC[0].icell.PDM XA.XIR[5].XIC[0].icell.Ien 0.04854f
C1470 XThR.Tn[9] XA.XIR[10].XIC[5].icell.PDM 0.04035f
C1471 XA.XIR[12].XIC[5].icell.Ien Vbias 0.19161f
C1472 XA.XIR[6].XIC[8].icell.Ien VPWR 0.18829f
C1473 XThC.Tn[7] XThR.Tn[6] 0.40738f
C1474 XThC.Tn[0] XA.XIR[12].XIC[0].icell.Ien 0.04604f
C1475 XThC.Tn[2] XA.XIR[13].XIC[2].icell.Ien 0.04604f
C1476 XThC.XTBN.A XThC.Tn[9] 0.12399f
C1477 XThC.XTBN.Y a_10915_9569# 0.21503f
C1478 XThC.Tn[0] XThR.Tn[11] 0.4074f
C1479 XA.XIR[3].XIC[3].icell.PDM VPWR 0.01171f
C1480 XA.XIR[8].XIC[5].icell.PDM VPWR 0.01171f
C1481 XA.XIR[14].XIC[2].icell.Ien VPWR 0.18883f
C1482 XA.XIR[15].XIC[11].icell.Ien Vbias 0.15966f
C1483 XA.XIR[13].XIC[0].icell.PDM XA.XIR[13].XIC[0].icell.Ien 0.04854f
C1484 XThC.XTB4.Y Vbias 0.01644f
C1485 XThC.XTB7.A XThC.XTB7.B 0.35844f
C1486 XA.XIR[2].XIC[9].icell.PDM VPWR 0.01171f
C1487 XA.XIR[13].XIC[4].icell.Ien VPWR 0.18829f
C1488 XA.XIR[12].XIC[1].icell.Ien XA.XIR[13].XIC[1].icell.PDM 0.02104f
C1489 XA.XIR[2].XIC[12].icell.Ien Iout 0.06801f
C1490 XThC.Tn[5] Iout 0.22432f
C1491 XA.XIR[1].XIC[14].icell.Ien Iout 0.06801f
C1492 XThC.Tn[1] XA.XIR[7].XIC[1].icell.Ien 0.04604f
C1493 XThC.Tn[9] XA.XIR[6].XIC[9].icell.PDM 0.02601f
C1494 XA.XIR[15].XIC_dummy_right.icell.Iout VPWR 0.21463f
C1495 XA.XIR[10].XIC_15.icell.PUM VPWR 0.01655f
C1496 XA.XIR[4].XIC[5].icell.Ien XA.XIR[5].XIC[5].icell.PDM 0.02104f
C1497 XA.XIR[1].XIC[9].icell.PDM XA.XIR[1].XIC[9].icell.Ien 0.04854f
C1498 VPWR data[0] 0.52929f
C1499 XA.XIR[11].XIC[7].icell.Ien VPWR 0.18829f
C1500 XThR.Tn[11] XA.XIR[12].XIC[9].icell.PDM 0.04035f
C1501 XA.XIR[9].XIC_15.icell.Ien XA.XIR[10].XIC_15.icell.PDM 0.02104f
C1502 XThC.XTB6.Y XThC.Tn[5] 0.20249f
C1503 XA.XIR[3].XIC_dummy_left.icell.Iout Iout 0.03553f
C1504 XThR.XTB6.Y XThR.Tn[13] 0.32265f
C1505 XA.XIR[10].XIC[9].icell.Ien VPWR 0.18829f
C1506 XThC.Tn[13] XThR.Tn[13] 0.40739f
C1507 XA.XIR[12].XIC[1].icell.Ien Iout 0.06801f
C1508 XThC.Tn[3] XThR.Tn[1] 0.40744f
C1509 a_n997_2667# VPWR 0.01642f
C1510 XA.XIR[2].XIC[11].icell.PDM XA.XIR[2].XIC[11].icell.Ien 0.04854f
C1511 XThC.Tn[4] XA.XIR[6].XIC[4].icell.Ien 0.04604f
C1512 XA.XIR[12].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1513 XThR.XTB5.A XThR.XTB1.Y 0.1098f
C1514 XThR.Tn[0] XA.XIR[1].XIC[7].icell.PDM 0.04035f
C1515 XThC.Tn[3] XThR.Tn[12] 0.40738f
C1516 XA.XIR[5].XIC[2].icell.Ien Iout 0.06801f
C1517 XThC.Tn[12] XThR.Tn[8] 0.40738f
C1518 XThC.Tn[10] XA.XIR[3].XIC[10].icell.Ien 0.04604f
C1519 XA.XIR[15].XIC_dummy_left.icell.Ien VPWR 0.38522f
C1520 XThR.Tn[1] XA.XIR[2].XIC[6].icell.PDM 0.04035f
C1521 XA.XIR[2].XIC[11].icell.Ien VPWR 0.18829f
C1522 XThC.Tn[5] XA.XIR[12].XIC[5].icell.Ien 0.04604f
C1523 XThC.XTBN.Y XThC.Tn[1] 0.49539f
C1524 XA.XIR[1].XIC[13].icell.Ien VPWR 0.18829f
C1525 XA.XIR[7].XIC[8].icell.PDM Vbias 0.03928f
C1526 XThR.Tn[7] XA.XIR[8].XIC[11].icell.PDM 0.04035f
C1527 XThR.Tn[8] XA.XIR[8].XIC[8].icell.Ien 0.14211f
C1528 XA.XIR[9].XIC[1].icell.Ien Vbias 0.19161f
C1529 XA.XIR[11].XIC[2].icell.PDM XA.XIR[11].XIC[2].icell.Ien 0.04854f
C1530 XThC.Tn[7] XThR.Tn[4] 0.40738f
C1531 XA.XIR[6].XIC_15.icell.PDM Vbias 0.03927f
C1532 XA.XIR[4].XIC[3].icell.Ien Vbias 0.19161f
C1533 XA.XIR[15].XIC[6].icell.PDM Vbias 0.03928f
C1534 XThR.Tn[6] XA.XIR[6].XIC_dummy_left.icell.Iout 0.03777f
C1535 XThC.Tn[2] XThR.Tn[10] 0.40738f
C1536 XA.XIR[5].XIC[14].icell.PDM XA.XIR[5].XIC[14].icell.Ien 0.04854f
C1537 XA.XIR[12].XIC[0].icell.Ien VPWR 0.18829f
C1538 XThC.XTB6.Y a_10051_9569# 0.07626f
C1539 XThR.Tn[11] VPWR 9.00382f
C1540 XThR.Tn[5] XA.XIR[5].XIC[7].icell.Ien 0.14211f
C1541 XA.XIR[9].XIC[4].icell.PDM Vbias 0.03928f
C1542 XThR.Tn[3] XA.XIR[4].XIC[12].icell.PDM 0.04035f
C1543 XA.XIR[7].XIC[9].icell.PDM VPWR 0.01171f
C1544 XThC.XTB2.Y Vbias 0.01484f
C1545 XThC.XTB5.A XThC.XTB7.B 0.30355f
C1546 XA.XIR[9].XIC[6].icell.Ien Vbias 0.19161f
C1547 XA.XIR[15].XIC[7].icell.PDM VPWR 0.01512f
C1548 XA.XIR[6].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1549 XA.XIR[6].XIC[14].icell.Ien Iout 0.06801f
C1550 XThR.Tn[1] XA.XIR[1].XIC[12].icell.Ien 0.14211f
C1551 XA.XIR[1].XIC[9].icell.PDM Vbias 0.03928f
C1552 XThR.XTB5.Y XThR.Tn[9] 0.01732f
C1553 XA.XIR[9].XIC[5].icell.PDM VPWR 0.01171f
C1554 XA.XIR[14].XIC[8].icell.Ien Iout 0.06801f
C1555 XA.XIR[4].XIC[9].icell.PDM Vbias 0.03928f
C1556 XA.XIR[1].XIC[2].icell.PDM XA.XIR[1].XIC[2].icell.Ien 0.04854f
C1557 XA.XIR[5].XIC_15.icell.Ien Vbias 0.19195f
C1558 XA.XIR[7].XIC[2].icell.Ien Vbias 0.19161f
C1559 XThC.Tn[8] XA.XIR[10].XIC[8].icell.Ien 0.04604f
C1560 XThR.XTBN.A a_n997_3979# 0.02087f
C1561 XA.XIR[12].XIC_15.icell.PDM Vbias 0.03927f
C1562 XThC.Tn[1] XA.XIR[8].XIC[1].icell.Ien 0.04604f
C1563 XA.XIR[2].XIC[4].icell.PDM XA.XIR[2].XIC[4].icell.Ien 0.04854f
C1564 XA.XIR[12].XIC[14].icell.Ien XA.XIR[13].XIC[14].icell.PDM 0.02104f
C1565 XA.XIR[15].XIC_dummy_right.icell.PDM XA.XIR[15].XIC_dummy_right.icell.Ien 0.04854f
C1566 XThC.Tn[0] XThR.Tn[14] 0.40739f
C1567 XThR.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.04035f
C1568 XThC.Tn[0] XA.XIR[11].XIC[0].icell.PDM 0.02601f
C1569 XA.XIR[14].XIC[0].icell.Ien XA.XIR[15].XIC[0].icell.PDM 0.02104f
C1570 XA.XIR[1].XIC[10].icell.PDM VPWR 0.01171f
C1571 XThC.Tn[11] XA.XIR[5].XIC[11].icell.Ien 0.04604f
C1572 XA.XIR[6].XIC[13].icell.Ien VPWR 0.18829f
C1573 XA.XIR[10].XIC[14].icell.Ien VPWR 0.18835f
C1574 XA.XIR[5].XIC_dummy_right.icell.PUM VPWR 0.01691f
C1575 XA.XIR[4].XIC[10].icell.PDM VPWR 0.01171f
C1576 XThC.Tn[4] XA.XIR[6].XIC[4].icell.PDM 0.02601f
C1577 XThR.Tn[13] XA.XIR[14].XIC[6].icell.PDM 0.04035f
C1578 XThC.Tn[11] XA.XIR[2].XIC[11].icell.PDM 0.02602f
C1579 XThC.Tn[1] XA.XIR[3].XIC[1].icell.PDM 0.02601f
C1580 XThR.Tn[9] Vbias 1.39532f
C1581 XThC.XTB7.B data[0] 0.0138f
C1582 XA.XIR[13].XIC_15.icell.PUM VPWR 0.01655f
C1583 XA.XIR[14].XIC[7].icell.Ien VPWR 0.18883f
C1584 XA.XIR[12].XIC_dummy_right.icell.PDM VPWR 0.08209f
C1585 XThR.Tn[8] XA.XIR[9].XIC[9].icell.PDM 0.04035f
C1586 XA.XIR[13].XIC[9].icell.Ien VPWR 0.18829f
C1587 XThC.Tn[11] VPWR 4.57828f
C1588 XThC.Tn[12] XA.XIR[15].XIC[12].icell.Ien 0.04292f
C1589 XA.XIR[5].XIC[7].icell.PDM XA.XIR[5].XIC[7].icell.Ien 0.04854f
C1590 XA.XIR[15].XIC_dummy_left.icell.PUM VPWR 0.01604f
C1591 XThC.XTBN.A XThC.Tn[7] 0.01451f
C1592 XThR.Tn[13] XA.XIR[13].XIC_dummy_left.icell.Iout 0.03385f
C1593 XThR.Tn[12] XA.XIR[12].XIC[13].icell.Ien 0.14211f
C1594 XThR.XTB6.A data[5] 0.37233f
C1595 XA.XIR[15].XIC[0].icell.Ien Vbias 0.15953f
C1596 XThR.Tn[5] XA.XIR[6].XIC[6].icell.PDM 0.04035f
C1597 XThR.XTBN.A XThR.Tn[7] 0.01439f
C1598 XThR.XTBN.A a_n997_2891# 0.01719f
C1599 VPWR bias[2] 1.67895f
C1600 XThR.Tn[6] XThR.Tn[7] 0.11401f
C1601 XA.XIR[10].XIC[3].icell.PDM Vbias 0.03928f
C1602 XThC.Tn[4] Vbias 0.84011f
C1603 XThC.Tn[9] XA.XIR[9].XIC[9].icell.Ien 0.04604f
C1604 XA.XIR[5].XIC[7].icell.Ien Iout 0.06801f
C1605 XThR.Tn[10] XA.XIR[11].XIC[14].icell.PDM 0.04056f
C1606 XThR.Tn[6] XA.XIR[7].XIC[5].icell.PDM 0.04035f
C1607 XA.XIR[12].XIC[3].icell.PDM XA.XIR[12].XIC[3].icell.Ien 0.04854f
C1608 XThC.Tn[2] XThR.Tn[13] 0.40738f
C1609 XA.XIR[5].XIC[1].icell.Ien VPWR 0.18829f
C1610 XA.XIR[15].XIC[5].icell.Ien Vbias 0.15966f
C1611 XThR.Tn[8] XA.XIR[8].XIC[13].icell.Ien 0.14211f
C1612 XThR.Tn[14] VPWR 9.25423f
C1613 XThC.Tn[10] XA.XIR[1].XIC[10].icell.Ien 0.04606f
C1614 XA.XIR[11].XIC[0].icell.PDM VPWR 0.01171f
C1615 XA.XIR[4].XIC[8].icell.Ien Vbias 0.19161f
C1616 XThC.Tn[5] XThR.Tn[9] 0.40738f
C1617 XA.XIR[12].XIC[2].icell.Ien Iout 0.06801f
C1618 XThC.Tn[1] XThR.Tn[8] 0.40738f
C1619 XA.XIR[10].XIC[4].icell.PDM VPWR 0.01171f
C1620 XThR.XTB2.Y a_n1335_8107# 0.01006f
C1621 XA.XIR[10].XIC[12].icell.Ien VPWR 0.18829f
C1622 XA.XIR[14].XIC[13].icell.PDM XA.XIR[14].XIC[13].icell.Ien 0.04854f
C1623 XA.XIR[8].XIC[2].icell.Ien Vbias 0.19161f
C1624 XThC.Tn[11] XA.XIR[7].XIC[11].icell.PDM 0.02601f
C1625 XThC.Tn[1] XA.XIR[11].XIC[1].icell.Ien 0.04604f
C1626 XA.XIR[14].XIC[9].icell.PDM XA.XIR[14].XIC[9].icell.Ien 0.04854f
C1627 XThR.Tn[5] XA.XIR[5].XIC[12].icell.Ien 0.14211f
C1628 XThC.XTB6.Y XThC.XTB7.Y 2.05133f
C1629 XA.XIR[0].XIC[11].icell.PDM Vbias 0.03945f
C1630 XA.XIR[5].XIC[6].icell.Ien VPWR 0.18829f
C1631 XThC.XTB7.B a_8739_9569# 0.0168f
C1632 XA.XIR[9].XIC[11].icell.Ien Vbias 0.19161f
C1633 XThC.Tn[14] XA.XIR[7].XIC[14].icell.Ien 0.04604f
C1634 XA.XIR[12].XIC[14].icell.PDM Vbias 0.03928f
C1635 XThC.Tn[8] XA.XIR[13].XIC[8].icell.Ien 0.04604f
C1636 XA.XIR[0].XIC[4].icell.Ien Vbias 0.19213f
C1637 XThR.Tn[12] XA.XIR[12].XIC[11].icell.Ien 0.14211f
C1638 XA.XIR[15].XIC_15.icell.PDM Vbias 0.03927f
C1639 XA.XIR[15].XIC_dummy_right.icell.Ien VPWR 0.3367f
C1640 XThC.Tn[4] XThC.Tn[5] 0.31867f
C1641 XThR.XTB2.Y a_n1049_7787# 0.2342f
C1642 XThC.Tn[0] XA.XIR[14].XIC[0].icell.PDM 0.02601f
C1643 XA.XIR[2].XIC_dummy_left.icell.Iout VPWR 0.10954f
C1644 XA.XIR[0].XIC[12].icell.PDM VPWR 0.01451f
C1645 XA.XIR[7].XIC[7].icell.Ien Vbias 0.19161f
C1646 XA.XIR[13].XIC[14].icell.Ien VPWR 0.18835f
C1647 XThC.Tn[5] XA.XIR[15].XIC[5].icell.Ien 0.04292f
C1648 XThC.Tn[6] XA.XIR[2].XIC[6].icell.PDM 0.02602f
C1649 XThR.Tn[4] XA.XIR[4].XIC[2].icell.Ien 0.14211f
C1650 XA.XIR[0].XIC[10].icell.PDM XA.XIR[0].XIC[10].icell.Ien 0.04854f
C1651 XThR.Tn[10] XA.XIR[11].XIC[8].icell.PDM 0.04035f
C1652 XThC.XTB4.Y XThC.XTB7.Y 0.03475f
C1653 XThR.Tn[0] Iout 1.12768f
C1654 XThR.XTB6.Y XThR.Tn[7] 0.01462f
C1655 XA.XIR[11].XIC[11].icell.PDM XA.XIR[11].XIC[11].icell.Ien 0.04854f
C1656 XThR.Tn[14] XA.XIR[15].XIC[9].icell.PDM 0.04035f
C1657 XThC.Tn[13] XThR.Tn[7] 0.40739f
C1658 XA.XIR[15].XIC_dummy_right.icell.PDM VPWR 0.0824f
C1659 XA.XIR[12].XIC_15.icell.Ien XA.XIR[13].XIC_15.icell.PDM 0.02104f
C1660 XThC.Tn[6] XA.XIR[11].XIC[6].icell.Ien 0.04604f
C1661 XThC.XTB7.B XThC.Tn[11] 0.03651f
C1662 XThC.Tn[10] XA.XIR[6].XIC[10].icell.Ien 0.04604f
C1663 data[2] data[3] 0.04128f
C1664 XA.XIR[2].XIC[0].icell.Ien XA.XIR[3].XIC[0].icell.PDM 0.02104f
C1665 XA.XIR[10].XIC[10].icell.Ien VPWR 0.18829f
C1666 a_6243_9615# Vbias 0.01011f
C1667 XA.XIR[6].XIC[2].icell.PDM Vbias 0.03928f
C1668 XA.XIR[5].XIC[9].icell.Ien XA.XIR[6].XIC[9].icell.PDM 0.02104f
C1669 XA.XIR[5].XIC[9].icell.PDM Vbias 0.03928f
C1670 XThR.Tn[10] XA.XIR[11].XIC[13].icell.PDM 0.0404f
C1671 XThR.Tn[3] XA.XIR[3].XIC[5].icell.Ien 0.14211f
C1672 a_3773_9615# XThC.Tn[2] 0.01043f
C1673 XA.XIR[9].XIC[3].icell.Ien Iout 0.06801f
C1674 XA.XIR[13].XIC[3].icell.PDM Vbias 0.03928f
C1675 XA.XIR[14].XIC[2].icell.PDM XA.XIR[14].XIC[2].icell.Ien 0.04854f
C1676 XThR.XTB3.Y VPWR 1.07975f
C1677 XA.XIR[12].XIC[8].icell.PDM Vbias 0.03928f
C1678 XThR.XTB5.A XThR.XTB6.A 1.80461f
C1679 XThC.Tn[12] XThR.Tn[3] 0.40738f
C1680 XA.XIR[11].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1681 XThC.Tn[0] VPWR 3.67891f
C1682 XA.XIR[6].XIC[3].icell.PDM VPWR 0.01171f
C1683 XThR.Tn[2] XA.XIR[3].XIC[13].icell.PDM 0.0404f
C1684 XA.XIR[14].XIC[0].icell.PDM VPWR 0.01171f
C1685 XA.XIR[5].XIC[10].icell.PDM VPWR 0.01171f
C1686 XA.XIR[5].XIC[12].icell.Ien Iout 0.06801f
C1687 XA.XIR[10].XIC[13].icell.Ien Vbias 0.19161f
C1688 XThC.Tn[8] XThR.Tn[5] 0.40738f
C1689 XA.XIR[3].XIC[4].icell.Ien Vbias 0.19161f
C1690 XA.XIR[13].XIC[4].icell.PDM VPWR 0.01171f
C1691 XA.XIR[13].XIC[12].icell.Ien VPWR 0.18829f
C1692 XThC.Tn[14] XA.XIR[8].XIC[14].icell.Ien 0.04604f
C1693 XThC.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.02601f
C1694 XA.XIR[12].XIC[9].icell.PDM VPWR 0.01171f
C1695 XA.XIR[11].XIC[8].icell.Ien XA.XIR[12].XIC[8].icell.PDM 0.02104f
C1696 XThC.Tn[1] XA.XIR[14].XIC[1].icell.Ien 0.04604f
C1697 XThC.XTB6.A XThC.XTB6.Y 0.10153f
C1698 XThC.XTB2.Y XThC.XTB7.Y 0.0437f
C1699 XA.XIR[9].XIC[2].icell.Ien VPWR 0.18829f
C1700 XA.XIR[3].XIC[4].icell.PDM Vbias 0.03928f
C1701 XA.XIR[4].XIC[13].icell.Ien Vbias 0.19161f
C1702 XA.XIR[12].XIC[13].icell.PDM Vbias 0.03928f
C1703 XA.XIR[12].XIC[7].icell.Ien Iout 0.06801f
C1704 XA.XIR[8].XIC[6].icell.PDM Vbias 0.03928f
C1705 XA.XIR[0].XIC[3].icell.PDM XA.XIR[0].XIC[3].icell.Ien 0.04854f
C1706 XA.XIR[2].XIC[10].icell.PDM Vbias 0.03928f
C1707 XA.XIR[8].XIC[7].icell.Ien Vbias 0.19161f
C1708 XA.XIR[15].XIC[14].icell.PDM Vbias 0.03928f
C1709 XThR.Tn[9] XA.XIR[10].XIC[7].icell.PDM 0.04035f
C1710 XA.XIR[5].XIC[11].icell.Ien VPWR 0.18829f
C1711 XA.XIR[8].XIC[7].icell.PDM VPWR 0.01171f
C1712 XA.XIR[3].XIC[5].icell.PDM VPWR 0.01171f
C1713 XThR.XTB7.B data[6] 0.07481f
C1714 XA.XIR[3].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.PDM 0.02104f
C1715 XA.XIR[0].XIC[9].icell.Ien Vbias 0.19213f
C1716 XA.XIR[2].XIC[11].icell.PDM VPWR 0.01171f
C1717 XThR.Tn[12] XA.XIR[13].XIC[1].icell.PDM 0.04035f
C1718 XA.XIR[5].XIC[2].icell.Ien XA.XIR[6].XIC[2].icell.PDM 0.02104f
C1719 XThC.Tn[14] XThR.Tn[2] 0.40744f
C1720 XA.XIR[1].XIC[0].icell.Ien Iout 0.06795f
C1721 XThC.XTB6.A XThC.XTB4.Y 0.04137f
C1722 XA.XIR[12].XIC[6].icell.Ien VPWR 0.18829f
C1723 XThC.Tn[1] XA.XIR[2].XIC[1].icell.Ien 0.04605f
C1724 XA.XIR[4].XIC[0].icell.Ien Iout 0.06795f
C1725 XA.XIR[10].XIC_15.icell.Ien VPWR 0.26829f
C1726 XThR.Tn[1] Iout 1.12765f
C1727 XThR.XTB6.Y a_n997_1579# 0.07626f
C1728 XA.XIR[7].XIC[12].icell.Ien Vbias 0.19161f
C1729 XThC.Tn[6] XA.XIR[14].XIC[6].icell.Ien 0.04604f
C1730 XA.XIR[2].XIC[10].icell.Ien XA.XIR[3].XIC[10].icell.PDM 0.02104f
C1731 XThR.Tn[4] XA.XIR[4].XIC[7].icell.Ien 0.14211f
C1732 XThR.Tn[12] Iout 1.12762f
C1733 XA.XIR[7].XIC[11].icell.Ien XA.XIR[8].XIC[11].icell.PDM 0.02104f
C1734 XA.XIR[11].XIC_dummy_right.icell.PDM XA.XIR[11].XIC_dummy_right.icell.Ien 0.04854f
C1735 XA.XIR[10].XIC[11].icell.Ien Vbias 0.19161f
C1736 XA.XIR[3].XIC[1].icell.Ien Vbias 0.19161f
C1737 XA.XIR[13].XIC[10].icell.Ien VPWR 0.18829f
C1738 XThR.Tn[10] XA.XIR[11].XIC[12].icell.PDM 0.04035f
C1739 XThR.Tn[0] XA.XIR[1].XIC[9].icell.PDM 0.04035f
C1740 XA.XIR[1].XIC[13].icell.Ien XA.XIR[2].XIC[13].icell.PDM 0.02104f
C1741 XA.XIR[15].XIC[2].icell.Ien Iout 0.07192f
C1742 XThR.Tn[11] XA.XIR[12].XIC_dummy_left.icell.Iout 0.02485f
C1743 XThC.Tn[10] XThR.Tn[6] 0.40738f
C1744 XThR.Tn[1] XA.XIR[2].XIC[8].icell.PDM 0.04035f
C1745 XA.XIR[4].XIC[5].icell.Ien Iout 0.06801f
C1746 XA.XIR[12].XIC[12].icell.Ien XA.XIR[13].XIC[12].icell.PDM 0.02104f
C1747 XThC.Tn[12] XThR.Tn[11] 0.40738f
C1748 XA.XIR[10].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1749 XThR.Tn[7] XA.XIR[8].XIC[13].icell.PDM 0.0404f
C1750 XA.XIR[6].XIC[11].icell.PDM XA.XIR[6].XIC[11].icell.Ien 0.04854f
C1751 XA.XIR[7].XIC[10].icell.PDM Vbias 0.03928f
C1752 XThC.Tn[2] XThR.Tn[7] 0.40738f
C1753 XThR.Tn[13] XA.XIR[14].XIC[14].icell.PDM 0.04056f
C1754 XA.XIR[15].XIC[8].icell.PDM Vbias 0.03928f
C1755 XThR.Tn[12] XA.XIR[12].XIC[5].icell.Ien 0.14211f
C1756 XThC.Tn[8] Iout 0.22393f
C1757 XA.XIR[14].XIC_dummy_left.icell.PDM VPWR 0.08221f
C1758 XA.XIR[10].XIC[4].icell.Ien XA.XIR[11].XIC[4].icell.PDM 0.02104f
C1759 XThR.Tn[3] XA.XIR[3].XIC[10].icell.Ien 0.14211f
C1760 XA.XIR[9].XIC[10].icell.Ien XA.XIR[10].XIC[10].icell.PDM 0.02104f
C1761 XA.XIR[10].XIC[5].icell.PDM XA.XIR[10].XIC[5].icell.Ien 0.04854f
C1762 XA.XIR[9].XIC[8].icell.Ien Iout 0.06801f
C1763 XThC.Tn[2] XA.XIR[4].XIC[2].icell.Ien 0.04604f
C1764 XThC.XTB6.Y XThC.Tn[8] 0.02463f
C1765 XThR.Tn[3] XA.XIR[4].XIC[14].icell.PDM 0.04056f
C1766 XA.XIR[9].XIC[6].icell.PDM Vbias 0.03928f
C1767 XA.XIR[6].XIC_dummy_left.icell.PDM XA.XIR[6].XIC_dummy_left.icell.Ien 0.04854f
C1768 XA.XIR[13].XIC[13].icell.Ien Vbias 0.19161f
C1769 XThR.XTB7.Y a_n1319_5317# 0.01283f
C1770 XA.XIR[7].XIC[11].icell.PDM VPWR 0.01171f
C1771 XThR.Tn[2] XA.XIR[2].XIC[5].icell.Ien 0.14211f
C1772 XA.XIR[12].XIC[12].icell.PDM Vbias 0.03928f
C1773 XThC.Tn[1] XA.XIR[6].XIC[1].icell.PDM 0.02601f
C1774 XThC.XTB2.Y XThC.XTB6.A 0.18237f
C1775 XA.XIR[4].XIC[4].icell.Ien VPWR 0.18829f
C1776 XA.XIR[15].XIC[9].icell.PDM VPWR 0.01512f
C1777 XThC.Tn[8] XA.XIR[2].XIC[8].icell.PDM 0.02602f
C1778 XA.XIR[15].XIC[13].icell.PDM Vbias 0.03928f
C1779 XA.XIR[7].XIC[4].icell.Ien Iout 0.06801f
C1780 XA.XIR[3].XIC[9].icell.Ien Vbias 0.19161f
C1781 XA.XIR[1].XIC[11].icell.PDM Vbias 0.03928f
C1782 XThC.Tn[1] XThR.Tn[3] 0.40738f
C1783 XA.XIR[9].XIC[7].icell.PDM VPWR 0.01171f
C1784 XThC.Tn[10] XThR.Tn[4] 0.40738f
C1785 XThC.XTBN.Y XThC.Tn[13] 0.41509f
C1786 XA.XIR[2].XIC[2].icell.Ien Vbias 0.19161f
C1787 XA.XIR[4].XIC[11].icell.PDM Vbias 0.03928f
C1788 XA.XIR[9].XIC[14].icell.PDM XA.XIR[9].XIC[14].icell.Ien 0.04854f
C1789 XA.XIR[7].XIC[12].icell.PDM XA.XIR[7].XIC[12].icell.Ien 0.04854f
C1790 XThC.XTB6.A data[1] 0.37233f
C1791 XA.XIR[9].XIC[7].icell.Ien VPWR 0.18829f
C1792 XA.XIR[1].XIC[4].icell.Ien Vbias 0.19173f
C1793 XThC.XTB4.Y XThC.Tn[8] 0.01307f
C1794 XA.XIR[2].XIC[3].icell.Ien XA.XIR[3].XIC[3].icell.PDM 0.02104f
C1795 XA.XIR[4].XIC[13].icell.PDM XA.XIR[4].XIC[13].icell.Ien 0.04854f
C1796 XA.XIR[7].XIC[4].icell.Ien XA.XIR[8].XIC[4].icell.PDM 0.02104f
C1797 XThR.Tn[9] XA.XIR[9].XIC[3].icell.Ien 0.14211f
C1798 XA.XIR[10].XIC[0].icell.Ien XA.XIR[11].XIC[0].icell.PDM 0.02104f
C1799 XThC.Tn[14] XThR.Tn[10] 0.40742f
C1800 XThC.Tn[4] XThR.Tn[0] 0.40763f
C1801 XThC.Tn[10] XA.XIR[10].XIC[10].icell.PDM 0.02601f
C1802 XThR.Tn[4] XA.XIR[5].XIC[6].icell.PDM 0.04035f
C1803 XThC.Tn[6] XThR.Tn[5] 0.40738f
C1804 XA.XIR[8].XIC[12].icell.Ien Vbias 0.19161f
C1805 XA.XIR[1].XIC[12].icell.PDM VPWR 0.01171f
C1806 XA.XIR[1].XIC[6].icell.Ien XA.XIR[2].XIC[6].icell.PDM 0.02104f
C1807 XA.XIR[10].XIC[1].icell.PDM XA.XIR[10].XIC[1].icell.Ien 0.04854f
C1808 XThC.Tn[7] XA.XIR[0].XIC[7].icell.Ien 0.04658f
C1809 XThC.Tn[11] XThC.Tn[12] 0.12311f
C1810 XA.XIR[8].XIC[11].icell.PDM XA.XIR[8].XIC[11].icell.Ien 0.04854f
C1811 XA.XIR[7].XIC[3].icell.Ien VPWR 0.18829f
C1812 XA.XIR[4].XIC[12].icell.PDM VPWR 0.01171f
C1813 XThR.Tn[13] XA.XIR[14].XIC[8].icell.PDM 0.04035f
C1814 XA.XIR[7].XIC_dummy_right.icell.PDM XA.XIR[7].XIC_dummy_right.icell.Ien 0.04854f
C1815 XThC.XTB7.B VPWR 1.33508f
C1816 XA.XIR[0].XIC[10].icell.Ien XA.XIR[1].XIC[10].icell.PDM 0.02104f
C1817 XA.XIR[14].XIC[11].icell.PDM XA.XIR[14].XIC[11].icell.Ien 0.04854f
C1818 XA.XIR[13].XIC_15.icell.Ien VPWR 0.26829f
C1819 XA.XIR[6].XIC[4].icell.PDM XA.XIR[6].XIC[4].icell.Ien 0.04854f
C1820 XA.XIR[15].XIC[3].icell.PDM XA.XIR[15].XIC[3].icell.Ien 0.04854f
C1821 XA.XIR[0].XIC[14].icell.Ien Vbias 0.19213f
C1822 XThR.Tn[8] XA.XIR[9].XIC[11].icell.PDM 0.04035f
C1823 XThR.Tn[10] XA.XIR[11].XIC[11].icell.PDM 0.04035f
C1824 XThC.XTBN.A XThC.XTB5.Y 0.10854f
C1825 XThC.Tn[0] XA.XIR[0].XIC[0].icell.Ien 0.04657f
C1826 XA.XIR[13].XIC[11].icell.Ien Vbias 0.19161f
C1827 XA.XIR[9].XIC[3].icell.Ien XA.XIR[10].XIC[3].icell.PDM 0.02104f
C1828 XThR.Tn[7] XA.XIR[7].XIC[0].icell.Ien 0.14211f
C1829 XThR.XTBN.A XThR.Tn[8] 0.1369f
C1830 XThC.Tn[8] XA.XIR[7].XIC[8].icell.PDM 0.02601f
C1831 XThR.Tn[5] XA.XIR[6].XIC[8].icell.PDM 0.04035f
C1832 XThC.Tn[3] XThR.Tn[2] 0.40741f
C1833 XThR.Tn[4] XA.XIR[4].XIC[12].icell.Ien 0.14211f
C1834 XThR.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.0404f
C1835 XThC.XTB7.Y a_6243_9615# 0.27822f
C1836 XA.XIR[11].XIC[1].icell.PDM Vbias 0.03928f
C1837 XA.XIR[0].XIC_15.icell.PUM VPWR 0.01577f
C1838 XThR.Tn[0] XA.XIR[0].XIC[4].icell.Ien 0.14211f
C1839 XThR.Tn[2] XA.XIR[3].XIC[0].icell.PDM 0.0404f
C1840 XA.XIR[13].XIC_dummy_right.icell.Iout VPWR 0.11567f
C1841 XThR.Tn[10] XA.XIR[10].XIC[3].icell.Ien 0.14211f
C1842 XThC.Tn[12] XThR.Tn[14] 0.40738f
C1843 XA.XIR[10].XIC[5].icell.PDM Vbias 0.03928f
C1844 XA.XIR[15].XIC[7].icell.Ien Iout 0.07192f
C1845 XThC.Tn[14] XA.XIR[8].XIC[14].icell.PDM 0.02601f
C1846 XThC.XTBN.A XThC.XTBN.Y 0.77125f
C1847 XThR.Tn[6] XA.XIR[7].XIC[7].icell.PDM 0.04035f
C1848 XThC.Tn[12] XA.XIR[10].XIC[12].icell.Ien 0.04604f
C1849 XA.XIR[6].XIC[4].icell.Ien Vbias 0.19161f
C1850 XA.XIR[4].XIC[10].icell.Ien Iout 0.06801f
C1851 XThR.Tn[7] XA.XIR[7].XIC[5].icell.Ien 0.14211f
C1852 XA.XIR[6].XIC[13].icell.Ien XA.XIR[7].XIC[13].icell.PDM 0.02104f
C1853 XA.XIR[15].XIC[1].icell.Ien VPWR 0.31713f
C1854 XA.XIR[5].XIC_dummy_left.icell.Iout VPWR 0.11011f
C1855 XA.XIR[0].XIC[1].icell.Ien Iout 0.0675f
C1856 XThC.Tn[10] XA.XIR[11].XIC[10].icell.Ien 0.04604f
C1857 XA.XIR[7].XIC[5].icell.PDM XA.XIR[7].XIC[5].icell.Ien 0.04854f
C1858 XA.XIR[9].XIC[7].icell.PDM XA.XIR[9].XIC[7].icell.Ien 0.04854f
C1859 XA.XIR[12].XIC[11].icell.PDM Vbias 0.03928f
C1860 XA.XIR[11].XIC[2].icell.PDM VPWR 0.01171f
C1861 XA.XIR[8].XIC[4].icell.Ien Iout 0.06801f
C1862 XA.XIR[4].XIC[6].icell.PDM XA.XIR[4].XIC[6].icell.Ien 0.04854f
C1863 XA.XIR[10].XIC[6].icell.PDM VPWR 0.01171f
C1864 XA.XIR[15].XIC[12].icell.PDM Vbias 0.03928f
C1865 XThC.Tn[3] XA.XIR[2].XIC[3].icell.PDM 0.02602f
C1866 XThR.Tn[3] XA.XIR[3].XIC_15.icell.Ien 0.13564f
C1867 XThC.XTBN.A XThC.Tn[10] 0.12208f
C1868 XA.XIR[14].XIC[8].icell.Ien XA.XIR[15].XIC[8].icell.PDM 0.02104f
C1869 XA.XIR[9].XIC[13].icell.Ien Iout 0.06801f
C1870 XThC.Tn[6] XA.XIR[12].XIC[6].icell.PDM 0.02601f
C1871 XThC.Tn[1] XThR.Tn[11] 0.40738f
C1872 XA.XIR[15].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.Iout 0.06446f
C1873 XA.XIR[8].XIC[4].icell.PDM XA.XIR[8].XIC[4].icell.Ien 0.04854f
C1874 XA.XIR[15].XIC[6].icell.Ien VPWR 0.31713f
C1875 XA.XIR[0].XIC[13].icell.PDM Vbias 0.03945f
C1876 XThC.Tn[7] XA.XIR[3].XIC[7].icell.Ien 0.04604f
C1877 XA.XIR[11].XIC[3].icell.Ien Vbias 0.19161f
C1878 XA.XIR[0].XIC[6].icell.Ien Iout 0.0675f
C1879 XThR.Tn[2] XA.XIR[2].XIC[10].icell.Ien 0.14211f
C1880 XThC.Tn[12] XA.XIR[0].XIC[12].icell.PDM 0.0279f
C1881 XA.XIR[0].XIC[3].icell.Ien XA.XIR[1].XIC[3].icell.PDM 0.02104f
C1882 XA.XIR[4].XIC[9].icell.Ien VPWR 0.18829f
C1883 XThC.XTB3.Y XThC.XTB5.Y 0.04438f
C1884 XThC.Tn[14] XA.XIR[2].XIC[14].icell.Ien 0.04605f
C1885 XA.XIR[10].XIC[5].icell.Ien Vbias 0.19161f
C1886 XA.XIR[0].XIC[0].icell.Ien VPWR 0.18776f
C1887 XThC.Tn[6] Iout 0.22423f
C1888 XThC.Tn[0] XA.XIR[10].XIC[0].icell.Ien 0.04604f
C1889 XA.XIR[8].XIC[11].icell.Ien XA.XIR[9].XIC[11].icell.PDM 0.02104f
C1890 XA.XIR[8].XIC[3].icell.Ien VPWR 0.18829f
C1891 XA.XIR[7].XIC[9].icell.Ien Iout 0.06801f
C1892 XA.XIR[8].XIC_dummy_left.icell.PDM XA.XIR[8].XIC_dummy_left.icell.Ien 0.04854f
C1893 XThC.XTB6.Y XThC.Tn[6] 0.01038f
C1894 XA.XIR[10].XIC[14].icell.PDM XA.XIR[10].XIC[14].icell.Ien 0.04854f
C1895 XA.XIR[3].XIC[14].icell.Ien Vbias 0.19161f
C1896 XThC.Tn[5] XA.XIR[10].XIC[5].icell.PDM 0.02601f
C1897 XA.XIR[3].XIC[10].icell.Ien XA.XIR[4].XIC[10].icell.PDM 0.02104f
C1898 XThC.Tn[14] XThR.Tn[13] 0.40742f
C1899 XThC.Tn[10] XA.XIR[13].XIC[10].icell.PDM 0.02601f
C1900 XA.XIR[0].XIC[14].icell.PDM VPWR 0.01141f
C1901 XA.XIR[3].XIC[12].icell.PDM XA.XIR[3].XIC[12].icell.Ien 0.04854f
C1902 XThC.Tn[4] XThR.Tn[1] 0.40744f
C1903 XA.XIR[2].XIC[7].icell.Ien Vbias 0.19161f
C1904 XThC.Tn[8] XThR.Tn[9] 0.40738f
C1905 XA.XIR[9].XIC[12].icell.Ien VPWR 0.18829f
C1906 XThR.XTB6.Y XThR.Tn[8] 0.02461f
C1907 XThR.XTBN.A data[4] 0.02581f
C1908 XA.XIR[1].XIC[9].icell.Ien Vbias 0.19173f
C1909 XThC.Tn[4] XThR.Tn[12] 0.40738f
C1910 XThC.Tn[13] XThR.Tn[8] 0.40739f
C1911 XA.XIR[2].XIC[0].icell.Ien Iout 0.06795f
C1912 XThR.Tn[9] XA.XIR[9].XIC[8].icell.Ien 0.14211f
C1913 XA.XIR[0].XIC[5].icell.Ien VPWR 0.18797f
C1914 XThC.XTB3.Y XThC.XTBN.Y 0.17246f
C1915 XThR.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.04035f
C1916 XThR.XTBN.A a_n997_3755# 0.01939f
C1917 XThR.XTB2.Y XThR.XTBN.A 0.04716f
C1918 XA.XIR[3].XIC_15.icell.PUM VPWR 0.01655f
C1919 XThC.XTBN.Y XThC.Tn[2] 0.49723f
C1920 XA.XIR[10].XIC[1].icell.Ien Iout 0.06801f
C1921 XThR.XTB7.A XThR.Tn[5] 0.02751f
C1922 XA.XIR[7].XIC[8].icell.Ien VPWR 0.18829f
C1923 XA.XIR[10].XIC_dummy_right.icell.Ien VPWR 0.35722f
C1924 XA.XIR[3].XIC_dummy_right.icell.PDM XA.XIR[3].XIC_dummy_right.icell.Ien 0.04854f
C1925 XA.XIR[6].XIC[6].icell.Ien XA.XIR[7].XIC[6].icell.PDM 0.02104f
C1926 XA.XIR[14].XIC_dummy_right.icell.PDM XA.XIR[14].XIC_dummy_right.icell.Ien 0.04854f
C1927 XThC.Tn[3] XA.XIR[7].XIC[3].icell.PDM 0.02601f
C1928 XThR.Tn[7] XA.XIR[8].XIC[0].icell.PDM 0.0404f
C1929 XThR.Tn[13] XA.XIR[14].XIC[12].icell.PDM 0.04035f
C1930 XThC.Tn[3] XThR.Tn[10] 0.40738f
C1931 XThC.Tn[14] XA.XIR[9].XIC[14].icell.PDM 0.02601f
C1932 XThC.XTB3.Y XThC.Tn[10] 0.29566f
C1933 XA.XIR[6].XIC[4].icell.PDM Vbias 0.03928f
C1934 XThC.Tn[5] XA.XIR[10].XIC[5].icell.Ien 0.04604f
C1935 XA.XIR[14].XIC[1].icell.PDM Vbias 0.03928f
C1936 XA.XIR[5].XIC[11].icell.PDM Vbias 0.03928f
C1937 XThR.XTB7.A data[5] 0.06538f
C1938 a_n1049_8581# VPWR 0.72063f
C1939 XA.XIR[13].XIC[5].icell.PDM Vbias 0.03928f
C1940 XA.XIR[4].XIC[13].icell.Ien XA.XIR[5].XIC[13].icell.PDM 0.02104f
C1941 XThR.Tn[11] XA.XIR[11].XIC[4].icell.Ien 0.14211f
C1942 XThC.XTB1.Y XThC.XTB5.Y 0.05054f
C1943 XThR.Tn[3] XA.XIR[4].XIC[1].icell.PDM 0.04035f
C1944 XThC.Tn[12] XA.XIR[13].XIC[12].icell.Ien 0.04604f
C1945 XA.XIR[11].XIC[13].icell.Ien Iout 0.06801f
C1946 XA.XIR[12].XIC[10].icell.PDM Vbias 0.03928f
C1947 XA.XIR[13].XIC[4].icell.Ien XA.XIR[14].XIC[4].icell.PDM 0.02104f
C1948 XA.XIR[10].XIC[0].icell.Ien VPWR 0.18829f
C1949 XA.XIR[10].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.Iout 0.06446f
C1950 XThC.Tn[8] XA.XIR[4].XIC[8].icell.Ien 0.04604f
C1951 XThR.XTB1.Y XThR.XTB5.Y 0.05054f
C1952 XA.XIR[3].XIC[6].icell.Ien Iout 0.06801f
C1953 XThR.Tn[0] XA.XIR[0].XIC[9].icell.Ien 0.14211f
C1954 XA.XIR[13].XIC[5].icell.PDM XA.XIR[13].XIC[5].icell.Ien 0.04854f
C1955 XA.XIR[6].XIC[5].icell.PDM VPWR 0.01171f
C1956 XThC.Tn[10] XA.XIR[14].XIC[10].icell.Ien 0.04604f
C1957 XThR.Tn[10] XA.XIR[10].XIC[8].icell.Ien 0.14211f
C1958 XA.XIR[15].XIC[11].icell.PDM Vbias 0.03928f
C1959 XThR.Tn[6] XA.XIR[6].XIC[3].icell.Ien 0.14211f
C1960 XA.XIR[5].XIC[12].icell.PDM VPWR 0.01171f
C1961 XA.XIR[14].XIC[2].icell.PDM VPWR 0.01171f
C1962 XA.XIR[12].XIC[6].icell.Ien XA.XIR[13].XIC[6].icell.PDM 0.02104f
C1963 XA.XIR[8].XIC[4].icell.Ien XA.XIR[9].XIC[4].icell.PDM 0.02104f
C1964 XThC.Tn[4] XA.XIR[7].XIC[4].icell.Ien 0.04604f
C1965 XA.XIR[13].XIC[6].icell.PDM VPWR 0.01171f
C1966 XA.XIR[3].XIC[3].icell.Ien XA.XIR[4].XIC[3].icell.PDM 0.02104f
C1967 XThR.Tn[7] XA.XIR[7].XIC[10].icell.Ien 0.14211f
C1968 XA.XIR[4].XIC_15.icell.Ien Iout 0.0694f
C1969 XA.XIR[6].XIC[9].icell.Ien Vbias 0.19161f
C1970 XThC.Tn[1] XA.XIR[5].XIC[1].icell.Ien 0.04604f
C1971 XA.XIR[3].XIC[5].icell.PDM XA.XIR[3].XIC[5].icell.Ien 0.04854f
C1972 XThC.XTB1.Y XThC.XTBN.Y 0.1979f
C1973 XThC.Tn[6] XA.XIR[15].XIC[6].icell.PDM 0.02601f
C1974 XThC.Tn[1] XThR.Tn[14] 0.40738f
C1975 XA.XIR[8].XIC[9].icell.Ien Iout 0.06801f
C1976 XA.XIR[12].XIC_dummy_left.icell.Ien XThR.Tn[12] 0.01244f
C1977 XA.XIR[8].XIC_dummy_left.icell.Ien XA.XIR[9].XIC_dummy_left.icell.PDM 0.02104f
C1978 XA.XIR[8].XIC[8].icell.PDM Vbias 0.03928f
C1979 XA.XIR[3].XIC[6].icell.PDM Vbias 0.03928f
C1980 XThR.XTB2.Y a_n1049_7493# 0.02133f
C1981 XA.XIR[14].XIC[3].icell.Ien Vbias 0.19161f
C1982 XThC.Tn[7] XA.XIR[0].XIC[7].icell.PDM 0.02803f
C1983 XA.XIR[2].XIC[12].icell.PDM Vbias 0.03928f
C1984 XA.XIR[13].XIC[5].icell.Ien Vbias 0.19161f
C1985 XA.XIR[12].XIC[10].icell.Ien XA.XIR[13].XIC[10].icell.PDM 0.02104f
C1986 XThR.Tn[6] XA.XIR[7].XIC_dummy_left.icell.Iout 0.01728f
C1987 XA.XIR[3].XIC[5].icell.Ien VPWR 0.18829f
C1988 XA.XIR[12].XIC_dummy_left.icell.Iout VPWR 0.10997f
C1989 XThR.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.04035f
C1990 XThC.Tn[0] XA.XIR[13].XIC[0].icell.Ien 0.04604f
C1991 XThR.XTB2.Y XThR.XTB6.Y 0.04959f
C1992 XThC.Tn[5] XA.XIR[13].XIC[5].icell.PDM 0.02601f
C1993 XA.XIR[11].XIC[8].icell.Ien Vbias 0.19161f
C1994 XThC.Tn[6] XA.XIR[9].XIC[6].icell.Ien 0.04604f
C1995 XA.XIR[0].XIC[11].icell.Ien Iout 0.0675f
C1996 XThR.Tn[2] XA.XIR[2].XIC_15.icell.Ien 0.13564f
C1997 XA.XIR[4].XIC_dummy_right.icell.Iout Iout 0.01732f
C1998 XA.XIR[13].XIC[0].icell.Ien XA.XIR[14].XIC[0].icell.PDM 0.02104f
C1999 XThC.Tn[12] VPWR 4.5561f
C2000 XThC.Tn[13] XA.XIR[0].XIC[13].icell.Ien 0.04662f
C2001 XThR.Tn[14] XA.XIR[15].XIC_dummy_left.icell.Iout 0.0203f
C2002 XA.XIR[3].XIC[7].icell.PDM VPWR 0.01171f
C2003 XA.XIR[4].XIC[14].icell.Ien VPWR 0.18835f
C2004 XA.XIR[8].XIC[9].icell.PDM VPWR 0.01171f
C2005 XA.XIR[13].XIC[1].icell.PDM XA.XIR[13].XIC[1].icell.Ien 0.04854f
C2006 XThC.XTBN.A a_7651_9569# 0.02087f
C2007 XA.XIR[2].XIC[13].icell.PDM VPWR 0.01171f
C2008 XThR.Tn[12] XA.XIR[13].XIC[3].icell.PDM 0.04035f
C2009 XThC.Tn[7] XA.XIR[1].XIC[7].icell.Ien 0.04606f
C2010 XA.XIR[7].XIC[14].icell.Ien Iout 0.06801f
C2011 XA.XIR[8].XIC[8].icell.Ien VPWR 0.18829f
C2012 XThR.XTB6.Y a_n1049_5611# 0.26831f
C2013 XA.XIR[11].XIC[11].icell.Ien Iout 0.06801f
C2014 XA.XIR[10].XIC_15.icell.PDM XA.XIR[10].XIC_15.icell.Ien 0.04854f
C2015 XA.XIR[10].XIC_15.icell.PDM VPWR 0.07527f
C2016 XA.XIR[1].XIC[10].icell.PDM XA.XIR[1].XIC[10].icell.Ien 0.04854f
C2017 XA.XIR[2].XIC[12].icell.Ien Vbias 0.19161f
C2018 XA.XIR[4].XIC[6].icell.Ien XA.XIR[5].XIC[6].icell.PDM 0.02104f
C2019 XA.XIR[13].XIC[1].icell.Ien Iout 0.06801f
C2020 XA.XIR[0].XIC_dummy_left.icell.Ien VPWR 0.38924f
C2021 XThR.Tn[13] XA.XIR[14].XIC[11].icell.PDM 0.04035f
C2022 XA.XIR[1].XIC[14].icell.Ien Vbias 0.19173f
C2023 XThC.Tn[5] Vbias 0.82298f
C2024 XA.XIR[13].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2025 XThR.Tn[9] XA.XIR[9].XIC[13].icell.Ien 0.14211f
C2026 XA.XIR[0].XIC[10].icell.Ien VPWR 0.18776f
C2027 XA.XIR[2].XIC[12].icell.PDM XA.XIR[2].XIC[12].icell.Ien 0.04854f
C2028 XThC.Tn[3] XThR.Tn[13] 0.40738f
C2029 XThR.Tn[0] XA.XIR[1].XIC[11].icell.PDM 0.04035f
C2030 XA.XIR[12].XIC[1].icell.Ien Vbias 0.19161f
C2031 XThC.Tn[5] XA.XIR[13].XIC[5].icell.Ien 0.04604f
C2032 XThR.Tn[1] XA.XIR[2].XIC[10].icell.PDM 0.04035f
C2033 XA.XIR[7].XIC[13].icell.Ien VPWR 0.18829f
C2034 XThC.Tn[6] XThR.Tn[9] 0.40738f
C2035 XThC.Tn[8] XA.XIR[12].XIC[8].icell.PDM 0.02601f
C2036 XThC.Tn[2] XThR.Tn[8] 0.40738f
C2037 XThR.Tn[13] XA.XIR[13].XIC[3].icell.Ien 0.14211f
C2038 XA.XIR[1].XIC_15.icell.PUM VPWR 0.01655f
C2039 XA.XIR[5].XIC[2].icell.Ien Vbias 0.19161f
C2040 XA.XIR[7].XIC[12].icell.PDM Vbias 0.03928f
C2041 XThC.Tn[4] XA.XIR[8].XIC[4].icell.Ien 0.04604f
C2042 XA.XIR[11].XIC[3].icell.PDM XA.XIR[11].XIC[3].icell.Ien 0.04854f
C2043 XA.XIR[14].XIC[13].icell.Ien Iout 0.06801f
C2044 XA.XIR[15].XIC[10].icell.PDM Vbias 0.03928f
C2045 XA.XIR[2].XIC_dummy_right.icell.PDM XA.XIR[2].XIC_dummy_right.icell.Ien 0.04854f
C2046 XA.XIR[13].XIC[0].icell.Ien VPWR 0.18829f
C2047 XThC.XTBN.Y a_2979_9615# 0.0607f
C2048 XA.XIR[5].XIC_15.icell.PDM XA.XIR[5].XIC_15.icell.Ien 0.04854f
C2049 XA.XIR[1].XIC[1].icell.Ien Iout 0.06801f
C2050 XThR.XTB7.Y XThR.XTBN.A 1.11559f
C2051 XA.XIR[10].XIC[2].icell.Ien Iout 0.06801f
C2052 XA.XIR[9].XIC[8].icell.PDM Vbias 0.03928f
C2053 a_10051_9569# Vbias 0.0105f
C2054 XThR.Tn[11] XA.XIR[11].XIC[9].icell.Ien 0.14211f
C2055 XThR.XTB5.A XThR.XTB7.A 0.07862f
C2056 XA.XIR[0].XIC[0].icell.PDM Vbias 0.03934f
C2057 XA.XIR[7].XIC[13].icell.PDM VPWR 0.01171f
C2058 XThR.XTB7.Y XThR.Tn[6] 0.21438f
C2059 a_9827_9569# XThC.Tn[12] 0.20217f
C2060 XThC.Tn[0] XThC.Tn[1] 0.88262f
C2061 XThC.Tn[7] XA.XIR[6].XIC[7].icell.Ien 0.04604f
C2062 XA.XIR[3].XIC[11].icell.Ien Iout 0.06801f
C2063 XThR.Tn[0] XA.XIR[0].XIC[14].icell.Ien 0.144f
C2064 XThC.Tn[13] XA.XIR[3].XIC[13].icell.Ien 0.04604f
C2065 XThR.Tn[6] XA.XIR[6].XIC[8].icell.Ien 0.14211f
C2066 XA.XIR[2].XIC[4].icell.Ien Iout 0.06801f
C2067 a_n1049_7787# VPWR 0.72195f
C2068 XA.XIR[1].XIC[13].icell.PDM Vbias 0.03928f
C2069 XA.XIR[6].XIC[14].icell.Ien Vbias 0.19161f
C2070 XA.XIR[1].XIC[6].icell.Ien Iout 0.06801f
C2071 XThR.Tn[7] XA.XIR[7].XIC_15.icell.Ien 0.13564f
C2072 XA.XIR[9].XIC[9].icell.PDM VPWR 0.01171f
C2073 XThC.Tn[12] XA.XIR[1].XIC[12].icell.PDM 0.02602f
C2074 XA.XIR[0].XIC[1].icell.PDM VPWR 0.01132f
C2075 XA.XIR[1].XIC[3].icell.PDM XA.XIR[1].XIC[3].icell.Ien 0.04854f
C2076 XA.XIR[4].XIC[13].icell.PDM Vbias 0.03928f
C2077 XA.XIR[9].XIC[0].icell.PDM XA.XIR[9].XIC[0].icell.Ien 0.04854f
C2078 XThC.Tn[0] XA.XIR[6].XIC[0].icell.Ien 0.04604f
C2079 XA.XIR[8].XIC[14].icell.Ien Iout 0.06801f
C2080 XThC.Tn[12] XA.XIR[4].XIC[12].icell.PDM 0.02601f
C2081 XThC.Tn[14] XThR.Tn[7] 0.40742f
C2082 XA.XIR[13].XIC[14].icell.PDM XA.XIR[13].XIC[14].icell.Ien 0.04854f
C2083 XThC.XTB5.A a_7331_10587# 0.01243f
C2084 XA.XIR[14].XIC[8].icell.Ien Vbias 0.19161f
C2085 XA.XIR[2].XIC[5].icell.PDM XA.XIR[2].XIC[5].icell.Ien 0.04854f
C2086 XThR.XTBN.Y XThR.Tn[5] 0.59911f
C2087 XThR.Tn[4] XA.XIR[5].XIC[8].icell.PDM 0.04035f
C2088 XA.XIR[3].XIC[10].icell.Ien VPWR 0.18829f
C2089 XA.XIR[1].XIC[14].icell.PDM VPWR 0.0118f
C2090 XA.XIR[10].XIC[14].icell.PDM VPWR 0.0118f
C2091 XA.XIR[11].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.Iout 0.06446f
C2092 XA.XIR[6].XIC_15.icell.PUM VPWR 0.01655f
C2093 XThR.Tn[3] XThR.Tn[4] 0.1175f
C2094 XThR.XTBN.A a_n997_2667# 0.01679f
C2095 XThC.Tn[11] XA.XIR[8].XIC[11].icell.PDM 0.02601f
C2096 XA.XIR[2].XIC[3].icell.Ien VPWR 0.18829f
C2097 XA.XIR[4].XIC[14].icell.PDM VPWR 0.0118f
C2098 XA.XIR[0].XIC_dummy_left.icell.PUM VPWR 0.015f
C2099 XThR.Tn[13] XA.XIR[14].XIC[10].icell.PDM 0.04035f
C2100 XA.XIR[14].XIC[11].icell.Ien Iout 0.06801f
C2101 XA.XIR[13].XIC_15.icell.PDM VPWR 0.07527f
C2102 XA.XIR[1].XIC[5].icell.Ien VPWR 0.18829f
C2103 XA.XIR[6].XIC[1].icell.Ien Iout 0.06801f
C2104 XThR.Tn[8] XA.XIR[9].XIC[13].icell.PDM 0.0404f
C2105 XA.XIR[8].XIC[13].icell.Ien VPWR 0.18829f
C2106 XA.XIR[5].XIC[8].icell.PDM XA.XIR[5].XIC[8].icell.Ien 0.04854f
C2107 XThC.Tn[13] XThR.Tn[3] 0.40739f
C2108 XThR.Tn[2] Iout 1.12764f
C2109 XThC.XTB7.A XThC.XTBN.A 0.197f
C2110 XThC.Tn[0] XA.XIR[2].XIC[0].icell.PDM 0.02602f
C2111 XThC.XTB1.Y a_7651_9569# 0.06353f
C2112 XThC.Tn[1] VPWR 3.60376f
C2113 XThR.XTB6.Y XThR.XTB7.Y 2.05133f
C2114 XThC.Tn[3] XA.XIR[12].XIC[3].icell.PDM 0.02601f
C2115 XThR.Tn[5] XA.XIR[6].XIC[10].icell.PDM 0.04035f
C2116 XA.XIR[10].XIC[12].icell.PDM XA.XIR[10].XIC[12].icell.Ien 0.04854f
C2117 XThR.XTBN.A XThR.Tn[11] 0.11968f
C2118 XThC.Tn[8] XA.XIR[15].XIC[8].icell.PDM 0.02601f
C2119 XThC.Tn[9] XThR.Tn[5] 0.40738f
C2120 XA.XIR[11].XIC[3].icell.PDM Vbias 0.03928f
C2121 XA.XIR[0].XIC_15.icell.Ien VPWR 0.26622f
C2122 XThC.Tn[14] XA.XIR[5].XIC[14].icell.Ien 0.04604f
C2123 XA.XIR[6].XIC[6].icell.Ien Iout 0.06801f
C2124 XThR.Tn[2] XA.XIR[3].XIC[2].icell.PDM 0.04035f
C2125 XThC.Tn[9] XA.XIR[0].XIC[9].icell.PDM 0.02801f
C2126 XThR.Tn[14] XA.XIR[14].XIC[4].icell.Ien 0.14211f
C2127 XA.XIR[10].XIC[7].icell.PDM Vbias 0.03928f
C2128 XThR.Tn[11] XA.XIR[11].XIC[14].icell.Ien 0.144f
C2129 XThR.Tn[1] XA.XIR[1].XIC[4].icell.Ien 0.14211f
C2130 XThC.Tn[14] XA.XIR[3].XIC[14].icell.PDM 0.02601f
C2131 XA.XIR[4].XIC_dummy_right.icell.Iout XA.XIR[5].XIC_dummy_right.icell.Iout 0.04047f
C2132 XA.XIR[13].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.Iout 0.06446f
C2133 XThR.Tn[6] XA.XIR[7].XIC[9].icell.PDM 0.04035f
C2134 XA.XIR[6].XIC[0].icell.Ien VPWR 0.18829f
C2135 XA.XIR[12].XIC[4].icell.PDM XA.XIR[12].XIC[4].icell.Ien 0.04854f
C2136 XThR.XTB5.A XThR.XTB7.B 0.30355f
C2137 XThC.Tn[2] XA.XIR[10].XIC[2].icell.PDM 0.02601f
C2138 XA.XIR[15].XIC_dummy_left.icell.Iout VPWR 0.24997f
C2139 XThR.Tn[13] XA.XIR[13].XIC[8].icell.Ien 0.14211f
C2140 XThC.Tn[10] XA.XIR[7].XIC[10].icell.Ien 0.04604f
C2141 XA.XIR[0].XIC_dummy_left.icell.Iout Iout 0.03553f
C2142 a_6243_9615# XThC.Tn[6] 0.26385f
C2143 XA.XIR[5].XIC[7].icell.Ien Vbias 0.19161f
C2144 XA.XIR[13].XIC[2].icell.Ien Iout 0.06801f
C2145 XA.XIR[11].XIC[4].icell.PDM VPWR 0.01171f
C2146 XA.XIR[10].XIC[8].icell.PDM VPWR 0.01171f
C2147 XA.XIR[0].XIC_dummy_right.icell.Iout VPWR 0.12361f
C2148 XA.XIR[11].XIC_dummy_right.icell.Iout XA.XIR[12].XIC_dummy_right.icell.Iout 0.04047f
C2149 XA.XIR[11].XIC[5].icell.Ien Iout 0.06801f
C2150 XThR.XTB6.A XThR.XTB5.Y 0.01866f
C2151 XA.XIR[12].XIC[2].icell.Ien Vbias 0.19161f
C2152 XA.XIR[6].XIC[5].icell.Ien VPWR 0.18829f
C2153 XA.XIR[10].XIC[7].icell.Ien Iout 0.06801f
C2154 XA.XIR[0].XIC_15.icell.PDM Vbias 0.03947f
C2155 XThC.XTB7.Y Vbias 0.01962f
C2156 XThC.Tn[7] XA.XIR[1].XIC[7].icell.PDM 0.02602f
C2157 XThC.Tn[11] XA.XIR[10].XIC[11].icell.PDM 0.02601f
C2158 bias[2] bias[1] 0.67657f
C2159 XThC.Tn[7] XA.XIR[4].XIC[7].icell.PDM 0.02601f
C2160 XThC.Tn[12] XA.XIR[9].XIC[12].icell.Ien 0.04604f
C2161 XThC.XTB5.A XThC.XTBN.A 0.06305f
C2162 XThR.Tn[6] XA.XIR[6].XIC[13].icell.Ien 0.14211f
C2163 XA.XIR[2].XIC[0].icell.PDM VPWR 0.01171f
C2164 XThC.XTB7.A XThC.XTB3.Y 0.57441f
C2165 XThC.Tn[0] XA.XIR[7].XIC[0].icell.PDM 0.02601f
C2166 XThC.Tn[2] XA.XIR[11].XIC[2].icell.Ien 0.04604f
C2167 XThC.Tn[11] XA.XIR[9].XIC[11].icell.PDM 0.02601f
C2168 XA.XIR[6].XIC_dummy_left.icell.PUM VPWR 0.01669f
C2169 XA.XIR[2].XIC[9].icell.Ien Iout 0.06801f
C2170 XThC.XTB7.A XThC.Tn[2] 0.1255f
C2171 XA.XIR[10].XIC[13].icell.PDM VPWR 0.01171f
C2172 XA.XIR[12].XIC[0].icell.PDM XA.XIR[12].XIC[0].icell.Ien 0.04854f
C2173 XA.XIR[1].XIC[11].icell.Ien Iout 0.06801f
C2174 XA.XIR[0].XIC_dummy_right.icell.PDM VPWR 0.08055f
C2175 XThC.Tn[13] XA.XIR[1].XIC[13].icell.Ien 0.04606f
C2176 XA.XIR[11].XIC[4].icell.Ien VPWR 0.18829f
C2177 XThR.Tn[11] XA.XIR[12].XIC[0].icell.PDM 0.04042f
C2178 XThC.Tn[6] XA.XIR[8].XIC[6].icell.PDM 0.02601f
C2179 XA.XIR[13].XIC[14].icell.PDM VPWR 0.0118f
C2180 XA.XIR[10].XIC[6].icell.Ien VPWR 0.18829f
C2181 XThR.Tn[11] XA.XIR[11].XIC[12].icell.Ien 0.14211f
C2182 XThC.Tn[11] XThR.Tn[6] 0.40738f
C2183 XA.XIR[0].XIC[11].icell.PDM XA.XIR[0].XIC[11].icell.Ien 0.04854f
C2184 XA.XIR[13].XIC_15.icell.PDM XA.XIR[13].XIC_15.icell.Ien 0.04854f
C2185 XA.XIR[3].XIC_15.icell.Ien VPWR 0.26829f
C2186 XThR.XTB6.Y XThR.Tn[11] 0.02465f
C2187 XThC.Tn[13] XThR.Tn[11] 0.40739f
C2188 XThR.Tn[10] Iout 1.12758f
C2189 XA.XIR[1].XIC_dummy_left.icell.Ien VPWR 0.39039f
C2190 XThR.XTB1.Y XThR.XTB6.A 0.01609f
C2191 XA.XIR[2].XIC[8].icell.Ien VPWR 0.18829f
C2192 XThR.Tn[0] Vbias 1.39647f
C2193 XThC.Tn[3] XThR.Tn[7] 0.40738f
C2194 XThC.Tn[9] Iout 0.22393f
C2195 XThR.Tn[10] XA.XIR[11].XIC_dummy_left.icell.Iout 0.01758f
C2196 XA.XIR[4].XIC_dummy_left.icell.Ien VPWR 0.38912f
C2197 XA.XIR[1].XIC[10].icell.Ien VPWR 0.18829f
C2198 XThR.Tn[8] XA.XIR[8].XIC[5].icell.Ien 0.14211f
C2199 XThR.Tn[7] XA.XIR[8].XIC[2].icell.PDM 0.04035f
C2200 XThC.XTB6.Y XThC.Tn[9] 0.0246f
C2201 XA.XIR[6].XIC[6].icell.PDM Vbias 0.03928f
C2202 XThC.Tn[3] XA.XIR[15].XIC[3].icell.PDM 0.02601f
C2203 XA.XIR[5].XIC[10].icell.Ien XA.XIR[6].XIC[10].icell.PDM 0.02104f
C2204 XThC.XTBN.A data[0] 0.02545f
C2205 XThR.XTB1.Y XThR.Tn[0] 0.1837f
C2206 XThC.Tn[4] XA.XIR[0].XIC[4].icell.PDM 0.02803f
C2207 XA.XIR[5].XIC[13].icell.PDM Vbias 0.03928f
C2208 XA.XIR[14].XIC[3].icell.PDM Vbias 0.03928f
C2209 XThC.Tn[10] XA.XIR[8].XIC[10].icell.Ien 0.04604f
C2210 XThC.Tn[14] XA.XIR[12].XIC[14].icell.Ien 0.04604f
C2211 XThC.Tn[12] XA.XIR[5].XIC[12].icell.PDM 0.02601f
C2212 XA.XIR[3].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2213 XA.XIR[13].XIC[7].icell.PDM Vbias 0.03928f
C2214 XA.XIR[14].XIC[3].icell.PDM XA.XIR[14].XIC[3].icell.Ien 0.04854f
C2215 XThR.Tn[5] XA.XIR[5].XIC[4].icell.Ien 0.14211f
C2216 XThR.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.04035f
C2217 XThR.XTB7.B XThR.Tn[9] 0.0565f
C2218 XA.XIR[7].XIC[0].icell.PDM VPWR 0.01171f
C2219 XThC.XTB5.A XThC.XTB3.Y 0.01156f
C2220 XThC.XTB1.Y XThC.XTB7.A 0.48957f
C2221 XA.XIR[9].XIC[3].icell.Ien Vbias 0.19161f
C2222 XThC.Tn[2] XA.XIR[13].XIC[2].icell.PDM 0.02601f
C2223 XA.XIR[6].XIC[7].icell.PDM VPWR 0.01171f
C2224 XA.XIR[6].XIC[11].icell.Ien Iout 0.06801f
C2225 XThC.Tn[2] XThR.Tn[3] 0.40738f
C2226 XThR.Tn[14] XA.XIR[14].XIC[9].icell.Ien 0.14211f
C2227 XA.XIR[14].XIC[4].icell.PDM VPWR 0.01171f
C2228 XThC.XTBN.Y XThC.Tn[14] 0.42645f
C2229 XThR.Tn[1] XA.XIR[1].XIC[9].icell.Ien 0.14211f
C2230 XThC.Tn[11] XThR.Tn[4] 0.40738f
C2231 XThC.Tn[13] XA.XIR[6].XIC[13].icell.Ien 0.04604f
C2232 XA.XIR[5].XIC[14].icell.PDM VPWR 0.0118f
C2233 XThC.Tn[4] XA.XIR[2].XIC[4].icell.Ien 0.04605f
C2234 XThR.XTB5.A XThR.XTB4.Y 0.02767f
C2235 XA.XIR[1].XIC[0].icell.PDM Vbias 0.03915f
C2236 XA.XIR[11].XIC[13].icell.Ien XA.XIR[12].XIC[13].icell.PDM 0.02104f
C2237 XA.XIR[13].XIC[8].icell.PDM VPWR 0.01171f
C2238 XThC.XTB4.Y XThC.Tn[9] 0.01318f
C2239 XThC.Tn[1] XA.XIR[15].XIC[1].icell.Ien 0.04292f
C2240 XA.XIR[14].XIC[5].icell.Ien Iout 0.06801f
C2241 XThC.XTB7.Y a_10051_9569# 0.013f
C2242 XThR.Tn[11] XA.XIR[11].XIC[10].icell.Ien 0.14211f
C2243 XA.XIR[11].XIC[9].icell.Ien XA.XIR[12].XIC[9].icell.PDM 0.02104f
C2244 XA.XIR[4].XIC[0].icell.PDM Vbias 0.03915f
C2245 XThC.Tn[5] XThR.Tn[0] 0.40765f
C2246 XA.XIR[5].XIC[12].icell.Ien Vbias 0.19161f
C2247 XA.XIR[13].XIC[7].icell.Ien Iout 0.06801f
C2248 XA.XIR[8].XIC[0].icell.Ien XThR.Tn[8] 0.14211f
C2249 XThC.Tn[7] XThR.Tn[5] 0.40738f
C2250 XA.XIR[3].XIC[8].icell.PDM Vbias 0.03928f
C2251 XA.XIR[8].XIC[10].icell.PDM Vbias 0.03928f
C2252 XA.XIR[2].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2253 XA.XIR[0].XIC[4].icell.PDM XA.XIR[0].XIC[4].icell.Ien 0.04854f
C2254 XA.XIR[2].XIC[14].icell.PDM Vbias 0.03928f
C2255 XThC.Tn[11] XA.XIR[13].XIC[11].icell.PDM 0.02601f
C2256 XA.XIR[10].XIC[12].icell.PDM VPWR 0.01171f
C2257 XThC.Tn[6] XA.XIR[9].XIC[6].icell.PDM 0.02601f
C2258 XA.XIR[1].XIC[1].icell.PDM VPWR 0.01171f
C2259 XA.XIR[5].XIC[1].icell.PDM XA.XIR[5].XIC[1].icell.Ien 0.04854f
C2260 XA.XIR[6].XIC[10].icell.Ien VPWR 0.18829f
C2261 XThC.Tn[2] XA.XIR[14].XIC[2].icell.Ien 0.04604f
C2262 XA.XIR[12].XIC[7].icell.Ien Vbias 0.19161f
C2263 XA.XIR[11].XIC[0].icell.Ien XThR.Tn[11] 0.14211f
C2264 XA.XIR[13].XIC[13].icell.PDM VPWR 0.01171f
C2265 XA.XIR[4].XIC[1].icell.PDM VPWR 0.01171f
C2266 XA.XIR[3].XIC[9].icell.PDM VPWR 0.01171f
C2267 XThC.XTB3.Y data[0] 0.03253f
C2268 XA.XIR[14].XIC[4].icell.Ien VPWR 0.18883f
C2269 XA.XIR[8].XIC[11].icell.PDM VPWR 0.01171f
C2270 XThR.XTB5.Y XThR.Tn[12] 0.32095f
C2271 XA.XIR[2].XIC_15.icell.PDM VPWR 0.07527f
C2272 XThC.XTBN.A a_8739_9569# 0.01719f
C2273 XA.XIR[13].XIC[6].icell.Ien VPWR 0.18829f
C2274 XThR.Tn[8] XA.XIR[9].XIC[0].icell.PDM 0.0404f
C2275 XA.XIR[2].XIC[14].icell.Ien Iout 0.06801f
C2276 XThR.Tn[12] XA.XIR[13].XIC[5].icell.PDM 0.04035f
C2277 XA.XIR[5].XIC[3].icell.Ien XA.XIR[6].XIC[3].icell.PDM 0.02104f
C2278 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.Iout 0.06446f
C2279 XA.XIR[11].XIC_15.icell.PUM VPWR 0.01655f
C2280 XThC.Tn[4] XThR.Tn[2] 0.40741f
C2281 XA.XIR[1].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2282 XA.XIR[14].XIC[0].icell.Ien Iout 0.06795f
C2283 XThC.XTB5.A XThC.XTB1.Y 0.1098f
C2284 XA.XIR[11].XIC[9].icell.Ien VPWR 0.18829f
C2285 XThC.Tn[13] XThR.Tn[14] 0.40739f
C2286 XA.XIR[1].XIC[0].icell.Ien Vbias 0.1916f
C2287 XA.XIR[4].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2288 XThR.Tn[13] Iout 1.12765f
C2289 XA.XIR[2].XIC[11].icell.Ien XA.XIR[3].XIC[11].icell.PDM 0.02104f
C2290 XA.XIR[7].XIC[12].icell.Ien XA.XIR[8].XIC[12].icell.PDM 0.02104f
C2291 XA.XIR[4].XIC[0].icell.Ien Vbias 0.19149f
C2292 XThR.XTB3.Y XThR.XTBN.A 0.03907f
C2293 XThR.Tn[1] Vbias 1.39531f
C2294 a_7875_9569# XThC.Tn[9] 0.19271f
C2295 XThC.XTB2.Y XThC.Tn[9] 0.292f
C2296 XThR.Tn[0] XA.XIR[1].XIC[13].icell.PDM 0.0404f
C2297 XA.XIR[1].XIC[14].icell.Ien XA.XIR[2].XIC[14].icell.PDM 0.02104f
C2298 XThR.Tn[5] XA.XIR[6].XIC_dummy_left.icell.Iout 0.01728f
C2299 XA.XIR[5].XIC[4].icell.Ien Iout 0.06801f
C2300 XThR.Tn[12] Vbias 1.39531f
C2301 XThR.Tn[1] XA.XIR[2].XIC[12].icell.PDM 0.04035f
C2302 XA.XIR[13].XIC[12].icell.PDM XA.XIR[13].XIC[12].icell.Ien 0.04854f
C2303 XA.XIR[2].XIC[13].icell.Ien VPWR 0.18829f
C2304 XThR.XTBN.Y XThR.Tn[9] 0.48067f
C2305 XThC.Tn[7] XA.XIR[5].XIC[7].icell.PDM 0.02601f
C2306 XThC.Tn[0] XThR.Tn[6] 0.40736f
C2307 XA.XIR[7].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2308 XA.XIR[1].XIC_15.icell.Ien VPWR 0.26829f
C2309 XA.XIR[15].XIC[2].icell.Ien Vbias 0.15966f
C2310 XA.XIR[11].XIC[2].icell.Ien XA.XIR[12].XIC[2].icell.PDM 0.02104f
C2311 XThC.XTBN.A XThC.Tn[11] 0.11997f
C2312 XThR.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.144f
C2313 XA.XIR[7].XIC[14].icell.PDM Vbias 0.03928f
C2314 XThR.Tn[8] XA.XIR[8].XIC[10].icell.Ien 0.14211f
C2315 XA.XIR[6].XIC[12].icell.PDM XA.XIR[6].XIC[12].icell.Ien 0.04854f
C2316 XThC.Tn[9] XA.XIR[1].XIC[9].icell.PDM 0.02602f
C2317 XA.XIR[7].XIC_dummy_right.icell.Ien XA.XIR[8].XIC_dummy_right.icell.PDM 0.02104f
C2318 XThC.Tn[2] XThR.Tn[11] 0.40738f
C2319 XA.XIR[4].XIC[5].icell.Ien Vbias 0.19161f
C2320 XA.XIR[0].XIC_dummy_right.icell.Ien VPWR 0.35555f
C2321 XThC.Tn[9] XA.XIR[4].XIC[9].icell.PDM 0.02601f
C2322 XThC.XTBN.Y a_4067_9615# 0.08456f
C2323 XA.XIR[10].XIC[5].icell.Ien XA.XIR[11].XIC[5].icell.PDM 0.02104f
C2324 XThR.Tn[11] XA.XIR[11].XIC_15.icell.Ien 0.13564f
C2325 VPWR bias[1] 1.65687f
C2326 XA.XIR[10].XIC[6].icell.PDM XA.XIR[10].XIC[6].icell.Ien 0.04854f
C2327 XA.XIR[1].XIC_dummy_left.icell.Iout Iout 0.03553f
C2328 XA.XIR[9].XIC[10].icell.PDM Vbias 0.03928f
C2329 XThC.Tn[7] Iout 0.22453f
C2330 XThC.XTB1.Y data[0] 0.06453f
C2331 XThR.Tn[5] XA.XIR[5].XIC[9].icell.Ien 0.14211f
C2332 XThC.Tn[8] Vbias 0.79784f
C2333 XThR.XTB4.Y XThR.Tn[9] 0.01318f
C2334 XA.XIR[0].XIC[2].icell.PDM Vbias 0.03945f
C2335 XA.XIR[5].XIC[3].icell.Ien VPWR 0.18829f
C2336 XA.XIR[7].XIC_15.icell.PDM VPWR 0.07527f
C2337 XA.XIR[15].XIC_dummy_left.icell.PDM XA.XIR[15].XIC_dummy_left.icell.Ien 0.04854f
C2338 XThC.XTB3.Y a_8739_9569# 0.07285f
C2339 XThC.Tn[8] XA.XIR[8].XIC[8].icell.PDM 0.02601f
C2340 XA.XIR[6].XIC_dummy_right.icell.PDM XA.XIR[6].XIC_dummy_right.icell.Ien 0.04854f
C2341 XThC.XTB6.Y XThC.Tn[7] 0.01474f
C2342 XA.XIR[9].XIC[8].icell.Ien Vbias 0.19161f
C2343 XThR.Tn[9] XThR.Tn[10] 0.12586f
C2344 XA.XIR[1].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2345 XThC.Tn[5] XThR.Tn[1] 0.40744f
C2346 XThR.Tn[1] XA.XIR[1].XIC[14].icell.Ien 0.144f
C2347 XThC.Tn[3] XA.XIR[0].XIC[3].icell.Ien 0.04658f
C2348 XA.XIR[10].XIC[11].icell.PDM VPWR 0.01171f
C2349 XThC.Tn[9] XThR.Tn[9] 0.40738f
C2350 XA.XIR[1].XIC_15.icell.PDM Vbias 0.03927f
C2351 XA.XIR[10].XIC[10].icell.PDM XA.XIR[10].XIC[10].icell.Ien 0.04854f
C2352 XA.XIR[9].XIC[11].icell.PDM VPWR 0.01171f
C2353 XThC.Tn[5] XThR.Tn[12] 0.40738f
C2354 XThC.Tn[8] XA.XIR[11].XIC[8].icell.Ien 0.04604f
C2355 XThC.Tn[14] XThR.Tn[8] 0.40742f
C2356 XA.XIR[13].XIC[12].icell.PDM VPWR 0.01171f
C2357 XA.XIR[0].XIC[3].icell.PDM VPWR 0.01132f
C2358 XA.XIR[7].XIC[4].icell.Ien Vbias 0.19161f
C2359 XA.XIR[9].XIC_15.icell.PDM XA.XIR[9].XIC_15.icell.Ien 0.04854f
C2360 XA.XIR[4].XIC_15.icell.PDM Vbias 0.03927f
C2361 XThC.XTB6.Y a_5949_10571# 0.01283f
C2362 XA.XIR[7].XIC[13].icell.PDM XA.XIR[7].XIC[13].icell.Ien 0.04854f
C2363 XThR.XTB3.Y a_n1049_7493# 0.23056f
C2364 XThC.XTBN.Y XThC.Tn[3] 0.49586f
C2365 XA.XIR[2].XIC[4].icell.Ien XA.XIR[3].XIC[4].icell.PDM 0.02104f
C2366 XA.XIR[4].XIC[14].icell.PDM XA.XIR[4].XIC[14].icell.Ien 0.04854f
C2367 XA.XIR[11].XIC[0].icell.PDM XA.XIR[11].XIC[0].icell.Ien 0.04854f
C2368 XThC.Tn[0] XThR.Tn[4] 0.40739f
C2369 XThR.XTBN.A VPWR 0.90694f
C2370 XThC.Tn[10] XA.XIR[11].XIC[10].icell.PDM 0.02601f
C2371 XA.XIR[7].XIC[5].icell.Ien XA.XIR[8].XIC[5].icell.PDM 0.02104f
C2372 XThC.Tn[0] XA.XIR[12].XIC[0].icell.PDM 0.02601f
C2373 XA.XIR[12].XIC[1].icell.Ien XThR.Tn[12] 0.14211f
C2374 XA.XIR[10].XIC[1].icell.Ien XA.XIR[11].XIC[1].icell.PDM 0.02104f
C2375 XThR.XTB5.Y a_n1049_6405# 0.24821f
C2376 XThR.Tn[4] XA.XIR[5].XIC[10].icell.PDM 0.04035f
C2377 XThC.Tn[5] XA.XIR[4].XIC[5].icell.Ien 0.04604f
C2378 XThR.Tn[14] XA.XIR[15].XIC[0].icell.PDM 0.04042f
C2379 XA.XIR[11].XIC[14].icell.Ien VPWR 0.18835f
C2380 XThR.Tn[6] VPWR 7.9997f
C2381 XA.XIR[1].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2382 XThR.XTB3.Y XThR.XTB6.Y 0.04428f
C2383 XThC.Tn[14] XA.XIR[6].XIC[14].icell.PDM 0.02601f
C2384 XThC.XTB4.Y XThC.Tn[7] 0.01805f
C2385 XA.XIR[1].XIC[7].icell.Ien XA.XIR[2].XIC[7].icell.PDM 0.02104f
C2386 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Ien 0.01532f
C2387 XA.XIR[6].XIC_15.icell.Ien VPWR 0.26829f
C2388 XThC.Tn[4] XThR.Tn[10] 0.40738f
C2389 XA.XIR[8].XIC[12].icell.PDM XA.XIR[8].XIC[12].icell.Ien 0.04854f
C2390 XThR.Tn[14] XA.XIR[14].XIC[12].icell.Ien 0.14211f
C2391 XThC.Tn[11] XA.XIR[3].XIC[11].icell.PDM 0.02601f
C2392 XA.XIR[14].XIC_15.icell.PUM VPWR 0.01655f
C2393 XA.XIR[4].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2394 XThC.Tn[14] XA.XIR[15].XIC[14].icell.Ien 0.04292f
C2395 XA.XIR[0].XIC[11].icell.Ien XA.XIR[1].XIC[11].icell.PDM 0.02104f
C2396 XA.XIR[14].XIC[9].icell.Ien VPWR 0.18883f
C2397 XA.XIR[6].XIC[5].icell.PDM XA.XIR[6].XIC[5].icell.Ien 0.04854f
C2398 a_4861_9615# XThC.Tn[3] 0.26251f
C2399 XA.XIR[15].XIC[4].icell.PDM XA.XIR[15].XIC[4].icell.Ien 0.04854f
C2400 XA.XIR[6].XIC_dummy_left.icell.Iout Iout 0.03553f
C2401 XA.XIR[2].XIC_dummy_left.icell.Ien VPWR 0.38902f
C2402 XA.XIR[3].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2403 XThR.Tn[3] XA.XIR[3].XIC[2].icell.Ien 0.14211f
C2404 XA.XIR[5].XIC[0].icell.PDM Vbias 0.03915f
C2405 XThR.Tn[13] XA.XIR[14].XIC_dummy_left.icell.Iout 0.0222f
C2406 XA.XIR[9].XIC[4].icell.Ien XA.XIR[10].XIC[4].icell.PDM 0.02104f
C2407 XA.XIR[8].XIC_dummy_right.icell.PDM XA.XIR[8].XIC_dummy_right.icell.Ien 0.04854f
C2408 XA.XIR[6].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2409 XThR.Tn[5] XA.XIR[6].XIC[12].icell.PDM 0.04035f
C2410 XA.XIR[14].XIC_dummy_right.icell.Iout XA.XIR[15].XIC_dummy_right.icell.Iout 0.04047f
C2411 XA.XIR[11].XIC[5].icell.PDM Vbias 0.03928f
C2412 XThC.Tn[4] XA.XIR[1].XIC[4].icell.PDM 0.02602f
C2413 XThR.Tn[2] XA.XIR[3].XIC[4].icell.PDM 0.04035f
C2414 XA.XIR[9].XIC_dummy_left.icell.Ien XA.XIR[10].XIC_dummy_left.icell.PDM 0.02104f
C2415 XA.XIR[10].XIC[9].icell.PDM Vbias 0.03928f
C2416 XA.XIR[5].XIC[1].icell.PDM VPWR 0.01171f
C2417 XA.XIR[5].XIC[9].icell.Ien Iout 0.06801f
C2418 XThC.Tn[4] XA.XIR[4].XIC[4].icell.PDM 0.02601f
C2419 XThC.Tn[2] XThR.Tn[14] 0.40738f
C2420 XThC.Tn[3] XA.XIR[3].XIC[3].icell.Ien 0.04604f
C2421 XThC.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.02601f
C2422 XThR.Tn[6] XA.XIR[7].XIC[11].icell.PDM 0.04035f
C2423 XThR.Tn[4] VPWR 8.03623f
C2424 XA.XIR[6].XIC[14].icell.Ien XA.XIR[7].XIC[14].icell.PDM 0.02104f
C2425 XThC.Tn[10] XA.XIR[2].XIC[10].icell.Ien 0.04605f
C2426 XA.XIR[12].XIC[0].icell.PDM VPWR 0.01171f
C2427 XA.XIR[15].XIC[7].icell.Ien Vbias 0.15966f
C2428 XA.XIR[9].XIC[8].icell.PDM XA.XIR[9].XIC[8].icell.Ien 0.04854f
C2429 XThR.Tn[8] XA.XIR[8].XIC_15.icell.Ien 0.13564f
C2430 a_n1049_7493# VPWR 0.72084f
C2431 XA.XIR[7].XIC[6].icell.PDM XA.XIR[7].XIC[6].icell.Ien 0.04854f
C2432 XA.XIR[11].XIC[6].icell.PDM VPWR 0.01171f
C2433 XA.XIR[11].XIC[12].icell.Ien VPWR 0.18829f
C2434 XA.XIR[14].XIC[13].icell.Ien XA.XIR[15].XIC[13].icell.PDM 0.02104f
C2435 XThC.Tn[3] XA.XIR[8].XIC[3].icell.PDM 0.02601f
C2436 XA.XIR[4].XIC[7].icell.PDM XA.XIR[4].XIC[7].icell.Ien 0.04854f
C2437 XA.XIR[4].XIC[10].icell.Ien Vbias 0.19161f
C2438 XA.XIR[12].XIC[4].icell.Ien Iout 0.06801f
C2439 XA.XIR[0].XIC[1].icell.Ien Vbias 0.19213f
C2440 XA.XIR[10].XIC[10].icell.PDM VPWR 0.01171f
C2441 XA.XIR[2].XIC[1].icell.PDM Vbias 0.03928f
C2442 XThR.Tn[14] XA.XIR[14].XIC[10].icell.Ien 0.14211f
C2443 XA.XIR[14].XIC[9].icell.Ien XA.XIR[15].XIC[9].icell.PDM 0.02104f
C2444 XThR.XTB6.Y VPWR 1.05512f
C2445 XA.XIR[8].XIC[4].icell.Ien Vbias 0.19161f
C2446 XThC.Tn[13] VPWR 4.60106f
C2447 XA.XIR[13].XIC[11].icell.PDM VPWR 0.01171f
C2448 XThR.Tn[5] XA.XIR[5].XIC[14].icell.Ien 0.144f
C2449 XA.XIR[9].XIC[12].icell.Ien XA.XIR[10].XIC[12].icell.PDM 0.02104f
C2450 XA.XIR[8].XIC[5].icell.PDM XA.XIR[8].XIC[5].icell.Ien 0.04854f
C2451 XA.XIR[5].XIC[8].icell.Ien VPWR 0.18829f
C2452 XA.XIR[8].XIC_dummy_right.icell.Iout XA.XIR[9].XIC_dummy_right.icell.Iout 0.04047f
C2453 XA.XIR[10].XIC_dummy_left.icell.Iout VPWR 0.11161f
C2454 XThC.Tn[8] XA.XIR[14].XIC[8].icell.Ien 0.04604f
C2455 XA.XIR[9].XIC[13].icell.Ien Vbias 0.19161f
C2456 XThC.Tn[0] XA.XIR[11].XIC[0].icell.Ien 0.04604f
C2457 XA.XIR[0].XIC[4].icell.Ien XA.XIR[1].XIC[4].icell.PDM 0.02104f
C2458 XThC.XTB6.A XThC.XTB7.Y 0.01596f
C2459 XA.XIR[10].XIC[14].icell.Ien XA.XIR[11].XIC[14].icell.PDM 0.02104f
C2460 XA.XIR[0].XIC[6].icell.Ien Vbias 0.19213f
C2461 XA.XIR[8].XIC[12].icell.Ien XA.XIR[9].XIC[12].icell.PDM 0.02104f
C2462 XA.XIR[2].XIC[2].icell.PDM VPWR 0.01171f
C2463 XThC.Tn[5] XA.XIR[11].XIC[5].icell.PDM 0.02601f
C2464 XThC.Tn[10] XA.XIR[14].XIC[10].icell.PDM 0.02601f
C2465 XA.XIR[3].XIC[11].icell.Ien XA.XIR[4].XIC[11].icell.PDM 0.02104f
C2466 XThC.Tn[0] XA.XIR[15].XIC[0].icell.PDM 0.02601f
C2467 XA.XIR[12].XIC[3].icell.Ien VPWR 0.18829f
C2468 XThC.Tn[6] Vbias 0.81928f
C2469 XThC.Tn[1] XA.XIR[0].XIC[1].icell.PDM 0.02803f
C2470 XA.XIR[14].XIC[14].icell.Ien VPWR 0.1889f
C2471 XA.XIR[3].XIC[13].icell.PDM XA.XIR[3].XIC[13].icell.Ien 0.04854f
C2472 XA.XIR[7].XIC[9].icell.Ien Vbias 0.19161f
C2473 XThC.Tn[6] XA.XIR[3].XIC[6].icell.PDM 0.02601f
C2474 XThR.Tn[11] XA.XIR[12].XIC[2].icell.PDM 0.04035f
C2475 XThC.Tn[4] XThR.Tn[13] 0.40738f
C2476 XThC.Tn[9] XA.XIR[5].XIC[9].icell.PDM 0.02601f
C2477 XThR.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.14211f
C2478 XA.XIR[11].XIC[11].icell.Ien XA.XIR[12].XIC[11].icell.PDM 0.02104f
C2479 XThC.XTB2.Y a_3773_9615# 0.2342f
C2480 XThR.Tn[7] Iout 1.1276f
C2481 XA.XIR[8].XIC_dummy_right.icell.Ien XA.XIR[9].XIC_dummy_right.icell.PDM 0.02104f
C2482 XThC.Tn[7] XThR.Tn[9] 0.40738f
C2483 XThC.Tn[3] XThR.Tn[8] 0.40738f
C2484 XThR.Tn[0] XA.XIR[1].XIC[0].icell.PDM 0.0404f
C2485 XThC.Tn[4] XA.XIR[5].XIC[4].icell.Ien 0.04604f
C2486 XA.XIR[2].XIC[0].icell.Ien Vbias 0.19149f
C2487 XA.XIR[3].XIC[0].icell.PDM XA.XIR[3].XIC[0].icell.Ien 0.04854f
C2488 XThR.Tn[10] XA.XIR[10].XIC[13].icell.Ien 0.14211f
C2489 XA.XIR[4].XIC[2].icell.Ien Iout 0.06801f
C2490 XA.XIR[6].XIC[7].icell.Ien XA.XIR[7].XIC[7].icell.PDM 0.02104f
C2491 XA.XIR[11].XIC[10].icell.Ien VPWR 0.18829f
C2492 XThR.Tn[7] XA.XIR[8].XIC[4].icell.PDM 0.04035f
C2493 XA.XIR[10].XIC[1].icell.Ien Vbias 0.19161f
C2494 XA.XIR[7].XIC[1].icell.PDM Vbias 0.03928f
C2495 XA.XIR[6].XIC[8].icell.PDM Vbias 0.03928f
C2496 XThC.XTBN.A VPWR 0.88815f
C2497 XThR.Tn[12] XA.XIR[12].XIC[2].icell.Ien 0.14211f
C2498 XA.XIR[14].XIC[5].icell.PDM Vbias 0.03928f
C2499 XThR.Tn[3] XA.XIR[3].XIC[7].icell.Ien 0.14211f
C2500 XA.XIR[5].XIC_15.icell.PDM Vbias 0.03927f
C2501 XA.XIR[14].XIC[2].icell.Ien XA.XIR[15].XIC[2].icell.PDM 0.02104f
C2502 XA.XIR[9].XIC[5].icell.Ien Iout 0.06801f
C2503 XA.XIR[13].XIC[9].icell.PDM Vbias 0.03928f
C2504 XA.XIR[4].XIC[14].icell.Ien XA.XIR[5].XIC[14].icell.PDM 0.02104f
C2505 XA.XIR[11].XIC[0].icell.Ien VPWR 0.18829f
C2506 XA.XIR[12].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2507 XThC.Tn[5] XThC.Tn[6] 0.14629f
C2508 XThR.Tn[3] XA.XIR[4].XIC[5].icell.PDM 0.04035f
C2509 XThC.Tn[3] XA.XIR[9].XIC[3].icell.PDM 0.02601f
C2510 XA.XIR[7].XIC[2].icell.PDM VPWR 0.01171f
C2511 XA.XIR[13].XIC[5].icell.Ien XA.XIR[14].XIC[5].icell.PDM 0.02104f
C2512 XThR.Tn[2] XA.XIR[2].XIC[2].icell.Ien 0.14211f
C2513 XA.XIR[1].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2514 XThR.Tn[14] XA.XIR[14].XIC_15.icell.Ien 0.13564f
C2515 XA.XIR[5].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.PDM 0.02104f
C2516 XA.XIR[15].XIC[0].icell.PDM VPWR 0.01512f
C2517 XA.XIR[6].XIC[9].icell.PDM VPWR 0.01171f
C2518 XA.XIR[13].XIC[6].icell.PDM XA.XIR[13].XIC[6].icell.Ien 0.04854f
C2519 XA.XIR[11].XIC[13].icell.Ien Vbias 0.19161f
C2520 XA.XIR[14].XIC[6].icell.PDM VPWR 0.01171f
C2521 XA.XIR[5].XIC_dummy_right.icell.PDM VPWR 0.08209f
C2522 XA.XIR[8].XIC[5].icell.Ien XA.XIR[9].XIC[5].icell.PDM 0.02104f
C2523 XA.XIR[14].XIC[12].icell.Ien VPWR 0.18883f
C2524 XA.XIR[12].XIC[7].icell.Ien XA.XIR[13].XIC[7].icell.PDM 0.02104f
C2525 XA.XIR[5].XIC[14].icell.Ien Iout 0.06801f
C2526 XA.XIR[3].XIC[6].icell.Ien Vbias 0.19161f
C2527 XThC.Tn[2] XA.XIR[9].XIC[2].icell.Ien 0.04604f
C2528 XA.XIR[3].XIC[4].icell.Ien XA.XIR[4].XIC[4].icell.PDM 0.02104f
C2529 XA.XIR[13].XIC[10].icell.PDM VPWR 0.01171f
C2530 XA.XIR[1].XIC[2].icell.PDM Vbias 0.03928f
C2531 XThC.Tn[12] XA.XIR[10].XIC[12].icell.PDM 0.02601f
C2532 XThC.Tn[9] XA.XIR[0].XIC[9].icell.Ien 0.04656f
C2533 XThC.XTB7.Y XThC.Tn[8] 0.07809f
C2534 XA.XIR[3].XIC[6].icell.PDM XA.XIR[3].XIC[6].icell.Ien 0.04854f
C2535 XA.XIR[4].XIC[2].icell.PDM Vbias 0.03928f
C2536 XA.XIR[9].XIC[4].icell.Ien VPWR 0.18829f
C2537 XThR.Tn[0] XThR.Tn[1] 0.27134f
C2538 XA.XIR[3].XIC[10].icell.PDM Vbias 0.03928f
C2539 XThC.Tn[3] XA.XIR[1].XIC[3].icell.Ien 0.04607f
C2540 XA.XIR[8].XIC[12].icell.PDM Vbias 0.03928f
C2541 XA.XIR[12].XIC[9].icell.Ien Iout 0.06801f
C2542 XA.XIR[4].XIC_15.icell.Ien Vbias 0.19195f
C2543 XA.XIR[13].XIC[10].icell.PDM XA.XIR[13].XIC[10].icell.Ien 0.04854f
C2544 XA.XIR[13].XIC_dummy_left.icell.Iout VPWR 0.11047f
C2545 XThR.Tn[10] XA.XIR[10].XIC[11].icell.Ien 0.14211f
C2546 XA.XIR[8].XIC[9].icell.Ien Vbias 0.19161f
C2547 XThR.XTB7.A XThR.XTB5.Y 0.11935f
C2548 XA.XIR[1].XIC[3].icell.PDM VPWR 0.01171f
C2549 XThC.Tn[5] XA.XIR[14].XIC[5].icell.PDM 0.02601f
C2550 XA.XIR[9].XIC[0].icell.Ien Iout 0.06795f
C2551 XThC.Tn[11] XA.XIR[4].XIC[11].icell.Ien 0.04604f
C2552 XA.XIR[5].XIC[13].icell.Ien VPWR 0.18829f
C2553 XThR.Tn[4] XA.XIR[5].XIC_dummy_left.icell.Iout 0.01728f
C2554 XA.XIR[4].XIC[3].icell.PDM VPWR 0.01171f
C2555 XA.XIR[13].XIC[1].icell.Ien XA.XIR[14].XIC[1].icell.PDM 0.02104f
C2556 XThC.XTB3.Y VPWR 1.07064f
C2557 XA.XIR[4].XIC_dummy_right.icell.PUM VPWR 0.01691f
C2558 XThR.Tn[3] XA.XIR[4].XIC_dummy_left.icell.Iout 0.01728f
C2559 XA.XIR[3].XIC[11].icell.PDM VPWR 0.01171f
C2560 XThC.Tn[14] XThR.Tn[3] 0.40742f
C2561 XThC.XTB1.Y XThC.Tn[0] 0.1842f
C2562 XThC.Tn[4] XA.XIR[5].XIC[4].icell.PDM 0.02601f
C2563 XA.XIR[8].XIC[13].icell.PDM VPWR 0.01171f
C2564 XThC.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.04604f
C2565 XThC.XTBN.A a_9827_9569# 0.09118f
C2566 XA.XIR[0].XIC[11].icell.Ien Vbias 0.19213f
C2567 XThC.Tn[2] VPWR 3.64821f
C2568 XThR.Tn[8] XA.XIR[9].XIC[2].icell.PDM 0.04035f
C2569 XThR.Tn[12] XA.XIR[13].XIC[7].icell.PDM 0.04035f
C2570 XA.XIR[10].XIC_15.icell.Ien XA.XIR[11].XIC_15.icell.PDM 0.02104f
C2571 XA.XIR[11].XIC_15.icell.PDM VPWR 0.07527f
C2572 XA.XIR[11].XIC_15.icell.Ien VPWR 0.26829f
C2573 XA.XIR[12].XIC[8].icell.Ien VPWR 0.18829f
C2574 XA.XIR[1].XIC[0].icell.PDM XA.XIR[1].XIC[0].icell.Ien 0.04854f
C2575 XThC.Tn[8] XThR.Tn[0] 0.40759f
C2576 XA.XIR[6].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2577 XThC.Tn[10] XThR.Tn[5] 0.40738f
C2578 XA.XIR[4].XIC[7].icell.Ien XA.XIR[5].XIC[7].icell.PDM 0.02104f
C2579 XA.XIR[1].XIC[11].icell.PDM XA.XIR[1].XIC[11].icell.Ien 0.04854f
C2580 XA.XIR[7].XIC[14].icell.Ien Vbias 0.19161f
C2581 XA.XIR[9].XIC[1].icell.PDM XA.XIR[9].XIC[1].icell.Ien 0.04854f
C2582 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[12].XIC_dummy_right.icell.PDM 0.02104f
C2583 XA.XIR[11].XIC[11].icell.Ien Vbias 0.19161f
C2584 XThR.Tn[4] XA.XIR[4].XIC[9].icell.Ien 0.14211f
C2585 XThC.Tn[0] XA.XIR[7].XIC[0].icell.Ien 0.04604f
C2586 XA.XIR[14].XIC[10].icell.Ien VPWR 0.18883f
C2587 XA.XIR[4].XIC[0].icell.PDM XA.XIR[4].XIC[0].icell.Ien 0.04854f
C2588 XThC.XTB5.Y a_5155_9615# 0.24821f
C2589 XA.XIR[2].XIC[13].icell.PDM XA.XIR[2].XIC[13].icell.Ien 0.04854f
C2590 XA.XIR[13].XIC[1].icell.Ien Vbias 0.19161f
C2591 XThC.XTB7.A a_4067_9615# 0.0127f
C2592 XThR.XTB1.Y XThR.XTB7.A 0.48957f
C2593 XA.XIR[15].XIC[4].icell.Ien Iout 0.07192f
C2594 XThC.XTBN.A XThC.XTB7.B 0.35142f
C2595 XThR.Tn[1] XA.XIR[2].XIC[14].icell.PDM 0.04056f
C2596 XA.XIR[7].XIC_15.icell.PUM VPWR 0.01655f
C2597 XA.XIR[11].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2598 XA.XIR[4].XIC[7].icell.Ien Iout 0.06801f
C2599 XThC.Tn[3] XA.XIR[6].XIC[3].icell.Ien 0.04604f
C2600 XThR.Tn[7] XA.XIR[7].XIC[2].icell.Ien 0.14211f
C2601 XThC.Tn[9] XA.XIR[3].XIC[9].icell.Ien 0.04604f
C2602 XA.XIR[15].XIC_dummy_left.icell.PDM VPWR 0.08252f
C2603 XA.XIR[4].XIC[1].icell.Ien VPWR 0.18829f
C2604 XA.XIR[11].XIC[4].icell.PDM XA.XIR[11].XIC[4].icell.Ien 0.04854f
C2605 XThC.Tn[4] XA.XIR[12].XIC[4].icell.Ien 0.04604f
C2606 XThR.Tn[12] XA.XIR[12].XIC[7].icell.Ien 0.14211f
C2607 XThC.XTBN.Y a_5155_9615# 0.07602f
C2608 XA.XIR[7].XIC[1].icell.Ien Iout 0.06801f
C2609 XThR.Tn[3] XA.XIR[3].XIC[12].icell.Ien 0.14211f
C2610 XA.XIR[14].XIC[13].icell.Ien Vbias 0.19161f
C2611 XA.XIR[9].XIC[10].icell.Ien Iout 0.06801f
C2612 XThC.XTB1.Y VPWR 1.11809f
C2613 XA.XIR[9].XIC[12].icell.PDM Vbias 0.03928f
C2614 XA.XIR[12].XIC[14].icell.Ien Iout 0.06801f
C2615 XThC.XTB5.Y XThC.XTB6.Y 2.12831f
C2616 XA.XIR[0].XIC[4].icell.PDM Vbias 0.03945f
C2617 XA.XIR[15].XIC[3].icell.Ien VPWR 0.31713f
C2618 XThC.Tn[11] XA.XIR[6].XIC[11].icell.PDM 0.02601f
C2619 XA.XIR[0].XIC[3].icell.Ien Iout 0.0675f
C2620 XA.XIR[10].XIC_dummy_right.icell.Iout XA.XIR[11].XIC_dummy_right.icell.Iout 0.04047f
C2621 XThC.Tn[8] XA.XIR[3].XIC[8].icell.PDM 0.02601f
C2622 XThR.Tn[2] XA.XIR[2].XIC[7].icell.Ien 0.14211f
C2623 XThC.Tn[12] XA.XIR[13].XIC[12].icell.PDM 0.02601f
C2624 XA.XIR[1].XIC[1].icell.Ien Vbias 0.19173f
C2625 XA.XIR[4].XIC[6].icell.Ien VPWR 0.18829f
C2626 XThC.XTB7.A XThC.Tn[3] 0.0337f
C2627 XA.XIR[10].XIC[2].icell.Ien Vbias 0.19161f
C2628 XA.XIR[14].XIC_dummy_left.icell.Ien XThR.Tn[14] 0.01244f
C2629 XThR.Tn[1] XA.XIR[1].XIC[0].icell.Ien 0.14251f
C2630 XThR.XTB7.B XThR.XTB5.Y 0.30227f
C2631 XA.XIR[7].XIC[6].icell.Ien Iout 0.06801f
C2632 a_2979_9615# XThC.Tn[0] 0.27729f
C2633 XA.XIR[3].XIC[11].icell.Ien Vbias 0.19161f
C2634 XA.XIR[9].XIC[13].icell.PDM VPWR 0.01171f
C2635 XThC.Tn[12] XThR.Tn[6] 0.40738f
C2636 XA.XIR[7].XIC[0].icell.Ien VPWR 0.18829f
C2637 XA.XIR[1].XIC[4].icell.PDM XA.XIR[1].XIC[4].icell.Ien 0.04854f
C2638 XA.XIR[6].XIC[0].icell.Ien XA.XIR[7].XIC[0].icell.PDM 0.02104f
C2639 XA.XIR[0].XIC[5].icell.PDM VPWR 0.01261f
C2640 XThC.Tn[7] XA.XIR[8].XIC[7].icell.Ien 0.04604f
C2641 XA.XIR[2].XIC[4].icell.Ien Vbias 0.19161f
C2642 XA.XIR[13].XIC[14].icell.Ien XA.XIR[14].XIC[14].icell.PDM 0.02104f
C2643 XThC.XTB6.Y XThC.XTBN.Y 0.18947f
C2644 XA.XIR[9].XIC[9].icell.Ien VPWR 0.18829f
C2645 XA.XIR[1].XIC[6].icell.Ien Vbias 0.19173f
C2646 XThC.Tn[14] XThR.Tn[11] 0.40742f
C2647 XThR.Tn[9] XA.XIR[9].XIC[5].icell.Ien 0.14211f
C2648 XA.XIR[0].XIC[2].icell.Ien VPWR 0.18776f
C2649 XThR.Tn[10] XA.XIR[11].XIC[1].icell.PDM 0.04035f
C2650 XThC.XTB3.Y XThC.XTB7.B 0.23315f
C2651 XThC.XTB4.Y XThC.XTB5.Y 2.06459f
C2652 XThC.Tn[4] XThR.Tn[7] 0.40738f
C2653 XA.XIR[2].XIC[6].icell.PDM XA.XIR[2].XIC[6].icell.Ien 0.04854f
C2654 XA.XIR[11].XIC[14].icell.PDM VPWR 0.0118f
C2655 XThR.Tn[4] XA.XIR[5].XIC[12].icell.PDM 0.04035f
C2656 XA.XIR[8].XIC[14].icell.Ien Vbias 0.19161f
C2657 XThR.Tn[14] XA.XIR[15].XIC[2].icell.PDM 0.04035f
C2658 XThC.Tn[10] Iout 0.22426f
C2659 XThC.Tn[1] XA.XIR[1].XIC[1].icell.PDM 0.02602f
C2660 XThC.XTB7.Y XThC.Tn[6] 0.2182f
C2661 XThC.Tn[1] XA.XIR[4].XIC[1].icell.PDM 0.02601f
C2662 XA.XIR[14].XIC_15.icell.PDM VPWR 0.07527f
C2663 XA.XIR[14].XIC[11].icell.Ien XA.XIR[15].XIC[11].icell.PDM 0.02104f
C2664 XA.XIR[7].XIC[5].icell.Ien VPWR 0.18829f
C2665 XA.XIR[14].XIC_15.icell.Ien VPWR 0.26861f
C2666 XThC.XTB6.Y XThC.Tn[10] 0.02478f
C2667 XThC.Tn[10] XA.XIR[5].XIC[10].icell.Ien 0.04604f
C2668 XThC.Tn[8] XThR.Tn[1] 0.40744f
C2669 XThR.Tn[0] XA.XIR[0].XIC[1].icell.Ien 0.14211f
C2670 XA.XIR[14].XIC[11].icell.Ien Vbias 0.19161f
C2671 XThR.Tn[13] XA.XIR[13].XIC[13].icell.Ien 0.14211f
C2672 XA.XIR[8].XIC_15.icell.PUM VPWR 0.01655f
C2673 XThR.XTB7.B XThR.XTB1.Y 1.61695f
C2674 XThC.Tn[8] XThR.Tn[12] 0.40738f
C2675 XThC.XTB4.Y XThC.XTBN.Y 0.15636f
C2676 XThC.Tn[0] XA.XIR[8].XIC[0].icell.PDM 0.02601f
C2677 XA.XIR[5].XIC[2].icell.PDM Vbias 0.03928f
C2678 XA.XIR[5].XIC[9].icell.PDM XA.XIR[5].XIC[9].icell.Ien 0.04854f
C2679 XA.XIR[12].XIC[12].icell.Ien Iout 0.06801f
C2680 XA.XIR[6].XIC[1].icell.Ien Vbias 0.19161f
C2681 XThC.Tn[3] XThR.Tn[3] 0.40738f
C2682 XA.XIR[10].XIC[12].icell.Ien XA.XIR[11].XIC[12].icell.PDM 0.02104f
C2683 XA.XIR[12].XIC[1].icell.PDM Vbias 0.03928f
C2684 XThC.Tn[12] XThR.Tn[4] 0.40738f
C2685 XA.XIR[8].XIC[1].icell.Ien Iout 0.06801f
C2686 XA.XIR[14].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2687 XThR.Tn[2] Vbias 1.39527f
C2688 XThR.Tn[5] XA.XIR[6].XIC[14].icell.PDM 0.04056f
C2689 XThR.Tn[4] XA.XIR[4].XIC[14].icell.Ien 0.144f
C2690 XThC.Tn[14] XA.XIR[10].XIC[14].icell.Ien 0.04604f
C2691 a_2979_9615# VPWR 0.70527f
C2692 XA.XIR[11].XIC[7].icell.PDM Vbias 0.03928f
C2693 XA.XIR[3].XIC[3].icell.Ien Iout 0.06801f
C2694 XA.XIR[9].XIC[0].icell.Ien XThR.Tn[9] 0.14211f
C2695 XThR.Tn[0] XA.XIR[0].XIC[6].icell.Ien 0.14211f
C2696 XThR.Tn[10] XA.XIR[10].XIC[5].icell.Ien 0.14211f
C2697 XThC.XTB4.Y XThC.Tn[10] 0.01405f
C2698 XThR.Tn[2] XA.XIR[3].XIC[6].icell.PDM 0.04035f
C2699 XThC.Tn[12] XA.XIR[11].XIC[12].icell.Ien 0.04604f
C2700 XA.XIR[5].XIC[3].icell.PDM VPWR 0.01171f
C2701 XA.XIR[15].XIC[9].icell.Ien Iout 0.07192f
C2702 XThC.Tn[6] XThR.Tn[0] 0.40767f
C2703 XThC.XTB4.Y a_4861_9615# 0.23756f
C2704 XThC.Tn[2] XA.XIR[11].XIC[2].icell.PDM 0.02601f
C2705 XThR.Tn[6] XA.XIR[7].XIC[13].icell.PDM 0.0404f
C2706 XA.XIR[12].XIC[5].icell.PDM XA.XIR[12].XIC[5].icell.Ien 0.04854f
C2707 XA.XIR[6].XIC[6].icell.Ien Vbias 0.19161f
C2708 XA.XIR[4].XIC[12].icell.Ien Iout 0.06801f
C2709 XThR.Tn[7] XA.XIR[7].XIC[7].icell.Ien 0.14211f
C2710 XThC.Tn[12] XThC.Tn[13] 0.17915f
C2711 XA.XIR[12].XIC[2].icell.PDM VPWR 0.01171f
C2712 XThC.Tn[8] XA.XIR[9].XIC[8].icell.Ien 0.04604f
C2713 XThC.XTB2.Y XThC.XTB5.Y 0.0451f
C2714 XThC.Tn[6] XA.XIR[6].XIC[6].icell.PDM 0.02601f
C2715 XThC.XTB1.Y XThC.XTB7.B 1.61695f
C2716 XA.XIR[8].XIC[6].icell.Ien Iout 0.06801f
C2717 XThC.Tn[13] XA.XIR[2].XIC[13].icell.PDM 0.02602f
C2718 XA.XIR[11].XIC[8].icell.PDM VPWR 0.01171f
C2719 XThC.Tn[3] XA.XIR[3].XIC[3].icell.PDM 0.02601f
C2720 XThR.XTBN.Y XThR.XTB5.Y 0.16186f
C2721 XA.XIR[2].XIC[3].icell.PDM Vbias 0.03928f
C2722 XA.XIR[13].XIC[2].icell.Ien Vbias 0.19161f
C2723 XThC.Tn[9] XA.XIR[1].XIC[9].icell.Ien 0.04606f
C2724 XThR.Tn[9] XA.XIR[10].XIC[0].icell.PDM 0.04042f
C2725 XA.XIR[3].XIC[2].icell.Ien VPWR 0.18829f
C2726 XA.XIR[9].XIC_15.icell.Ien Iout 0.0694f
C2727 XThC.Tn[0] XA.XIR[8].XIC[0].icell.Ien 0.04604f
C2728 XA.XIR[4].XIC[0].icell.Ien XA.XIR[5].XIC[0].icell.PDM 0.02104f
C2729 XA.XIR[15].XIC[8].icell.Ien VPWR 0.31713f
C2730 XThC.Tn[11] XA.XIR[11].XIC[11].icell.PDM 0.02601f
C2731 XA.XIR[0].XIC[8].icell.Ien Iout 0.0675f
C2732 XA.XIR[11].XIC[5].icell.Ien Vbias 0.19161f
C2733 XThR.Tn[2] XA.XIR[2].XIC[12].icell.Ien 0.14211f
C2734 XThC.XTBN.Y a_7875_9569# 0.229f
C2735 XThR.Tn[13] XA.XIR[13].XIC[11].icell.Ien 0.14211f
C2736 XA.XIR[10].XIC[7].icell.Ien Vbias 0.19161f
C2737 XA.XIR[8].XIC[0].icell.PDM VPWR 0.01171f
C2738 XA.XIR[4].XIC[11].icell.Ien VPWR 0.18829f
C2739 XThC.XTB2.Y XThC.XTBN.Y 0.2075f
C2740 XA.XIR[1].XIC_dummy_left.icell.Ien XA.XIR[2].XIC_dummy_left.icell.PDM 0.02104f
C2741 XThC.Tn[5] XThR.Tn[2] 0.40741f
C2742 XThR.XTB4.Y XThR.XTB5.Y 2.06459f
C2743 XA.XIR[12].XIC[10].icell.Ien Iout 0.06801f
C2744 XA.XIR[11].XIC[13].icell.PDM VPWR 0.01171f
C2745 XA.XIR[2].XIC[4].icell.PDM VPWR 0.01171f
C2746 XA.XIR[8].XIC[5].icell.Ien VPWR 0.18829f
C2747 XThC.Tn[14] XThR.Tn[14] 0.40742f
C2748 XA.XIR[7].XIC[11].icell.Ien Iout 0.06801f
C2749 XThR.Tn[2] XA.XIR[3].XIC_dummy_left.icell.Iout 0.01728f
C2750 XThR.XTB5.Y XThR.Tn[10] 0.01742f
C2751 XA.XIR[5].XIC[2].icell.PDM XA.XIR[5].XIC[2].icell.Ien 0.04854f
C2752 XThC.Tn[13] XA.XIR[7].XIC[13].icell.Ien 0.04604f
C2753 XA.XIR[12].XIC[1].icell.PDM XA.XIR[12].XIC[1].icell.Ien 0.04854f
C2754 XA.XIR[14].XIC[14].icell.PDM VPWR 0.0118f
C2755 XThR.Tn[11] XA.XIR[12].XIC[4].icell.PDM 0.04035f
C2756 XA.XIR[2].XIC[9].icell.Ien Vbias 0.19161f
C2757 XA.XIR[9].XIC_dummy_right.icell.Iout Iout 0.01732f
C2758 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[0].XIC_dummy_right.icell.Iout 0.06446f
C2759 XA.XIR[3].XIC[0].icell.Ien Iout 0.06795f
C2760 XA.XIR[9].XIC[14].icell.Ien VPWR 0.18835f
C2761 XThR.Tn[8] Iout 1.12761f
C2762 XA.XIR[13].XIC_15.icell.Ien XA.XIR[14].XIC_15.icell.PDM 0.02104f
C2763 XA.XIR[1].XIC[11].icell.Ien Vbias 0.19173f
C2764 XThC.Tn[0] XA.XIR[9].XIC[0].icell.PDM 0.02601f
C2765 XThR.Tn[9] XA.XIR[9].XIC[10].icell.Ien 0.14211f
C2766 XThR.XTB1.Y XThR.XTBN.Y 0.20262f
C2767 XA.XIR[0].XIC[12].icell.PDM XA.XIR[0].XIC[12].icell.Ien 0.04854f
C2768 XA.XIR[0].XIC[7].icell.Ien VPWR 0.18776f
C2769 XThC.Tn[1] XThR.Tn[6] 0.40738f
C2770 XA.XIR[11].XIC[1].icell.Ien Iout 0.06801f
C2771 XThR.Tn[0] XA.XIR[1].XIC[2].icell.PDM 0.04035f
C2772 data[5] data[4] 0.64735f
C2773 XThC.Tn[4] XA.XIR[15].XIC[4].icell.Ien 0.04292f
C2774 XThC.XTBN.A XThC.Tn[12] 0.22871f
C2775 XA.XIR[11].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2776 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[15].XIC_dummy_right.icell.PDM 0.02104f
C2777 XThR.Tn[1] XA.XIR[2].XIC[1].icell.PDM 0.04035f
C2778 XThR.Tn[5] a_n1049_5611# 0.27042f
C2779 XThC.Tn[13] XA.XIR[7].XIC[13].icell.PDM 0.02601f
C2780 XA.XIR[7].XIC[10].icell.Ien VPWR 0.18829f
C2781 XA.XIR[0].XIC_dummy_right.icell.Iout XA.XIR[1].XIC_dummy_right.icell.Iout 0.04047f
C2782 XThC.Tn[3] XThR.Tn[11] 0.40738f
C2783 XThR.XTB2.Y data[5] 0.017f
C2784 XA.XIR[14].XIC_dummy_left.icell.Ien VPWR 0.38902f
C2785 XThR.Tn[7] XA.XIR[8].XIC[6].icell.PDM 0.04035f
C2786 XA.XIR[7].XIC[3].icell.PDM Vbias 0.03928f
C2787 XThR.Tn[10] Vbias 1.39532f
C2788 XThC.Tn[5] XA.XIR[11].XIC[5].icell.Ien 0.04604f
C2789 XA.XIR[15].XIC[14].icell.Ien Iout 0.07192f
C2790 XThC.Tn[9] XA.XIR[6].XIC[9].icell.Ien 0.04604f
C2791 XA.XIR[6].XIC[10].icell.PDM Vbias 0.03928f
C2792 XA.XIR[15].XIC[1].icell.PDM Vbias 0.03928f
C2793 XThR.XTB1.Y XThR.XTB4.Y 0.05121f
C2794 XA.XIR[5].XIC[11].icell.Ien XA.XIR[6].XIC[11].icell.PDM 0.02104f
C2795 XA.XIR[0].XIC_dummy_right.icell.PDM XA.XIR[0].XIC_dummy_right.icell.Ien 0.04854f
C2796 XThR.Tn[6] XA.XIR[6].XIC[0].icell.Ien 0.14211f
C2797 XThC.Tn[14] XA.XIR[13].XIC[14].icell.Ien 0.04604f
C2798 XA.XIR[8].XIC[0].icell.Ien VPWR 0.18829f
C2799 XThC.Tn[9] Vbias 0.79809f
C2800 XA.XIR[14].XIC[7].icell.PDM Vbias 0.03928f
C2801 XThC.XTB5.Y XThC.Tn[4] 0.20108f
C2802 XThC.Tn[12] XA.XIR[14].XIC[12].icell.Ien 0.04604f
C2803 XThR.Tn[11] XA.XIR[11].XIC[6].icell.Ien 0.14211f
C2804 XA.XIR[14].XIC[4].icell.PDM XA.XIR[14].XIC[4].icell.Ien 0.04854f
C2805 XThR.Tn[3] XA.XIR[4].XIC[7].icell.PDM 0.04035f
C2806 XThC.Tn[2] XA.XIR[14].XIC[2].icell.PDM 0.02601f
C2807 XA.XIR[7].XIC[4].icell.PDM VPWR 0.01171f
C2808 XThC.Tn[6] XThR.Tn[1] 0.40744f
C2809 XThR.XTB6.A XThR.XTB7.A 0.44014f
C2810 XA.XIR[12].XIC_dummy_left.icell.Iout XA.XIR[13].XIC_dummy_left.icell.Iout 0.03665f
C2811 XThC.Tn[10] XThR.Tn[9] 0.40738f
C2812 XA.XIR[3].XIC[8].icell.Ien Iout 0.06801f
C2813 XA.XIR[15].XIC[2].icell.PDM VPWR 0.01512f
C2814 XA.XIR[6].XIC[11].icell.PDM VPWR 0.01171f
C2815 XThR.Tn[0] XA.XIR[0].XIC[11].icell.Ien 0.14211f
C2816 XThC.Tn[6] XThR.Tn[12] 0.40738f
C2817 XThC.Tn[1] XA.XIR[5].XIC[1].icell.PDM 0.02601f
C2818 XThR.Tn[6] XA.XIR[6].XIC[5].icell.Ien 0.14211f
C2819 XA.XIR[14].XIC[8].icell.PDM VPWR 0.01171f
C2820 XA.XIR[14].XIC_dummy_left.icell.PDM XA.XIR[14].XIC_dummy_left.icell.Ien 0.04854f
C2821 XThR.XTB5.Y a_n997_1803# 0.06458f
C2822 XA.XIR[13].XIC_dummy_right.icell.Iout XA.XIR[14].XIC_dummy_right.icell.Iout 0.04047f
C2823 XA.XIR[1].XIC[4].icell.PDM Vbias 0.03928f
C2824 XA.XIR[6].XIC[11].icell.Ien Vbias 0.19161f
C2825 XA.XIR[1].XIC[3].icell.Ien Iout 0.06801f
C2826 XThR.Tn[7] XA.XIR[7].XIC[12].icell.Ien 0.14211f
C2827 XThC.XTBN.Y XThC.Tn[4] 0.49752f
C2828 XThC.Tn[1] XThR.Tn[4] 0.40738f
C2829 XA.XIR[9].XIC[0].icell.PDM VPWR 0.01171f
C2830 XA.XIR[4].XIC[4].icell.PDM Vbias 0.03928f
C2831 XA.XIR[12].XIC_15.icell.Ien Iout 0.0694f
C2832 XA.XIR[8].XIC[11].icell.Ien Iout 0.06801f
C2833 XA.XIR[8].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2834 XA.XIR[3].XIC[12].icell.PDM Vbias 0.03928f
C2835 XThC.Tn[11] XA.XIR[14].XIC[11].icell.PDM 0.02601f
C2836 XA.XIR[14].XIC[5].icell.Ien Vbias 0.19161f
C2837 XA.XIR[8].XIC[14].icell.PDM Vbias 0.03928f
C2838 XThC.Tn[5] XThR.Tn[10] 0.40738f
C2839 XThC.Tn[0] XA.XIR[5].XIC[0].icell.Ien 0.04604f
C2840 XThC.Tn[13] XA.XIR[8].XIC[13].icell.Ien 0.04604f
C2841 XA.XIR[11].XIC[12].icell.PDM VPWR 0.01171f
C2842 XA.XIR[0].XIC[5].icell.PDM XA.XIR[0].XIC[5].icell.Ien 0.04854f
C2843 XA.XIR[13].XIC[7].icell.Ien Vbias 0.19161f
C2844 XA.XIR[3].XIC[7].icell.Ien VPWR 0.18829f
C2845 XA.XIR[1].XIC[5].icell.PDM VPWR 0.01171f
C2846 XA.XIR[12].XIC[14].icell.PDM XA.XIR[12].XIC[14].icell.Ien 0.04854f
C2847 XA.XIR[14].XIC[13].icell.PDM VPWR 0.01171f
C2848 XA.XIR[15].XIC[12].icell.Ien Iout 0.07192f
C2849 XA.XIR[0].XIC[13].icell.Ien Iout 0.0675f
C2850 XA.XIR[4].XIC[5].icell.PDM VPWR 0.01171f
C2851 XThR.Tn[13] XA.XIR[14].XIC[1].icell.PDM 0.04035f
C2852 XA.XIR[1].XIC[2].icell.Ien VPWR 0.18829f
C2853 XA.XIR[8].XIC_15.icell.PDM VPWR 0.07527f
C2854 XA.XIR[3].XIC[13].icell.PDM VPWR 0.01171f
C2855 XA.XIR[12].XIC_dummy_right.icell.Iout Iout 0.01732f
C2856 XThC.Tn[7] XA.XIR[2].XIC[7].icell.Ien 0.04605f
C2857 XThR.Tn[8] XA.XIR[9].XIC[4].icell.PDM 0.04035f
C2858 XA.XIR[5].XIC[4].icell.Ien XA.XIR[6].XIC[4].icell.PDM 0.02104f
C2859 XThR.Tn[12] XA.XIR[13].XIC[9].icell.PDM 0.04035f
C2860 XA.XIR[8].XIC[10].icell.Ien VPWR 0.18829f
C2861 XA.XIR[14].XIC[1].icell.Ien Iout 0.06801f
C2862 XA.XIR[2].XIC[14].icell.Ien Vbias 0.19161f
C2863 XA.XIR[14].XIC_dummy_left.icell.PUM VPWR 0.01604f
C2864 XA.XIR[14].XIC_dummy_right.icell.Ien VPWR 0.35722f
C2865 XThR.Tn[5] XA.XIR[6].XIC[1].icell.PDM 0.04035f
C2866 XA.XIR[7].XIC[13].icell.Ien XA.XIR[8].XIC[13].icell.PDM 0.02104f
C2867 XA.XIR[2].XIC[12].icell.Ien XA.XIR[3].XIC[12].icell.PDM 0.02104f
C2868 XA.XIR[14].XIC[0].icell.Ien Vbias 0.19149f
C2869 XThC.Tn[3] XThR.Tn[14] 0.40738f
C2870 XThC.Tn[8] XA.XIR[6].XIC[8].icell.PDM 0.02601f
C2871 XThR.Tn[9] XA.XIR[9].XIC_15.icell.Ien 0.13564f
C2872 XA.XIR[0].XIC[12].icell.Ien VPWR 0.1902f
C2873 XA.XIR[6].XIC[3].icell.Ien Iout 0.06801f
C2874 XThC.Tn[5] XA.XIR[14].XIC[5].icell.Ien 0.04604f
C2875 XThR.Tn[13] Vbias 1.39532f
C2876 XThC.XTB7.A a_5155_9615# 0.02287f
C2877 XA.XIR[13].XIC[12].icell.Ien XA.XIR[14].XIC[12].icell.PDM 0.02104f
C2878 XA.XIR[1].XIC_15.icell.Ien XA.XIR[2].XIC_15.icell.PDM 0.02104f
C2879 XThR.XTB5.A data[4] 0.14415f
C2880 XThR.Tn[6] XA.XIR[7].XIC[0].icell.PDM 0.04039f
C2881 XA.XIR[7].XIC_15.icell.Ien VPWR 0.26829f
C2882 XA.XIR[2].XIC_15.icell.PUM VPWR 0.01655f
C2883 XThR.Tn[13] XA.XIR[13].XIC[5].icell.Ien 0.14211f
C2884 XA.XIR[5].XIC[0].icell.Ien VPWR 0.18829f
C2885 XA.XIR[11].XIC[3].icell.Ien XA.XIR[12].XIC[3].icell.PDM 0.02104f
C2886 XThR.XTB5.A XThR.XTB2.Y 0.02203f
C2887 XThR.XTB7.B XThR.XTB6.A 1.47641f
C2888 XA.XIR[5].XIC[4].icell.Ien Vbias 0.19161f
C2889 XA.XIR[6].XIC[13].icell.PDM XA.XIR[6].XIC[13].icell.Ien 0.04854f
C2890 XA.XIR[4].XIC_dummy_left.icell.Iout VPWR 0.10954f
C2891 XA.XIR[2].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.PDM 0.02104f
C2892 XThC.Tn[14] VPWR 4.55561f
C2893 XThC.XTBN.Y a_6243_9615# 0.07767f
C2894 XThC.Tn[13] XA.XIR[10].XIC[13].icell.PDM 0.02601f
C2895 XA.XIR[2].XIC[1].icell.Ien Iout 0.06801f
C2896 XA.XIR[10].XIC[6].icell.Ien XA.XIR[11].XIC[6].icell.PDM 0.02104f
C2897 XA.XIR[7].XIC_dummy_left.icell.Iout Iout 0.03553f
C2898 XA.XIR[11].XIC[2].icell.Ien Iout 0.06801f
C2899 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[3].XIC_dummy_right.icell.Iout 0.06446f
C2900 XA.XIR[15].XIC[10].icell.Ien Iout 0.07192f
C2901 XA.XIR[10].XIC[7].icell.PDM XA.XIR[10].XIC[7].icell.Ien 0.04854f
C2902 XThR.Tn[8] XThR.Tn[9] 0.10569f
C2903 XA.XIR[9].XIC_dummy_left.icell.PDM VPWR 0.08221f
C2904 XA.XIR[10].XIC[4].icell.Ien Iout 0.06801f
C2905 XA.XIR[6].XIC[2].icell.Ien VPWR 0.18829f
C2906 XA.XIR[9].XIC[14].icell.PDM Vbias 0.03928f
C2907 XA.XIR[0].XIC[6].icell.PDM Vbias 0.03945f
C2908 XA.XIR[7].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2909 XThC.XTB7.A XThC.XTB6.Y 0.19112f
C2910 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Ien 0.01546f
C2911 XA.XIR[10].XIC_dummy_left.icell.Ien XThR.Tn[10] 0.01244f
C2912 XA.XIR[3].XIC[13].icell.Ien Iout 0.06801f
C2913 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Ien 0.01597f
C2914 XA.XIR[11].XIC[11].icell.PDM VPWR 0.01171f
C2915 XThC.Tn[7] Vbias 0.82088f
C2916 VPWR data[6] 0.21221f
C2917 XThR.Tn[6] XA.XIR[6].XIC[10].icell.Ien 0.14211f
C2918 XA.XIR[2].XIC[6].icell.Ien Iout 0.06801f
C2919 XA.XIR[10].XIC[10].icell.Ien XA.XIR[11].XIC[10].icell.PDM 0.02104f
C2920 XThC.Tn[5] XThR.Tn[13] 0.40738f
C2921 XA.XIR[14].XIC[12].icell.PDM VPWR 0.01171f
C2922 XA.XIR[1].XIC[8].icell.Ien Iout 0.06801f
C2923 XA.XIR[9].XIC_15.icell.PDM VPWR 0.07527f
C2924 XA.XIR[0].XIC[7].icell.PDM VPWR 0.01132f
C2925 XA.XIR[2].XIC_dummy_left.icell.PDM XA.XIR[2].XIC_dummy_left.icell.Ien 0.04854f
C2926 XA.XIR[7].XIC[14].icell.PDM XA.XIR[7].XIC[14].icell.Ien 0.04854f
C2927 XThC.Tn[4] XThR.Tn[8] 0.40738f
C2928 XA.XIR[10].XIC[3].icell.Ien VPWR 0.18829f
C2929 XA.XIR[2].XIC[5].icell.Ien XA.XIR[3].XIC[5].icell.PDM 0.02104f
C2930 XA.XIR[4].XIC_15.icell.PDM XA.XIR[4].XIC_15.icell.Ien 0.04854f
C2931 XA.XIR[7].XIC[6].icell.Ien XA.XIR[8].XIC[6].icell.PDM 0.02104f
C2932 bias[2] bias[0] 0.04602f
C2933 XThR.Tn[10] XA.XIR[11].XIC[3].icell.PDM 0.04035f
C2934 XThR.Tn[4] XA.XIR[5].XIC[14].icell.PDM 0.04056f
C2935 XThC.XTB7.A XThC.XTB4.Y 0.14536f
C2936 XThR.Tn[14] XA.XIR[15].XIC[4].icell.PDM 0.04035f
C2937 XA.XIR[3].XIC[12].icell.Ien VPWR 0.18829f
C2938 XA.XIR[1].XIC[8].icell.Ien XA.XIR[2].XIC[8].icell.PDM 0.02104f
C2939 XA.XIR[8].XIC[13].icell.PDM XA.XIR[8].XIC[13].icell.Ien 0.04854f
C2940 XA.XIR[12].XIC_15.icell.PDM XA.XIR[12].XIC_15.icell.Ien 0.04854f
C2941 XA.XIR[2].XIC[5].icell.Ien VPWR 0.18829f
C2942 XA.XIR[0].XIC[12].icell.Ien XA.XIR[1].XIC[12].icell.PDM 0.02104f
C2943 XThC.XTB6.Y a_5949_9615# 0.26831f
C2944 XA.XIR[1].XIC[7].icell.Ien VPWR 0.18829f
C2945 XThR.Tn[8] XA.XIR[8].XIC[2].icell.Ien 0.14211f
C2946 XA.XIR[6].XIC[6].icell.PDM XA.XIR[6].XIC[6].icell.Ien 0.04854f
C2947 XThC.Tn[6] XA.XIR[0].XIC[6].icell.Ien 0.04659f
C2948 XThC.Tn[1] XThC.Tn[2] 0.71417f
C2949 XThR.Tn[0] XA.XIR[0].XIC_dummy_left.icell.Iout 0.03838f
C2950 a_3773_9615# Vbias 0.01444f
C2951 XThC.Tn[3] XA.XIR[6].XIC[3].icell.PDM 0.02601f
C2952 XA.XIR[15].XIC[5].icell.PDM XA.XIR[15].XIC[5].icell.Ien 0.04854f
C2953 XA.XIR[8].XIC_15.icell.Ien VPWR 0.26829f
C2954 XThR.Tn[3] Iout 1.12764f
C2955 XThR.Tn[1] XA.XIR[1].XIC[1].icell.Ien 0.14211f
C2956 XThC.Tn[10] XA.XIR[2].XIC[10].icell.PDM 0.02602f
C2957 XThC.Tn[0] XA.XIR[3].XIC[0].icell.PDM 0.02601f
C2958 XA.XIR[5].XIC[4].icell.PDM Vbias 0.03928f
C2959 XThR.XTB7.A a_n1049_5317# 0.02018f
C2960 XA.XIR[9].XIC[5].icell.Ien XA.XIR[10].XIC[5].icell.PDM 0.02104f
C2961 XThR.XTBN.Y XThR.XTB6.A 0.03867f
C2962 XA.XIR[12].XIC[3].icell.PDM Vbias 0.03928f
C2963 XA.XIR[8].XIC_dummy_left.icell.Iout Iout 0.03553f
C2964 XA.XIR[0].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.PDM 0.02104f
C2965 a_4067_9615# VPWR 0.70663f
C2966 XA.XIR[11].XIC[9].icell.PDM Vbias 0.03928f
C2967 XA.XIR[15].XIC_15.icell.Ien Iout 0.0733f
C2968 a_n997_3755# XThR.Tn[9] 0.19352f
C2969 XThR.XTB2.Y XThR.Tn[9] 0.292f
C2970 XA.XIR[6].XIC[8].icell.Ien Iout 0.06801f
C2971 XThR.Tn[2] XA.XIR[3].XIC[8].icell.PDM 0.04035f
C2972 XThC.XTB7.Y XThC.Tn[9] 0.07413f
C2973 XThR.Tn[1] XA.XIR[1].XIC[6].icell.Ien 0.14211f
C2974 XThR.Tn[14] XA.XIR[14].XIC[6].icell.Ien 0.14211f
C2975 XThC.Tn[11] XA.XIR[12].XIC[11].icell.Ien 0.04604f
C2976 XA.XIR[5].XIC[5].icell.PDM VPWR 0.01171f
C2977 XThR.XTBN.Y XThR.Tn[0] 0.55717f
C2978 XA.XIR[8].XIC_dummy_right.icell.Iout VPWR 0.11567f
C2979 XThC.Tn[13] XA.XIR[13].XIC[13].icell.PDM 0.02601f
C2980 XA.XIR[14].XIC[2].icell.Ien Iout 0.06801f
C2981 XA.XIR[6].XIC_15.icell.Ien XA.XIR[7].XIC_15.icell.PDM 0.02104f
C2982 XThR.XTB6.A XThR.XTB4.Y 0.04137f
C2983 XA.XIR[12].XIC[4].icell.PDM VPWR 0.01171f
C2984 XA.XIR[5].XIC[9].icell.Ien Vbias 0.19161f
C2985 XA.XIR[13].XIC[4].icell.Ien Iout 0.06801f
C2986 XA.XIR[9].XIC[9].icell.PDM XA.XIR[9].XIC[9].icell.Ien 0.04854f
C2987 XA.XIR[7].XIC[7].icell.PDM XA.XIR[7].XIC[7].icell.Ien 0.04854f
C2988 XThC.Tn[1] XA.XIR[4].XIC[1].icell.Ien 0.04604f
C2989 XA.XIR[11].XIC[10].icell.PDM VPWR 0.01171f
C2990 XA.XIR[8].XIC[1].icell.PDM Vbias 0.03928f
C2991 XThC.XTB2.Y XThC.XTB7.A 0.2319f
C2992 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[13].XIC_dummy_left.icell.PDM 0.02104f
C2993 XThC.XTB5.A XThC.XTB4.Y 0.02767f
C2994 XA.XIR[4].XIC[8].icell.PDM XA.XIR[4].XIC[8].icell.Ien 0.04854f
C2995 XA.XIR[2].XIC[5].icell.PDM Vbias 0.03928f
C2996 XA.XIR[15].XIC_dummy_right.icell.Iout Iout 0.01732f
C2997 XA.XIR[11].XIC[7].icell.Ien Iout 0.06801f
C2998 XA.XIR[14].XIC[11].icell.PDM VPWR 0.01171f
C2999 XThR.Tn[9] XA.XIR[10].XIC[2].icell.PDM 0.04035f
C3000 XA.XIR[12].XIC[4].icell.Ien Vbias 0.19161f
C3001 XA.XIR[10].XIC[9].icell.Ien Iout 0.06801f
C3002 XThC.XTB1.Y XThC.Tn[1] 0.01068f
C3003 XA.XIR[6].XIC[7].icell.Ien VPWR 0.18829f
C3004 XA.XIR[8].XIC[6].icell.PDM XA.XIR[8].XIC[6].icell.Ien 0.04854f
C3005 XThR.XTB7.A a_n1049_6405# 0.02287f
C3006 XThC.Tn[3] VPWR 3.60513f
C3007 XThC.XTBN.Y a_8963_9569# 0.22784f
C3008 XThC.XTB7.A data[1] 0.06544f
C3009 XThC.Tn[10] XA.XIR[7].XIC[10].icell.PDM 0.02601f
C3010 XA.XIR[0].XIC[5].icell.Ien XA.XIR[1].XIC[5].icell.PDM 0.02104f
C3011 XA.XIR[3].XIC[0].icell.PDM VPWR 0.01171f
C3012 XA.XIR[8].XIC[2].icell.PDM VPWR 0.01171f
C3013 XA.XIR[4].XIC_dummy_left.icell.Iout XA.XIR[5].XIC_dummy_left.icell.Iout 0.03665f
C3014 XThC.Tn[9] XThR.Tn[0] 0.40759f
C3015 XThC.Tn[11] XThR.Tn[5] 0.40738f
C3016 XThR.Tn[6] XA.XIR[6].XIC_15.icell.Ien 0.13564f
C3017 XThR.Tn[1] XThR.Tn[2] 0.15279f
C3018 XThC.Tn[6] XA.XIR[3].XIC[6].icell.Ien 0.04604f
C3019 XA.XIR[2].XIC[6].icell.PDM VPWR 0.01171f
C3020 XA.XIR[8].XIC[13].icell.Ien XA.XIR[9].XIC[13].icell.PDM 0.02104f
C3021 XA.XIR[13].XIC[3].icell.Ien VPWR 0.18829f
C3022 XA.XIR[2].XIC[11].icell.Ien Iout 0.06801f
C3023 XThR.XTB1.Y a_n997_3979# 0.06353f
C3024 XA.XIR[3].XIC[12].icell.Ien XA.XIR[4].XIC[12].icell.PDM 0.02104f
C3025 XThC.Tn[13] XA.XIR[2].XIC[13].icell.Ien 0.04605f
C3026 XA.XIR[1].XIC[13].icell.Ien Iout 0.06801f
C3027 XA.XIR[3].XIC[14].icell.PDM XA.XIR[3].XIC[14].icell.Ien 0.04854f
C3028 XA.XIR[11].XIC[6].icell.Ien VPWR 0.18829f
C3029 XA.XIR[9].XIC_dummy_left.icell.Ien VPWR 0.38914f
C3030 XThR.Tn[11] XA.XIR[12].XIC[6].icell.PDM 0.04035f
C3031 XA.XIR[10].XIC[8].icell.Ien VPWR 0.18829f
C3032 XA.XIR[12].XIC[0].icell.Ien Iout 0.06795f
C3033 XThR.Tn[11] Iout 1.12764f
C3034 XThR.XTB7.B a_n1049_5317# 0.01743f
C3035 XThR.Tn[0] XA.XIR[1].XIC[4].icell.PDM 0.04035f
C3036 XThC.Tn[5] XA.XIR[2].XIC[5].icell.PDM 0.02602f
C3037 XA.XIR[3].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.PDM 0.02104f
C3038 XA.XIR[3].XIC[1].icell.PDM XA.XIR[3].XIC[1].icell.Ien 0.04854f
C3039 XThR.Tn[1] XA.XIR[2].XIC[3].icell.PDM 0.04035f
C3040 XThR.Tn[7] Vbias 1.39526f
C3041 XThR.Tn[5] XA.XIR[5].XIC[1].icell.Ien 0.14211f
C3042 XThR.Tn[11] XA.XIR[11].XIC_dummy_left.icell.Iout 0.03385f
C3043 XA.XIR[2].XIC[10].icell.Ien VPWR 0.18829f
C3044 XA.XIR[6].XIC[8].icell.Ien XA.XIR[7].XIC[8].icell.PDM 0.02104f
C3045 XThC.XTB5.A XThC.XTB2.Y 0.02203f
C3046 XThC.Tn[8] XThR.Tn[2] 0.40741f
C3047 XA.XIR[1].XIC[12].icell.Ien VPWR 0.18829f
C3048 XThR.Tn[8] XA.XIR[8].XIC[7].icell.Ien 0.14211f
C3049 XA.XIR[7].XIC[5].icell.PDM Vbias 0.03928f
C3050 XThR.Tn[7] XA.XIR[8].XIC[8].icell.PDM 0.04035f
C3051 XA.XIR[9].XIC[2].icell.PDM XA.XIR[9].XIC[2].icell.Ien 0.04854f
C3052 XA.XIR[12].XIC[12].icell.PDM XA.XIR[12].XIC[12].icell.Ien 0.04854f
C3053 XThC.Tn[14] XA.XIR[0].XIC[14].icell.PDM 0.02792f
C3054 XA.XIR[15].XIC[3].icell.PDM Vbias 0.03928f
C3055 XA.XIR[4].XIC[2].icell.Ien Vbias 0.19161f
C3056 XA.XIR[6].XIC[12].icell.PDM Vbias 0.03928f
C3057 XA.XIR[14].XIC[9].icell.PDM Vbias 0.03928f
C3058 XA.XIR[14].XIC[3].icell.Ien XA.XIR[15].XIC[3].icell.PDM 0.02104f
C3059 XThC.XTB5.A data[1] 0.11102f
C3060 XThC.XTB7.A XThC.Tn[4] 0.02779f
C3061 XThC.Tn[7] XA.XIR[10].XIC[7].icell.PDM 0.02601f
C3062 XThC.Tn[4] XA.XIR[10].XIC[4].icell.Ien 0.04604f
C3063 XA.XIR[4].XIC_15.icell.Ien XA.XIR[5].XIC_15.icell.PDM 0.02104f
C3064 XThR.Tn[3] XA.XIR[4].XIC[9].icell.PDM 0.04035f
C3065 XThR.Tn[5] XA.XIR[5].XIC[6].icell.Ien 0.14211f
C3066 XA.XIR[9].XIC[1].icell.PDM Vbias 0.03928f
C3067 XA.XIR[7].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3068 XThR.XTB6.Y XThR.XTBN.A 0.06405f
C3069 XThR.XTBN.Y XThR.Tn[1] 0.61094f
C3070 XA.XIR[7].XIC[6].icell.PDM VPWR 0.01171f
C3071 XA.XIR[13].XIC[6].icell.Ien XA.XIR[14].XIC[6].icell.PDM 0.02104f
C3072 XA.XIR[9].XIC[5].icell.Ien Vbias 0.19161f
C3073 XA.XIR[6].XIC[13].icell.PDM VPWR 0.01171f
C3074 XA.XIR[15].XIC[14].icell.PDM XA.XIR[15].XIC[14].icell.Ien 0.04854f
C3075 XA.XIR[15].XIC[4].icell.PDM VPWR 0.01512f
C3076 XA.XIR[13].XIC[7].icell.PDM XA.XIR[13].XIC[7].icell.Ien 0.04854f
C3077 XA.XIR[6].XIC[13].icell.Ien Iout 0.06801f
C3078 XThC.Tn[13] XThR.Tn[6] 0.40739f
C3079 XThC.Tn[7] XA.XIR[5].XIC[7].icell.Ien 0.04604f
C3080 VPWR data[2] 0.21031f
C3081 XA.XIR[10].XIC[14].icell.Ien Iout 0.06801f
C3082 XThR.XTBN.Y XThR.Tn[12] 0.50762f
C3083 XThR.Tn[1] XA.XIR[1].XIC[11].icell.Ien 0.14211f
C3084 XA.XIR[8].XIC[6].icell.Ien XA.XIR[9].XIC[6].icell.PDM 0.02104f
C3085 XA.XIR[12].XIC[8].icell.Ien XA.XIR[13].XIC[8].icell.PDM 0.02104f
C3086 XA.XIR[14].XIC[10].icell.PDM VPWR 0.01171f
C3087 XThC.Tn[12] XA.XIR[11].XIC[12].icell.PDM 0.02601f
C3088 XA.XIR[1].XIC[1].icell.Ien XA.XIR[2].XIC[1].icell.PDM 0.02104f
C3089 XA.XIR[3].XIC[5].icell.Ien XA.XIR[4].XIC[5].icell.PDM 0.02104f
C3090 XA.XIR[13].XIC_dummy_left.icell.Ien XThR.Tn[13] 0.01244f
C3091 XA.XIR[1].XIC[6].icell.PDM Vbias 0.03928f
C3092 VPWR bias[0] 2.91967f
C3093 XA.XIR[9].XIC[2].icell.PDM VPWR 0.01171f
C3094 XA.XIR[14].XIC[7].icell.Ien Iout 0.06801f
C3095 XA.XIR[3].XIC[7].icell.PDM XA.XIR[3].XIC[7].icell.Ien 0.04854f
C3096 XThC.Tn[5] XThR.Tn[7] 0.40738f
C3097 XA.XIR[4].XIC[6].icell.PDM Vbias 0.03928f
C3098 XThC.Tn[3] XA.XIR[7].XIC[3].icell.Ien 0.04604f
C3099 XA.XIR[5].XIC[14].icell.Ien Vbias 0.19161f
C3100 XA.XIR[13].XIC[9].icell.Ien Iout 0.06801f
C3101 XA.XIR[13].XIC[10].icell.Ien XA.XIR[14].XIC[10].icell.PDM 0.02104f
C3102 XA.XIR[12].XIC[13].icell.Ien VPWR 0.18829f
C3103 XA.XIR[3].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3104 XThC.Tn[11] Iout 0.22485f
C3105 XA.XIR[3].XIC[14].icell.PDM Vbias 0.03928f
C3106 XThC.Tn[5] XA.XIR[7].XIC[5].icell.PDM 0.02601f
C3107 XThC.XTB7.Y XThC.Tn[7] 0.08399f
C3108 XThC.XTB6.Y XThC.Tn[11] 0.02473f
C3109 XThR.XTB7.Y XThR.Tn[9] 0.07413f
C3110 XThR.Tn[4] XA.XIR[5].XIC[1].icell.PDM 0.04035f
C3111 XA.XIR[1].XIC[7].icell.PDM VPWR 0.01171f
C3112 XThR.Tn[8] XA.XIR[9].XIC_dummy_left.icell.Iout 0.01728f
C3113 XA.XIR[6].XIC[12].icell.Ien VPWR 0.18829f
C3114 XA.XIR[12].XIC[9].icell.Ien Vbias 0.19161f
C3115 XThC.Tn[9] XThR.Tn[1] 0.40744f
C3116 data[1] data[0] 0.64735f
C3117 XA.XIR[9].XIC[14].icell.Ien XA.XIR[10].XIC[14].icell.PDM 0.02104f
C3118 XA.XIR[4].XIC[7].icell.PDM VPWR 0.01171f
C3119 XA.XIR[5].XIC_15.icell.PUM VPWR 0.01655f
C3120 XThR.Tn[13] XA.XIR[14].XIC[3].icell.PDM 0.04035f
C3121 XThC.Tn[9] XThR.Tn[12] 0.40738f
C3122 XA.XIR[9].XIC[0].icell.Ien Vbias 0.19149f
C3123 XA.XIR[3].XIC_15.icell.PDM VPWR 0.07527f
C3124 XA.XIR[14].XIC[6].icell.Ien VPWR 0.18883f
C3125 XThC.Tn[5] XA.XIR[9].XIC[5].icell.Ien 0.04604f
C3126 XThR.XTBN.Y a_n1049_5317# 0.07731f
C3127 XThR.Tn[8] XA.XIR[9].XIC[6].icell.PDM 0.04035f
C3128 XA.XIR[13].XIC[8].icell.Ien VPWR 0.18829f
C3129 XThC.Tn[4] XThR.Tn[3] 0.40738f
C3130 XA.XIR[1].XIC_dummy_right.icell.Ien XA.XIR[1].XIC_dummy_right.icell.Iout 0.06446f
C3131 XThC.Tn[12] XA.XIR[0].XIC[12].icell.Ien 0.04662f
C3132 XA.XIR[5].XIC[1].icell.Ien Iout 0.06801f
C3133 XThC.Tn[13] XThR.Tn[4] 0.40739f
C3134 XThR.Tn[14] Iout 1.12763f
C3135 XThC.Tn[11] XA.XIR[15].XIC[11].icell.Ien 0.04292f
C3136 XA.XIR[1].XIC[12].icell.PDM XA.XIR[1].XIC[12].icell.Ien 0.04854f
C3137 XA.XIR[4].XIC[8].icell.Ien XA.XIR[5].XIC[8].icell.PDM 0.02104f
C3138 XThC.Tn[6] XA.XIR[1].XIC[6].icell.Ien 0.04606f
C3139 XThC.XTB4.Y XThC.Tn[11] 0.30457f
C3140 XThC.Tn[8] XThR.Tn[10] 0.40738f
C3141 XThR.Tn[0] XA.XIR[1].XIC_dummy_left.icell.Iout 0.01728f
C3142 XThC.Tn[0] XThR.Tn[5] 0.40739f
C3143 XA.XIR[7].XIC[0].icell.PDM XA.XIR[7].XIC[0].icell.Ien 0.04854f
C3144 XA.XIR[10].XIC[12].icell.Ien Iout 0.06801f
C3145 XThR.Tn[5] XA.XIR[6].XIC[3].icell.PDM 0.04035f
C3146 XThC.Tn[7] XThR.Tn[0] 0.40759f
C3147 XThC.Tn[8] XThC.Tn[9] 0.0619f
C3148 XA.XIR[4].XIC[1].icell.PDM XA.XIR[4].XIC[1].icell.Ien 0.04854f
C3149 XA.XIR[2].XIC[14].icell.PDM XA.XIR[2].XIC[14].icell.Ien 0.04854f
C3150 XThC.XTB7.A a_6243_9615# 0.02018f
C3151 XA.XIR[10].XIC[0].icell.PDM Vbias 0.03915f
C3152 XA.XIR[8].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3153 XThC.Tn[14] XA.XIR[4].XIC[14].icell.Ien 0.04604f
C3154 XA.XIR[5].XIC[6].icell.Ien Iout 0.06801f
C3155 XThR.Tn[6] XA.XIR[7].XIC[2].icell.PDM 0.04035f
C3156 XA.XIR[2].XIC_15.icell.Ien VPWR 0.26829f
C3157 XA.XIR[12].XIC[11].icell.Ien VPWR 0.18829f
C3158 XA.XIR[1].XIC_dummy_right.icell.PDM XA.XIR[1].XIC_dummy_right.icell.Ien 0.04854f
C3159 XA.XIR[15].XIC[4].icell.Ien Vbias 0.15966f
C3160 XThR.Tn[8] XA.XIR[8].XIC[12].icell.Ien 0.14211f
C3161 XThC.Tn[4] XA.XIR[13].XIC[4].icell.Ien 0.04604f
C3162 XThC.Tn[7] XA.XIR[13].XIC[7].icell.PDM 0.02601f
C3163 XA.XIR[11].XIC[5].icell.PDM XA.XIR[11].XIC[5].icell.Ien 0.04854f
C3164 XA.XIR[4].XIC[7].icell.Ien Vbias 0.19161f
C3165 XA.XIR[10].XIC[1].icell.PDM VPWR 0.01171f
C3166 XA.XIR[2].XIC_dummy_left.icell.Iout Iout 0.03553f
C3167 XThC.Tn[3] XA.XIR[8].XIC[3].icell.Ien 0.04604f
C3168 XThC.XTB7.B data[2] 0.07481f
C3169 XThR.Tn[12] a_n997_1803# 0.18719f
C3170 XThR.XTBN.Y a_n1049_6405# 0.07602f
C3171 XA.XIR[13].XIC[14].icell.Ien Iout 0.06801f
C3172 XThR.Tn[5] XA.XIR[5].XIC[11].icell.Ien 0.14211f
C3173 XThC.Tn[6] XThR.Tn[2] 0.40741f
C3174 XThC.Tn[12] XA.XIR[14].XIC[12].icell.PDM 0.02601f
C3175 XA.XIR[7].XIC[1].icell.Ien Vbias 0.19161f
C3176 XA.XIR[0].XIC[8].icell.PDM Vbias 0.03945f
C3177 XA.XIR[5].XIC[5].icell.Ien VPWR 0.18829f
C3178 XThC.XTB5.Y Vbias 0.01606f
C3179 XA.XIR[2].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3180 XA.XIR[9].XIC[10].icell.Ien Vbias 0.19161f
C3181 XA.XIR[12].XIC[14].icell.Ien Vbias 0.19161f
C3182 XA.XIR[15].XIC_15.icell.PDM XA.XIR[15].XIC_15.icell.Ien 0.04854f
C3183 XA.XIR[0].XIC[3].icell.Ien Vbias 0.19213f
C3184 XThC.Tn[6] XA.XIR[6].XIC[6].icell.Ien 0.04604f
C3185 XThC.Tn[0] XA.XIR[6].XIC[0].icell.PDM 0.02601f
C3186 XThR.XTB4.Y a_n1049_6405# 0.01546f
C3187 XThR.Tn[5] VPWR 8.03417f
C3188 XThC.Tn[12] XA.XIR[3].XIC[12].icell.Ien 0.04604f
C3189 XA.XIR[10].XIC[10].icell.Ien Iout 0.06801f
C3190 XA.XIR[0].XIC[9].icell.PDM VPWR 0.01451f
C3191 XThR.Tn[2] XA.XIR[2].XIC[0].icell.Ien 0.14251f
C3192 XA.XIR[6].XIC[1].icell.Ien XA.XIR[7].XIC[1].icell.PDM 0.02104f
C3193 XA.XIR[1].XIC[5].icell.PDM XA.XIR[1].XIC[5].icell.Ien 0.04854f
C3194 XA.XIR[11].XIC[0].icell.Ien XA.XIR[12].XIC[0].icell.PDM 0.02104f
C3195 XA.XIR[7].XIC[6].icell.Ien Vbias 0.19161f
C3196 XThC.Tn[7] XA.XIR[12].XIC[7].icell.Ien 0.04604f
C3197 XThC.Tn[10] XA.XIR[12].XIC[10].icell.PDM 0.02601f
C3198 XThC.Tn[2] XThR.Tn[6] 0.40738f
C3199 XThR.Tn[12] XThR.Tn[13] 0.11103f
C3200 XThC.XTBN.Y Vbias 0.22975f
C3201 XA.XIR[11].XIC[1].icell.PDM XA.XIR[11].XIC[1].icell.Ien 0.04854f
C3202 XA.XIR[2].XIC[7].icell.PDM XA.XIR[2].XIC[7].icell.Ien 0.04854f
C3203 XThR.Tn[10] XA.XIR[11].XIC[5].icell.PDM 0.04035f
C3204 XThC.Tn[4] XThR.Tn[11] 0.40738f
C3205 XThR.Tn[14] XA.XIR[15].XIC[6].icell.PDM 0.04035f
C3206 VPWR data[5] 0.4402f
C3207 XThC.Tn[0] Iout 0.07042f
C3208 XThC.Tn[9] XA.XIR[10].XIC[9].icell.PDM 0.02601f
C3209 XThC.Tn[10] Vbias 0.81591f
C3210 XThC.XTB5.Y XThC.Tn[5] 0.01168f
C3211 a_10915_9569# XThC.Tn[14] 0.20879f
C3212 XA.XIR[3].XIC_dummy_left.icell.Ien VPWR 0.38998f
C3213 XThC.Tn[8] XThR.Tn[13] 0.40738f
C3214 XThR.Tn[14] XA.XIR[14].XIC_dummy_left.icell.Iout 0.03385f
C3215 XA.XIR[13].XIC[12].icell.Ien Iout 0.06801f
C3216 XThR.Tn[1] XA.XIR[1].XIC_dummy_left.icell.Iout 0.03842f
C3217 XA.XIR[5].XIC[6].icell.PDM Vbias 0.03928f
C3218 XThC.Tn[7] XThR.Tn[1] 0.40744f
C3219 XThR.Tn[3] XA.XIR[3].XIC[4].icell.Ien 0.14211f
C3220 XA.XIR[5].XIC[10].icell.PDM XA.XIR[5].XIC[10].icell.Ien 0.04854f
C3221 XThC.Tn[11] XThR.Tn[9] 0.40738f
C3222 XA.XIR[9].XIC[2].icell.Ien Iout 0.06801f
C3223 XA.XIR[13].XIC[0].icell.PDM Vbias 0.03915f
C3224 XA.XIR[6].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.Iout 0.06446f
C3225 XA.XIR[12].XIC[5].icell.PDM Vbias 0.03928f
C3226 XThC.Tn[7] XThR.Tn[12] 0.40738f
C3227 XThC.Tn[14] XA.XIR[1].XIC[14].icell.PDM 0.02602f
C3228 XThC.Tn[14] XA.XIR[10].XIC[14].icell.PDM 0.02601f
C3229 XA.XIR[12].XIC[12].icell.Ien Vbias 0.19161f
C3230 XThR.Tn[11] XA.XIR[12].XIC[14].icell.PDM 0.04056f
C3231 a_5155_9615# VPWR 0.7051f
C3232 XThC.Tn[14] XA.XIR[4].XIC[14].icell.PDM 0.02601f
C3233 XA.XIR[6].XIC[0].icell.PDM VPWR 0.01171f
C3234 XThC.XTBN.Y XThC.Tn[5] 0.49425f
C3235 XThC.Tn[2] XThR.Tn[4] 0.40738f
C3236 XThR.Tn[2] XA.XIR[3].XIC[10].icell.PDM 0.04035f
C3237 XA.XIR[15].XIC[13].icell.Ien VPWR 0.31713f
C3238 XA.XIR[5].XIC[7].icell.PDM VPWR 0.01171f
C3239 XA.XIR[8].XIC[1].icell.Ien Vbias 0.19161f
C3240 XA.XIR[5].XIC[11].icell.Ien Iout 0.06801f
C3241 XA.XIR[3].XIC[3].icell.Ien Vbias 0.19161f
C3242 XA.XIR[13].XIC[1].icell.PDM VPWR 0.01171f
C3243 XThC.Tn[13] XA.XIR[5].XIC[13].icell.Ien 0.04604f
C3244 XA.XIR[12].XIC[6].icell.PDM XA.XIR[12].XIC[6].icell.Ien 0.04854f
C3245 XThC.Tn[6] XThR.Tn[10] 0.40738f
C3246 XThR.XTB5.A XThR.XTB3.Y 0.01152f
C3247 XThR.XTB7.B XThR.XTB7.A 0.35833f
C3248 XA.XIR[12].XIC[6].icell.PDM VPWR 0.01171f
C3249 XA.XIR[15].XIC[9].icell.Ien Vbias 0.15966f
C3250 XThC.Tn[13] XA.XIR[8].XIC[13].icell.PDM 0.02601f
C3251 XThC.Tn[7] XThC.Tn[8] 0.06603f
C3252 XA.XIR[3].XIC[1].icell.PDM Vbias 0.03928f
C3253 XA.XIR[8].XIC[3].icell.PDM Vbias 0.03928f
C3254 XA.XIR[4].XIC[12].icell.Ien Vbias 0.19161f
C3255 XA.XIR[12].XIC[6].icell.Ien Iout 0.06801f
C3256 XThC.Tn[9] XA.XIR[7].XIC[9].icell.Ien 0.04604f
C3257 XA.XIR[6].XIC_dummy_left.icell.Ien XA.XIR[6].XIC_dummy_left.icell.Iout 0.06446f
C3258 XA.XIR[10].XIC_15.icell.Ien Iout 0.0694f
C3259 VPWR Iout 57.8523f
C3260 XA.XIR[2].XIC[7].icell.PDM Vbias 0.03928f
C3261 XA.XIR[8].XIC[6].icell.Ien Vbias 0.19161f
C3262 XThR.Tn[9] XA.XIR[10].XIC[4].icell.PDM 0.04035f
C3263 XThC.XTB6.Y VPWR 1.03165f
C3264 XA.XIR[12].XIC[10].icell.PDM XA.XIR[12].XIC[10].icell.Ien 0.04854f
C3265 XA.XIR[4].XIC[1].icell.Ien XA.XIR[5].XIC[1].icell.PDM 0.02104f
C3266 XA.XIR[11].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3267 XThC.Tn[2] XA.XIR[2].XIC[2].icell.PDM 0.02602f
C3268 XA.XIR[5].XIC[10].icell.Ien VPWR 0.18829f
C3269 XThC.XTBN.Y a_10051_9569# 0.23006f
C3270 XA.XIR[9].XIC_15.icell.Ien Vbias 0.19195f
C3271 XThR.XTB5.Y XThR.Tn[8] 0.01728f
C3272 XThR.XTB7.A XThR.Tn[2] 0.12549f
C3273 XA.XIR[13].XIC[10].icell.Ien Iout 0.06801f
C3274 XA.XIR[3].XIC[2].icell.PDM VPWR 0.01171f
C3275 XA.XIR[11].XIC[14].icell.PDM XA.XIR[11].XIC[14].icell.Ien 0.04854f
C3276 XThC.Tn[5] XA.XIR[12].XIC[5].icell.PDM 0.02601f
C3277 XThR.Tn[4] XA.XIR[4].XIC[1].icell.Ien 0.14211f
C3278 XA.XIR[8].XIC[4].icell.PDM VPWR 0.01171f
C3279 XA.XIR[10].XIC[1].icell.Ien XThR.Tn[10] 0.14211f
C3280 XThC.Tn[10] XA.XIR[15].XIC[10].icell.PDM 0.02601f
C3281 XA.XIR[0].XIC[8].icell.Ien Vbias 0.19213f
C3282 XA.XIR[2].XIC[8].icell.PDM VPWR 0.01171f
C3283 XThR.Tn[3] XA.XIR[3].XIC[1].icell.Ien 0.14211f
C3284 XThC.Tn[11] XA.XIR[0].XIC[11].icell.PDM 0.0279f
C3285 XA.XIR[10].XIC_dummy_right.icell.Iout Iout 0.01732f
C3286 XA.XIR[12].XIC[5].icell.Ien VPWR 0.18829f
C3287 XA.XIR[5].XIC[3].icell.PDM XA.XIR[5].XIC[3].icell.Ien 0.04854f
C3288 XA.XIR[12].XIC[10].icell.Ien Vbias 0.19161f
C3289 XThC.Tn[11] XA.XIR[9].XIC[11].icell.Ien 0.04604f
C3290 XA.XIR[15].XIC[12].icell.PDM XA.XIR[15].XIC[12].icell.Ien 0.04854f
C3291 XThC.Tn[4] XThR.Tn[14] 0.40738f
C3292 XA.XIR[7].XIC[11].icell.Ien Vbias 0.19161f
C3293 XThR.Tn[11] XA.XIR[12].XIC[8].icell.PDM 0.04035f
C3294 XThC.Tn[4] XA.XIR[10].XIC[4].icell.PDM 0.02601f
C3295 XA.XIR[9].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3296 XA.XIR[15].XIC[11].icell.Ien VPWR 0.31713f
C3297 XThR.Tn[4] XA.XIR[4].XIC[6].icell.Ien 0.14211f
C3298 XThC.Tn[9] XA.XIR[13].XIC[9].icell.PDM 0.02601f
C3299 XThC.XTB4.Y VPWR 0.91479f
C3300 XThC.Tn[12] XA.XIR[1].XIC[12].icell.Ien 0.04606f
C3301 XA.XIR[0].XIC[13].icell.PDM XA.XIR[0].XIC[13].icell.Ien 0.04854f
C3302 XA.XIR[3].XIC[0].icell.Ien Vbias 0.19149f
C3303 XThR.Tn[8] Vbias 1.39526f
C3304 XThR.Tn[0] XA.XIR[1].XIC[6].icell.PDM 0.04035f
C3305 XA.XIR[8].XIC_dummy_left.icell.Iout XA.XIR[9].XIC_dummy_left.icell.Iout 0.03665f
C3306 XThC.XTB3.Y XThC.XTBN.A 0.03907f
C3307 XA.XIR[4].XIC_dummy_right.icell.Ien XA.XIR[4].XIC_dummy_right.icell.Iout 0.06446f
C3308 XThR.Tn[1] XA.XIR[2].XIC[5].icell.PDM 0.04035f
C3309 XThR.XTB5.A VPWR 0.83234f
C3310 XThR.Tn[5] XA.XIR[5].XIC_dummy_left.icell.Iout 0.03935f
C3311 XA.XIR[11].XIC[1].icell.Ien Vbias 0.19161f
C3312 XA.XIR[4].XIC[4].icell.Ien Iout 0.06801f
C3313 XA.XIR[7].XIC[7].icell.PDM Vbias 0.03928f
C3314 XThR.XTB1.Y XThR.Tn[8] 0.29191f
C3315 XThR.Tn[7] XA.XIR[8].XIC[10].icell.PDM 0.04035f
C3316 XThR.Tn[11] XA.XIR[12].XIC[13].icell.PDM 0.0404f
C3317 XA.XIR[6].XIC_dummy_left.icell.PDM VPWR 0.08221f
C3318 XA.XIR[6].XIC[14].icell.PDM Vbias 0.03928f
C3319 XA.XIR[15].XIC[5].icell.PDM Vbias 0.03928f
C3320 XA.XIR[5].XIC[12].icell.Ien XA.XIR[6].XIC[12].icell.PDM 0.02104f
C3321 XThC.Tn[14] XA.XIR[13].XIC[14].icell.PDM 0.02601f
C3322 XThR.Tn[12] XA.XIR[12].XIC[4].icell.Ien 0.14211f
C3323 XThC.Tn[2] XA.XIR[7].XIC[2].icell.PDM 0.02601f
C3324 XThR.Tn[3] XA.XIR[3].XIC[9].icell.Ien 0.14211f
C3325 XThC.Tn[13] XA.XIR[9].XIC[13].icell.PDM 0.02601f
C3326 XA.XIR[15].XIC[14].icell.Ien Vbias 0.15966f
C3327 XA.XIR[9].XIC[7].icell.Ien Iout 0.06801f
C3328 XThR.XTBN.Y XThR.XTB7.A 0.59539f
C3329 XA.XIR[14].XIC[5].icell.PDM XA.XIR[14].XIC[5].icell.Ien 0.04854f
C3330 XA.XIR[9].XIC[3].icell.PDM Vbias 0.03928f
C3331 XThR.Tn[3] XA.XIR[4].XIC[11].icell.PDM 0.04035f
C3332 XA.XIR[2].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3333 XThC.Tn[9] XA.XIR[8].XIC[9].icell.Ien 0.04604f
C3334 XA.XIR[7].XIC[8].icell.PDM VPWR 0.01171f
C3335 XThR.Tn[2] XA.XIR[2].XIC[4].icell.Ien 0.14211f
C3336 XA.XIR[9].XIC[1].icell.Ien VPWR 0.18829f
C3337 XThC.Tn[6] XThR.Tn[13] 0.40738f
C3338 XA.XIR[4].XIC[3].icell.Ien VPWR 0.18829f
C3339 XA.XIR[15].XIC[6].icell.PDM VPWR 0.01512f
C3340 XA.XIR[6].XIC_15.icell.PDM VPWR 0.07527f
C3341 XThC.Tn[7] XA.XIR[15].XIC[7].icell.Ien 0.04292f
C3342 XA.XIR[4].XIC_dummy_left.icell.Ien XA.XIR[4].XIC_dummy_left.icell.Iout 0.06446f
C3343 XA.XIR[5].XIC_dummy_right.icell.Ien XA.XIR[6].XIC_dummy_right.icell.PDM 0.02104f
C3344 XA.XIR[10].XIC_dummy_left.icell.PDM XA.XIR[10].XIC_dummy_left.icell.Ien 0.04854f
C3345 XThC.Tn[0] XThR.Tn[9] 0.40738f
C3346 XA.XIR[7].XIC[3].icell.Ien Iout 0.06801f
C3347 XThC.Tn[5] XThR.Tn[8] 0.40738f
C3348 XA.XIR[3].XIC[8].icell.Ien Vbias 0.19161f
C3349 XA.XIR[1].XIC[8].icell.PDM Vbias 0.03928f
C3350 XThR.XTB2.Y XThR.XTB5.Y 0.0451f
C3351 XThR.XTB7.A XThR.XTB4.Y 0.14536f
C3352 XA.XIR[13].XIC_15.icell.Ien Iout 0.0694f
C3353 XA.XIR[9].XIC[4].icell.PDM VPWR 0.01171f
C3354 XThC.Tn[12] XA.XIR[6].XIC[12].icell.Ien 0.04604f
C3355 XThC.Tn[3] XA.XIR[2].XIC[3].icell.Ien 0.04605f
C3356 XA.XIR[4].XIC[8].icell.PDM Vbias 0.03928f
C3357 XThC.XTB2.Y VPWR 0.97668f
C3358 XThC.XTB5.Y XThC.XTB7.Y 0.036f
C3359 XThC.XTB7.B XThC.XTB6.Y 0.30244f
C3360 XA.XIR[14].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3361 XA.XIR[9].XIC[6].icell.Ien VPWR 0.18829f
C3362 XA.XIR[1].XIC[3].icell.Ien Vbias 0.19173f
C3363 XThC.Tn[0] XA.XIR[15].XIC[0].icell.Ien 0.04292f
C3364 XThR.Tn[9] XA.XIR[9].XIC[2].icell.Ien 0.14211f
C3365 XA.XIR[12].XIC_15.icell.Ien Vbias 0.19195f
C3366 XA.XIR[0].XIC[6].icell.PDM XA.XIR[0].XIC[6].icell.Ien 0.04854f
C3367 XThC.XTB1.Y XThC.XTBN.A 0.12307f
C3368 XThC.Tn[5] XA.XIR[15].XIC[5].icell.PDM 0.02601f
C3369 XThR.Tn[4] XA.XIR[5].XIC[3].icell.PDM 0.04035f
C3370 XA.XIR[8].XIC[11].icell.Ien Vbias 0.19161f
C3371 XA.XIR[1].XIC[9].icell.PDM VPWR 0.01171f
C3372 XThC.XTB3.Y XThC.Tn[2] 0.18399f
C3373 XThC.Tn[6] XA.XIR[0].XIC[6].icell.PDM 0.02803f
C3374 XA.XIR[14].XIC[1].icell.PDM XA.XIR[14].XIC[1].icell.Ien 0.04854f
C3375 VPWR data[1] 0.44103f
C3376 XA.XIR[4].XIC[9].icell.PDM VPWR 0.01171f
C3377 XThC.Tn[14] XA.XIR[5].XIC[14].icell.PDM 0.02601f
C3378 XA.XIR[5].XIC_15.icell.Ien VPWR 0.26829f
C3379 XA.XIR[7].XIC[2].icell.Ien VPWR 0.18829f
C3380 XA.XIR[13].XIC_dummy_right.icell.Iout Iout 0.01732f
C3381 XThR.Tn[13] XA.XIR[14].XIC[5].icell.PDM 0.04035f
C3382 XThC.Tn[6] XThC.Tn[7] 0.0974f
C3383 XThC.XTB7.Y XThC.XTBN.Y 0.50018f
C3384 XA.XIR[12].XIC_15.icell.PDM VPWR 0.07527f
C3385 XA.XIR[11].XIC_15.icell.PDM XA.XIR[11].XIC_15.icell.Ien 0.04854f
C3386 XThC.Tn[4] XA.XIR[13].XIC[4].icell.PDM 0.02601f
C3387 XA.XIR[0].XIC[13].icell.Ien Vbias 0.19213f
C3388 XA.XIR[12].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3389 XA.XIR[15].XIC[12].icell.Ien Vbias 0.15966f
C3390 XThR.Tn[8] XA.XIR[9].XIC[8].icell.PDM 0.04035f
C3391 XA.XIR[5].XIC[5].icell.Ien XA.XIR[6].XIC[5].icell.PDM 0.02104f
C3392 XThR.XTB1.Y data[4] 0.06453f
C3393 XA.XIR[15].XIC[1].icell.Ien Iout 0.07192f
C3394 XThC.XTB4.Y XThC.XTB7.B 0.33064f
C3395 XA.XIR[5].XIC_dummy_left.icell.Iout Iout 0.03553f
C3396 XThC.Tn[8] XThR.Tn[7] 0.40738f
C3397 XThR.XTB1.Y XThR.XTB2.Y 2.14864f
C3398 XThC.XTB7.Y XThC.Tn[10] 0.07427f
C3399 XThR.Tn[9] VPWR 8.97014f
C3400 XThR.Tn[11] XA.XIR[12].XIC[12].icell.PDM 0.04035f
C3401 XA.XIR[5].XIC_dummy_right.icell.Iout VPWR 0.11567f
C3402 XA.XIR[2].XIC[13].icell.Ien XA.XIR[3].XIC[13].icell.PDM 0.02104f
C3403 XThR.Tn[5] XA.XIR[6].XIC[5].icell.PDM 0.04035f
C3404 XThR.Tn[4] XA.XIR[4].XIC[11].icell.Ien 0.14211f
C3405 XA.XIR[7].XIC[14].icell.Ien XA.XIR[8].XIC[14].icell.PDM 0.02104f
C3406 XA.XIR[14].XIC[1].icell.Ien Vbias 0.19161f
C3407 XThR.Tn[0] XA.XIR[0].XIC[3].icell.Ien 0.14211f
C3408 XThR.Tn[10] XA.XIR[10].XIC[2].icell.Ien 0.14211f
C3409 XA.XIR[10].XIC[2].icell.PDM Vbias 0.03928f
C3410 XA.XIR[15].XIC[6].icell.Ien Iout 0.07192f
C3411 XThR.XTB7.B XThR.XTBN.Y 0.3875f
C3412 XThR.Tn[6] XA.XIR[7].XIC[4].icell.PDM 0.04035f
C3413 XThR.Tn[14] XA.XIR[15].XIC[14].icell.PDM 0.04056f
C3414 XThR.Tn[7] XA.XIR[7].XIC[4].icell.Ien 0.14211f
C3415 XA.XIR[6].XIC[3].icell.Ien Vbias 0.19161f
C3416 XA.XIR[4].XIC[9].icell.Ien Iout 0.06801f
C3417 XA.XIR[15].XIC[0].icell.Ien VPWR 0.31713f
C3418 XA.XIR[0].XIC[0].icell.Ien Iout 0.06743f
C3419 XThC.Tn[11] XA.XIR[10].XIC[11].icell.Ien 0.04604f
C3420 XA.XIR[11].XIC[4].icell.Ien XA.XIR[12].XIC[4].icell.PDM 0.02104f
C3421 XThC.XTB1.Y XThC.XTB3.Y 0.04033f
C3422 XA.XIR[6].XIC[14].icell.PDM XA.XIR[6].XIC[14].icell.Ien 0.04854f
C3423 XA.XIR[8].XIC[3].icell.Ien Iout 0.06801f
C3424 XThC.Tn[13] XA.XIR[11].XIC[13].icell.PDM 0.02601f
C3425 XThR.Tn[12] XA.XIR[12].XIC[9].icell.Ien 0.14211f
C3426 XA.XIR[10].XIC[3].icell.PDM VPWR 0.01171f
C3427 XA.XIR[10].XIC[7].icell.Ien XA.XIR[11].XIC[7].icell.PDM 0.02104f
C3428 XThC.Tn[4] VPWR 3.6464f
C3429 XThR.Tn[3] XA.XIR[3].XIC[14].icell.Ien 0.144f
C3430 XA.XIR[10].XIC[8].icell.PDM XA.XIR[10].XIC[8].icell.Ien 0.04854f
C3431 XThR.XTB7.B XThR.XTB4.Y 0.33064f
C3432 XA.XIR[9].XIC[12].icell.Ien Iout 0.06801f
C3433 XThR.XTBN.Y XThR.Tn[2] 0.6189f
C3434 XA.XIR[2].XIC[1].icell.Ien Vbias 0.19161f
C3435 XThC.Tn[10] XThR.Tn[0] 0.40762f
C3436 XA.XIR[0].XIC[10].icell.PDM Vbias 0.03945f
C3437 XA.XIR[15].XIC[5].icell.Ien VPWR 0.31713f
C3438 XThC.Tn[12] XThR.Tn[5] 0.40738f
C3439 XA.XIR[11].XIC[2].icell.Ien Vbias 0.19161f
C3440 XA.XIR[0].XIC[5].icell.Ien Iout 0.0675f
C3441 XThR.XTB7.B XThR.Tn[10] 0.06102f
C3442 XThR.Tn[2] XA.XIR[2].XIC[9].icell.Ien 0.14211f
C3443 XThC.XTB7.B a_7875_9569# 0.01174f
C3444 XA.XIR[15].XIC[10].icell.Ien Vbias 0.15966f
C3445 XThC.XTB7.A Vbias 0.0148f
C3446 XA.XIR[10].XIC[4].icell.Ien Vbias 0.19161f
C3447 XA.XIR[4].XIC[8].icell.Ien VPWR 0.18829f
C3448 XThC.XTB2.Y XThC.XTB7.B 0.22599f
C3449 XThC.XTB6.A XThC.XTB5.Y 0.01866f
C3450 a_8963_9569# XThC.Tn[11] 0.1927f
C3451 XA.XIR[7].XIC[8].icell.Ien Iout 0.06801f
C3452 XA.XIR[8].XIC[2].icell.Ien VPWR 0.18829f
C3453 XA.XIR[3].XIC[13].icell.Ien Vbias 0.19161f
C3454 XA.XIR[14].XIC[14].icell.PDM XA.XIR[14].XIC[14].icell.Ien 0.04854f
C3455 XA.XIR[13].XIC[1].icell.Ien XThR.Tn[13] 0.14211f
C3456 XThC.Tn[2] XA.XIR[0].XIC[2].icell.Ien 0.04658f
C3457 XA.XIR[0].XIC[11].icell.PDM VPWR 0.01132f
C3458 XA.XIR[2].XIC[6].icell.Ien Vbias 0.19161f
C3459 XA.XIR[7].XIC_15.icell.PDM XA.XIR[7].XIC_15.icell.Ien 0.04854f
C3460 XA.XIR[9].XIC[11].icell.Ien VPWR 0.18829f
C3461 XA.XIR[1].XIC[8].icell.Ien Vbias 0.19173f
C3462 XA.XIR[2].XIC[6].icell.Ien XA.XIR[3].XIC[6].icell.PDM 0.02104f
C3463 XA.XIR[7].XIC[7].icell.Ien XA.XIR[8].XIC[7].icell.PDM 0.02104f
C3464 XA.XIR[12].XIC[14].icell.PDM VPWR 0.0118f
C3465 XThC.Tn[11] XA.XIR[1].XIC[11].icell.PDM 0.02602f
C3466 XThR.Tn[9] XA.XIR[9].XIC[7].icell.Ien 0.14211f
C3467 XThR.Tn[10] XA.XIR[11].XIC[7].icell.PDM 0.04035f
C3468 XA.XIR[0].XIC[4].icell.Ien VPWR 0.18788f
C3469 XThC.XTB6.A XThC.XTBN.Y 0.03867f
C3470 XThR.Tn[14] XA.XIR[15].XIC[8].icell.PDM 0.04035f
C3471 XThC.Tn[9] XThR.Tn[2] 0.40741f
C3472 XA.XIR[15].XIC_15.icell.PDM VPWR 0.07867f
C3473 XThC.Tn[11] XA.XIR[4].XIC[11].icell.PDM 0.02601f
C3474 XA.XIR[1].XIC[9].icell.Ien XA.XIR[2].XIC[9].icell.PDM 0.02104f
C3475 XA.XIR[10].XIC[0].icell.Ien Iout 0.06795f
C3476 XA.XIR[8].XIC[14].icell.PDM XA.XIR[8].XIC[14].icell.Ien 0.04854f
C3477 XA.XIR[7].XIC[7].icell.Ien VPWR 0.18829f
C3478 XThC.Tn[4] XA.XIR[4].XIC[4].icell.Ien 0.04604f
C3479 XThR.XTB5.Y XThR.XTB7.Y 0.036f
C3480 XThR.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.04035f
C3481 XA.XIR[0].XIC[13].icell.Ien XA.XIR[1].XIC[13].icell.PDM 0.02104f
C3482 XA.XIR[7].XIC_dummy_left.icell.Ien XThR.Tn[7] 0.01256f
C3483 XA.XIR[6].XIC[7].icell.PDM XA.XIR[6].XIC[7].icell.Ien 0.04854f
C3484 XThC.Tn[10] XA.XIR[8].XIC[10].icell.PDM 0.02601f
C3485 XA.XIR[15].XIC[6].icell.PDM XA.XIR[15].XIC[6].icell.Ien 0.04854f
C3486 XThC.XTB7.A XThC.Tn[5] 0.02777f
C3487 XA.XIR[6].XIC[1].icell.PDM Vbias 0.03928f
C3488 XA.XIR[12].XIC_dummy_left.icell.Ien VPWR 0.38922f
C3489 XA.XIR[5].XIC[8].icell.PDM Vbias 0.03928f
C3490 XA.XIR[11].XIC[12].icell.PDM XA.XIR[11].XIC[12].icell.Ien 0.04854f
C3491 XA.XIR[9].XIC[6].icell.Ien XA.XIR[10].XIC[6].icell.PDM 0.02104f
C3492 XThR.Tn[14] XA.XIR[15].XIC[13].icell.PDM 0.0404f
C3493 XA.XIR[13].XIC[2].icell.PDM Vbias 0.03928f
C3494 XThR.Tn[11] XA.XIR[11].XIC[3].icell.Ien 0.14211f
C3495 XThR.Tn[3] Vbias 1.39527f
C3496 XThC.Tn[14] XA.XIR[11].XIC[14].icell.Ien 0.04604f
C3497 XThC.Tn[14] XThR.Tn[6] 0.40742f
C3498 XA.XIR[12].XIC[7].icell.PDM Vbias 0.03928f
C3499 XThR.Tn[12] XA.XIR[12].XIC[14].icell.Ien 0.144f
C3500 a_6243_9615# VPWR 0.7055f
C3501 XA.XIR[12].XIC_dummy_left.icell.Iout Iout 0.03553f
C3502 XThR.Tn[0] XA.XIR[0].XIC[8].icell.Ien 0.14211f
C3503 XA.XIR[3].XIC[5].icell.Ien Iout 0.06801f
C3504 XA.XIR[6].XIC[2].icell.PDM VPWR 0.01171f
C3505 XThC.Tn[11] XA.XIR[13].XIC[11].icell.Ien 0.04604f
C3506 XThR.Tn[10] XA.XIR[10].XIC[7].icell.Ien 0.14211f
C3507 XThR.Tn[2] XA.XIR[3].XIC[12].icell.PDM 0.04035f
C3508 XA.XIR[15].XIC[10].icell.PDM XA.XIR[15].XIC[10].icell.Ien 0.04854f
C3509 XA.XIR[5].XIC_dummy_left.icell.PDM XA.XIR[5].XIC_dummy_left.icell.Ien 0.04854f
C3510 XThR.Tn[6] XA.XIR[6].XIC[2].icell.Ien 0.14211f
C3511 XThC.Tn[2] XA.XIR[12].XIC[2].icell.PDM 0.02601f
C3512 XA.XIR[5].XIC[9].icell.PDM VPWR 0.01171f
C3513 XThR.XTBN.Y XThR.XTB4.Y 0.15627f
C3514 XThC.Tn[13] XA.XIR[14].XIC[13].icell.PDM 0.02601f
C3515 XThC.Tn[6] XThR.Tn[7] 0.40738f
C3516 XA.XIR[11].XIC_dummy_left.icell.Iout XA.XIR[12].XIC_dummy_left.icell.Iout 0.03665f
C3517 XThC.Tn[12] Iout 0.2243f
C3518 XA.XIR[15].XIC_15.icell.Ien Vbias 0.15966f
C3519 XA.XIR[13].XIC[3].icell.PDM VPWR 0.01171f
C3520 XA.XIR[6].XIC[8].icell.Ien Vbias 0.19161f
C3521 XThC.Tn[8] XA.XIR[0].XIC[8].icell.PDM 0.02805f
C3522 XA.XIR[4].XIC[14].icell.Ien Iout 0.06801f
C3523 XThR.Tn[7] XA.XIR[7].XIC[9].icell.Ien 0.14211f
C3524 XThR.XTBN.Y XThR.Tn[10] 0.46535f
C3525 XThC.XTB5.Y XThC.Tn[8] 0.0173f
C3526 XA.XIR[12].XIC[8].icell.PDM VPWR 0.01171f
C3527 XThC.Tn[13] XA.XIR[3].XIC[13].icell.PDM 0.02601f
C3528 XThR.XTB1.Y XThR.XTB7.Y 0.05211f
C3529 XA.XIR[9].XIC[10].icell.PDM XA.XIR[9].XIC[10].icell.Ien 0.04854f
C3530 XA.XIR[13].XIC_dummy_left.icell.PDM XA.XIR[13].XIC_dummy_left.icell.Ien 0.04854f
C3531 XThC.XTB6.Y XThC.Tn[12] 0.0253f
C3532 XA.XIR[7].XIC[8].icell.PDM XA.XIR[7].XIC[8].icell.Ien 0.04854f
C3533 XThC.Tn[2] XA.XIR[3].XIC[2].icell.Ien 0.04604f
C3534 XA.XIR[8].XIC[8].icell.Ien Iout 0.06801f
C3535 XA.XIR[3].XIC[3].icell.PDM Vbias 0.03928f
C3536 XA.XIR[8].XIC[5].icell.PDM Vbias 0.03928f
C3537 XA.XIR[14].XIC[2].icell.Ien Vbias 0.19161f
C3538 XA.XIR[4].XIC[9].icell.PDM XA.XIR[4].XIC[9].icell.Ien 0.04854f
C3539 XThC.Tn[10] XThR.Tn[1] 0.40744f
C3540 XThC.Tn[1] XA.XIR[10].XIC[1].icell.PDM 0.02601f
C3541 XThC.Tn[9] XA.XIR[2].XIC[9].icell.Ien 0.04605f
C3542 a_5949_9615# XThC.Tn[5] 0.26251f
C3543 XA.XIR[2].XIC[9].icell.PDM Vbias 0.03928f
C3544 XA.XIR[13].XIC[4].icell.Ien Vbias 0.19161f
C3545 XA.XIR[15].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3546 XA.XIR[10].XIC[13].icell.Ien VPWR 0.18829f
C3547 XThR.Tn[9] XA.XIR[10].XIC[6].icell.PDM 0.04035f
C3548 XA.XIR[3].XIC[4].icell.Ien VPWR 0.18829f
C3549 XThC.Tn[10] XThR.Tn[12] 0.40738f
C3550 XThC.Tn[11] XA.XIR[12].XIC[11].icell.PDM 0.02601f
C3551 XA.XIR[1].XIC[2].icell.Ien XA.XIR[2].XIC[2].icell.PDM 0.02104f
C3552 XA.XIR[8].XIC[7].icell.PDM XA.XIR[8].XIC[7].icell.Ien 0.04854f
C3553 XThR.XTB4.Y XThR.Tn[10] 0.01391f
C3554 XA.XIR[0].XIC[10].icell.Ien Iout 0.0675f
C3555 XA.XIR[11].XIC[7].icell.Ien Vbias 0.19161f
C3556 XThR.Tn[2] XA.XIR[2].XIC[14].icell.Ien 0.144f
C3557 XThC.XTBN.Y XThC.Tn[8] 0.41222f
C3558 XThC.Tn[5] XThR.Tn[3] 0.40738f
C3559 XA.XIR[6].XIC_dummy_right.icell.Iout XA.XIR[7].XIC_dummy_right.icell.Iout 0.04047f
C3560 XA.XIR[0].XIC[6].icell.Ien XA.XIR[1].XIC[6].icell.PDM 0.02104f
C3561 XA.XIR[3].XIC[4].icell.PDM VPWR 0.01171f
C3562 XA.XIR[4].XIC[13].icell.Ien VPWR 0.18829f
C3563 XA.XIR[8].XIC[6].icell.PDM VPWR 0.01171f
C3564 XA.XIR[10].XIC[9].icell.Ien Vbias 0.19161f
C3565 XThR.Tn[4] XA.XIR[4].XIC_dummy_left.icell.Iout 0.03908f
C3566 XA.XIR[12].XIC[13].icell.PDM VPWR 0.01171f
C3567 XThC.XTB1.Y a_2979_9615# 0.21263f
C3568 XThC.Tn[14] XThR.Tn[4] 0.40742f
C3569 XA.XIR[8].XIC[14].icell.Ien XA.XIR[9].XIC[14].icell.PDM 0.02104f
C3570 XThR.Tn[3] XA.XIR[3].XIC_dummy_left.icell.Iout 0.03843f
C3571 XA.XIR[2].XIC[10].icell.PDM VPWR 0.01171f
C3572 XThC.Tn[6] XA.XIR[1].XIC[6].icell.PDM 0.02602f
C3573 XThR.Tn[12] XA.XIR[13].XIC[0].icell.PDM 0.04041f
C3574 XThR.XTB5.Y XThR.Tn[11] 0.02067f
C3575 XA.XIR[7].XIC[13].icell.Ien Iout 0.06801f
C3576 XA.XIR[8].XIC[7].icell.Ien VPWR 0.18829f
C3577 XA.XIR[15].XIC[14].icell.PDM VPWR 0.01521f
C3578 XThC.Tn[9] XThR.Tn[10] 0.40738f
C3579 XThC.Tn[1] XThR.Tn[5] 0.40738f
C3580 XA.XIR[3].XIC[13].icell.Ien XA.XIR[4].XIC[13].icell.PDM 0.02104f
C3581 XThC.Tn[6] XA.XIR[4].XIC[6].icell.PDM 0.02601f
C3582 XThR.Tn[12] XA.XIR[12].XIC[12].icell.Ien 0.14211f
C3583 XA.XIR[3].XIC_15.icell.PDM XA.XIR[3].XIC_15.icell.Ien 0.04854f
C3584 XA.XIR[14].XIC_15.icell.PDM XA.XIR[14].XIC_15.icell.Ien 0.04854f
C3585 XA.XIR[2].XIC[11].icell.Ien Vbias 0.19161f
C3586 XThC.Tn[10] XA.XIR[9].XIC[10].icell.PDM 0.02601f
C3587 XThR.Tn[11] XA.XIR[12].XIC[10].icell.PDM 0.04035f
C3588 XA.XIR[5].XIC_dummy_right.icell.Ien VPWR 0.35722f
C3589 XA.XIR[13].XIC[0].icell.Ien Iout 0.06795f
C3590 XThC.Tn[13] XThC.Tn[14] 0.3543f
C3591 XA.XIR[1].XIC[13].icell.Ien Vbias 0.19173f
C3592 XThR.Tn[9] XA.XIR[9].XIC[12].icell.Ien 0.14211f
C3593 XA.XIR[0].XIC[9].icell.Ien VPWR 0.18925f
C3594 XA.XIR[12].XIC_dummy_left.icell.PUM VPWR 0.01604f
C3595 XThC.Tn[5] XA.XIR[8].XIC[5].icell.PDM 0.02601f
C3596 XA.XIR[3].XIC[0].icell.Ien XA.XIR[4].XIC[0].icell.PDM 0.02104f
C3597 XThR.Tn[0] XA.XIR[1].XIC[8].icell.PDM 0.04035f
C3598 XThR.Tn[14] XA.XIR[15].XIC[12].icell.PDM 0.04035f
C3599 XA.XIR[12].XIC[0].icell.Ien Vbias 0.19149f
C3600 XThR.XTBN.Y a_n997_1803# 0.22873f
C3601 XThR.Tn[1] XA.XIR[2].XIC[7].icell.PDM 0.04035f
C3602 XA.XIR[7].XIC[12].icell.Ien VPWR 0.18829f
C3603 XThR.Tn[11] Vbias 1.39532f
C3604 XA.XIR[6].XIC[9].icell.Ien XA.XIR[7].XIC[9].icell.PDM 0.02104f
C3605 XThR.XTB6.A data[4] 0.48493f
C3606 XThR.Tn[13] XA.XIR[13].XIC[2].icell.Ien 0.14211f
C3607 XA.XIR[9].XIC[3].icell.PDM XA.XIR[9].XIC[3].icell.Ien 0.04854f
C3608 XA.XIR[7].XIC[9].icell.PDM Vbias 0.03928f
C3609 XThC.Tn[3] XA.XIR[5].XIC[3].icell.Ien 0.04604f
C3610 XThR.Tn[7] XA.XIR[8].XIC[12].icell.PDM 0.04035f
C3611 XThC.Tn[14] XA.XIR[14].XIC[14].icell.Ien 0.04604f
C3612 XThR.XTB6.A XThR.XTB2.Y 0.18237f
C3613 XA.XIR[15].XIC[7].icell.PDM Vbias 0.03928f
C3614 XA.XIR[4].XIC[2].icell.PDM XA.XIR[4].XIC[2].icell.Ien 0.04854f
C3615 XA.XIR[10].XIC[11].icell.Ien VPWR 0.18829f
C3616 XA.XIR[3].XIC[1].icell.Ien VPWR 0.18829f
C3617 XThC.Tn[7] XThR.Tn[2] 0.40741f
C3618 XThC.XTB7.B a_6243_9615# 0.01743f
C3619 XThC.Tn[7] XA.XIR[11].XIC[7].icell.PDM 0.02601f
C3620 XA.XIR[14].XIC[4].icell.Ien XA.XIR[15].XIC[4].icell.PDM 0.02104f
C3621 XA.XIR[11].XIC_dummy_right.icell.Ien XA.XIR[11].XIC_dummy_right.icell.Iout 0.06446f
C3622 XThC.Tn[2] XA.XIR[15].XIC[2].icell.PDM 0.02601f
C3623 XThR.Tn[11] XA.XIR[11].XIC[8].icell.Ien 0.14211f
C3624 XA.XIR[9].XIC[5].icell.PDM Vbias 0.03928f
C3625 XThR.Tn[3] XA.XIR[4].XIC[13].icell.PDM 0.0404f
C3626 XThC.Tn[3] XA.XIR[0].XIC[3].icell.PDM 0.02804f
C3627 XA.XIR[7].XIC[10].icell.PDM VPWR 0.01171f
C3628 XA.XIR[13].XIC[7].icell.Ien XA.XIR[14].XIC[7].icell.PDM 0.02104f
C3629 XA.XIR[9].XIC_dummy_left.icell.Iout VPWR 0.10954f
C3630 XThR.XTBN.Y XThR.Tn[13] 0.56841f
C3631 XThC.Tn[11] XA.XIR[5].XIC[11].icell.PDM 0.02601f
C3632 XA.XIR[3].XIC[10].icell.Ien Iout 0.06801f
C3633 XA.XIR[7].XIC[0].icell.Ien XA.XIR[8].XIC[0].icell.PDM 0.02104f
C3634 XThR.Tn[0] XA.XIR[0].XIC[13].icell.Ien 0.14211f
C3635 XA.XIR[12].XIC[13].icell.Ien XA.XIR[13].XIC[13].icell.PDM 0.02104f
C3636 XA.XIR[15].XIC[8].icell.PDM VPWR 0.01512f
C3637 XA.XIR[13].XIC[8].icell.PDM XA.XIR[13].XIC[8].icell.Ien 0.04854f
C3638 XA.XIR[14].XIC_dummy_left.icell.Ien XA.XIR[15].XIC_dummy_left.icell.PDM 0.02104f
C3639 XThR.Tn[6] XA.XIR[6].XIC[7].icell.Ien 0.14211f
C3640 XA.XIR[8].XIC[7].icell.Ien XA.XIR[9].XIC[7].icell.PDM 0.02104f
C3641 XThR.Tn[12] XA.XIR[12].XIC[10].icell.Ien 0.14211f
C3642 XA.XIR[2].XIC[3].icell.Ien Iout 0.06801f
C3643 XA.XIR[12].XIC[9].icell.Ien XA.XIR[13].XIC[9].icell.PDM 0.02104f
C3644 XA.XIR[0].XIC_dummy_left.icell.Iout XA.XIR[1].XIC_dummy_left.icell.Iout 0.03665f
C3645 XThC.Tn[3] XThR.Tn[6] 0.40738f
C3646 XThC.Tn[1] XA.XIR[13].XIC[1].icell.PDM 0.02601f
C3647 XA.XIR[1].XIC[10].icell.PDM Vbias 0.03928f
C3648 XA.XIR[3].XIC[6].icell.Ien XA.XIR[4].XIC[6].icell.PDM 0.02104f
C3649 XA.XIR[1].XIC[5].icell.Ien Iout 0.06801f
C3650 XThR.Tn[7] XA.XIR[7].XIC[14].icell.Ien 0.144f
C3651 XA.XIR[6].XIC[13].icell.Ien Vbias 0.19161f
C3652 XA.XIR[9].XIC[6].icell.PDM VPWR 0.01171f
C3653 XA.XIR[10].XIC[14].icell.Ien Vbias 0.19161f
C3654 XA.XIR[3].XIC[8].icell.PDM XA.XIR[3].XIC[8].icell.Ien 0.04854f
C3655 XA.XIR[13].XIC[13].icell.Ien VPWR 0.18829f
C3656 XA.XIR[4].XIC[10].icell.PDM Vbias 0.03928f
C3657 XThC.Tn[11] XA.XIR[15].XIC[11].icell.PDM 0.02601f
C3658 XThC.Tn[5] XThR.Tn[11] 0.40738f
C3659 XA.XIR[12].XIC[12].icell.PDM VPWR 0.01171f
C3660 XA.XIR[8].XIC[13].icell.Ien Iout 0.06801f
C3661 XA.XIR[6].XIC[0].icell.PDM XA.XIR[6].XIC[0].icell.Ien 0.04854f
C3662 XA.XIR[14].XIC[7].icell.Ien Vbias 0.19161f
C3663 XThC.XTB7.A XThC.XTB7.Y 0.37429f
C3664 XThC.Tn[8] XA.XIR[0].XIC[8].icell.Ien 0.04654f
C3665 XThC.Tn[1] Iout 0.22482f
C3666 XA.XIR[13].XIC[9].icell.Ien Vbias 0.19161f
C3667 XA.XIR[15].XIC[13].icell.PDM VPWR 0.01512f
C3668 XThC.Tn[7] XA.XIR[10].XIC[7].icell.Ien 0.04604f
C3669 XThR.Tn[4] XA.XIR[5].XIC[5].icell.PDM 0.04035f
C3670 XA.XIR[3].XIC[9].icell.Ien VPWR 0.18829f
C3671 XThC.Tn[11] Vbias 0.82596f
C3672 XA.XIR[1].XIC[11].icell.PDM VPWR 0.01171f
C3673 XThC.Tn[2] XA.XIR[1].XIC[2].icell.Ien 0.04606f
C3674 XThC.Tn[9] XThR.Tn[13] 0.40738f
C3675 XA.XIR[0].XIC_15.icell.Ien Iout 0.06774f
C3676 XA.XIR[2].XIC[2].icell.Ien VPWR 0.18829f
C3677 XA.XIR[4].XIC[11].icell.PDM VPWR 0.01171f
C3678 XA.XIR[6].XIC[2].icell.Ien XA.XIR[7].XIC[2].icell.PDM 0.02104f
C3679 XA.XIR[2].XIC_dummy_right.icell.Iout XA.XIR[3].XIC_dummy_right.icell.Iout 0.04047f
C3680 XThR.Tn[13] XA.XIR[14].XIC[7].icell.PDM 0.04035f
C3681 XThC.Tn[5] XA.XIR[9].XIC[5].icell.PDM 0.02601f
C3682 XA.XIR[1].XIC[4].icell.Ien VPWR 0.18829f
C3683 XThC.Tn[10] XA.XIR[4].XIC[10].icell.Ien 0.04604f
C3684 XThC.Tn[12] XThR.Tn[9] 0.40738f
C3685 XA.XIR[6].XIC[0].icell.Ien Iout 0.06795f
C3686 XThC.Tn[8] XThR.Tn[8] 0.40738f
C3687 XThR.Tn[8] XA.XIR[9].XIC[10].icell.PDM 0.04035f
C3688 XA.XIR[8].XIC[12].icell.Ien VPWR 0.18829f
C3689 bias[1] bias[0] 0.6046f
C3690 XA.XIR[15].XIC_dummy_left.icell.Iout Iout 0.03553f
C3691 bias[2] Vbias 0.4026f
C3692 XThR.Tn[14] XA.XIR[15].XIC[11].icell.PDM 0.04035f
C3693 XThC.Tn[6] XA.XIR[7].XIC[6].icell.Ien 0.04604f
C3694 XA.XIR[1].XIC[13].icell.PDM XA.XIR[1].XIC[13].icell.Ien 0.04854f
C3695 XA.XIR[4].XIC[9].icell.Ien XA.XIR[5].XIC[9].icell.PDM 0.02104f
C3696 XThC.Tn[3] XThR.Tn[4] 0.40738f
C3697 XThR.XTB7.B a_n997_3979# 0.01152f
C3698 XThC.XTBN.Y XThC.Tn[6] 0.49549f
C3699 XA.XIR[5].XIC[1].icell.Ien Vbias 0.19161f
C3700 XA.XIR[7].XIC[1].icell.PDM XA.XIR[7].XIC[1].icell.Ien 0.04854f
C3701 XThR.Tn[5] XA.XIR[6].XIC[7].icell.PDM 0.04035f
C3702 XA.XIR[0].XIC_dummy_right.icell.Iout Iout 0.01732f
C3703 XThR.Tn[14] Vbias 1.39537f
C3704 XA.XIR[11].XIC[0].icell.PDM Vbias 0.03915f
C3705 XA.XIR[14].XIC[12].icell.PDM XA.XIR[14].XIC[12].icell.Ien 0.04854f
C3706 XA.XIR[0].XIC[14].icell.Ien VPWR 0.18783f
C3707 XA.XIR[2].XIC_15.icell.PDM XA.XIR[2].XIC_15.icell.Ien 0.04854f
C3708 XA.XIR[6].XIC[5].icell.Ien Iout 0.06801f
C3709 XThC.Tn[7] XThR.Tn[10] 0.40738f
C3710 XA.XIR[10].XIC[4].icell.PDM Vbias 0.03928f
C3711 XThR.Tn[14] XA.XIR[14].XIC[3].icell.Ien 0.14211f
C3712 XThR.Tn[1] XA.XIR[1].XIC[3].icell.Ien 0.14211f
C3713 XA.XIR[10].XIC[12].icell.Ien Vbias 0.19161f
C3714 XA.XIR[12].XIC[2].icell.Ien XA.XIR[13].XIC[2].icell.PDM 0.02104f
C3715 XA.XIR[13].XIC[11].icell.Ien VPWR 0.18829f
C3716 XThR.Tn[6] XA.XIR[7].XIC[6].icell.PDM 0.04035f
C3717 a_7651_9569# XThC.Tn[8] 0.1927f
C3718 XThC.Tn[7] XA.XIR[14].XIC[7].icell.PDM 0.02601f
C3719 XThR.Tn[13] XA.XIR[13].XIC[7].icell.Ien 0.14211f
C3720 XA.XIR[5].XIC[6].icell.Ien Vbias 0.19161f
C3721 XThR.Tn[12] XA.XIR[12].XIC_15.icell.Ien 0.13564f
C3722 XA.XIR[11].XIC[6].icell.PDM XA.XIR[11].XIC[6].icell.Ien 0.04854f
C3723 XA.XIR[11].XIC[1].icell.PDM VPWR 0.01171f
C3724 XThC.Tn[2] XA.XIR[6].XIC[2].icell.Ien 0.04604f
C3725 XThC.Tn[6] XA.XIR[5].XIC[6].icell.PDM 0.02601f
C3726 XThR.XTB2.Y XThR.Tn[1] 0.17876f
C3727 XA.XIR[10].XIC[5].icell.PDM VPWR 0.01171f
C3728 XThC.Tn[8] XA.XIR[3].XIC[8].icell.Ien 0.04604f
C3729 XA.XIR[11].XIC[4].icell.Ien Iout 0.06801f
C3730 XThC.Tn[8] XA.XIR[1].XIC[8].icell.PDM 0.02602f
C3731 XA.XIR[6].XIC[4].icell.Ien VPWR 0.18829f
C3732 XThR.XTB7.B XThR.Tn[7] 0.07415f
C3733 XThC.Tn[3] XA.XIR[12].XIC[3].icell.Ien 0.04604f
C3734 XA.XIR[10].XIC[6].icell.Ien Iout 0.06801f
C3735 XThR.XTB7.B a_n997_2891# 0.0168f
C3736 XThC.Tn[8] XA.XIR[4].XIC[8].icell.PDM 0.02601f
C3737 XA.XIR[0].XIC[12].icell.PDM Vbias 0.03945f
C3738 XThC.Tn[1] XA.XIR[9].XIC[1].icell.Ien 0.04604f
C3739 XA.XIR[12].XIC[11].icell.PDM VPWR 0.01171f
C3740 XThC.XTB7.B a_8963_9569# 0.02071f
C3741 XA.XIR[13].XIC[14].icell.Ien Vbias 0.19161f
C3742 XA.XIR[3].XIC_15.icell.Ien Iout 0.0694f
C3743 XA.XIR[11].XIC[10].icell.PDM XA.XIR[11].XIC[10].icell.Ien 0.04854f
C3744 XThC.Tn[5] XThR.Tn[14] 0.40738f
C3745 XA.XIR[15].XIC[12].icell.PDM VPWR 0.01512f
C3746 XThC.XTB6.A XThC.XTB7.A 0.44014f
C3747 XThR.Tn[6] XA.XIR[6].XIC[12].icell.Ien 0.14211f
C3748 XA.XIR[2].XIC[8].icell.Ien Iout 0.06801f
C3749 XThR.XTB6.A XThR.XTB7.Y 0.01596f
C3750 XThR.XTB3.Y XThR.XTB5.Y 0.04438f
C3751 XA.XIR[1].XIC[10].icell.Ien Iout 0.06801f
C3752 XA.XIR[2].XIC_dummy_left.icell.Ien XA.XIR[3].XIC_dummy_left.icell.PDM 0.02104f
C3753 XThC.Tn[7] XA.XIR[13].XIC[7].icell.Ien 0.04604f
C3754 XA.XIR[1].XIC[6].icell.PDM XA.XIR[1].XIC[6].icell.Ien 0.04854f
C3755 XA.XIR[0].XIC[13].icell.PDM VPWR 0.01132f
C3756 XA.XIR[4].XIC[2].icell.Ien XA.XIR[5].XIC[2].icell.PDM 0.02104f
C3757 XThC.XTB2.Y XThC.Tn[1] 0.18085f
C3758 XA.XIR[11].XIC[3].icell.Ien VPWR 0.18829f
C3759 XA.XIR[10].XIC[5].icell.Ien VPWR 0.18829f
C3760 XA.XIR[12].XIC_dummy_left.icell.Ien XA.XIR[12].XIC_dummy_left.icell.Iout 0.06446f
C3761 XA.XIR[10].XIC[10].icell.Ien Vbias 0.19161f
C3762 XThC.Tn[6] XA.XIR[8].XIC[6].icell.Ien 0.04604f
C3763 XA.XIR[3].XIC_dummy_right.icell.Iout Iout 0.01732f
C3764 XThR.Tn[10] XA.XIR[11].XIC[9].icell.PDM 0.04035f
C3765 XA.XIR[2].XIC[8].icell.PDM XA.XIR[2].XIC[8].icell.Ien 0.04854f
C3766 XThR.Tn[14] XA.XIR[15].XIC[10].icell.PDM 0.04035f
C3767 XA.XIR[3].XIC[14].icell.Ien VPWR 0.18835f
C3768 XThC.Tn[9] XA.XIR[11].XIC[9].icell.PDM 0.02601f
C3769 XThR.XTBN.Y a_n997_3979# 0.23021f
C3770 XA.XIR[8].XIC[0].icell.PDM XA.XIR[8].XIC[0].icell.Ien 0.04854f
C3771 XA.XIR[2].XIC[7].icell.Ien VPWR 0.18829f
C3772 XThR.Tn[9] XA.XIR[10].XIC[14].icell.PDM 0.04056f
C3773 XA.XIR[9].XIC_dummy_right.icell.Ien XA.XIR[10].XIC_dummy_right.icell.PDM 0.02104f
C3774 XA.XIR[1].XIC[9].icell.Ien VPWR 0.18829f
C3775 XThC.Tn[13] XA.XIR[6].XIC[13].icell.PDM 0.02601f
C3776 XThR.Tn[8] XA.XIR[8].XIC[4].icell.Ien 0.14211f
C3777 XA.XIR[14].XIC_dummy_left.icell.Iout XA.XIR[15].XIC_dummy_left.icell.Iout 0.03665f
C3778 XThC.Tn[10] XA.XIR[3].XIC[10].icell.PDM 0.02601f
C3779 XThC.Tn[0] Vbias 0.27091f
C3780 XA.XIR[6].XIC[3].icell.PDM Vbias 0.03928f
C3781 XA.XIR[2].XIC_dummy_left.icell.Iout XA.XIR[3].XIC_dummy_left.icell.Iout 0.03665f
C3782 XThC.Tn[9] XA.XIR[5].XIC[9].icell.Ien 0.04604f
C3783 XA.XIR[1].XIC_dummy_right.icell.Iout XA.XIR[2].XIC_dummy_right.icell.Iout 0.04047f
C3784 XThC.XTB3.Y a_4067_9615# 0.23056f
C3785 XThR.XTB1.Y XThR.XTB3.Y 0.04033f
C3786 XA.XIR[5].XIC[10].icell.PDM Vbias 0.03928f
C3787 XA.XIR[14].XIC[0].icell.PDM Vbias 0.03915f
C3788 XA.XIR[5].XIC[11].icell.PDM XA.XIR[5].XIC[11].icell.Ien 0.04854f
C3789 a_4067_9615# XThC.Tn[2] 0.27296f
C3790 XThC.Tn[7] XThR.Tn[13] 0.40738f
C3791 XA.XIR[13].XIC[4].icell.PDM Vbias 0.03928f
C3792 XA.XIR[13].XIC[12].icell.Ien Vbias 0.19161f
C3793 XThC.Tn[14] XA.XIR[11].XIC[14].icell.PDM 0.02601f
C3794 XThR.Tn[5] XA.XIR[5].XIC[3].icell.Ien 0.14211f
C3795 XThR.Tn[3] XA.XIR[4].XIC[0].icell.PDM 0.0404f
C3796 XThC.Tn[13] XA.XIR[12].XIC[13].icell.Ien 0.04604f
C3797 XA.XIR[12].XIC[9].icell.PDM Vbias 0.03928f
C3798 XThC.Tn[1] XThR.Tn[9] 0.40738f
C3799 XThC.XTB5.A XThC.XTB6.A 1.80461f
C3800 XA.XIR[9].XIC[2].icell.Ien Vbias 0.19161f
C3801 XA.XIR[14].XIC_dummy_right.icell.Ien XA.XIR[14].XIC_dummy_right.icell.Iout 0.06446f
C3802 XThC.Tn[6] XThR.Tn[8] 0.40738f
C3803 XA.XIR[6].XIC[4].icell.PDM VPWR 0.01171f
C3804 XThR.Tn[2] XA.XIR[3].XIC[14].icell.PDM 0.04056f
C3805 XThR.XTB7.A a_n1049_6699# 0.02294f
C3806 XA.XIR[6].XIC[10].icell.Ien Iout 0.06801f
C3807 XThR.Tn[1] XA.XIR[1].XIC[8].icell.Ien 0.14211f
C3808 XThR.Tn[14] XA.XIR[14].XIC[8].icell.Ien 0.14211f
C3809 XA.XIR[14].XIC[1].icell.PDM VPWR 0.01171f
C3810 XA.XIR[5].XIC[11].icell.PDM VPWR 0.01171f
C3811 XThR.XTB5.Y VPWR 1.0269f
C3812 XThR.XTBN.Y XThR.Tn[7] 0.89994f
C3813 XThR.XTBN.Y a_n997_2891# 0.22804f
C3814 XA.XIR[12].XIC[7].icell.PDM XA.XIR[12].XIC[7].icell.Ien 0.04854f
C3815 XThC.Tn[3] XA.XIR[1].XIC[3].icell.PDM 0.02602f
C3816 XA.XIR[13].XIC[5].icell.PDM VPWR 0.01171f
C3817 XA.XIR[14].XIC[4].icell.Ien Iout 0.06801f
C3818 XA.XIR[12].XIC[10].icell.PDM VPWR 0.01171f
C3819 XA.XIR[5].XIC[11].icell.Ien Vbias 0.19161f
C3820 XThC.Tn[3] XA.XIR[4].XIC[3].icell.PDM 0.02601f
C3821 XA.XIR[13].XIC[6].icell.Ien Iout 0.06801f
C3822 XThC.XTB3.Y XThC.Tn[3] 0.01335f
C3823 XA.XIR[3].XIC[5].icell.PDM Vbias 0.03928f
C3824 XA.XIR[8].XIC[7].icell.PDM Vbias 0.03928f
C3825 XA.XIR[15].XIC[11].icell.PDM VPWR 0.01512f
C3826 XThR.Tn[5] XThR.Tn[6] 0.11432f
C3827 XA.XIR[2].XIC[11].icell.PDM Vbias 0.03928f
C3828 XThC.Tn[2] XThC.Tn[3] 0.59596f
C3829 XA.XIR[11].XIC[9].icell.Ien Iout 0.06801f
C3830 XThR.XTB4.Y XThR.Tn[7] 0.01797f
C3831 XThR.Tn[9] XA.XIR[10].XIC[8].icell.PDM 0.04035f
C3832 XThC.Tn[2] XA.XIR[8].XIC[2].icell.PDM 0.02601f
C3833 XA.XIR[6].XIC[9].icell.Ien VPWR 0.18829f
C3834 XA.XIR[12].XIC[6].icell.Ien Vbias 0.19161f
C3835 XA.XIR[10].XIC_15.icell.Ien Vbias 0.19195f
C3836 VPWR Vbias 98.8642f
C3837 XThC.Tn[8] XA.XIR[1].XIC[8].icell.Ien 0.04606f
C3838 XThR.Tn[10] a_n997_2891# 0.1927f
C3839 XThR.XTBN.A data[5] 0.0148f
C3840 XThC.XTB6.A data[0] 0.48493f
C3841 XA.XIR[8].XIC[8].icell.PDM VPWR 0.01171f
C3842 XA.XIR[3].XIC[6].icell.PDM VPWR 0.01171f
C3843 XA.XIR[14].XIC[3].icell.Ien VPWR 0.18883f
C3844 XThC.Tn[9] XThR.Tn[7] 0.40738f
C3845 XA.XIR[2].XIC[12].icell.PDM VPWR 0.01171f
C3846 XA.XIR[8].XIC[0].icell.Ien XA.XIR[9].XIC[0].icell.PDM 0.02104f
C3847 XA.XIR[2].XIC[13].icell.Ien Iout 0.06801f
C3848 XA.XIR[13].XIC[5].icell.Ien VPWR 0.18829f
C3849 XThR.Tn[12] XA.XIR[13].XIC[2].icell.PDM 0.04035f
C3850 XThR.XTB1.Y VPWR 1.13458f
C3851 XA.XIR[13].XIC[10].icell.Ien Vbias 0.19161f
C3852 XThC.XTB2.Y a_3523_10575# 0.01006f
C3853 XThC.XTB7.Y XThC.Tn[11] 0.07422f
C3854 XThR.XTB6.Y a_n1319_5611# 0.01283f
C3855 XA.XIR[1].XIC_15.icell.Ien Iout 0.0694f
C3856 XA.XIR[5].XIC[4].icell.PDM XA.XIR[5].XIC[4].icell.Ien 0.04854f
C3857 XA.XIR[12].XIC[11].icell.Ien XA.XIR[13].XIC[11].icell.PDM 0.02104f
C3858 XA.XIR[10].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3859 XThR.Tn[9] XA.XIR[10].XIC[13].icell.PDM 0.0404f
C3860 XThC.Tn[4] XA.XIR[11].XIC[4].icell.PDM 0.02601f
C3861 XA.XIR[11].XIC[8].icell.Ien VPWR 0.18829f
C3862 XThC.Tn[9] XA.XIR[14].XIC[9].icell.PDM 0.02601f
C3863 XThR.XTB7.Y XThR.Tn[12] 0.07066f
C3864 XThC.Tn[12] XA.XIR[7].XIC[12].icell.Ien 0.04604f
C3865 XThC.Tn[0] XA.XIR[0].XIC[0].icell.PDM 0.02804f
C3866 XA.XIR[0].XIC[14].icell.PDM XA.XIR[0].XIC[14].icell.Ien 0.04854f
C3867 XThC.Tn[5] XA.XIR[3].XIC[5].icell.PDM 0.02601f
C3868 XThC.Tn[8] XA.XIR[5].XIC[8].icell.PDM 0.02601f
C3869 XThR.Tn[0] XA.XIR[1].XIC[10].icell.PDM 0.04035f
C3870 XA.XIR[5].XIC[3].icell.Ien Iout 0.06801f
C3871 XThR.Tn[4] XThR.Tn[5] 0.12171f
C3872 XThR.Tn[1] XA.XIR[2].XIC[9].icell.PDM 0.04035f
C3873 XThC.Tn[8] XThR.Tn[3] 0.40738f
C3874 XA.XIR[2].XIC[12].icell.Ien VPWR 0.18829f
C3875 XA.XIR[1].XIC_dummy_right.icell.Iout Iout 0.01732f
C3876 XThC.Tn[3] XA.XIR[15].XIC[3].icell.Ien 0.04292f
C3877 XThR.Tn[7] XA.XIR[8].XIC[14].icell.PDM 0.04056f
C3878 XA.XIR[1].XIC[14].icell.Ien VPWR 0.18835f
C3879 XA.XIR[7].XIC[11].icell.PDM Vbias 0.03928f
C3880 XThC.Tn[5] VPWR 3.59867f
C3881 XThR.Tn[8] XA.XIR[8].XIC[9].icell.Ien 0.14211f
C3882 XThC.Tn[14] XA.XIR[14].XIC[14].icell.PDM 0.02601f
C3883 XA.XIR[15].XIC[9].icell.PDM Vbias 0.03928f
C3884 XA.XIR[4].XIC[4].icell.Ien Vbias 0.19161f
C3885 XA.XIR[5].XIC[13].icell.Ien XA.XIR[6].XIC[13].icell.PDM 0.02104f
C3886 XA.XIR[3].XIC_dummy_left.icell.Iout VPWR 0.11229f
C3887 XThR.XTB6.Y XThR.Tn[5] 0.20186f
C3888 XThC.Tn[14] XA.XIR[9].XIC[14].icell.Ien 0.04604f
C3889 XThC.Tn[11] XThR.Tn[0] 0.40763f
C3890 XThC.Tn[13] XThR.Tn[5] 0.40739f
C3891 XThC.Tn[4] XA.XIR[11].XIC[4].icell.Ien 0.04604f
C3892 XA.XIR[12].XIC[1].icell.Ien VPWR 0.18829f
C3893 XThC.Tn[8] XA.XIR[6].XIC[8].icell.Ien 0.04604f
C3894 XThR.Tn[5] XA.XIR[5].XIC[8].icell.Ien 0.14211f
C3895 XA.XIR[14].XIC[6].icell.PDM XA.XIR[14].XIC[6].icell.Ien 0.04854f
C3896 XA.XIR[9].XIC[7].icell.PDM Vbias 0.03928f
C3897 XThR.XTBN.Y a_n997_1579# 0.23006f
C3898 XA.XIR[5].XIC[2].icell.Ien VPWR 0.18829f
C3899 XA.XIR[7].XIC[12].icell.PDM VPWR 0.01171f
C3900 XThR.XTB7.Y a_n1049_5317# 0.27822f
C3901 XThC.Tn[9] XA.XIR[12].XIC[9].icell.Ien 0.04604f
C3902 XA.XIR[7].XIC_dummy_left.icell.Ien XA.XIR[7].XIC_dummy_left.icell.Iout 0.06446f
C3903 XThR.Tn[6] Iout 1.12758f
C3904 XA.XIR[11].XIC[14].icell.Ien Iout 0.06801f
C3905 XA.XIR[10].XIC_dummy_left.icell.Ien XA.XIR[11].XIC_dummy_left.icell.PDM 0.02104f
C3906 XA.XIR[9].XIC[7].icell.Ien Vbias 0.19161f
C3907 XA.XIR[15].XIC[10].icell.PDM VPWR 0.01512f
C3908 XThC.Tn[2] XA.XIR[9].XIC[2].icell.PDM 0.02601f
C3909 XA.XIR[6].XIC_15.icell.Ien Iout 0.0694f
C3910 XThC.Tn[12] XA.XIR[12].XIC[12].icell.PDM 0.02601f
C3911 XA.XIR[2].XIC[1].icell.PDM XA.XIR[2].XIC[1].icell.Ien 0.04854f
C3912 XThR.Tn[1] XA.XIR[1].XIC[13].icell.Ien 0.14211f
C3913 XA.XIR[1].XIC[12].icell.PDM Vbias 0.03928f
C3914 XA.XIR[9].XIC[8].icell.PDM VPWR 0.01171f
C3915 XA.XIR[14].XIC[9].icell.Ien Iout 0.06801f
C3916 XThC.Tn[8] data[0] 0.01744f
C3917 XA.XIR[0].XIC[0].icell.PDM VPWR 0.01132f
C3918 XA.XIR[14].XIC[10].icell.PDM XA.XIR[14].XIC[10].icell.Ien 0.04854f
C3919 XA.XIR[7].XIC[3].icell.Ien Vbias 0.19161f
C3920 XA.XIR[4].XIC[12].icell.PDM Vbias 0.03928f
C3921 XThC.XTB7.B Vbias 0.12116f
C3922 XThC.Tn[10] XThR.Tn[2] 0.40741f
C3923 XA.XIR[13].XIC_15.icell.Ien Vbias 0.19195f
C3924 XA.XIR[12].XIC[0].icell.Ien XThR.Tn[12] 0.14211f
C3925 XA.XIR[0].XIC[7].icell.PDM XA.XIR[0].XIC[7].icell.Ien 0.04854f
C3926 XThR.Tn[4] XA.XIR[5].XIC[7].icell.PDM 0.04035f
C3927 XA.XIR[6].XIC_dummy_right.icell.Iout Iout 0.01732f
C3928 XThR.Tn[11] XThR.Tn[12] 0.1626f
C3929 XA.XIR[1].XIC[13].icell.PDM VPWR 0.01171f
C3930 XA.XIR[6].XIC[14].icell.Ien VPWR 0.18835f
C3931 XThC.Tn[12] XA.XIR[8].XIC[12].icell.Ien 0.04604f
C3932 XThR.Tn[9] XA.XIR[10].XIC[12].icell.PDM 0.04035f
C3933 XA.XIR[4].XIC[13].icell.PDM VPWR 0.01171f
C3934 XThC.XTB7.A XThC.Tn[6] 0.10502f
C3935 XThR.Tn[13] XA.XIR[14].XIC[9].icell.PDM 0.04035f
C3936 XThC.Tn[4] XA.XIR[14].XIC[4].icell.PDM 0.02601f
C3937 XA.XIR[13].XIC_dummy_right.icell.PUM VPWR 0.01691f
C3938 XA.XIR[14].XIC[8].icell.Ien VPWR 0.18883f
C3939 XThR.XTB5.A XThR.XTBN.A 0.06303f
C3940 XThC.Tn[13] XA.XIR[15].XIC[13].icell.Ien 0.04292f
C3941 XThR.Tn[8] XA.XIR[9].XIC[12].icell.PDM 0.04035f
C3942 XA.XIR[5].XIC[6].icell.Ien XA.XIR[6].XIC[6].icell.PDM 0.02104f
C3943 XThR.Tn[4] Iout 1.12761f
C3944 XThC.Tn[3] XA.XIR[5].XIC[3].icell.PDM 0.02601f
C3945 XA.XIR[12].XIC_dummy_right.icell.Ien XA.XIR[13].XIC_dummy_right.icell.PDM 0.02104f
C3946 XThC.Tn[6] XA.XIR[2].XIC[6].icell.Ien 0.04605f
C3947 XThC.Tn[8] XThR.Tn[11] 0.40738f
C3948 XA.XIR[11].XIC[12].icell.Ien Iout 0.06801f
C3949 XA.XIR[10].XIC_dummy_left.icell.Ien VPWR 0.39005f
C3950 XA.XIR[15].XIC[1].icell.Ien Vbias 0.15966f
C3951 data[7] VGND 0.49949f
C3952 data[6] VGND 0.47974f
C3953 data[4] VGND 0.59317f
C3954 data[5] VGND 1.17814f
C3955 Iout VGND 0.32108p
C3956 data[3] VGND 0.49926f
C3957 data[2] VGND 0.48064f
C3958 data[0] VGND 0.59269f
C3959 data[1] VGND 1.17844f
C3960 Vbias VGND 0.17164p
C3961 bias[0] VGND 1.39569f
C3962 bias[1] VGND 0.46888f
C3963 bias[2] VGND 0.40015f
C3964 VPWR VGND 0.37401p
C3965 a_n997_715# VGND 0.5638f
C3966 XA.XIR[15].XIC_dummy_right.icell.Iout VGND 0.7524f
C3967 XA.XIR[15].XIC_dummy_right.icell.SM VGND 0.01013f
C3968 XA.XIR[15].XIC_dummy_right.icell.Ien VGND 0.64532f
C3969 XA.XIR[15].XIC_15.icell.Ien VGND 0.44493f
C3970 XA.XIR[15].XIC[14].icell.Ien VGND 0.4451f
C3971 XA.XIR[15].XIC[13].icell.Ien VGND 0.44506f
C3972 XA.XIR[15].XIC[12].icell.Ien VGND 0.44506f
C3973 XA.XIR[15].XIC[11].icell.Ien VGND 0.44506f
C3974 XA.XIR[15].XIC[10].icell.Ien VGND 0.44506f
C3975 XA.XIR[15].XIC[9].icell.Ien VGND 0.44506f
C3976 XA.XIR[15].XIC[8].icell.Ien VGND 0.44506f
C3977 XA.XIR[15].XIC[7].icell.Ien VGND 0.44506f
C3978 XA.XIR[15].XIC[6].icell.Ien VGND 0.44506f
C3979 XA.XIR[15].XIC[5].icell.Ien VGND 0.44506f
C3980 XA.XIR[15].XIC[4].icell.Ien VGND 0.44506f
C3981 XA.XIR[15].XIC[3].icell.Ien VGND 0.44506f
C3982 XA.XIR[15].XIC[2].icell.Ien VGND 0.44506f
C3983 XA.XIR[15].XIC_dummy_left.icell.Iout VGND 0.70682f
C3984 XA.XIR[15].XIC[1].icell.Ien VGND 0.44506f
C3985 XA.XIR[15].XIC[0].icell.Ien VGND 0.44521f
C3986 XA.XIR[15].XIC_dummy_left.icell.SM VGND 0.01033f
C3987 XA.XIR[15].XIC_dummy_left.icell.Ien VGND 0.6116f
C3988 XA.XIR[15].XIC_dummy_right.icell.PDM VGND 0.23278f
C3989 XA.XIR[15].XIC_15.icell.PDM VGND 0.18786f
C3990 XA.XIR[15].XIC[14].icell.PDM VGND 0.18744f
C3991 XA.XIR[15].XIC[13].icell.PDM VGND 0.18744f
C3992 XA.XIR[15].XIC[12].icell.PDM VGND 0.18744f
C3993 XA.XIR[15].XIC[11].icell.PDM VGND 0.18744f
C3994 XA.XIR[15].XIC[10].icell.PDM VGND 0.18744f
C3995 XA.XIR[15].XIC[9].icell.PDM VGND 0.18744f
C3996 XA.XIR[15].XIC[8].icell.PDM VGND 0.18744f
C3997 XA.XIR[15].XIC[7].icell.PDM VGND 0.18744f
C3998 XA.XIR[15].XIC[6].icell.PDM VGND 0.18744f
C3999 XA.XIR[15].XIC[5].icell.PDM VGND 0.18744f
C4000 XA.XIR[15].XIC[4].icell.PDM VGND 0.18744f
C4001 XA.XIR[15].XIC[3].icell.PDM VGND 0.18744f
C4002 XA.XIR[15].XIC[2].icell.PDM VGND 0.18744f
C4003 XA.XIR[15].XIC[1].icell.PDM VGND 0.18744f
C4004 XA.XIR[15].XIC[0].icell.PDM VGND 0.1876f
C4005 XA.XIR[15].XIC_dummy_left.icell.PDM VGND 0.22703f
C4006 XA.XIR[14].XIC_dummy_right.icell.Iout VGND 0.85788f
C4007 XA.XIR[14].XIC_dummy_right.icell.SM VGND 0.01013f
C4008 XA.XIR[14].XIC_dummy_right.icell.Ien VGND 0.60818f
C4009 XA.XIR[14].XIC_15.icell.Ien VGND 0.37264f
C4010 XA.XIR[14].XIC[14].icell.Ien VGND 0.37333f
C4011 XA.XIR[14].XIC[13].icell.Ien VGND 0.3733f
C4012 XA.XIR[14].XIC[12].icell.Ien VGND 0.3733f
C4013 XA.XIR[14].XIC[11].icell.Ien VGND 0.3733f
C4014 XA.XIR[14].XIC[10].icell.Ien VGND 0.3733f
C4015 XA.XIR[14].XIC[9].icell.Ien VGND 0.3733f
C4016 XA.XIR[14].XIC[8].icell.Ien VGND 0.3733f
C4017 XA.XIR[14].XIC[7].icell.Ien VGND 0.3733f
C4018 XA.XIR[14].XIC[6].icell.Ien VGND 0.3733f
C4019 XA.XIR[14].XIC[5].icell.Ien VGND 0.3733f
C4020 XA.XIR[14].XIC[4].icell.Ien VGND 0.3733f
C4021 XA.XIR[14].XIC[3].icell.Ien VGND 0.3733f
C4022 XA.XIR[14].XIC[2].icell.Ien VGND 0.3733f
C4023 XA.XIR[14].XIC_dummy_left.icell.Iout VGND 0.8066f
C4024 XThR.Tn[14] VGND 13.06755f
C4025 XA.XIR[14].XIC[1].icell.Ien VGND 0.3733f
C4026 a_n997_1579# VGND 0.54776f
C4027 XA.XIR[14].XIC[0].icell.Ien VGND 0.37345f
C4028 XA.XIR[14].XIC_dummy_left.icell.SM VGND 0.01033f
C4029 XA.XIR[14].XIC_dummy_left.icell.Ien VGND 0.57576f
C4030 a_n997_1803# VGND 0.53619f
C4031 XA.XIR[14].XIC_dummy_right.icell.PDM VGND 0.23384f
C4032 XA.XIR[14].XIC_15.icell.PDM VGND 0.18862f
C4033 XA.XIR[14].XIC[14].icell.PDM VGND 0.1882f
C4034 XA.XIR[14].XIC[13].icell.PDM VGND 0.1882f
C4035 XA.XIR[14].XIC[12].icell.PDM VGND 0.1882f
C4036 XA.XIR[14].XIC[11].icell.PDM VGND 0.1882f
C4037 XA.XIR[14].XIC[10].icell.PDM VGND 0.1882f
C4038 XA.XIR[14].XIC[9].icell.PDM VGND 0.1882f
C4039 XA.XIR[14].XIC[8].icell.PDM VGND 0.1882f
C4040 XA.XIR[14].XIC[7].icell.PDM VGND 0.1882f
C4041 XA.XIR[14].XIC[6].icell.PDM VGND 0.1882f
C4042 XA.XIR[14].XIC[5].icell.PDM VGND 0.1882f
C4043 XA.XIR[14].XIC[4].icell.PDM VGND 0.1882f
C4044 XA.XIR[14].XIC[3].icell.PDM VGND 0.1882f
C4045 XA.XIR[14].XIC[2].icell.PDM VGND 0.1882f
C4046 XA.XIR[14].XIC[1].icell.PDM VGND 0.1882f
C4047 XA.XIR[14].XIC[0].icell.PDM VGND 0.18836f
C4048 XA.XIR[14].XIC_dummy_left.icell.PDM VGND 0.22809f
C4049 XA.XIR[13].XIC_dummy_right.icell.Iout VGND 0.85788f
C4050 XA.XIR[13].XIC_dummy_right.icell.SM VGND 0.01013f
C4051 XA.XIR[13].XIC_dummy_right.icell.Ien VGND 0.60818f
C4052 XA.XIR[13].XIC_15.icell.Ien VGND 0.37264f
C4053 XA.XIR[13].XIC[14].icell.Ien VGND 0.37333f
C4054 XA.XIR[13].XIC[13].icell.Ien VGND 0.3733f
C4055 XA.XIR[13].XIC[12].icell.Ien VGND 0.3733f
C4056 XA.XIR[13].XIC[11].icell.Ien VGND 0.3733f
C4057 XA.XIR[13].XIC[10].icell.Ien VGND 0.3733f
C4058 XA.XIR[13].XIC[9].icell.Ien VGND 0.3733f
C4059 XA.XIR[13].XIC[8].icell.Ien VGND 0.3733f
C4060 XA.XIR[13].XIC[7].icell.Ien VGND 0.3733f
C4061 XA.XIR[13].XIC[6].icell.Ien VGND 0.3733f
C4062 XA.XIR[13].XIC[5].icell.Ien VGND 0.3733f
C4063 XA.XIR[13].XIC[4].icell.Ien VGND 0.3733f
C4064 XA.XIR[13].XIC[3].icell.Ien VGND 0.3733f
C4065 XA.XIR[13].XIC[2].icell.Ien VGND 0.3733f
C4066 XA.XIR[13].XIC_dummy_left.icell.Iout VGND 0.80664f
C4067 XThR.Tn[13] VGND 12.91167f
C4068 XA.XIR[13].XIC[1].icell.Ien VGND 0.3733f
C4069 XA.XIR[13].XIC[0].icell.Ien VGND 0.37345f
C4070 XA.XIR[13].XIC_dummy_left.icell.SM VGND 0.01033f
C4071 XA.XIR[13].XIC_dummy_left.icell.Ien VGND 0.57422f
C4072 XA.XIR[13].XIC_dummy_right.icell.PDM VGND 0.23384f
C4073 XA.XIR[13].XIC_15.icell.PDM VGND 0.18862f
C4074 XA.XIR[13].XIC[14].icell.PDM VGND 0.1882f
C4075 XA.XIR[13].XIC[13].icell.PDM VGND 0.1882f
C4076 XA.XIR[13].XIC[12].icell.PDM VGND 0.1882f
C4077 XA.XIR[13].XIC[11].icell.PDM VGND 0.1882f
C4078 XA.XIR[13].XIC[10].icell.PDM VGND 0.1882f
C4079 XA.XIR[13].XIC[9].icell.PDM VGND 0.1882f
C4080 XA.XIR[13].XIC[8].icell.PDM VGND 0.1882f
C4081 XA.XIR[13].XIC[7].icell.PDM VGND 0.1882f
C4082 XA.XIR[13].XIC[6].icell.PDM VGND 0.1882f
C4083 XA.XIR[13].XIC[5].icell.PDM VGND 0.1882f
C4084 XA.XIR[13].XIC[4].icell.PDM VGND 0.1882f
C4085 XA.XIR[13].XIC[3].icell.PDM VGND 0.1882f
C4086 XA.XIR[13].XIC[2].icell.PDM VGND 0.1882f
C4087 XA.XIR[13].XIC[1].icell.PDM VGND 0.1882f
C4088 XA.XIR[13].XIC[0].icell.PDM VGND 0.18836f
C4089 XA.XIR[13].XIC_dummy_left.icell.PDM VGND 0.22809f
C4090 XA.XIR[12].XIC_dummy_right.icell.Iout VGND 0.85788f
C4091 XA.XIR[12].XIC_dummy_right.icell.SM VGND 0.01013f
C4092 XA.XIR[12].XIC_dummy_right.icell.Ien VGND 0.60818f
C4093 XA.XIR[12].XIC_15.icell.Ien VGND 0.37264f
C4094 XA.XIR[12].XIC[14].icell.Ien VGND 0.37333f
C4095 XA.XIR[12].XIC[13].icell.Ien VGND 0.3733f
C4096 XA.XIR[12].XIC[12].icell.Ien VGND 0.3733f
C4097 XA.XIR[12].XIC[11].icell.Ien VGND 0.3733f
C4098 XA.XIR[12].XIC[10].icell.Ien VGND 0.3733f
C4099 XA.XIR[12].XIC[9].icell.Ien VGND 0.3733f
C4100 XA.XIR[12].XIC[8].icell.Ien VGND 0.3733f
C4101 XA.XIR[12].XIC[7].icell.Ien VGND 0.3733f
C4102 XA.XIR[12].XIC[6].icell.Ien VGND 0.3733f
C4103 XA.XIR[12].XIC[5].icell.Ien VGND 0.3733f
C4104 XA.XIR[12].XIC[4].icell.Ien VGND 0.3733f
C4105 XA.XIR[12].XIC[3].icell.Ien VGND 0.3733f
C4106 XA.XIR[12].XIC[2].icell.Ien VGND 0.3733f
C4107 XA.XIR[12].XIC_dummy_left.icell.Iout VGND 0.80529f
C4108 XThR.Tn[12] VGND 12.80173f
C4109 XA.XIR[12].XIC[1].icell.Ien VGND 0.3733f
C4110 XA.XIR[12].XIC[0].icell.Ien VGND 0.37345f
C4111 XA.XIR[12].XIC_dummy_left.icell.SM VGND 0.01033f
C4112 XA.XIR[12].XIC_dummy_left.icell.Ien VGND 0.5728f
C4113 a_n997_2667# VGND 0.5457f
C4114 XA.XIR[12].XIC_dummy_right.icell.PDM VGND 0.23384f
C4115 XA.XIR[12].XIC_15.icell.PDM VGND 0.18862f
C4116 XA.XIR[12].XIC[14].icell.PDM VGND 0.1882f
C4117 XA.XIR[12].XIC[13].icell.PDM VGND 0.1882f
C4118 XA.XIR[12].XIC[12].icell.PDM VGND 0.1882f
C4119 XA.XIR[12].XIC[11].icell.PDM VGND 0.1882f
C4120 XA.XIR[12].XIC[10].icell.PDM VGND 0.1882f
C4121 XA.XIR[12].XIC[9].icell.PDM VGND 0.1882f
C4122 XA.XIR[12].XIC[8].icell.PDM VGND 0.1882f
C4123 XA.XIR[12].XIC[7].icell.PDM VGND 0.1882f
C4124 XA.XIR[12].XIC[6].icell.PDM VGND 0.1882f
C4125 XA.XIR[12].XIC[5].icell.PDM VGND 0.1882f
C4126 XA.XIR[12].XIC[4].icell.PDM VGND 0.1882f
C4127 XA.XIR[12].XIC[3].icell.PDM VGND 0.1882f
C4128 XA.XIR[12].XIC[2].icell.PDM VGND 0.1882f
C4129 XA.XIR[12].XIC[1].icell.PDM VGND 0.1882f
C4130 XA.XIR[12].XIC[0].icell.PDM VGND 0.18836f
C4131 XA.XIR[12].XIC_dummy_left.icell.PDM VGND 0.22809f
C4132 XA.XIR[11].XIC_dummy_right.icell.Iout VGND 0.85788f
C4133 XA.XIR[11].XIC_dummy_right.icell.SM VGND 0.01013f
C4134 XA.XIR[11].XIC_dummy_right.icell.Ien VGND 0.60818f
C4135 XA.XIR[11].XIC_15.icell.Ien VGND 0.37264f
C4136 XA.XIR[11].XIC[14].icell.Ien VGND 0.37333f
C4137 XA.XIR[11].XIC[13].icell.Ien VGND 0.3733f
C4138 XA.XIR[11].XIC[12].icell.Ien VGND 0.3733f
C4139 XA.XIR[11].XIC[11].icell.Ien VGND 0.3733f
C4140 XA.XIR[11].XIC[10].icell.Ien VGND 0.3733f
C4141 XA.XIR[11].XIC[9].icell.Ien VGND 0.3733f
C4142 XA.XIR[11].XIC[8].icell.Ien VGND 0.3733f
C4143 XA.XIR[11].XIC[7].icell.Ien VGND 0.3733f
C4144 XA.XIR[11].XIC[6].icell.Ien VGND 0.3733f
C4145 XA.XIR[11].XIC[5].icell.Ien VGND 0.3733f
C4146 XA.XIR[11].XIC[4].icell.Ien VGND 0.3733f
C4147 XA.XIR[11].XIC[3].icell.Ien VGND 0.3733f
C4148 XA.XIR[11].XIC[2].icell.Ien VGND 0.3733f
C4149 XA.XIR[11].XIC_dummy_left.icell.Iout VGND 0.80765f
C4150 XThR.Tn[11] VGND 12.86402f
C4151 XA.XIR[11].XIC[1].icell.Ien VGND 0.3733f
C4152 a_n997_2891# VGND 0.54795f
C4153 XA.XIR[11].XIC[0].icell.Ien VGND 0.37345f
C4154 XA.XIR[11].XIC_dummy_left.icell.SM VGND 0.01033f
C4155 XA.XIR[11].XIC_dummy_left.icell.Ien VGND 0.57294f
C4156 XA.XIR[11].XIC_dummy_right.icell.PDM VGND 0.23384f
C4157 XA.XIR[11].XIC_15.icell.PDM VGND 0.18862f
C4158 XA.XIR[11].XIC[14].icell.PDM VGND 0.1882f
C4159 XA.XIR[11].XIC[13].icell.PDM VGND 0.1882f
C4160 XA.XIR[11].XIC[12].icell.PDM VGND 0.1882f
C4161 XA.XIR[11].XIC[11].icell.PDM VGND 0.1882f
C4162 XA.XIR[11].XIC[10].icell.PDM VGND 0.1882f
C4163 XA.XIR[11].XIC[9].icell.PDM VGND 0.1882f
C4164 XA.XIR[11].XIC[8].icell.PDM VGND 0.1882f
C4165 XA.XIR[11].XIC[7].icell.PDM VGND 0.1882f
C4166 XA.XIR[11].XIC[6].icell.PDM VGND 0.1882f
C4167 XA.XIR[11].XIC[5].icell.PDM VGND 0.1882f
C4168 XA.XIR[11].XIC[4].icell.PDM VGND 0.1882f
C4169 XA.XIR[11].XIC[3].icell.PDM VGND 0.1882f
C4170 XA.XIR[11].XIC[2].icell.PDM VGND 0.1882f
C4171 XA.XIR[11].XIC[1].icell.PDM VGND 0.1882f
C4172 XA.XIR[11].XIC[0].icell.PDM VGND 0.18836f
C4173 XA.XIR[11].XIC_dummy_left.icell.PDM VGND 0.22809f
C4174 XA.XIR[10].XIC_dummy_right.icell.Iout VGND 0.85788f
C4175 XA.XIR[10].XIC_dummy_right.icell.SM VGND 0.01013f
C4176 XA.XIR[10].XIC_dummy_right.icell.Ien VGND 0.60818f
C4177 XA.XIR[10].XIC_15.icell.Ien VGND 0.37264f
C4178 XA.XIR[10].XIC[14].icell.Ien VGND 0.37333f
C4179 XA.XIR[10].XIC[13].icell.Ien VGND 0.3733f
C4180 XA.XIR[10].XIC[12].icell.Ien VGND 0.3733f
C4181 XA.XIR[10].XIC[11].icell.Ien VGND 0.3733f
C4182 XA.XIR[10].XIC[10].icell.Ien VGND 0.3733f
C4183 XA.XIR[10].XIC[9].icell.Ien VGND 0.3733f
C4184 XA.XIR[10].XIC[8].icell.Ien VGND 0.3733f
C4185 XA.XIR[10].XIC[7].icell.Ien VGND 0.3733f
C4186 XA.XIR[10].XIC[6].icell.Ien VGND 0.3733f
C4187 XA.XIR[10].XIC[5].icell.Ien VGND 0.3733f
C4188 XA.XIR[10].XIC[4].icell.Ien VGND 0.3733f
C4189 XA.XIR[10].XIC[3].icell.Ien VGND 0.3733f
C4190 XA.XIR[10].XIC[2].icell.Ien VGND 0.3733f
C4191 XA.XIR[10].XIC_dummy_left.icell.Iout VGND 0.80648f
C4192 XThR.Tn[10] VGND 12.83941f
C4193 XA.XIR[10].XIC[1].icell.Ien VGND 0.3733f
C4194 XA.XIR[10].XIC[0].icell.Ien VGND 0.37345f
C4195 XA.XIR[10].XIC_dummy_left.icell.SM VGND 0.01033f
C4196 XA.XIR[10].XIC_dummy_left.icell.Ien VGND 0.57422f
C4197 XA.XIR[10].XIC_dummy_right.icell.PDM VGND 0.23384f
C4198 XA.XIR[10].XIC_15.icell.PDM VGND 0.18862f
C4199 XA.XIR[10].XIC[14].icell.PDM VGND 0.1882f
C4200 XA.XIR[10].XIC[13].icell.PDM VGND 0.1882f
C4201 XA.XIR[10].XIC[12].icell.PDM VGND 0.1882f
C4202 XA.XIR[10].XIC[11].icell.PDM VGND 0.1882f
C4203 XA.XIR[10].XIC[10].icell.PDM VGND 0.1882f
C4204 XA.XIR[10].XIC[9].icell.PDM VGND 0.1882f
C4205 XA.XIR[10].XIC[8].icell.PDM VGND 0.1882f
C4206 XA.XIR[10].XIC[7].icell.PDM VGND 0.1882f
C4207 XA.XIR[10].XIC[6].icell.PDM VGND 0.1882f
C4208 XA.XIR[10].XIC[5].icell.PDM VGND 0.1882f
C4209 XA.XIR[10].XIC[4].icell.PDM VGND 0.1882f
C4210 XA.XIR[10].XIC[3].icell.PDM VGND 0.1882f
C4211 XA.XIR[10].XIC[2].icell.PDM VGND 0.1882f
C4212 XA.XIR[10].XIC[1].icell.PDM VGND 0.1882f
C4213 XA.XIR[10].XIC[0].icell.PDM VGND 0.18836f
C4214 XA.XIR[10].XIC_dummy_left.icell.PDM VGND 0.22809f
C4215 XA.XIR[9].XIC_dummy_right.icell.Iout VGND 0.85788f
C4216 XA.XIR[9].XIC_dummy_right.icell.SM VGND 0.01013f
C4217 XA.XIR[9].XIC_dummy_right.icell.Ien VGND 0.60818f
C4218 XA.XIR[9].XIC_15.icell.Ien VGND 0.37264f
C4219 XA.XIR[9].XIC[14].icell.Ien VGND 0.37333f
C4220 XA.XIR[9].XIC[13].icell.Ien VGND 0.3733f
C4221 XA.XIR[9].XIC[12].icell.Ien VGND 0.3733f
C4222 XA.XIR[9].XIC[11].icell.Ien VGND 0.3733f
C4223 XA.XIR[9].XIC[10].icell.Ien VGND 0.3733f
C4224 XA.XIR[9].XIC[9].icell.Ien VGND 0.3733f
C4225 XA.XIR[9].XIC[8].icell.Ien VGND 0.3733f
C4226 XA.XIR[9].XIC[7].icell.Ien VGND 0.3733f
C4227 XA.XIR[9].XIC[6].icell.Ien VGND 0.3733f
C4228 XA.XIR[9].XIC[5].icell.Ien VGND 0.3733f
C4229 XA.XIR[9].XIC[4].icell.Ien VGND 0.3733f
C4230 XA.XIR[9].XIC[3].icell.Ien VGND 0.3733f
C4231 XA.XIR[9].XIC[2].icell.Ien VGND 0.3733f
C4232 XA.XIR[9].XIC_dummy_left.icell.Iout VGND 0.80834f
C4233 XA.XIR[9].XIC[1].icell.Ien VGND 0.3733f
C4234 XThR.Tn[9] VGND 12.8472f
C4235 a_n997_3755# VGND 0.54861f
C4236 XA.XIR[9].XIC[0].icell.Ien VGND 0.37345f
C4237 XA.XIR[9].XIC_dummy_left.icell.SM VGND 0.01033f
C4238 XA.XIR[9].XIC_dummy_left.icell.Ien VGND 0.5732f
C4239 a_n997_3979# VGND 0.54721f
C4240 XA.XIR[9].XIC_dummy_right.icell.PDM VGND 0.23384f
C4241 XA.XIR[9].XIC_15.icell.PDM VGND 0.18862f
C4242 XA.XIR[9].XIC[14].icell.PDM VGND 0.1882f
C4243 XA.XIR[9].XIC[13].icell.PDM VGND 0.1882f
C4244 XA.XIR[9].XIC[12].icell.PDM VGND 0.1882f
C4245 XA.XIR[9].XIC[11].icell.PDM VGND 0.1882f
C4246 XA.XIR[9].XIC[10].icell.PDM VGND 0.1882f
C4247 XA.XIR[9].XIC[9].icell.PDM VGND 0.1882f
C4248 XA.XIR[9].XIC[8].icell.PDM VGND 0.1882f
C4249 XA.XIR[9].XIC[7].icell.PDM VGND 0.1882f
C4250 XA.XIR[9].XIC[6].icell.PDM VGND 0.1882f
C4251 XA.XIR[9].XIC[5].icell.PDM VGND 0.1882f
C4252 XA.XIR[9].XIC[4].icell.PDM VGND 0.1882f
C4253 XA.XIR[9].XIC[3].icell.PDM VGND 0.1882f
C4254 XA.XIR[9].XIC[2].icell.PDM VGND 0.1882f
C4255 XA.XIR[9].XIC[1].icell.PDM VGND 0.1882f
C4256 XA.XIR[9].XIC[0].icell.PDM VGND 0.18836f
C4257 XA.XIR[9].XIC_dummy_left.icell.PDM VGND 0.22809f
C4258 XA.XIR[8].XIC_dummy_right.icell.Iout VGND 0.85788f
C4259 XA.XIR[8].XIC_dummy_right.icell.SM VGND 0.01013f
C4260 XA.XIR[8].XIC_dummy_right.icell.Ien VGND 0.60818f
C4261 XA.XIR[8].XIC_15.icell.Ien VGND 0.37264f
C4262 XA.XIR[8].XIC[14].icell.Ien VGND 0.37333f
C4263 XA.XIR[8].XIC[13].icell.Ien VGND 0.3733f
C4264 XA.XIR[8].XIC[12].icell.Ien VGND 0.3733f
C4265 XA.XIR[8].XIC[11].icell.Ien VGND 0.3733f
C4266 XA.XIR[8].XIC[10].icell.Ien VGND 0.3733f
C4267 XA.XIR[8].XIC[9].icell.Ien VGND 0.3733f
C4268 XA.XIR[8].XIC[8].icell.Ien VGND 0.3733f
C4269 XA.XIR[8].XIC[7].icell.Ien VGND 0.3733f
C4270 XA.XIR[8].XIC[6].icell.Ien VGND 0.3733f
C4271 XA.XIR[8].XIC[5].icell.Ien VGND 0.3733f
C4272 XA.XIR[8].XIC[4].icell.Ien VGND 0.3733f
C4273 XA.XIR[8].XIC[3].icell.Ien VGND 0.3733f
C4274 XA.XIR[8].XIC[2].icell.Ien VGND 0.3733f
C4275 XA.XIR[8].XIC_dummy_left.icell.Iout VGND 0.80566f
C4276 XA.XIR[8].XIC[1].icell.Ien VGND 0.3733f
C4277 XThR.Tn[8] VGND 12.78722f
C4278 XA.XIR[8].XIC[0].icell.Ien VGND 0.37345f
C4279 XA.XIR[8].XIC_dummy_left.icell.SM VGND 0.01033f
C4280 XA.XIR[8].XIC_dummy_left.icell.Ien VGND 0.57308f
C4281 XA.XIR[8].XIC_dummy_right.icell.PDM VGND 0.23384f
C4282 XA.XIR[8].XIC_15.icell.PDM VGND 0.18862f
C4283 XA.XIR[8].XIC[14].icell.PDM VGND 0.1882f
C4284 XA.XIR[8].XIC[13].icell.PDM VGND 0.1882f
C4285 XA.XIR[8].XIC[12].icell.PDM VGND 0.1882f
C4286 XA.XIR[8].XIC[11].icell.PDM VGND 0.1882f
C4287 XA.XIR[8].XIC[10].icell.PDM VGND 0.1882f
C4288 XA.XIR[8].XIC[9].icell.PDM VGND 0.1882f
C4289 XA.XIR[8].XIC[8].icell.PDM VGND 0.1882f
C4290 XA.XIR[8].XIC[7].icell.PDM VGND 0.1882f
C4291 XA.XIR[8].XIC[6].icell.PDM VGND 0.1882f
C4292 XA.XIR[8].XIC[5].icell.PDM VGND 0.1882f
C4293 XA.XIR[8].XIC[4].icell.PDM VGND 0.1882f
C4294 XA.XIR[8].XIC[3].icell.PDM VGND 0.1882f
C4295 XA.XIR[8].XIC[2].icell.PDM VGND 0.1882f
C4296 XA.XIR[8].XIC[1].icell.PDM VGND 0.1882f
C4297 XA.XIR[8].XIC[0].icell.PDM VGND 0.18836f
C4298 XA.XIR[8].XIC_dummy_left.icell.PDM VGND 0.22809f
C4299 XA.XIR[7].XIC_dummy_right.icell.Iout VGND 0.85788f
C4300 XA.XIR[7].XIC_dummy_right.icell.SM VGND 0.01013f
C4301 XA.XIR[7].XIC_dummy_right.icell.Ien VGND 0.60818f
C4302 XA.XIR[7].XIC_15.icell.Ien VGND 0.37264f
C4303 XA.XIR[7].XIC[14].icell.Ien VGND 0.37333f
C4304 XA.XIR[7].XIC[13].icell.Ien VGND 0.3733f
C4305 XA.XIR[7].XIC[12].icell.Ien VGND 0.3733f
C4306 XA.XIR[7].XIC[11].icell.Ien VGND 0.3733f
C4307 XA.XIR[7].XIC[10].icell.Ien VGND 0.3733f
C4308 XA.XIR[7].XIC[9].icell.Ien VGND 0.3733f
C4309 XA.XIR[7].XIC[8].icell.Ien VGND 0.3733f
C4310 XA.XIR[7].XIC[7].icell.Ien VGND 0.3733f
C4311 XA.XIR[7].XIC[6].icell.Ien VGND 0.3733f
C4312 XA.XIR[7].XIC[5].icell.Ien VGND 0.3733f
C4313 XA.XIR[7].XIC[4].icell.Ien VGND 0.3733f
C4314 XA.XIR[7].XIC[3].icell.Ien VGND 0.3733f
C4315 XA.XIR[7].XIC[2].icell.Ien VGND 0.3733f
C4316 XA.XIR[7].XIC_dummy_left.icell.Iout VGND 0.80598f
C4317 XA.XIR[7].XIC[1].icell.Ien VGND 0.3733f
C4318 XA.XIR[7].XIC[0].icell.Ien VGND 0.37345f
C4319 XA.XIR[7].XIC_dummy_left.icell.SM VGND 0.01033f
C4320 XThR.Tn[7] VGND 13.23029f
C4321 XThR.XTBN.A VGND 1.22814f
C4322 XA.XIR[7].XIC_dummy_left.icell.Ien VGND 0.57576f
C4323 XA.XIR[7].XIC_dummy_right.icell.PDM VGND 0.23384f
C4324 XA.XIR[7].XIC_15.icell.PDM VGND 0.18862f
C4325 XA.XIR[7].XIC[14].icell.PDM VGND 0.1882f
C4326 XA.XIR[7].XIC[13].icell.PDM VGND 0.1882f
C4327 XA.XIR[7].XIC[12].icell.PDM VGND 0.1882f
C4328 XA.XIR[7].XIC[11].icell.PDM VGND 0.1882f
C4329 XA.XIR[7].XIC[10].icell.PDM VGND 0.1882f
C4330 XA.XIR[7].XIC[9].icell.PDM VGND 0.1882f
C4331 XA.XIR[7].XIC[8].icell.PDM VGND 0.1882f
C4332 XA.XIR[7].XIC[7].icell.PDM VGND 0.1882f
C4333 XA.XIR[7].XIC[6].icell.PDM VGND 0.1882f
C4334 XA.XIR[7].XIC[5].icell.PDM VGND 0.1882f
C4335 XA.XIR[7].XIC[4].icell.PDM VGND 0.1882f
C4336 XA.XIR[7].XIC[3].icell.PDM VGND 0.1882f
C4337 XA.XIR[7].XIC[2].icell.PDM VGND 0.1882f
C4338 XA.XIR[7].XIC[1].icell.PDM VGND 0.1882f
C4339 XA.XIR[7].XIC[0].icell.PDM VGND 0.18836f
C4340 XA.XIR[7].XIC_dummy_left.icell.PDM VGND 0.22809f
C4341 XA.XIR[6].XIC_dummy_right.icell.Iout VGND 0.85788f
C4342 XA.XIR[6].XIC_dummy_right.icell.SM VGND 0.01013f
C4343 XA.XIR[6].XIC_dummy_right.icell.Ien VGND 0.60818f
C4344 XA.XIR[6].XIC_15.icell.Ien VGND 0.37264f
C4345 XA.XIR[6].XIC[14].icell.Ien VGND 0.37333f
C4346 XA.XIR[6].XIC[13].icell.Ien VGND 0.3733f
C4347 XA.XIR[6].XIC[12].icell.Ien VGND 0.3733f
C4348 XA.XIR[6].XIC[11].icell.Ien VGND 0.3733f
C4349 XA.XIR[6].XIC[10].icell.Ien VGND 0.3733f
C4350 XA.XIR[6].XIC[9].icell.Ien VGND 0.3733f
C4351 XA.XIR[6].XIC[8].icell.Ien VGND 0.3733f
C4352 XA.XIR[6].XIC[7].icell.Ien VGND 0.3733f
C4353 XA.XIR[6].XIC[6].icell.Ien VGND 0.3733f
C4354 XA.XIR[6].XIC[5].icell.Ien VGND 0.3733f
C4355 XA.XIR[6].XIC[4].icell.Ien VGND 0.3733f
C4356 XA.XIR[6].XIC[3].icell.Ien VGND 0.3733f
C4357 XA.XIR[6].XIC[2].icell.Ien VGND 0.3733f
C4358 XA.XIR[6].XIC_dummy_left.icell.Iout VGND 0.80693f
C4359 XA.XIR[6].XIC[1].icell.Ien VGND 0.3733f
C4360 XA.XIR[6].XIC[0].icell.Ien VGND 0.37345f
C4361 XA.XIR[6].XIC_dummy_left.icell.SM VGND 0.01033f
C4362 XA.XIR[6].XIC_dummy_left.icell.Ien VGND 0.57422f
C4363 XThR.Tn[6] VGND 12.9018f
C4364 a_n1049_5317# VGND 0.02283f
C4365 XThR.XTB7.Y VGND 1.36132f
C4366 XA.XIR[6].XIC_dummy_right.icell.PDM VGND 0.23384f
C4367 XA.XIR[6].XIC_15.icell.PDM VGND 0.18862f
C4368 XA.XIR[6].XIC[14].icell.PDM VGND 0.1882f
C4369 XA.XIR[6].XIC[13].icell.PDM VGND 0.1882f
C4370 XA.XIR[6].XIC[12].icell.PDM VGND 0.1882f
C4371 XA.XIR[6].XIC[11].icell.PDM VGND 0.1882f
C4372 XA.XIR[6].XIC[10].icell.PDM VGND 0.1882f
C4373 XA.XIR[6].XIC[9].icell.PDM VGND 0.1882f
C4374 XA.XIR[6].XIC[8].icell.PDM VGND 0.1882f
C4375 XA.XIR[6].XIC[7].icell.PDM VGND 0.1882f
C4376 XA.XIR[6].XIC[6].icell.PDM VGND 0.1882f
C4377 XA.XIR[6].XIC[5].icell.PDM VGND 0.1882f
C4378 XA.XIR[6].XIC[4].icell.PDM VGND 0.1882f
C4379 XA.XIR[6].XIC[3].icell.PDM VGND 0.1882f
C4380 XA.XIR[6].XIC[2].icell.PDM VGND 0.1882f
C4381 XA.XIR[6].XIC[1].icell.PDM VGND 0.1882f
C4382 XA.XIR[6].XIC[0].icell.PDM VGND 0.18836f
C4383 XA.XIR[6].XIC_dummy_left.icell.PDM VGND 0.22809f
C4384 XA.XIR[5].XIC_dummy_right.icell.Iout VGND 0.85788f
C4385 XA.XIR[5].XIC_dummy_right.icell.SM VGND 0.01013f
C4386 XA.XIR[5].XIC_dummy_right.icell.Ien VGND 0.60818f
C4387 XA.XIR[5].XIC_15.icell.Ien VGND 0.37264f
C4388 XA.XIR[5].XIC[14].icell.Ien VGND 0.37333f
C4389 XA.XIR[5].XIC[13].icell.Ien VGND 0.3733f
C4390 XA.XIR[5].XIC[12].icell.Ien VGND 0.3733f
C4391 XA.XIR[5].XIC[11].icell.Ien VGND 0.3733f
C4392 XA.XIR[5].XIC[10].icell.Ien VGND 0.3733f
C4393 XA.XIR[5].XIC[9].icell.Ien VGND 0.3733f
C4394 XA.XIR[5].XIC[8].icell.Ien VGND 0.3733f
C4395 XA.XIR[5].XIC[7].icell.Ien VGND 0.3733f
C4396 XA.XIR[5].XIC[6].icell.Ien VGND 0.3733f
C4397 XA.XIR[5].XIC[5].icell.Ien VGND 0.3733f
C4398 XA.XIR[5].XIC[4].icell.Ien VGND 0.3733f
C4399 XA.XIR[5].XIC[3].icell.Ien VGND 0.3733f
C4400 XA.XIR[5].XIC[2].icell.Ien VGND 0.3733f
C4401 XA.XIR[5].XIC_dummy_left.icell.Iout VGND 0.80562f
C4402 XA.XIR[5].XIC[1].icell.Ien VGND 0.3733f
C4403 a_n1049_5611# VGND 0.02888f
C4404 XA.XIR[5].XIC[0].icell.Ien VGND 0.37345f
C4405 XA.XIR[5].XIC_dummy_left.icell.SM VGND 0.01033f
C4406 XA.XIR[5].XIC_dummy_left.icell.Ien VGND 0.57288f
C4407 XThR.Tn[5] VGND 12.89248f
C4408 XThR.XTB6.Y VGND 1.38212f
C4409 XA.XIR[5].XIC_dummy_right.icell.PDM VGND 0.23384f
C4410 XA.XIR[5].XIC_15.icell.PDM VGND 0.18862f
C4411 XA.XIR[5].XIC[14].icell.PDM VGND 0.1882f
C4412 XA.XIR[5].XIC[13].icell.PDM VGND 0.1882f
C4413 XA.XIR[5].XIC[12].icell.PDM VGND 0.1882f
C4414 XA.XIR[5].XIC[11].icell.PDM VGND 0.1882f
C4415 XA.XIR[5].XIC[10].icell.PDM VGND 0.1882f
C4416 XA.XIR[5].XIC[9].icell.PDM VGND 0.1882f
C4417 XA.XIR[5].XIC[8].icell.PDM VGND 0.1882f
C4418 XA.XIR[5].XIC[7].icell.PDM VGND 0.1882f
C4419 XA.XIR[5].XIC[6].icell.PDM VGND 0.1882f
C4420 XA.XIR[5].XIC[5].icell.PDM VGND 0.1882f
C4421 XA.XIR[5].XIC[4].icell.PDM VGND 0.1882f
C4422 XA.XIR[5].XIC[3].icell.PDM VGND 0.1882f
C4423 XA.XIR[5].XIC[2].icell.PDM VGND 0.1882f
C4424 XA.XIR[5].XIC[1].icell.PDM VGND 0.1882f
C4425 XA.XIR[5].XIC[0].icell.PDM VGND 0.18836f
C4426 XA.XIR[5].XIC_dummy_left.icell.PDM VGND 0.22809f
C4427 XA.XIR[4].XIC_dummy_right.icell.Iout VGND 0.85788f
C4428 XA.XIR[4].XIC_dummy_right.icell.SM VGND 0.01013f
C4429 XA.XIR[4].XIC_dummy_right.icell.Ien VGND 0.60818f
C4430 XA.XIR[4].XIC_15.icell.Ien VGND 0.37264f
C4431 XA.XIR[4].XIC[14].icell.Ien VGND 0.37333f
C4432 XA.XIR[4].XIC[13].icell.Ien VGND 0.3733f
C4433 XA.XIR[4].XIC[12].icell.Ien VGND 0.3733f
C4434 XA.XIR[4].XIC[11].icell.Ien VGND 0.3733f
C4435 XA.XIR[4].XIC[10].icell.Ien VGND 0.3733f
C4436 XA.XIR[4].XIC[9].icell.Ien VGND 0.3733f
C4437 XA.XIR[4].XIC[8].icell.Ien VGND 0.3733f
C4438 XA.XIR[4].XIC[7].icell.Ien VGND 0.3733f
C4439 XA.XIR[4].XIC[6].icell.Ien VGND 0.3733f
C4440 XA.XIR[4].XIC[5].icell.Ien VGND 0.3733f
C4441 XA.XIR[4].XIC[4].icell.Ien VGND 0.3733f
C4442 XA.XIR[4].XIC[3].icell.Ien VGND 0.3733f
C4443 XA.XIR[4].XIC[2].icell.Ien VGND 0.3733f
C4444 XA.XIR[4].XIC_dummy_left.icell.Iout VGND 0.80734f
C4445 XA.XIR[4].XIC[1].icell.Ien VGND 0.3733f
C4446 XA.XIR[4].XIC[0].icell.Ien VGND 0.37345f
C4447 XA.XIR[4].XIC_dummy_left.icell.SM VGND 0.01033f
C4448 XA.XIR[4].XIC_dummy_left.icell.Ien VGND 0.57333f
C4449 XA.XIR[4].XIC_dummy_right.icell.PDM VGND 0.23384f
C4450 XA.XIR[4].XIC_15.icell.PDM VGND 0.18862f
C4451 XA.XIR[4].XIC[14].icell.PDM VGND 0.1882f
C4452 XA.XIR[4].XIC[13].icell.PDM VGND 0.1882f
C4453 XA.XIR[4].XIC[12].icell.PDM VGND 0.1882f
C4454 XA.XIR[4].XIC[11].icell.PDM VGND 0.1882f
C4455 XA.XIR[4].XIC[10].icell.PDM VGND 0.1882f
C4456 XA.XIR[4].XIC[9].icell.PDM VGND 0.1882f
C4457 XA.XIR[4].XIC[8].icell.PDM VGND 0.1882f
C4458 XA.XIR[4].XIC[7].icell.PDM VGND 0.1882f
C4459 XA.XIR[4].XIC[6].icell.PDM VGND 0.1882f
C4460 XA.XIR[4].XIC[5].icell.PDM VGND 0.1882f
C4461 XA.XIR[4].XIC[4].icell.PDM VGND 0.1882f
C4462 XA.XIR[4].XIC[3].icell.PDM VGND 0.1882f
C4463 XA.XIR[4].XIC[2].icell.PDM VGND 0.1882f
C4464 XA.XIR[4].XIC[1].icell.PDM VGND 0.1882f
C4465 XA.XIR[4].XIC[0].icell.PDM VGND 0.18836f
C4466 XA.XIR[4].XIC_dummy_left.icell.PDM VGND 0.22809f
C4467 XThR.Tn[4] VGND 12.95212f
C4468 a_n1049_6405# VGND 0.02935f
C4469 XA.XIR[3].XIC_dummy_right.icell.Iout VGND 0.85788f
C4470 XA.XIR[3].XIC_dummy_right.icell.SM VGND 0.01013f
C4471 XA.XIR[3].XIC_dummy_right.icell.Ien VGND 0.60818f
C4472 XA.XIR[3].XIC_15.icell.Ien VGND 0.37264f
C4473 XA.XIR[3].XIC[14].icell.Ien VGND 0.37333f
C4474 XA.XIR[3].XIC[13].icell.Ien VGND 0.3733f
C4475 XA.XIR[3].XIC[12].icell.Ien VGND 0.3733f
C4476 XA.XIR[3].XIC[11].icell.Ien VGND 0.3733f
C4477 XA.XIR[3].XIC[10].icell.Ien VGND 0.3733f
C4478 XA.XIR[3].XIC[9].icell.Ien VGND 0.3733f
C4479 XA.XIR[3].XIC[8].icell.Ien VGND 0.3733f
C4480 XA.XIR[3].XIC[7].icell.Ien VGND 0.3733f
C4481 XA.XIR[3].XIC[6].icell.Ien VGND 0.3733f
C4482 XA.XIR[3].XIC[5].icell.Ien VGND 0.3733f
C4483 XA.XIR[3].XIC[4].icell.Ien VGND 0.3733f
C4484 XA.XIR[3].XIC[3].icell.Ien VGND 0.3733f
C4485 XA.XIR[3].XIC[2].icell.Ien VGND 0.3733f
C4486 XThR.XTB5.Y VGND 1.32753f
C4487 XA.XIR[3].XIC_dummy_left.icell.Iout VGND 0.80575f
C4488 XA.XIR[3].XIC[1].icell.Ien VGND 0.3733f
C4489 XA.XIR[3].XIC[0].icell.Ien VGND 0.37345f
C4490 XA.XIR[3].XIC_dummy_left.icell.SM VGND 0.01033f
C4491 XA.XIR[3].XIC_dummy_left.icell.Ien VGND 0.57422f
C4492 a_n1049_6699# VGND 0.02979f
C4493 XA.XIR[3].XIC_dummy_right.icell.PDM VGND 0.23384f
C4494 XA.XIR[3].XIC_15.icell.PDM VGND 0.18862f
C4495 XA.XIR[3].XIC[14].icell.PDM VGND 0.1882f
C4496 XA.XIR[3].XIC[13].icell.PDM VGND 0.1882f
C4497 XA.XIR[3].XIC[12].icell.PDM VGND 0.1882f
C4498 XA.XIR[3].XIC[11].icell.PDM VGND 0.1882f
C4499 XA.XIR[3].XIC[10].icell.PDM VGND 0.1882f
C4500 XA.XIR[3].XIC[9].icell.PDM VGND 0.1882f
C4501 XA.XIR[3].XIC[8].icell.PDM VGND 0.1882f
C4502 XA.XIR[3].XIC[7].icell.PDM VGND 0.1882f
C4503 XA.XIR[3].XIC[6].icell.PDM VGND 0.1882f
C4504 XA.XIR[3].XIC[5].icell.PDM VGND 0.1882f
C4505 XA.XIR[3].XIC[4].icell.PDM VGND 0.1882f
C4506 XA.XIR[3].XIC[3].icell.PDM VGND 0.1882f
C4507 XA.XIR[3].XIC[2].icell.PDM VGND 0.1882f
C4508 XA.XIR[3].XIC[1].icell.PDM VGND 0.1882f
C4509 XA.XIR[3].XIC[0].icell.PDM VGND 0.18836f
C4510 XA.XIR[3].XIC_dummy_left.icell.PDM VGND 0.22809f
C4511 XA.XIR[2].XIC_dummy_right.icell.Iout VGND 0.85788f
C4512 XA.XIR[2].XIC_dummy_right.icell.SM VGND 0.01013f
C4513 XA.XIR[2].XIC_dummy_right.icell.Ien VGND 0.60818f
C4514 XA.XIR[2].XIC_15.icell.Ien VGND 0.37264f
C4515 XA.XIR[2].XIC[14].icell.Ien VGND 0.37333f
C4516 XA.XIR[2].XIC[13].icell.Ien VGND 0.3733f
C4517 XA.XIR[2].XIC[12].icell.Ien VGND 0.3733f
C4518 XA.XIR[2].XIC[11].icell.Ien VGND 0.3733f
C4519 XA.XIR[2].XIC[10].icell.Ien VGND 0.3733f
C4520 XA.XIR[2].XIC[9].icell.Ien VGND 0.3733f
C4521 XA.XIR[2].XIC[8].icell.Ien VGND 0.3733f
C4522 XA.XIR[2].XIC[7].icell.Ien VGND 0.3733f
C4523 XA.XIR[2].XIC[6].icell.Ien VGND 0.3733f
C4524 XA.XIR[2].XIC[5].icell.Ien VGND 0.3733f
C4525 XA.XIR[2].XIC[4].icell.Ien VGND 0.3733f
C4526 XA.XIR[2].XIC[3].icell.Ien VGND 0.3733f
C4527 XA.XIR[2].XIC[2].icell.Ien VGND 0.3733f
C4528 XA.XIR[2].XIC_dummy_left.icell.Iout VGND 0.80789f
C4529 XA.XIR[2].XIC[1].icell.Ien VGND 0.3733f
C4530 XThR.Tn[3] VGND 12.94485f
C4531 XThR.XTB4.Y VGND 1.48815f
C4532 XA.XIR[2].XIC[0].icell.Ien VGND 0.37345f
C4533 XA.XIR[2].XIC_dummy_left.icell.SM VGND 0.01033f
C4534 XA.XIR[2].XIC_dummy_left.icell.Ien VGND 0.57556f
C4535 XA.XIR[2].XIC_dummy_right.icell.PDM VGND 0.23384f
C4536 XA.XIR[2].XIC_15.icell.PDM VGND 0.18862f
C4537 XA.XIR[2].XIC[14].icell.PDM VGND 0.1882f
C4538 XA.XIR[2].XIC[13].icell.PDM VGND 0.1882f
C4539 XA.XIR[2].XIC[12].icell.PDM VGND 0.1882f
C4540 XA.XIR[2].XIC[11].icell.PDM VGND 0.1882f
C4541 XA.XIR[2].XIC[10].icell.PDM VGND 0.1882f
C4542 XA.XIR[2].XIC[9].icell.PDM VGND 0.1882f
C4543 XA.XIR[2].XIC[8].icell.PDM VGND 0.1882f
C4544 XA.XIR[2].XIC[7].icell.PDM VGND 0.1882f
C4545 XA.XIR[2].XIC[6].icell.PDM VGND 0.1882f
C4546 XA.XIR[2].XIC[5].icell.PDM VGND 0.1882f
C4547 XA.XIR[2].XIC[4].icell.PDM VGND 0.1882f
C4548 XA.XIR[2].XIC[3].icell.PDM VGND 0.1882f
C4549 XA.XIR[2].XIC[2].icell.PDM VGND 0.1882f
C4550 XA.XIR[2].XIC[1].icell.PDM VGND 0.1882f
C4551 XA.XIR[2].XIC[0].icell.PDM VGND 0.18836f
C4552 XA.XIR[2].XIC_dummy_left.icell.PDM VGND 0.22809f
C4553 XA.XIR[1].XIC_dummy_right.icell.Iout VGND 0.85788f
C4554 XA.XIR[1].XIC_dummy_right.icell.SM VGND 0.01013f
C4555 XA.XIR[1].XIC_dummy_right.icell.Ien VGND 0.60818f
C4556 XA.XIR[1].XIC_15.icell.Ien VGND 0.37264f
C4557 XA.XIR[1].XIC[14].icell.Ien VGND 0.37333f
C4558 XA.XIR[1].XIC[13].icell.Ien VGND 0.3733f
C4559 XA.XIR[1].XIC[12].icell.Ien VGND 0.3733f
C4560 XA.XIR[1].XIC[11].icell.Ien VGND 0.3733f
C4561 XA.XIR[1].XIC[10].icell.Ien VGND 0.3733f
C4562 XA.XIR[1].XIC[9].icell.Ien VGND 0.3733f
C4563 XA.XIR[1].XIC[8].icell.Ien VGND 0.3733f
C4564 XA.XIR[1].XIC[7].icell.Ien VGND 0.3733f
C4565 XA.XIR[1].XIC[6].icell.Ien VGND 0.3733f
C4566 XA.XIR[1].XIC[5].icell.Ien VGND 0.3733f
C4567 XA.XIR[1].XIC[4].icell.Ien VGND 0.3733f
C4568 XA.XIR[1].XIC[3].icell.Ien VGND 0.3733f
C4569 XA.XIR[1].XIC[2].icell.Ien VGND 0.3733f
C4570 XA.XIR[1].XIC_dummy_left.icell.Iout VGND 0.80575f
C4571 XA.XIR[1].XIC[1].icell.Ien VGND 0.3733f
C4572 XThR.Tn[2] VGND 12.94933f
C4573 a_n1049_7493# VGND 0.02484f
C4574 XThR.XTB3.Y VGND 2.09162f
C4575 XThR.XTB7.A VGND 1.95537f
C4576 XA.XIR[1].XIC[0].icell.Ien VGND 0.37345f
C4577 XA.XIR[1].XIC_dummy_left.icell.SM VGND 0.01033f
C4578 XA.XIR[1].XIC_dummy_left.icell.Ien VGND 0.57375f
C4579 XA.XIR[1].XIC_dummy_right.icell.PDM VGND 0.23384f
C4580 XA.XIR[1].XIC_15.icell.PDM VGND 0.18862f
C4581 XA.XIR[1].XIC[14].icell.PDM VGND 0.1882f
C4582 XA.XIR[1].XIC[13].icell.PDM VGND 0.1882f
C4583 XA.XIR[1].XIC[12].icell.PDM VGND 0.1882f
C4584 XA.XIR[1].XIC[11].icell.PDM VGND 0.1882f
C4585 XA.XIR[1].XIC[10].icell.PDM VGND 0.1882f
C4586 XA.XIR[1].XIC[9].icell.PDM VGND 0.1882f
C4587 XA.XIR[1].XIC[8].icell.PDM VGND 0.1882f
C4588 XA.XIR[1].XIC[7].icell.PDM VGND 0.1882f
C4589 XA.XIR[1].XIC[6].icell.PDM VGND 0.1882f
C4590 XA.XIR[1].XIC[5].icell.PDM VGND 0.1882f
C4591 XA.XIR[1].XIC[4].icell.PDM VGND 0.1882f
C4592 XA.XIR[1].XIC[3].icell.PDM VGND 0.1882f
C4593 XA.XIR[1].XIC[2].icell.PDM VGND 0.1882f
C4594 XA.XIR[1].XIC[1].icell.PDM VGND 0.1882f
C4595 XA.XIR[1].XIC[0].icell.PDM VGND 0.18836f
C4596 XA.XIR[1].XIC_dummy_left.icell.PDM VGND 0.22809f
C4597 a_n1049_7787# VGND 0.03396f
C4598 XA.XIR[0].XIC_dummy_right.icell.Iout VGND 0.87403f
C4599 XA.XIR[0].XIC_dummy_right.icell.SM VGND 0.01013f
C4600 XA.XIR[0].XIC_dummy_right.icell.Ien VGND 0.61797f
C4601 XA.XIR[0].XIC_15.icell.Ien VGND 0.37874f
C4602 XA.XIR[0].XIC[14].icell.Ien VGND 0.39158f
C4603 XA.XIR[0].XIC[13].icell.Ien VGND 0.39155f
C4604 XA.XIR[0].XIC[12].icell.Ien VGND 0.38822f
C4605 XA.XIR[0].XIC[11].icell.Ien VGND 0.3889f
C4606 XA.XIR[0].XIC[10].icell.Ien VGND 0.39022f
C4607 XA.XIR[0].XIC[9].icell.Ien VGND 0.3885f
C4608 XA.XIR[0].XIC[8].icell.Ien VGND 0.38898f
C4609 XA.XIR[0].XIC[7].icell.Ien VGND 0.38927f
C4610 XA.XIR[0].XIC[6].icell.Ien VGND 0.38927f
C4611 XA.XIR[0].XIC[5].icell.Ien VGND 0.38822f
C4612 XA.XIR[0].XIC[4].icell.Ien VGND 0.38827f
C4613 XA.XIR[0].XIC[3].icell.Ien VGND 0.38951f
C4614 XA.XIR[0].XIC[2].icell.Ien VGND 0.39155f
C4615 XA.XIR[0].XIC_dummy_left.icell.Iout VGND 0.83189f
C4616 XA.XIR[0].XIC[1].icell.Ien VGND 0.39155f
C4617 XA.XIR[0].XIC[0].icell.Ien VGND 0.39085f
C4618 XA.XIR[0].XIC_dummy_left.icell.SM VGND 0.01033f
C4619 XThR.Tn[1] VGND 12.98858f
C4620 XThR.XTB2.Y VGND 1.4743f
C4621 XThR.XTB6.A VGND 0.95418f
C4622 XA.XIR[0].XIC_dummy_left.icell.Ien VGND 0.58648f
C4623 XA.XIR[0].XIC_dummy_right.icell.PDM VGND 0.251f
C4624 XA.XIR[0].XIC_15.icell.PDM VGND 0.20773f
C4625 XA.XIR[0].XIC[14].icell.PDM VGND 0.24601f
C4626 XA.XIR[0].XIC[13].icell.PDM VGND 0.24585f
C4627 XA.XIR[0].XIC[12].icell.PDM VGND 0.24146f
C4628 XA.XIR[0].XIC[11].icell.PDM VGND 0.24184f
C4629 XA.XIR[0].XIC[10].icell.PDM VGND 0.24174f
C4630 XA.XIR[0].XIC[9].icell.PDM VGND 0.24147f
C4631 XA.XIR[0].XIC[8].icell.PDM VGND 0.24147f
C4632 XA.XIR[0].XIC[7].icell.PDM VGND 0.2442f
C4633 XA.XIR[0].XIC[6].icell.PDM VGND 0.24156f
C4634 XA.XIR[0].XIC[5].icell.PDM VGND 0.24321f
C4635 XA.XIR[0].XIC[4].icell.PDM VGND 0.24159f
C4636 XA.XIR[0].XIC[3].icell.PDM VGND 0.24451f
C4637 XA.XIR[0].XIC[2].icell.PDM VGND 0.2458f
C4638 XA.XIR[0].XIC[1].icell.PDM VGND 0.2458f
C4639 XA.XIR[0].XIC[0].icell.PDM VGND 0.24486f
C4640 XA.XIR[0].XIC_dummy_left.icell.PDM VGND 0.25065f
C4641 XThR.Tn[0] VGND 13.29109f
C4642 a_n1049_8581# VGND 0.0432f
C4643 XThR.XTBN.Y VGND 7.77528f
C4644 XThR.XTB1.Y VGND 1.80882f
C4645 XThR.XTB7.B VGND 2.60708f
C4646 XThR.XTB5.A VGND 1.75667f
C4647 XThC.Tn[14] VGND 5.52615f
C4648 XThC.Tn[13] VGND 5.16689f
C4649 XThC.Tn[12] VGND 5.1562f
C4650 XThC.Tn[11] VGND 5.52379f
C4651 XThC.Tn[10] VGND 5.0515f
C4652 XThC.Tn[9] VGND 5.34336f
C4653 XThC.Tn[8] VGND 4.89287f
C4654 a_10915_9569# VGND 0.55912f
C4655 a_10051_9569# VGND 0.55747f
C4656 a_9827_9569# VGND 0.54584f
C4657 a_8963_9569# VGND 0.55439f
C4658 a_8739_9569# VGND 0.553f
C4659 a_7875_9569# VGND 0.55432f
C4660 a_7651_9569# VGND 0.55717f
C4661 XThC.Tn[7] VGND 5.47379f
C4662 XThC.Tn[6] VGND 5.48958f
C4663 XThC.Tn[5] VGND 5.60438f
C4664 XThC.Tn[4] VGND 5.55465f
C4665 XThC.Tn[3] VGND 5.88113f
C4666 XThC.Tn[2] VGND 5.58434f
C4667 XThC.Tn[1] VGND 5.71884f
C4668 XThC.Tn[0] VGND 6.85356f
C4669 a_6243_9615# VGND 0.03028f
C4670 a_5949_9615# VGND 0.03456f
C4671 a_5155_9615# VGND 0.03624f
C4672 a_4861_9615# VGND 0.03647f
C4673 a_4067_9615# VGND 0.03118f
C4674 a_3773_9615# VGND 0.03896f
C4675 a_2979_9615# VGND 0.04122f
C4676 XThC.XTBN.Y VGND 8.71712f
C4677 XThC.XTB7.Y VGND 1.35988f
C4678 XThC.XTB6.Y VGND 1.3794f
C4679 XThC.XTB7.B VGND 2.83799f
C4680 XThC.XTB5.Y VGND 1.32558f
C4681 XThC.XTBN.A VGND 1.2246f
C4682 XThC.XTB4.Y VGND 1.6934f
C4683 XThC.XTB3.Y VGND 1.96717f
C4684 XThC.XTB7.A VGND 1.94951f
C4685 XThC.XTB6.A VGND 0.95452f
C4686 XThC.XTB2.Y VGND 1.4752f
C4687 XThC.XTB1.Y VGND 1.77643f
C4688 XThC.XTB5.A VGND 1.75974f
C4689 bias[0].t0 VGND 0.86609f
C4690 bias[0].n0 VGND 0.31538f
C4691 bias[0].n1 VGND 0.22269f
C4692 bias[0].t1 VGND 0.86609f
C4693 bias[0].n2 VGND 0.33687f
C4694 XThR.XTB3.Y.t1 VGND 0.06176f
C4695 XThR.XTB3.Y.n0 VGND 0.01521f
C4696 XThR.XTB3.Y.t8 VGND 0.04903f
C4697 XThR.XTB3.Y.t15 VGND 0.02889f
C4698 XThR.XTB3.Y.t13 VGND 0.04903f
C4699 XThR.XTB3.Y.t6 VGND 0.02889f
C4700 XThR.XTB3.Y.t9 VGND 0.04903f
C4701 XThR.XTB3.Y.t17 VGND 0.02889f
C4702 XThR.XTB3.Y.n1 VGND 0.08226f
C4703 XThR.XTB3.Y.n2 VGND 0.08688f
C4704 XThR.XTB3.Y.n3 VGND 0.03573f
C4705 XThR.XTB3.Y.n4 VGND 0.0707f
C4706 XThR.XTB3.Y.t12 VGND 0.04903f
C4707 XThR.XTB3.Y.t4 VGND 0.02889f
C4708 XThR.XTB3.Y.n5 VGND 0.06608f
C4709 XThR.XTB3.Y.n6 VGND 0.03236f
C4710 XThR.XTB3.Y.n7 VGND 0.02685f
C4711 XThR.XTB3.Y.t18 VGND 0.04903f
C4712 XThR.XTB3.Y.t5 VGND 0.02889f
C4713 XThR.XTB3.Y.n8 VGND 0.03005f
C4714 XThR.XTB3.Y.t7 VGND 0.04903f
C4715 XThR.XTB3.Y.t10 VGND 0.02889f
C4716 XThR.XTB3.Y.n9 VGND 0.05992f
C4717 XThR.XTB3.Y.t11 VGND 0.04903f
C4718 XThR.XTB3.Y.t16 VGND 0.02889f
C4719 XThR.XTB3.Y.n10 VGND 0.06454f
C4720 XThR.XTB3.Y.n11 VGND 0.03645f
C4721 XThR.XTB3.Y.n12 VGND 0.06034f
C4722 XThR.XTB3.Y.n13 VGND 0.03128f
C4723 XThR.XTB3.Y.n14 VGND 0.02851f
C4724 XThR.XTB3.Y.n15 VGND 0.06454f
C4725 XThR.XTB3.Y.t14 VGND 0.04903f
C4726 XThR.XTB3.Y.t3 VGND 0.02889f
C4727 XThR.XTB3.Y.n16 VGND 0.05838f
C4728 XThR.XTB3.Y.n17 VGND 0.03236f
C4729 XThR.XTB3.Y.n18 VGND 0.04707f
C4730 XThR.XTB3.Y.n19 VGND 1.31347f
C4731 XThR.XTB3.Y.t0 VGND 0.03152f
C4732 XThR.XTB3.Y.t2 VGND 0.03152f
C4733 XThR.XTB3.Y.n20 VGND 0.06766f
C4734 XThR.XTB3.Y.n21 VGND 0.157f
C4735 XThR.XTB3.Y.n22 VGND 0.03296f
C4736 XThR.XTB1.Y.t1 VGND 0.03165f
C4737 XThR.XTB1.Y.t8 VGND 0.02512f
C4738 XThR.XTB1.Y.t15 VGND 0.0148f
C4739 XThR.XTB1.Y.t14 VGND 0.02512f
C4740 XThR.XTB1.Y.t7 VGND 0.0148f
C4741 XThR.XTB1.Y.t10 VGND 0.02512f
C4742 XThR.XTB1.Y.t18 VGND 0.0148f
C4743 XThR.XTB1.Y.n1 VGND 0.04215f
C4744 XThR.XTB1.Y.n2 VGND 0.04452f
C4745 XThR.XTB1.Y.n3 VGND 0.01831f
C4746 XThR.XTB1.Y.n4 VGND 0.03623f
C4747 XThR.XTB1.Y.t13 VGND 0.02512f
C4748 XThR.XTB1.Y.t4 VGND 0.0148f
C4749 XThR.XTB1.Y.n5 VGND 0.03386f
C4750 XThR.XTB1.Y.n6 VGND 0.01658f
C4751 XThR.XTB1.Y.n7 VGND 0.01376f
C4752 XThR.XTB1.Y.t6 VGND 0.02512f
C4753 XThR.XTB1.Y.t11 VGND 0.0148f
C4754 XThR.XTB1.Y.n8 VGND 0.0154f
C4755 XThR.XTB1.Y.t12 VGND 0.02512f
C4756 XThR.XTB1.Y.t16 VGND 0.0148f
C4757 XThR.XTB1.Y.n9 VGND 0.0307f
C4758 XThR.XTB1.Y.t17 VGND 0.02512f
C4759 XThR.XTB1.Y.t5 VGND 0.0148f
C4760 XThR.XTB1.Y.n10 VGND 0.03307f
C4761 XThR.XTB1.Y.n11 VGND 0.01868f
C4762 XThR.XTB1.Y.n12 VGND 0.03092f
C4763 XThR.XTB1.Y.n13 VGND 0.01603f
C4764 XThR.XTB1.Y.n14 VGND 0.01461f
C4765 XThR.XTB1.Y.n15 VGND 0.03307f
C4766 XThR.XTB1.Y.t3 VGND 0.02512f
C4767 XThR.XTB1.Y.t9 VGND 0.0148f
C4768 XThR.XTB1.Y.n16 VGND 0.02991f
C4769 XThR.XTB1.Y.n17 VGND 0.01658f
C4770 XThR.XTB1.Y.n18 VGND 0.02412f
C4771 XThR.XTB1.Y.n19 VGND 0.75219f
C4772 XThR.XTB1.Y.t0 VGND 0.01615f
C4773 XThR.XTB1.Y.t2 VGND 0.01615f
C4774 XThR.XTB1.Y.n20 VGND 0.03467f
C4775 XThR.XTB1.Y.n21 VGND 0.08068f
C4776 XThR.XTB1.Y.n22 VGND 0.01689f
C4777 XThR.Tn[13].t2 VGND 0.01241f
C4778 XThR.Tn[13].t0 VGND 0.01241f
C4779 XThR.Tn[13].n0 VGND 0.02481f
C4780 XThR.Tn[13].t3 VGND 0.01241f
C4781 XThR.Tn[13].t1 VGND 0.01241f
C4782 XThR.Tn[13].n1 VGND 0.03094f
C4783 XThR.Tn[13].n2 VGND 0.06242f
C4784 XThR.Tn[13].t9 VGND 0.01909f
C4785 XThR.Tn[13].t11 VGND 0.01909f
C4786 XThR.Tn[13].n3 VGND 0.05796f
C4787 XThR.Tn[13].t10 VGND 0.01909f
C4788 XThR.Tn[13].t8 VGND 0.01909f
C4789 XThR.Tn[13].n4 VGND 0.04243f
C4790 XThR.Tn[13].n5 VGND 0.19293f
C4791 XThR.Tn[13].t6 VGND 0.01909f
C4792 XThR.Tn[13].t4 VGND 0.01909f
C4793 XThR.Tn[13].n6 VGND 0.04124f
C4794 XThR.Tn[13].t7 VGND 0.01909f
C4795 XThR.Tn[13].t5 VGND 0.01909f
C4796 XThR.Tn[13].n7 VGND 0.06277f
C4797 XThR.Tn[13].n8 VGND 0.17429f
C4798 XThR.Tn[13].n9 VGND 0.02334f
C4799 XThR.Tn[13].t72 VGND 0.01492f
C4800 XThR.Tn[13].t64 VGND 0.01633f
C4801 XThR.Tn[13].n10 VGND 0.03989f
C4802 XThR.Tn[13].n11 VGND 0.07663f
C4803 XThR.Tn[13].t28 VGND 0.01492f
C4804 XThR.Tn[13].t21 VGND 0.01633f
C4805 XThR.Tn[13].n12 VGND 0.03989f
C4806 XThR.Tn[13].t44 VGND 0.01487f
C4807 XThR.Tn[13].t12 VGND 0.01628f
C4808 XThR.Tn[13].n13 VGND 0.0415f
C4809 XThR.Tn[13].n14 VGND 0.02916f
C4810 XThR.Tn[13].n16 VGND 0.09357f
C4811 XThR.Tn[13].t65 VGND 0.01492f
C4812 XThR.Tn[13].t57 VGND 0.01633f
C4813 XThR.Tn[13].n17 VGND 0.03989f
C4814 XThR.Tn[13].t19 VGND 0.01487f
C4815 XThR.Tn[13].t52 VGND 0.01628f
C4816 XThR.Tn[13].n18 VGND 0.0415f
C4817 XThR.Tn[13].n19 VGND 0.02916f
C4818 XThR.Tn[13].n21 VGND 0.09357f
C4819 XThR.Tn[13].t22 VGND 0.01492f
C4820 XThR.Tn[13].t14 VGND 0.01633f
C4821 XThR.Tn[13].n22 VGND 0.03989f
C4822 XThR.Tn[13].t34 VGND 0.01487f
C4823 XThR.Tn[13].t70 VGND 0.01628f
C4824 XThR.Tn[13].n23 VGND 0.0415f
C4825 XThR.Tn[13].n24 VGND 0.02916f
C4826 XThR.Tn[13].n26 VGND 0.09357f
C4827 XThR.Tn[13].t49 VGND 0.01492f
C4828 XThR.Tn[13].t39 VGND 0.01633f
C4829 XThR.Tn[13].n27 VGND 0.03989f
C4830 XThR.Tn[13].t66 VGND 0.01487f
C4831 XThR.Tn[13].t35 VGND 0.01628f
C4832 XThR.Tn[13].n28 VGND 0.0415f
C4833 XThR.Tn[13].n29 VGND 0.02916f
C4834 XThR.Tn[13].n31 VGND 0.09357f
C4835 XThR.Tn[13].t24 VGND 0.01492f
C4836 XThR.Tn[13].t16 VGND 0.01633f
C4837 XThR.Tn[13].n32 VGND 0.03989f
C4838 XThR.Tn[13].t37 VGND 0.01487f
C4839 XThR.Tn[13].t71 VGND 0.01628f
C4840 XThR.Tn[13].n33 VGND 0.0415f
C4841 XThR.Tn[13].n34 VGND 0.02916f
C4842 XThR.Tn[13].n36 VGND 0.09357f
C4843 XThR.Tn[13].t60 VGND 0.01492f
C4844 XThR.Tn[13].t30 VGND 0.01633f
C4845 XThR.Tn[13].n37 VGND 0.03989f
C4846 XThR.Tn[13].t13 VGND 0.01487f
C4847 XThR.Tn[13].t26 VGND 0.01628f
C4848 XThR.Tn[13].n38 VGND 0.0415f
C4849 XThR.Tn[13].n39 VGND 0.02916f
C4850 XThR.Tn[13].n41 VGND 0.09357f
C4851 XThR.Tn[13].t29 VGND 0.01492f
C4852 XThR.Tn[13].t25 VGND 0.01633f
C4853 XThR.Tn[13].n42 VGND 0.03989f
C4854 XThR.Tn[13].t43 VGND 0.01487f
C4855 XThR.Tn[13].t18 VGND 0.01628f
C4856 XThR.Tn[13].n43 VGND 0.0415f
C4857 XThR.Tn[13].n44 VGND 0.02916f
C4858 XThR.Tn[13].n46 VGND 0.09357f
C4859 XThR.Tn[13].t32 VGND 0.01492f
C4860 XThR.Tn[13].t38 VGND 0.01633f
C4861 XThR.Tn[13].n47 VGND 0.03989f
C4862 XThR.Tn[13].t48 VGND 0.01487f
C4863 XThR.Tn[13].t33 VGND 0.01628f
C4864 XThR.Tn[13].n48 VGND 0.0415f
C4865 XThR.Tn[13].n49 VGND 0.02916f
C4866 XThR.Tn[13].n51 VGND 0.09357f
C4867 XThR.Tn[13].t51 VGND 0.01492f
C4868 XThR.Tn[13].t59 VGND 0.01633f
C4869 XThR.Tn[13].n52 VGND 0.03989f
C4870 XThR.Tn[13].t68 VGND 0.01487f
C4871 XThR.Tn[13].t53 VGND 0.01628f
C4872 XThR.Tn[13].n53 VGND 0.0415f
C4873 XThR.Tn[13].n54 VGND 0.02916f
C4874 XThR.Tn[13].n56 VGND 0.09357f
C4875 XThR.Tn[13].t41 VGND 0.01492f
C4876 XThR.Tn[13].t17 VGND 0.01633f
C4877 XThR.Tn[13].n57 VGND 0.03989f
C4878 XThR.Tn[13].t58 VGND 0.01487f
C4879 XThR.Tn[13].t73 VGND 0.01628f
C4880 XThR.Tn[13].n58 VGND 0.0415f
C4881 XThR.Tn[13].n59 VGND 0.02916f
C4882 XThR.Tn[13].n61 VGND 0.09357f
C4883 XThR.Tn[13].t63 VGND 0.01492f
C4884 XThR.Tn[13].t55 VGND 0.01633f
C4885 XThR.Tn[13].n62 VGND 0.03989f
C4886 XThR.Tn[13].t15 VGND 0.01487f
C4887 XThR.Tn[13].t45 VGND 0.01628f
C4888 XThR.Tn[13].n63 VGND 0.0415f
C4889 XThR.Tn[13].n64 VGND 0.02916f
C4890 XThR.Tn[13].n66 VGND 0.09357f
C4891 XThR.Tn[13].t31 VGND 0.01492f
C4892 XThR.Tn[13].t27 VGND 0.01633f
C4893 XThR.Tn[13].n67 VGND 0.03989f
C4894 XThR.Tn[13].t46 VGND 0.01487f
C4895 XThR.Tn[13].t20 VGND 0.01628f
C4896 XThR.Tn[13].n68 VGND 0.0415f
C4897 XThR.Tn[13].n69 VGND 0.02916f
C4898 XThR.Tn[13].n71 VGND 0.09357f
C4899 XThR.Tn[13].t50 VGND 0.01492f
C4900 XThR.Tn[13].t40 VGND 0.01633f
C4901 XThR.Tn[13].n72 VGND 0.03989f
C4902 XThR.Tn[13].t67 VGND 0.01487f
C4903 XThR.Tn[13].t36 VGND 0.01628f
C4904 XThR.Tn[13].n73 VGND 0.0415f
C4905 XThR.Tn[13].n74 VGND 0.02916f
C4906 XThR.Tn[13].n76 VGND 0.09357f
C4907 XThR.Tn[13].t69 VGND 0.01492f
C4908 XThR.Tn[13].t62 VGND 0.01633f
C4909 XThR.Tn[13].n77 VGND 0.03989f
C4910 XThR.Tn[13].t23 VGND 0.01487f
C4911 XThR.Tn[13].t54 VGND 0.01628f
C4912 XThR.Tn[13].n78 VGND 0.0415f
C4913 XThR.Tn[13].n79 VGND 0.02916f
C4914 XThR.Tn[13].n81 VGND 0.09357f
C4915 XThR.Tn[13].t42 VGND 0.01492f
C4916 XThR.Tn[13].t56 VGND 0.01633f
C4917 XThR.Tn[13].n82 VGND 0.03989f
C4918 XThR.Tn[13].t61 VGND 0.01487f
C4919 XThR.Tn[13].t47 VGND 0.01628f
C4920 XThR.Tn[13].n83 VGND 0.0415f
C4921 XThR.Tn[13].n84 VGND 0.02916f
C4922 XThR.Tn[13].n86 VGND 0.09357f
C4923 XThR.Tn[13].n87 VGND 0.08503f
C4924 XThR.Tn[13].n88 VGND 0.33338f
C4925 XThC.XTB3.Y.t1 VGND 0.06296f
C4926 XThC.XTB3.Y.n0 VGND 0.04069f
C4927 XThC.XTB3.Y.n1 VGND 0.05192f
C4928 XThC.XTB3.Y.t2 VGND 0.03159f
C4929 XThC.XTB3.Y.t0 VGND 0.03159f
C4930 XThC.XTB3.Y.n2 VGND 0.06782f
C4931 XThC.XTB3.Y.t10 VGND 0.04914f
C4932 XThC.XTB3.Y.t17 VGND 0.02896f
C4933 XThC.XTB3.Y.n3 VGND 0.05852f
C4934 XThC.XTB3.Y.t14 VGND 0.04914f
C4935 XThC.XTB3.Y.t5 VGND 0.02896f
C4936 XThC.XTB3.Y.n4 VGND 0.03012f
C4937 XThC.XTB3.Y.t15 VGND 0.04914f
C4938 XThC.XTB3.Y.t6 VGND 0.02896f
C4939 XThC.XTB3.Y.n5 VGND 0.06469f
C4940 XThC.XTB3.Y.t3 VGND 0.04914f
C4941 XThC.XTB3.Y.t9 VGND 0.02896f
C4942 XThC.XTB3.Y.n6 VGND 0.06006f
C4943 XThC.XTB3.Y.n7 VGND 0.03654f
C4944 XThC.XTB3.Y.n8 VGND 0.06049f
C4945 XThC.XTB3.Y.n9 VGND 0.0234f
C4946 XThC.XTB3.Y.n10 VGND 0.02857f
C4947 XThC.XTB3.Y.n11 VGND 0.06469f
C4948 XThC.XTB3.Y.n12 VGND 0.03243f
C4949 XThC.XTB3.Y.n13 VGND 0.05514f
C4950 XThC.XTB3.Y.t16 VGND 0.04914f
C4951 XThC.XTB3.Y.t7 VGND 0.02896f
C4952 XThC.XTB3.Y.n14 VGND 0.06624f
C4953 XThC.XTB3.Y.t4 VGND 0.04914f
C4954 XThC.XTB3.Y.t13 VGND 0.02896f
C4955 XThC.XTB3.Y.t12 VGND 0.04914f
C4956 XThC.XTB3.Y.t18 VGND 0.02896f
C4957 XThC.XTB3.Y.t11 VGND 0.04914f
C4958 XThC.XTB3.Y.t8 VGND 0.02896f
C4959 XThC.XTB3.Y.n15 VGND 0.08245f
C4960 XThC.XTB3.Y.n16 VGND 0.08709f
C4961 XThC.XTB3.Y.n17 VGND 0.03356f
C4962 XThC.XTB3.Y.n18 VGND 0.07087f
C4963 XThC.XTB3.Y.n19 VGND 0.03243f
C4964 XThC.XTB3.Y.n20 VGND 0.02691f
C4965 XThC.XTB3.Y.n21 VGND 1.39635f
C4966 XThC.XTB3.Y.n22 VGND 0.14933f
C4967 XThR.Tn[8].t6 VGND 0.01919f
C4968 XThR.Tn[8].t4 VGND 0.01919f
C4969 XThR.Tn[8].n0 VGND 0.05828f
C4970 XThR.Tn[8].t7 VGND 0.01919f
C4971 XThR.Tn[8].t5 VGND 0.01919f
C4972 XThR.Tn[8].n1 VGND 0.04267f
C4973 XThR.Tn[8].n2 VGND 0.19401f
C4974 XThR.Tn[8].t3 VGND 0.01248f
C4975 XThR.Tn[8].t8 VGND 0.01248f
C4976 XThR.Tn[8].n3 VGND 0.03112f
C4977 XThR.Tn[8].t11 VGND 0.01248f
C4978 XThR.Tn[8].t9 VGND 0.01248f
C4979 XThR.Tn[8].n4 VGND 0.02495f
C4980 XThR.Tn[8].n5 VGND 0.05754f
C4981 XThR.Tn[8].t39 VGND 0.015f
C4982 XThR.Tn[8].t33 VGND 0.01643f
C4983 XThR.Tn[8].n6 VGND 0.04011f
C4984 XThR.Tn[8].n7 VGND 0.07706f
C4985 XThR.Tn[8].t59 VGND 0.015f
C4986 XThR.Tn[8].t49 VGND 0.01643f
C4987 XThR.Tn[8].n8 VGND 0.04011f
C4988 XThR.Tn[8].t13 VGND 0.01495f
C4989 XThR.Tn[8].t45 VGND 0.01637f
C4990 XThR.Tn[8].n9 VGND 0.04174f
C4991 XThR.Tn[8].n10 VGND 0.02932f
C4992 XThR.Tn[8].n12 VGND 0.09409f
C4993 XThR.Tn[8].t34 VGND 0.015f
C4994 XThR.Tn[8].t26 VGND 0.01643f
C4995 XThR.Tn[8].n13 VGND 0.04011f
C4996 XThR.Tn[8].t53 VGND 0.01495f
C4997 XThR.Tn[8].t22 VGND 0.01637f
C4998 XThR.Tn[8].n14 VGND 0.04174f
C4999 XThR.Tn[8].n15 VGND 0.02932f
C5000 XThR.Tn[8].n17 VGND 0.09409f
C5001 XThR.Tn[8].t50 VGND 0.015f
C5002 XThR.Tn[8].t43 VGND 0.01643f
C5003 XThR.Tn[8].n18 VGND 0.04011f
C5004 XThR.Tn[8].t65 VGND 0.01495f
C5005 XThR.Tn[8].t40 VGND 0.01637f
C5006 XThR.Tn[8].n19 VGND 0.04174f
C5007 XThR.Tn[8].n20 VGND 0.02932f
C5008 XThR.Tn[8].n22 VGND 0.09409f
C5009 XThR.Tn[8].t12 VGND 0.015f
C5010 XThR.Tn[8].t70 VGND 0.01643f
C5011 XThR.Tn[8].n23 VGND 0.04011f
C5012 XThR.Tn[8].t36 VGND 0.01495f
C5013 XThR.Tn[8].t66 VGND 0.01637f
C5014 XThR.Tn[8].n24 VGND 0.04174f
C5015 XThR.Tn[8].n25 VGND 0.02932f
C5016 XThR.Tn[8].n27 VGND 0.09409f
C5017 XThR.Tn[8].t52 VGND 0.015f
C5018 XThR.Tn[8].t44 VGND 0.01643f
C5019 XThR.Tn[8].n28 VGND 0.04011f
C5020 XThR.Tn[8].t68 VGND 0.01495f
C5021 XThR.Tn[8].t41 VGND 0.01637f
C5022 XThR.Tn[8].n29 VGND 0.04174f
C5023 XThR.Tn[8].n30 VGND 0.02932f
C5024 XThR.Tn[8].n32 VGND 0.09409f
C5025 XThR.Tn[8].t28 VGND 0.015f
C5026 XThR.Tn[8].t61 VGND 0.01643f
C5027 XThR.Tn[8].n33 VGND 0.04011f
C5028 XThR.Tn[8].t47 VGND 0.01495f
C5029 XThR.Tn[8].t58 VGND 0.01637f
C5030 XThR.Tn[8].n34 VGND 0.04174f
C5031 XThR.Tn[8].n35 VGND 0.02932f
C5032 XThR.Tn[8].n37 VGND 0.09409f
C5033 XThR.Tn[8].t60 VGND 0.015f
C5034 XThR.Tn[8].t56 VGND 0.01643f
C5035 XThR.Tn[8].n38 VGND 0.04011f
C5036 XThR.Tn[8].t14 VGND 0.01495f
C5037 XThR.Tn[8].t51 VGND 0.01637f
C5038 XThR.Tn[8].n39 VGND 0.04174f
C5039 XThR.Tn[8].n40 VGND 0.02932f
C5040 XThR.Tn[8].n42 VGND 0.09409f
C5041 XThR.Tn[8].t63 VGND 0.015f
C5042 XThR.Tn[8].t69 VGND 0.01643f
C5043 XThR.Tn[8].n43 VGND 0.04011f
C5044 XThR.Tn[8].t20 VGND 0.01495f
C5045 XThR.Tn[8].t64 VGND 0.01637f
C5046 XThR.Tn[8].n44 VGND 0.04174f
C5047 XThR.Tn[8].n45 VGND 0.02932f
C5048 XThR.Tn[8].n47 VGND 0.09409f
C5049 XThR.Tn[8].t17 VGND 0.015f
C5050 XThR.Tn[8].t27 VGND 0.01643f
C5051 XThR.Tn[8].n48 VGND 0.04011f
C5052 XThR.Tn[8].t38 VGND 0.01495f
C5053 XThR.Tn[8].t24 VGND 0.01637f
C5054 XThR.Tn[8].n49 VGND 0.04174f
C5055 XThR.Tn[8].n50 VGND 0.02932f
C5056 XThR.Tn[8].n52 VGND 0.09409f
C5057 XThR.Tn[8].t72 VGND 0.015f
C5058 XThR.Tn[8].t46 VGND 0.01643f
C5059 XThR.Tn[8].n53 VGND 0.04011f
C5060 XThR.Tn[8].t31 VGND 0.01495f
C5061 XThR.Tn[8].t42 VGND 0.01637f
C5062 XThR.Tn[8].n54 VGND 0.04174f
C5063 XThR.Tn[8].n55 VGND 0.02932f
C5064 XThR.Tn[8].n57 VGND 0.09409f
C5065 XThR.Tn[8].t30 VGND 0.015f
C5066 XThR.Tn[8].t21 VGND 0.01643f
C5067 XThR.Tn[8].n58 VGND 0.04011f
C5068 XThR.Tn[8].t48 VGND 0.01495f
C5069 XThR.Tn[8].t16 VGND 0.01637f
C5070 XThR.Tn[8].n59 VGND 0.04174f
C5071 XThR.Tn[8].n60 VGND 0.02932f
C5072 XThR.Tn[8].n62 VGND 0.09409f
C5073 XThR.Tn[8].t62 VGND 0.015f
C5074 XThR.Tn[8].t57 VGND 0.01643f
C5075 XThR.Tn[8].n63 VGND 0.04011f
C5076 XThR.Tn[8].t18 VGND 0.01495f
C5077 XThR.Tn[8].t54 VGND 0.01637f
C5078 XThR.Tn[8].n64 VGND 0.04174f
C5079 XThR.Tn[8].n65 VGND 0.02932f
C5080 XThR.Tn[8].n67 VGND 0.09409f
C5081 XThR.Tn[8].t15 VGND 0.015f
C5082 XThR.Tn[8].t71 VGND 0.01643f
C5083 XThR.Tn[8].n68 VGND 0.04011f
C5084 XThR.Tn[8].t37 VGND 0.01495f
C5085 XThR.Tn[8].t67 VGND 0.01637f
C5086 XThR.Tn[8].n69 VGND 0.04174f
C5087 XThR.Tn[8].n70 VGND 0.02932f
C5088 XThR.Tn[8].n72 VGND 0.09409f
C5089 XThR.Tn[8].t35 VGND 0.015f
C5090 XThR.Tn[8].t29 VGND 0.01643f
C5091 XThR.Tn[8].n73 VGND 0.04011f
C5092 XThR.Tn[8].t55 VGND 0.01495f
C5093 XThR.Tn[8].t25 VGND 0.01637f
C5094 XThR.Tn[8].n74 VGND 0.04174f
C5095 XThR.Tn[8].n75 VGND 0.02932f
C5096 XThR.Tn[8].n77 VGND 0.09409f
C5097 XThR.Tn[8].t73 VGND 0.015f
C5098 XThR.Tn[8].t23 VGND 0.01643f
C5099 XThR.Tn[8].n78 VGND 0.04011f
C5100 XThR.Tn[8].t32 VGND 0.01495f
C5101 XThR.Tn[8].t19 VGND 0.01637f
C5102 XThR.Tn[8].n79 VGND 0.04174f
C5103 XThR.Tn[8].n80 VGND 0.02932f
C5104 XThR.Tn[8].n82 VGND 0.09409f
C5105 XThR.Tn[8].n83 VGND 0.08551f
C5106 XThR.Tn[8].n84 VGND 0.26201f
C5107 XThR.Tn[8].t0 VGND 0.01919f
C5108 XThR.Tn[8].t2 VGND 0.01919f
C5109 XThR.Tn[8].n85 VGND 0.04147f
C5110 XThR.Tn[8].t10 VGND 0.01919f
C5111 XThR.Tn[8].t1 VGND 0.01919f
C5112 XThR.Tn[8].n86 VGND 0.06312f
C5113 XThR.Tn[8].n87 VGND 0.17526f
C5114 XThR.Tn[0].t3 VGND 0.01769f
C5115 XThR.Tn[0].t4 VGND 0.01769f
C5116 XThR.Tn[0].n0 VGND 0.03571f
C5117 XThR.Tn[0].t2 VGND 0.01769f
C5118 XThR.Tn[0].t1 VGND 0.01769f
C5119 XThR.Tn[0].n1 VGND 0.04178f
C5120 XThR.Tn[0].n2 VGND 0.12532f
C5121 XThR.Tn[0].t6 VGND 0.0115f
C5122 XThR.Tn[0].t7 VGND 0.0115f
C5123 XThR.Tn[0].n3 VGND 0.02618f
C5124 XThR.Tn[0].t5 VGND 0.0115f
C5125 XThR.Tn[0].t8 VGND 0.0115f
C5126 XThR.Tn[0].n4 VGND 0.02618f
C5127 XThR.Tn[0].t11 VGND 0.0115f
C5128 XThR.Tn[0].t9 VGND 0.0115f
C5129 XThR.Tn[0].n5 VGND 0.02618f
C5130 XThR.Tn[0].t0 VGND 0.0115f
C5131 XThR.Tn[0].t10 VGND 0.0115f
C5132 XThR.Tn[0].n6 VGND 0.04363f
C5133 XThR.Tn[0].n7 VGND 0.12469f
C5134 XThR.Tn[0].n8 VGND 0.07708f
C5135 XThR.Tn[0].n9 VGND 0.08699f
C5136 XThR.Tn[0].t48 VGND 0.01383f
C5137 XThR.Tn[0].t40 VGND 0.01514f
C5138 XThR.Tn[0].n10 VGND 0.03697f
C5139 XThR.Tn[0].n11 VGND 0.07101f
C5140 XThR.Tn[0].t67 VGND 0.01383f
C5141 XThR.Tn[0].t58 VGND 0.01514f
C5142 XThR.Tn[0].n12 VGND 0.03697f
C5143 XThR.Tn[0].t24 VGND 0.01378f
C5144 XThR.Tn[0].t50 VGND 0.01509f
C5145 XThR.Tn[0].n13 VGND 0.03846f
C5146 XThR.Tn[0].n14 VGND 0.02702f
C5147 XThR.Tn[0].n16 VGND 0.08671f
C5148 XThR.Tn[0].t41 VGND 0.01383f
C5149 XThR.Tn[0].t33 VGND 0.01514f
C5150 XThR.Tn[0].n17 VGND 0.03697f
C5151 XThR.Tn[0].t61 VGND 0.01378f
C5152 XThR.Tn[0].t26 VGND 0.01509f
C5153 XThR.Tn[0].n18 VGND 0.03846f
C5154 XThR.Tn[0].n19 VGND 0.02702f
C5155 XThR.Tn[0].n21 VGND 0.08671f
C5156 XThR.Tn[0].t59 VGND 0.01383f
C5157 XThR.Tn[0].t51 VGND 0.01514f
C5158 XThR.Tn[0].n22 VGND 0.03697f
C5159 XThR.Tn[0].t12 VGND 0.01378f
C5160 XThR.Tn[0].t44 VGND 0.01509f
C5161 XThR.Tn[0].n23 VGND 0.03846f
C5162 XThR.Tn[0].n24 VGND 0.02702f
C5163 XThR.Tn[0].n26 VGND 0.08671f
C5164 XThR.Tn[0].t21 VGND 0.01383f
C5165 XThR.Tn[0].t15 VGND 0.01514f
C5166 XThR.Tn[0].n27 VGND 0.03697f
C5167 XThR.Tn[0].t43 VGND 0.01378f
C5168 XThR.Tn[0].t72 VGND 0.01509f
C5169 XThR.Tn[0].n28 VGND 0.03846f
C5170 XThR.Tn[0].n29 VGND 0.02702f
C5171 XThR.Tn[0].n31 VGND 0.08671f
C5172 XThR.Tn[0].t60 VGND 0.01383f
C5173 XThR.Tn[0].t52 VGND 0.01514f
C5174 XThR.Tn[0].n32 VGND 0.03697f
C5175 XThR.Tn[0].t13 VGND 0.01378f
C5176 XThR.Tn[0].t46 VGND 0.01509f
C5177 XThR.Tn[0].n33 VGND 0.03846f
C5178 XThR.Tn[0].n34 VGND 0.02702f
C5179 XThR.Tn[0].n36 VGND 0.08671f
C5180 XThR.Tn[0].t35 VGND 0.01383f
C5181 XThR.Tn[0].t68 VGND 0.01514f
C5182 XThR.Tn[0].n37 VGND 0.03697f
C5183 XThR.Tn[0].t54 VGND 0.01378f
C5184 XThR.Tn[0].t64 VGND 0.01509f
C5185 XThR.Tn[0].n38 VGND 0.03846f
C5186 XThR.Tn[0].n39 VGND 0.02702f
C5187 XThR.Tn[0].n41 VGND 0.08671f
C5188 XThR.Tn[0].t66 VGND 0.01383f
C5189 XThR.Tn[0].t63 VGND 0.01514f
C5190 XThR.Tn[0].n42 VGND 0.03697f
C5191 XThR.Tn[0].t23 VGND 0.01378f
C5192 XThR.Tn[0].t55 VGND 0.01509f
C5193 XThR.Tn[0].n43 VGND 0.03846f
C5194 XThR.Tn[0].n44 VGND 0.02702f
C5195 XThR.Tn[0].n46 VGND 0.08671f
C5196 XThR.Tn[0].t70 VGND 0.01383f
C5197 XThR.Tn[0].t14 VGND 0.01514f
C5198 XThR.Tn[0].n47 VGND 0.03697f
C5199 XThR.Tn[0].t28 VGND 0.01378f
C5200 XThR.Tn[0].t71 VGND 0.01509f
C5201 XThR.Tn[0].n48 VGND 0.03846f
C5202 XThR.Tn[0].n49 VGND 0.02702f
C5203 XThR.Tn[0].n51 VGND 0.08671f
C5204 XThR.Tn[0].t25 VGND 0.01383f
C5205 XThR.Tn[0].t34 VGND 0.01514f
C5206 XThR.Tn[0].n52 VGND 0.03697f
C5207 XThR.Tn[0].t47 VGND 0.01378f
C5208 XThR.Tn[0].t29 VGND 0.01509f
C5209 XThR.Tn[0].n53 VGND 0.03846f
C5210 XThR.Tn[0].n54 VGND 0.02702f
C5211 XThR.Tn[0].n56 VGND 0.08671f
C5212 XThR.Tn[0].t17 VGND 0.01383f
C5213 XThR.Tn[0].t53 VGND 0.01514f
C5214 XThR.Tn[0].n57 VGND 0.03697f
C5215 XThR.Tn[0].t38 VGND 0.01378f
C5216 XThR.Tn[0].t49 VGND 0.01509f
C5217 XThR.Tn[0].n58 VGND 0.03846f
C5218 XThR.Tn[0].n59 VGND 0.02702f
C5219 XThR.Tn[0].n61 VGND 0.08671f
C5220 XThR.Tn[0].t37 VGND 0.01383f
C5221 XThR.Tn[0].t31 VGND 0.01514f
C5222 XThR.Tn[0].n62 VGND 0.03697f
C5223 XThR.Tn[0].t56 VGND 0.01378f
C5224 XThR.Tn[0].t19 VGND 0.01509f
C5225 XThR.Tn[0].n63 VGND 0.03846f
C5226 XThR.Tn[0].n64 VGND 0.02702f
C5227 XThR.Tn[0].n66 VGND 0.08671f
C5228 XThR.Tn[0].t69 VGND 0.01383f
C5229 XThR.Tn[0].t65 VGND 0.01514f
C5230 XThR.Tn[0].n67 VGND 0.03697f
C5231 XThR.Tn[0].t27 VGND 0.01378f
C5232 XThR.Tn[0].t57 VGND 0.01509f
C5233 XThR.Tn[0].n68 VGND 0.03846f
C5234 XThR.Tn[0].n69 VGND 0.02702f
C5235 XThR.Tn[0].n71 VGND 0.08671f
C5236 XThR.Tn[0].t22 VGND 0.01383f
C5237 XThR.Tn[0].t16 VGND 0.01514f
C5238 XThR.Tn[0].n72 VGND 0.03697f
C5239 XThR.Tn[0].t45 VGND 0.01378f
C5240 XThR.Tn[0].t73 VGND 0.01509f
C5241 XThR.Tn[0].n73 VGND 0.03846f
C5242 XThR.Tn[0].n74 VGND 0.02702f
C5243 XThR.Tn[0].n76 VGND 0.08671f
C5244 XThR.Tn[0].t42 VGND 0.01383f
C5245 XThR.Tn[0].t36 VGND 0.01514f
C5246 XThR.Tn[0].n77 VGND 0.03697f
C5247 XThR.Tn[0].t62 VGND 0.01378f
C5248 XThR.Tn[0].t30 VGND 0.01509f
C5249 XThR.Tn[0].n78 VGND 0.03846f
C5250 XThR.Tn[0].n79 VGND 0.02702f
C5251 XThR.Tn[0].n81 VGND 0.08671f
C5252 XThR.Tn[0].t18 VGND 0.01383f
C5253 XThR.Tn[0].t32 VGND 0.01514f
C5254 XThR.Tn[0].n82 VGND 0.03697f
C5255 XThR.Tn[0].t39 VGND 0.01378f
C5256 XThR.Tn[0].t20 VGND 0.01509f
C5257 XThR.Tn[0].n83 VGND 0.03846f
C5258 XThR.Tn[0].n84 VGND 0.02702f
C5259 XThR.Tn[0].n86 VGND 0.08671f
C5260 XThR.Tn[0].n87 VGND 0.0788f
C5261 XThR.Tn[0].n88 VGND 0.22563f
C5262 XThR.Tn[7].t2 VGND 0.0118f
C5263 XThR.Tn[7].t1 VGND 0.0118f
C5264 XThR.Tn[7].n0 VGND 0.02606f
C5265 XThR.Tn[7].t3 VGND 0.0118f
C5266 XThR.Tn[7].t0 VGND 0.0118f
C5267 XThR.Tn[7].n1 VGND 0.03641f
C5268 XThR.Tn[7].n2 VGND 0.13363f
C5269 XThR.Tn[7].t6 VGND 0.01815f
C5270 XThR.Tn[7].t7 VGND 0.01815f
C5271 XThR.Tn[7].n3 VGND 0.05527f
C5272 XThR.Tn[7].t5 VGND 0.01815f
C5273 XThR.Tn[7].t4 VGND 0.01815f
C5274 XThR.Tn[7].n4 VGND 0.04021f
C5275 XThR.Tn[7].n5 VGND 0.17693f
C5276 XThR.Tn[7].n6 VGND 0.02205f
C5277 XThR.Tn[7].t53 VGND 0.01419f
C5278 XThR.Tn[7].t45 VGND 0.01553f
C5279 XThR.Tn[7].n7 VGND 0.03793f
C5280 XThR.Tn[7].n8 VGND 0.07287f
C5281 XThR.Tn[7].t8 VGND 0.01419f
C5282 XThR.Tn[7].t60 VGND 0.01553f
C5283 XThR.Tn[7].n9 VGND 0.03793f
C5284 XThR.Tn[7].t26 VGND 0.01414f
C5285 XThR.Tn[7].t38 VGND 0.01548f
C5286 XThR.Tn[7].n10 VGND 0.03947f
C5287 XThR.Tn[7].n11 VGND 0.02773f
C5288 XThR.Tn[7].n13 VGND 0.08897f
C5289 XThR.Tn[7].t47 VGND 0.01419f
C5290 XThR.Tn[7].t37 VGND 0.01553f
C5291 XThR.Tn[7].n14 VGND 0.03793f
C5292 XThR.Tn[7].t66 VGND 0.01414f
C5293 XThR.Tn[7].t15 VGND 0.01548f
C5294 XThR.Tn[7].n15 VGND 0.03947f
C5295 XThR.Tn[7].n16 VGND 0.02773f
C5296 XThR.Tn[7].n18 VGND 0.08897f
C5297 XThR.Tn[7].t62 VGND 0.01419f
C5298 XThR.Tn[7].t55 VGND 0.01553f
C5299 XThR.Tn[7].n19 VGND 0.03793f
C5300 XThR.Tn[7].t18 VGND 0.01414f
C5301 XThR.Tn[7].t32 VGND 0.01548f
C5302 XThR.Tn[7].n20 VGND 0.03947f
C5303 XThR.Tn[7].n21 VGND 0.02773f
C5304 XThR.Tn[7].n23 VGND 0.08897f
C5305 XThR.Tn[7].t25 VGND 0.01419f
C5306 XThR.Tn[7].t21 VGND 0.01553f
C5307 XThR.Tn[7].n24 VGND 0.03793f
C5308 XThR.Tn[7].t50 VGND 0.01414f
C5309 XThR.Tn[7].t63 VGND 0.01548f
C5310 XThR.Tn[7].n25 VGND 0.03947f
C5311 XThR.Tn[7].n26 VGND 0.02773f
C5312 XThR.Tn[7].n28 VGND 0.08897f
C5313 XThR.Tn[7].t65 VGND 0.01419f
C5314 XThR.Tn[7].t56 VGND 0.01553f
C5315 XThR.Tn[7].n29 VGND 0.03793f
C5316 XThR.Tn[7].t19 VGND 0.01414f
C5317 XThR.Tn[7].t34 VGND 0.01548f
C5318 XThR.Tn[7].n30 VGND 0.03947f
C5319 XThR.Tn[7].n31 VGND 0.02773f
C5320 XThR.Tn[7].n33 VGND 0.08897f
C5321 XThR.Tn[7].t40 VGND 0.01419f
C5322 XThR.Tn[7].t11 VGND 0.01553f
C5323 XThR.Tn[7].n34 VGND 0.03793f
C5324 XThR.Tn[7].t58 VGND 0.01414f
C5325 XThR.Tn[7].t54 VGND 0.01548f
C5326 XThR.Tn[7].n35 VGND 0.03947f
C5327 XThR.Tn[7].n36 VGND 0.02773f
C5328 XThR.Tn[7].n38 VGND 0.08897f
C5329 XThR.Tn[7].t9 VGND 0.01419f
C5330 XThR.Tn[7].t68 VGND 0.01553f
C5331 XThR.Tn[7].n39 VGND 0.03793f
C5332 XThR.Tn[7].t27 VGND 0.01414f
C5333 XThR.Tn[7].t46 VGND 0.01548f
C5334 XThR.Tn[7].n40 VGND 0.03947f
C5335 XThR.Tn[7].n41 VGND 0.02773f
C5336 XThR.Tn[7].n43 VGND 0.08897f
C5337 XThR.Tn[7].t14 VGND 0.01419f
C5338 XThR.Tn[7].t20 VGND 0.01553f
C5339 XThR.Tn[7].n44 VGND 0.03793f
C5340 XThR.Tn[7].t31 VGND 0.01414f
C5341 XThR.Tn[7].t61 VGND 0.01548f
C5342 XThR.Tn[7].n45 VGND 0.03947f
C5343 XThR.Tn[7].n46 VGND 0.02773f
C5344 XThR.Tn[7].n48 VGND 0.08897f
C5345 XThR.Tn[7].t29 VGND 0.01419f
C5346 XThR.Tn[7].t39 VGND 0.01553f
C5347 XThR.Tn[7].n49 VGND 0.03793f
C5348 XThR.Tn[7].t52 VGND 0.01414f
C5349 XThR.Tn[7].t16 VGND 0.01548f
C5350 XThR.Tn[7].n50 VGND 0.03947f
C5351 XThR.Tn[7].n51 VGND 0.02773f
C5352 XThR.Tn[7].n53 VGND 0.08897f
C5353 XThR.Tn[7].t23 VGND 0.01419f
C5354 XThR.Tn[7].t57 VGND 0.01553f
C5355 XThR.Tn[7].n54 VGND 0.03793f
C5356 XThR.Tn[7].t43 VGND 0.01414f
C5357 XThR.Tn[7].t36 VGND 0.01548f
C5358 XThR.Tn[7].n55 VGND 0.03947f
C5359 XThR.Tn[7].n56 VGND 0.02773f
C5360 XThR.Tn[7].n58 VGND 0.08897f
C5361 XThR.Tn[7].t42 VGND 0.01419f
C5362 XThR.Tn[7].t33 VGND 0.01553f
C5363 XThR.Tn[7].n59 VGND 0.03793f
C5364 XThR.Tn[7].t59 VGND 0.01414f
C5365 XThR.Tn[7].t10 VGND 0.01548f
C5366 XThR.Tn[7].n60 VGND 0.03947f
C5367 XThR.Tn[7].n61 VGND 0.02773f
C5368 XThR.Tn[7].n63 VGND 0.08897f
C5369 XThR.Tn[7].t12 VGND 0.01419f
C5370 XThR.Tn[7].t69 VGND 0.01553f
C5371 XThR.Tn[7].n64 VGND 0.03793f
C5372 XThR.Tn[7].t30 VGND 0.01414f
C5373 XThR.Tn[7].t48 VGND 0.01548f
C5374 XThR.Tn[7].n65 VGND 0.03947f
C5375 XThR.Tn[7].n66 VGND 0.02773f
C5376 XThR.Tn[7].n68 VGND 0.08897f
C5377 XThR.Tn[7].t28 VGND 0.01419f
C5378 XThR.Tn[7].t22 VGND 0.01553f
C5379 XThR.Tn[7].n69 VGND 0.03793f
C5380 XThR.Tn[7].t51 VGND 0.01414f
C5381 XThR.Tn[7].t64 VGND 0.01548f
C5382 XThR.Tn[7].n70 VGND 0.03947f
C5383 XThR.Tn[7].n71 VGND 0.02773f
C5384 XThR.Tn[7].n73 VGND 0.08897f
C5385 XThR.Tn[7].t49 VGND 0.01419f
C5386 XThR.Tn[7].t41 VGND 0.01553f
C5387 XThR.Tn[7].n74 VGND 0.03793f
C5388 XThR.Tn[7].t67 VGND 0.01414f
C5389 XThR.Tn[7].t17 VGND 0.01548f
C5390 XThR.Tn[7].n75 VGND 0.03947f
C5391 XThR.Tn[7].n76 VGND 0.02773f
C5392 XThR.Tn[7].n78 VGND 0.08897f
C5393 XThR.Tn[7].t24 VGND 0.01419f
C5394 XThR.Tn[7].t35 VGND 0.01553f
C5395 XThR.Tn[7].n79 VGND 0.03793f
C5396 XThR.Tn[7].t44 VGND 0.01414f
C5397 XThR.Tn[7].t13 VGND 0.01548f
C5398 XThR.Tn[7].n80 VGND 0.03947f
C5399 XThR.Tn[7].n81 VGND 0.02773f
C5400 XThR.Tn[7].n83 VGND 0.08897f
C5401 XThR.Tn[7].n84 VGND 0.08086f
C5402 XThR.Tn[7].n85 VGND 0.32824f
C5403 XThR.Tn[11].t2 VGND 0.01248f
C5404 XThR.Tn[11].t0 VGND 0.01248f
C5405 XThR.Tn[11].n0 VGND 0.02496f
C5406 XThR.Tn[11].t3 VGND 0.01248f
C5407 XThR.Tn[11].t1 VGND 0.01248f
C5408 XThR.Tn[11].n1 VGND 0.03112f
C5409 XThR.Tn[11].n2 VGND 0.06279f
C5410 XThR.Tn[11].t8 VGND 0.0192f
C5411 XThR.Tn[11].t10 VGND 0.0192f
C5412 XThR.Tn[11].n3 VGND 0.05829f
C5413 XThR.Tn[11].t9 VGND 0.0192f
C5414 XThR.Tn[11].t11 VGND 0.0192f
C5415 XThR.Tn[11].n4 VGND 0.04268f
C5416 XThR.Tn[11].n5 VGND 0.19406f
C5417 XThR.Tn[11].t4 VGND 0.0192f
C5418 XThR.Tn[11].t6 VGND 0.0192f
C5419 XThR.Tn[11].n6 VGND 0.04148f
C5420 XThR.Tn[11].t5 VGND 0.0192f
C5421 XThR.Tn[11].t7 VGND 0.0192f
C5422 XThR.Tn[11].n7 VGND 0.06313f
C5423 XThR.Tn[11].n8 VGND 0.1753f
C5424 XThR.Tn[11].n9 VGND 0.02347f
C5425 XThR.Tn[11].t56 VGND 0.015f
C5426 XThR.Tn[11].t48 VGND 0.01643f
C5427 XThR.Tn[11].n10 VGND 0.04012f
C5428 XThR.Tn[11].n11 VGND 0.07707f
C5429 XThR.Tn[11].t12 VGND 0.015f
C5430 XThR.Tn[11].t67 VGND 0.01643f
C5431 XThR.Tn[11].n12 VGND 0.04012f
C5432 XThR.Tn[11].t27 VGND 0.01496f
C5433 XThR.Tn[11].t58 VGND 0.01638f
C5434 XThR.Tn[11].n13 VGND 0.04174f
C5435 XThR.Tn[11].n14 VGND 0.02933f
C5436 XThR.Tn[11].n16 VGND 0.09411f
C5437 XThR.Tn[11].t49 VGND 0.015f
C5438 XThR.Tn[11].t41 VGND 0.01643f
C5439 XThR.Tn[11].n17 VGND 0.04012f
C5440 XThR.Tn[11].t65 VGND 0.01496f
C5441 XThR.Tn[11].t36 VGND 0.01638f
C5442 XThR.Tn[11].n18 VGND 0.04174f
C5443 XThR.Tn[11].n19 VGND 0.02933f
C5444 XThR.Tn[11].n21 VGND 0.09411f
C5445 XThR.Tn[11].t68 VGND 0.015f
C5446 XThR.Tn[11].t60 VGND 0.01643f
C5447 XThR.Tn[11].n22 VGND 0.04012f
C5448 XThR.Tn[11].t18 VGND 0.01496f
C5449 XThR.Tn[11].t54 VGND 0.01638f
C5450 XThR.Tn[11].n23 VGND 0.04174f
C5451 XThR.Tn[11].n24 VGND 0.02933f
C5452 XThR.Tn[11].n26 VGND 0.09411f
C5453 XThR.Tn[11].t33 VGND 0.015f
C5454 XThR.Tn[11].t23 VGND 0.01643f
C5455 XThR.Tn[11].n27 VGND 0.04012f
C5456 XThR.Tn[11].t50 VGND 0.01496f
C5457 XThR.Tn[11].t19 VGND 0.01638f
C5458 XThR.Tn[11].n28 VGND 0.04174f
C5459 XThR.Tn[11].n29 VGND 0.02933f
C5460 XThR.Tn[11].n31 VGND 0.09411f
C5461 XThR.Tn[11].t70 VGND 0.015f
C5462 XThR.Tn[11].t62 VGND 0.01643f
C5463 XThR.Tn[11].n32 VGND 0.04012f
C5464 XThR.Tn[11].t21 VGND 0.01496f
C5465 XThR.Tn[11].t55 VGND 0.01638f
C5466 XThR.Tn[11].n33 VGND 0.04174f
C5467 XThR.Tn[11].n34 VGND 0.02933f
C5468 XThR.Tn[11].n36 VGND 0.09411f
C5469 XThR.Tn[11].t44 VGND 0.015f
C5470 XThR.Tn[11].t14 VGND 0.01643f
C5471 XThR.Tn[11].n37 VGND 0.04012f
C5472 XThR.Tn[11].t59 VGND 0.01496f
C5473 XThR.Tn[11].t72 VGND 0.01638f
C5474 XThR.Tn[11].n38 VGND 0.04174f
C5475 XThR.Tn[11].n39 VGND 0.02933f
C5476 XThR.Tn[11].n41 VGND 0.09411f
C5477 XThR.Tn[11].t13 VGND 0.015f
C5478 XThR.Tn[11].t71 VGND 0.01643f
C5479 XThR.Tn[11].n42 VGND 0.04012f
C5480 XThR.Tn[11].t28 VGND 0.01496f
C5481 XThR.Tn[11].t64 VGND 0.01638f
C5482 XThR.Tn[11].n43 VGND 0.04174f
C5483 XThR.Tn[11].n44 VGND 0.02933f
C5484 XThR.Tn[11].n46 VGND 0.09411f
C5485 XThR.Tn[11].t16 VGND 0.015f
C5486 XThR.Tn[11].t22 VGND 0.01643f
C5487 XThR.Tn[11].n47 VGND 0.04012f
C5488 XThR.Tn[11].t32 VGND 0.01496f
C5489 XThR.Tn[11].t17 VGND 0.01638f
C5490 XThR.Tn[11].n48 VGND 0.04174f
C5491 XThR.Tn[11].n49 VGND 0.02933f
C5492 XThR.Tn[11].n51 VGND 0.09411f
C5493 XThR.Tn[11].t35 VGND 0.015f
C5494 XThR.Tn[11].t43 VGND 0.01643f
C5495 XThR.Tn[11].n52 VGND 0.04012f
C5496 XThR.Tn[11].t52 VGND 0.01496f
C5497 XThR.Tn[11].t37 VGND 0.01638f
C5498 XThR.Tn[11].n53 VGND 0.04174f
C5499 XThR.Tn[11].n54 VGND 0.02933f
C5500 XThR.Tn[11].n56 VGND 0.09411f
C5501 XThR.Tn[11].t25 VGND 0.015f
C5502 XThR.Tn[11].t63 VGND 0.01643f
C5503 XThR.Tn[11].n57 VGND 0.04012f
C5504 XThR.Tn[11].t42 VGND 0.01496f
C5505 XThR.Tn[11].t57 VGND 0.01638f
C5506 XThR.Tn[11].n58 VGND 0.04174f
C5507 XThR.Tn[11].n59 VGND 0.02933f
C5508 XThR.Tn[11].n61 VGND 0.09411f
C5509 XThR.Tn[11].t47 VGND 0.015f
C5510 XThR.Tn[11].t39 VGND 0.01643f
C5511 XThR.Tn[11].n62 VGND 0.04012f
C5512 XThR.Tn[11].t61 VGND 0.01496f
C5513 XThR.Tn[11].t29 VGND 0.01638f
C5514 XThR.Tn[11].n63 VGND 0.04174f
C5515 XThR.Tn[11].n64 VGND 0.02933f
C5516 XThR.Tn[11].n66 VGND 0.09411f
C5517 XThR.Tn[11].t15 VGND 0.015f
C5518 XThR.Tn[11].t73 VGND 0.01643f
C5519 XThR.Tn[11].n67 VGND 0.04012f
C5520 XThR.Tn[11].t30 VGND 0.01496f
C5521 XThR.Tn[11].t66 VGND 0.01638f
C5522 XThR.Tn[11].n68 VGND 0.04174f
C5523 XThR.Tn[11].n69 VGND 0.02933f
C5524 XThR.Tn[11].n71 VGND 0.09411f
C5525 XThR.Tn[11].t34 VGND 0.015f
C5526 XThR.Tn[11].t24 VGND 0.01643f
C5527 XThR.Tn[11].n72 VGND 0.04012f
C5528 XThR.Tn[11].t51 VGND 0.01496f
C5529 XThR.Tn[11].t20 VGND 0.01638f
C5530 XThR.Tn[11].n73 VGND 0.04174f
C5531 XThR.Tn[11].n74 VGND 0.02933f
C5532 XThR.Tn[11].n76 VGND 0.09411f
C5533 XThR.Tn[11].t53 VGND 0.015f
C5534 XThR.Tn[11].t46 VGND 0.01643f
C5535 XThR.Tn[11].n77 VGND 0.04012f
C5536 XThR.Tn[11].t69 VGND 0.01496f
C5537 XThR.Tn[11].t38 VGND 0.01638f
C5538 XThR.Tn[11].n78 VGND 0.04174f
C5539 XThR.Tn[11].n79 VGND 0.02933f
C5540 XThR.Tn[11].n81 VGND 0.09411f
C5541 XThR.Tn[11].t26 VGND 0.015f
C5542 XThR.Tn[11].t40 VGND 0.01643f
C5543 XThR.Tn[11].n82 VGND 0.04012f
C5544 XThR.Tn[11].t45 VGND 0.01496f
C5545 XThR.Tn[11].t31 VGND 0.01638f
C5546 XThR.Tn[11].n83 VGND 0.04174f
C5547 XThR.Tn[11].n84 VGND 0.02933f
C5548 XThR.Tn[11].n86 VGND 0.09411f
C5549 XThR.Tn[11].n87 VGND 0.08553f
C5550 XThR.Tn[11].n88 VGND 0.30653f
C5551 XThR.Tn[4].t1 VGND 0.01806f
C5552 XThR.Tn[4].t2 VGND 0.01806f
C5553 XThR.Tn[4].n0 VGND 0.03645f
C5554 XThR.Tn[4].t0 VGND 0.01806f
C5555 XThR.Tn[4].t3 VGND 0.01806f
C5556 XThR.Tn[4].n1 VGND 0.04265f
C5557 XThR.Tn[4].n2 VGND 0.12794f
C5558 XThR.Tn[4].t8 VGND 0.01174f
C5559 XThR.Tn[4].t9 VGND 0.01174f
C5560 XThR.Tn[4].n3 VGND 0.04454f
C5561 XThR.Tn[4].t11 VGND 0.01174f
C5562 XThR.Tn[4].t10 VGND 0.01174f
C5563 XThR.Tn[4].n4 VGND 0.02673f
C5564 XThR.Tn[4].n5 VGND 0.1273f
C5565 XThR.Tn[4].t6 VGND 0.01174f
C5566 XThR.Tn[4].t5 VGND 0.01174f
C5567 XThR.Tn[4].n6 VGND 0.02673f
C5568 XThR.Tn[4].n7 VGND 0.0787f
C5569 XThR.Tn[4].t7 VGND 0.01174f
C5570 XThR.Tn[4].t4 VGND 0.01174f
C5571 XThR.Tn[4].n8 VGND 0.02673f
C5572 XThR.Tn[4].n9 VGND 0.08881f
C5573 XThR.Tn[4].t44 VGND 0.01411f
C5574 XThR.Tn[4].t38 VGND 0.01545f
C5575 XThR.Tn[4].n10 VGND 0.03774f
C5576 XThR.Tn[4].n11 VGND 0.0725f
C5577 XThR.Tn[4].t65 VGND 0.01411f
C5578 XThR.Tn[4].t54 VGND 0.01545f
C5579 XThR.Tn[4].n12 VGND 0.03774f
C5580 XThR.Tn[4].t19 VGND 0.01407f
C5581 XThR.Tn[4].t50 VGND 0.01541f
C5582 XThR.Tn[4].n13 VGND 0.03927f
C5583 XThR.Tn[4].n14 VGND 0.02759f
C5584 XThR.Tn[4].n16 VGND 0.08853f
C5585 XThR.Tn[4].t39 VGND 0.01411f
C5586 XThR.Tn[4].t31 VGND 0.01545f
C5587 XThR.Tn[4].n17 VGND 0.03774f
C5588 XThR.Tn[4].t58 VGND 0.01407f
C5589 XThR.Tn[4].t27 VGND 0.01541f
C5590 XThR.Tn[4].n18 VGND 0.03927f
C5591 XThR.Tn[4].n19 VGND 0.02759f
C5592 XThR.Tn[4].n21 VGND 0.08853f
C5593 XThR.Tn[4].t55 VGND 0.01411f
C5594 XThR.Tn[4].t48 VGND 0.01545f
C5595 XThR.Tn[4].n22 VGND 0.03774f
C5596 XThR.Tn[4].t70 VGND 0.01407f
C5597 XThR.Tn[4].t45 VGND 0.01541f
C5598 XThR.Tn[4].n23 VGND 0.03927f
C5599 XThR.Tn[4].n24 VGND 0.02759f
C5600 XThR.Tn[4].n26 VGND 0.08853f
C5601 XThR.Tn[4].t17 VGND 0.01411f
C5602 XThR.Tn[4].t13 VGND 0.01545f
C5603 XThR.Tn[4].n27 VGND 0.03774f
C5604 XThR.Tn[4].t41 VGND 0.01407f
C5605 XThR.Tn[4].t71 VGND 0.01541f
C5606 XThR.Tn[4].n28 VGND 0.03927f
C5607 XThR.Tn[4].n29 VGND 0.02759f
C5608 XThR.Tn[4].n31 VGND 0.08853f
C5609 XThR.Tn[4].t57 VGND 0.01411f
C5610 XThR.Tn[4].t49 VGND 0.01545f
C5611 XThR.Tn[4].n32 VGND 0.03774f
C5612 XThR.Tn[4].t73 VGND 0.01407f
C5613 XThR.Tn[4].t46 VGND 0.01541f
C5614 XThR.Tn[4].n33 VGND 0.03927f
C5615 XThR.Tn[4].n34 VGND 0.02759f
C5616 XThR.Tn[4].n36 VGND 0.08853f
C5617 XThR.Tn[4].t33 VGND 0.01411f
C5618 XThR.Tn[4].t66 VGND 0.01545f
C5619 XThR.Tn[4].n37 VGND 0.03774f
C5620 XThR.Tn[4].t52 VGND 0.01407f
C5621 XThR.Tn[4].t63 VGND 0.01541f
C5622 XThR.Tn[4].n38 VGND 0.03927f
C5623 XThR.Tn[4].n39 VGND 0.02759f
C5624 XThR.Tn[4].n41 VGND 0.08853f
C5625 XThR.Tn[4].t64 VGND 0.01411f
C5626 XThR.Tn[4].t61 VGND 0.01545f
C5627 XThR.Tn[4].n42 VGND 0.03774f
C5628 XThR.Tn[4].t18 VGND 0.01407f
C5629 XThR.Tn[4].t56 VGND 0.01541f
C5630 XThR.Tn[4].n43 VGND 0.03927f
C5631 XThR.Tn[4].n44 VGND 0.02759f
C5632 XThR.Tn[4].n46 VGND 0.08853f
C5633 XThR.Tn[4].t68 VGND 0.01411f
C5634 XThR.Tn[4].t12 VGND 0.01545f
C5635 XThR.Tn[4].n47 VGND 0.03774f
C5636 XThR.Tn[4].t25 VGND 0.01407f
C5637 XThR.Tn[4].t69 VGND 0.01541f
C5638 XThR.Tn[4].n48 VGND 0.03927f
C5639 XThR.Tn[4].n49 VGND 0.02759f
C5640 XThR.Tn[4].n51 VGND 0.08853f
C5641 XThR.Tn[4].t22 VGND 0.01411f
C5642 XThR.Tn[4].t32 VGND 0.01545f
C5643 XThR.Tn[4].n52 VGND 0.03774f
C5644 XThR.Tn[4].t43 VGND 0.01407f
C5645 XThR.Tn[4].t29 VGND 0.01541f
C5646 XThR.Tn[4].n53 VGND 0.03927f
C5647 XThR.Tn[4].n54 VGND 0.02759f
C5648 XThR.Tn[4].n56 VGND 0.08853f
C5649 XThR.Tn[4].t15 VGND 0.01411f
C5650 XThR.Tn[4].t51 VGND 0.01545f
C5651 XThR.Tn[4].n57 VGND 0.03774f
C5652 XThR.Tn[4].t36 VGND 0.01407f
C5653 XThR.Tn[4].t47 VGND 0.01541f
C5654 XThR.Tn[4].n58 VGND 0.03927f
C5655 XThR.Tn[4].n59 VGND 0.02759f
C5656 XThR.Tn[4].n61 VGND 0.08853f
C5657 XThR.Tn[4].t35 VGND 0.01411f
C5658 XThR.Tn[4].t26 VGND 0.01545f
C5659 XThR.Tn[4].n62 VGND 0.03774f
C5660 XThR.Tn[4].t53 VGND 0.01407f
C5661 XThR.Tn[4].t21 VGND 0.01541f
C5662 XThR.Tn[4].n63 VGND 0.03927f
C5663 XThR.Tn[4].n64 VGND 0.02759f
C5664 XThR.Tn[4].n66 VGND 0.08853f
C5665 XThR.Tn[4].t67 VGND 0.01411f
C5666 XThR.Tn[4].t62 VGND 0.01545f
C5667 XThR.Tn[4].n67 VGND 0.03774f
C5668 XThR.Tn[4].t23 VGND 0.01407f
C5669 XThR.Tn[4].t59 VGND 0.01541f
C5670 XThR.Tn[4].n68 VGND 0.03927f
C5671 XThR.Tn[4].n69 VGND 0.02759f
C5672 XThR.Tn[4].n71 VGND 0.08853f
C5673 XThR.Tn[4].t20 VGND 0.01411f
C5674 XThR.Tn[4].t14 VGND 0.01545f
C5675 XThR.Tn[4].n72 VGND 0.03774f
C5676 XThR.Tn[4].t42 VGND 0.01407f
C5677 XThR.Tn[4].t72 VGND 0.01541f
C5678 XThR.Tn[4].n73 VGND 0.03927f
C5679 XThR.Tn[4].n74 VGND 0.02759f
C5680 XThR.Tn[4].n76 VGND 0.08853f
C5681 XThR.Tn[4].t40 VGND 0.01411f
C5682 XThR.Tn[4].t34 VGND 0.01545f
C5683 XThR.Tn[4].n77 VGND 0.03774f
C5684 XThR.Tn[4].t60 VGND 0.01407f
C5685 XThR.Tn[4].t30 VGND 0.01541f
C5686 XThR.Tn[4].n78 VGND 0.03927f
C5687 XThR.Tn[4].n79 VGND 0.02759f
C5688 XThR.Tn[4].n81 VGND 0.08853f
C5689 XThR.Tn[4].t16 VGND 0.01411f
C5690 XThR.Tn[4].t28 VGND 0.01545f
C5691 XThR.Tn[4].n82 VGND 0.03774f
C5692 XThR.Tn[4].t37 VGND 0.01407f
C5693 XThR.Tn[4].t24 VGND 0.01541f
C5694 XThR.Tn[4].n83 VGND 0.03927f
C5695 XThR.Tn[4].n84 VGND 0.02759f
C5696 XThR.Tn[4].n86 VGND 0.08853f
C5697 XThR.Tn[4].n87 VGND 0.08045f
C5698 XThR.Tn[4].n88 VGND 0.15199f
C5699 XThC.Tn[7].t4 VGND 0.01305f
C5700 XThC.Tn[7].t7 VGND 0.01305f
C5701 XThC.Tn[7].n0 VGND 0.0281f
C5702 XThC.Tn[7].t6 VGND 0.01305f
C5703 XThC.Tn[7].t5 VGND 0.01305f
C5704 XThC.Tn[7].n1 VGND 0.04266f
C5705 XThC.Tn[7].n2 VGND 0.12542f
C5706 XThC.Tn[7].t8 VGND 0.01034f
C5707 XThC.Tn[7].t11 VGND 0.01129f
C5708 XThC.Tn[7].n3 VGND 0.02522f
C5709 XThC.Tn[7].n4 VGND 0.01441f
C5710 XThC.Tn[7].n5 VGND 0.01753f
C5711 XThC.Tn[7].t25 VGND 0.01034f
C5712 XThC.Tn[7].t30 VGND 0.01129f
C5713 XThC.Tn[7].n6 VGND 0.02522f
C5714 XThC.Tn[7].n7 VGND 0.01441f
C5715 XThC.Tn[7].n8 VGND 0.08328f
C5716 XThC.Tn[7].t27 VGND 0.01034f
C5717 XThC.Tn[7].t34 VGND 0.01129f
C5718 XThC.Tn[7].n9 VGND 0.02522f
C5719 XThC.Tn[7].n10 VGND 0.01441f
C5720 XThC.Tn[7].n11 VGND 0.08328f
C5721 XThC.Tn[7].t29 VGND 0.01034f
C5722 XThC.Tn[7].t35 VGND 0.01129f
C5723 XThC.Tn[7].n12 VGND 0.02522f
C5724 XThC.Tn[7].n13 VGND 0.01441f
C5725 XThC.Tn[7].n14 VGND 0.08328f
C5726 XThC.Tn[7].t18 VGND 0.01034f
C5727 XThC.Tn[7].t22 VGND 0.01129f
C5728 XThC.Tn[7].n15 VGND 0.02522f
C5729 XThC.Tn[7].n16 VGND 0.01441f
C5730 XThC.Tn[7].n17 VGND 0.08328f
C5731 XThC.Tn[7].t20 VGND 0.01034f
C5732 XThC.Tn[7].t23 VGND 0.01129f
C5733 XThC.Tn[7].n18 VGND 0.02522f
C5734 XThC.Tn[7].n19 VGND 0.01441f
C5735 XThC.Tn[7].n20 VGND 0.08328f
C5736 XThC.Tn[7].t33 VGND 0.01034f
C5737 XThC.Tn[7].t39 VGND 0.01129f
C5738 XThC.Tn[7].n21 VGND 0.02522f
C5739 XThC.Tn[7].n22 VGND 0.01441f
C5740 XThC.Tn[7].n23 VGND 0.08328f
C5741 XThC.Tn[7].t10 VGND 0.01034f
C5742 XThC.Tn[7].t14 VGND 0.01129f
C5743 XThC.Tn[7].n24 VGND 0.02522f
C5744 XThC.Tn[7].n25 VGND 0.01441f
C5745 XThC.Tn[7].n26 VGND 0.08328f
C5746 XThC.Tn[7].t12 VGND 0.01034f
C5747 XThC.Tn[7].t16 VGND 0.01129f
C5748 XThC.Tn[7].n27 VGND 0.02522f
C5749 XThC.Tn[7].n28 VGND 0.01441f
C5750 XThC.Tn[7].n29 VGND 0.08328f
C5751 XThC.Tn[7].t31 VGND 0.01034f
C5752 XThC.Tn[7].t36 VGND 0.01129f
C5753 XThC.Tn[7].n30 VGND 0.02522f
C5754 XThC.Tn[7].n31 VGND 0.01441f
C5755 XThC.Tn[7].n32 VGND 0.08328f
C5756 XThC.Tn[7].t32 VGND 0.01034f
C5757 XThC.Tn[7].t38 VGND 0.01129f
C5758 XThC.Tn[7].n33 VGND 0.02522f
C5759 XThC.Tn[7].n34 VGND 0.01441f
C5760 XThC.Tn[7].n35 VGND 0.08328f
C5761 XThC.Tn[7].t13 VGND 0.01034f
C5762 XThC.Tn[7].t17 VGND 0.01129f
C5763 XThC.Tn[7].n36 VGND 0.02522f
C5764 XThC.Tn[7].n37 VGND 0.01441f
C5765 XThC.Tn[7].n38 VGND 0.08328f
C5766 XThC.Tn[7].t21 VGND 0.01034f
C5767 XThC.Tn[7].t26 VGND 0.01129f
C5768 XThC.Tn[7].n39 VGND 0.02522f
C5769 XThC.Tn[7].n40 VGND 0.01441f
C5770 XThC.Tn[7].n41 VGND 0.08328f
C5771 XThC.Tn[7].t24 VGND 0.01034f
C5772 XThC.Tn[7].t28 VGND 0.01129f
C5773 XThC.Tn[7].n42 VGND 0.02522f
C5774 XThC.Tn[7].n43 VGND 0.01441f
C5775 XThC.Tn[7].n44 VGND 0.08328f
C5776 XThC.Tn[7].t37 VGND 0.01034f
C5777 XThC.Tn[7].t9 VGND 0.01129f
C5778 XThC.Tn[7].n45 VGND 0.02522f
C5779 XThC.Tn[7].n46 VGND 0.01441f
C5780 XThC.Tn[7].n47 VGND 0.08328f
C5781 XThC.Tn[7].t15 VGND 0.01034f
C5782 XThC.Tn[7].t19 VGND 0.01129f
C5783 XThC.Tn[7].n48 VGND 0.02522f
C5784 XThC.Tn[7].n49 VGND 0.01441f
C5785 XThC.Tn[7].n50 VGND 0.08328f
C5786 XThC.Tn[7].n51 VGND 0.52699f
C5787 XThC.Tn[7].n52 VGND 0.03388f
C5788 XThC.Tn[7].n53 VGND 0.02617f
C5789 XThC.Tn[7].n54 VGND 0.01873f
C5790 XThC.Tn[7].n55 VGND 0.09263f
C5791 XThC.Tn[7].n56 VGND 0.01561f
C5792 XThR.Tn[1].t11 VGND 0.01166f
C5793 XThR.Tn[1].t8 VGND 0.01166f
C5794 XThR.Tn[1].n0 VGND 0.04425f
C5795 XThR.Tn[1].t10 VGND 0.01166f
C5796 XThR.Tn[1].t9 VGND 0.01166f
C5797 XThR.Tn[1].n1 VGND 0.02656f
C5798 XThR.Tn[1].n2 VGND 0.12648f
C5799 XThR.Tn[1].t6 VGND 0.01166f
C5800 XThR.Tn[1].t5 VGND 0.01166f
C5801 XThR.Tn[1].n3 VGND 0.02656f
C5802 XThR.Tn[1].n4 VGND 0.07819f
C5803 XThR.Tn[1].t7 VGND 0.01166f
C5804 XThR.Tn[1].t4 VGND 0.01166f
C5805 XThR.Tn[1].n5 VGND 0.02656f
C5806 XThR.Tn[1].n6 VGND 0.08824f
C5807 XThR.Tn[1].t24 VGND 0.01402f
C5808 XThR.Tn[1].t18 VGND 0.01536f
C5809 XThR.Tn[1].n7 VGND 0.0375f
C5810 XThR.Tn[1].n8 VGND 0.07203f
C5811 XThR.Tn[1].t44 VGND 0.01402f
C5812 XThR.Tn[1].t34 VGND 0.01536f
C5813 XThR.Tn[1].n9 VGND 0.0375f
C5814 XThR.Tn[1].t61 VGND 0.01398f
C5815 XThR.Tn[1].t30 VGND 0.01531f
C5816 XThR.Tn[1].n10 VGND 0.03901f
C5817 XThR.Tn[1].n11 VGND 0.02741f
C5818 XThR.Tn[1].n13 VGND 0.08795f
C5819 XThR.Tn[1].t19 VGND 0.01402f
C5820 XThR.Tn[1].t73 VGND 0.01536f
C5821 XThR.Tn[1].n14 VGND 0.0375f
C5822 XThR.Tn[1].t38 VGND 0.01398f
C5823 XThR.Tn[1].t69 VGND 0.01531f
C5824 XThR.Tn[1].n15 VGND 0.03901f
C5825 XThR.Tn[1].n16 VGND 0.02741f
C5826 XThR.Tn[1].n18 VGND 0.08795f
C5827 XThR.Tn[1].t35 VGND 0.01402f
C5828 XThR.Tn[1].t28 VGND 0.01536f
C5829 XThR.Tn[1].n19 VGND 0.0375f
C5830 XThR.Tn[1].t50 VGND 0.01398f
C5831 XThR.Tn[1].t25 VGND 0.01531f
C5832 XThR.Tn[1].n20 VGND 0.03901f
C5833 XThR.Tn[1].n21 VGND 0.02741f
C5834 XThR.Tn[1].n23 VGND 0.08795f
C5835 XThR.Tn[1].t59 VGND 0.01402f
C5836 XThR.Tn[1].t55 VGND 0.01536f
C5837 XThR.Tn[1].n24 VGND 0.0375f
C5838 XThR.Tn[1].t21 VGND 0.01398f
C5839 XThR.Tn[1].t51 VGND 0.01531f
C5840 XThR.Tn[1].n25 VGND 0.03901f
C5841 XThR.Tn[1].n26 VGND 0.02741f
C5842 XThR.Tn[1].n28 VGND 0.08795f
C5843 XThR.Tn[1].t37 VGND 0.01402f
C5844 XThR.Tn[1].t29 VGND 0.01536f
C5845 XThR.Tn[1].n29 VGND 0.0375f
C5846 XThR.Tn[1].t53 VGND 0.01398f
C5847 XThR.Tn[1].t26 VGND 0.01531f
C5848 XThR.Tn[1].n30 VGND 0.03901f
C5849 XThR.Tn[1].n31 VGND 0.02741f
C5850 XThR.Tn[1].n33 VGND 0.08795f
C5851 XThR.Tn[1].t13 VGND 0.01402f
C5852 XThR.Tn[1].t46 VGND 0.01536f
C5853 XThR.Tn[1].n34 VGND 0.0375f
C5854 XThR.Tn[1].t32 VGND 0.01398f
C5855 XThR.Tn[1].t43 VGND 0.01531f
C5856 XThR.Tn[1].n35 VGND 0.03901f
C5857 XThR.Tn[1].n36 VGND 0.02741f
C5858 XThR.Tn[1].n38 VGND 0.08795f
C5859 XThR.Tn[1].t45 VGND 0.01402f
C5860 XThR.Tn[1].t41 VGND 0.01536f
C5861 XThR.Tn[1].n39 VGND 0.0375f
C5862 XThR.Tn[1].t60 VGND 0.01398f
C5863 XThR.Tn[1].t36 VGND 0.01531f
C5864 XThR.Tn[1].n40 VGND 0.03901f
C5865 XThR.Tn[1].n41 VGND 0.02741f
C5866 XThR.Tn[1].n43 VGND 0.08795f
C5867 XThR.Tn[1].t48 VGND 0.01402f
C5868 XThR.Tn[1].t54 VGND 0.01536f
C5869 XThR.Tn[1].n44 VGND 0.0375f
C5870 XThR.Tn[1].t67 VGND 0.01398f
C5871 XThR.Tn[1].t49 VGND 0.01531f
C5872 XThR.Tn[1].n45 VGND 0.03901f
C5873 XThR.Tn[1].n46 VGND 0.02741f
C5874 XThR.Tn[1].n48 VGND 0.08795f
C5875 XThR.Tn[1].t64 VGND 0.01402f
C5876 XThR.Tn[1].t12 VGND 0.01536f
C5877 XThR.Tn[1].n49 VGND 0.0375f
C5878 XThR.Tn[1].t23 VGND 0.01398f
C5879 XThR.Tn[1].t71 VGND 0.01531f
C5880 XThR.Tn[1].n50 VGND 0.03901f
C5881 XThR.Tn[1].n51 VGND 0.02741f
C5882 XThR.Tn[1].n53 VGND 0.08795f
C5883 XThR.Tn[1].t57 VGND 0.01402f
C5884 XThR.Tn[1].t31 VGND 0.01536f
C5885 XThR.Tn[1].n54 VGND 0.0375f
C5886 XThR.Tn[1].t16 VGND 0.01398f
C5887 XThR.Tn[1].t27 VGND 0.01531f
C5888 XThR.Tn[1].n55 VGND 0.03901f
C5889 XThR.Tn[1].n56 VGND 0.02741f
C5890 XThR.Tn[1].n58 VGND 0.08795f
C5891 XThR.Tn[1].t15 VGND 0.01402f
C5892 XThR.Tn[1].t68 VGND 0.01536f
C5893 XThR.Tn[1].n59 VGND 0.0375f
C5894 XThR.Tn[1].t33 VGND 0.01398f
C5895 XThR.Tn[1].t63 VGND 0.01531f
C5896 XThR.Tn[1].n60 VGND 0.03901f
C5897 XThR.Tn[1].n61 VGND 0.02741f
C5898 XThR.Tn[1].n63 VGND 0.08795f
C5899 XThR.Tn[1].t47 VGND 0.01402f
C5900 XThR.Tn[1].t42 VGND 0.01536f
C5901 XThR.Tn[1].n64 VGND 0.0375f
C5902 XThR.Tn[1].t65 VGND 0.01398f
C5903 XThR.Tn[1].t39 VGND 0.01531f
C5904 XThR.Tn[1].n65 VGND 0.03901f
C5905 XThR.Tn[1].n66 VGND 0.02741f
C5906 XThR.Tn[1].n68 VGND 0.08795f
C5907 XThR.Tn[1].t62 VGND 0.01402f
C5908 XThR.Tn[1].t56 VGND 0.01536f
C5909 XThR.Tn[1].n69 VGND 0.0375f
C5910 XThR.Tn[1].t22 VGND 0.01398f
C5911 XThR.Tn[1].t52 VGND 0.01531f
C5912 XThR.Tn[1].n70 VGND 0.03901f
C5913 XThR.Tn[1].n71 VGND 0.02741f
C5914 XThR.Tn[1].n73 VGND 0.08795f
C5915 XThR.Tn[1].t20 VGND 0.01402f
C5916 XThR.Tn[1].t14 VGND 0.01536f
C5917 XThR.Tn[1].n74 VGND 0.0375f
C5918 XThR.Tn[1].t40 VGND 0.01398f
C5919 XThR.Tn[1].t72 VGND 0.01531f
C5920 XThR.Tn[1].n75 VGND 0.03901f
C5921 XThR.Tn[1].n76 VGND 0.02741f
C5922 XThR.Tn[1].n78 VGND 0.08795f
C5923 XThR.Tn[1].t58 VGND 0.01402f
C5924 XThR.Tn[1].t70 VGND 0.01536f
C5925 XThR.Tn[1].n79 VGND 0.0375f
C5926 XThR.Tn[1].t17 VGND 0.01398f
C5927 XThR.Tn[1].t66 VGND 0.01531f
C5928 XThR.Tn[1].n80 VGND 0.03901f
C5929 XThR.Tn[1].n81 VGND 0.02741f
C5930 XThR.Tn[1].n83 VGND 0.08795f
C5931 XThR.Tn[1].n84 VGND 0.07993f
C5932 XThR.Tn[1].n85 VGND 0.23008f
C5933 XThR.Tn[1].t0 VGND 0.01794f
C5934 XThR.Tn[1].t1 VGND 0.01794f
C5935 XThR.Tn[1].n86 VGND 0.03622f
C5936 XThR.Tn[1].t3 VGND 0.01794f
C5937 XThR.Tn[1].t2 VGND 0.01794f
C5938 XThR.Tn[1].n87 VGND 0.04238f
C5939 XThR.Tn[1].n88 VGND 0.11863f
C5940 XThR.Tn[1].n89 VGND 0.03755f
C5941 XThC.Tn[8].n0 VGND 0.02379f
C5942 XThC.Tn[8].n1 VGND 0.01907f
C5943 XThC.Tn[8].n2 VGND 0.04799f
C5944 XThC.Tn[8].t5 VGND 0.01467f
C5945 XThC.Tn[8].t6 VGND 0.01467f
C5946 XThC.Tn[8].n3 VGND 0.0317f
C5947 XThC.Tn[8].t4 VGND 0.01467f
C5948 XThC.Tn[8].t7 VGND 0.01467f
C5949 XThC.Tn[8].n4 VGND 0.04825f
C5950 XThC.Tn[8].n5 VGND 0.13407f
C5951 XThC.Tn[8].t8 VGND 0.01467f
C5952 XThC.Tn[8].t11 VGND 0.01467f
C5953 XThC.Tn[8].n6 VGND 0.04455f
C5954 XThC.Tn[8].t10 VGND 0.01467f
C5955 XThC.Tn[8].t9 VGND 0.01467f
C5956 XThC.Tn[8].n7 VGND 0.03262f
C5957 XThC.Tn[8].n8 VGND 0.14517f
C5958 XThC.Tn[8].n9 VGND 0.02108f
C5959 XThC.Tn[8].t43 VGND 0.01163f
C5960 XThC.Tn[8].t41 VGND 0.0127f
C5961 XThC.Tn[8].n10 VGND 0.02837f
C5962 XThC.Tn[8].n11 VGND 0.01621f
C5963 XThC.Tn[8].n12 VGND 0.01972f
C5964 XThC.Tn[8].t29 VGND 0.01163f
C5965 XThC.Tn[8].t26 VGND 0.0127f
C5966 XThC.Tn[8].n13 VGND 0.02837f
C5967 XThC.Tn[8].n14 VGND 0.01621f
C5968 XThC.Tn[8].n15 VGND 0.09367f
C5969 XThC.Tn[8].t34 VGND 0.01163f
C5970 XThC.Tn[8].t28 VGND 0.0127f
C5971 XThC.Tn[8].n16 VGND 0.02837f
C5972 XThC.Tn[8].n17 VGND 0.01621f
C5973 XThC.Tn[8].n18 VGND 0.09367f
C5974 XThC.Tn[8].t35 VGND 0.01163f
C5975 XThC.Tn[8].t30 VGND 0.0127f
C5976 XThC.Tn[8].n19 VGND 0.02837f
C5977 XThC.Tn[8].n20 VGND 0.01621f
C5978 XThC.Tn[8].n21 VGND 0.09367f
C5979 XThC.Tn[8].t22 VGND 0.01163f
C5980 XThC.Tn[8].t19 VGND 0.0127f
C5981 XThC.Tn[8].n22 VGND 0.02837f
C5982 XThC.Tn[8].n23 VGND 0.01621f
C5983 XThC.Tn[8].n24 VGND 0.09367f
C5984 XThC.Tn[8].t23 VGND 0.01163f
C5985 XThC.Tn[8].t20 VGND 0.0127f
C5986 XThC.Tn[8].n25 VGND 0.02837f
C5987 XThC.Tn[8].n26 VGND 0.01621f
C5988 XThC.Tn[8].n27 VGND 0.09367f
C5989 XThC.Tn[8].t39 VGND 0.01163f
C5990 XThC.Tn[8].t33 VGND 0.0127f
C5991 XThC.Tn[8].n28 VGND 0.02837f
C5992 XThC.Tn[8].n29 VGND 0.01621f
C5993 XThC.Tn[8].n30 VGND 0.09367f
C5994 XThC.Tn[8].t14 VGND 0.01163f
C5995 XThC.Tn[8].t42 VGND 0.0127f
C5996 XThC.Tn[8].n31 VGND 0.02837f
C5997 XThC.Tn[8].n32 VGND 0.01621f
C5998 XThC.Tn[8].n33 VGND 0.09367f
C5999 XThC.Tn[8].t16 VGND 0.01163f
C6000 XThC.Tn[8].t12 VGND 0.0127f
C6001 XThC.Tn[8].n34 VGND 0.02837f
C6002 XThC.Tn[8].n35 VGND 0.01621f
C6003 XThC.Tn[8].n36 VGND 0.09367f
C6004 XThC.Tn[8].t36 VGND 0.01163f
C6005 XThC.Tn[8].t31 VGND 0.0127f
C6006 XThC.Tn[8].n37 VGND 0.02837f
C6007 XThC.Tn[8].n38 VGND 0.01621f
C6008 XThC.Tn[8].n39 VGND 0.09367f
C6009 XThC.Tn[8].t38 VGND 0.01163f
C6010 XThC.Tn[8].t32 VGND 0.0127f
C6011 XThC.Tn[8].n40 VGND 0.02837f
C6012 XThC.Tn[8].n41 VGND 0.01621f
C6013 XThC.Tn[8].n42 VGND 0.09367f
C6014 XThC.Tn[8].t17 VGND 0.01163f
C6015 XThC.Tn[8].t13 VGND 0.0127f
C6016 XThC.Tn[8].n43 VGND 0.02837f
C6017 XThC.Tn[8].n44 VGND 0.01621f
C6018 XThC.Tn[8].n45 VGND 0.09367f
C6019 XThC.Tn[8].t25 VGND 0.01163f
C6020 XThC.Tn[8].t21 VGND 0.0127f
C6021 XThC.Tn[8].n46 VGND 0.02837f
C6022 XThC.Tn[8].n47 VGND 0.01621f
C6023 XThC.Tn[8].n48 VGND 0.09367f
C6024 XThC.Tn[8].t27 VGND 0.01163f
C6025 XThC.Tn[8].t24 VGND 0.0127f
C6026 XThC.Tn[8].n49 VGND 0.02837f
C6027 XThC.Tn[8].n50 VGND 0.01621f
C6028 XThC.Tn[8].n51 VGND 0.09367f
C6029 XThC.Tn[8].t40 VGND 0.01163f
C6030 XThC.Tn[8].t37 VGND 0.0127f
C6031 XThC.Tn[8].n52 VGND 0.02837f
C6032 XThC.Tn[8].n53 VGND 0.01621f
C6033 XThC.Tn[8].n54 VGND 0.09367f
C6034 XThC.Tn[8].t18 VGND 0.01163f
C6035 XThC.Tn[8].t15 VGND 0.0127f
C6036 XThC.Tn[8].n55 VGND 0.02837f
C6037 XThC.Tn[8].n56 VGND 0.01621f
C6038 XThC.Tn[8].n57 VGND 0.09367f
C6039 XThC.Tn[8].n58 VGND 0.04332f
C6040 XThC.Tn[8].n59 VGND 0.41007f
C6041 XThC.Tn[8].n60 VGND 0.03291f
C6042 XThC.XTB1.Y.t1 VGND 0.03224f
C6043 XThC.XTB1.Y.n0 VGND 0.02084f
C6044 XThC.XTB1.Y.n1 VGND 0.02659f
C6045 XThC.XTB1.Y.t2 VGND 0.01618f
C6046 XThC.XTB1.Y.t0 VGND 0.01618f
C6047 XThC.XTB1.Y.n2 VGND 0.03473f
C6048 XThC.XTB1.Y.t17 VGND 0.02517f
C6049 XThC.XTB1.Y.t5 VGND 0.01483f
C6050 XThC.XTB1.Y.n3 VGND 0.02997f
C6051 XThC.XTB1.Y.t6 VGND 0.02517f
C6052 XThC.XTB1.Y.t12 VGND 0.01483f
C6053 XThC.XTB1.Y.n4 VGND 0.01542f
C6054 XThC.XTB1.Y.t8 VGND 0.02517f
C6055 XThC.XTB1.Y.t13 VGND 0.01483f
C6056 XThC.XTB1.Y.n5 VGND 0.03313f
C6057 XThC.XTB1.Y.t11 VGND 0.02517f
C6058 XThC.XTB1.Y.t16 VGND 0.01483f
C6059 XThC.XTB1.Y.n6 VGND 0.03076f
C6060 XThC.XTB1.Y.n7 VGND 0.01871f
C6061 XThC.XTB1.Y.n8 VGND 0.03098f
C6062 XThC.XTB1.Y.n9 VGND 0.01198f
C6063 XThC.XTB1.Y.n10 VGND 0.01463f
C6064 XThC.XTB1.Y.n11 VGND 0.03313f
C6065 XThC.XTB1.Y.n12 VGND 0.01661f
C6066 XThC.XTB1.Y.n13 VGND 0.02824f
C6067 XThC.XTB1.Y.t18 VGND 0.02517f
C6068 XThC.XTB1.Y.t9 VGND 0.01483f
C6069 XThC.XTB1.Y.n14 VGND 0.03392f
C6070 XThC.XTB1.Y.t7 VGND 0.02517f
C6071 XThC.XTB1.Y.t15 VGND 0.01483f
C6072 XThC.XTB1.Y.t14 VGND 0.02517f
C6073 XThC.XTB1.Y.t3 VGND 0.01483f
C6074 XThC.XTB1.Y.t10 VGND 0.02517f
C6075 XThC.XTB1.Y.t4 VGND 0.01483f
C6076 XThC.XTB1.Y.n15 VGND 0.04223f
C6077 XThC.XTB1.Y.n16 VGND 0.0446f
C6078 XThC.XTB1.Y.n17 VGND 0.01719f
C6079 XThC.XTB1.Y.n18 VGND 0.0363f
C6080 XThC.XTB1.Y.n19 VGND 0.01661f
C6081 XThC.XTB1.Y.n20 VGND 0.01378f
C6082 XThC.XTB1.Y.n21 VGND 0.77148f
C6083 XThC.XTB1.Y.n22 VGND 0.07634f
C6084 XThC.Tn[14].n0 VGND 0.02301f
C6085 XThC.Tn[14].n1 VGND 0.01845f
C6086 XThC.Tn[14].n2 VGND 0.04642f
C6087 XThC.Tn[14].t4 VGND 0.01419f
C6088 XThC.Tn[14].t5 VGND 0.01419f
C6089 XThC.Tn[14].n3 VGND 0.03067f
C6090 XThC.Tn[14].t7 VGND 0.01419f
C6091 XThC.Tn[14].t6 VGND 0.01419f
C6092 XThC.Tn[14].n4 VGND 0.04667f
C6093 XThC.Tn[14].n5 VGND 0.12968f
C6094 XThC.Tn[14].t11 VGND 0.01419f
C6095 XThC.Tn[14].t10 VGND 0.01419f
C6096 XThC.Tn[14].n6 VGND 0.04309f
C6097 XThC.Tn[14].t9 VGND 0.01419f
C6098 XThC.Tn[14].t8 VGND 0.01419f
C6099 XThC.Tn[14].n7 VGND 0.03155f
C6100 XThC.Tn[14].n8 VGND 0.14042f
C6101 XThC.Tn[14].n9 VGND 0.02039f
C6102 XThC.Tn[14].t43 VGND 0.01125f
C6103 XThC.Tn[14].t38 VGND 0.01229f
C6104 XThC.Tn[14].n10 VGND 0.02744f
C6105 XThC.Tn[14].n11 VGND 0.01568f
C6106 XThC.Tn[14].n12 VGND 0.01907f
C6107 XThC.Tn[14].t29 VGND 0.01125f
C6108 XThC.Tn[14].t22 VGND 0.01229f
C6109 XThC.Tn[14].n13 VGND 0.02744f
C6110 XThC.Tn[14].n14 VGND 0.01568f
C6111 XThC.Tn[14].n15 VGND 0.09061f
C6112 XThC.Tn[14].t32 VGND 0.01125f
C6113 XThC.Tn[14].t25 VGND 0.01229f
C6114 XThC.Tn[14].n16 VGND 0.02744f
C6115 XThC.Tn[14].n17 VGND 0.01568f
C6116 XThC.Tn[14].n18 VGND 0.09061f
C6117 XThC.Tn[14].t34 VGND 0.01125f
C6118 XThC.Tn[14].t26 VGND 0.01229f
C6119 XThC.Tn[14].n19 VGND 0.02744f
C6120 XThC.Tn[14].n20 VGND 0.01568f
C6121 XThC.Tn[14].n21 VGND 0.09061f
C6122 XThC.Tn[14].t20 VGND 0.01125f
C6123 XThC.Tn[14].t14 VGND 0.01229f
C6124 XThC.Tn[14].n22 VGND 0.02744f
C6125 XThC.Tn[14].n23 VGND 0.01568f
C6126 XThC.Tn[14].n24 VGND 0.09061f
C6127 XThC.Tn[14].t23 VGND 0.01125f
C6128 XThC.Tn[14].t17 VGND 0.01229f
C6129 XThC.Tn[14].n25 VGND 0.02744f
C6130 XThC.Tn[14].n26 VGND 0.01568f
C6131 XThC.Tn[14].n27 VGND 0.09061f
C6132 XThC.Tn[14].t37 VGND 0.01125f
C6133 XThC.Tn[14].t31 VGND 0.01229f
C6134 XThC.Tn[14].n28 VGND 0.02744f
C6135 XThC.Tn[14].n29 VGND 0.01568f
C6136 XThC.Tn[14].n30 VGND 0.09061f
C6137 XThC.Tn[14].t13 VGND 0.01125f
C6138 XThC.Tn[14].t39 VGND 0.01229f
C6139 XThC.Tn[14].n31 VGND 0.02744f
C6140 XThC.Tn[14].n32 VGND 0.01568f
C6141 XThC.Tn[14].n33 VGND 0.09061f
C6142 XThC.Tn[14].t15 VGND 0.01125f
C6143 XThC.Tn[14].t41 VGND 0.01229f
C6144 XThC.Tn[14].n34 VGND 0.02744f
C6145 XThC.Tn[14].n35 VGND 0.01568f
C6146 XThC.Tn[14].n36 VGND 0.09061f
C6147 XThC.Tn[14].t35 VGND 0.01125f
C6148 XThC.Tn[14].t27 VGND 0.01229f
C6149 XThC.Tn[14].n37 VGND 0.02744f
C6150 XThC.Tn[14].n38 VGND 0.01568f
C6151 XThC.Tn[14].n39 VGND 0.09061f
C6152 XThC.Tn[14].t36 VGND 0.01125f
C6153 XThC.Tn[14].t30 VGND 0.01229f
C6154 XThC.Tn[14].n40 VGND 0.02744f
C6155 XThC.Tn[14].n41 VGND 0.01568f
C6156 XThC.Tn[14].n42 VGND 0.09061f
C6157 XThC.Tn[14].t16 VGND 0.01125f
C6158 XThC.Tn[14].t42 VGND 0.01229f
C6159 XThC.Tn[14].n43 VGND 0.02744f
C6160 XThC.Tn[14].n44 VGND 0.01568f
C6161 XThC.Tn[14].n45 VGND 0.09061f
C6162 XThC.Tn[14].t24 VGND 0.01125f
C6163 XThC.Tn[14].t19 VGND 0.01229f
C6164 XThC.Tn[14].n46 VGND 0.02744f
C6165 XThC.Tn[14].n47 VGND 0.01568f
C6166 XThC.Tn[14].n48 VGND 0.09061f
C6167 XThC.Tn[14].t28 VGND 0.01125f
C6168 XThC.Tn[14].t21 VGND 0.01229f
C6169 XThC.Tn[14].n49 VGND 0.02744f
C6170 XThC.Tn[14].n50 VGND 0.01568f
C6171 XThC.Tn[14].n51 VGND 0.09061f
C6172 XThC.Tn[14].t40 VGND 0.01125f
C6173 XThC.Tn[14].t33 VGND 0.01229f
C6174 XThC.Tn[14].n52 VGND 0.02744f
C6175 XThC.Tn[14].n53 VGND 0.01568f
C6176 XThC.Tn[14].n54 VGND 0.09061f
C6177 XThC.Tn[14].t18 VGND 0.01125f
C6178 XThC.Tn[14].t12 VGND 0.01229f
C6179 XThC.Tn[14].n55 VGND 0.02744f
C6180 XThC.Tn[14].n56 VGND 0.01568f
C6181 XThC.Tn[14].n57 VGND 0.09061f
C6182 XThC.Tn[14].n58 VGND 0.54091f
C6183 XThC.Tn[14].n59 VGND 0.03454f
C6184 XThR.Tn[10].t4 VGND 0.01941f
C6185 XThR.Tn[10].t2 VGND 0.01941f
C6186 XThR.Tn[10].n0 VGND 0.05892f
C6187 XThR.Tn[10].t5 VGND 0.01941f
C6188 XThR.Tn[10].t3 VGND 0.01941f
C6189 XThR.Tn[10].n1 VGND 0.04314f
C6190 XThR.Tn[10].n2 VGND 0.19615f
C6191 XThR.Tn[10].t6 VGND 0.01941f
C6192 XThR.Tn[10].t10 VGND 0.01941f
C6193 XThR.Tn[10].n3 VGND 0.04193f
C6194 XThR.Tn[10].t7 VGND 0.01941f
C6195 XThR.Tn[10].t9 VGND 0.01941f
C6196 XThR.Tn[10].n4 VGND 0.06382f
C6197 XThR.Tn[10].n5 VGND 0.1772f
C6198 XThR.Tn[10].t54 VGND 0.01517f
C6199 XThR.Tn[10].t47 VGND 0.01661f
C6200 XThR.Tn[10].n7 VGND 0.04056f
C6201 XThR.Tn[10].n8 VGND 0.07791f
C6202 XThR.Tn[10].t13 VGND 0.01517f
C6203 XThR.Tn[10].t63 VGND 0.01661f
C6204 XThR.Tn[10].n9 VGND 0.04056f
C6205 XThR.Tn[10].t50 VGND 0.01512f
C6206 XThR.Tn[10].t60 VGND 0.01655f
C6207 XThR.Tn[10].n10 VGND 0.0422f
C6208 XThR.Tn[10].n11 VGND 0.02964f
C6209 XThR.Tn[10].n13 VGND 0.09513f
C6210 XThR.Tn[10].t48 VGND 0.01517f
C6211 XThR.Tn[10].t41 VGND 0.01661f
C6212 XThR.Tn[10].n14 VGND 0.04056f
C6213 XThR.Tn[10].t23 VGND 0.01512f
C6214 XThR.Tn[10].t36 VGND 0.01655f
C6215 XThR.Tn[10].n15 VGND 0.0422f
C6216 XThR.Tn[10].n16 VGND 0.02964f
C6217 XThR.Tn[10].n18 VGND 0.09513f
C6218 XThR.Tn[10].t65 VGND 0.01517f
C6219 XThR.Tn[10].t58 VGND 0.01661f
C6220 XThR.Tn[10].n19 VGND 0.04056f
C6221 XThR.Tn[10].t40 VGND 0.01512f
C6222 XThR.Tn[10].t55 VGND 0.01655f
C6223 XThR.Tn[10].n20 VGND 0.0422f
C6224 XThR.Tn[10].n21 VGND 0.02964f
C6225 XThR.Tn[10].n23 VGND 0.09513f
C6226 XThR.Tn[10].t30 VGND 0.01517f
C6227 XThR.Tn[10].t26 VGND 0.01661f
C6228 XThR.Tn[10].n24 VGND 0.04056f
C6229 XThR.Tn[10].t70 VGND 0.01512f
C6230 XThR.Tn[10].t21 VGND 0.01655f
C6231 XThR.Tn[10].n25 VGND 0.0422f
C6232 XThR.Tn[10].n26 VGND 0.02964f
C6233 XThR.Tn[10].n28 VGND 0.09513f
C6234 XThR.Tn[10].t67 VGND 0.01517f
C6235 XThR.Tn[10].t59 VGND 0.01661f
C6236 XThR.Tn[10].n29 VGND 0.04056f
C6237 XThR.Tn[10].t42 VGND 0.01512f
C6238 XThR.Tn[10].t56 VGND 0.01655f
C6239 XThR.Tn[10].n30 VGND 0.0422f
C6240 XThR.Tn[10].n31 VGND 0.02964f
C6241 XThR.Tn[10].n33 VGND 0.09513f
C6242 XThR.Tn[10].t44 VGND 0.01517f
C6243 XThR.Tn[10].t15 VGND 0.01661f
C6244 XThR.Tn[10].n34 VGND 0.04056f
C6245 XThR.Tn[10].t18 VGND 0.01512f
C6246 XThR.Tn[10].t12 VGND 0.01655f
C6247 XThR.Tn[10].n35 VGND 0.0422f
C6248 XThR.Tn[10].n36 VGND 0.02964f
C6249 XThR.Tn[10].n38 VGND 0.09513f
C6250 XThR.Tn[10].t14 VGND 0.01517f
C6251 XThR.Tn[10].t69 VGND 0.01661f
C6252 XThR.Tn[10].n39 VGND 0.04056f
C6253 XThR.Tn[10].t51 VGND 0.01512f
C6254 XThR.Tn[10].t66 VGND 0.01655f
C6255 XThR.Tn[10].n40 VGND 0.0422f
C6256 XThR.Tn[10].n41 VGND 0.02964f
C6257 XThR.Tn[10].n43 VGND 0.09513f
C6258 XThR.Tn[10].t17 VGND 0.01517f
C6259 XThR.Tn[10].t24 VGND 0.01661f
C6260 XThR.Tn[10].n44 VGND 0.04056f
C6261 XThR.Tn[10].t53 VGND 0.01512f
C6262 XThR.Tn[10].t20 VGND 0.01655f
C6263 XThR.Tn[10].n45 VGND 0.0422f
C6264 XThR.Tn[10].n46 VGND 0.02964f
C6265 XThR.Tn[10].n48 VGND 0.09513f
C6266 XThR.Tn[10].t33 VGND 0.01517f
C6267 XThR.Tn[10].t43 VGND 0.01661f
C6268 XThR.Tn[10].n49 VGND 0.04056f
C6269 XThR.Tn[10].t73 VGND 0.01512f
C6270 XThR.Tn[10].t38 VGND 0.01655f
C6271 XThR.Tn[10].n50 VGND 0.0422f
C6272 XThR.Tn[10].n51 VGND 0.02964f
C6273 XThR.Tn[10].n53 VGND 0.09513f
C6274 XThR.Tn[10].t28 VGND 0.01517f
C6275 XThR.Tn[10].t61 VGND 0.01661f
C6276 XThR.Tn[10].n54 VGND 0.04056f
C6277 XThR.Tn[10].t62 VGND 0.01512f
C6278 XThR.Tn[10].t57 VGND 0.01655f
C6279 XThR.Tn[10].n55 VGND 0.0422f
C6280 XThR.Tn[10].n56 VGND 0.02964f
C6281 XThR.Tn[10].n58 VGND 0.09513f
C6282 XThR.Tn[10].t46 VGND 0.01517f
C6283 XThR.Tn[10].t35 VGND 0.01661f
C6284 XThR.Tn[10].n59 VGND 0.04056f
C6285 XThR.Tn[10].t19 VGND 0.01512f
C6286 XThR.Tn[10].t32 VGND 0.01655f
C6287 XThR.Tn[10].n60 VGND 0.0422f
C6288 XThR.Tn[10].n61 VGND 0.02964f
C6289 XThR.Tn[10].n63 VGND 0.09513f
C6290 XThR.Tn[10].t16 VGND 0.01517f
C6291 XThR.Tn[10].t72 VGND 0.01661f
C6292 XThR.Tn[10].n64 VGND 0.04056f
C6293 XThR.Tn[10].t52 VGND 0.01512f
C6294 XThR.Tn[10].t68 VGND 0.01655f
C6295 XThR.Tn[10].n65 VGND 0.0422f
C6296 XThR.Tn[10].n66 VGND 0.02964f
C6297 XThR.Tn[10].n68 VGND 0.09513f
C6298 XThR.Tn[10].t31 VGND 0.01517f
C6299 XThR.Tn[10].t27 VGND 0.01661f
C6300 XThR.Tn[10].n69 VGND 0.04056f
C6301 XThR.Tn[10].t71 VGND 0.01512f
C6302 XThR.Tn[10].t22 VGND 0.01655f
C6303 XThR.Tn[10].n70 VGND 0.0422f
C6304 XThR.Tn[10].n71 VGND 0.02964f
C6305 XThR.Tn[10].n73 VGND 0.09513f
C6306 XThR.Tn[10].t49 VGND 0.01517f
C6307 XThR.Tn[10].t45 VGND 0.01661f
C6308 XThR.Tn[10].n74 VGND 0.04056f
C6309 XThR.Tn[10].t25 VGND 0.01512f
C6310 XThR.Tn[10].t39 VGND 0.01655f
C6311 XThR.Tn[10].n75 VGND 0.0422f
C6312 XThR.Tn[10].n76 VGND 0.02964f
C6313 XThR.Tn[10].n78 VGND 0.09513f
C6314 XThR.Tn[10].t29 VGND 0.01517f
C6315 XThR.Tn[10].t37 VGND 0.01661f
C6316 XThR.Tn[10].n79 VGND 0.04056f
C6317 XThR.Tn[10].t64 VGND 0.01512f
C6318 XThR.Tn[10].t34 VGND 0.01655f
C6319 XThR.Tn[10].n80 VGND 0.0422f
C6320 XThR.Tn[10].n81 VGND 0.02964f
C6321 XThR.Tn[10].n83 VGND 0.09513f
C6322 XThR.Tn[10].n84 VGND 0.08645f
C6323 XThR.Tn[10].n85 VGND 0.26614f
C6324 XThR.Tn[10].t11 VGND 0.01261f
C6325 XThR.Tn[10].t1 VGND 0.01261f
C6326 XThR.Tn[10].n86 VGND 0.03146f
C6327 XThR.Tn[10].t0 VGND 0.01261f
C6328 XThR.Tn[10].t8 VGND 0.01261f
C6329 XThR.Tn[10].n87 VGND 0.02523f
C6330 XThR.Tn[10].n88 VGND 0.05817f
C6331 XThC.Tn[3].t5 VGND 0.01185f
C6332 XThC.Tn[3].t4 VGND 0.01185f
C6333 XThC.Tn[3].n0 VGND 0.02391f
C6334 XThC.Tn[3].t7 VGND 0.01185f
C6335 XThC.Tn[3].t6 VGND 0.01185f
C6336 XThC.Tn[3].n1 VGND 0.02797f
C6337 XThC.Tn[3].n2 VGND 0.08391f
C6338 XThC.Tn[3].n3 VGND 0.01753f
C6339 XThC.Tn[3].n4 VGND 0.02921f
C6340 XThC.Tn[3].n5 VGND 0.01753f
C6341 XThC.Tn[3].n6 VGND 0.0835f
C6342 XThC.Tn[3].n7 VGND 0.01753f
C6343 XThC.Tn[3].n8 VGND 0.05162f
C6344 XThC.Tn[3].n9 VGND 0.05825f
C6345 XThC.Tn[3].t42 VGND 0.01025f
C6346 XThC.Tn[3].n10 VGND 0.0229f
C6347 XThC.Tn[3].n11 VGND 0.01309f
C6348 XThC.Tn[3].n12 VGND 0.01592f
C6349 XThC.Tn[3].t27 VGND 0.01025f
C6350 XThC.Tn[3].n13 VGND 0.0229f
C6351 XThC.Tn[3].n14 VGND 0.01309f
C6352 XThC.Tn[3].n15 VGND 0.07562f
C6353 XThC.Tn[3].t29 VGND 0.01025f
C6354 XThC.Tn[3].n16 VGND 0.0229f
C6355 XThC.Tn[3].n17 VGND 0.01309f
C6356 XThC.Tn[3].n18 VGND 0.07562f
C6357 XThC.Tn[3].t31 VGND 0.01025f
C6358 XThC.Tn[3].n19 VGND 0.0229f
C6359 XThC.Tn[3].n20 VGND 0.01309f
C6360 XThC.Tn[3].n21 VGND 0.07562f
C6361 XThC.Tn[3].t20 VGND 0.01025f
C6362 XThC.Tn[3].n22 VGND 0.0229f
C6363 XThC.Tn[3].n23 VGND 0.01309f
C6364 XThC.Tn[3].n24 VGND 0.07562f
C6365 XThC.Tn[3].t21 VGND 0.01025f
C6366 XThC.Tn[3].n25 VGND 0.0229f
C6367 XThC.Tn[3].n26 VGND 0.01309f
C6368 XThC.Tn[3].n27 VGND 0.07562f
C6369 XThC.Tn[3].t34 VGND 0.01025f
C6370 XThC.Tn[3].n28 VGND 0.0229f
C6371 XThC.Tn[3].n29 VGND 0.01309f
C6372 XThC.Tn[3].n30 VGND 0.07562f
C6373 XThC.Tn[3].t43 VGND 0.01025f
C6374 XThC.Tn[3].n31 VGND 0.0229f
C6375 XThC.Tn[3].n32 VGND 0.01309f
C6376 XThC.Tn[3].n33 VGND 0.07562f
C6377 XThC.Tn[3].t13 VGND 0.01025f
C6378 XThC.Tn[3].n34 VGND 0.0229f
C6379 XThC.Tn[3].n35 VGND 0.01309f
C6380 XThC.Tn[3].n36 VGND 0.07562f
C6381 XThC.Tn[3].t32 VGND 0.01025f
C6382 XThC.Tn[3].n37 VGND 0.0229f
C6383 XThC.Tn[3].n38 VGND 0.01309f
C6384 XThC.Tn[3].n39 VGND 0.07562f
C6385 XThC.Tn[3].t33 VGND 0.01025f
C6386 XThC.Tn[3].n40 VGND 0.0229f
C6387 XThC.Tn[3].n41 VGND 0.01309f
C6388 XThC.Tn[3].n42 VGND 0.07562f
C6389 XThC.Tn[3].t14 VGND 0.01025f
C6390 XThC.Tn[3].n43 VGND 0.0229f
C6391 XThC.Tn[3].n44 VGND 0.01309f
C6392 XThC.Tn[3].n45 VGND 0.07562f
C6393 XThC.Tn[3].t22 VGND 0.01025f
C6394 XThC.Tn[3].n46 VGND 0.0229f
C6395 XThC.Tn[3].n47 VGND 0.01309f
C6396 XThC.Tn[3].n48 VGND 0.07562f
C6397 XThC.Tn[3].t25 VGND 0.01025f
C6398 XThC.Tn[3].n49 VGND 0.0229f
C6399 XThC.Tn[3].n50 VGND 0.01309f
C6400 XThC.Tn[3].n51 VGND 0.07562f
C6401 XThC.Tn[3].t38 VGND 0.01025f
C6402 XThC.Tn[3].n52 VGND 0.0229f
C6403 XThC.Tn[3].n53 VGND 0.01309f
C6404 XThC.Tn[3].n54 VGND 0.07562f
C6405 XThC.Tn[3].t16 VGND 0.01025f
C6406 XThC.Tn[3].n55 VGND 0.0229f
C6407 XThC.Tn[3].n56 VGND 0.01309f
C6408 XThC.Tn[3].n57 VGND 0.07562f
C6409 XThC.Tn[3].n58 VGND 0.03994f
C6410 XThC.Tn[1].t11 VGND 0.0116f
C6411 XThC.Tn[1].t10 VGND 0.0116f
C6412 XThC.Tn[1].n0 VGND 0.02342f
C6413 XThC.Tn[1].t9 VGND 0.0116f
C6414 XThC.Tn[1].t8 VGND 0.0116f
C6415 XThC.Tn[1].n1 VGND 0.02741f
C6416 XThC.Tn[1].n2 VGND 0.08221f
C6417 XThC.Tn[1].n3 VGND 0.01718f
C6418 XThC.Tn[1].n4 VGND 0.01718f
C6419 XThC.Tn[1].n5 VGND 0.01718f
C6420 XThC.Tn[1].n6 VGND 0.02862f
C6421 XThC.Tn[1].n7 VGND 0.0818f
C6422 XThC.Tn[1].n8 VGND 0.05057f
C6423 XThC.Tn[1].n9 VGND 0.05707f
C6424 XThC.Tn[1].t29 VGND 0.01005f
C6425 XThC.Tn[1].n10 VGND 0.02244f
C6426 XThC.Tn[1].n11 VGND 0.01282f
C6427 XThC.Tn[1].n12 VGND 0.01559f
C6428 XThC.Tn[1].t14 VGND 0.01005f
C6429 XThC.Tn[1].n13 VGND 0.02244f
C6430 XThC.Tn[1].n14 VGND 0.01282f
C6431 XThC.Tn[1].n15 VGND 0.07408f
C6432 XThC.Tn[1].t16 VGND 0.01005f
C6433 XThC.Tn[1].n16 VGND 0.02244f
C6434 XThC.Tn[1].n17 VGND 0.01282f
C6435 XThC.Tn[1].n18 VGND 0.07408f
C6436 XThC.Tn[1].t18 VGND 0.01005f
C6437 XThC.Tn[1].n19 VGND 0.02244f
C6438 XThC.Tn[1].n20 VGND 0.01282f
C6439 XThC.Tn[1].n21 VGND 0.07408f
C6440 XThC.Tn[1].t39 VGND 0.01005f
C6441 XThC.Tn[1].n22 VGND 0.02244f
C6442 XThC.Tn[1].n23 VGND 0.01282f
C6443 XThC.Tn[1].n24 VGND 0.07408f
C6444 XThC.Tn[1].t40 VGND 0.01005f
C6445 XThC.Tn[1].n25 VGND 0.02244f
C6446 XThC.Tn[1].n26 VGND 0.01282f
C6447 XThC.Tn[1].n27 VGND 0.07408f
C6448 XThC.Tn[1].t21 VGND 0.01005f
C6449 XThC.Tn[1].n28 VGND 0.02244f
C6450 XThC.Tn[1].n29 VGND 0.01282f
C6451 XThC.Tn[1].n30 VGND 0.07408f
C6452 XThC.Tn[1].t30 VGND 0.01005f
C6453 XThC.Tn[1].n31 VGND 0.02244f
C6454 XThC.Tn[1].n32 VGND 0.01282f
C6455 XThC.Tn[1].n33 VGND 0.07408f
C6456 XThC.Tn[1].t32 VGND 0.01005f
C6457 XThC.Tn[1].n34 VGND 0.02244f
C6458 XThC.Tn[1].n35 VGND 0.01282f
C6459 XThC.Tn[1].n36 VGND 0.07408f
C6460 XThC.Tn[1].t19 VGND 0.01005f
C6461 XThC.Tn[1].n37 VGND 0.02244f
C6462 XThC.Tn[1].n38 VGND 0.01282f
C6463 XThC.Tn[1].n39 VGND 0.07408f
C6464 XThC.Tn[1].t20 VGND 0.01005f
C6465 XThC.Tn[1].n40 VGND 0.02244f
C6466 XThC.Tn[1].n41 VGND 0.01282f
C6467 XThC.Tn[1].n42 VGND 0.07408f
C6468 XThC.Tn[1].t33 VGND 0.01005f
C6469 XThC.Tn[1].n43 VGND 0.02244f
C6470 XThC.Tn[1].n44 VGND 0.01282f
C6471 XThC.Tn[1].n45 VGND 0.07408f
C6472 XThC.Tn[1].t41 VGND 0.01005f
C6473 XThC.Tn[1].n46 VGND 0.02244f
C6474 XThC.Tn[1].n47 VGND 0.01282f
C6475 XThC.Tn[1].n48 VGND 0.07408f
C6476 XThC.Tn[1].t12 VGND 0.01005f
C6477 XThC.Tn[1].n49 VGND 0.02244f
C6478 XThC.Tn[1].n50 VGND 0.01282f
C6479 XThC.Tn[1].n51 VGND 0.07408f
C6480 XThC.Tn[1].t25 VGND 0.01005f
C6481 XThC.Tn[1].n52 VGND 0.02244f
C6482 XThC.Tn[1].n53 VGND 0.01282f
C6483 XThC.Tn[1].n54 VGND 0.07408f
C6484 XThC.Tn[1].t35 VGND 0.01005f
C6485 XThC.Tn[1].n55 VGND 0.02244f
C6486 XThC.Tn[1].n56 VGND 0.01282f
C6487 XThC.Tn[1].n57 VGND 0.07408f
C6488 XThC.Tn[1].n58 VGND 0.27353f
C6489 XThC.Tn[1].n59 VGND 0.0276f
C6490 Vbias.t266 VGND 0.1745f
C6491 Vbias.n0 VGND 0.18997f
C6492 Vbias.t85 VGND 0.1745f
C6493 Vbias.n1 VGND 0.1903f
C6494 Vbias.n2 VGND 0.1262f
C6495 Vbias.t180 VGND 0.1745f
C6496 Vbias.n3 VGND 0.1903f
C6497 Vbias.n4 VGND 0.1262f
C6498 Vbias.t188 VGND 0.1745f
C6499 Vbias.n5 VGND 0.1903f
C6500 Vbias.n6 VGND 0.1262f
C6501 Vbias.t21 VGND 0.1745f
C6502 Vbias.n7 VGND 0.1903f
C6503 Vbias.n8 VGND 0.1262f
C6504 Vbias.t107 VGND 0.1745f
C6505 Vbias.n9 VGND 0.1903f
C6506 Vbias.n10 VGND 0.1262f
C6507 Vbias.t190 VGND 0.1745f
C6508 Vbias.n11 VGND 0.1903f
C6509 Vbias.n12 VGND 0.1262f
C6510 Vbias.t25 VGND 0.1745f
C6511 Vbias.n13 VGND 0.1903f
C6512 Vbias.n14 VGND 0.1262f
C6513 Vbias.t45 VGND 0.1745f
C6514 Vbias.n15 VGND 0.1903f
C6515 Vbias.n16 VGND 0.1262f
C6516 Vbias.t117 VGND 0.1745f
C6517 Vbias.n17 VGND 0.1903f
C6518 Vbias.n18 VGND 0.1262f
C6519 Vbias.t208 VGND 0.1745f
C6520 Vbias.n19 VGND 0.1903f
C6521 Vbias.n20 VGND 0.1262f
C6522 Vbias.t229 VGND 0.1745f
C6523 Vbias.n21 VGND 0.1903f
C6524 Vbias.n22 VGND 0.1262f
C6525 Vbias.t120 VGND 0.1745f
C6526 Vbias.n23 VGND 0.1903f
C6527 Vbias.n24 VGND 0.1262f
C6528 Vbias.t148 VGND 0.1745f
C6529 Vbias.n25 VGND 0.1903f
C6530 Vbias.n26 VGND 0.1262f
C6531 Vbias.t157 VGND 0.1745f
C6532 Vbias.n27 VGND 0.1903f
C6533 Vbias.n28 VGND 0.1262f
C6534 Vbias.t67 VGND 0.1745f
C6535 Vbias.n29 VGND 0.1903f
C6536 Vbias.n30 VGND 0.1262f
C6537 Vbias.n31 VGND 0.5296f
C6538 Vbias.t146 VGND 0.1745f
C6539 Vbias.n32 VGND 0.18997f
C6540 Vbias.t222 VGND 0.1745f
C6541 Vbias.n33 VGND 0.1903f
C6542 Vbias.n34 VGND 0.1262f
C6543 Vbias.t65 VGND 0.1745f
C6544 Vbias.n35 VGND 0.1903f
C6545 Vbias.n36 VGND 0.1262f
C6546 Vbias.t73 VGND 0.1745f
C6547 Vbias.n37 VGND 0.1903f
C6548 Vbias.n38 VGND 0.1262f
C6549 Vbias.t158 VGND 0.1745f
C6550 Vbias.n39 VGND 0.1903f
C6551 Vbias.n40 VGND 0.1262f
C6552 Vbias.t251 VGND 0.1745f
C6553 Vbias.n41 VGND 0.1903f
C6554 Vbias.n42 VGND 0.1262f
C6555 Vbias.t78 VGND 0.1745f
C6556 Vbias.n43 VGND 0.1903f
C6557 Vbias.n44 VGND 0.1262f
C6558 Vbias.t164 VGND 0.1745f
C6559 Vbias.n45 VGND 0.1903f
C6560 Vbias.n46 VGND 0.1262f
C6561 Vbias.t184 VGND 0.1745f
C6562 Vbias.n47 VGND 0.1903f
C6563 Vbias.n48 VGND 0.1262f
C6564 Vbias.t260 VGND 0.1745f
C6565 Vbias.n49 VGND 0.1903f
C6566 Vbias.n50 VGND 0.1262f
C6567 Vbias.t90 VGND 0.1745f
C6568 Vbias.n51 VGND 0.1903f
C6569 Vbias.n52 VGND 0.1262f
C6570 Vbias.t112 VGND 0.1745f
C6571 Vbias.n53 VGND 0.1903f
C6572 Vbias.n54 VGND 0.1262f
C6573 Vbias.t265 VGND 0.1745f
C6574 Vbias.n55 VGND 0.1903f
C6575 Vbias.n56 VGND 0.1262f
C6576 Vbias.t32 VGND 0.1745f
C6577 Vbias.n57 VGND 0.1903f
C6578 Vbias.n58 VGND 0.1262f
C6579 Vbias.t41 VGND 0.1745f
C6580 Vbias.n59 VGND 0.1903f
C6581 Vbias.n60 VGND 0.1262f
C6582 Vbias.t200 VGND 0.1745f
C6583 Vbias.n61 VGND 0.1903f
C6584 Vbias.n62 VGND 0.1262f
C6585 Vbias.n63 VGND 0.54484f
C6586 Vbias.t221 VGND 0.1745f
C6587 Vbias.n64 VGND 0.18997f
C6588 Vbias.t37 VGND 0.1745f
C6589 Vbias.n65 VGND 0.1903f
C6590 Vbias.n66 VGND 0.1262f
C6591 Vbias.t138 VGND 0.1745f
C6592 Vbias.n67 VGND 0.1903f
C6593 Vbias.n68 VGND 0.1262f
C6594 Vbias.t145 VGND 0.1745f
C6595 Vbias.n69 VGND 0.1903f
C6596 Vbias.n70 VGND 0.1262f
C6597 Vbias.t230 VGND 0.1745f
C6598 Vbias.n71 VGND 0.1903f
C6599 Vbias.n72 VGND 0.1262f
C6600 Vbias.t64 VGND 0.1745f
C6601 Vbias.n73 VGND 0.1903f
C6602 Vbias.n74 VGND 0.1262f
C6603 Vbias.t151 VGND 0.1745f
C6604 Vbias.n75 VGND 0.1903f
C6605 Vbias.n76 VGND 0.1262f
C6606 Vbias.t236 VGND 0.1745f
C6607 Vbias.n77 VGND 0.1903f
C6608 Vbias.n78 VGND 0.1262f
C6609 Vbias.t259 VGND 0.1745f
C6610 Vbias.n79 VGND 0.1903f
C6611 Vbias.n80 VGND 0.1262f
C6612 Vbias.t77 VGND 0.1745f
C6613 Vbias.n81 VGND 0.1903f
C6614 Vbias.n82 VGND 0.1262f
C6615 Vbias.t163 VGND 0.1745f
C6616 Vbias.n83 VGND 0.1903f
C6617 Vbias.n84 VGND 0.1262f
C6618 Vbias.t183 VGND 0.1745f
C6619 Vbias.n85 VGND 0.1903f
C6620 Vbias.n86 VGND 0.1262f
C6621 Vbias.t83 VGND 0.1745f
C6622 Vbias.n87 VGND 0.1903f
C6623 Vbias.n88 VGND 0.1262f
C6624 Vbias.t103 VGND 0.1745f
C6625 Vbias.n89 VGND 0.1903f
C6626 Vbias.n90 VGND 0.1262f
C6627 Vbias.t110 VGND 0.1745f
C6628 Vbias.n91 VGND 0.1903f
C6629 Vbias.n92 VGND 0.1262f
C6630 Vbias.t19 VGND 0.1745f
C6631 Vbias.n93 VGND 0.1903f
C6632 Vbias.n94 VGND 0.1262f
C6633 Vbias.n95 VGND 0.54484f
C6634 Vbias.t36 VGND 0.1745f
C6635 Vbias.n96 VGND 0.18997f
C6636 Vbias.t106 VGND 0.1745f
C6637 Vbias.n97 VGND 0.1903f
C6638 Vbias.n98 VGND 0.1262f
C6639 Vbias.t209 VGND 0.1745f
C6640 Vbias.n99 VGND 0.1903f
C6641 Vbias.n100 VGND 0.1262f
C6642 Vbias.t220 VGND 0.1745f
C6643 Vbias.n101 VGND 0.1903f
C6644 Vbias.n102 VGND 0.1262f
C6645 Vbias.t44 VGND 0.1745f
C6646 Vbias.n103 VGND 0.1903f
C6647 Vbias.n104 VGND 0.1262f
C6648 Vbias.t137 VGND 0.1745f
C6649 Vbias.n105 VGND 0.1903f
C6650 Vbias.n106 VGND 0.1262f
C6651 Vbias.t224 VGND 0.1745f
C6652 Vbias.n107 VGND 0.1903f
C6653 Vbias.n108 VGND 0.1262f
C6654 Vbias.t48 VGND 0.1745f
C6655 Vbias.n109 VGND 0.1903f
C6656 Vbias.n110 VGND 0.1262f
C6657 Vbias.t76 VGND 0.1745f
C6658 Vbias.n111 VGND 0.1903f
C6659 Vbias.n112 VGND 0.1262f
C6660 Vbias.t149 VGND 0.1745f
C6661 Vbias.n113 VGND 0.1903f
C6662 Vbias.n114 VGND 0.1262f
C6663 Vbias.t234 VGND 0.1745f
C6664 Vbias.n115 VGND 0.1903f
C6665 Vbias.n116 VGND 0.1262f
C6666 Vbias.t258 VGND 0.1745f
C6667 Vbias.n117 VGND 0.1903f
C6668 Vbias.n118 VGND 0.1262f
C6669 Vbias.t154 VGND 0.1745f
C6670 Vbias.n119 VGND 0.1903f
C6671 Vbias.n120 VGND 0.1262f
C6672 Vbias.t176 VGND 0.1745f
C6673 Vbias.n121 VGND 0.1903f
C6674 Vbias.n122 VGND 0.1262f
C6675 Vbias.t181 VGND 0.1745f
C6676 Vbias.n123 VGND 0.1903f
C6677 Vbias.n124 VGND 0.1262f
C6678 Vbias.t92 VGND 0.1745f
C6679 Vbias.n125 VGND 0.1903f
C6680 Vbias.n126 VGND 0.1262f
C6681 Vbias.n127 VGND 0.54484f
C6682 Vbias.t192 VGND 0.1745f
C6683 Vbias.n128 VGND 0.18997f
C6684 Vbias.t12 VGND 0.1745f
C6685 Vbias.n129 VGND 0.1903f
C6686 Vbias.n130 VGND 0.1262f
C6687 Vbias.t109 VGND 0.1745f
C6688 Vbias.n131 VGND 0.1903f
C6689 Vbias.n132 VGND 0.1262f
C6690 Vbias.t121 VGND 0.1745f
C6691 Vbias.n133 VGND 0.1903f
C6692 Vbias.n134 VGND 0.1262f
C6693 Vbias.t212 VGND 0.1745f
C6694 Vbias.n135 VGND 0.1903f
C6695 Vbias.n136 VGND 0.1262f
C6696 Vbias.t40 VGND 0.1745f
C6697 Vbias.n137 VGND 0.1903f
C6698 Vbias.n138 VGND 0.1262f
C6699 Vbias.t122 VGND 0.1745f
C6700 Vbias.n139 VGND 0.1903f
C6701 Vbias.n140 VGND 0.1262f
C6702 Vbias.t215 VGND 0.1745f
C6703 Vbias.n141 VGND 0.1903f
C6704 Vbias.n142 VGND 0.1262f
C6705 Vbias.t237 VGND 0.1745f
C6706 Vbias.n143 VGND 0.1903f
C6707 Vbias.n144 VGND 0.1262f
C6708 Vbias.t49 VGND 0.1745f
C6709 Vbias.n145 VGND 0.1903f
C6710 Vbias.n146 VGND 0.1262f
C6711 Vbias.t140 VGND 0.1745f
C6712 Vbias.n147 VGND 0.1903f
C6713 Vbias.n148 VGND 0.1262f
C6714 Vbias.t165 VGND 0.1745f
C6715 Vbias.n149 VGND 0.1903f
C6716 Vbias.n150 VGND 0.1262f
C6717 Vbias.t53 VGND 0.1745f
C6718 Vbias.n151 VGND 0.1903f
C6719 Vbias.n152 VGND 0.1262f
C6720 Vbias.t84 VGND 0.1745f
C6721 Vbias.n153 VGND 0.1903f
C6722 Vbias.n154 VGND 0.1262f
C6723 Vbias.t91 VGND 0.1745f
C6724 Vbias.n155 VGND 0.1903f
C6725 Vbias.n156 VGND 0.1262f
C6726 Vbias.t255 VGND 0.1745f
C6727 Vbias.n157 VGND 0.1903f
C6728 Vbias.n158 VGND 0.1262f
C6729 Vbias.n159 VGND 0.54484f
C6730 Vbias.t61 VGND 0.1745f
C6731 Vbias.n160 VGND 0.18997f
C6732 Vbias.t134 VGND 0.1745f
C6733 Vbias.n161 VGND 0.1903f
C6734 Vbias.n162 VGND 0.1262f
C6735 Vbias.t232 VGND 0.1745f
C6736 Vbias.n163 VGND 0.1903f
C6737 Vbias.n164 VGND 0.1262f
C6738 Vbias.t247 VGND 0.1745f
C6739 Vbias.n165 VGND 0.1903f
C6740 Vbias.n166 VGND 0.1262f
C6741 Vbias.t72 VGND 0.1745f
C6742 Vbias.n167 VGND 0.1903f
C6743 Vbias.n168 VGND 0.1262f
C6744 Vbias.t161 VGND 0.1745f
C6745 Vbias.n169 VGND 0.1903f
C6746 Vbias.n170 VGND 0.1262f
C6747 Vbias.t250 VGND 0.1745f
C6748 Vbias.n171 VGND 0.1903f
C6749 Vbias.n172 VGND 0.1262f
C6750 Vbias.t80 VGND 0.1745f
C6751 Vbias.n173 VGND 0.1903f
C6752 Vbias.n174 VGND 0.1262f
C6753 Vbias.t100 VGND 0.1745f
C6754 Vbias.n175 VGND 0.1903f
C6755 Vbias.n176 VGND 0.1262f
C6756 Vbias.t173 VGND 0.1745f
C6757 Vbias.n177 VGND 0.1903f
C6758 Vbias.n178 VGND 0.1262f
C6759 Vbias.t262 VGND 0.1745f
C6760 Vbias.n179 VGND 0.1903f
C6761 Vbias.n180 VGND 0.1262f
C6762 Vbias.t28 VGND 0.1745f
C6763 Vbias.n181 VGND 0.1903f
C6764 Vbias.n182 VGND 0.1262f
C6765 Vbias.t178 VGND 0.1745f
C6766 Vbias.n183 VGND 0.1903f
C6767 Vbias.n184 VGND 0.1262f
C6768 Vbias.t197 VGND 0.1745f
C6769 Vbias.n185 VGND 0.1903f
C6770 Vbias.n186 VGND 0.1262f
C6771 Vbias.t213 VGND 0.1745f
C6772 Vbias.n187 VGND 0.1903f
C6773 Vbias.n188 VGND 0.1262f
C6774 Vbias.t115 VGND 0.1745f
C6775 Vbias.n189 VGND 0.1903f
C6776 Vbias.n190 VGND 0.1262f
C6777 Vbias.n191 VGND 0.54484f
C6778 Vbias.t195 VGND 0.1745f
C6779 Vbias.n192 VGND 0.18997f
C6780 Vbias.t16 VGND 0.1745f
C6781 Vbias.n193 VGND 0.1903f
C6782 Vbias.n194 VGND 0.1262f
C6783 Vbias.t114 VGND 0.1745f
C6784 Vbias.n195 VGND 0.1903f
C6785 Vbias.n196 VGND 0.1262f
C6786 Vbias.t123 VGND 0.1745f
C6787 Vbias.n197 VGND 0.1903f
C6788 Vbias.n198 VGND 0.1262f
C6789 Vbias.t214 VGND 0.1745f
C6790 Vbias.n199 VGND 0.1903f
C6791 Vbias.n200 VGND 0.1262f
C6792 Vbias.t42 VGND 0.1745f
C6793 Vbias.n201 VGND 0.1903f
C6794 Vbias.n202 VGND 0.1262f
C6795 Vbias.t126 VGND 0.1745f
C6796 Vbias.n203 VGND 0.1903f
C6797 Vbias.n204 VGND 0.1262f
C6798 Vbias.t218 VGND 0.1745f
C6799 Vbias.n205 VGND 0.1903f
C6800 Vbias.n206 VGND 0.1262f
C6801 Vbias.t240 VGND 0.1745f
C6802 Vbias.n207 VGND 0.1903f
C6803 Vbias.n208 VGND 0.1262f
C6804 Vbias.t52 VGND 0.1745f
C6805 Vbias.n209 VGND 0.1903f
C6806 Vbias.n210 VGND 0.1262f
C6807 Vbias.t142 VGND 0.1745f
C6808 Vbias.n211 VGND 0.1903f
C6809 Vbias.n212 VGND 0.1262f
C6810 Vbias.t168 VGND 0.1745f
C6811 Vbias.n213 VGND 0.1903f
C6812 Vbias.n214 VGND 0.1262f
C6813 Vbias.t57 VGND 0.1745f
C6814 Vbias.n215 VGND 0.1903f
C6815 Vbias.n216 VGND 0.1262f
C6816 Vbias.t86 VGND 0.1745f
C6817 Vbias.n217 VGND 0.1903f
C6818 Vbias.n218 VGND 0.1262f
C6819 Vbias.t95 VGND 0.1745f
C6820 Vbias.n219 VGND 0.1903f
C6821 Vbias.n220 VGND 0.1262f
C6822 Vbias.t256 VGND 0.1745f
C6823 Vbias.n221 VGND 0.1903f
C6824 Vbias.n222 VGND 0.1262f
C6825 Vbias.n223 VGND 0.54484f
C6826 Vbias.t15 VGND 0.1745f
C6827 Vbias.n224 VGND 0.18997f
C6828 Vbias.t89 VGND 0.1745f
C6829 Vbias.n225 VGND 0.1903f
C6830 Vbias.n226 VGND 0.1262f
C6831 Vbias.t186 VGND 0.1745f
C6832 Vbias.n227 VGND 0.1903f
C6833 Vbias.n228 VGND 0.1262f
C6834 Vbias.t194 VGND 0.1745f
C6835 Vbias.n229 VGND 0.1903f
C6836 Vbias.n230 VGND 0.1262f
C6837 Vbias.t29 VGND 0.1745f
C6838 Vbias.n231 VGND 0.1903f
C6839 Vbias.n232 VGND 0.1262f
C6840 Vbias.t113 VGND 0.1745f
C6841 Vbias.n233 VGND 0.1903f
C6842 Vbias.n234 VGND 0.1262f
C6843 Vbias.t198 VGND 0.1745f
C6844 Vbias.n235 VGND 0.1903f
C6845 Vbias.n236 VGND 0.1262f
C6846 Vbias.t34 VGND 0.1745f
C6847 Vbias.n237 VGND 0.1903f
C6848 Vbias.n238 VGND 0.1262f
C6849 Vbias.t51 VGND 0.1745f
C6850 Vbias.n239 VGND 0.1903f
C6851 Vbias.n240 VGND 0.1262f
C6852 Vbias.t125 VGND 0.1745f
C6853 Vbias.n241 VGND 0.1903f
C6854 Vbias.n242 VGND 0.1262f
C6855 Vbias.t217 VGND 0.1745f
C6856 Vbias.n243 VGND 0.1903f
C6857 Vbias.n244 VGND 0.1262f
C6858 Vbias.t239 VGND 0.1745f
C6859 Vbias.n245 VGND 0.1903f
C6860 Vbias.n246 VGND 0.1262f
C6861 Vbias.t129 VGND 0.1745f
C6862 Vbias.n247 VGND 0.1903f
C6863 Vbias.n248 VGND 0.1262f
C6864 Vbias.t155 VGND 0.1745f
C6865 Vbias.n249 VGND 0.1903f
C6866 Vbias.n250 VGND 0.1262f
C6867 Vbias.t167 VGND 0.1745f
C6868 Vbias.n251 VGND 0.1903f
C6869 Vbias.n252 VGND 0.1262f
C6870 Vbias.t70 VGND 0.1745f
C6871 Vbias.n253 VGND 0.1903f
C6872 Vbias.n254 VGND 0.1262f
C6873 Vbias.n255 VGND 0.54484f
C6874 Vbias.t88 VGND 0.1745f
C6875 Vbias.n256 VGND 0.18997f
C6876 Vbias.t160 VGND 0.1745f
C6877 Vbias.n257 VGND 0.1903f
C6878 Vbias.n258 VGND 0.1262f
C6879 Vbias.t263 VGND 0.1745f
C6880 Vbias.n259 VGND 0.1903f
C6881 Vbias.n260 VGND 0.1262f
C6882 Vbias.t14 VGND 0.1745f
C6883 Vbias.n261 VGND 0.1903f
C6884 Vbias.n262 VGND 0.1262f
C6885 Vbias.t99 VGND 0.1745f
C6886 Vbias.n263 VGND 0.1903f
C6887 Vbias.n264 VGND 0.1262f
C6888 Vbias.t185 VGND 0.1745f
C6889 Vbias.n265 VGND 0.1903f
C6890 Vbias.n266 VGND 0.1262f
C6891 Vbias.t17 VGND 0.1745f
C6892 Vbias.n267 VGND 0.1903f
C6893 Vbias.n268 VGND 0.1262f
C6894 Vbias.t104 VGND 0.1745f
C6895 Vbias.n269 VGND 0.1903f
C6896 Vbias.n270 VGND 0.1262f
C6897 Vbias.t124 VGND 0.1745f
C6898 Vbias.n271 VGND 0.1903f
C6899 Vbias.n272 VGND 0.1262f
C6900 Vbias.t196 VGND 0.1745f
C6901 Vbias.n273 VGND 0.1903f
C6902 Vbias.n274 VGND 0.1262f
C6903 Vbias.t33 VGND 0.1745f
C6904 Vbias.n275 VGND 0.1903f
C6905 Vbias.n276 VGND 0.1262f
C6906 Vbias.t50 VGND 0.1745f
C6907 Vbias.n277 VGND 0.1903f
C6908 Vbias.n278 VGND 0.1262f
C6909 Vbias.t203 VGND 0.1745f
C6910 Vbias.n279 VGND 0.1903f
C6911 Vbias.n280 VGND 0.1262f
C6912 Vbias.t226 VGND 0.1745f
C6913 Vbias.n281 VGND 0.1903f
C6914 Vbias.n282 VGND 0.1262f
C6915 Vbias.t238 VGND 0.1745f
C6916 Vbias.n283 VGND 0.1903f
C6917 Vbias.n284 VGND 0.1262f
C6918 Vbias.t143 VGND 0.1745f
C6919 Vbias.n285 VGND 0.1903f
C6920 Vbias.n286 VGND 0.1262f
C6921 Vbias.n287 VGND 0.54484f
C6922 Vbias.t55 VGND 0.1745f
C6923 Vbias.n288 VGND 0.18997f
C6924 Vbias.t128 VGND 0.1745f
C6925 Vbias.n289 VGND 0.1903f
C6926 Vbias.n290 VGND 0.1262f
C6927 Vbias.t228 VGND 0.1745f
C6928 Vbias.n291 VGND 0.1903f
C6929 Vbias.n292 VGND 0.1262f
C6930 Vbias.t241 VGND 0.1745f
C6931 Vbias.n293 VGND 0.1903f
C6932 Vbias.n294 VGND 0.1262f
C6933 Vbias.t69 VGND 0.1745f
C6934 Vbias.n295 VGND 0.1903f
C6935 Vbias.n296 VGND 0.1262f
C6936 Vbias.t156 VGND 0.1745f
C6937 Vbias.n297 VGND 0.1903f
C6938 Vbias.n298 VGND 0.1262f
C6939 Vbias.t243 VGND 0.1745f
C6940 Vbias.n299 VGND 0.1903f
C6941 Vbias.n300 VGND 0.1262f
C6942 Vbias.t74 VGND 0.1745f
C6943 Vbias.n301 VGND 0.1903f
C6944 Vbias.n302 VGND 0.1262f
C6945 Vbias.t97 VGND 0.1745f
C6946 Vbias.n303 VGND 0.1903f
C6947 Vbias.n304 VGND 0.1262f
C6948 Vbias.t170 VGND 0.1745f
C6949 Vbias.n305 VGND 0.1903f
C6950 Vbias.n306 VGND 0.1262f
C6951 Vbias.t257 VGND 0.1745f
C6952 Vbias.n307 VGND 0.1903f
C6953 Vbias.n308 VGND 0.1262f
C6954 Vbias.t27 VGND 0.1745f
C6955 Vbias.n309 VGND 0.1903f
C6956 Vbias.n310 VGND 0.1262f
C6957 Vbias.t174 VGND 0.1745f
C6958 Vbias.n311 VGND 0.1903f
C6959 Vbias.n312 VGND 0.1262f
C6960 Vbias.t193 VGND 0.1745f
C6961 Vbias.n313 VGND 0.1903f
C6962 Vbias.n314 VGND 0.1262f
C6963 Vbias.t210 VGND 0.1745f
C6964 Vbias.n315 VGND 0.1903f
C6965 Vbias.n316 VGND 0.1262f
C6966 Vbias.t111 VGND 0.1745f
C6967 Vbias.n317 VGND 0.1903f
C6968 Vbias.n318 VGND 0.1262f
C6969 Vbias.n319 VGND 0.54484f
C6970 Vbias.t127 VGND 0.1745f
C6971 Vbias.n320 VGND 0.18997f
C6972 Vbias.t201 VGND 0.1745f
C6973 Vbias.n321 VGND 0.1903f
C6974 Vbias.n322 VGND 0.1262f
C6975 Vbias.t43 VGND 0.1745f
C6976 Vbias.n323 VGND 0.1903f
C6977 Vbias.n324 VGND 0.1262f
C6978 Vbias.t54 VGND 0.1745f
C6979 Vbias.n325 VGND 0.1903f
C6980 Vbias.n326 VGND 0.1262f
C6981 Vbias.t141 VGND 0.1745f
C6982 Vbias.n327 VGND 0.1903f
C6983 Vbias.n328 VGND 0.1262f
C6984 Vbias.t227 VGND 0.1745f
C6985 Vbias.n329 VGND 0.1903f
C6986 Vbias.n330 VGND 0.1262f
C6987 Vbias.t56 VGND 0.1745f
C6988 Vbias.n331 VGND 0.1903f
C6989 Vbias.n332 VGND 0.1262f
C6990 Vbias.t144 VGND 0.1745f
C6991 Vbias.n333 VGND 0.1903f
C6992 Vbias.n334 VGND 0.1262f
C6993 Vbias.t169 VGND 0.1745f
C6994 Vbias.n335 VGND 0.1903f
C6995 Vbias.n336 VGND 0.1262f
C6996 Vbias.t242 VGND 0.1745f
C6997 Vbias.n337 VGND 0.1903f
C6998 Vbias.n338 VGND 0.1262f
C6999 Vbias.t71 VGND 0.1745f
C7000 Vbias.n339 VGND 0.1903f
C7001 Vbias.n340 VGND 0.1262f
C7002 Vbias.t96 VGND 0.1745f
C7003 Vbias.n341 VGND 0.1903f
C7004 Vbias.n342 VGND 0.1262f
C7005 Vbias.t249 VGND 0.1745f
C7006 Vbias.n343 VGND 0.1903f
C7007 Vbias.n344 VGND 0.1262f
C7008 Vbias.t13 VGND 0.1745f
C7009 Vbias.n345 VGND 0.1903f
C7010 Vbias.n346 VGND 0.1262f
C7011 Vbias.t26 VGND 0.1745f
C7012 Vbias.n347 VGND 0.1903f
C7013 Vbias.n348 VGND 0.1262f
C7014 Vbias.t182 VGND 0.1745f
C7015 Vbias.n349 VGND 0.1903f
C7016 Vbias.n350 VGND 0.1262f
C7017 Vbias.n351 VGND 0.54484f
C7018 Vbias.t204 VGND 0.1745f
C7019 Vbias.n352 VGND 0.18997f
C7020 Vbias.t23 VGND 0.1745f
C7021 Vbias.n353 VGND 0.1903f
C7022 Vbias.n354 VGND 0.1262f
C7023 Vbias.t119 VGND 0.1745f
C7024 Vbias.n355 VGND 0.1903f
C7025 Vbias.n356 VGND 0.1262f
C7026 Vbias.t130 VGND 0.1745f
C7027 Vbias.n357 VGND 0.1903f
C7028 Vbias.n358 VGND 0.1262f
C7029 Vbias.t219 VGND 0.1745f
C7030 Vbias.n359 VGND 0.1903f
C7031 Vbias.n360 VGND 0.1262f
C7032 Vbias.t46 VGND 0.1745f
C7033 Vbias.n361 VGND 0.1903f
C7034 Vbias.n362 VGND 0.1262f
C7035 Vbias.t133 VGND 0.1745f
C7036 Vbias.n363 VGND 0.1903f
C7037 Vbias.n364 VGND 0.1262f
C7038 Vbias.t225 VGND 0.1745f
C7039 Vbias.n365 VGND 0.1903f
C7040 Vbias.n366 VGND 0.1262f
C7041 Vbias.t246 VGND 0.1745f
C7042 Vbias.n367 VGND 0.1903f
C7043 Vbias.n368 VGND 0.1262f
C7044 Vbias.t60 VGND 0.1745f
C7045 Vbias.n369 VGND 0.1903f
C7046 Vbias.n370 VGND 0.1262f
C7047 Vbias.t150 VGND 0.1745f
C7048 Vbias.n371 VGND 0.1903f
C7049 Vbias.n372 VGND 0.1262f
C7050 Vbias.t172 VGND 0.1745f
C7051 Vbias.n373 VGND 0.1903f
C7052 Vbias.n374 VGND 0.1262f
C7053 Vbias.t68 VGND 0.1745f
C7054 Vbias.n375 VGND 0.1903f
C7055 Vbias.n376 VGND 0.1262f
C7056 Vbias.t87 VGND 0.1745f
C7057 Vbias.n377 VGND 0.1903f
C7058 Vbias.n378 VGND 0.1262f
C7059 Vbias.t98 VGND 0.1745f
C7060 Vbias.n379 VGND 0.1903f
C7061 Vbias.n380 VGND 0.1262f
C7062 Vbias.t261 VGND 0.1745f
C7063 Vbias.n381 VGND 0.1903f
C7064 Vbias.n382 VGND 0.1262f
C7065 Vbias.n383 VGND 0.54484f
C7066 Vbias.t22 VGND 0.1745f
C7067 Vbias.n384 VGND 0.18997f
C7068 Vbias.t94 VGND 0.1745f
C7069 Vbias.n385 VGND 0.1903f
C7070 Vbias.n386 VGND 0.1262f
C7071 Vbias.t191 VGND 0.1745f
C7072 Vbias.n387 VGND 0.1903f
C7073 Vbias.n388 VGND 0.1262f
C7074 Vbias.t202 VGND 0.1745f
C7075 Vbias.n389 VGND 0.1903f
C7076 Vbias.n390 VGND 0.1262f
C7077 Vbias.t35 VGND 0.1745f
C7078 Vbias.n391 VGND 0.1903f
C7079 Vbias.n392 VGND 0.1262f
C7080 Vbias.t118 VGND 0.1745f
C7081 Vbias.n393 VGND 0.1903f
C7082 Vbias.n394 VGND 0.1262f
C7083 Vbias.t206 VGND 0.1745f
C7084 Vbias.n395 VGND 0.1903f
C7085 Vbias.n396 VGND 0.1262f
C7086 Vbias.t39 VGND 0.1745f
C7087 Vbias.n397 VGND 0.1903f
C7088 Vbias.n398 VGND 0.1262f
C7089 Vbias.t59 VGND 0.1745f
C7090 Vbias.n399 VGND 0.1903f
C7091 Vbias.n400 VGND 0.1262f
C7092 Vbias.t132 VGND 0.1745f
C7093 Vbias.n401 VGND 0.1903f
C7094 Vbias.n402 VGND 0.1262f
C7095 Vbias.t223 VGND 0.1745f
C7096 Vbias.n403 VGND 0.1903f
C7097 Vbias.n404 VGND 0.1262f
C7098 Vbias.t245 VGND 0.1745f
C7099 Vbias.n405 VGND 0.1903f
C7100 Vbias.n406 VGND 0.1262f
C7101 Vbias.t139 VGND 0.1745f
C7102 Vbias.n407 VGND 0.1903f
C7103 Vbias.n408 VGND 0.1262f
C7104 Vbias.t159 VGND 0.1745f
C7105 Vbias.n409 VGND 0.1903f
C7106 Vbias.n410 VGND 0.1262f
C7107 Vbias.t171 VGND 0.1745f
C7108 Vbias.n411 VGND 0.1903f
C7109 Vbias.n412 VGND 0.1262f
C7110 Vbias.t79 VGND 0.1745f
C7111 Vbias.n413 VGND 0.1903f
C7112 Vbias.n414 VGND 0.1262f
C7113 Vbias.n415 VGND 0.54484f
C7114 Vbias.t93 VGND 0.1745f
C7115 Vbias.n416 VGND 0.18997f
C7116 Vbias.t166 VGND 0.1745f
C7117 Vbias.n417 VGND 0.1903f
C7118 Vbias.n418 VGND 0.1262f
C7119 Vbias.t267 VGND 0.1745f
C7120 Vbias.n419 VGND 0.1903f
C7121 Vbias.n420 VGND 0.1262f
C7122 Vbias.t20 VGND 0.1745f
C7123 Vbias.n421 VGND 0.1903f
C7124 Vbias.n422 VGND 0.1262f
C7125 Vbias.t105 VGND 0.1745f
C7126 Vbias.n423 VGND 0.1903f
C7127 Vbias.n424 VGND 0.1262f
C7128 Vbias.t189 VGND 0.1745f
C7129 Vbias.n425 VGND 0.1903f
C7130 Vbias.n426 VGND 0.1262f
C7131 Vbias.t24 VGND 0.1745f
C7132 Vbias.n427 VGND 0.1903f
C7133 Vbias.n428 VGND 0.1262f
C7134 Vbias.t108 VGND 0.1745f
C7135 Vbias.n429 VGND 0.1903f
C7136 Vbias.n430 VGND 0.1262f
C7137 Vbias.t131 VGND 0.1745f
C7138 Vbias.n431 VGND 0.1903f
C7139 Vbias.n432 VGND 0.1262f
C7140 Vbias.t205 VGND 0.1745f
C7141 Vbias.n433 VGND 0.1903f
C7142 Vbias.n434 VGND 0.1262f
C7143 Vbias.t38 VGND 0.1745f
C7144 Vbias.n435 VGND 0.1903f
C7145 Vbias.n436 VGND 0.1262f
C7146 Vbias.t58 VGND 0.1745f
C7147 Vbias.n437 VGND 0.1903f
C7148 Vbias.n438 VGND 0.1262f
C7149 Vbias.t211 VGND 0.1745f
C7150 Vbias.n439 VGND 0.1903f
C7151 Vbias.n440 VGND 0.1262f
C7152 Vbias.t231 VGND 0.1745f
C7153 Vbias.n441 VGND 0.1903f
C7154 Vbias.n442 VGND 0.1262f
C7155 Vbias.t244 VGND 0.1745f
C7156 Vbias.n443 VGND 0.1903f
C7157 Vbias.n444 VGND 0.1262f
C7158 Vbias.t152 VGND 0.1745f
C7159 Vbias.n445 VGND 0.1903f
C7160 Vbias.n446 VGND 0.1262f
C7161 Vbias.n447 VGND 0.54484f
C7162 Vbias.t63 VGND 0.1745f
C7163 Vbias.n448 VGND 0.18997f
C7164 Vbias.t136 VGND 0.1745f
C7165 Vbias.n449 VGND 0.1903f
C7166 Vbias.n450 VGND 0.1262f
C7167 Vbias.t235 VGND 0.1745f
C7168 Vbias.n451 VGND 0.1903f
C7169 Vbias.n452 VGND 0.1262f
C7170 Vbias.t248 VGND 0.1745f
C7171 Vbias.n453 VGND 0.1903f
C7172 Vbias.n454 VGND 0.1262f
C7173 Vbias.t75 VGND 0.1745f
C7174 Vbias.n455 VGND 0.1903f
C7175 Vbias.n456 VGND 0.1262f
C7176 Vbias.t162 VGND 0.1745f
C7177 Vbias.n457 VGND 0.1903f
C7178 Vbias.n458 VGND 0.1262f
C7179 Vbias.t253 VGND 0.1745f
C7180 Vbias.n459 VGND 0.1903f
C7181 Vbias.n460 VGND 0.1262f
C7182 Vbias.t82 VGND 0.1745f
C7183 Vbias.n461 VGND 0.1903f
C7184 Vbias.n462 VGND 0.1262f
C7185 Vbias.t102 VGND 0.1745f
C7186 Vbias.n463 VGND 0.1903f
C7187 Vbias.n464 VGND 0.1262f
C7188 Vbias.t177 VGND 0.1745f
C7189 Vbias.n465 VGND 0.1903f
C7190 Vbias.n466 VGND 0.1262f
C7191 Vbias.t264 VGND 0.1745f
C7192 Vbias.n467 VGND 0.1903f
C7193 Vbias.n468 VGND 0.1262f
C7194 Vbias.t31 VGND 0.1745f
C7195 Vbias.n469 VGND 0.1903f
C7196 Vbias.n470 VGND 0.1262f
C7197 Vbias.t179 VGND 0.1745f
C7198 Vbias.n471 VGND 0.1903f
C7199 Vbias.n472 VGND 0.1262f
C7200 Vbias.t199 VGND 0.1745f
C7201 Vbias.n473 VGND 0.1903f
C7202 Vbias.n474 VGND 0.1262f
C7203 Vbias.t216 VGND 0.1745f
C7204 Vbias.n475 VGND 0.1903f
C7205 Vbias.n476 VGND 0.1262f
C7206 Vbias.t116 VGND 0.1745f
C7207 Vbias.n477 VGND 0.1903f
C7208 Vbias.n478 VGND 0.1262f
C7209 Vbias.n479 VGND 0.54484f
C7210 Vbias.t135 VGND 0.1745f
C7211 Vbias.n480 VGND 0.18997f
C7212 Vbias.t207 VGND 0.1745f
C7213 Vbias.n481 VGND 0.1903f
C7214 Vbias.n482 VGND 0.1262f
C7215 Vbias.t47 VGND 0.1745f
C7216 Vbias.n483 VGND 0.1903f
C7217 Vbias.n484 VGND 0.1262f
C7218 Vbias.t62 VGND 0.1745f
C7219 Vbias.n485 VGND 0.1903f
C7220 Vbias.n486 VGND 0.1262f
C7221 Vbias.t147 VGND 0.1745f
C7222 Vbias.n487 VGND 0.1903f
C7223 Vbias.n488 VGND 0.1262f
C7224 Vbias.t233 VGND 0.1745f
C7225 Vbias.n489 VGND 0.1903f
C7226 Vbias.n490 VGND 0.1262f
C7227 Vbias.t66 VGND 0.1745f
C7228 Vbias.n491 VGND 0.1903f
C7229 Vbias.n492 VGND 0.1262f
C7230 Vbias.t153 VGND 0.1745f
C7231 Vbias.n493 VGND 0.1903f
C7232 Vbias.n494 VGND 0.1262f
C7233 Vbias.t175 VGND 0.1745f
C7234 Vbias.n495 VGND 0.1903f
C7235 Vbias.n496 VGND 0.1262f
C7236 Vbias.t252 VGND 0.1745f
C7237 Vbias.n497 VGND 0.1903f
C7238 Vbias.n498 VGND 0.1262f
C7239 Vbias.t81 VGND 0.1745f
C7240 Vbias.n499 VGND 0.1903f
C7241 Vbias.n500 VGND 0.1262f
C7242 Vbias.t101 VGND 0.1745f
C7243 Vbias.n501 VGND 0.1903f
C7244 Vbias.n502 VGND 0.1262f
C7245 Vbias.t254 VGND 0.1745f
C7246 Vbias.n503 VGND 0.1903f
C7247 Vbias.n504 VGND 0.1262f
C7248 Vbias.t18 VGND 0.1745f
C7249 Vbias.n505 VGND 0.1903f
C7250 Vbias.n506 VGND 0.1262f
C7251 Vbias.t30 VGND 0.1745f
C7252 Vbias.n507 VGND 0.1903f
C7253 Vbias.n508 VGND 0.1262f
C7254 Vbias.t187 VGND 0.1745f
C7255 Vbias.n509 VGND 0.1903f
C7256 Vbias.n510 VGND 0.1262f
C7257 Vbias.n511 VGND 0.63367f
C7258 Vbias.t5 VGND 0.17357f
C7259 Vbias.n512 VGND 0.58869f
C7260 Vbias.t9 VGND 0.02547f
C7261 Vbias.t0 VGND 0.02547f
C7262 Vbias.n513 VGND 0.05413f
C7263 Vbias.t2 VGND 0.01606f
C7264 Vbias.t8 VGND 0.01606f
C7265 Vbias.n514 VGND 0.03416f
C7266 Vbias.n515 VGND 2.28043f
C7267 Vbias.t4 VGND 0.33466f
C7268 Vbias.n516 VGND 0.38359f
C7269 Vbias.n517 VGND 0.21155f
C7270 Vbias.t7 VGND 0.17357f
C7271 Vbias.n518 VGND 0.54497f
C7272 Vbias.t3 VGND 0.02547f
C7273 Vbias.t11 VGND 0.02547f
C7274 Vbias.n519 VGND 0.05413f
C7275 Vbias.t1 VGND 0.01606f
C7276 Vbias.t10 VGND 0.01606f
C7277 Vbias.n520 VGND 0.03416f
C7278 Vbias.n521 VGND 2.28043f
C7279 Vbias.t6 VGND 0.33461f
C7280 Vbias.n522 VGND 0.38359f
C7281 Vbias.n523 VGND 0.19521f
C7282 Vbias.n524 VGND 1.81716f
C7283 XThC.Tn[2].t7 VGND 0.01169f
C7284 XThC.Tn[2].t6 VGND 0.01169f
C7285 XThC.Tn[2].n0 VGND 0.02361f
C7286 XThC.Tn[2].t5 VGND 0.01169f
C7287 XThC.Tn[2].t4 VGND 0.01169f
C7288 XThC.Tn[2].n1 VGND 0.02762f
C7289 XThC.Tn[2].n2 VGND 0.07732f
C7290 XThC.Tn[2].n3 VGND 0.01731f
C7291 XThC.Tn[2].n4 VGND 0.01731f
C7292 XThC.Tn[2].n5 VGND 0.01731f
C7293 XThC.Tn[2].n6 VGND 0.02884f
C7294 XThC.Tn[2].n7 VGND 0.08243f
C7295 XThC.Tn[2].n8 VGND 0.05096f
C7296 XThC.Tn[2].n9 VGND 0.05751f
C7297 XThC.Tn[2].t18 VGND 0.01012f
C7298 XThC.Tn[2].n10 VGND 0.02261f
C7299 XThC.Tn[2].n11 VGND 0.01292f
C7300 XThC.Tn[2].n12 VGND 0.01571f
C7301 XThC.Tn[2].t35 VGND 0.01012f
C7302 XThC.Tn[2].n13 VGND 0.02261f
C7303 XThC.Tn[2].n14 VGND 0.01292f
C7304 XThC.Tn[2].n15 VGND 0.07465f
C7305 XThC.Tn[2].t37 VGND 0.01012f
C7306 XThC.Tn[2].n16 VGND 0.02261f
C7307 XThC.Tn[2].n17 VGND 0.01292f
C7308 XThC.Tn[2].n18 VGND 0.07465f
C7309 XThC.Tn[2].t39 VGND 0.01012f
C7310 XThC.Tn[2].n19 VGND 0.02261f
C7311 XThC.Tn[2].n20 VGND 0.01292f
C7312 XThC.Tn[2].n21 VGND 0.07465f
C7313 XThC.Tn[2].t28 VGND 0.01012f
C7314 XThC.Tn[2].n22 VGND 0.02261f
C7315 XThC.Tn[2].n23 VGND 0.01292f
C7316 XThC.Tn[2].n24 VGND 0.07465f
C7317 XThC.Tn[2].t29 VGND 0.01012f
C7318 XThC.Tn[2].n25 VGND 0.02261f
C7319 XThC.Tn[2].n26 VGND 0.01292f
C7320 XThC.Tn[2].n27 VGND 0.07465f
C7321 XThC.Tn[2].t42 VGND 0.01012f
C7322 XThC.Tn[2].n28 VGND 0.02261f
C7323 XThC.Tn[2].n29 VGND 0.01292f
C7324 XThC.Tn[2].n30 VGND 0.07465f
C7325 XThC.Tn[2].t19 VGND 0.01012f
C7326 XThC.Tn[2].n31 VGND 0.02261f
C7327 XThC.Tn[2].n32 VGND 0.01292f
C7328 XThC.Tn[2].n33 VGND 0.07465f
C7329 XThC.Tn[2].t21 VGND 0.01012f
C7330 XThC.Tn[2].n34 VGND 0.02261f
C7331 XThC.Tn[2].n35 VGND 0.01292f
C7332 XThC.Tn[2].n36 VGND 0.07465f
C7333 XThC.Tn[2].t40 VGND 0.01012f
C7334 XThC.Tn[2].n37 VGND 0.02261f
C7335 XThC.Tn[2].n38 VGND 0.01292f
C7336 XThC.Tn[2].n39 VGND 0.07465f
C7337 XThC.Tn[2].t41 VGND 0.01012f
C7338 XThC.Tn[2].n40 VGND 0.02261f
C7339 XThC.Tn[2].n41 VGND 0.01292f
C7340 XThC.Tn[2].n42 VGND 0.07465f
C7341 XThC.Tn[2].t22 VGND 0.01012f
C7342 XThC.Tn[2].n43 VGND 0.02261f
C7343 XThC.Tn[2].n44 VGND 0.01292f
C7344 XThC.Tn[2].n45 VGND 0.07465f
C7345 XThC.Tn[2].t30 VGND 0.01012f
C7346 XThC.Tn[2].n46 VGND 0.02261f
C7347 XThC.Tn[2].n47 VGND 0.01292f
C7348 XThC.Tn[2].n48 VGND 0.07465f
C7349 XThC.Tn[2].t33 VGND 0.01012f
C7350 XThC.Tn[2].n49 VGND 0.02261f
C7351 XThC.Tn[2].n50 VGND 0.01292f
C7352 XThC.Tn[2].n51 VGND 0.07465f
C7353 XThC.Tn[2].t14 VGND 0.01012f
C7354 XThC.Tn[2].n52 VGND 0.02261f
C7355 XThC.Tn[2].n53 VGND 0.01292f
C7356 XThC.Tn[2].n54 VGND 0.07465f
C7357 XThC.Tn[2].t24 VGND 0.01012f
C7358 XThC.Tn[2].n55 VGND 0.02261f
C7359 XThC.Tn[2].n56 VGND 0.01292f
C7360 XThC.Tn[2].n57 VGND 0.07465f
C7361 XThC.Tn[2].n58 VGND 0.27153f
C7362 XThC.Tn[2].n59 VGND 0.0441f
C7363 XThC.Tn[2].n60 VGND 0.02447f
C7364 XThC.Tn[4].t9 VGND 0.01194f
C7365 XThC.Tn[4].t8 VGND 0.01194f
C7366 XThC.Tn[4].n0 VGND 0.02411f
C7367 XThC.Tn[4].t11 VGND 0.01194f
C7368 XThC.Tn[4].t10 VGND 0.01194f
C7369 XThC.Tn[4].n1 VGND 0.02821f
C7370 XThC.Tn[4].n2 VGND 0.07897f
C7371 XThC.Tn[4].n3 VGND 0.01768f
C7372 XThC.Tn[4].n4 VGND 0.01768f
C7373 XThC.Tn[4].n5 VGND 0.01768f
C7374 XThC.Tn[4].n6 VGND 0.02946f
C7375 XThC.Tn[4].n7 VGND 0.0842f
C7376 XThC.Tn[4].n8 VGND 0.05205f
C7377 XThC.Tn[4].n9 VGND 0.05874f
C7378 XThC.Tn[4].t26 VGND 0.01034f
C7379 XThC.Tn[4].n10 VGND 0.02309f
C7380 XThC.Tn[4].n11 VGND 0.0132f
C7381 XThC.Tn[4].n12 VGND 0.01605f
C7382 XThC.Tn[4].t43 VGND 0.01034f
C7383 XThC.Tn[4].n13 VGND 0.02309f
C7384 XThC.Tn[4].n14 VGND 0.0132f
C7385 XThC.Tn[4].n15 VGND 0.07625f
C7386 XThC.Tn[4].t13 VGND 0.01034f
C7387 XThC.Tn[4].n16 VGND 0.02309f
C7388 XThC.Tn[4].n17 VGND 0.0132f
C7389 XThC.Tn[4].n18 VGND 0.07625f
C7390 XThC.Tn[4].t15 VGND 0.01034f
C7391 XThC.Tn[4].n19 VGND 0.02309f
C7392 XThC.Tn[4].n20 VGND 0.0132f
C7393 XThC.Tn[4].n21 VGND 0.07625f
C7394 XThC.Tn[4].t36 VGND 0.01034f
C7395 XThC.Tn[4].n22 VGND 0.02309f
C7396 XThC.Tn[4].n23 VGND 0.0132f
C7397 XThC.Tn[4].n24 VGND 0.07625f
C7398 XThC.Tn[4].t37 VGND 0.01034f
C7399 XThC.Tn[4].n25 VGND 0.02309f
C7400 XThC.Tn[4].n26 VGND 0.0132f
C7401 XThC.Tn[4].n27 VGND 0.07625f
C7402 XThC.Tn[4].t18 VGND 0.01034f
C7403 XThC.Tn[4].n28 VGND 0.02309f
C7404 XThC.Tn[4].n29 VGND 0.0132f
C7405 XThC.Tn[4].n30 VGND 0.07625f
C7406 XThC.Tn[4].t27 VGND 0.01034f
C7407 XThC.Tn[4].n31 VGND 0.02309f
C7408 XThC.Tn[4].n32 VGND 0.0132f
C7409 XThC.Tn[4].n33 VGND 0.07625f
C7410 XThC.Tn[4].t29 VGND 0.01034f
C7411 XThC.Tn[4].n34 VGND 0.02309f
C7412 XThC.Tn[4].n35 VGND 0.0132f
C7413 XThC.Tn[4].n36 VGND 0.07625f
C7414 XThC.Tn[4].t16 VGND 0.01034f
C7415 XThC.Tn[4].n37 VGND 0.02309f
C7416 XThC.Tn[4].n38 VGND 0.0132f
C7417 XThC.Tn[4].n39 VGND 0.07625f
C7418 XThC.Tn[4].t17 VGND 0.01034f
C7419 XThC.Tn[4].n40 VGND 0.02309f
C7420 XThC.Tn[4].n41 VGND 0.0132f
C7421 XThC.Tn[4].n42 VGND 0.07625f
C7422 XThC.Tn[4].t30 VGND 0.01034f
C7423 XThC.Tn[4].n43 VGND 0.02309f
C7424 XThC.Tn[4].n44 VGND 0.0132f
C7425 XThC.Tn[4].n45 VGND 0.07625f
C7426 XThC.Tn[4].t38 VGND 0.01034f
C7427 XThC.Tn[4].n46 VGND 0.02309f
C7428 XThC.Tn[4].n47 VGND 0.0132f
C7429 XThC.Tn[4].n48 VGND 0.07625f
C7430 XThC.Tn[4].t41 VGND 0.01034f
C7431 XThC.Tn[4].n49 VGND 0.02309f
C7432 XThC.Tn[4].n50 VGND 0.0132f
C7433 XThC.Tn[4].n51 VGND 0.07625f
C7434 XThC.Tn[4].t22 VGND 0.01034f
C7435 XThC.Tn[4].n52 VGND 0.02309f
C7436 XThC.Tn[4].n53 VGND 0.0132f
C7437 XThC.Tn[4].n54 VGND 0.07625f
C7438 XThC.Tn[4].t32 VGND 0.01034f
C7439 XThC.Tn[4].n55 VGND 0.02309f
C7440 XThC.Tn[4].n56 VGND 0.0132f
C7441 XThC.Tn[4].n57 VGND 0.07625f
C7442 XThC.Tn[4].n58 VGND 0.23757f
C7443 XThC.Tn[4].n59 VGND 0.04514f
C7444 XThC.Tn[4].n60 VGND 0.025f
C7445 XThR.Tn[5].t6 VGND 0.01808f
C7446 XThR.Tn[5].t7 VGND 0.01808f
C7447 XThR.Tn[5].n0 VGND 0.03649f
C7448 XThR.Tn[5].t5 VGND 0.01808f
C7449 XThR.Tn[5].t4 VGND 0.01808f
C7450 XThR.Tn[5].n1 VGND 0.04269f
C7451 XThR.Tn[5].n2 VGND 0.11952f
C7452 XThR.Tn[5].t11 VGND 0.01175f
C7453 XThR.Tn[5].t8 VGND 0.01175f
C7454 XThR.Tn[5].n3 VGND 0.02676f
C7455 XThR.Tn[5].t10 VGND 0.01175f
C7456 XThR.Tn[5].t9 VGND 0.01175f
C7457 XThR.Tn[5].n4 VGND 0.02676f
C7458 XThR.Tn[5].t0 VGND 0.01175f
C7459 XThR.Tn[5].t1 VGND 0.01175f
C7460 XThR.Tn[5].n5 VGND 0.04459f
C7461 XThR.Tn[5].t3 VGND 0.01175f
C7462 XThR.Tn[5].t2 VGND 0.01175f
C7463 XThR.Tn[5].n6 VGND 0.02676f
C7464 XThR.Tn[5].n7 VGND 0.12743f
C7465 XThR.Tn[5].n8 VGND 0.07877f
C7466 XThR.Tn[5].n9 VGND 0.0889f
C7467 XThR.Tn[5].t17 VGND 0.01413f
C7468 XThR.Tn[5].t72 VGND 0.01547f
C7469 XThR.Tn[5].n10 VGND 0.03778f
C7470 XThR.Tn[5].n11 VGND 0.07257f
C7471 XThR.Tn[5].t39 VGND 0.01413f
C7472 XThR.Tn[5].t26 VGND 0.01547f
C7473 XThR.Tn[5].n12 VGND 0.03778f
C7474 XThR.Tn[5].t13 VGND 0.01408f
C7475 XThR.Tn[5].t23 VGND 0.01542f
C7476 XThR.Tn[5].n13 VGND 0.03931f
C7477 XThR.Tn[5].n14 VGND 0.02761f
C7478 XThR.Tn[5].n16 VGND 0.08862f
C7479 XThR.Tn[5].t73 VGND 0.01413f
C7480 XThR.Tn[5].t66 VGND 0.01547f
C7481 XThR.Tn[5].n17 VGND 0.03778f
C7482 XThR.Tn[5].t48 VGND 0.01408f
C7483 XThR.Tn[5].t61 VGND 0.01542f
C7484 XThR.Tn[5].n18 VGND 0.03931f
C7485 XThR.Tn[5].n19 VGND 0.02761f
C7486 XThR.Tn[5].n21 VGND 0.08862f
C7487 XThR.Tn[5].t28 VGND 0.01413f
C7488 XThR.Tn[5].t21 VGND 0.01547f
C7489 XThR.Tn[5].n22 VGND 0.03778f
C7490 XThR.Tn[5].t65 VGND 0.01408f
C7491 XThR.Tn[5].t18 VGND 0.01542f
C7492 XThR.Tn[5].n23 VGND 0.03931f
C7493 XThR.Tn[5].n24 VGND 0.02761f
C7494 XThR.Tn[5].n26 VGND 0.08862f
C7495 XThR.Tn[5].t55 VGND 0.01413f
C7496 XThR.Tn[5].t51 VGND 0.01547f
C7497 XThR.Tn[5].n27 VGND 0.03778f
C7498 XThR.Tn[5].t33 VGND 0.01408f
C7499 XThR.Tn[5].t46 VGND 0.01542f
C7500 XThR.Tn[5].n28 VGND 0.03931f
C7501 XThR.Tn[5].n29 VGND 0.02761f
C7502 XThR.Tn[5].n31 VGND 0.08862f
C7503 XThR.Tn[5].t30 VGND 0.01413f
C7504 XThR.Tn[5].t22 VGND 0.01547f
C7505 XThR.Tn[5].n32 VGND 0.03778f
C7506 XThR.Tn[5].t67 VGND 0.01408f
C7507 XThR.Tn[5].t19 VGND 0.01542f
C7508 XThR.Tn[5].n33 VGND 0.03931f
C7509 XThR.Tn[5].n34 VGND 0.02761f
C7510 XThR.Tn[5].n36 VGND 0.08862f
C7511 XThR.Tn[5].t69 VGND 0.01413f
C7512 XThR.Tn[5].t40 VGND 0.01547f
C7513 XThR.Tn[5].n37 VGND 0.03778f
C7514 XThR.Tn[5].t43 VGND 0.01408f
C7515 XThR.Tn[5].t37 VGND 0.01542f
C7516 XThR.Tn[5].n38 VGND 0.03931f
C7517 XThR.Tn[5].n39 VGND 0.02761f
C7518 XThR.Tn[5].n41 VGND 0.08862f
C7519 XThR.Tn[5].t38 VGND 0.01413f
C7520 XThR.Tn[5].t32 VGND 0.01547f
C7521 XThR.Tn[5].n42 VGND 0.03778f
C7522 XThR.Tn[5].t14 VGND 0.01408f
C7523 XThR.Tn[5].t29 VGND 0.01542f
C7524 XThR.Tn[5].n43 VGND 0.03931f
C7525 XThR.Tn[5].n44 VGND 0.02761f
C7526 XThR.Tn[5].n46 VGND 0.08862f
C7527 XThR.Tn[5].t42 VGND 0.01413f
C7528 XThR.Tn[5].t49 VGND 0.01547f
C7529 XThR.Tn[5].n47 VGND 0.03778f
C7530 XThR.Tn[5].t16 VGND 0.01408f
C7531 XThR.Tn[5].t45 VGND 0.01542f
C7532 XThR.Tn[5].n48 VGND 0.03931f
C7533 XThR.Tn[5].n49 VGND 0.02761f
C7534 XThR.Tn[5].n51 VGND 0.08862f
C7535 XThR.Tn[5].t58 VGND 0.01413f
C7536 XThR.Tn[5].t68 VGND 0.01547f
C7537 XThR.Tn[5].n52 VGND 0.03778f
C7538 XThR.Tn[5].t36 VGND 0.01408f
C7539 XThR.Tn[5].t63 VGND 0.01542f
C7540 XThR.Tn[5].n53 VGND 0.03931f
C7541 XThR.Tn[5].n54 VGND 0.02761f
C7542 XThR.Tn[5].n56 VGND 0.08862f
C7543 XThR.Tn[5].t53 VGND 0.01413f
C7544 XThR.Tn[5].t24 VGND 0.01547f
C7545 XThR.Tn[5].n57 VGND 0.03778f
C7546 XThR.Tn[5].t25 VGND 0.01408f
C7547 XThR.Tn[5].t20 VGND 0.01542f
C7548 XThR.Tn[5].n58 VGND 0.03931f
C7549 XThR.Tn[5].n59 VGND 0.02761f
C7550 XThR.Tn[5].n61 VGND 0.08862f
C7551 XThR.Tn[5].t71 VGND 0.01413f
C7552 XThR.Tn[5].t60 VGND 0.01547f
C7553 XThR.Tn[5].n62 VGND 0.03778f
C7554 XThR.Tn[5].t44 VGND 0.01408f
C7555 XThR.Tn[5].t57 VGND 0.01542f
C7556 XThR.Tn[5].n63 VGND 0.03931f
C7557 XThR.Tn[5].n64 VGND 0.02761f
C7558 XThR.Tn[5].n66 VGND 0.08862f
C7559 XThR.Tn[5].t41 VGND 0.01413f
C7560 XThR.Tn[5].t35 VGND 0.01547f
C7561 XThR.Tn[5].n67 VGND 0.03778f
C7562 XThR.Tn[5].t15 VGND 0.01408f
C7563 XThR.Tn[5].t31 VGND 0.01542f
C7564 XThR.Tn[5].n68 VGND 0.03931f
C7565 XThR.Tn[5].n69 VGND 0.02761f
C7566 XThR.Tn[5].n71 VGND 0.08862f
C7567 XThR.Tn[5].t56 VGND 0.01413f
C7568 XThR.Tn[5].t52 VGND 0.01547f
C7569 XThR.Tn[5].n72 VGND 0.03778f
C7570 XThR.Tn[5].t34 VGND 0.01408f
C7571 XThR.Tn[5].t47 VGND 0.01542f
C7572 XThR.Tn[5].n73 VGND 0.03931f
C7573 XThR.Tn[5].n74 VGND 0.02761f
C7574 XThR.Tn[5].n76 VGND 0.08862f
C7575 XThR.Tn[5].t12 VGND 0.01413f
C7576 XThR.Tn[5].t70 VGND 0.01547f
C7577 XThR.Tn[5].n77 VGND 0.03778f
C7578 XThR.Tn[5].t50 VGND 0.01408f
C7579 XThR.Tn[5].t64 VGND 0.01542f
C7580 XThR.Tn[5].n78 VGND 0.03931f
C7581 XThR.Tn[5].n79 VGND 0.02761f
C7582 XThR.Tn[5].n81 VGND 0.08862f
C7583 XThR.Tn[5].t54 VGND 0.01413f
C7584 XThR.Tn[5].t62 VGND 0.01547f
C7585 XThR.Tn[5].n82 VGND 0.03778f
C7586 XThR.Tn[5].t27 VGND 0.01408f
C7587 XThR.Tn[5].t59 VGND 0.01542f
C7588 XThR.Tn[5].n83 VGND 0.03931f
C7589 XThR.Tn[5].n84 VGND 0.02761f
C7590 XThR.Tn[5].n86 VGND 0.08862f
C7591 XThR.Tn[5].n87 VGND 0.08053f
C7592 XThR.Tn[5].n88 VGND 0.15597f
C7593 XThR.Tn[5].n89 VGND 0.03783f
C7594 XThR.Tn[3].t9 VGND 0.01821f
C7595 XThR.Tn[3].t10 VGND 0.01821f
C7596 XThR.Tn[3].n0 VGND 0.03675f
C7597 XThR.Tn[3].t8 VGND 0.01821f
C7598 XThR.Tn[3].t11 VGND 0.01821f
C7599 XThR.Tn[3].n1 VGND 0.043f
C7600 XThR.Tn[3].n2 VGND 0.12037f
C7601 XThR.Tn[3].t7 VGND 0.01183f
C7602 XThR.Tn[3].t4 VGND 0.01183f
C7603 XThR.Tn[3].n3 VGND 0.02695f
C7604 XThR.Tn[3].t6 VGND 0.01183f
C7605 XThR.Tn[3].t5 VGND 0.01183f
C7606 XThR.Tn[3].n4 VGND 0.02695f
C7607 XThR.Tn[3].t0 VGND 0.01183f
C7608 XThR.Tn[3].t1 VGND 0.01183f
C7609 XThR.Tn[3].n5 VGND 0.0449f
C7610 XThR.Tn[3].t3 VGND 0.01183f
C7611 XThR.Tn[3].t2 VGND 0.01183f
C7612 XThR.Tn[3].n6 VGND 0.02695f
C7613 XThR.Tn[3].n7 VGND 0.12834f
C7614 XThR.Tn[3].n8 VGND 0.07933f
C7615 XThR.Tn[3].n9 VGND 0.08953f
C7616 XThR.Tn[3].t64 VGND 0.01423f
C7617 XThR.Tn[3].t57 VGND 0.01558f
C7618 XThR.Tn[3].n10 VGND 0.03805f
C7619 XThR.Tn[3].n11 VGND 0.07309f
C7620 XThR.Tn[3].t18 VGND 0.01423f
C7621 XThR.Tn[3].t70 VGND 0.01558f
C7622 XThR.Tn[3].n12 VGND 0.03805f
C7623 XThR.Tn[3].t24 VGND 0.01418f
C7624 XThR.Tn[3].t55 VGND 0.01553f
C7625 XThR.Tn[3].n13 VGND 0.03959f
C7626 XThR.Tn[3].n14 VGND 0.02781f
C7627 XThR.Tn[3].n16 VGND 0.08925f
C7628 XThR.Tn[3].t59 VGND 0.01423f
C7629 XThR.Tn[3].t49 VGND 0.01558f
C7630 XThR.Tn[3].n17 VGND 0.03805f
C7631 XThR.Tn[3].t62 VGND 0.01418f
C7632 XThR.Tn[3].t29 VGND 0.01553f
C7633 XThR.Tn[3].n18 VGND 0.03959f
C7634 XThR.Tn[3].n19 VGND 0.02781f
C7635 XThR.Tn[3].n21 VGND 0.08925f
C7636 XThR.Tn[3].t71 VGND 0.01423f
C7637 XThR.Tn[3].t67 VGND 0.01558f
C7638 XThR.Tn[3].n22 VGND 0.03805f
C7639 XThR.Tn[3].t12 VGND 0.01418f
C7640 XThR.Tn[3].t47 VGND 0.01553f
C7641 XThR.Tn[3].n23 VGND 0.03959f
C7642 XThR.Tn[3].n24 VGND 0.02781f
C7643 XThR.Tn[3].n26 VGND 0.08925f
C7644 XThR.Tn[3].t39 VGND 0.01423f
C7645 XThR.Tn[3].t33 VGND 0.01558f
C7646 XThR.Tn[3].n27 VGND 0.03805f
C7647 XThR.Tn[3].t42 VGND 0.01418f
C7648 XThR.Tn[3].t13 VGND 0.01553f
C7649 XThR.Tn[3].n28 VGND 0.03959f
C7650 XThR.Tn[3].n29 VGND 0.02781f
C7651 XThR.Tn[3].n31 VGND 0.08925f
C7652 XThR.Tn[3].t72 VGND 0.01423f
C7653 XThR.Tn[3].t68 VGND 0.01558f
C7654 XThR.Tn[3].n32 VGND 0.03805f
C7655 XThR.Tn[3].t16 VGND 0.01418f
C7656 XThR.Tn[3].t48 VGND 0.01553f
C7657 XThR.Tn[3].n33 VGND 0.03959f
C7658 XThR.Tn[3].n34 VGND 0.02781f
C7659 XThR.Tn[3].n36 VGND 0.08925f
C7660 XThR.Tn[3].t52 VGND 0.01423f
C7661 XThR.Tn[3].t20 VGND 0.01558f
C7662 XThR.Tn[3].n37 VGND 0.03805f
C7663 XThR.Tn[3].t56 VGND 0.01418f
C7664 XThR.Tn[3].t66 VGND 0.01553f
C7665 XThR.Tn[3].n38 VGND 0.03959f
C7666 XThR.Tn[3].n39 VGND 0.02781f
C7667 XThR.Tn[3].n41 VGND 0.08925f
C7668 XThR.Tn[3].t19 VGND 0.01423f
C7669 XThR.Tn[3].t14 VGND 0.01558f
C7670 XThR.Tn[3].n42 VGND 0.03805f
C7671 XThR.Tn[3].t23 VGND 0.01418f
C7672 XThR.Tn[3].t61 VGND 0.01553f
C7673 XThR.Tn[3].n43 VGND 0.03959f
C7674 XThR.Tn[3].n44 VGND 0.02781f
C7675 XThR.Tn[3].n46 VGND 0.08925f
C7676 XThR.Tn[3].t22 VGND 0.01423f
C7677 XThR.Tn[3].t31 VGND 0.01558f
C7678 XThR.Tn[3].n47 VGND 0.03805f
C7679 XThR.Tn[3].t28 VGND 0.01418f
C7680 XThR.Tn[3].t73 VGND 0.01553f
C7681 XThR.Tn[3].n48 VGND 0.03959f
C7682 XThR.Tn[3].n49 VGND 0.02781f
C7683 XThR.Tn[3].n51 VGND 0.08925f
C7684 XThR.Tn[3].t41 VGND 0.01423f
C7685 XThR.Tn[3].t51 VGND 0.01558f
C7686 XThR.Tn[3].n52 VGND 0.03805f
C7687 XThR.Tn[3].t45 VGND 0.01418f
C7688 XThR.Tn[3].t30 VGND 0.01553f
C7689 XThR.Tn[3].n53 VGND 0.03959f
C7690 XThR.Tn[3].n54 VGND 0.02781f
C7691 XThR.Tn[3].n56 VGND 0.08925f
C7692 XThR.Tn[3].t35 VGND 0.01423f
C7693 XThR.Tn[3].t69 VGND 0.01558f
C7694 XThR.Tn[3].n57 VGND 0.03805f
C7695 XThR.Tn[3].t37 VGND 0.01418f
C7696 XThR.Tn[3].t50 VGND 0.01553f
C7697 XThR.Tn[3].n58 VGND 0.03959f
C7698 XThR.Tn[3].n59 VGND 0.02781f
C7699 XThR.Tn[3].n61 VGND 0.08925f
C7700 XThR.Tn[3].t54 VGND 0.01423f
C7701 XThR.Tn[3].t44 VGND 0.01558f
C7702 XThR.Tn[3].n62 VGND 0.03805f
C7703 XThR.Tn[3].t58 VGND 0.01418f
C7704 XThR.Tn[3].t25 VGND 0.01553f
C7705 XThR.Tn[3].n63 VGND 0.03959f
C7706 XThR.Tn[3].n64 VGND 0.02781f
C7707 XThR.Tn[3].n66 VGND 0.08925f
C7708 XThR.Tn[3].t21 VGND 0.01423f
C7709 XThR.Tn[3].t17 VGND 0.01558f
C7710 XThR.Tn[3].n67 VGND 0.03805f
C7711 XThR.Tn[3].t26 VGND 0.01418f
C7712 XThR.Tn[3].t63 VGND 0.01553f
C7713 XThR.Tn[3].n68 VGND 0.03959f
C7714 XThR.Tn[3].n69 VGND 0.02781f
C7715 XThR.Tn[3].n71 VGND 0.08925f
C7716 XThR.Tn[3].t40 VGND 0.01423f
C7717 XThR.Tn[3].t34 VGND 0.01558f
C7718 XThR.Tn[3].n72 VGND 0.03805f
C7719 XThR.Tn[3].t43 VGND 0.01418f
C7720 XThR.Tn[3].t15 VGND 0.01553f
C7721 XThR.Tn[3].n73 VGND 0.03959f
C7722 XThR.Tn[3].n74 VGND 0.02781f
C7723 XThR.Tn[3].n76 VGND 0.08925f
C7724 XThR.Tn[3].t60 VGND 0.01423f
C7725 XThR.Tn[3].t53 VGND 0.01558f
C7726 XThR.Tn[3].n77 VGND 0.03805f
C7727 XThR.Tn[3].t65 VGND 0.01418f
C7728 XThR.Tn[3].t32 VGND 0.01553f
C7729 XThR.Tn[3].n78 VGND 0.03959f
C7730 XThR.Tn[3].n79 VGND 0.02781f
C7731 XThR.Tn[3].n81 VGND 0.08925f
C7732 XThR.Tn[3].t36 VGND 0.01423f
C7733 XThR.Tn[3].t46 VGND 0.01558f
C7734 XThR.Tn[3].n82 VGND 0.03805f
C7735 XThR.Tn[3].t38 VGND 0.01418f
C7736 XThR.Tn[3].t27 VGND 0.01553f
C7737 XThR.Tn[3].n83 VGND 0.03959f
C7738 XThR.Tn[3].n84 VGND 0.02781f
C7739 XThR.Tn[3].n86 VGND 0.08925f
C7740 XThR.Tn[3].n87 VGND 0.0811f
C7741 XThR.Tn[3].n88 VGND 0.17963f
C7742 XThR.Tn[3].n89 VGND 0.0381f
C7743 XThC.XTB4.Y.t1 VGND 0.12238f
C7744 XThC.XTB4.Y.n0 VGND 0.16166f
C7745 XThC.XTB4.Y.t4 VGND 0.02956f
C7746 XThC.XTB4.Y.t13 VGND 0.05016f
C7747 XThC.XTB4.Y.n1 VGND 0.05972f
C7748 XThC.XTB4.Y.t7 VGND 0.02956f
C7749 XThC.XTB4.Y.t17 VGND 0.05016f
C7750 XThC.XTB4.Y.n2 VGND 0.03074f
C7751 XThC.XTB4.Y.t10 VGND 0.02956f
C7752 XThC.XTB4.Y.t2 VGND 0.05016f
C7753 XThC.XTB4.Y.n3 VGND 0.06603f
C7754 XThC.XTB4.Y.t14 VGND 0.02956f
C7755 XThC.XTB4.Y.t3 VGND 0.05016f
C7756 XThC.XTB4.Y.n4 VGND 0.0613f
C7757 XThC.XTB4.Y.n5 VGND 0.03729f
C7758 XThC.XTB4.Y.n6 VGND 0.06174f
C7759 XThC.XTB4.Y.n7 VGND 0.02389f
C7760 XThC.XTB4.Y.n8 VGND 0.02916f
C7761 XThC.XTB4.Y.n9 VGND 0.06603f
C7762 XThC.XTB4.Y.n10 VGND 0.0331f
C7763 XThC.XTB4.Y.n11 VGND 0.06459f
C7764 XThC.XTB4.Y.t5 VGND 0.02956f
C7765 XThC.XTB4.Y.t16 VGND 0.05016f
C7766 XThC.XTB4.Y.n12 VGND 0.06761f
C7767 XThC.XTB4.Y.t9 VGND 0.02956f
C7768 XThC.XTB4.Y.t6 VGND 0.05016f
C7769 XThC.XTB4.Y.t15 VGND 0.02956f
C7770 XThC.XTB4.Y.t12 VGND 0.05016f
C7771 XThC.XTB4.Y.t11 VGND 0.02956f
C7772 XThC.XTB4.Y.t8 VGND 0.05016f
C7773 XThC.XTB4.Y.n13 VGND 0.08416f
C7774 XThC.XTB4.Y.n14 VGND 0.08889f
C7775 XThC.XTB4.Y.n15 VGND 0.03426f
C7776 XThC.XTB4.Y.n16 VGND 0.07234f
C7777 XThC.XTB4.Y.n17 VGND 0.0331f
C7778 XThC.XTB4.Y.n18 VGND 0.02701f
C7779 XThC.XTB4.Y.n19 VGND 0.63971f
C7780 XThC.XTB4.Y.n20 VGND 1.29767f
C7781 XThC.XTB4.Y.n21 VGND 0.08408f
C7782 XThC.XTB4.Y.t0 VGND 0.06491f
C7783 XThC.XTB4.Y.n22 VGND 0.04329f
C7784 XThC.Tn[0].t4 VGND 0.0118f
C7785 XThC.Tn[0].t3 VGND 0.0118f
C7786 XThC.Tn[0].n0 VGND 0.02383f
C7787 XThC.Tn[0].t6 VGND 0.0118f
C7788 XThC.Tn[0].t5 VGND 0.0118f
C7789 XThC.Tn[0].n1 VGND 0.02788f
C7790 XThC.Tn[0].n2 VGND 0.07804f
C7791 XThC.Tn[0].n3 VGND 0.01747f
C7792 XThC.Tn[0].n4 VGND 0.01747f
C7793 XThC.Tn[0].n5 VGND 0.01747f
C7794 XThC.Tn[0].n6 VGND 0.02911f
C7795 XThC.Tn[0].n7 VGND 0.0832f
C7796 XThC.Tn[0].n8 VGND 0.05143f
C7797 XThC.Tn[0].n9 VGND 0.05805f
C7798 XThC.Tn[0].t22 VGND 0.01022f
C7799 XThC.Tn[0].n10 VGND 0.02282f
C7800 XThC.Tn[0].n11 VGND 0.01304f
C7801 XThC.Tn[0].n12 VGND 0.01586f
C7802 XThC.Tn[0].t41 VGND 0.01022f
C7803 XThC.Tn[0].n13 VGND 0.02282f
C7804 XThC.Tn[0].n14 VGND 0.01304f
C7805 XThC.Tn[0].n15 VGND 0.07535f
C7806 XThC.Tn[0].t12 VGND 0.01022f
C7807 XThC.Tn[0].n16 VGND 0.02282f
C7808 XThC.Tn[0].n17 VGND 0.01304f
C7809 XThC.Tn[0].n18 VGND 0.07535f
C7810 XThC.Tn[0].t13 VGND 0.01022f
C7811 XThC.Tn[0].n19 VGND 0.02282f
C7812 XThC.Tn[0].n20 VGND 0.01304f
C7813 XThC.Tn[0].n21 VGND 0.07535f
C7814 XThC.Tn[0].t32 VGND 0.01022f
C7815 XThC.Tn[0].n22 VGND 0.02282f
C7816 XThC.Tn[0].n23 VGND 0.01304f
C7817 XThC.Tn[0].n24 VGND 0.07535f
C7818 XThC.Tn[0].t34 VGND 0.01022f
C7819 XThC.Tn[0].n25 VGND 0.02282f
C7820 XThC.Tn[0].n26 VGND 0.01304f
C7821 XThC.Tn[0].n27 VGND 0.07535f
C7822 XThC.Tn[0].t17 VGND 0.01022f
C7823 XThC.Tn[0].n28 VGND 0.02282f
C7824 XThC.Tn[0].n29 VGND 0.01304f
C7825 XThC.Tn[0].n30 VGND 0.07535f
C7826 XThC.Tn[0].t25 VGND 0.01022f
C7827 XThC.Tn[0].n31 VGND 0.02282f
C7828 XThC.Tn[0].n32 VGND 0.01304f
C7829 XThC.Tn[0].n33 VGND 0.07535f
C7830 XThC.Tn[0].t26 VGND 0.01022f
C7831 XThC.Tn[0].n34 VGND 0.02282f
C7832 XThC.Tn[0].n35 VGND 0.01304f
C7833 XThC.Tn[0].n36 VGND 0.07535f
C7834 XThC.Tn[0].t15 VGND 0.01022f
C7835 XThC.Tn[0].n37 VGND 0.02282f
C7836 XThC.Tn[0].n38 VGND 0.01304f
C7837 XThC.Tn[0].n39 VGND 0.07535f
C7838 XThC.Tn[0].t16 VGND 0.01022f
C7839 XThC.Tn[0].n40 VGND 0.02282f
C7840 XThC.Tn[0].n41 VGND 0.01304f
C7841 XThC.Tn[0].n42 VGND 0.07535f
C7842 XThC.Tn[0].t27 VGND 0.01022f
C7843 XThC.Tn[0].n43 VGND 0.02282f
C7844 XThC.Tn[0].n44 VGND 0.01304f
C7845 XThC.Tn[0].n45 VGND 0.07535f
C7846 XThC.Tn[0].t36 VGND 0.01022f
C7847 XThC.Tn[0].n46 VGND 0.02282f
C7848 XThC.Tn[0].n47 VGND 0.01304f
C7849 XThC.Tn[0].n48 VGND 0.07535f
C7850 XThC.Tn[0].t38 VGND 0.01022f
C7851 XThC.Tn[0].n49 VGND 0.02282f
C7852 XThC.Tn[0].n50 VGND 0.01304f
C7853 XThC.Tn[0].n51 VGND 0.07535f
C7854 XThC.Tn[0].t19 VGND 0.01022f
C7855 XThC.Tn[0].n52 VGND 0.02282f
C7856 XThC.Tn[0].n53 VGND 0.01304f
C7857 XThC.Tn[0].n54 VGND 0.07535f
C7858 XThC.Tn[0].t29 VGND 0.01022f
C7859 XThC.Tn[0].n55 VGND 0.02282f
C7860 XThC.Tn[0].n56 VGND 0.01304f
C7861 XThC.Tn[0].n57 VGND 0.07535f
C7862 XThC.Tn[0].n58 VGND 0.13474f
C7863 XThC.Tn[0].n59 VGND 0.03416f
C7864 XThC.Tn[0].n60 VGND 0.0247f
C7865 XThC.Tn[13].t6 VGND 0.01445f
C7866 XThC.Tn[13].t5 VGND 0.01445f
C7867 XThC.Tn[13].n0 VGND 0.03122f
C7868 XThC.Tn[13].t4 VGND 0.01445f
C7869 XThC.Tn[13].t7 VGND 0.01445f
C7870 XThC.Tn[13].n1 VGND 0.04921f
C7871 XThC.Tn[13].n2 VGND 0.13032f
C7872 XThC.Tn[13].t9 VGND 0.01445f
C7873 XThC.Tn[13].t8 VGND 0.01445f
C7874 XThC.Tn[13].n3 VGND 0.04387f
C7875 XThC.Tn[13].t11 VGND 0.01445f
C7876 XThC.Tn[13].t10 VGND 0.01445f
C7877 XThC.Tn[13].n4 VGND 0.03212f
C7878 XThC.Tn[13].n5 VGND 0.14294f
C7879 XThC.Tn[13].t29 VGND 0.01145f
C7880 XThC.Tn[13].t27 VGND 0.01251f
C7881 XThC.Tn[13].n7 VGND 0.02793f
C7882 XThC.Tn[13].n8 VGND 0.01596f
C7883 XThC.Tn[13].n9 VGND 0.01941f
C7884 XThC.Tn[13].t15 VGND 0.01145f
C7885 XThC.Tn[13].t12 VGND 0.01251f
C7886 XThC.Tn[13].n10 VGND 0.02793f
C7887 XThC.Tn[13].n11 VGND 0.01596f
C7888 XThC.Tn[13].n12 VGND 0.09223f
C7889 XThC.Tn[13].t20 VGND 0.01145f
C7890 XThC.Tn[13].t14 VGND 0.01251f
C7891 XThC.Tn[13].n13 VGND 0.02793f
C7892 XThC.Tn[13].n14 VGND 0.01596f
C7893 XThC.Tn[13].n15 VGND 0.09223f
C7894 XThC.Tn[13].t21 VGND 0.01145f
C7895 XThC.Tn[13].t16 VGND 0.01251f
C7896 XThC.Tn[13].n16 VGND 0.02793f
C7897 XThC.Tn[13].n17 VGND 0.01596f
C7898 XThC.Tn[13].n18 VGND 0.09223f
C7899 XThC.Tn[13].t40 VGND 0.01145f
C7900 XThC.Tn[13].t37 VGND 0.01251f
C7901 XThC.Tn[13].n19 VGND 0.02793f
C7902 XThC.Tn[13].n20 VGND 0.01596f
C7903 XThC.Tn[13].n21 VGND 0.09223f
C7904 XThC.Tn[13].t41 VGND 0.01145f
C7905 XThC.Tn[13].t38 VGND 0.01251f
C7906 XThC.Tn[13].n22 VGND 0.02793f
C7907 XThC.Tn[13].n23 VGND 0.01596f
C7908 XThC.Tn[13].n24 VGND 0.09223f
C7909 XThC.Tn[13].t25 VGND 0.01145f
C7910 XThC.Tn[13].t19 VGND 0.01251f
C7911 XThC.Tn[13].n25 VGND 0.02793f
C7912 XThC.Tn[13].n26 VGND 0.01596f
C7913 XThC.Tn[13].n27 VGND 0.09223f
C7914 XThC.Tn[13].t32 VGND 0.01145f
C7915 XThC.Tn[13].t28 VGND 0.01251f
C7916 XThC.Tn[13].n28 VGND 0.02793f
C7917 XThC.Tn[13].n29 VGND 0.01596f
C7918 XThC.Tn[13].n30 VGND 0.09223f
C7919 XThC.Tn[13].t34 VGND 0.01145f
C7920 XThC.Tn[13].t30 VGND 0.01251f
C7921 XThC.Tn[13].n31 VGND 0.02793f
C7922 XThC.Tn[13].n32 VGND 0.01596f
C7923 XThC.Tn[13].n33 VGND 0.09223f
C7924 XThC.Tn[13].t22 VGND 0.01145f
C7925 XThC.Tn[13].t17 VGND 0.01251f
C7926 XThC.Tn[13].n34 VGND 0.02793f
C7927 XThC.Tn[13].n35 VGND 0.01596f
C7928 XThC.Tn[13].n36 VGND 0.09223f
C7929 XThC.Tn[13].t24 VGND 0.01145f
C7930 XThC.Tn[13].t18 VGND 0.01251f
C7931 XThC.Tn[13].n37 VGND 0.02793f
C7932 XThC.Tn[13].n38 VGND 0.01596f
C7933 XThC.Tn[13].n39 VGND 0.09223f
C7934 XThC.Tn[13].t35 VGND 0.01145f
C7935 XThC.Tn[13].t31 VGND 0.01251f
C7936 XThC.Tn[13].n40 VGND 0.02793f
C7937 XThC.Tn[13].n41 VGND 0.01596f
C7938 XThC.Tn[13].n42 VGND 0.09223f
C7939 XThC.Tn[13].t43 VGND 0.01145f
C7940 XThC.Tn[13].t39 VGND 0.01251f
C7941 XThC.Tn[13].n43 VGND 0.02793f
C7942 XThC.Tn[13].n44 VGND 0.01596f
C7943 XThC.Tn[13].n45 VGND 0.09223f
C7944 XThC.Tn[13].t13 VGND 0.01145f
C7945 XThC.Tn[13].t42 VGND 0.01251f
C7946 XThC.Tn[13].n46 VGND 0.02793f
C7947 XThC.Tn[13].n47 VGND 0.01596f
C7948 XThC.Tn[13].n48 VGND 0.09223f
C7949 XThC.Tn[13].t26 VGND 0.01145f
C7950 XThC.Tn[13].t23 VGND 0.01251f
C7951 XThC.Tn[13].n49 VGND 0.02793f
C7952 XThC.Tn[13].n50 VGND 0.01596f
C7953 XThC.Tn[13].n51 VGND 0.09223f
C7954 XThC.Tn[13].t36 VGND 0.01145f
C7955 XThC.Tn[13].t33 VGND 0.01251f
C7956 XThC.Tn[13].n52 VGND 0.02793f
C7957 XThC.Tn[13].n53 VGND 0.01596f
C7958 XThC.Tn[13].n54 VGND 0.09223f
C7959 XThC.Tn[13].n55 VGND 0.51097f
C7960 XThC.Tn[13].n56 VGND 0.04181f
C7961 XThC.Tn[13].n57 VGND 0.01878f
C7962 XThC.Tn[13].n58 VGND 0.02342f
C7963 XThC.Tn[13].n59 VGND 0.04331f
C7964 XThC.Tn[12].n0 VGND 0.01883f
C7965 XThC.Tn[12].n1 VGND 0.02348f
C7966 XThC.Tn[12].n2 VGND 0.04736f
C7967 XThC.Tn[12].t5 VGND 0.01448f
C7968 XThC.Tn[12].t6 VGND 0.01448f
C7969 XThC.Tn[12].n3 VGND 0.03129f
C7970 XThC.Tn[12].t4 VGND 0.01448f
C7971 XThC.Tn[12].t7 VGND 0.01448f
C7972 XThC.Tn[12].n4 VGND 0.04762f
C7973 XThC.Tn[12].n5 VGND 0.13232f
C7974 XThC.Tn[12].t9 VGND 0.01448f
C7975 XThC.Tn[12].t8 VGND 0.01448f
C7976 XThC.Tn[12].n6 VGND 0.04397f
C7977 XThC.Tn[12].t11 VGND 0.01448f
C7978 XThC.Tn[12].t10 VGND 0.01448f
C7979 XThC.Tn[12].n7 VGND 0.03219f
C7980 XThC.Tn[12].n8 VGND 0.14328f
C7981 XThC.Tn[12].n9 VGND 0.02081f
C7982 XThC.Tn[12].t37 VGND 0.01148f
C7983 XThC.Tn[12].t35 VGND 0.01254f
C7984 XThC.Tn[12].n10 VGND 0.028f
C7985 XThC.Tn[12].n11 VGND 0.016f
C7986 XThC.Tn[12].n12 VGND 0.01946f
C7987 XThC.Tn[12].t23 VGND 0.01148f
C7988 XThC.Tn[12].t20 VGND 0.01254f
C7989 XThC.Tn[12].n13 VGND 0.028f
C7990 XThC.Tn[12].n14 VGND 0.016f
C7991 XThC.Tn[12].n15 VGND 0.09245f
C7992 XThC.Tn[12].t28 VGND 0.01148f
C7993 XThC.Tn[12].t22 VGND 0.01254f
C7994 XThC.Tn[12].n16 VGND 0.028f
C7995 XThC.Tn[12].n17 VGND 0.016f
C7996 XThC.Tn[12].n18 VGND 0.09245f
C7997 XThC.Tn[12].t29 VGND 0.01148f
C7998 XThC.Tn[12].t24 VGND 0.01254f
C7999 XThC.Tn[12].n19 VGND 0.028f
C8000 XThC.Tn[12].n20 VGND 0.016f
C8001 XThC.Tn[12].n21 VGND 0.09245f
C8002 XThC.Tn[12].t16 VGND 0.01148f
C8003 XThC.Tn[12].t13 VGND 0.01254f
C8004 XThC.Tn[12].n22 VGND 0.028f
C8005 XThC.Tn[12].n23 VGND 0.016f
C8006 XThC.Tn[12].n24 VGND 0.09245f
C8007 XThC.Tn[12].t17 VGND 0.01148f
C8008 XThC.Tn[12].t14 VGND 0.01254f
C8009 XThC.Tn[12].n25 VGND 0.028f
C8010 XThC.Tn[12].n26 VGND 0.016f
C8011 XThC.Tn[12].n27 VGND 0.09245f
C8012 XThC.Tn[12].t33 VGND 0.01148f
C8013 XThC.Tn[12].t27 VGND 0.01254f
C8014 XThC.Tn[12].n28 VGND 0.028f
C8015 XThC.Tn[12].n29 VGND 0.016f
C8016 XThC.Tn[12].n30 VGND 0.09245f
C8017 XThC.Tn[12].t40 VGND 0.01148f
C8018 XThC.Tn[12].t36 VGND 0.01254f
C8019 XThC.Tn[12].n31 VGND 0.028f
C8020 XThC.Tn[12].n32 VGND 0.016f
C8021 XThC.Tn[12].n33 VGND 0.09245f
C8022 XThC.Tn[12].t42 VGND 0.01148f
C8023 XThC.Tn[12].t38 VGND 0.01254f
C8024 XThC.Tn[12].n34 VGND 0.028f
C8025 XThC.Tn[12].n35 VGND 0.016f
C8026 XThC.Tn[12].n36 VGND 0.09245f
C8027 XThC.Tn[12].t30 VGND 0.01148f
C8028 XThC.Tn[12].t25 VGND 0.01254f
C8029 XThC.Tn[12].n37 VGND 0.028f
C8030 XThC.Tn[12].n38 VGND 0.016f
C8031 XThC.Tn[12].n39 VGND 0.09245f
C8032 XThC.Tn[12].t32 VGND 0.01148f
C8033 XThC.Tn[12].t26 VGND 0.01254f
C8034 XThC.Tn[12].n40 VGND 0.028f
C8035 XThC.Tn[12].n41 VGND 0.016f
C8036 XThC.Tn[12].n42 VGND 0.09245f
C8037 XThC.Tn[12].t43 VGND 0.01148f
C8038 XThC.Tn[12].t39 VGND 0.01254f
C8039 XThC.Tn[12].n43 VGND 0.028f
C8040 XThC.Tn[12].n44 VGND 0.016f
C8041 XThC.Tn[12].n45 VGND 0.09245f
C8042 XThC.Tn[12].t19 VGND 0.01148f
C8043 XThC.Tn[12].t15 VGND 0.01254f
C8044 XThC.Tn[12].n46 VGND 0.028f
C8045 XThC.Tn[12].n47 VGND 0.016f
C8046 XThC.Tn[12].n48 VGND 0.09245f
C8047 XThC.Tn[12].t21 VGND 0.01148f
C8048 XThC.Tn[12].t18 VGND 0.01254f
C8049 XThC.Tn[12].n49 VGND 0.028f
C8050 XThC.Tn[12].n50 VGND 0.016f
C8051 XThC.Tn[12].n51 VGND 0.09245f
C8052 XThC.Tn[12].t34 VGND 0.01148f
C8053 XThC.Tn[12].t31 VGND 0.01254f
C8054 XThC.Tn[12].n52 VGND 0.028f
C8055 XThC.Tn[12].n53 VGND 0.016f
C8056 XThC.Tn[12].n54 VGND 0.09245f
C8057 XThC.Tn[12].t12 VGND 0.01148f
C8058 XThC.Tn[12].t41 VGND 0.01254f
C8059 XThC.Tn[12].n55 VGND 0.028f
C8060 XThC.Tn[12].n56 VGND 0.016f
C8061 XThC.Tn[12].n57 VGND 0.09245f
C8062 XThC.Tn[12].n58 VGND 0.5067f
C8063 XThC.Tn[12].n59 VGND 0.03519f
C8064 XThC.Tn[11].t11 VGND 0.01474f
C8065 XThC.Tn[11].t8 VGND 0.01474f
C8066 XThC.Tn[11].n0 VGND 0.03186f
C8067 XThC.Tn[11].t3 VGND 0.01474f
C8068 XThC.Tn[11].t1 VGND 0.01474f
C8069 XThC.Tn[11].n1 VGND 0.05022f
C8070 XThC.Tn[11].n2 VGND 0.13299f
C8071 XThC.Tn[11].t4 VGND 0.01474f
C8072 XThC.Tn[11].t7 VGND 0.01474f
C8073 XThC.Tn[11].n3 VGND 0.04477f
C8074 XThC.Tn[11].t6 VGND 0.01474f
C8075 XThC.Tn[11].t5 VGND 0.01474f
C8076 XThC.Tn[11].n4 VGND 0.03278f
C8077 XThC.Tn[11].n5 VGND 0.14588f
C8078 XThC.Tn[11].t20 VGND 0.01169f
C8079 XThC.Tn[11].t18 VGND 0.01277f
C8080 XThC.Tn[11].n7 VGND 0.02851f
C8081 XThC.Tn[11].n8 VGND 0.01629f
C8082 XThC.Tn[11].n9 VGND 0.01981f
C8083 XThC.Tn[11].t38 VGND 0.01169f
C8084 XThC.Tn[11].t35 VGND 0.01277f
C8085 XThC.Tn[11].n10 VGND 0.02851f
C8086 XThC.Tn[11].n11 VGND 0.01629f
C8087 XThC.Tn[11].n12 VGND 0.09412f
C8088 XThC.Tn[11].t43 VGND 0.01169f
C8089 XThC.Tn[11].t37 VGND 0.01277f
C8090 XThC.Tn[11].n13 VGND 0.02851f
C8091 XThC.Tn[11].n14 VGND 0.01629f
C8092 XThC.Tn[11].n15 VGND 0.09412f
C8093 XThC.Tn[11].t12 VGND 0.01169f
C8094 XThC.Tn[11].t39 VGND 0.01277f
C8095 XThC.Tn[11].n16 VGND 0.02851f
C8096 XThC.Tn[11].n17 VGND 0.01629f
C8097 XThC.Tn[11].n18 VGND 0.09412f
C8098 XThC.Tn[11].t31 VGND 0.01169f
C8099 XThC.Tn[11].t28 VGND 0.01277f
C8100 XThC.Tn[11].n19 VGND 0.02851f
C8101 XThC.Tn[11].n20 VGND 0.01629f
C8102 XThC.Tn[11].n21 VGND 0.09412f
C8103 XThC.Tn[11].t32 VGND 0.01169f
C8104 XThC.Tn[11].t29 VGND 0.01277f
C8105 XThC.Tn[11].n22 VGND 0.02851f
C8106 XThC.Tn[11].n23 VGND 0.01629f
C8107 XThC.Tn[11].n24 VGND 0.09412f
C8108 XThC.Tn[11].t16 VGND 0.01169f
C8109 XThC.Tn[11].t42 VGND 0.01277f
C8110 XThC.Tn[11].n25 VGND 0.02851f
C8111 XThC.Tn[11].n26 VGND 0.01629f
C8112 XThC.Tn[11].n27 VGND 0.09412f
C8113 XThC.Tn[11].t23 VGND 0.01169f
C8114 XThC.Tn[11].t19 VGND 0.01277f
C8115 XThC.Tn[11].n28 VGND 0.02851f
C8116 XThC.Tn[11].n29 VGND 0.01629f
C8117 XThC.Tn[11].n30 VGND 0.09412f
C8118 XThC.Tn[11].t25 VGND 0.01169f
C8119 XThC.Tn[11].t21 VGND 0.01277f
C8120 XThC.Tn[11].n31 VGND 0.02851f
C8121 XThC.Tn[11].n32 VGND 0.01629f
C8122 XThC.Tn[11].n33 VGND 0.09412f
C8123 XThC.Tn[11].t13 VGND 0.01169f
C8124 XThC.Tn[11].t40 VGND 0.01277f
C8125 XThC.Tn[11].n34 VGND 0.02851f
C8126 XThC.Tn[11].n35 VGND 0.01629f
C8127 XThC.Tn[11].n36 VGND 0.09412f
C8128 XThC.Tn[11].t15 VGND 0.01169f
C8129 XThC.Tn[11].t41 VGND 0.01277f
C8130 XThC.Tn[11].n37 VGND 0.02851f
C8131 XThC.Tn[11].n38 VGND 0.01629f
C8132 XThC.Tn[11].n39 VGND 0.09412f
C8133 XThC.Tn[11].t26 VGND 0.01169f
C8134 XThC.Tn[11].t22 VGND 0.01277f
C8135 XThC.Tn[11].n40 VGND 0.02851f
C8136 XThC.Tn[11].n41 VGND 0.01629f
C8137 XThC.Tn[11].n42 VGND 0.09412f
C8138 XThC.Tn[11].t34 VGND 0.01169f
C8139 XThC.Tn[11].t30 VGND 0.01277f
C8140 XThC.Tn[11].n43 VGND 0.02851f
C8141 XThC.Tn[11].n44 VGND 0.01629f
C8142 XThC.Tn[11].n45 VGND 0.09412f
C8143 XThC.Tn[11].t36 VGND 0.01169f
C8144 XThC.Tn[11].t33 VGND 0.01277f
C8145 XThC.Tn[11].n46 VGND 0.02851f
C8146 XThC.Tn[11].n47 VGND 0.01629f
C8147 XThC.Tn[11].n48 VGND 0.09412f
C8148 XThC.Tn[11].t17 VGND 0.01169f
C8149 XThC.Tn[11].t14 VGND 0.01277f
C8150 XThC.Tn[11].n49 VGND 0.02851f
C8151 XThC.Tn[11].n50 VGND 0.01629f
C8152 XThC.Tn[11].n51 VGND 0.09412f
C8153 XThC.Tn[11].t27 VGND 0.01169f
C8154 XThC.Tn[11].t24 VGND 0.01277f
C8155 XThC.Tn[11].n52 VGND 0.02851f
C8156 XThC.Tn[11].n53 VGND 0.01629f
C8157 XThC.Tn[11].n54 VGND 0.09412f
C8158 XThC.Tn[11].n55 VGND 0.04302f
C8159 XThC.Tn[11].n56 VGND 0.01917f
C8160 XThC.Tn[11].n57 VGND 0.0239f
C8161 XThC.Tn[11].n58 VGND 0.0442f
C8162 XThC.Tn[9].n0 VGND 0.02381f
C8163 XThC.Tn[9].n1 VGND 0.0191f
C8164 XThC.Tn[9].n2 VGND 0.04403f
C8165 XThC.Tn[9].t26 VGND 0.01164f
C8166 XThC.Tn[9].t12 VGND 0.01272f
C8167 XThC.Tn[9].n3 VGND 0.0284f
C8168 XThC.Tn[9].n4 VGND 0.01623f
C8169 XThC.Tn[9].n5 VGND 0.01974f
C8170 XThC.Tn[9].t13 VGND 0.01164f
C8171 XThC.Tn[9].t30 VGND 0.01272f
C8172 XThC.Tn[9].n6 VGND 0.0284f
C8173 XThC.Tn[9].n7 VGND 0.01623f
C8174 XThC.Tn[9].n8 VGND 0.09378f
C8175 XThC.Tn[9].t15 VGND 0.01164f
C8176 XThC.Tn[9].t34 VGND 0.01272f
C8177 XThC.Tn[9].n9 VGND 0.0284f
C8178 XThC.Tn[9].n10 VGND 0.01623f
C8179 XThC.Tn[9].n11 VGND 0.09378f
C8180 XThC.Tn[9].t17 VGND 0.01164f
C8181 XThC.Tn[9].t35 VGND 0.01272f
C8182 XThC.Tn[9].n12 VGND 0.0284f
C8183 XThC.Tn[9].n13 VGND 0.01623f
C8184 XThC.Tn[9].n14 VGND 0.09378f
C8185 XThC.Tn[9].t39 VGND 0.01164f
C8186 XThC.Tn[9].t24 VGND 0.01272f
C8187 XThC.Tn[9].n15 VGND 0.0284f
C8188 XThC.Tn[9].n16 VGND 0.01623f
C8189 XThC.Tn[9].n17 VGND 0.09378f
C8190 XThC.Tn[9].t40 VGND 0.01164f
C8191 XThC.Tn[9].t25 VGND 0.01272f
C8192 XThC.Tn[9].n18 VGND 0.0284f
C8193 XThC.Tn[9].n19 VGND 0.01623f
C8194 XThC.Tn[9].n20 VGND 0.09378f
C8195 XThC.Tn[9].t22 VGND 0.01164f
C8196 XThC.Tn[9].t38 VGND 0.01272f
C8197 XThC.Tn[9].n21 VGND 0.0284f
C8198 XThC.Tn[9].n22 VGND 0.01623f
C8199 XThC.Tn[9].n23 VGND 0.09378f
C8200 XThC.Tn[9].t28 VGND 0.01164f
C8201 XThC.Tn[9].t14 VGND 0.01272f
C8202 XThC.Tn[9].n24 VGND 0.0284f
C8203 XThC.Tn[9].n25 VGND 0.01623f
C8204 XThC.Tn[9].n26 VGND 0.09378f
C8205 XThC.Tn[9].t31 VGND 0.01164f
C8206 XThC.Tn[9].t16 VGND 0.01272f
C8207 XThC.Tn[9].n27 VGND 0.0284f
C8208 XThC.Tn[9].n28 VGND 0.01623f
C8209 XThC.Tn[9].n29 VGND 0.09378f
C8210 XThC.Tn[9].t19 VGND 0.01164f
C8211 XThC.Tn[9].t36 VGND 0.01272f
C8212 XThC.Tn[9].n30 VGND 0.0284f
C8213 XThC.Tn[9].n31 VGND 0.01623f
C8214 XThC.Tn[9].n32 VGND 0.09378f
C8215 XThC.Tn[9].t21 VGND 0.01164f
C8216 XThC.Tn[9].t37 VGND 0.01272f
C8217 XThC.Tn[9].n33 VGND 0.0284f
C8218 XThC.Tn[9].n34 VGND 0.01623f
C8219 XThC.Tn[9].n35 VGND 0.09378f
C8220 XThC.Tn[9].t32 VGND 0.01164f
C8221 XThC.Tn[9].t18 VGND 0.01272f
C8222 XThC.Tn[9].n36 VGND 0.0284f
C8223 XThC.Tn[9].n37 VGND 0.01623f
C8224 XThC.Tn[9].n38 VGND 0.09378f
C8225 XThC.Tn[9].t42 VGND 0.01164f
C8226 XThC.Tn[9].t27 VGND 0.01272f
C8227 XThC.Tn[9].n39 VGND 0.0284f
C8228 XThC.Tn[9].n40 VGND 0.01623f
C8229 XThC.Tn[9].n41 VGND 0.09378f
C8230 XThC.Tn[9].t43 VGND 0.01164f
C8231 XThC.Tn[9].t29 VGND 0.01272f
C8232 XThC.Tn[9].n42 VGND 0.0284f
C8233 XThC.Tn[9].n43 VGND 0.01623f
C8234 XThC.Tn[9].n44 VGND 0.09378f
C8235 XThC.Tn[9].t23 VGND 0.01164f
C8236 XThC.Tn[9].t41 VGND 0.01272f
C8237 XThC.Tn[9].n45 VGND 0.0284f
C8238 XThC.Tn[9].n46 VGND 0.01623f
C8239 XThC.Tn[9].n47 VGND 0.09378f
C8240 XThC.Tn[9].t33 VGND 0.01164f
C8241 XThC.Tn[9].t20 VGND 0.01272f
C8242 XThC.Tn[9].n48 VGND 0.0284f
C8243 XThC.Tn[9].n49 VGND 0.01623f
C8244 XThC.Tn[9].n50 VGND 0.09378f
C8245 XThC.Tn[9].n51 VGND 0.04286f
C8246 XThC.Tn[9].t0 VGND 0.01469f
C8247 XThC.Tn[9].t3 VGND 0.01469f
C8248 XThC.Tn[9].n52 VGND 0.03174f
C8249 XThC.Tn[9].t2 VGND 0.01469f
C8250 XThC.Tn[9].t1 VGND 0.01469f
C8251 XThC.Tn[9].n53 VGND 0.05003f
C8252 XThC.Tn[9].n54 VGND 0.1325f
C8253 XThC.Tn[9].t9 VGND 0.01469f
C8254 XThC.Tn[9].t8 VGND 0.01469f
C8255 XThC.Tn[9].n56 VGND 0.0446f
C8256 XThC.Tn[9].t11 VGND 0.01469f
C8257 XThC.Tn[9].t10 VGND 0.01469f
C8258 XThC.Tn[9].n57 VGND 0.03266f
C8259 XThC.Tn[9].n58 VGND 0.14534f
C8260 XThC.Tn[5].t11 VGND 0.0121f
C8261 XThC.Tn[5].t10 VGND 0.0121f
C8262 XThC.Tn[5].n0 VGND 0.02443f
C8263 XThC.Tn[5].t9 VGND 0.0121f
C8264 XThC.Tn[5].t8 VGND 0.0121f
C8265 XThC.Tn[5].n1 VGND 0.02858f
C8266 XThC.Tn[5].n2 VGND 0.08573f
C8267 XThC.Tn[5].n3 VGND 0.01791f
C8268 XThC.Tn[5].n4 VGND 0.01791f
C8269 XThC.Tn[5].n5 VGND 0.01791f
C8270 XThC.Tn[5].n6 VGND 0.02985f
C8271 XThC.Tn[5].n7 VGND 0.0853f
C8272 XThC.Tn[5].n8 VGND 0.05273f
C8273 XThC.Tn[5].n9 VGND 0.05951f
C8274 XThC.Tn[5].t33 VGND 0.01048f
C8275 XThC.Tn[5].n10 VGND 0.0234f
C8276 XThC.Tn[5].n11 VGND 0.01337f
C8277 XThC.Tn[5].n12 VGND 0.01626f
C8278 XThC.Tn[5].t19 VGND 0.01048f
C8279 XThC.Tn[5].n13 VGND 0.0234f
C8280 XThC.Tn[5].n14 VGND 0.01337f
C8281 XThC.Tn[5].n15 VGND 0.07725f
C8282 XThC.Tn[5].t23 VGND 0.01048f
C8283 XThC.Tn[5].n16 VGND 0.0234f
C8284 XThC.Tn[5].n17 VGND 0.01337f
C8285 XThC.Tn[5].n18 VGND 0.07725f
C8286 XThC.Tn[5].t24 VGND 0.01048f
C8287 XThC.Tn[5].n19 VGND 0.0234f
C8288 XThC.Tn[5].n20 VGND 0.01337f
C8289 XThC.Tn[5].n21 VGND 0.07725f
C8290 XThC.Tn[5].t13 VGND 0.01048f
C8291 XThC.Tn[5].n22 VGND 0.0234f
C8292 XThC.Tn[5].n23 VGND 0.01337f
C8293 XThC.Tn[5].n24 VGND 0.07725f
C8294 XThC.Tn[5].t14 VGND 0.01048f
C8295 XThC.Tn[5].n25 VGND 0.0234f
C8296 XThC.Tn[5].n26 VGND 0.01337f
C8297 XThC.Tn[5].n27 VGND 0.07725f
C8298 XThC.Tn[5].t27 VGND 0.01048f
C8299 XThC.Tn[5].n28 VGND 0.0234f
C8300 XThC.Tn[5].n29 VGND 0.01337f
C8301 XThC.Tn[5].n30 VGND 0.07725f
C8302 XThC.Tn[5].t35 VGND 0.01048f
C8303 XThC.Tn[5].n31 VGND 0.0234f
C8304 XThC.Tn[5].n32 VGND 0.01337f
C8305 XThC.Tn[5].n33 VGND 0.07725f
C8306 XThC.Tn[5].t37 VGND 0.01048f
C8307 XThC.Tn[5].n34 VGND 0.0234f
C8308 XThC.Tn[5].n35 VGND 0.01337f
C8309 XThC.Tn[5].n36 VGND 0.07725f
C8310 XThC.Tn[5].t25 VGND 0.01048f
C8311 XThC.Tn[5].n37 VGND 0.0234f
C8312 XThC.Tn[5].n38 VGND 0.01337f
C8313 XThC.Tn[5].n39 VGND 0.07725f
C8314 XThC.Tn[5].t26 VGND 0.01048f
C8315 XThC.Tn[5].n40 VGND 0.0234f
C8316 XThC.Tn[5].n41 VGND 0.01337f
C8317 XThC.Tn[5].n42 VGND 0.07725f
C8318 XThC.Tn[5].t39 VGND 0.01048f
C8319 XThC.Tn[5].n43 VGND 0.0234f
C8320 XThC.Tn[5].n44 VGND 0.01337f
C8321 XThC.Tn[5].n45 VGND 0.07725f
C8322 XThC.Tn[5].t16 VGND 0.01048f
C8323 XThC.Tn[5].n46 VGND 0.0234f
C8324 XThC.Tn[5].n47 VGND 0.01337f
C8325 XThC.Tn[5].n48 VGND 0.07725f
C8326 XThC.Tn[5].t18 VGND 0.01048f
C8327 XThC.Tn[5].n49 VGND 0.0234f
C8328 XThC.Tn[5].n50 VGND 0.01337f
C8329 XThC.Tn[5].n51 VGND 0.07725f
C8330 XThC.Tn[5].t30 VGND 0.01048f
C8331 XThC.Tn[5].n52 VGND 0.0234f
C8332 XThC.Tn[5].n53 VGND 0.01337f
C8333 XThC.Tn[5].n54 VGND 0.07725f
C8334 XThC.Tn[5].t41 VGND 0.01048f
C8335 XThC.Tn[5].n55 VGND 0.0234f
C8336 XThC.Tn[5].n56 VGND 0.01337f
C8337 XThC.Tn[5].n57 VGND 0.07725f
C8338 XThC.Tn[5].n58 VGND 0.2186f
C8339 XThC.Tn[5].n59 VGND 0.04035f
C8340 XThR.Tn[9].t2 VGND 0.01931f
C8341 XThR.Tn[9].t0 VGND 0.01931f
C8342 XThR.Tn[9].n0 VGND 0.05863f
C8343 XThR.Tn[9].t3 VGND 0.01931f
C8344 XThR.Tn[9].t1 VGND 0.01931f
C8345 XThR.Tn[9].n1 VGND 0.04293f
C8346 XThR.Tn[9].n2 VGND 0.19519f
C8347 XThR.Tn[9].t5 VGND 0.01255f
C8348 XThR.Tn[9].t7 VGND 0.01255f
C8349 XThR.Tn[9].n3 VGND 0.03131f
C8350 XThR.Tn[9].t4 VGND 0.01255f
C8351 XThR.Tn[9].t6 VGND 0.01255f
C8352 XThR.Tn[9].n4 VGND 0.0251f
C8353 XThR.Tn[9].n5 VGND 0.06315f
C8354 XThR.Tn[9].t17 VGND 0.01509f
C8355 XThR.Tn[9].t71 VGND 0.01653f
C8356 XThR.Tn[9].n6 VGND 0.04036f
C8357 XThR.Tn[9].n7 VGND 0.07752f
C8358 XThR.Tn[9].t35 VGND 0.01509f
C8359 XThR.Tn[9].t28 VGND 0.01653f
C8360 XThR.Tn[9].n8 VGND 0.04036f
C8361 XThR.Tn[9].t50 VGND 0.01504f
C8362 XThR.Tn[9].t19 VGND 0.01647f
C8363 XThR.Tn[9].n9 VGND 0.04199f
C8364 XThR.Tn[9].n10 VGND 0.0295f
C8365 XThR.Tn[9].n12 VGND 0.09466f
C8366 XThR.Tn[9].t72 VGND 0.01509f
C8367 XThR.Tn[9].t64 VGND 0.01653f
C8368 XThR.Tn[9].n13 VGND 0.04036f
C8369 XThR.Tn[9].t26 VGND 0.01504f
C8370 XThR.Tn[9].t59 VGND 0.01647f
C8371 XThR.Tn[9].n14 VGND 0.04199f
C8372 XThR.Tn[9].n15 VGND 0.0295f
C8373 XThR.Tn[9].n17 VGND 0.09466f
C8374 XThR.Tn[9].t29 VGND 0.01509f
C8375 XThR.Tn[9].t21 VGND 0.01653f
C8376 XThR.Tn[9].n18 VGND 0.04036f
C8377 XThR.Tn[9].t41 VGND 0.01504f
C8378 XThR.Tn[9].t15 VGND 0.01647f
C8379 XThR.Tn[9].n19 VGND 0.04199f
C8380 XThR.Tn[9].n20 VGND 0.0295f
C8381 XThR.Tn[9].n22 VGND 0.09466f
C8382 XThR.Tn[9].t56 VGND 0.01509f
C8383 XThR.Tn[9].t46 VGND 0.01653f
C8384 XThR.Tn[9].n23 VGND 0.04036f
C8385 XThR.Tn[9].t73 VGND 0.01504f
C8386 XThR.Tn[9].t42 VGND 0.01647f
C8387 XThR.Tn[9].n24 VGND 0.04199f
C8388 XThR.Tn[9].n25 VGND 0.0295f
C8389 XThR.Tn[9].n27 VGND 0.09466f
C8390 XThR.Tn[9].t31 VGND 0.01509f
C8391 XThR.Tn[9].t23 VGND 0.01653f
C8392 XThR.Tn[9].n28 VGND 0.04036f
C8393 XThR.Tn[9].t44 VGND 0.01504f
C8394 XThR.Tn[9].t16 VGND 0.01647f
C8395 XThR.Tn[9].n29 VGND 0.04199f
C8396 XThR.Tn[9].n30 VGND 0.0295f
C8397 XThR.Tn[9].n32 VGND 0.09466f
C8398 XThR.Tn[9].t67 VGND 0.01509f
C8399 XThR.Tn[9].t37 VGND 0.01653f
C8400 XThR.Tn[9].n33 VGND 0.04036f
C8401 XThR.Tn[9].t20 VGND 0.01504f
C8402 XThR.Tn[9].t33 VGND 0.01647f
C8403 XThR.Tn[9].n34 VGND 0.04199f
C8404 XThR.Tn[9].n35 VGND 0.0295f
C8405 XThR.Tn[9].n37 VGND 0.09466f
C8406 XThR.Tn[9].t36 VGND 0.01509f
C8407 XThR.Tn[9].t32 VGND 0.01653f
C8408 XThR.Tn[9].n38 VGND 0.04036f
C8409 XThR.Tn[9].t51 VGND 0.01504f
C8410 XThR.Tn[9].t25 VGND 0.01647f
C8411 XThR.Tn[9].n39 VGND 0.04199f
C8412 XThR.Tn[9].n40 VGND 0.0295f
C8413 XThR.Tn[9].n42 VGND 0.09466f
C8414 XThR.Tn[9].t39 VGND 0.01509f
C8415 XThR.Tn[9].t45 VGND 0.01653f
C8416 XThR.Tn[9].n43 VGND 0.04036f
C8417 XThR.Tn[9].t55 VGND 0.01504f
C8418 XThR.Tn[9].t40 VGND 0.01647f
C8419 XThR.Tn[9].n44 VGND 0.04199f
C8420 XThR.Tn[9].n45 VGND 0.0295f
C8421 XThR.Tn[9].n47 VGND 0.09466f
C8422 XThR.Tn[9].t58 VGND 0.01509f
C8423 XThR.Tn[9].t66 VGND 0.01653f
C8424 XThR.Tn[9].n48 VGND 0.04036f
C8425 XThR.Tn[9].t13 VGND 0.01504f
C8426 XThR.Tn[9].t60 VGND 0.01647f
C8427 XThR.Tn[9].n49 VGND 0.04199f
C8428 XThR.Tn[9].n50 VGND 0.0295f
C8429 XThR.Tn[9].n52 VGND 0.09466f
C8430 XThR.Tn[9].t48 VGND 0.01509f
C8431 XThR.Tn[9].t24 VGND 0.01653f
C8432 XThR.Tn[9].n53 VGND 0.04036f
C8433 XThR.Tn[9].t65 VGND 0.01504f
C8434 XThR.Tn[9].t18 VGND 0.01647f
C8435 XThR.Tn[9].n54 VGND 0.04199f
C8436 XThR.Tn[9].n55 VGND 0.0295f
C8437 XThR.Tn[9].n57 VGND 0.09466f
C8438 XThR.Tn[9].t70 VGND 0.01509f
C8439 XThR.Tn[9].t62 VGND 0.01653f
C8440 XThR.Tn[9].n58 VGND 0.04036f
C8441 XThR.Tn[9].t22 VGND 0.01504f
C8442 XThR.Tn[9].t52 VGND 0.01647f
C8443 XThR.Tn[9].n59 VGND 0.04199f
C8444 XThR.Tn[9].n60 VGND 0.0295f
C8445 XThR.Tn[9].n62 VGND 0.09466f
C8446 XThR.Tn[9].t38 VGND 0.01509f
C8447 XThR.Tn[9].t34 VGND 0.01653f
C8448 XThR.Tn[9].n63 VGND 0.04036f
C8449 XThR.Tn[9].t53 VGND 0.01504f
C8450 XThR.Tn[9].t27 VGND 0.01647f
C8451 XThR.Tn[9].n64 VGND 0.04199f
C8452 XThR.Tn[9].n65 VGND 0.0295f
C8453 XThR.Tn[9].n67 VGND 0.09466f
C8454 XThR.Tn[9].t57 VGND 0.01509f
C8455 XThR.Tn[9].t47 VGND 0.01653f
C8456 XThR.Tn[9].n68 VGND 0.04036f
C8457 XThR.Tn[9].t12 VGND 0.01504f
C8458 XThR.Tn[9].t43 VGND 0.01647f
C8459 XThR.Tn[9].n69 VGND 0.04199f
C8460 XThR.Tn[9].n70 VGND 0.0295f
C8461 XThR.Tn[9].n72 VGND 0.09466f
C8462 XThR.Tn[9].t14 VGND 0.01509f
C8463 XThR.Tn[9].t69 VGND 0.01653f
C8464 XThR.Tn[9].n73 VGND 0.04036f
C8465 XThR.Tn[9].t30 VGND 0.01504f
C8466 XThR.Tn[9].t61 VGND 0.01647f
C8467 XThR.Tn[9].n74 VGND 0.04199f
C8468 XThR.Tn[9].n75 VGND 0.0295f
C8469 XThR.Tn[9].n77 VGND 0.09466f
C8470 XThR.Tn[9].t49 VGND 0.01509f
C8471 XThR.Tn[9].t63 VGND 0.01653f
C8472 XThR.Tn[9].n78 VGND 0.04036f
C8473 XThR.Tn[9].t68 VGND 0.01504f
C8474 XThR.Tn[9].t54 VGND 0.01647f
C8475 XThR.Tn[9].n79 VGND 0.04199f
C8476 XThR.Tn[9].n80 VGND 0.0295f
C8477 XThR.Tn[9].n82 VGND 0.09466f
C8478 XThR.Tn[9].n83 VGND 0.08603f
C8479 XThR.Tn[9].n84 VGND 0.27907f
C8480 XThR.Tn[9].t10 VGND 0.01931f
C8481 XThR.Tn[9].t8 VGND 0.01931f
C8482 XThR.Tn[9].n85 VGND 0.04172f
C8483 XThR.Tn[9].t11 VGND 0.01931f
C8484 XThR.Tn[9].t9 VGND 0.01931f
C8485 XThR.Tn[9].n86 VGND 0.0635f
C8486 XThR.Tn[9].n87 VGND 0.17633f
C8487 XThR.Tn[9].n88 VGND 0.02361f
C8488 XThC.Tn[6].t7 VGND 0.01221f
C8489 XThC.Tn[6].t6 VGND 0.01221f
C8490 XThC.Tn[6].n0 VGND 0.02464f
C8491 XThC.Tn[6].t5 VGND 0.01221f
C8492 XThC.Tn[6].t4 VGND 0.01221f
C8493 XThC.Tn[6].n1 VGND 0.02883f
C8494 XThC.Tn[6].n2 VGND 0.0807f
C8495 XThC.Tn[6].n3 VGND 0.01807f
C8496 XThC.Tn[6].n4 VGND 0.01807f
C8497 XThC.Tn[6].n5 VGND 0.01807f
C8498 XThC.Tn[6].n6 VGND 0.0301f
C8499 XThC.Tn[6].n7 VGND 0.08604f
C8500 XThC.Tn[6].n8 VGND 0.05319f
C8501 XThC.Tn[6].n9 VGND 0.06003f
C8502 XThC.Tn[6].t26 VGND 0.01057f
C8503 XThC.Tn[6].n10 VGND 0.0236f
C8504 XThC.Tn[6].n11 VGND 0.01349f
C8505 XThC.Tn[6].n12 VGND 0.0164f
C8506 XThC.Tn[6].t13 VGND 0.01057f
C8507 XThC.Tn[6].n13 VGND 0.0236f
C8508 XThC.Tn[6].n14 VGND 0.01349f
C8509 XThC.Tn[6].n15 VGND 0.07792f
C8510 XThC.Tn[6].t17 VGND 0.01057f
C8511 XThC.Tn[6].n16 VGND 0.0236f
C8512 XThC.Tn[6].n17 VGND 0.01349f
C8513 XThC.Tn[6].n18 VGND 0.07792f
C8514 XThC.Tn[6].t18 VGND 0.01057f
C8515 XThC.Tn[6].n19 VGND 0.0236f
C8516 XThC.Tn[6].n20 VGND 0.01349f
C8517 XThC.Tn[6].n21 VGND 0.07792f
C8518 XThC.Tn[6].t37 VGND 0.01057f
C8519 XThC.Tn[6].n22 VGND 0.0236f
C8520 XThC.Tn[6].n23 VGND 0.01349f
C8521 XThC.Tn[6].n24 VGND 0.07792f
C8522 XThC.Tn[6].t38 VGND 0.01057f
C8523 XThC.Tn[6].n25 VGND 0.0236f
C8524 XThC.Tn[6].n26 VGND 0.01349f
C8525 XThC.Tn[6].n27 VGND 0.07792f
C8526 XThC.Tn[6].t22 VGND 0.01057f
C8527 XThC.Tn[6].n28 VGND 0.0236f
C8528 XThC.Tn[6].n29 VGND 0.01349f
C8529 XThC.Tn[6].n30 VGND 0.07792f
C8530 XThC.Tn[6].t29 VGND 0.01057f
C8531 XThC.Tn[6].n31 VGND 0.0236f
C8532 XThC.Tn[6].n32 VGND 0.01349f
C8533 XThC.Tn[6].n33 VGND 0.07792f
C8534 XThC.Tn[6].t31 VGND 0.01057f
C8535 XThC.Tn[6].n34 VGND 0.0236f
C8536 XThC.Tn[6].n35 VGND 0.01349f
C8537 XThC.Tn[6].n36 VGND 0.07792f
C8538 XThC.Tn[6].t19 VGND 0.01057f
C8539 XThC.Tn[6].n37 VGND 0.0236f
C8540 XThC.Tn[6].n38 VGND 0.01349f
C8541 XThC.Tn[6].n39 VGND 0.07792f
C8542 XThC.Tn[6].t21 VGND 0.01057f
C8543 XThC.Tn[6].n40 VGND 0.0236f
C8544 XThC.Tn[6].n41 VGND 0.01349f
C8545 XThC.Tn[6].n42 VGND 0.07792f
C8546 XThC.Tn[6].t32 VGND 0.01057f
C8547 XThC.Tn[6].n43 VGND 0.0236f
C8548 XThC.Tn[6].n44 VGND 0.01349f
C8549 XThC.Tn[6].n45 VGND 0.07792f
C8550 XThC.Tn[6].t41 VGND 0.01057f
C8551 XThC.Tn[6].n46 VGND 0.0236f
C8552 XThC.Tn[6].n47 VGND 0.01349f
C8553 XThC.Tn[6].n48 VGND 0.07792f
C8554 XThC.Tn[6].t43 VGND 0.01057f
C8555 XThC.Tn[6].n49 VGND 0.0236f
C8556 XThC.Tn[6].n50 VGND 0.01349f
C8557 XThC.Tn[6].n51 VGND 0.07792f
C8558 XThC.Tn[6].t24 VGND 0.01057f
C8559 XThC.Tn[6].n52 VGND 0.0236f
C8560 XThC.Tn[6].n53 VGND 0.01349f
C8561 XThC.Tn[6].n54 VGND 0.07792f
C8562 XThC.Tn[6].t34 VGND 0.01057f
C8563 XThC.Tn[6].n55 VGND 0.0236f
C8564 XThC.Tn[6].n56 VGND 0.01349f
C8565 XThC.Tn[6].n57 VGND 0.07792f
C8566 XThC.Tn[6].n58 VGND 0.20284f
C8567 XThC.Tn[6].n59 VGND 0.04609f
C8568 XThC.Tn[6].n60 VGND 0.02554f
C8569 XThC.XTBN.Y.n0 VGND 0.01531f
C8570 XThC.XTBN.Y.t50 VGND 0.01024f
C8571 XThC.XTBN.Y.t18 VGND 0.01024f
C8572 XThC.XTBN.Y.n1 VGND 0.01477f
C8573 XThC.XTBN.Y.t120 VGND 0.01024f
C8574 XThC.XTBN.Y.t114 VGND 0.01024f
C8575 XThC.XTBN.Y.n3 VGND 0.0138f
C8576 XThC.XTBN.Y.n5 VGND 0.01477f
C8577 XThC.XTBN.Y.n10 VGND 0.02164f
C8578 XThC.XTBN.Y.t79 VGND 0.01024f
C8579 XThC.XTBN.Y.t36 VGND 0.01024f
C8580 XThC.XTBN.Y.n13 VGND 0.01477f
C8581 XThC.XTBN.Y.t26 VGND 0.01024f
C8582 XThC.XTBN.Y.t21 VGND 0.01024f
C8583 XThC.XTBN.Y.n15 VGND 0.0138f
C8584 XThC.XTBN.Y.n17 VGND 0.01477f
C8585 XThC.XTBN.Y.n22 VGND 0.02164f
C8586 XThC.XTBN.Y.n25 VGND 0.11789f
C8587 XThC.XTBN.Y.t106 VGND 0.01024f
C8588 XThC.XTBN.Y.t70 VGND 0.01024f
C8589 XThC.XTBN.Y.n26 VGND 0.01477f
C8590 XThC.XTBN.Y.t56 VGND 0.01024f
C8591 XThC.XTBN.Y.t48 VGND 0.01024f
C8592 XThC.XTBN.Y.n28 VGND 0.0138f
C8593 XThC.XTBN.Y.n30 VGND 0.01477f
C8594 XThC.XTBN.Y.n35 VGND 0.02164f
C8595 XThC.XTBN.Y.n38 VGND 0.07443f
C8596 XThC.XTBN.Y.t39 VGND 0.01024f
C8597 XThC.XTBN.Y.t122 VGND 0.01024f
C8598 XThC.XTBN.Y.n39 VGND 0.01477f
C8599 XThC.XTBN.Y.t109 VGND 0.01024f
C8600 XThC.XTBN.Y.t102 VGND 0.01024f
C8601 XThC.XTBN.Y.n41 VGND 0.0138f
C8602 XThC.XTBN.Y.n43 VGND 0.01477f
C8603 XThC.XTBN.Y.n48 VGND 0.02164f
C8604 XThC.XTBN.Y.n51 VGND 0.07443f
C8605 XThC.XTBN.Y.t47 VGND 0.01024f
C8606 XThC.XTBN.Y.t17 VGND 0.01024f
C8607 XThC.XTBN.Y.n52 VGND 0.01477f
C8608 XThC.XTBN.Y.t116 VGND 0.01024f
C8609 XThC.XTBN.Y.t111 VGND 0.01024f
C8610 XThC.XTBN.Y.n54 VGND 0.0138f
C8611 XThC.XTBN.Y.n56 VGND 0.01477f
C8612 XThC.XTBN.Y.n61 VGND 0.02164f
C8613 XThC.XTBN.Y.n64 VGND 0.07443f
C8614 XThC.XTBN.Y.t101 VGND 0.01024f
C8615 XThC.XTBN.Y.t63 VGND 0.01024f
C8616 XThC.XTBN.Y.n65 VGND 0.01477f
C8617 XThC.XTBN.Y.t52 VGND 0.01024f
C8618 XThC.XTBN.Y.t44 VGND 0.01024f
C8619 XThC.XTBN.Y.n67 VGND 0.0138f
C8620 XThC.XTBN.Y.n69 VGND 0.01477f
C8621 XThC.XTBN.Y.n74 VGND 0.02164f
C8622 XThC.XTBN.Y.n77 VGND 0.07443f
C8623 XThC.XTBN.Y.t25 VGND 0.01024f
C8624 XThC.XTBN.Y.t100 VGND 0.01024f
C8625 XThC.XTBN.Y.n78 VGND 0.01477f
C8626 XThC.XTBN.Y.t93 VGND 0.01024f
C8627 XThC.XTBN.Y.t90 VGND 0.01024f
C8628 XThC.XTBN.Y.n80 VGND 0.0138f
C8629 XThC.XTBN.Y.n82 VGND 0.01477f
C8630 XThC.XTBN.Y.n87 VGND 0.02164f
C8631 XThC.XTBN.Y.n90 VGND 0.06646f
C8632 XThC.XTBN.Y.t46 VGND 0.01024f
C8633 XThC.XTBN.Y.t6 VGND 0.01024f
C8634 XThC.XTBN.Y.n92 VGND 0.01243f
C8635 XThC.XTBN.Y.t12 VGND 0.01024f
C8636 XThC.XTBN.Y.n93 VGND 0.01348f
C8637 XThC.XTBN.Y.n95 VGND 0.01252f
C8638 XThC.XTBN.Y.n98 VGND 0.01348f
C8639 XThC.XTBN.Y.t54 VGND 0.01024f
C8640 XThC.XTBN.Y.n99 VGND 0.01227f
C8641 XThC.XTBN.Y.n101 VGND 0.01009f
C8642 XThC.XTBN.Y.t38 VGND 0.01024f
C8643 XThC.XTBN.Y.t113 VGND 0.01024f
C8644 XThC.XTBN.Y.n103 VGND 0.01243f
C8645 XThC.XTBN.Y.t119 VGND 0.01024f
C8646 XThC.XTBN.Y.n104 VGND 0.01348f
C8647 XThC.XTBN.Y.n106 VGND 0.01252f
C8648 XThC.XTBN.Y.n109 VGND 0.01348f
C8649 XThC.XTBN.Y.t42 VGND 0.01024f
C8650 XThC.XTBN.Y.n110 VGND 0.01227f
C8651 XThC.XTBN.Y.n113 VGND 0.11256f
C8652 XThC.XTBN.Y.t30 VGND 0.01024f
C8653 XThC.XTBN.Y.t98 VGND 0.01024f
C8654 XThC.XTBN.Y.n115 VGND 0.01243f
C8655 XThC.XTBN.Y.t103 VGND 0.01024f
C8656 XThC.XTBN.Y.n116 VGND 0.01348f
C8657 XThC.XTBN.Y.n118 VGND 0.01252f
C8658 XThC.XTBN.Y.n121 VGND 0.01348f
C8659 XThC.XTBN.Y.t34 VGND 0.01024f
C8660 XThC.XTBN.Y.n122 VGND 0.01227f
C8661 XThC.XTBN.Y.n125 VGND 0.07521f
C8662 XThC.XTBN.Y.t96 VGND 0.01024f
C8663 XThC.XTBN.Y.t51 VGND 0.01024f
C8664 XThC.XTBN.Y.n127 VGND 0.01243f
C8665 XThC.XTBN.Y.t58 VGND 0.01024f
C8666 XThC.XTBN.Y.n128 VGND 0.01348f
C8667 XThC.XTBN.Y.n130 VGND 0.01252f
C8668 XThC.XTBN.Y.n133 VGND 0.01348f
C8669 XThC.XTBN.Y.t99 VGND 0.01024f
C8670 XThC.XTBN.Y.n134 VGND 0.01227f
C8671 XThC.XTBN.Y.n137 VGND 0.07521f
C8672 XThC.XTBN.Y.t88 VGND 0.01024f
C8673 XThC.XTBN.Y.t37 VGND 0.01024f
C8674 XThC.XTBN.Y.n139 VGND 0.01243f
C8675 XThC.XTBN.Y.t40 VGND 0.01024f
C8676 XThC.XTBN.Y.n140 VGND 0.01348f
C8677 XThC.XTBN.Y.n142 VGND 0.01252f
C8678 XThC.XTBN.Y.n145 VGND 0.01348f
C8679 XThC.XTBN.Y.t91 VGND 0.01024f
C8680 XThC.XTBN.Y.n146 VGND 0.01227f
C8681 XThC.XTBN.Y.n149 VGND 0.07534f
C8682 XThC.XTBN.Y.t7 VGND 0.01024f
C8683 XThC.XTBN.Y.t81 VGND 0.01024f
C8684 XThC.XTBN.Y.n151 VGND 0.01243f
C8685 XThC.XTBN.Y.t86 VGND 0.01024f
C8686 XThC.XTBN.Y.n152 VGND 0.01348f
C8687 XThC.XTBN.Y.n154 VGND 0.01252f
C8688 XThC.XTBN.Y.n157 VGND 0.01348f
C8689 XThC.XTBN.Y.t13 VGND 0.01024f
C8690 XThC.XTBN.Y.n158 VGND 0.01227f
C8691 XThC.XTBN.Y.n161 VGND 0.07521f
C8692 XThC.XTBN.Y.t23 VGND 0.01024f
C8693 XThC.XTBN.Y.t95 VGND 0.01024f
C8694 XThC.XTBN.Y.n163 VGND 0.01243f
C8695 XThC.XTBN.Y.t97 VGND 0.01024f
C8696 XThC.XTBN.Y.n164 VGND 0.01348f
C8697 XThC.XTBN.Y.n166 VGND 0.01252f
C8698 XThC.XTBN.Y.n169 VGND 0.01348f
C8699 XThC.XTBN.Y.t28 VGND 0.01024f
C8700 XThC.XTBN.Y.n170 VGND 0.01227f
C8701 XThC.XTBN.Y.n173 VGND 0.08751f
C8702 XThC.XTBN.Y.n174 VGND 0.11019f
C8703 XThC.XTBN.Y.t75 VGND 0.01024f
C8704 XThC.XTBN.Y.t33 VGND 0.01024f
C8705 XThC.XTBN.Y.n175 VGND 0.01477f
C8706 XThC.XTBN.Y.t27 VGND 0.01024f
C8707 XThC.XTBN.Y.n176 VGND 0.02293f
C8708 XThC.XTBN.Y.n181 VGND 0.01477f
C8709 XThC.XTBN.Y.t9 VGND 0.01024f
C8710 XThC.XTBN.Y.n182 VGND 0.0138f
C8711 XThC.XTBN.Y.n186 VGND 0.11129f
C8712 XThC.XTBN.Y.n187 VGND 0.02169f
C8713 XThC.XTBN.Y.n188 VGND 0.01513f
C8714 XThC.XTBN.Y.n189 VGND 0.0307f
C8715 XThR.Tn[12].t0 VGND 0.01931f
C8716 XThR.Tn[12].t2 VGND 0.01931f
C8717 XThR.Tn[12].n0 VGND 0.04293f
C8718 XThR.Tn[12].t3 VGND 0.01931f
C8719 XThR.Tn[12].t1 VGND 0.01931f
C8720 XThR.Tn[12].n1 VGND 0.05864f
C8721 XThR.Tn[12].n2 VGND 0.1952f
C8722 XThR.Tn[12].t7 VGND 0.01255f
C8723 XThR.Tn[12].t5 VGND 0.01255f
C8724 XThR.Tn[12].n3 VGND 0.03131f
C8725 XThR.Tn[12].t6 VGND 0.01255f
C8726 XThR.Tn[12].t4 VGND 0.01255f
C8727 XThR.Tn[12].n4 VGND 0.0251f
C8728 XThR.Tn[12].n5 VGND 0.05789f
C8729 XThR.Tn[12].t36 VGND 0.01509f
C8730 XThR.Tn[12].t28 VGND 0.01653f
C8731 XThR.Tn[12].n6 VGND 0.04036f
C8732 XThR.Tn[12].n7 VGND 0.07753f
C8733 XThR.Tn[12].t53 VGND 0.01509f
C8734 XThR.Tn[12].t43 VGND 0.01653f
C8735 XThR.Tn[12].n8 VGND 0.04036f
C8736 XThR.Tn[12].t71 VGND 0.01504f
C8737 XThR.Tn[12].t21 VGND 0.01647f
C8738 XThR.Tn[12].n9 VGND 0.04199f
C8739 XThR.Tn[12].n10 VGND 0.0295f
C8740 XThR.Tn[12].n12 VGND 0.09466f
C8741 XThR.Tn[12].t30 VGND 0.01509f
C8742 XThR.Tn[12].t20 VGND 0.01653f
C8743 XThR.Tn[12].n13 VGND 0.04036f
C8744 XThR.Tn[12].t49 VGND 0.01504f
C8745 XThR.Tn[12].t60 VGND 0.01647f
C8746 XThR.Tn[12].n14 VGND 0.04199f
C8747 XThR.Tn[12].n15 VGND 0.0295f
C8748 XThR.Tn[12].n17 VGND 0.09466f
C8749 XThR.Tn[12].t45 VGND 0.01509f
C8750 XThR.Tn[12].t38 VGND 0.01653f
C8751 XThR.Tn[12].n18 VGND 0.04036f
C8752 XThR.Tn[12].t63 VGND 0.01504f
C8753 XThR.Tn[12].t15 VGND 0.01647f
C8754 XThR.Tn[12].n19 VGND 0.04199f
C8755 XThR.Tn[12].n20 VGND 0.0295f
C8756 XThR.Tn[12].n22 VGND 0.09466f
C8757 XThR.Tn[12].t70 VGND 0.01509f
C8758 XThR.Tn[12].t66 VGND 0.01653f
C8759 XThR.Tn[12].n23 VGND 0.04036f
C8760 XThR.Tn[12].t33 VGND 0.01504f
C8761 XThR.Tn[12].t46 VGND 0.01647f
C8762 XThR.Tn[12].n24 VGND 0.04199f
C8763 XThR.Tn[12].n25 VGND 0.0295f
C8764 XThR.Tn[12].n27 VGND 0.09466f
C8765 XThR.Tn[12].t48 VGND 0.01509f
C8766 XThR.Tn[12].t39 VGND 0.01653f
C8767 XThR.Tn[12].n28 VGND 0.04036f
C8768 XThR.Tn[12].t64 VGND 0.01504f
C8769 XThR.Tn[12].t17 VGND 0.01647f
C8770 XThR.Tn[12].n29 VGND 0.04199f
C8771 XThR.Tn[12].n30 VGND 0.0295f
C8772 XThR.Tn[12].n32 VGND 0.09466f
C8773 XThR.Tn[12].t23 VGND 0.01509f
C8774 XThR.Tn[12].t56 VGND 0.01653f
C8775 XThR.Tn[12].n33 VGND 0.04036f
C8776 XThR.Tn[12].t41 VGND 0.01504f
C8777 XThR.Tn[12].t37 VGND 0.01647f
C8778 XThR.Tn[12].n34 VGND 0.04199f
C8779 XThR.Tn[12].n35 VGND 0.0295f
C8780 XThR.Tn[12].n37 VGND 0.09466f
C8781 XThR.Tn[12].t54 VGND 0.01509f
C8782 XThR.Tn[12].t51 VGND 0.01653f
C8783 XThR.Tn[12].n38 VGND 0.04036f
C8784 XThR.Tn[12].t72 VGND 0.01504f
C8785 XThR.Tn[12].t29 VGND 0.01647f
C8786 XThR.Tn[12].n39 VGND 0.04199f
C8787 XThR.Tn[12].n40 VGND 0.0295f
C8788 XThR.Tn[12].n42 VGND 0.09466f
C8789 XThR.Tn[12].t59 VGND 0.01509f
C8790 XThR.Tn[12].t65 VGND 0.01653f
C8791 XThR.Tn[12].n43 VGND 0.04036f
C8792 XThR.Tn[12].t14 VGND 0.01504f
C8793 XThR.Tn[12].t44 VGND 0.01647f
C8794 XThR.Tn[12].n44 VGND 0.04199f
C8795 XThR.Tn[12].n45 VGND 0.0295f
C8796 XThR.Tn[12].n47 VGND 0.09466f
C8797 XThR.Tn[12].t12 VGND 0.01509f
C8798 XThR.Tn[12].t22 VGND 0.01653f
C8799 XThR.Tn[12].n48 VGND 0.04036f
C8800 XThR.Tn[12].t35 VGND 0.01504f
C8801 XThR.Tn[12].t61 VGND 0.01647f
C8802 XThR.Tn[12].n49 VGND 0.04199f
C8803 XThR.Tn[12].n50 VGND 0.0295f
C8804 XThR.Tn[12].n52 VGND 0.09466f
C8805 XThR.Tn[12].t68 VGND 0.01509f
C8806 XThR.Tn[12].t40 VGND 0.01653f
C8807 XThR.Tn[12].n53 VGND 0.04036f
C8808 XThR.Tn[12].t26 VGND 0.01504f
C8809 XThR.Tn[12].t19 VGND 0.01647f
C8810 XThR.Tn[12].n54 VGND 0.04199f
C8811 XThR.Tn[12].n55 VGND 0.0295f
C8812 XThR.Tn[12].n57 VGND 0.09466f
C8813 XThR.Tn[12].t25 VGND 0.01509f
C8814 XThR.Tn[12].t16 VGND 0.01653f
C8815 XThR.Tn[12].n58 VGND 0.04036f
C8816 XThR.Tn[12].t42 VGND 0.01504f
C8817 XThR.Tn[12].t55 VGND 0.01647f
C8818 XThR.Tn[12].n59 VGND 0.04199f
C8819 XThR.Tn[12].n60 VGND 0.0295f
C8820 XThR.Tn[12].n62 VGND 0.09466f
C8821 XThR.Tn[12].t57 VGND 0.01509f
C8822 XThR.Tn[12].t52 VGND 0.01653f
C8823 XThR.Tn[12].n63 VGND 0.04036f
C8824 XThR.Tn[12].t13 VGND 0.01504f
C8825 XThR.Tn[12].t31 VGND 0.01647f
C8826 XThR.Tn[12].n64 VGND 0.04199f
C8827 XThR.Tn[12].n65 VGND 0.0295f
C8828 XThR.Tn[12].n67 VGND 0.09466f
C8829 XThR.Tn[12].t73 VGND 0.01509f
C8830 XThR.Tn[12].t67 VGND 0.01653f
C8831 XThR.Tn[12].n68 VGND 0.04036f
C8832 XThR.Tn[12].t34 VGND 0.01504f
C8833 XThR.Tn[12].t47 VGND 0.01647f
C8834 XThR.Tn[12].n69 VGND 0.04199f
C8835 XThR.Tn[12].n70 VGND 0.0295f
C8836 XThR.Tn[12].n72 VGND 0.09466f
C8837 XThR.Tn[12].t32 VGND 0.01509f
C8838 XThR.Tn[12].t24 VGND 0.01653f
C8839 XThR.Tn[12].n73 VGND 0.04036f
C8840 XThR.Tn[12].t50 VGND 0.01504f
C8841 XThR.Tn[12].t62 VGND 0.01647f
C8842 XThR.Tn[12].n74 VGND 0.04199f
C8843 XThR.Tn[12].n75 VGND 0.0295f
C8844 XThR.Tn[12].n77 VGND 0.09466f
C8845 XThR.Tn[12].t69 VGND 0.01509f
C8846 XThR.Tn[12].t18 VGND 0.01653f
C8847 XThR.Tn[12].n78 VGND 0.04036f
C8848 XThR.Tn[12].t27 VGND 0.01504f
C8849 XThR.Tn[12].t58 VGND 0.01647f
C8850 XThR.Tn[12].n79 VGND 0.04199f
C8851 XThR.Tn[12].n80 VGND 0.0295f
C8852 XThR.Tn[12].n82 VGND 0.09466f
C8853 XThR.Tn[12].n83 VGND 0.08603f
C8854 XThR.Tn[12].n84 VGND 0.29341f
C8855 XThR.Tn[12].t10 VGND 0.01931f
C8856 XThR.Tn[12].t8 VGND 0.01931f
C8857 XThR.Tn[12].n85 VGND 0.04172f
C8858 XThR.Tn[12].t11 VGND 0.01931f
C8859 XThR.Tn[12].t9 VGND 0.01931f
C8860 XThR.Tn[12].n86 VGND 0.06351f
C8861 XThR.Tn[12].n87 VGND 0.17633f
C8862 XThR.Tn[14].t0 VGND 0.0197f
C8863 XThR.Tn[14].t1 VGND 0.0197f
C8864 XThR.Tn[14].n0 VGND 0.0598f
C8865 XThR.Tn[14].t2 VGND 0.0197f
C8866 XThR.Tn[14].t3 VGND 0.0197f
C8867 XThR.Tn[14].n1 VGND 0.04378f
C8868 XThR.Tn[14].n2 VGND 0.19909f
C8869 XThR.Tn[14].t6 VGND 0.0128f
C8870 XThR.Tn[14].t7 VGND 0.0128f
C8871 XThR.Tn[14].n3 VGND 0.03193f
C8872 XThR.Tn[14].t4 VGND 0.0128f
C8873 XThR.Tn[14].t5 VGND 0.0128f
C8874 XThR.Tn[14].n4 VGND 0.02561f
C8875 XThR.Tn[14].n5 VGND 0.05904f
C8876 XThR.Tn[14].t69 VGND 0.01539f
C8877 XThR.Tn[14].t62 VGND 0.01686f
C8878 XThR.Tn[14].n6 VGND 0.04116f
C8879 XThR.Tn[14].n7 VGND 0.07907f
C8880 XThR.Tn[14].t24 VGND 0.01539f
C8881 XThR.Tn[14].t13 VGND 0.01686f
C8882 XThR.Tn[14].n8 VGND 0.04116f
C8883 XThR.Tn[14].t28 VGND 0.01534f
C8884 XThR.Tn[14].t60 VGND 0.0168f
C8885 XThR.Tn[14].n9 VGND 0.04283f
C8886 XThR.Tn[14].n10 VGND 0.03009f
C8887 XThR.Tn[14].n12 VGND 0.09655f
C8888 XThR.Tn[14].t64 VGND 0.01539f
C8889 XThR.Tn[14].t54 VGND 0.01686f
C8890 XThR.Tn[14].n13 VGND 0.04116f
C8891 XThR.Tn[14].t67 VGND 0.01534f
C8892 XThR.Tn[14].t34 VGND 0.0168f
C8893 XThR.Tn[14].n14 VGND 0.04283f
C8894 XThR.Tn[14].n15 VGND 0.03009f
C8895 XThR.Tn[14].n17 VGND 0.09655f
C8896 XThR.Tn[14].t14 VGND 0.01539f
C8897 XThR.Tn[14].t72 VGND 0.01686f
C8898 XThR.Tn[14].n18 VGND 0.04116f
C8899 XThR.Tn[14].t17 VGND 0.01534f
C8900 XThR.Tn[14].t52 VGND 0.0168f
C8901 XThR.Tn[14].n19 VGND 0.04283f
C8902 XThR.Tn[14].n20 VGND 0.03009f
C8903 XThR.Tn[14].n22 VGND 0.09655f
C8904 XThR.Tn[14].t44 VGND 0.01539f
C8905 XThR.Tn[14].t38 VGND 0.01686f
C8906 XThR.Tn[14].n23 VGND 0.04116f
C8907 XThR.Tn[14].t47 VGND 0.01534f
C8908 XThR.Tn[14].t18 VGND 0.0168f
C8909 XThR.Tn[14].n24 VGND 0.04283f
C8910 XThR.Tn[14].n25 VGND 0.03009f
C8911 XThR.Tn[14].n27 VGND 0.09655f
C8912 XThR.Tn[14].t15 VGND 0.01539f
C8913 XThR.Tn[14].t73 VGND 0.01686f
C8914 XThR.Tn[14].n28 VGND 0.04116f
C8915 XThR.Tn[14].t21 VGND 0.01534f
C8916 XThR.Tn[14].t53 VGND 0.0168f
C8917 XThR.Tn[14].n29 VGND 0.04283f
C8918 XThR.Tn[14].n30 VGND 0.03009f
C8919 XThR.Tn[14].n32 VGND 0.09655f
C8920 XThR.Tn[14].t57 VGND 0.01539f
C8921 XThR.Tn[14].t25 VGND 0.01686f
C8922 XThR.Tn[14].n33 VGND 0.04116f
C8923 XThR.Tn[14].t61 VGND 0.01534f
C8924 XThR.Tn[14].t71 VGND 0.0168f
C8925 XThR.Tn[14].n34 VGND 0.04283f
C8926 XThR.Tn[14].n35 VGND 0.03009f
C8927 XThR.Tn[14].n37 VGND 0.09655f
C8928 XThR.Tn[14].t23 VGND 0.01539f
C8929 XThR.Tn[14].t19 VGND 0.01686f
C8930 XThR.Tn[14].n38 VGND 0.04116f
C8931 XThR.Tn[14].t29 VGND 0.01534f
C8932 XThR.Tn[14].t66 VGND 0.0168f
C8933 XThR.Tn[14].n39 VGND 0.04283f
C8934 XThR.Tn[14].n40 VGND 0.03009f
C8935 XThR.Tn[14].n42 VGND 0.09655f
C8936 XThR.Tn[14].t27 VGND 0.01539f
C8937 XThR.Tn[14].t36 VGND 0.01686f
C8938 XThR.Tn[14].n43 VGND 0.04116f
C8939 XThR.Tn[14].t33 VGND 0.01534f
C8940 XThR.Tn[14].t16 VGND 0.0168f
C8941 XThR.Tn[14].n44 VGND 0.04283f
C8942 XThR.Tn[14].n45 VGND 0.03009f
C8943 XThR.Tn[14].n47 VGND 0.09655f
C8944 XThR.Tn[14].t46 VGND 0.01539f
C8945 XThR.Tn[14].t56 VGND 0.01686f
C8946 XThR.Tn[14].n48 VGND 0.04116f
C8947 XThR.Tn[14].t50 VGND 0.01534f
C8948 XThR.Tn[14].t35 VGND 0.0168f
C8949 XThR.Tn[14].n49 VGND 0.04283f
C8950 XThR.Tn[14].n50 VGND 0.03009f
C8951 XThR.Tn[14].n52 VGND 0.09655f
C8952 XThR.Tn[14].t40 VGND 0.01539f
C8953 XThR.Tn[14].t12 VGND 0.01686f
C8954 XThR.Tn[14].n53 VGND 0.04116f
C8955 XThR.Tn[14].t42 VGND 0.01534f
C8956 XThR.Tn[14].t55 VGND 0.0168f
C8957 XThR.Tn[14].n54 VGND 0.04283f
C8958 XThR.Tn[14].n55 VGND 0.03009f
C8959 XThR.Tn[14].n57 VGND 0.09655f
C8960 XThR.Tn[14].t59 VGND 0.01539f
C8961 XThR.Tn[14].t49 VGND 0.01686f
C8962 XThR.Tn[14].n58 VGND 0.04116f
C8963 XThR.Tn[14].t63 VGND 0.01534f
C8964 XThR.Tn[14].t30 VGND 0.0168f
C8965 XThR.Tn[14].n59 VGND 0.04283f
C8966 XThR.Tn[14].n60 VGND 0.03009f
C8967 XThR.Tn[14].n62 VGND 0.09655f
C8968 XThR.Tn[14].t26 VGND 0.01539f
C8969 XThR.Tn[14].t22 VGND 0.01686f
C8970 XThR.Tn[14].n63 VGND 0.04116f
C8971 XThR.Tn[14].t31 VGND 0.01534f
C8972 XThR.Tn[14].t68 VGND 0.0168f
C8973 XThR.Tn[14].n64 VGND 0.04283f
C8974 XThR.Tn[14].n65 VGND 0.03009f
C8975 XThR.Tn[14].n67 VGND 0.09655f
C8976 XThR.Tn[14].t45 VGND 0.01539f
C8977 XThR.Tn[14].t39 VGND 0.01686f
C8978 XThR.Tn[14].n68 VGND 0.04116f
C8979 XThR.Tn[14].t48 VGND 0.01534f
C8980 XThR.Tn[14].t20 VGND 0.0168f
C8981 XThR.Tn[14].n69 VGND 0.04283f
C8982 XThR.Tn[14].n70 VGND 0.03009f
C8983 XThR.Tn[14].n72 VGND 0.09655f
C8984 XThR.Tn[14].t65 VGND 0.01539f
C8985 XThR.Tn[14].t58 VGND 0.01686f
C8986 XThR.Tn[14].n73 VGND 0.04116f
C8987 XThR.Tn[14].t70 VGND 0.01534f
C8988 XThR.Tn[14].t37 VGND 0.0168f
C8989 XThR.Tn[14].n74 VGND 0.04283f
C8990 XThR.Tn[14].n75 VGND 0.03009f
C8991 XThR.Tn[14].n77 VGND 0.09655f
C8992 XThR.Tn[14].t41 VGND 0.01539f
C8993 XThR.Tn[14].t51 VGND 0.01686f
C8994 XThR.Tn[14].n78 VGND 0.04116f
C8995 XThR.Tn[14].t43 VGND 0.01534f
C8996 XThR.Tn[14].t32 VGND 0.0168f
C8997 XThR.Tn[14].n79 VGND 0.04283f
C8998 XThR.Tn[14].n80 VGND 0.03009f
C8999 XThR.Tn[14].n82 VGND 0.09655f
C9000 XThR.Tn[14].n83 VGND 0.08774f
C9001 XThR.Tn[14].n84 VGND 0.35247f
C9002 XThR.Tn[14].t10 VGND 0.0197f
C9003 XThR.Tn[14].t11 VGND 0.0197f
C9004 XThR.Tn[14].n85 VGND 0.04256f
C9005 XThR.Tn[14].t8 VGND 0.0197f
C9006 XThR.Tn[14].t9 VGND 0.0197f
C9007 XThR.Tn[14].n86 VGND 0.06477f
C9008 XThR.Tn[14].n87 VGND 0.17985f
C9009 XThR.Tn[6].t2 VGND 0.01813f
C9010 XThR.Tn[6].t1 VGND 0.01813f
C9011 XThR.Tn[6].n0 VGND 0.04282f
C9012 XThR.Tn[6].t3 VGND 0.01813f
C9013 XThR.Tn[6].t0 VGND 0.01813f
C9014 XThR.Tn[6].n1 VGND 0.0366f
C9015 XThR.Tn[6].n2 VGND 0.12845f
C9016 XThR.Tn[6].t8 VGND 0.01179f
C9017 XThR.Tn[6].t9 VGND 0.01179f
C9018 XThR.Tn[6].n3 VGND 0.04472f
C9019 XThR.Tn[6].t11 VGND 0.01179f
C9020 XThR.Tn[6].t10 VGND 0.01179f
C9021 XThR.Tn[6].n4 VGND 0.02684f
C9022 XThR.Tn[6].n5 VGND 0.12781f
C9023 XThR.Tn[6].t7 VGND 0.01179f
C9024 XThR.Tn[6].t6 VGND 0.01179f
C9025 XThR.Tn[6].n6 VGND 0.02684f
C9026 XThR.Tn[6].n7 VGND 0.07901f
C9027 XThR.Tn[6].t4 VGND 0.01179f
C9028 XThR.Tn[6].t5 VGND 0.01179f
C9029 XThR.Tn[6].n8 VGND 0.02684f
C9030 XThR.Tn[6].n9 VGND 0.08917f
C9031 XThR.Tn[6].t62 VGND 0.01417f
C9032 XThR.Tn[6].t56 VGND 0.01552f
C9033 XThR.Tn[6].n10 VGND 0.03789f
C9034 XThR.Tn[6].n11 VGND 0.07279f
C9035 XThR.Tn[6].t20 VGND 0.01417f
C9036 XThR.Tn[6].t72 VGND 0.01552f
C9037 XThR.Tn[6].n12 VGND 0.03789f
C9038 XThR.Tn[6].t36 VGND 0.01412f
C9039 XThR.Tn[6].t68 VGND 0.01547f
C9040 XThR.Tn[6].n13 VGND 0.03943f
C9041 XThR.Tn[6].n14 VGND 0.0277f
C9042 XThR.Tn[6].n16 VGND 0.08888f
C9043 XThR.Tn[6].t57 VGND 0.01417f
C9044 XThR.Tn[6].t49 VGND 0.01552f
C9045 XThR.Tn[6].n17 VGND 0.03789f
C9046 XThR.Tn[6].t14 VGND 0.01412f
C9047 XThR.Tn[6].t45 VGND 0.01547f
C9048 XThR.Tn[6].n18 VGND 0.03943f
C9049 XThR.Tn[6].n19 VGND 0.0277f
C9050 XThR.Tn[6].n21 VGND 0.08888f
C9051 XThR.Tn[6].t73 VGND 0.01417f
C9052 XThR.Tn[6].t66 VGND 0.01552f
C9053 XThR.Tn[6].n22 VGND 0.03789f
C9054 XThR.Tn[6].t26 VGND 0.01412f
C9055 XThR.Tn[6].t63 VGND 0.01547f
C9056 XThR.Tn[6].n23 VGND 0.03943f
C9057 XThR.Tn[6].n24 VGND 0.0277f
C9058 XThR.Tn[6].n26 VGND 0.08888f
C9059 XThR.Tn[6].t35 VGND 0.01417f
C9060 XThR.Tn[6].t31 VGND 0.01552f
C9061 XThR.Tn[6].n27 VGND 0.03789f
C9062 XThR.Tn[6].t59 VGND 0.01412f
C9063 XThR.Tn[6].t27 VGND 0.01547f
C9064 XThR.Tn[6].n28 VGND 0.03943f
C9065 XThR.Tn[6].n29 VGND 0.0277f
C9066 XThR.Tn[6].n31 VGND 0.08888f
C9067 XThR.Tn[6].t13 VGND 0.01417f
C9068 XThR.Tn[6].t67 VGND 0.01552f
C9069 XThR.Tn[6].n32 VGND 0.03789f
C9070 XThR.Tn[6].t29 VGND 0.01412f
C9071 XThR.Tn[6].t64 VGND 0.01547f
C9072 XThR.Tn[6].n33 VGND 0.03943f
C9073 XThR.Tn[6].n34 VGND 0.0277f
C9074 XThR.Tn[6].n36 VGND 0.08888f
C9075 XThR.Tn[6].t51 VGND 0.01417f
C9076 XThR.Tn[6].t22 VGND 0.01552f
C9077 XThR.Tn[6].n37 VGND 0.03789f
C9078 XThR.Tn[6].t70 VGND 0.01412f
C9079 XThR.Tn[6].t19 VGND 0.01547f
C9080 XThR.Tn[6].n38 VGND 0.03943f
C9081 XThR.Tn[6].n39 VGND 0.0277f
C9082 XThR.Tn[6].n41 VGND 0.08888f
C9083 XThR.Tn[6].t21 VGND 0.01417f
C9084 XThR.Tn[6].t17 VGND 0.01552f
C9085 XThR.Tn[6].n42 VGND 0.03789f
C9086 XThR.Tn[6].t37 VGND 0.01412f
C9087 XThR.Tn[6].t12 VGND 0.01547f
C9088 XThR.Tn[6].n43 VGND 0.03943f
C9089 XThR.Tn[6].n44 VGND 0.0277f
C9090 XThR.Tn[6].n46 VGND 0.08888f
C9091 XThR.Tn[6].t24 VGND 0.01417f
C9092 XThR.Tn[6].t30 VGND 0.01552f
C9093 XThR.Tn[6].n47 VGND 0.03789f
C9094 XThR.Tn[6].t43 VGND 0.01412f
C9095 XThR.Tn[6].t25 VGND 0.01547f
C9096 XThR.Tn[6].n48 VGND 0.03943f
C9097 XThR.Tn[6].n49 VGND 0.0277f
C9098 XThR.Tn[6].n51 VGND 0.08888f
C9099 XThR.Tn[6].t40 VGND 0.01417f
C9100 XThR.Tn[6].t50 VGND 0.01552f
C9101 XThR.Tn[6].n52 VGND 0.03789f
C9102 XThR.Tn[6].t61 VGND 0.01412f
C9103 XThR.Tn[6].t47 VGND 0.01547f
C9104 XThR.Tn[6].n53 VGND 0.03943f
C9105 XThR.Tn[6].n54 VGND 0.0277f
C9106 XThR.Tn[6].n56 VGND 0.08888f
C9107 XThR.Tn[6].t33 VGND 0.01417f
C9108 XThR.Tn[6].t69 VGND 0.01552f
C9109 XThR.Tn[6].n57 VGND 0.03789f
C9110 XThR.Tn[6].t54 VGND 0.01412f
C9111 XThR.Tn[6].t65 VGND 0.01547f
C9112 XThR.Tn[6].n58 VGND 0.03943f
C9113 XThR.Tn[6].n59 VGND 0.0277f
C9114 XThR.Tn[6].n61 VGND 0.08888f
C9115 XThR.Tn[6].t53 VGND 0.01417f
C9116 XThR.Tn[6].t44 VGND 0.01552f
C9117 XThR.Tn[6].n62 VGND 0.03789f
C9118 XThR.Tn[6].t71 VGND 0.01412f
C9119 XThR.Tn[6].t39 VGND 0.01547f
C9120 XThR.Tn[6].n63 VGND 0.03943f
C9121 XThR.Tn[6].n64 VGND 0.0277f
C9122 XThR.Tn[6].n66 VGND 0.08888f
C9123 XThR.Tn[6].t23 VGND 0.01417f
C9124 XThR.Tn[6].t18 VGND 0.01552f
C9125 XThR.Tn[6].n67 VGND 0.03789f
C9126 XThR.Tn[6].t41 VGND 0.01412f
C9127 XThR.Tn[6].t15 VGND 0.01547f
C9128 XThR.Tn[6].n68 VGND 0.03943f
C9129 XThR.Tn[6].n69 VGND 0.0277f
C9130 XThR.Tn[6].n71 VGND 0.08888f
C9131 XThR.Tn[6].t38 VGND 0.01417f
C9132 XThR.Tn[6].t32 VGND 0.01552f
C9133 XThR.Tn[6].n72 VGND 0.03789f
C9134 XThR.Tn[6].t60 VGND 0.01412f
C9135 XThR.Tn[6].t28 VGND 0.01547f
C9136 XThR.Tn[6].n73 VGND 0.03943f
C9137 XThR.Tn[6].n74 VGND 0.0277f
C9138 XThR.Tn[6].n76 VGND 0.08888f
C9139 XThR.Tn[6].t58 VGND 0.01417f
C9140 XThR.Tn[6].t52 VGND 0.01552f
C9141 XThR.Tn[6].n77 VGND 0.03789f
C9142 XThR.Tn[6].t16 VGND 0.01412f
C9143 XThR.Tn[6].t48 VGND 0.01547f
C9144 XThR.Tn[6].n78 VGND 0.03943f
C9145 XThR.Tn[6].n79 VGND 0.0277f
C9146 XThR.Tn[6].n81 VGND 0.08888f
C9147 XThR.Tn[6].t34 VGND 0.01417f
C9148 XThR.Tn[6].t46 VGND 0.01552f
C9149 XThR.Tn[6].n82 VGND 0.03789f
C9150 XThR.Tn[6].t55 VGND 0.01412f
C9151 XThR.Tn[6].t42 VGND 0.01547f
C9152 XThR.Tn[6].n83 VGND 0.03943f
C9153 XThR.Tn[6].n84 VGND 0.0277f
C9154 XThR.Tn[6].n86 VGND 0.08888f
C9155 XThR.Tn[6].n87 VGND 0.08078f
C9156 XThR.Tn[6].n88 VGND 0.13446f
C9157 XThR.XTBN.Y.t60 VGND 0.01124f
C9158 XThR.XTBN.Y.n1 VGND 0.01347f
C9159 XThR.XTBN.Y.t12 VGND 0.01124f
C9160 XThR.XTBN.Y.t81 VGND 0.01124f
C9161 XThR.XTBN.Y.n2 VGND 0.01479f
C9162 XThR.XTBN.Y.t121 VGND 0.01124f
C9163 XThR.XTBN.Y.n3 VGND 0.01365f
C9164 XThR.XTBN.Y.n5 VGND 0.01304f
C9165 XThR.XTBN.Y.n8 VGND 0.01479f
C9166 XThR.XTBN.Y.n10 VGND 0.0122f
C9167 XThR.XTBN.Y.t115 VGND 0.01124f
C9168 XThR.XTBN.Y.n12 VGND 0.01347f
C9169 XThR.XTBN.Y.t65 VGND 0.01124f
C9170 XThR.XTBN.Y.t21 VGND 0.01124f
C9171 XThR.XTBN.Y.n13 VGND 0.01479f
C9172 XThR.XTBN.Y.t57 VGND 0.01124f
C9173 XThR.XTBN.Y.n14 VGND 0.01365f
C9174 XThR.XTBN.Y.n16 VGND 0.01304f
C9175 XThR.XTBN.Y.n19 VGND 0.01479f
C9176 XThR.XTBN.Y.n22 VGND 0.12354f
C9177 XThR.XTBN.Y.t27 VGND 0.01124f
C9178 XThR.XTBN.Y.n24 VGND 0.01347f
C9179 XThR.XTBN.Y.t96 VGND 0.01124f
C9180 XThR.XTBN.Y.t46 VGND 0.01124f
C9181 XThR.XTBN.Y.n25 VGND 0.01479f
C9182 XThR.XTBN.Y.t89 VGND 0.01124f
C9183 XThR.XTBN.Y.n26 VGND 0.01365f
C9184 XThR.XTBN.Y.n28 VGND 0.01304f
C9185 XThR.XTBN.Y.n31 VGND 0.01479f
C9186 XThR.XTBN.Y.n34 VGND 0.08255f
C9187 XThR.XTBN.Y.t80 VGND 0.01124f
C9188 XThR.XTBN.Y.n36 VGND 0.01347f
C9189 XThR.XTBN.Y.t31 VGND 0.01124f
C9190 XThR.XTBN.Y.t102 VGND 0.01124f
C9191 XThR.XTBN.Y.n37 VGND 0.01479f
C9192 XThR.XTBN.Y.t25 VGND 0.01124f
C9193 XThR.XTBN.Y.n38 VGND 0.01365f
C9194 XThR.XTBN.Y.n40 VGND 0.01304f
C9195 XThR.XTBN.Y.n43 VGND 0.01479f
C9196 XThR.XTBN.Y.n46 VGND 0.08255f
C9197 XThR.XTBN.Y.t85 VGND 0.01124f
C9198 XThR.XTBN.Y.n48 VGND 0.01347f
C9199 XThR.XTBN.Y.t33 VGND 0.01124f
C9200 XThR.XTBN.Y.t105 VGND 0.01124f
C9201 XThR.XTBN.Y.n49 VGND 0.01479f
C9202 XThR.XTBN.Y.t26 VGND 0.01124f
C9203 XThR.XTBN.Y.n50 VGND 0.01365f
C9204 XThR.XTBN.Y.n52 VGND 0.01304f
C9205 XThR.XTBN.Y.n55 VGND 0.01479f
C9206 XThR.XTBN.Y.n58 VGND 0.08269f
C9207 XThR.XTBN.Y.t54 VGND 0.01124f
C9208 XThR.XTBN.Y.n60 VGND 0.01347f
C9209 XThR.XTBN.Y.t5 VGND 0.01124f
C9210 XThR.XTBN.Y.t73 VGND 0.01124f
C9211 XThR.XTBN.Y.n61 VGND 0.01479f
C9212 XThR.XTBN.Y.t114 VGND 0.01124f
C9213 XThR.XTBN.Y.n62 VGND 0.01365f
C9214 XThR.XTBN.Y.n64 VGND 0.01304f
C9215 XThR.XTBN.Y.n67 VGND 0.01479f
C9216 XThR.XTBN.Y.n70 VGND 0.08255f
C9217 XThR.XTBN.Y.t49 VGND 0.01124f
C9218 XThR.XTBN.Y.n72 VGND 0.01347f
C9219 XThR.XTBN.Y.t119 VGND 0.01124f
C9220 XThR.XTBN.Y.t69 VGND 0.01124f
C9221 XThR.XTBN.Y.n73 VGND 0.01479f
C9222 XThR.XTBN.Y.t108 VGND 0.01124f
C9223 XThR.XTBN.Y.n74 VGND 0.01365f
C9224 XThR.XTBN.Y.n76 VGND 0.01304f
C9225 XThR.XTBN.Y.n79 VGND 0.01479f
C9226 XThR.XTBN.Y.n82 VGND 0.09424f
C9227 XThR.XTBN.Y.t99 VGND 0.01124f
C9228 XThR.XTBN.Y.t87 VGND 0.01124f
C9229 XThR.XTBN.Y.n83 VGND 0.01621f
C9230 XThR.XTBN.Y.t77 VGND 0.01124f
C9231 XThR.XTBN.Y.t68 VGND 0.01124f
C9232 XThR.XTBN.Y.n84 VGND 0.01515f
C9233 XThR.XTBN.Y.n87 VGND 0.01621f
C9234 XThR.XTBN.Y.n92 VGND 0.02375f
C9235 XThR.XTBN.Y.n93 VGND 0.01318f
C9236 XThR.XTBN.Y.t66 VGND 0.01124f
C9237 XThR.XTBN.Y.t23 VGND 0.01124f
C9238 XThR.XTBN.Y.n94 VGND 0.01621f
C9239 XThR.XTBN.Y.t59 VGND 0.01124f
C9240 XThR.XTBN.Y.t97 VGND 0.01124f
C9241 XThR.XTBN.Y.n95 VGND 0.01515f
C9242 XThR.XTBN.Y.n98 VGND 0.01621f
C9243 XThR.XTBN.Y.n103 VGND 0.02375f
C9244 XThR.XTBN.Y.n105 VGND 0.13142f
C9245 XThR.XTBN.Y.t15 VGND 0.01124f
C9246 XThR.XTBN.Y.t83 VGND 0.01124f
C9247 XThR.XTBN.Y.n106 VGND 0.01621f
C9248 XThR.XTBN.Y.t123 VGND 0.01124f
C9249 XThR.XTBN.Y.t39 VGND 0.01124f
C9250 XThR.XTBN.Y.n107 VGND 0.01515f
C9251 XThR.XTBN.Y.n110 VGND 0.01621f
C9252 XThR.XTBN.Y.n115 VGND 0.02375f
C9253 XThR.XTBN.Y.n117 VGND 0.08248f
C9254 XThR.XTBN.Y.t100 VGND 0.01124f
C9255 XThR.XTBN.Y.t50 VGND 0.01124f
C9256 XThR.XTBN.Y.n118 VGND 0.01621f
C9257 XThR.XTBN.Y.t92 VGND 0.01124f
C9258 XThR.XTBN.Y.t13 VGND 0.01124f
C9259 XThR.XTBN.Y.n119 VGND 0.01515f
C9260 XThR.XTBN.Y.n122 VGND 0.01621f
C9261 XThR.XTBN.Y.n127 VGND 0.02375f
C9262 XThR.XTBN.Y.n129 VGND 0.08248f
C9263 XThR.XTBN.Y.t45 VGND 0.01124f
C9264 XThR.XTBN.Y.t117 VGND 0.01124f
C9265 XThR.XTBN.Y.n130 VGND 0.01621f
C9266 XThR.XTBN.Y.t36 VGND 0.01124f
C9267 XThR.XTBN.Y.t75 VGND 0.01124f
C9268 XThR.XTBN.Y.n131 VGND 0.01515f
C9269 XThR.XTBN.Y.n134 VGND 0.01621f
C9270 XThR.XTBN.Y.n139 VGND 0.02375f
C9271 XThR.XTBN.Y.n141 VGND 0.08248f
C9272 XThR.XTBN.Y.t19 VGND 0.01124f
C9273 XThR.XTBN.Y.t86 VGND 0.01124f
C9274 XThR.XTBN.Y.n142 VGND 0.01621f
C9275 XThR.XTBN.Y.t6 VGND 0.01124f
C9276 XThR.XTBN.Y.t43 VGND 0.01124f
C9277 XThR.XTBN.Y.n143 VGND 0.01515f
C9278 XThR.XTBN.Y.n146 VGND 0.01621f
C9279 XThR.XTBN.Y.n151 VGND 0.02375f
C9280 XThR.XTBN.Y.n153 VGND 0.08248f
C9281 XThR.XTBN.Y.t41 VGND 0.01124f
C9282 XThR.XTBN.Y.t113 VGND 0.01124f
C9283 XThR.XTBN.Y.n154 VGND 0.01621f
C9284 XThR.XTBN.Y.t34 VGND 0.01124f
C9285 XThR.XTBN.Y.t72 VGND 0.01124f
C9286 XThR.XTBN.Y.n155 VGND 0.01515f
C9287 XThR.XTBN.Y.n158 VGND 0.01621f
C9288 XThR.XTBN.Y.n163 VGND 0.02375f
C9289 XThR.XTBN.Y.n165 VGND 0.07589f
C9290 XThR.XTBN.Y.n166 VGND 0.12019f
C9291 XThR.XTBN.Y.t106 VGND 0.01124f
C9292 XThR.XTBN.Y.t63 VGND 0.01124f
C9293 XThR.XTBN.Y.n167 VGND 0.01515f
C9294 XThR.XTBN.Y.n169 VGND 0.01621f
C9295 XThR.XTBN.Y.t56 VGND 0.01124f
C9296 XThR.XTBN.Y.t7 VGND 0.01124f
C9297 XThR.XTBN.Y.n170 VGND 0.02517f
C9298 XThR.XTBN.Y.n174 VGND 0.01621f
C9299 XThR.XTBN.Y.n178 VGND 0.12255f
C9300 XThR.XTBN.Y.n179 VGND 0.02242f
C9301 XThR.XTBN.Y.n180 VGND 0.01587f
C9302 XThR.XTBN.Y.n183 VGND 0.0112f
C9303 XThR.XTBN.Y.n184 VGND 0.022f
C9304 XThC.Tn[10].n0 VGND 0.02345f
C9305 XThC.Tn[10].n1 VGND 0.0188f
C9306 XThC.Tn[10].n2 VGND 0.0473f
C9307 XThC.Tn[10].t38 VGND 0.01146f
C9308 XThC.Tn[10].t36 VGND 0.01252f
C9309 XThC.Tn[10].n3 VGND 0.02796f
C9310 XThC.Tn[10].n4 VGND 0.01598f
C9311 XThC.Tn[10].n5 VGND 0.01943f
C9312 XThC.Tn[10].t24 VGND 0.01146f
C9313 XThC.Tn[10].t21 VGND 0.01252f
C9314 XThC.Tn[10].n6 VGND 0.02796f
C9315 XThC.Tn[10].n7 VGND 0.01598f
C9316 XThC.Tn[10].n8 VGND 0.09232f
C9317 XThC.Tn[10].t29 VGND 0.01146f
C9318 XThC.Tn[10].t23 VGND 0.01252f
C9319 XThC.Tn[10].n9 VGND 0.02796f
C9320 XThC.Tn[10].n10 VGND 0.01598f
C9321 XThC.Tn[10].n11 VGND 0.09232f
C9322 XThC.Tn[10].t30 VGND 0.01146f
C9323 XThC.Tn[10].t25 VGND 0.01252f
C9324 XThC.Tn[10].n12 VGND 0.02796f
C9325 XThC.Tn[10].n13 VGND 0.01598f
C9326 XThC.Tn[10].n14 VGND 0.09232f
C9327 XThC.Tn[10].t17 VGND 0.01146f
C9328 XThC.Tn[10].t14 VGND 0.01252f
C9329 XThC.Tn[10].n15 VGND 0.02796f
C9330 XThC.Tn[10].n16 VGND 0.01598f
C9331 XThC.Tn[10].n17 VGND 0.09232f
C9332 XThC.Tn[10].t18 VGND 0.01146f
C9333 XThC.Tn[10].t15 VGND 0.01252f
C9334 XThC.Tn[10].n18 VGND 0.02796f
C9335 XThC.Tn[10].n19 VGND 0.01598f
C9336 XThC.Tn[10].n20 VGND 0.09232f
C9337 XThC.Tn[10].t34 VGND 0.01146f
C9338 XThC.Tn[10].t28 VGND 0.01252f
C9339 XThC.Tn[10].n21 VGND 0.02796f
C9340 XThC.Tn[10].n22 VGND 0.01598f
C9341 XThC.Tn[10].n23 VGND 0.09232f
C9342 XThC.Tn[10].t41 VGND 0.01146f
C9343 XThC.Tn[10].t37 VGND 0.01252f
C9344 XThC.Tn[10].n24 VGND 0.02796f
C9345 XThC.Tn[10].n25 VGND 0.01598f
C9346 XThC.Tn[10].n26 VGND 0.09232f
C9347 XThC.Tn[10].t43 VGND 0.01146f
C9348 XThC.Tn[10].t39 VGND 0.01252f
C9349 XThC.Tn[10].n27 VGND 0.02796f
C9350 XThC.Tn[10].n28 VGND 0.01598f
C9351 XThC.Tn[10].n29 VGND 0.09232f
C9352 XThC.Tn[10].t31 VGND 0.01146f
C9353 XThC.Tn[10].t26 VGND 0.01252f
C9354 XThC.Tn[10].n30 VGND 0.02796f
C9355 XThC.Tn[10].n31 VGND 0.01598f
C9356 XThC.Tn[10].n32 VGND 0.09232f
C9357 XThC.Tn[10].t33 VGND 0.01146f
C9358 XThC.Tn[10].t27 VGND 0.01252f
C9359 XThC.Tn[10].n33 VGND 0.02796f
C9360 XThC.Tn[10].n34 VGND 0.01598f
C9361 XThC.Tn[10].n35 VGND 0.09232f
C9362 XThC.Tn[10].t12 VGND 0.01146f
C9363 XThC.Tn[10].t40 VGND 0.01252f
C9364 XThC.Tn[10].n36 VGND 0.02796f
C9365 XThC.Tn[10].n37 VGND 0.01598f
C9366 XThC.Tn[10].n38 VGND 0.09232f
C9367 XThC.Tn[10].t20 VGND 0.01146f
C9368 XThC.Tn[10].t16 VGND 0.01252f
C9369 XThC.Tn[10].n39 VGND 0.02796f
C9370 XThC.Tn[10].n40 VGND 0.01598f
C9371 XThC.Tn[10].n41 VGND 0.09232f
C9372 XThC.Tn[10].t22 VGND 0.01146f
C9373 XThC.Tn[10].t19 VGND 0.01252f
C9374 XThC.Tn[10].n42 VGND 0.02796f
C9375 XThC.Tn[10].n43 VGND 0.01598f
C9376 XThC.Tn[10].n44 VGND 0.09232f
C9377 XThC.Tn[10].t35 VGND 0.01146f
C9378 XThC.Tn[10].t32 VGND 0.01252f
C9379 XThC.Tn[10].n45 VGND 0.02796f
C9380 XThC.Tn[10].n46 VGND 0.01598f
C9381 XThC.Tn[10].n47 VGND 0.09232f
C9382 XThC.Tn[10].t13 VGND 0.01146f
C9383 XThC.Tn[10].t42 VGND 0.01252f
C9384 XThC.Tn[10].n48 VGND 0.02796f
C9385 XThC.Tn[10].n49 VGND 0.01598f
C9386 XThC.Tn[10].n50 VGND 0.09232f
C9387 XThC.Tn[10].n51 VGND 0.46113f
C9388 XThC.Tn[10].n52 VGND 0.03515f
C9389 XThC.Tn[10].t4 VGND 0.01446f
C9390 XThC.Tn[10].t3 VGND 0.01446f
C9391 XThC.Tn[10].n53 VGND 0.03125f
C9392 XThC.Tn[10].t6 VGND 0.01446f
C9393 XThC.Tn[10].t0 VGND 0.01446f
C9394 XThC.Tn[10].n54 VGND 0.04756f
C9395 XThC.Tn[10].n55 VGND 0.13215f
C9396 XThC.Tn[10].n56 VGND 0.02078f
C9397 XThC.Tn[10].t11 VGND 0.01446f
C9398 XThC.Tn[10].t10 VGND 0.01446f
C9399 XThC.Tn[10].n57 VGND 0.04391f
C9400 XThC.Tn[10].t9 VGND 0.01446f
C9401 XThC.Tn[10].t8 VGND 0.01446f
C9402 XThC.Tn[10].n58 VGND 0.03215f
C9403 XThC.Tn[10].n59 VGND 0.14309f
C9404 Iout.n0 VGND 0.22972f
C9405 Iout.n1 VGND 1.20114f
C9406 Iout.n2 VGND 0.22972f
C9407 Iout.n3 VGND 0.22972f
C9408 Iout.t119 VGND 0.02212f
C9409 Iout.n4 VGND 0.04919f
C9410 Iout.n5 VGND 0.19431f
C9411 Iout.n6 VGND 0.22972f
C9412 Iout.n7 VGND 1.20114f
C9413 Iout.n8 VGND 0.22972f
C9414 Iout.t238 VGND 0.02212f
C9415 Iout.n9 VGND 0.04919f
C9416 Iout.n10 VGND 0.19431f
C9417 Iout.n11 VGND 0.22972f
C9418 Iout.n12 VGND 1.20114f
C9419 Iout.n13 VGND 0.22972f
C9420 Iout.t183 VGND 0.02212f
C9421 Iout.n14 VGND 0.04919f
C9422 Iout.n15 VGND 0.19431f
C9423 Iout.n16 VGND 0.22972f
C9424 Iout.n17 VGND 1.20114f
C9425 Iout.n18 VGND 0.22972f
C9426 Iout.t16 VGND 0.02212f
C9427 Iout.n19 VGND 0.04919f
C9428 Iout.n20 VGND 0.19431f
C9429 Iout.n21 VGND 0.47625f
C9430 Iout.t139 VGND 0.02212f
C9431 Iout.n22 VGND 0.04919f
C9432 Iout.n23 VGND 0.28657f
C9433 Iout.n24 VGND 0.22972f
C9434 Iout.n25 VGND 0.22972f
C9435 Iout.n26 VGND 0.22972f
C9436 Iout.n27 VGND 0.22972f
C9437 Iout.n28 VGND 0.22972f
C9438 Iout.n29 VGND 0.22972f
C9439 Iout.n30 VGND 0.22972f
C9440 Iout.n31 VGND 0.22972f
C9441 Iout.n32 VGND 0.22972f
C9442 Iout.n33 VGND 0.22972f
C9443 Iout.n34 VGND 0.22972f
C9444 Iout.n35 VGND 0.22972f
C9445 Iout.n36 VGND 0.22972f
C9446 Iout.n37 VGND 0.22972f
C9447 Iout.t30 VGND 0.02212f
C9448 Iout.n38 VGND 0.04919f
C9449 Iout.n39 VGND 0.02502f
C9450 Iout.n40 VGND 0.22972f
C9451 Iout.n41 VGND 0.04584f
C9452 Iout.t71 VGND 0.02212f
C9453 Iout.n42 VGND 0.04919f
C9454 Iout.n43 VGND 0.02502f
C9455 Iout.t109 VGND 0.02212f
C9456 Iout.n44 VGND 0.04919f
C9457 Iout.n45 VGND 0.02502f
C9458 Iout.n46 VGND 0.22972f
C9459 Iout.t92 VGND 0.02212f
C9460 Iout.n47 VGND 0.04919f
C9461 Iout.n48 VGND 0.02502f
C9462 Iout.n49 VGND 0.22972f
C9463 Iout.t186 VGND 0.02212f
C9464 Iout.n50 VGND 0.04919f
C9465 Iout.n51 VGND 0.02502f
C9466 Iout.n52 VGND 0.22972f
C9467 Iout.t187 VGND 0.02212f
C9468 Iout.n53 VGND 0.04919f
C9469 Iout.n54 VGND 0.02502f
C9470 Iout.n55 VGND 0.22972f
C9471 Iout.t229 VGND 0.02212f
C9472 Iout.n56 VGND 0.04919f
C9473 Iout.n57 VGND 0.02502f
C9474 Iout.n58 VGND 0.22972f
C9475 Iout.t27 VGND 0.02212f
C9476 Iout.n59 VGND 0.04919f
C9477 Iout.n60 VGND 0.02502f
C9478 Iout.n61 VGND 0.22972f
C9479 Iout.t211 VGND 0.02212f
C9480 Iout.n62 VGND 0.04919f
C9481 Iout.n63 VGND 0.02502f
C9482 Iout.n64 VGND 0.22972f
C9483 Iout.t60 VGND 0.02212f
C9484 Iout.n65 VGND 0.04919f
C9485 Iout.n66 VGND 0.02502f
C9486 Iout.n67 VGND 0.22972f
C9487 Iout.t43 VGND 0.02212f
C9488 Iout.n68 VGND 0.04919f
C9489 Iout.n69 VGND 0.02502f
C9490 Iout.n70 VGND 0.22972f
C9491 Iout.t111 VGND 0.02212f
C9492 Iout.n71 VGND 0.04919f
C9493 Iout.n72 VGND 0.02502f
C9494 Iout.n73 VGND 0.22972f
C9495 Iout.t76 VGND 0.02212f
C9496 Iout.n74 VGND 0.04919f
C9497 Iout.n75 VGND 0.02502f
C9498 Iout.n76 VGND 0.22972f
C9499 Iout.t190 VGND 0.02212f
C9500 Iout.n77 VGND 0.04919f
C9501 Iout.n78 VGND 0.02502f
C9502 Iout.n79 VGND 0.22972f
C9503 Iout.n80 VGND 0.22972f
C9504 Iout.t131 VGND 0.02212f
C9505 Iout.n81 VGND 0.04919f
C9506 Iout.n82 VGND 0.02502f
C9507 Iout.n83 VGND 0.22972f
C9508 Iout.n84 VGND 0.04584f
C9509 Iout.t177 VGND 0.02212f
C9510 Iout.n85 VGND 0.04919f
C9511 Iout.n86 VGND 0.02502f
C9512 Iout.t21 VGND 0.02212f
C9513 Iout.n87 VGND 0.04919f
C9514 Iout.n88 VGND 0.02502f
C9515 Iout.n89 VGND 0.22972f
C9516 Iout.t95 VGND 0.02212f
C9517 Iout.n90 VGND 0.04919f
C9518 Iout.n91 VGND 0.02502f
C9519 Iout.n92 VGND 0.22972f
C9520 Iout.t29 VGND 0.02212f
C9521 Iout.n93 VGND 0.04919f
C9522 Iout.n94 VGND 0.02502f
C9523 Iout.n95 VGND 0.22972f
C9524 Iout.t94 VGND 0.02212f
C9525 Iout.n96 VGND 0.04919f
C9526 Iout.n97 VGND 0.02502f
C9527 Iout.n98 VGND 0.22972f
C9528 Iout.t55 VGND 0.02212f
C9529 Iout.n99 VGND 0.04919f
C9530 Iout.n100 VGND 0.02502f
C9531 Iout.n101 VGND 0.22972f
C9532 Iout.t33 VGND 0.02212f
C9533 Iout.n102 VGND 0.04919f
C9534 Iout.n103 VGND 0.02502f
C9535 Iout.n104 VGND 0.22972f
C9536 Iout.t157 VGND 0.02212f
C9537 Iout.n105 VGND 0.04919f
C9538 Iout.n106 VGND 0.02502f
C9539 Iout.n107 VGND 0.22972f
C9540 Iout.t145 VGND 0.02212f
C9541 Iout.n108 VGND 0.04919f
C9542 Iout.n109 VGND 0.02502f
C9543 Iout.n110 VGND 0.22972f
C9544 Iout.t155 VGND 0.02212f
C9545 Iout.n111 VGND 0.04919f
C9546 Iout.n112 VGND 0.02502f
C9547 Iout.n113 VGND 0.22972f
C9548 Iout.t168 VGND 0.02212f
C9549 Iout.n114 VGND 0.04919f
C9550 Iout.n115 VGND 0.02502f
C9551 Iout.n116 VGND 0.22972f
C9552 Iout.t152 VGND 0.02212f
C9553 Iout.n117 VGND 0.04919f
C9554 Iout.n118 VGND 0.02502f
C9555 Iout.n119 VGND 0.22972f
C9556 Iout.t189 VGND 0.02212f
C9557 Iout.n120 VGND 0.04919f
C9558 Iout.n121 VGND 0.02502f
C9559 Iout.n122 VGND 0.04584f
C9560 Iout.t161 VGND 0.02212f
C9561 Iout.n123 VGND 0.04919f
C9562 Iout.n124 VGND 0.02502f
C9563 Iout.n125 VGND 0.22972f
C9564 Iout.n126 VGND 0.22972f
C9565 Iout.t173 VGND 0.02212f
C9566 Iout.n127 VGND 0.04919f
C9567 Iout.n128 VGND 0.02502f
C9568 Iout.n129 VGND 0.04584f
C9569 Iout.t236 VGND 0.02212f
C9570 Iout.n130 VGND 0.04919f
C9571 Iout.n131 VGND 0.02502f
C9572 Iout.n132 VGND 0.22972f
C9573 Iout.t218 VGND 0.02212f
C9574 Iout.n133 VGND 0.04919f
C9575 Iout.n134 VGND 0.02502f
C9576 Iout.n135 VGND 0.04584f
C9577 Iout.t220 VGND 0.02212f
C9578 Iout.n136 VGND 0.04919f
C9579 Iout.n137 VGND 0.02502f
C9580 Iout.n138 VGND 0.22972f
C9581 Iout.n139 VGND 0.22972f
C9582 Iout.t80 VGND 0.02212f
C9583 Iout.n140 VGND 0.04919f
C9584 Iout.n141 VGND 0.02502f
C9585 Iout.n142 VGND 0.04584f
C9586 Iout.t14 VGND 0.02212f
C9587 Iout.n143 VGND 0.04919f
C9588 Iout.n144 VGND 0.02502f
C9589 Iout.n145 VGND 0.13561f
C9590 Iout.t170 VGND 0.02212f
C9591 Iout.n146 VGND 0.04919f
C9592 Iout.n147 VGND 0.02502f
C9593 Iout.n148 VGND 0.04584f
C9594 Iout.t17 VGND 0.02212f
C9595 Iout.n149 VGND 0.04919f
C9596 Iout.n150 VGND 0.02502f
C9597 Iout.n151 VGND 0.22972f
C9598 Iout.n152 VGND 0.13561f
C9599 Iout.n153 VGND 0.22972f
C9600 Iout.n154 VGND 0.22972f
C9601 Iout.n155 VGND 0.22972f
C9602 Iout.t205 VGND 0.02212f
C9603 Iout.n156 VGND 0.04919f
C9604 Iout.n157 VGND 0.02502f
C9605 Iout.n158 VGND 0.22972f
C9606 Iout.n159 VGND 0.22972f
C9607 Iout.n160 VGND 0.22972f
C9608 Iout.n161 VGND 0.22972f
C9609 Iout.n162 VGND 0.22972f
C9610 Iout.n163 VGND 0.22972f
C9611 Iout.n164 VGND 0.22972f
C9612 Iout.n165 VGND 0.22972f
C9613 Iout.n166 VGND 0.22972f
C9614 Iout.n167 VGND 0.22972f
C9615 Iout.t166 VGND 0.02212f
C9616 Iout.n168 VGND 0.04919f
C9617 Iout.n169 VGND 0.02502f
C9618 Iout.n170 VGND 0.22972f
C9619 Iout.n171 VGND 0.04584f
C9620 Iout.t53 VGND 0.02212f
C9621 Iout.n172 VGND 0.04919f
C9622 Iout.n173 VGND 0.02502f
C9623 Iout.t85 VGND 0.02212f
C9624 Iout.n174 VGND 0.04919f
C9625 Iout.n175 VGND 0.02502f
C9626 Iout.n176 VGND 0.22972f
C9627 Iout.t10 VGND 0.02212f
C9628 Iout.n177 VGND 0.04919f
C9629 Iout.n178 VGND 0.02502f
C9630 Iout.n179 VGND 0.22972f
C9631 Iout.t52 VGND 0.02212f
C9632 Iout.n180 VGND 0.04919f
C9633 Iout.n181 VGND 0.02502f
C9634 Iout.n182 VGND 0.22972f
C9635 Iout.t5 VGND 0.02212f
C9636 Iout.n183 VGND 0.04919f
C9637 Iout.n184 VGND 0.02502f
C9638 Iout.n185 VGND 0.22972f
C9639 Iout.t91 VGND 0.02212f
C9640 Iout.n186 VGND 0.04919f
C9641 Iout.n187 VGND 0.02502f
C9642 Iout.n188 VGND 0.22972f
C9643 Iout.t120 VGND 0.02212f
C9644 Iout.n189 VGND 0.04919f
C9645 Iout.n190 VGND 0.02502f
C9646 Iout.n191 VGND 0.13561f
C9647 Iout.t75 VGND 0.02212f
C9648 Iout.n192 VGND 0.04919f
C9649 Iout.n193 VGND 0.02502f
C9650 Iout.n194 VGND 0.04584f
C9651 Iout.t194 VGND 0.02212f
C9652 Iout.n195 VGND 0.04919f
C9653 Iout.n196 VGND 0.02502f
C9654 Iout.n197 VGND 0.13561f
C9655 Iout.n198 VGND 0.04584f
C9656 Iout.t118 VGND 0.02212f
C9657 Iout.n199 VGND 0.04919f
C9658 Iout.n200 VGND 0.02502f
C9659 Iout.n201 VGND 0.04584f
C9660 Iout.t87 VGND 0.02212f
C9661 Iout.n202 VGND 0.04919f
C9662 Iout.n203 VGND 0.02502f
C9663 Iout.n204 VGND 0.13561f
C9664 Iout.n205 VGND 0.04584f
C9665 Iout.t144 VGND 0.02212f
C9666 Iout.n206 VGND 0.04919f
C9667 Iout.n207 VGND 0.02502f
C9668 Iout.n208 VGND 0.13561f
C9669 Iout.n209 VGND 0.04584f
C9670 Iout.t141 VGND 0.02212f
C9671 Iout.n210 VGND 0.04919f
C9672 Iout.n211 VGND 0.02502f
C9673 Iout.n212 VGND 0.13561f
C9674 Iout.n213 VGND 0.04584f
C9675 Iout.t26 VGND 0.02212f
C9676 Iout.n214 VGND 0.04919f
C9677 Iout.n215 VGND 0.02502f
C9678 Iout.n216 VGND 0.13561f
C9679 Iout.n217 VGND 0.04584f
C9680 Iout.t156 VGND 0.02212f
C9681 Iout.n218 VGND 0.04919f
C9682 Iout.n219 VGND 0.02502f
C9683 Iout.n220 VGND 0.13561f
C9684 Iout.n221 VGND 0.04584f
C9685 Iout.t67 VGND 0.02212f
C9686 Iout.n222 VGND 0.04919f
C9687 Iout.n223 VGND 0.02502f
C9688 Iout.n224 VGND 0.13561f
C9689 Iout.n225 VGND 0.04584f
C9690 Iout.t180 VGND 0.02212f
C9691 Iout.n226 VGND 0.04919f
C9692 Iout.n227 VGND 0.02502f
C9693 Iout.n228 VGND 0.04584f
C9694 Iout.n229 VGND 0.13561f
C9695 Iout.n230 VGND 0.22972f
C9696 Iout.n231 VGND 0.04584f
C9697 Iout.t132 VGND 0.02212f
C9698 Iout.n232 VGND 0.04919f
C9699 Iout.n233 VGND 0.02502f
C9700 Iout.n234 VGND 0.04584f
C9701 Iout.t212 VGND 0.02212f
C9702 Iout.n235 VGND 0.04919f
C9703 Iout.n236 VGND 0.02502f
C9704 Iout.n237 VGND 0.04584f
C9705 Iout.t7 VGND 0.02212f
C9706 Iout.n238 VGND 0.04919f
C9707 Iout.n239 VGND 0.02502f
C9708 Iout.n240 VGND 0.04584f
C9709 Iout.t46 VGND 0.02212f
C9710 Iout.n241 VGND 0.04919f
C9711 Iout.n242 VGND 0.02502f
C9712 Iout.n243 VGND 0.04584f
C9713 Iout.t44 VGND 0.02212f
C9714 Iout.n244 VGND 0.04919f
C9715 Iout.n245 VGND 0.02502f
C9716 Iout.n246 VGND 0.04584f
C9717 Iout.t241 VGND 0.02212f
C9718 Iout.n247 VGND 0.04919f
C9719 Iout.n248 VGND 0.02502f
C9720 Iout.n249 VGND 0.04584f
C9721 Iout.t22 VGND 0.02212f
C9722 Iout.n250 VGND 0.04919f
C9723 Iout.n251 VGND 0.02502f
C9724 Iout.t114 VGND 0.02212f
C9725 Iout.n252 VGND 0.04919f
C9726 Iout.n253 VGND 0.02502f
C9727 Iout.n254 VGND 0.04584f
C9728 Iout.t250 VGND 0.02212f
C9729 Iout.n255 VGND 0.04919f
C9730 Iout.n256 VGND 0.02502f
C9731 Iout.n257 VGND 0.04584f
C9732 Iout.n258 VGND 0.22972f
C9733 Iout.t223 VGND 0.02212f
C9734 Iout.n259 VGND 0.04919f
C9735 Iout.n260 VGND 0.02502f
C9736 Iout.n261 VGND 0.04584f
C9737 Iout.n262 VGND 0.22972f
C9738 Iout.n263 VGND 0.22972f
C9739 Iout.n264 VGND 0.04584f
C9740 Iout.t188 VGND 0.02212f
C9741 Iout.n265 VGND 0.04919f
C9742 Iout.n266 VGND 0.02502f
C9743 Iout.n267 VGND 0.04584f
C9744 Iout.n268 VGND 0.22972f
C9745 Iout.n269 VGND 0.22972f
C9746 Iout.n270 VGND 0.04584f
C9747 Iout.t225 VGND 0.02212f
C9748 Iout.n271 VGND 0.04919f
C9749 Iout.n272 VGND 0.02502f
C9750 Iout.n273 VGND 0.04584f
C9751 Iout.n274 VGND 0.22972f
C9752 Iout.n275 VGND 0.22972f
C9753 Iout.n276 VGND 0.04584f
C9754 Iout.t174 VGND 0.02212f
C9755 Iout.n277 VGND 0.04919f
C9756 Iout.n278 VGND 0.02502f
C9757 Iout.n279 VGND 0.04584f
C9758 Iout.n280 VGND 0.22972f
C9759 Iout.n281 VGND 0.22972f
C9760 Iout.n282 VGND 0.04584f
C9761 Iout.t127 VGND 0.02212f
C9762 Iout.n283 VGND 0.04919f
C9763 Iout.n284 VGND 0.02502f
C9764 Iout.n285 VGND 0.04584f
C9765 Iout.n286 VGND 0.22972f
C9766 Iout.n287 VGND 0.22972f
C9767 Iout.n288 VGND 0.04584f
C9768 Iout.t116 VGND 0.02212f
C9769 Iout.n289 VGND 0.04919f
C9770 Iout.n290 VGND 0.02502f
C9771 Iout.n291 VGND 0.04584f
C9772 Iout.n292 VGND 0.22972f
C9773 Iout.n293 VGND 0.22972f
C9774 Iout.n294 VGND 0.04584f
C9775 Iout.t252 VGND 0.02212f
C9776 Iout.n295 VGND 0.04919f
C9777 Iout.n296 VGND 0.02502f
C9778 Iout.n297 VGND 0.04584f
C9779 Iout.n298 VGND 0.22972f
C9780 Iout.n299 VGND 0.22972f
C9781 Iout.n300 VGND 0.04584f
C9782 Iout.t4 VGND 0.02212f
C9783 Iout.n301 VGND 0.04919f
C9784 Iout.n302 VGND 0.02502f
C9785 Iout.n303 VGND 0.04584f
C9786 Iout.n304 VGND 0.22972f
C9787 Iout.t216 VGND 0.02212f
C9788 Iout.n305 VGND 0.04919f
C9789 Iout.n306 VGND 0.02502f
C9790 Iout.n307 VGND 0.04584f
C9791 Iout.t193 VGND 0.02212f
C9792 Iout.n308 VGND 0.04919f
C9793 Iout.n309 VGND 0.02502f
C9794 Iout.n310 VGND 0.04584f
C9795 Iout.t25 VGND 0.02212f
C9796 Iout.n311 VGND 0.04919f
C9797 Iout.n312 VGND 0.02502f
C9798 Iout.n313 VGND 0.04584f
C9799 Iout.t154 VGND 0.02212f
C9800 Iout.n314 VGND 0.04919f
C9801 Iout.n315 VGND 0.02502f
C9802 Iout.n316 VGND 0.04584f
C9803 Iout.t143 VGND 0.02212f
C9804 Iout.n317 VGND 0.04919f
C9805 Iout.n318 VGND 0.02502f
C9806 Iout.n319 VGND 0.04584f
C9807 Iout.t113 VGND 0.02212f
C9808 Iout.n320 VGND 0.04919f
C9809 Iout.n321 VGND 0.02502f
C9810 Iout.n322 VGND 0.04584f
C9811 Iout.t213 VGND 0.02212f
C9812 Iout.n323 VGND 0.04919f
C9813 Iout.n324 VGND 0.02502f
C9814 Iout.n325 VGND 0.04584f
C9815 Iout.t230 VGND 0.02212f
C9816 Iout.n326 VGND 0.04919f
C9817 Iout.n327 VGND 0.02502f
C9818 Iout.n328 VGND 0.04584f
C9819 Iout.t47 VGND 0.02212f
C9820 Iout.n329 VGND 0.04919f
C9821 Iout.n330 VGND 0.02502f
C9822 Iout.n331 VGND 0.04584f
C9823 Iout.n332 VGND 0.22972f
C9824 Iout.t136 VGND 0.02212f
C9825 Iout.n333 VGND 0.04919f
C9826 Iout.n334 VGND 0.02502f
C9827 Iout.n335 VGND 0.04584f
C9828 Iout.t215 VGND 0.02212f
C9829 Iout.n336 VGND 0.04919f
C9830 Iout.n337 VGND 0.02502f
C9831 Iout.n338 VGND 0.04584f
C9832 Iout.t151 VGND 0.02212f
C9833 Iout.n339 VGND 0.04919f
C9834 Iout.n340 VGND 0.02502f
C9835 Iout.n341 VGND 0.04584f
C9836 Iout.t184 VGND 0.02212f
C9837 Iout.n342 VGND 0.04919f
C9838 Iout.n343 VGND 0.02502f
C9839 Iout.n344 VGND 0.04584f
C9840 Iout.t214 VGND 0.02212f
C9841 Iout.n345 VGND 0.04919f
C9842 Iout.n346 VGND 0.02502f
C9843 Iout.n347 VGND 0.04584f
C9844 Iout.t233 VGND 0.02212f
C9845 Iout.n348 VGND 0.04919f
C9846 Iout.n349 VGND 0.02502f
C9847 Iout.n350 VGND 0.04584f
C9848 Iout.t90 VGND 0.02212f
C9849 Iout.n351 VGND 0.04919f
C9850 Iout.n352 VGND 0.02502f
C9851 Iout.n353 VGND 0.04584f
C9852 Iout.t66 VGND 0.02212f
C9853 Iout.n354 VGND 0.04919f
C9854 Iout.n355 VGND 0.02502f
C9855 Iout.n356 VGND 0.04584f
C9856 Iout.t251 VGND 0.02212f
C9857 Iout.n357 VGND 0.04919f
C9858 Iout.n358 VGND 0.02502f
C9859 Iout.n359 VGND 0.04584f
C9860 Iout.t82 VGND 0.02212f
C9861 Iout.n360 VGND 0.04919f
C9862 Iout.n361 VGND 0.02502f
C9863 Iout.n362 VGND 0.04584f
C9864 Iout.t248 VGND 0.02212f
C9865 Iout.n363 VGND 0.04919f
C9866 Iout.n364 VGND 0.02502f
C9867 Iout.n365 VGND 0.04584f
C9868 Iout.t70 VGND 0.02212f
C9869 Iout.n366 VGND 0.04919f
C9870 Iout.n367 VGND 0.02502f
C9871 Iout.n368 VGND 0.04584f
C9872 Iout.n369 VGND 0.22972f
C9873 Iout.t62 VGND 0.02212f
C9874 Iout.n370 VGND 0.04919f
C9875 Iout.n371 VGND 0.02502f
C9876 Iout.n372 VGND 0.04584f
C9877 Iout.n373 VGND 0.22972f
C9878 Iout.n374 VGND 0.22972f
C9879 Iout.n375 VGND 0.04584f
C9880 Iout.t72 VGND 0.02212f
C9881 Iout.n376 VGND 0.04919f
C9882 Iout.n377 VGND 0.02502f
C9883 Iout.t54 VGND 0.02212f
C9884 Iout.n378 VGND 0.04919f
C9885 Iout.n379 VGND 0.02502f
C9886 Iout.n380 VGND 0.04584f
C9887 Iout.n381 VGND 0.22972f
C9888 Iout.n382 VGND 0.22972f
C9889 Iout.n383 VGND 0.04584f
C9890 Iout.t175 VGND 0.02212f
C9891 Iout.n384 VGND 0.04919f
C9892 Iout.n385 VGND 0.02502f
C9893 Iout.t61 VGND 0.02212f
C9894 Iout.n386 VGND 0.04919f
C9895 Iout.n387 VGND 0.02502f
C9896 Iout.n388 VGND 0.04584f
C9897 Iout.n389 VGND 0.22972f
C9898 Iout.n390 VGND 0.22972f
C9899 Iout.n391 VGND 0.04584f
C9900 Iout.t237 VGND 0.02212f
C9901 Iout.n392 VGND 0.04919f
C9902 Iout.n393 VGND 0.02502f
C9903 Iout.t195 VGND 0.02212f
C9904 Iout.n394 VGND 0.04919f
C9905 Iout.n395 VGND 0.02502f
C9906 Iout.n396 VGND 0.04584f
C9907 Iout.n397 VGND 0.22972f
C9908 Iout.n398 VGND 0.22972f
C9909 Iout.n399 VGND 0.04584f
C9910 Iout.t181 VGND 0.02212f
C9911 Iout.n400 VGND 0.04919f
C9912 Iout.n401 VGND 0.02502f
C9913 Iout.t23 VGND 0.02212f
C9914 Iout.n402 VGND 0.04919f
C9915 Iout.n403 VGND 0.02502f
C9916 Iout.n404 VGND 0.04584f
C9917 Iout.n405 VGND 0.22972f
C9918 Iout.n406 VGND 0.22972f
C9919 Iout.n407 VGND 0.04584f
C9920 Iout.t11 VGND 0.02212f
C9921 Iout.n408 VGND 0.04919f
C9922 Iout.n409 VGND 0.02502f
C9923 Iout.t40 VGND 0.02212f
C9924 Iout.n410 VGND 0.04919f
C9925 Iout.n411 VGND 0.02502f
C9926 Iout.n412 VGND 0.04584f
C9927 Iout.n413 VGND 0.22972f
C9928 Iout.n414 VGND 0.22972f
C9929 Iout.n415 VGND 0.04584f
C9930 Iout.t142 VGND 0.02212f
C9931 Iout.n416 VGND 0.04919f
C9932 Iout.n417 VGND 0.02502f
C9933 Iout.t162 VGND 0.02212f
C9934 Iout.n418 VGND 0.04919f
C9935 Iout.n419 VGND 0.02502f
C9936 Iout.n420 VGND 0.04584f
C9937 Iout.n421 VGND 0.22972f
C9938 Iout.n422 VGND 0.22972f
C9939 Iout.n423 VGND 0.04584f
C9940 Iout.t88 VGND 0.02212f
C9941 Iout.n424 VGND 0.04919f
C9942 Iout.n425 VGND 0.02502f
C9943 Iout.t210 VGND 0.02212f
C9944 Iout.n426 VGND 0.04919f
C9945 Iout.n427 VGND 0.02502f
C9946 Iout.n428 VGND 0.04584f
C9947 Iout.n429 VGND 0.22972f
C9948 Iout.n430 VGND 0.22972f
C9949 Iout.n431 VGND 0.04584f
C9950 Iout.t58 VGND 0.02212f
C9951 Iout.n432 VGND 0.04919f
C9952 Iout.n433 VGND 0.02502f
C9953 Iout.t18 VGND 0.02212f
C9954 Iout.n434 VGND 0.04919f
C9955 Iout.n435 VGND 0.02502f
C9956 Iout.n436 VGND 0.22972f
C9957 Iout.n437 VGND 0.04584f
C9958 Iout.t172 VGND 0.02212f
C9959 Iout.n438 VGND 0.04919f
C9960 Iout.n439 VGND 0.02502f
C9961 Iout.n440 VGND 0.04584f
C9962 Iout.t68 VGND 0.02212f
C9963 Iout.n441 VGND 0.04919f
C9964 Iout.n442 VGND 0.02502f
C9965 Iout.n443 VGND 0.04584f
C9966 Iout.n444 VGND 0.22972f
C9967 Iout.n445 VGND 0.22972f
C9968 Iout.n446 VGND 0.04584f
C9969 Iout.t176 VGND 0.02212f
C9970 Iout.n447 VGND 0.04919f
C9971 Iout.n448 VGND 0.02502f
C9972 Iout.t129 VGND 0.02212f
C9973 Iout.n449 VGND 0.04919f
C9974 Iout.n450 VGND 0.02502f
C9975 Iout.n451 VGND 0.04584f
C9976 Iout.t243 VGND 0.02212f
C9977 Iout.n452 VGND 0.04919f
C9978 Iout.n453 VGND 0.02502f
C9979 Iout.n454 VGND 0.04584f
C9980 Iout.n455 VGND 0.22972f
C9981 Iout.n456 VGND 0.22972f
C9982 Iout.n457 VGND 0.04584f
C9983 Iout.t146 VGND 0.02212f
C9984 Iout.n458 VGND 0.04919f
C9985 Iout.n459 VGND 0.02502f
C9986 Iout.t56 VGND 0.02212f
C9987 Iout.n460 VGND 0.04919f
C9988 Iout.n461 VGND 0.02502f
C9989 Iout.n462 VGND 0.04584f
C9990 Iout.t79 VGND 0.02212f
C9991 Iout.n463 VGND 0.04919f
C9992 Iout.n464 VGND 0.02502f
C9993 Iout.n465 VGND 0.04584f
C9994 Iout.n466 VGND 0.22972f
C9995 Iout.n467 VGND 0.22972f
C9996 Iout.n468 VGND 0.04584f
C9997 Iout.t150 VGND 0.02212f
C9998 Iout.n469 VGND 0.04919f
C9999 Iout.n470 VGND 0.02502f
C10000 Iout.n471 VGND 0.04584f
C10001 Iout.t106 VGND 0.02212f
C10002 Iout.n472 VGND 0.04919f
C10003 Iout.n473 VGND 0.02502f
C10004 Iout.n474 VGND 0.04584f
C10005 Iout.n475 VGND 0.22972f
C10006 Iout.n476 VGND 0.22972f
C10007 Iout.n477 VGND 0.04584f
C10008 Iout.t117 VGND 0.02212f
C10009 Iout.n478 VGND 0.04919f
C10010 Iout.n479 VGND 0.02502f
C10011 Iout.t138 VGND 0.02212f
C10012 Iout.n480 VGND 0.04919f
C10013 Iout.n481 VGND 0.02502f
C10014 Iout.n482 VGND 0.04584f
C10015 Iout.t153 VGND 0.02212f
C10016 Iout.n483 VGND 0.04919f
C10017 Iout.n484 VGND 0.02502f
C10018 Iout.n485 VGND 0.04584f
C10019 Iout.n486 VGND 0.22972f
C10020 Iout.n487 VGND 0.22972f
C10021 Iout.n488 VGND 0.04584f
C10022 Iout.t36 VGND 0.02212f
C10023 Iout.n489 VGND 0.04919f
C10024 Iout.n490 VGND 0.02502f
C10025 Iout.t160 VGND 0.02212f
C10026 Iout.n491 VGND 0.04919f
C10027 Iout.n492 VGND 0.02502f
C10028 Iout.n493 VGND 0.04584f
C10029 Iout.t51 VGND 0.02212f
C10030 Iout.n494 VGND 0.04919f
C10031 Iout.n495 VGND 0.02502f
C10032 Iout.n496 VGND 0.04584f
C10033 Iout.n497 VGND 0.22972f
C10034 Iout.n498 VGND 0.13561f
C10035 Iout.n499 VGND 0.04584f
C10036 Iout.t219 VGND 0.02212f
C10037 Iout.n500 VGND 0.04919f
C10038 Iout.n501 VGND 0.02502f
C10039 Iout.n502 VGND 0.13561f
C10040 Iout.n503 VGND 0.04584f
C10041 Iout.t246 VGND 0.02212f
C10042 Iout.n504 VGND 0.04919f
C10043 Iout.n505 VGND 0.02502f
C10044 Iout.n506 VGND 0.04584f
C10045 Iout.t207 VGND 0.02212f
C10046 Iout.n507 VGND 0.04919f
C10047 Iout.n508 VGND 0.02502f
C10048 Iout.t185 VGND 0.02212f
C10049 Iout.n509 VGND 0.04919f
C10050 Iout.n510 VGND 0.02502f
C10051 Iout.n511 VGND 0.13561f
C10052 Iout.n512 VGND 0.04584f
C10053 Iout.t41 VGND 0.02212f
C10054 Iout.n513 VGND 0.04919f
C10055 Iout.n514 VGND 0.02502f
C10056 Iout.n515 VGND 0.04584f
C10057 Iout.n516 VGND 0.13561f
C10058 Iout.n517 VGND 0.22972f
C10059 Iout.n518 VGND 0.04584f
C10060 Iout.t24 VGND 0.02212f
C10061 Iout.n519 VGND 0.04919f
C10062 Iout.n520 VGND 0.02502f
C10063 Iout.n521 VGND 0.04584f
C10064 Iout.n522 VGND 0.22972f
C10065 Iout.n523 VGND 0.22972f
C10066 Iout.n524 VGND 0.04584f
C10067 Iout.t96 VGND 0.02212f
C10068 Iout.n525 VGND 0.04919f
C10069 Iout.n526 VGND 0.02502f
C10070 Iout.n527 VGND 0.04584f
C10071 Iout.n528 VGND 0.22972f
C10072 Iout.n529 VGND 0.22972f
C10073 Iout.n530 VGND 0.04584f
C10074 Iout.t171 VGND 0.02212f
C10075 Iout.n531 VGND 0.04919f
C10076 Iout.n532 VGND 0.02502f
C10077 Iout.n533 VGND 0.04584f
C10078 Iout.t217 VGND 0.02212f
C10079 Iout.n534 VGND 0.04919f
C10080 Iout.n535 VGND 0.02502f
C10081 Iout.t69 VGND 0.02212f
C10082 Iout.n536 VGND 0.04919f
C10083 Iout.n537 VGND 0.02502f
C10084 Iout.n538 VGND 0.04584f
C10085 Iout.n539 VGND 0.22972f
C10086 Iout.n540 VGND 0.22972f
C10087 Iout.n541 VGND 0.04584f
C10088 Iout.t226 VGND 0.02212f
C10089 Iout.n542 VGND 0.04919f
C10090 Iout.n543 VGND 0.02502f
C10091 Iout.n544 VGND 0.04584f
C10092 Iout.n545 VGND 0.22972f
C10093 Iout.n546 VGND 0.22972f
C10094 Iout.n547 VGND 0.04584f
C10095 Iout.t135 VGND 0.02212f
C10096 Iout.n548 VGND 0.04919f
C10097 Iout.n549 VGND 0.02502f
C10098 Iout.n550 VGND 0.04584f
C10099 Iout.n551 VGND 0.22972f
C10100 Iout.n552 VGND 0.22972f
C10101 Iout.n553 VGND 0.04584f
C10102 Iout.t49 VGND 0.02212f
C10103 Iout.n554 VGND 0.04919f
C10104 Iout.n555 VGND 0.02502f
C10105 Iout.n556 VGND 0.04584f
C10106 Iout.t209 VGND 0.02212f
C10107 Iout.n557 VGND 0.04919f
C10108 Iout.n558 VGND 0.02502f
C10109 Iout.t108 VGND 0.02212f
C10110 Iout.n559 VGND 0.04919f
C10111 Iout.n560 VGND 0.02502f
C10112 Iout.n561 VGND 0.04584f
C10113 Iout.n562 VGND 0.22972f
C10114 Iout.t48 VGND 0.02212f
C10115 Iout.n563 VGND 0.04919f
C10116 Iout.n564 VGND 0.02502f
C10117 Iout.n565 VGND 0.04584f
C10118 Iout.n566 VGND 0.22972f
C10119 Iout.n567 VGND 0.22972f
C10120 Iout.n568 VGND 0.04584f
C10121 Iout.t255 VGND 0.02212f
C10122 Iout.n569 VGND 0.04919f
C10123 Iout.n570 VGND 0.02502f
C10124 Iout.n571 VGND 0.04584f
C10125 Iout.n572 VGND 0.22972f
C10126 Iout.t15 VGND 0.02212f
C10127 Iout.n573 VGND 0.04919f
C10128 Iout.n574 VGND 0.02502f
C10129 Iout.n575 VGND 0.04584f
C10130 Iout.t197 VGND 0.02212f
C10131 Iout.n576 VGND 0.04919f
C10132 Iout.n577 VGND 0.02502f
C10133 Iout.n578 VGND 0.04584f
C10134 Iout.n579 VGND 0.22972f
C10135 Iout.n580 VGND 0.22972f
C10136 Iout.n581 VGND 0.04584f
C10137 Iout.t224 VGND 0.02212f
C10138 Iout.n582 VGND 0.04919f
C10139 Iout.n583 VGND 0.02502f
C10140 Iout.n584 VGND 0.04584f
C10141 Iout.n585 VGND 0.22972f
C10142 Iout.n586 VGND 0.22972f
C10143 Iout.n587 VGND 0.04584f
C10144 Iout.t81 VGND 0.02212f
C10145 Iout.n588 VGND 0.04919f
C10146 Iout.n589 VGND 0.02502f
C10147 Iout.n590 VGND 0.04584f
C10148 Iout.n591 VGND 0.22972f
C10149 Iout.n592 VGND 0.22972f
C10150 Iout.n593 VGND 0.04584f
C10151 Iout.t164 VGND 0.02212f
C10152 Iout.n594 VGND 0.04919f
C10153 Iout.n595 VGND 0.02502f
C10154 Iout.n596 VGND 0.04584f
C10155 Iout.n597 VGND 0.22972f
C10156 Iout.n598 VGND 0.22972f
C10157 Iout.n599 VGND 0.04584f
C10158 Iout.t137 VGND 0.02212f
C10159 Iout.n600 VGND 0.04919f
C10160 Iout.n601 VGND 0.02502f
C10161 Iout.n602 VGND 0.04584f
C10162 Iout.n603 VGND 0.22972f
C10163 Iout.n604 VGND 0.22972f
C10164 Iout.n605 VGND 0.04584f
C10165 Iout.t86 VGND 0.02212f
C10166 Iout.n606 VGND 0.04919f
C10167 Iout.n607 VGND 0.02502f
C10168 Iout.n608 VGND 0.04584f
C10169 Iout.n609 VGND 0.22972f
C10170 Iout.n610 VGND 0.22972f
C10171 Iout.n611 VGND 0.04584f
C10172 Iout.t244 VGND 0.02212f
C10173 Iout.n612 VGND 0.04919f
C10174 Iout.n613 VGND 0.02502f
C10175 Iout.n614 VGND 0.04584f
C10176 Iout.n615 VGND 0.22972f
C10177 Iout.n616 VGND 0.22972f
C10178 Iout.n617 VGND 0.04584f
C10179 Iout.t98 VGND 0.02212f
C10180 Iout.n618 VGND 0.04919f
C10181 Iout.n619 VGND 0.02502f
C10182 Iout.n620 VGND 0.04584f
C10183 Iout.n621 VGND 0.22972f
C10184 Iout.n622 VGND 0.22972f
C10185 Iout.n623 VGND 0.04584f
C10186 Iout.t239 VGND 0.02212f
C10187 Iout.n624 VGND 0.04919f
C10188 Iout.n625 VGND 0.02502f
C10189 Iout.n626 VGND 0.04584f
C10190 Iout.n627 VGND 0.22972f
C10191 Iout.n628 VGND 0.22972f
C10192 Iout.n629 VGND 0.04584f
C10193 Iout.t6 VGND 0.02212f
C10194 Iout.n630 VGND 0.04919f
C10195 Iout.n631 VGND 0.02502f
C10196 Iout.n632 VGND 0.04584f
C10197 Iout.n633 VGND 0.22972f
C10198 Iout.n634 VGND 0.22972f
C10199 Iout.n635 VGND 0.04584f
C10200 Iout.t201 VGND 0.02212f
C10201 Iout.n636 VGND 0.04919f
C10202 Iout.n637 VGND 0.02502f
C10203 Iout.n638 VGND 0.04584f
C10204 Iout.n639 VGND 0.22972f
C10205 Iout.n640 VGND 0.22972f
C10206 Iout.n641 VGND 0.04584f
C10207 Iout.t73 VGND 0.02212f
C10208 Iout.n642 VGND 0.04919f
C10209 Iout.n643 VGND 0.02502f
C10210 Iout.n644 VGND 0.04584f
C10211 Iout.n645 VGND 0.22972f
C10212 Iout.n646 VGND 0.22972f
C10213 Iout.n647 VGND 0.04584f
C10214 Iout.t228 VGND 0.02212f
C10215 Iout.n648 VGND 0.04919f
C10216 Iout.n649 VGND 0.02502f
C10217 Iout.n650 VGND 0.04584f
C10218 Iout.n651 VGND 0.22972f
C10219 Iout.n652 VGND 0.22972f
C10220 Iout.n653 VGND 0.04584f
C10221 Iout.t134 VGND 0.02212f
C10222 Iout.n654 VGND 0.04919f
C10223 Iout.n655 VGND 0.02502f
C10224 Iout.n656 VGND 0.04584f
C10225 Iout.t8 VGND 0.02212f
C10226 Iout.n657 VGND 0.04919f
C10227 Iout.n658 VGND 0.02502f
C10228 Iout.n659 VGND 0.04584f
C10229 Iout.t206 VGND 0.02212f
C10230 Iout.n660 VGND 0.04919f
C10231 Iout.n661 VGND 0.02502f
C10232 Iout.n662 VGND 0.04584f
C10233 Iout.t126 VGND 0.02212f
C10234 Iout.n663 VGND 0.04919f
C10235 Iout.n664 VGND 0.02502f
C10236 Iout.n665 VGND 0.04584f
C10237 Iout.t84 VGND 0.02212f
C10238 Iout.n666 VGND 0.04919f
C10239 Iout.n667 VGND 0.02502f
C10240 Iout.n668 VGND 0.04584f
C10241 Iout.t37 VGND 0.02212f
C10242 Iout.n669 VGND 0.04919f
C10243 Iout.n670 VGND 0.02502f
C10244 Iout.n671 VGND 0.04584f
C10245 Iout.t112 VGND 0.02212f
C10246 Iout.n672 VGND 0.04919f
C10247 Iout.n673 VGND 0.02502f
C10248 Iout.n674 VGND 0.04584f
C10249 Iout.t247 VGND 0.02212f
C10250 Iout.n675 VGND 0.04919f
C10251 Iout.n676 VGND 0.02502f
C10252 Iout.n677 VGND 0.04584f
C10253 Iout.t240 VGND 0.02212f
C10254 Iout.n678 VGND 0.04919f
C10255 Iout.n679 VGND 0.02502f
C10256 Iout.n680 VGND 0.04584f
C10257 Iout.t140 VGND 0.02212f
C10258 Iout.n681 VGND 0.04919f
C10259 Iout.n682 VGND 0.02502f
C10260 Iout.n683 VGND 0.04584f
C10261 Iout.t182 VGND 0.02212f
C10262 Iout.n684 VGND 0.04919f
C10263 Iout.n685 VGND 0.02502f
C10264 Iout.n686 VGND 0.04584f
C10265 Iout.t59 VGND 0.02212f
C10266 Iout.n687 VGND 0.04919f
C10267 Iout.n688 VGND 0.02502f
C10268 Iout.n689 VGND 0.04584f
C10269 Iout.t19 VGND 0.02212f
C10270 Iout.n690 VGND 0.04919f
C10271 Iout.n691 VGND 0.02502f
C10272 Iout.t198 VGND 0.02212f
C10273 Iout.n692 VGND 0.04919f
C10274 Iout.n693 VGND 0.02502f
C10275 Iout.n694 VGND 0.04584f
C10276 Iout.t34 VGND 0.02212f
C10277 Iout.n695 VGND 0.04919f
C10278 Iout.n696 VGND 0.02502f
C10279 Iout.n697 VGND 0.04584f
C10280 Iout.n698 VGND 0.22972f
C10281 Iout.t232 VGND 0.02212f
C10282 Iout.n699 VGND 0.04919f
C10283 Iout.n700 VGND 0.02502f
C10284 Iout.n701 VGND 0.04584f
C10285 Iout.n702 VGND 0.22972f
C10286 Iout.n703 VGND 0.22972f
C10287 Iout.n704 VGND 0.04584f
C10288 Iout.t234 VGND 0.02212f
C10289 Iout.n705 VGND 0.04919f
C10290 Iout.n706 VGND 0.02502f
C10291 Iout.n707 VGND 0.04584f
C10292 Iout.n708 VGND 0.22972f
C10293 Iout.n709 VGND 0.22972f
C10294 Iout.n710 VGND 0.04584f
C10295 Iout.t158 VGND 0.02212f
C10296 Iout.n711 VGND 0.04919f
C10297 Iout.n712 VGND 0.02502f
C10298 Iout.n713 VGND 0.04584f
C10299 Iout.n714 VGND 0.22972f
C10300 Iout.n715 VGND 0.22972f
C10301 Iout.n716 VGND 0.04584f
C10302 Iout.t202 VGND 0.02212f
C10303 Iout.n717 VGND 0.04919f
C10304 Iout.n718 VGND 0.02502f
C10305 Iout.n719 VGND 0.04584f
C10306 Iout.n720 VGND 0.22972f
C10307 Iout.n721 VGND 0.22972f
C10308 Iout.n722 VGND 0.04584f
C10309 Iout.t149 VGND 0.02212f
C10310 Iout.n723 VGND 0.04919f
C10311 Iout.n724 VGND 0.02502f
C10312 Iout.n725 VGND 0.04584f
C10313 Iout.n726 VGND 0.22972f
C10314 Iout.n727 VGND 0.22972f
C10315 Iout.n728 VGND 0.04584f
C10316 Iout.t192 VGND 0.02212f
C10317 Iout.n729 VGND 0.04919f
C10318 Iout.n730 VGND 0.02502f
C10319 Iout.n731 VGND 0.04584f
C10320 Iout.n732 VGND 0.22972f
C10321 Iout.n733 VGND 0.22972f
C10322 Iout.n734 VGND 0.04584f
C10323 Iout.t105 VGND 0.02212f
C10324 Iout.n735 VGND 0.04919f
C10325 Iout.n736 VGND 0.02502f
C10326 Iout.n737 VGND 0.04584f
C10327 Iout.n738 VGND 0.22972f
C10328 Iout.n739 VGND 0.22972f
C10329 Iout.n740 VGND 0.04584f
C10330 Iout.t101 VGND 0.02212f
C10331 Iout.n741 VGND 0.04919f
C10332 Iout.n742 VGND 0.02502f
C10333 Iout.n743 VGND 0.04584f
C10334 Iout.n744 VGND 0.22972f
C10335 Iout.n745 VGND 0.22972f
C10336 Iout.n746 VGND 0.04584f
C10337 Iout.t1 VGND 0.02212f
C10338 Iout.n747 VGND 0.04919f
C10339 Iout.n748 VGND 0.02502f
C10340 Iout.n749 VGND 0.04584f
C10341 Iout.n750 VGND 0.22972f
C10342 Iout.n751 VGND 0.22972f
C10343 Iout.n752 VGND 0.04584f
C10344 Iout.t3 VGND 0.02212f
C10345 Iout.n753 VGND 0.04919f
C10346 Iout.n754 VGND 0.02502f
C10347 Iout.n755 VGND 0.04584f
C10348 Iout.n756 VGND 0.22972f
C10349 Iout.n757 VGND 0.22972f
C10350 Iout.n758 VGND 0.04584f
C10351 Iout.t77 VGND 0.02212f
C10352 Iout.n759 VGND 0.04919f
C10353 Iout.n760 VGND 0.02502f
C10354 Iout.n761 VGND 0.04584f
C10355 Iout.n762 VGND 0.22972f
C10356 Iout.n763 VGND 0.22972f
C10357 Iout.n764 VGND 0.04584f
C10358 Iout.t254 VGND 0.02212f
C10359 Iout.n765 VGND 0.04919f
C10360 Iout.n766 VGND 0.02502f
C10361 Iout.n767 VGND 0.04584f
C10362 Iout.n768 VGND 0.22972f
C10363 Iout.n769 VGND 0.22972f
C10364 Iout.n770 VGND 0.04584f
C10365 Iout.t38 VGND 0.02212f
C10366 Iout.n771 VGND 0.04919f
C10367 Iout.n772 VGND 0.02502f
C10368 Iout.n773 VGND 0.04584f
C10369 Iout.n774 VGND 0.22972f
C10370 Iout.n775 VGND 0.22972f
C10371 Iout.n776 VGND 0.04584f
C10372 Iout.t42 VGND 0.02212f
C10373 Iout.n777 VGND 0.04919f
C10374 Iout.n778 VGND 0.02502f
C10375 Iout.n779 VGND 0.04584f
C10376 Iout.n780 VGND 0.22972f
C10377 Iout.t83 VGND 0.02212f
C10378 Iout.n781 VGND 0.04919f
C10379 Iout.n782 VGND 0.02502f
C10380 Iout.n783 VGND 0.04584f
C10381 Iout.t104 VGND 0.02212f
C10382 Iout.n784 VGND 0.04919f
C10383 Iout.n785 VGND 0.02502f
C10384 Iout.n786 VGND 0.04584f
C10385 Iout.t147 VGND 0.02212f
C10386 Iout.n787 VGND 0.04919f
C10387 Iout.n788 VGND 0.02502f
C10388 Iout.n789 VGND 0.04584f
C10389 Iout.t178 VGND 0.02212f
C10390 Iout.n790 VGND 0.04919f
C10391 Iout.n791 VGND 0.02502f
C10392 Iout.n792 VGND 0.04584f
C10393 Iout.t235 VGND 0.02212f
C10394 Iout.n793 VGND 0.04919f
C10395 Iout.n794 VGND 0.02502f
C10396 Iout.n795 VGND 0.04584f
C10397 Iout.t115 VGND 0.02212f
C10398 Iout.n796 VGND 0.04919f
C10399 Iout.n797 VGND 0.02502f
C10400 Iout.n798 VGND 0.04584f
C10401 Iout.t199 VGND 0.02212f
C10402 Iout.n799 VGND 0.04919f
C10403 Iout.n800 VGND 0.02502f
C10404 Iout.n801 VGND 0.04584f
C10405 Iout.t20 VGND 0.02212f
C10406 Iout.n802 VGND 0.04919f
C10407 Iout.n803 VGND 0.02502f
C10408 Iout.n804 VGND 0.04584f
C10409 Iout.t31 VGND 0.02212f
C10410 Iout.n805 VGND 0.04919f
C10411 Iout.n806 VGND 0.02502f
C10412 Iout.n807 VGND 0.04584f
C10413 Iout.t191 VGND 0.02212f
C10414 Iout.n808 VGND 0.04919f
C10415 Iout.n809 VGND 0.02502f
C10416 Iout.n810 VGND 0.04584f
C10417 Iout.t208 VGND 0.02212f
C10418 Iout.n811 VGND 0.04919f
C10419 Iout.n812 VGND 0.02502f
C10420 Iout.n813 VGND 0.04584f
C10421 Iout.t78 VGND 0.02212f
C10422 Iout.n814 VGND 0.04919f
C10423 Iout.n815 VGND 0.02502f
C10424 Iout.n816 VGND 0.04584f
C10425 Iout.t231 VGND 0.02212f
C10426 Iout.n817 VGND 0.04919f
C10427 Iout.n818 VGND 0.02502f
C10428 Iout.n819 VGND 0.04584f
C10429 Iout.t65 VGND 0.02212f
C10430 Iout.n820 VGND 0.04919f
C10431 Iout.n821 VGND 0.02502f
C10432 Iout.n822 VGND 0.04584f
C10433 Iout.t74 VGND 0.02212f
C10434 Iout.n823 VGND 0.04919f
C10435 Iout.n824 VGND 0.02502f
C10436 Iout.n825 VGND 0.04584f
C10437 Iout.n826 VGND 0.22972f
C10438 Iout.t227 VGND 0.02212f
C10439 Iout.n827 VGND 0.04919f
C10440 Iout.n828 VGND 0.02502f
C10441 Iout.n829 VGND 0.07841f
C10442 Iout.n830 VGND 0.47625f
C10443 Iout.n831 VGND 0.04584f
C10444 Iout.t196 VGND 0.02212f
C10445 Iout.n832 VGND 0.04919f
C10446 Iout.n833 VGND 0.02502f
C10447 Iout.t35 VGND 0.02212f
C10448 Iout.n834 VGND 0.04919f
C10449 Iout.n835 VGND 0.02502f
C10450 Iout.n836 VGND 0.04584f
C10451 Iout.n837 VGND 0.47625f
C10452 Iout.n838 VGND 0.07841f
C10453 Iout.t9 VGND 0.02212f
C10454 Iout.n839 VGND 0.04919f
C10455 Iout.n840 VGND 0.02502f
C10456 Iout.t249 VGND 0.02212f
C10457 Iout.n841 VGND 0.04919f
C10458 Iout.n842 VGND 0.02502f
C10459 Iout.n843 VGND 0.07841f
C10460 Iout.n844 VGND 0.47625f
C10461 Iout.n845 VGND 0.04584f
C10462 Iout.t130 VGND 0.02212f
C10463 Iout.n846 VGND 0.04919f
C10464 Iout.n847 VGND 0.02502f
C10465 Iout.t165 VGND 0.02212f
C10466 Iout.n848 VGND 0.04919f
C10467 Iout.n849 VGND 0.02502f
C10468 Iout.n850 VGND 0.04584f
C10469 Iout.n851 VGND 0.47625f
C10470 Iout.n852 VGND 0.07841f
C10471 Iout.t89 VGND 0.02212f
C10472 Iout.n853 VGND 0.04919f
C10473 Iout.n854 VGND 0.02502f
C10474 Iout.t125 VGND 0.02212f
C10475 Iout.n855 VGND 0.04919f
C10476 Iout.n856 VGND 0.02502f
C10477 Iout.n857 VGND 0.07841f
C10478 Iout.n858 VGND 0.47625f
C10479 Iout.n859 VGND 0.04584f
C10480 Iout.t12 VGND 0.02212f
C10481 Iout.n860 VGND 0.04919f
C10482 Iout.n861 VGND 0.02502f
C10483 Iout.t253 VGND 0.02212f
C10484 Iout.n862 VGND 0.04919f
C10485 Iout.n863 VGND 0.02502f
C10486 Iout.n864 VGND 0.04584f
C10487 Iout.n865 VGND 0.47625f
C10488 Iout.n866 VGND 0.07841f
C10489 Iout.t103 VGND 0.02212f
C10490 Iout.n867 VGND 0.04919f
C10491 Iout.n868 VGND 0.02502f
C10492 Iout.t133 VGND 0.02212f
C10493 Iout.n869 VGND 0.04919f
C10494 Iout.n870 VGND 0.02502f
C10495 Iout.n871 VGND 0.07841f
C10496 Iout.n872 VGND 0.47625f
C10497 Iout.n873 VGND 0.04584f
C10498 Iout.t128 VGND 0.02212f
C10499 Iout.n874 VGND 0.04919f
C10500 Iout.n875 VGND 0.02502f
C10501 Iout.t159 VGND 0.02212f
C10502 Iout.n876 VGND 0.04919f
C10503 Iout.n877 VGND 0.02502f
C10504 Iout.n878 VGND 0.04584f
C10505 Iout.n879 VGND 0.47625f
C10506 Iout.n880 VGND 0.07841f
C10507 Iout.t28 VGND 0.02212f
C10508 Iout.n881 VGND 0.04919f
C10509 Iout.n882 VGND 0.02502f
C10510 Iout.t13 VGND 0.02212f
C10511 Iout.n883 VGND 0.04919f
C10512 Iout.n884 VGND 0.02502f
C10513 Iout.n885 VGND 0.07841f
C10514 Iout.n886 VGND 0.47625f
C10515 Iout.n887 VGND 0.04584f
C10516 Iout.t102 VGND 0.02212f
C10517 Iout.n888 VGND 0.04919f
C10518 Iout.n889 VGND 0.02502f
C10519 Iout.t163 VGND 0.02212f
C10520 Iout.n890 VGND 0.04919f
C10521 Iout.n891 VGND 0.02502f
C10522 Iout.n892 VGND 0.04584f
C10523 Iout.n893 VGND 0.47625f
C10524 Iout.n894 VGND 0.07841f
C10525 Iout.t245 VGND 0.02212f
C10526 Iout.n895 VGND 0.04919f
C10527 Iout.n896 VGND 0.02502f
C10528 Iout.t122 VGND 0.02212f
C10529 Iout.n897 VGND 0.04919f
C10530 Iout.n898 VGND 0.02502f
C10531 Iout.n899 VGND 0.07841f
C10532 Iout.n900 VGND 0.47625f
C10533 Iout.n901 VGND 0.04584f
C10534 Iout.t200 VGND 0.02212f
C10535 Iout.n902 VGND 0.04919f
C10536 Iout.n903 VGND 0.02502f
C10537 Iout.t57 VGND 0.02212f
C10538 Iout.n904 VGND 0.04919f
C10539 Iout.n905 VGND 0.02502f
C10540 Iout.n906 VGND 0.04584f
C10541 Iout.n907 VGND 0.47625f
C10542 Iout.n908 VGND 0.07841f
C10543 Iout.t99 VGND 0.02212f
C10544 Iout.n909 VGND 0.04919f
C10545 Iout.n910 VGND 0.02502f
C10546 Iout.t64 VGND 0.02212f
C10547 Iout.n911 VGND 0.04919f
C10548 Iout.n912 VGND 0.02502f
C10549 Iout.n913 VGND 0.07841f
C10550 Iout.n914 VGND 0.47625f
C10551 Iout.n915 VGND 0.04584f
C10552 Iout.t221 VGND 0.02212f
C10553 Iout.n916 VGND 0.04919f
C10554 Iout.n917 VGND 0.02502f
C10555 Iout.t148 VGND 0.02212f
C10556 Iout.n918 VGND 0.04919f
C10557 Iout.n919 VGND 0.02502f
C10558 Iout.n920 VGND 0.04584f
C10559 Iout.n921 VGND 0.47625f
C10560 Iout.n922 VGND 0.07841f
C10561 Iout.t121 VGND 0.02212f
C10562 Iout.n923 VGND 0.04919f
C10563 Iout.n924 VGND 0.02502f
C10564 Iout.n925 VGND 0.07841f
C10565 Iout.t50 VGND 0.02212f
C10566 Iout.n926 VGND 0.04919f
C10567 Iout.n927 VGND 0.02502f
C10568 Iout.n928 VGND 0.07841f
C10569 Iout.n929 VGND 0.47625f
C10570 Iout.n930 VGND 0.04584f
C10571 Iout.t2 VGND 0.02212f
C10572 Iout.n931 VGND 0.04919f
C10573 Iout.n932 VGND 0.02502f
C10574 Iout.n933 VGND 0.04584f
C10575 Iout.t0 VGND 0.02212f
C10576 Iout.n934 VGND 0.04919f
C10577 Iout.n935 VGND 0.19431f
C10578 Iout.n936 VGND 2.54526f
C10579 Iout.n937 VGND 1.20114f
C10580 Iout.t169 VGND 0.02212f
C10581 Iout.n938 VGND 0.04919f
C10582 Iout.n939 VGND 0.19431f
C10583 Iout.n940 VGND 0.04584f
C10584 Iout.n941 VGND 0.22972f
C10585 Iout.n942 VGND 0.22972f
C10586 Iout.n943 VGND 0.04584f
C10587 Iout.t179 VGND 0.02212f
C10588 Iout.n944 VGND 0.04919f
C10589 Iout.n945 VGND 0.02502f
C10590 Iout.n946 VGND 0.04584f
C10591 Iout.n947 VGND 0.22972f
C10592 Iout.n948 VGND 0.22972f
C10593 Iout.n949 VGND 0.04584f
C10594 Iout.t110 VGND 0.02212f
C10595 Iout.n950 VGND 0.04919f
C10596 Iout.n951 VGND 0.02502f
C10597 Iout.n952 VGND 0.04584f
C10598 Iout.t32 VGND 0.02212f
C10599 Iout.n953 VGND 0.04919f
C10600 Iout.n954 VGND 0.19431f
C10601 Iout.n955 VGND 1.20114f
C10602 Iout.n956 VGND 1.20114f
C10603 Iout.t93 VGND 0.02212f
C10604 Iout.n957 VGND 0.04919f
C10605 Iout.n958 VGND 0.19431f
C10606 Iout.n959 VGND 0.04584f
C10607 Iout.n960 VGND 0.22972f
C10608 Iout.n961 VGND 0.22972f
C10609 Iout.n962 VGND 0.04584f
C10610 Iout.t39 VGND 0.02212f
C10611 Iout.n963 VGND 0.04919f
C10612 Iout.n964 VGND 0.02502f
C10613 Iout.n965 VGND 0.04584f
C10614 Iout.n966 VGND 0.22972f
C10615 Iout.n967 VGND 0.22972f
C10616 Iout.n968 VGND 0.04584f
C10617 Iout.t124 VGND 0.02212f
C10618 Iout.n969 VGND 0.04919f
C10619 Iout.n970 VGND 0.02502f
C10620 Iout.n971 VGND 0.04584f
C10621 Iout.t63 VGND 0.02212f
C10622 Iout.n972 VGND 0.04919f
C10623 Iout.n973 VGND 0.19431f
C10624 Iout.n974 VGND 1.20114f
C10625 Iout.n975 VGND 1.20114f
C10626 Iout.t204 VGND 0.02212f
C10627 Iout.n976 VGND 0.04919f
C10628 Iout.n977 VGND 0.19431f
C10629 Iout.n978 VGND 0.04584f
C10630 Iout.n979 VGND 0.22972f
C10631 Iout.n980 VGND 0.22972f
C10632 Iout.n981 VGND 0.04584f
C10633 Iout.t45 VGND 0.02212f
C10634 Iout.n982 VGND 0.04919f
C10635 Iout.n983 VGND 0.02502f
C10636 Iout.n984 VGND 0.04584f
C10637 Iout.n985 VGND 0.22972f
C10638 Iout.n986 VGND 0.22972f
C10639 Iout.n987 VGND 0.04584f
C10640 Iout.t107 VGND 0.02212f
C10641 Iout.n988 VGND 0.04919f
C10642 Iout.n989 VGND 0.02502f
C10643 Iout.n990 VGND 0.04584f
C10644 Iout.t167 VGND 0.02212f
C10645 Iout.n991 VGND 0.04919f
C10646 Iout.n992 VGND 0.19431f
C10647 Iout.n993 VGND 1.20114f
C10648 Iout.n994 VGND 1.20114f
C10649 Iout.t242 VGND 0.02212f
C10650 Iout.n995 VGND 0.04919f
C10651 Iout.n996 VGND 0.19431f
C10652 Iout.n997 VGND 0.04584f
C10653 Iout.n998 VGND 0.22972f
C10654 Iout.n999 VGND 0.22972f
C10655 Iout.n1000 VGND 0.04584f
C10656 Iout.t123 VGND 0.02212f
C10657 Iout.n1001 VGND 0.04919f
C10658 Iout.n1002 VGND 0.02502f
C10659 Iout.n1003 VGND 0.04584f
C10660 Iout.n1004 VGND 0.22972f
C10661 Iout.n1005 VGND 0.22972f
C10662 Iout.n1006 VGND 0.04584f
C10663 Iout.t222 VGND 0.02212f
C10664 Iout.n1007 VGND 0.04919f
C10665 Iout.n1008 VGND 0.02502f
C10666 Iout.n1009 VGND 0.04584f
C10667 Iout.t203 VGND 0.02212f
C10668 Iout.n1010 VGND 0.04919f
C10669 Iout.n1011 VGND 0.19431f
C10670 Iout.n1012 VGND 1.20114f
C10671 Iout.n1013 VGND 1.07853f
C10672 Iout.t97 VGND 0.02212f
C10673 Iout.n1014 VGND 0.04919f
C10674 Iout.n1015 VGND 0.19431f
C10675 Iout.n1016 VGND 0.04584f
C10676 Iout.n1017 VGND 0.22972f
C10677 Iout.n1018 VGND 0.13561f
C10678 Iout.n1019 VGND 0.04584f
C10679 Iout.t100 VGND 0.02212f
C10680 Iout.n1020 VGND 0.04919f
C10681 Iout.n1021 VGND 0.19431f
C10682 Iout.n1022 VGND 0.22314f
C10683 VPWR.n0 VGND 0.03455f
C10684 VPWR.t760 VGND 0.21849f
C10685 VPWR.t726 VGND 0.09669f
C10686 VPWR.t895 VGND 0.27876f
C10687 VPWR.t890 VGND 0.10548f
C10688 VPWR.t1366 VGND 0.10548f
C10689 VPWR.t1346 VGND 0.10548f
C10690 VPWR.t622 VGND 0.10548f
C10691 VPWR.t1833 VGND 0.10548f
C10692 VPWR.t1829 VGND 0.10548f
C10693 VPWR.t626 VGND 0.07409f
C10694 VPWR.n1 VGND 0.1346f
C10695 VPWR.n2 VGND 0.07122f
C10696 VPWR.t727 VGND 0.04214f
C10697 VPWR.t627 VGND 0.01056f
C10698 VPWR.t1830 VGND 0.01056f
C10699 VPWR.n4 VGND 0.02319f
C10700 VPWR.t1834 VGND 0.01056f
C10701 VPWR.t623 VGND 0.01056f
C10702 VPWR.n5 VGND 0.02315f
C10703 VPWR.n6 VGND 0.04755f
C10704 VPWR.n7 VGND 0.13403f
C10705 VPWR.n8 VGND 0.04244f
C10706 VPWR.n9 VGND 0.03117f
C10707 VPWR.n10 VGND 0.05587f
C10708 VPWR.n12 VGND 0.01202f
C10709 VPWR.n13 VGND 0.01408f
C10710 VPWR.n14 VGND 0.02065f
C10711 VPWR.n15 VGND 0.06252f
C10712 VPWR.t761 VGND 0.04212f
C10713 VPWR.n17 VGND 0.05418f
C10714 VPWR.n18 VGND 0.24742f
C10715 VPWR.n19 VGND 0.72146f
C10716 VPWR.n20 VGND 0.79671f
C10717 VPWR.n21 VGND 0.0873f
C10718 VPWR.n22 VGND 0.06682f
C10719 VPWR.n23 VGND 0.12196f
C10720 VPWR.n24 VGND 0.07937f
C10721 VPWR.n25 VGND 0.07719f
C10722 VPWR.n26 VGND 0.09048f
C10723 VPWR.t494 VGND 0.03559f
C10724 VPWR.n27 VGND 0.13411f
C10725 VPWR.n28 VGND 0.13411f
C10726 VPWR.t493 VGND 0.9453f
C10727 VPWR.n29 VGND 0.13411f
C10728 VPWR.n30 VGND 0.13411f
C10729 VPWR.n31 VGND 0.07971f
C10730 VPWR.t1797 VGND 0.03559f
C10731 VPWR.n32 VGND 0.01995f
C10732 VPWR.n33 VGND 0.01662f
C10733 VPWR.n34 VGND 0.01648f
C10734 VPWR.n35 VGND 0.07937f
C10735 VPWR.n36 VGND 0.17591f
C10736 VPWR.n37 VGND 0.71129f
C10737 VPWR.n38 VGND 1.06417f
C10738 VPWR.n39 VGND 0.23484f
C10739 VPWR.n40 VGND 0.7488f
C10740 VPWR.n41 VGND 0.10237f
C10741 VPWR.n42 VGND 0.02207f
C10742 VPWR.n43 VGND 0.05863f
C10743 VPWR.n44 VGND 0.02207f
C10744 VPWR.n45 VGND 0.118f
C10745 VPWR.n46 VGND 0.02207f
C10746 VPWR.n47 VGND 0.09401f
C10747 VPWR.n48 VGND 0.02207f
C10748 VPWR.n49 VGND 0.09401f
C10749 VPWR.n50 VGND 0.02207f
C10750 VPWR.n51 VGND 0.09401f
C10751 VPWR.n52 VGND 0.02207f
C10752 VPWR.n53 VGND 0.09401f
C10753 VPWR.n54 VGND 0.02207f
C10754 VPWR.n55 VGND 0.09401f
C10755 VPWR.n56 VGND 0.02207f
C10756 VPWR.n57 VGND 0.09401f
C10757 VPWR.n58 VGND 0.02207f
C10758 VPWR.n59 VGND 0.09401f
C10759 VPWR.n60 VGND 0.02207f
C10760 VPWR.n61 VGND 0.09401f
C10761 VPWR.n62 VGND 0.02207f
C10762 VPWR.n63 VGND 0.09401f
C10763 VPWR.n64 VGND 0.02207f
C10764 VPWR.n65 VGND 0.09401f
C10765 VPWR.n66 VGND 0.02207f
C10766 VPWR.n67 VGND 0.09401f
C10767 VPWR.n68 VGND 0.02207f
C10768 VPWR.n69 VGND 0.09401f
C10769 VPWR.n70 VGND 0.02207f
C10770 VPWR.n71 VGND 0.09401f
C10771 VPWR.n72 VGND 0.02207f
C10772 VPWR.n73 VGND 0.10179f
C10773 VPWR.n74 VGND 0.08498f
C10774 VPWR.t1559 VGND 0.02456f
C10775 VPWR.t1664 VGND 0.02183f
C10776 VPWR.n75 VGND 0.06746f
C10777 VPWR.t1427 VGND 0.06796f
C10778 VPWR.t1434 VGND 0.02456f
C10779 VPWR.t1428 VGND 0.02183f
C10780 VPWR.n76 VGND 0.06746f
C10781 VPWR.n77 VGND 0.02534f
C10782 VPWR.n78 VGND 0.10257f
C10783 VPWR.n79 VGND 0.10257f
C10784 VPWR.n80 VGND 0.02534f
C10785 VPWR.t1415 VGND 0.02456f
C10786 VPWR.t1788 VGND 0.02183f
C10787 VPWR.n81 VGND 0.06746f
C10788 VPWR.t1654 VGND 0.06796f
C10789 VPWR.t1565 VGND 0.02456f
C10790 VPWR.t1655 VGND 0.02183f
C10791 VPWR.n82 VGND 0.06746f
C10792 VPWR.n83 VGND 0.02534f
C10793 VPWR.n84 VGND 0.10257f
C10794 VPWR.n85 VGND 0.10257f
C10795 VPWR.n86 VGND 0.02534f
C10796 VPWR.t1535 VGND 0.02456f
C10797 VPWR.t1527 VGND 0.02183f
C10798 VPWR.n87 VGND 0.06746f
C10799 VPWR.t1508 VGND 0.06796f
C10800 VPWR.t1791 VGND 0.02456f
C10801 VPWR.t1509 VGND 0.02183f
C10802 VPWR.n88 VGND 0.06746f
C10803 VPWR.n89 VGND 0.02534f
C10804 VPWR.n90 VGND 0.10257f
C10805 VPWR.n91 VGND 0.10257f
C10806 VPWR.n92 VGND 0.02534f
C10807 VPWR.t1661 VGND 0.02456f
C10808 VPWR.t1697 VGND 0.02183f
C10809 VPWR.n93 VGND 0.06746f
C10810 VPWR.t1631 VGND 0.06796f
C10811 VPWR.t1645 VGND 0.02456f
C10812 VPWR.t1632 VGND 0.02183f
C10813 VPWR.n94 VGND 0.06746f
C10814 VPWR.n95 VGND 0.02534f
C10815 VPWR.n96 VGND 0.10257f
C10816 VPWR.n97 VGND 0.10257f
C10817 VPWR.n98 VGND 0.02534f
C10818 VPWR.t1485 VGND 0.02456f
C10819 VPWR.t1504 VGND 0.02183f
C10820 VPWR.n99 VGND 0.06746f
C10821 VPWR.t1468 VGND 0.06796f
C10822 VPWR.t1764 VGND 0.02456f
C10823 VPWR.t1469 VGND 0.02183f
C10824 VPWR.n100 VGND 0.06746f
C10825 VPWR.n101 VGND 0.02534f
C10826 VPWR.n102 VGND 0.10257f
C10827 VPWR.n103 VGND 0.10257f
C10828 VPWR.n104 VGND 0.02534f
C10829 VPWR.t1608 VGND 0.02456f
C10830 VPWR.t1745 VGND 0.02183f
C10831 VPWR.n105 VGND 0.06746f
C10832 VPWR.t1589 VGND 0.06796f
C10833 VPWR.t1596 VGND 0.02456f
C10834 VPWR.t1590 VGND 0.02183f
C10835 VPWR.n106 VGND 0.06746f
C10836 VPWR.n107 VGND 0.02534f
C10837 VPWR.n108 VGND 0.10257f
C10838 VPWR.n109 VGND 0.10257f
C10839 VPWR.n110 VGND 0.02534f
C10840 VPWR.t1488 VGND 0.02456f
C10841 VPWR.t1482 VGND 0.02183f
C10842 VPWR.n111 VGND 0.06746f
C10843 VPWR.t1699 VGND 0.06796f
C10844 VPWR.t1726 VGND 0.02456f
C10845 VPWR.t1700 VGND 0.02183f
C10846 VPWR.n112 VGND 0.06746f
C10847 VPWR.n113 VGND 0.02534f
C10848 VPWR.n114 VGND 0.10257f
C10849 VPWR.n115 VGND 0.10257f
C10850 VPWR.n116 VGND 0.02534f
C10851 VPWR.t1611 VGND 0.02456f
C10852 VPWR.t1708 VGND 0.02183f
C10853 VPWR.n117 VGND 0.06746f
C10854 VPWR.t1465 VGND 0.10698f
C10855 VPWR.t1441 VGND 0.05786f
C10856 VPWR.t1572 VGND 0.06796f
C10857 VPWR.t1466 VGND 0.02456f
C10858 VPWR.t1573 VGND 0.02183f
C10859 VPWR.n118 VGND 0.06746f
C10860 VPWR.n119 VGND 0.02206f
C10861 VPWR.n120 VGND 0.02421f
C10862 VPWR.n122 VGND 0.01343f
C10863 VPWR.n123 VGND 0.02206f
C10864 VPWR.n124 VGND 0.02421f
C10865 VPWR.n125 VGND 0.02297f
C10866 VPWR.n126 VGND 0.01452f
C10867 VPWR.n127 VGND 0.0204f
C10868 VPWR.n128 VGND 0.02077f
C10869 VPWR.n129 VGND 0.01309f
C10870 VPWR.n131 VGND 0.01343f
C10871 VPWR.n132 VGND 0.01957f
C10872 VPWR.n133 VGND 0.02206f
C10873 VPWR.n134 VGND 0.02421f
C10874 VPWR.n135 VGND 0.02297f
C10875 VPWR.n136 VGND 0.02723f
C10876 VPWR.n138 VGND 0.0204f
C10877 VPWR.n139 VGND 0.02077f
C10878 VPWR.n140 VGND 0.01309f
C10879 VPWR.n142 VGND 0.01343f
C10880 VPWR.n143 VGND 0.01873f
C10881 VPWR.n144 VGND 0.02206f
C10882 VPWR.n145 VGND 0.02421f
C10883 VPWR.n146 VGND 0.02297f
C10884 VPWR.n147 VGND 0.02723f
C10885 VPWR.n149 VGND 0.0204f
C10886 VPWR.n150 VGND 0.02077f
C10887 VPWR.n151 VGND 0.01309f
C10888 VPWR.n153 VGND 0.01343f
C10889 VPWR.n154 VGND 0.01757f
C10890 VPWR.n155 VGND 0.15601f
C10891 VPWR.n156 VGND 0.02206f
C10892 VPWR.n157 VGND 0.02421f
C10893 VPWR.n158 VGND 0.02297f
C10894 VPWR.n159 VGND 0.02723f
C10895 VPWR.n161 VGND 0.0204f
C10896 VPWR.n162 VGND 0.02077f
C10897 VPWR.n163 VGND 0.01309f
C10898 VPWR.n165 VGND 0.01343f
C10899 VPWR.n166 VGND 0.01757f
C10900 VPWR.n167 VGND 0.12963f
C10901 VPWR.n168 VGND 0.02206f
C10902 VPWR.n169 VGND 0.02421f
C10903 VPWR.n170 VGND 0.02297f
C10904 VPWR.n171 VGND 0.02723f
C10905 VPWR.n173 VGND 0.0204f
C10906 VPWR.n174 VGND 0.02077f
C10907 VPWR.n175 VGND 0.01309f
C10908 VPWR.n177 VGND 0.01343f
C10909 VPWR.n178 VGND 0.01757f
C10910 VPWR.n179 VGND 0.12963f
C10911 VPWR.n180 VGND 0.02206f
C10912 VPWR.n181 VGND 0.02421f
C10913 VPWR.n182 VGND 0.02297f
C10914 VPWR.n183 VGND 0.02723f
C10915 VPWR.n185 VGND 0.0204f
C10916 VPWR.n186 VGND 0.02077f
C10917 VPWR.n187 VGND 0.01309f
C10918 VPWR.n189 VGND 0.01343f
C10919 VPWR.n190 VGND 0.01757f
C10920 VPWR.n191 VGND 0.12963f
C10921 VPWR.n192 VGND 0.02206f
C10922 VPWR.n193 VGND 0.02421f
C10923 VPWR.n194 VGND 0.02297f
C10924 VPWR.n195 VGND 0.02723f
C10925 VPWR.n197 VGND 0.0204f
C10926 VPWR.n198 VGND 0.02077f
C10927 VPWR.n199 VGND 0.01309f
C10928 VPWR.n201 VGND 0.01343f
C10929 VPWR.n202 VGND 0.01757f
C10930 VPWR.n203 VGND 0.12963f
C10931 VPWR.n204 VGND 0.02206f
C10932 VPWR.n205 VGND 0.02421f
C10933 VPWR.n206 VGND 0.02297f
C10934 VPWR.n207 VGND 0.02723f
C10935 VPWR.n209 VGND 0.0204f
C10936 VPWR.n210 VGND 0.02077f
C10937 VPWR.n211 VGND 0.01309f
C10938 VPWR.n213 VGND 0.01343f
C10939 VPWR.n214 VGND 0.01757f
C10940 VPWR.n215 VGND 0.12963f
C10941 VPWR.n216 VGND 0.02206f
C10942 VPWR.n217 VGND 0.02421f
C10943 VPWR.n218 VGND 0.02297f
C10944 VPWR.n219 VGND 0.02723f
C10945 VPWR.n221 VGND 0.0204f
C10946 VPWR.n222 VGND 0.02077f
C10947 VPWR.n223 VGND 0.01309f
C10948 VPWR.n225 VGND 0.01343f
C10949 VPWR.n226 VGND 0.01757f
C10950 VPWR.n227 VGND 0.12963f
C10951 VPWR.n228 VGND 0.02206f
C10952 VPWR.n229 VGND 0.02421f
C10953 VPWR.n230 VGND 0.02297f
C10954 VPWR.n231 VGND 0.02723f
C10955 VPWR.n233 VGND 0.0204f
C10956 VPWR.n234 VGND 0.02077f
C10957 VPWR.n235 VGND 0.01309f
C10958 VPWR.n237 VGND 0.01343f
C10959 VPWR.n238 VGND 0.01757f
C10960 VPWR.n239 VGND 0.12963f
C10961 VPWR.n240 VGND 0.02206f
C10962 VPWR.n241 VGND 0.02421f
C10963 VPWR.n242 VGND 0.02297f
C10964 VPWR.n243 VGND 0.02723f
C10965 VPWR.n245 VGND 0.0204f
C10966 VPWR.n246 VGND 0.02077f
C10967 VPWR.n247 VGND 0.01309f
C10968 VPWR.n249 VGND 0.01343f
C10969 VPWR.n250 VGND 0.01757f
C10970 VPWR.n251 VGND 0.12963f
C10971 VPWR.n252 VGND 0.02206f
C10972 VPWR.n253 VGND 0.02421f
C10973 VPWR.n254 VGND 0.02297f
C10974 VPWR.n255 VGND 0.02723f
C10975 VPWR.n257 VGND 0.0204f
C10976 VPWR.n258 VGND 0.02077f
C10977 VPWR.n259 VGND 0.01309f
C10978 VPWR.n261 VGND 0.01343f
C10979 VPWR.n262 VGND 0.01757f
C10980 VPWR.n263 VGND 0.12963f
C10981 VPWR.n264 VGND 0.02206f
C10982 VPWR.n265 VGND 0.02421f
C10983 VPWR.n266 VGND 0.02297f
C10984 VPWR.n267 VGND 0.02723f
C10985 VPWR.n269 VGND 0.0204f
C10986 VPWR.n270 VGND 0.02077f
C10987 VPWR.n271 VGND 0.01309f
C10988 VPWR.n273 VGND 0.01343f
C10989 VPWR.n274 VGND 0.01757f
C10990 VPWR.n275 VGND 0.12963f
C10991 VPWR.n276 VGND 0.02206f
C10992 VPWR.n277 VGND 0.02421f
C10993 VPWR.n278 VGND 0.02297f
C10994 VPWR.n279 VGND 0.02723f
C10995 VPWR.n281 VGND 0.0204f
C10996 VPWR.n282 VGND 0.02077f
C10997 VPWR.n283 VGND 0.01309f
C10998 VPWR.n285 VGND 0.01343f
C10999 VPWR.n286 VGND 0.01757f
C11000 VPWR.n287 VGND 0.12963f
C11001 VPWR.n288 VGND 0.02206f
C11002 VPWR.n289 VGND 0.02421f
C11003 VPWR.n290 VGND 0.02297f
C11004 VPWR.n291 VGND 0.02723f
C11005 VPWR.n293 VGND 0.0204f
C11006 VPWR.n294 VGND 0.02077f
C11007 VPWR.n295 VGND 0.01309f
C11008 VPWR.n297 VGND 0.01343f
C11009 VPWR.n298 VGND 0.01757f
C11010 VPWR.n299 VGND 0.12963f
C11011 VPWR.n300 VGND 0.17489f
C11012 VPWR.n301 VGND 0.01757f
C11013 VPWR.n302 VGND 0.01309f
C11014 VPWR.n303 VGND 0.0204f
C11015 VPWR.n304 VGND 0.02077f
C11016 VPWR.n306 VGND 0.02297f
C11017 VPWR.n307 VGND 0.02723f
C11018 VPWR.n308 VGND 0.02534f
C11019 VPWR.t584 VGND 0.02456f
C11020 VPWR.t789 VGND 0.02183f
C11021 VPWR.n309 VGND 0.06746f
C11022 VPWR.t583 VGND 0.10698f
C11023 VPWR.t1218 VGND 0.05786f
C11024 VPWR.t788 VGND 0.06796f
C11025 VPWR.t1256 VGND 0.02456f
C11026 VPWR.t1772 VGND 0.02183f
C11027 VPWR.n310 VGND 0.06746f
C11028 VPWR.n311 VGND 0.01325f
C11029 VPWR.n312 VGND 0.05616f
C11030 VPWR.t1771 VGND 0.09829f
C11031 VPWR.t1214 VGND 0.05786f
C11032 VPWR.t1255 VGND 0.08814f
C11033 VPWR.t986 VGND 0.02456f
C11034 VPWR.t1226 VGND 0.02183f
C11035 VPWR.n313 VGND 0.06746f
C11036 VPWR.n314 VGND 0.01325f
C11037 VPWR.n316 VGND 0.07978f
C11038 VPWR.t1225 VGND 0.06796f
C11039 VPWR.t812 VGND 0.05786f
C11040 VPWR.t985 VGND 0.08814f
C11041 VPWR.t1309 VGND 0.02456f
C11042 VPWR.t992 VGND 0.02183f
C11043 VPWR.n317 VGND 0.06746f
C11044 VPWR.n318 VGND 0.01325f
C11045 VPWR.n320 VGND 0.07978f
C11046 VPWR.t991 VGND 0.06796f
C11047 VPWR.t741 VGND 0.05786f
C11048 VPWR.t1308 VGND 0.08814f
C11049 VPWR.t69 VGND 0.02456f
C11050 VPWR.t178 VGND 0.02183f
C11051 VPWR.n321 VGND 0.06746f
C11052 VPWR.n322 VGND 0.01325f
C11053 VPWR.n324 VGND 0.07978f
C11054 VPWR.t177 VGND 0.06796f
C11055 VPWR.t742 VGND 0.05786f
C11056 VPWR.t68 VGND 0.08814f
C11057 VPWR.t479 VGND 0.02456f
C11058 VPWR.t1026 VGND 0.02183f
C11059 VPWR.n325 VGND 0.06746f
C11060 VPWR.n326 VGND 0.01325f
C11061 VPWR.n328 VGND 0.07978f
C11062 VPWR.t1025 VGND 0.06796f
C11063 VPWR.t1219 VGND 0.05786f
C11064 VPWR.t478 VGND 0.08814f
C11065 VPWR.t388 VGND 0.02456f
C11066 VPWR.t485 VGND 0.02183f
C11067 VPWR.n329 VGND 0.06746f
C11068 VPWR.n330 VGND 0.01325f
C11069 VPWR.n332 VGND 0.07978f
C11070 VPWR.t484 VGND 0.06796f
C11071 VPWR.t809 VGND 0.05786f
C11072 VPWR.t387 VGND 0.08814f
C11073 VPWR.t668 VGND 0.02456f
C11074 VPWR.t361 VGND 0.02183f
C11075 VPWR.n333 VGND 0.06746f
C11076 VPWR.n334 VGND 0.01325f
C11077 VPWR.n336 VGND 0.07978f
C11078 VPWR.t360 VGND 0.06796f
C11079 VPWR.t745 VGND 0.05786f
C11080 VPWR.t667 VGND 0.08814f
C11081 VPWR.t546 VGND 0.02456f
C11082 VPWR.t1280 VGND 0.02183f
C11083 VPWR.n337 VGND 0.06746f
C11084 VPWR.n338 VGND 0.01325f
C11085 VPWR.n340 VGND 0.07978f
C11086 VPWR.t1279 VGND 0.06796f
C11087 VPWR.t1215 VGND 0.05786f
C11088 VPWR.t545 VGND 0.08814f
C11089 VPWR.t1377 VGND 0.02456f
C11090 VPWR.t613 VGND 0.02183f
C11091 VPWR.n341 VGND 0.06746f
C11092 VPWR.n342 VGND 0.01325f
C11093 VPWR.n344 VGND 0.07978f
C11094 VPWR.t612 VGND 0.06796f
C11095 VPWR.t1216 VGND 0.05786f
C11096 VPWR.t1376 VGND 0.08814f
C11097 VPWR.t1816 VGND 0.02456f
C11098 VPWR.t1383 VGND 0.02183f
C11099 VPWR.n345 VGND 0.06746f
C11100 VPWR.n346 VGND 0.01325f
C11101 VPWR.n348 VGND 0.07978f
C11102 VPWR.t1382 VGND 0.06796f
C11103 VPWR.t743 VGND 0.05786f
C11104 VPWR.t1815 VGND 0.08814f
C11105 VPWR.t1213 VGND 0.02456f
C11106 VPWR.t1822 VGND 0.02183f
C11107 VPWR.n349 VGND 0.06746f
C11108 VPWR.n350 VGND 0.01325f
C11109 VPWR.n352 VGND 0.07978f
C11110 VPWR.t1821 VGND 0.06796f
C11111 VPWR.t744 VGND 0.05786f
C11112 VPWR.t1212 VGND 0.08814f
C11113 VPWR.t9 VGND 0.02456f
C11114 VPWR.t902 VGND 0.02183f
C11115 VPWR.n353 VGND 0.06746f
C11116 VPWR.n354 VGND 0.01325f
C11117 VPWR.n356 VGND 0.07978f
C11118 VPWR.t901 VGND 0.06796f
C11119 VPWR.t1217 VGND 0.05786f
C11120 VPWR.t8 VGND 0.08814f
C11121 VPWR.t1068 VGND 0.02456f
C11122 VPWR.t674 VGND 0.02183f
C11123 VPWR.n357 VGND 0.06746f
C11124 VPWR.n358 VGND 0.01325f
C11125 VPWR.n360 VGND 0.07978f
C11126 VPWR.t673 VGND 0.06796f
C11127 VPWR.t810 VGND 0.05786f
C11128 VPWR.t1067 VGND 0.08814f
C11129 VPWR.t1272 VGND 0.02456f
C11130 VPWR.t1044 VGND 0.02183f
C11131 VPWR.n361 VGND 0.06746f
C11132 VPWR.n362 VGND 0.01325f
C11133 VPWR.n364 VGND 0.07978f
C11134 VPWR.t1043 VGND 0.06796f
C11135 VPWR.t811 VGND 0.05786f
C11136 VPWR.t1271 VGND 0.08814f
C11137 VPWR.t842 VGND 0.02456f
C11138 VPWR.t1113 VGND 0.02183f
C11139 VPWR.n365 VGND 0.06746f
C11140 VPWR.n366 VGND 0.01325f
C11141 VPWR.n368 VGND 0.07978f
C11142 VPWR.t1112 VGND 0.06796f
C11143 VPWR.t746 VGND 0.05786f
C11144 VPWR.t841 VGND 0.08814f
C11145 VPWR.n369 VGND 0.07978f
C11146 VPWR.n371 VGND 0.01325f
C11147 VPWR.n372 VGND 0.10257f
C11148 VPWR.n373 VGND 0.74411f
C11149 VPWR.n374 VGND 0.10257f
C11150 VPWR.t578 VGND 0.02456f
C11151 VPWR.t662 VGND 0.02183f
C11152 VPWR.n375 VGND 0.06746f
C11153 VPWR.t577 VGND 0.10698f
C11154 VPWR.t1362 VGND 0.05786f
C11155 VPWR.t661 VGND 0.06796f
C11156 VPWR.t1116 VGND 0.08814f
C11157 VPWR.t785 VGND 0.02456f
C11158 VPWR.t1335 VGND 0.02183f
C11159 VPWR.n376 VGND 0.06746f
C11160 VPWR.n377 VGND 0.10257f
C11161 VPWR.n378 VGND 0.10257f
C11162 VPWR.t1117 VGND 0.02456f
C11163 VPWR.t1036 VGND 0.02183f
C11164 VPWR.n379 VGND 0.06746f
C11165 VPWR.t883 VGND 0.05786f
C11166 VPWR.t1035 VGND 0.06796f
C11167 VPWR.t753 VGND 0.08814f
C11168 VPWR.t1060 VGND 0.02456f
C11169 VPWR.t1397 VGND 0.02183f
C11170 VPWR.n380 VGND 0.06746f
C11171 VPWR.n381 VGND 0.10257f
C11172 VPWR.n382 VGND 0.10257f
C11173 VPWR.t754 VGND 0.02456f
C11174 VPWR.t1146 VGND 0.02183f
C11175 VPWR.n383 VGND 0.06746f
C11176 VPWR.t1361 VGND 0.05786f
C11177 VPWR.t1145 VGND 0.06796f
C11178 VPWR.t1825 VGND 0.08814f
C11179 VPWR.t906 VGND 0.02456f
C11180 VPWR.t1802 VGND 0.02183f
C11181 VPWR.n384 VGND 0.06746f
C11182 VPWR.n385 VGND 0.10257f
C11183 VPWR.n386 VGND 0.10257f
C11184 VPWR.t1826 VGND 0.02456f
C11185 VPWR.t1393 VGND 0.02183f
C11186 VPWR.n387 VGND 0.06746f
C11187 VPWR.t887 VGND 0.05786f
C11188 VPWR.t1392 VGND 0.06796f
C11189 VPWR.t238 VGND 0.08814f
C11190 VPWR.t1387 VGND 0.02456f
C11191 VPWR.t939 VGND 0.02183f
C11192 VPWR.n388 VGND 0.06746f
C11193 VPWR.n389 VGND 0.10257f
C11194 VPWR.n390 VGND 0.10257f
C11195 VPWR.t239 VGND 0.02456f
C11196 VPWR.t296 VGND 0.02183f
C11197 VPWR.n391 VGND 0.06746f
C11198 VPWR.t1359 VGND 0.05786f
C11199 VPWR.t295 VGND 0.06796f
C11200 VPWR.t356 VGND 0.08814f
C11201 VPWR.t1284 VGND 0.02456f
C11202 VPWR.t367 VGND 0.02183f
C11203 VPWR.n392 VGND 0.06746f
C11204 VPWR.n393 VGND 0.10257f
C11205 VPWR.n394 VGND 0.10257f
C11206 VPWR.t357 VGND 0.02456f
C11207 VPWR.t1844 VGND 0.02183f
C11208 VPWR.n395 VGND 0.06746f
C11209 VPWR.t1208 VGND 0.05786f
C11210 VPWR.t1843 VGND 0.06796f
C11211 VPWR.t632 VGND 0.08814f
C11212 VPWR.t489 VGND 0.02456f
C11213 VPWR.t1885 VGND 0.02183f
C11214 VPWR.n396 VGND 0.06746f
C11215 VPWR.n397 VGND 0.10257f
C11216 VPWR.n398 VGND 0.10257f
C11217 VPWR.t633 VGND 0.02456f
C11218 VPWR.t188 VGND 0.02183f
C11219 VPWR.n399 VGND 0.06746f
C11220 VPWR.t886 VGND 0.05786f
C11221 VPWR.t187 VGND 0.06796f
C11222 VPWR.t987 VGND 0.08814f
C11223 VPWR.t1315 VGND 0.02456f
C11224 VPWR.t980 VGND 0.02183f
C11225 VPWR.n400 VGND 0.06746f
C11226 VPWR.n401 VGND 0.10257f
C11227 VPWR.n402 VGND 0.10257f
C11228 VPWR.t988 VGND 0.02456f
C11229 VPWR.t1238 VGND 0.02183f
C11230 VPWR.n403 VGND 0.06746f
C11231 VPWR.t884 VGND 0.05786f
C11232 VPWR.t1237 VGND 0.06796f
C11233 VPWR.t828 VGND 0.02456f
C11234 VPWR.t1735 VGND 0.02183f
C11235 VPWR.n404 VGND 0.06746f
C11236 VPWR.t1248 VGND 0.02456f
C11237 VPWR.t1447 VGND 0.02183f
C11238 VPWR.n405 VGND 0.06746f
C11239 VPWR.t587 VGND 0.10698f
C11240 VPWR.t923 VGND 0.05786f
C11241 VPWR.t837 VGND 0.06796f
C11242 VPWR.t588 VGND 0.02456f
C11243 VPWR.t838 VGND 0.02183f
C11244 VPWR.n406 VGND 0.06746f
C11245 VPWR.n407 VGND 0.01325f
C11246 VPWR.n409 VGND 0.07978f
C11247 VPWR.t74 VGND 0.08814f
C11248 VPWR.t1190 VGND 0.05786f
C11249 VPWR.t708 VGND 0.06796f
C11250 VPWR.t75 VGND 0.02456f
C11251 VPWR.t709 VGND 0.02183f
C11252 VPWR.n410 VGND 0.06746f
C11253 VPWR.n411 VGND 0.01325f
C11254 VPWR.n413 VGND 0.07978f
C11255 VPWR.t1155 VGND 0.08814f
C11256 VPWR.t706 VGND 0.05786f
C11257 VPWR.t1053 VGND 0.06796f
C11258 VPWR.t1156 VGND 0.02456f
C11259 VPWR.t1054 VGND 0.02183f
C11260 VPWR.n414 VGND 0.06746f
C11261 VPWR.n415 VGND 0.01325f
C11262 VPWR.n417 VGND 0.07978f
C11263 VPWR.t1077 VGND 0.08814f
C11264 VPWR.t705 VGND 0.05786f
C11265 VPWR.t757 VGND 0.06796f
C11266 VPWR.t1078 VGND 0.02456f
C11267 VPWR.t758 VGND 0.02183f
C11268 VPWR.n418 VGND 0.06746f
C11269 VPWR.n419 VGND 0.01325f
C11270 VPWR.n421 VGND 0.07978f
C11271 VPWR.t689 VGND 0.08814f
C11272 VPWR.t922 VGND 0.05786f
C11273 VPWR.t1182 VGND 0.06796f
C11274 VPWR.t690 VGND 0.02456f
C11275 VPWR.t1183 VGND 0.02183f
C11276 VPWR.n422 VGND 0.06746f
C11277 VPWR.n423 VGND 0.01325f
C11278 VPWR.n425 VGND 0.07978f
C11279 VPWR.t1327 VGND 0.08814f
C11280 VPWR.t915 VGND 0.05786f
C11281 VPWR.t847 VGND 0.06796f
C11282 VPWR.t1328 VGND 0.02456f
C11283 VPWR.t848 VGND 0.02183f
C11284 VPWR.n426 VGND 0.06746f
C11285 VPWR.n427 VGND 0.01325f
C11286 VPWR.n429 VGND 0.07978f
C11287 VPWR.t1103 VGND 0.08814f
C11288 VPWR.t914 VGND 0.05786f
C11289 VPWR.t1909 VGND 0.06796f
C11290 VPWR.t1104 VGND 0.02456f
C11291 VPWR.t1910 VGND 0.02183f
C11292 VPWR.n430 VGND 0.06746f
C11293 VPWR.n431 VGND 0.01325f
C11294 VPWR.n433 VGND 0.07978f
C11295 VPWR.t1903 VGND 0.08814f
C11296 VPWR.t921 VGND 0.05786f
C11297 VPWR.t232 VGND 0.06796f
C11298 VPWR.t1904 VGND 0.02456f
C11299 VPWR.t233 VGND 0.02183f
C11300 VPWR.n434 VGND 0.06746f
C11301 VPWR.n435 VGND 0.01325f
C11302 VPWR.n437 VGND 0.07978f
C11303 VPWR.t1925 VGND 0.08814f
C11304 VPWR.t920 VGND 0.05786f
C11305 VPWR.t156 VGND 0.06796f
C11306 VPWR.t1926 VGND 0.02456f
C11307 VPWR.t157 VGND 0.02183f
C11308 VPWR.n438 VGND 0.06746f
C11309 VPWR.n439 VGND 0.01325f
C11310 VPWR.n441 VGND 0.07978f
C11311 VPWR.t798 VGND 0.08814f
C11312 VPWR.t916 VGND 0.05786f
C11313 VPWR.t383 VGND 0.06796f
C11314 VPWR.t799 VGND 0.02456f
C11315 VPWR.t384 VGND 0.02183f
C11316 VPWR.n442 VGND 0.06746f
C11317 VPWR.n443 VGND 0.01325f
C11318 VPWR.n445 VGND 0.07978f
C11319 VPWR.t350 VGND 0.08814f
C11320 VPWR.t704 VGND 0.05786f
C11321 VPWR.t1126 VGND 0.06796f
C11322 VPWR.t351 VGND 0.02456f
C11323 VPWR.t1127 VGND 0.02183f
C11324 VPWR.n446 VGND 0.06746f
C11325 VPWR.n447 VGND 0.01325f
C11326 VPWR.n449 VGND 0.07978f
C11327 VPWR.t1120 VGND 0.08814f
C11328 VPWR.t703 VGND 0.05786f
C11329 VPWR.t1813 VGND 0.06796f
C11330 VPWR.t1121 VGND 0.02456f
C11331 VPWR.t1814 VGND 0.02183f
C11332 VPWR.n450 VGND 0.06746f
C11333 VPWR.n451 VGND 0.01325f
C11334 VPWR.n453 VGND 0.07978f
C11335 VPWR.t1807 VGND 0.08814f
C11336 VPWR.t913 VGND 0.05786f
C11337 VPWR.t399 VGND 0.06796f
C11338 VPWR.t1808 VGND 0.02456f
C11339 VPWR.t400 VGND 0.02183f
C11340 VPWR.n454 VGND 0.06746f
C11341 VPWR.n455 VGND 0.01325f
C11342 VPWR.n457 VGND 0.07978f
C11343 VPWR.t258 VGND 0.08814f
C11344 VPWR.t912 VGND 0.05786f
C11345 VPWR.t1199 VGND 0.06796f
C11346 VPWR.t259 VGND 0.02456f
C11347 VPWR.t1200 VGND 0.02183f
C11348 VPWR.n458 VGND 0.06746f
C11349 VPWR.n459 VGND 0.01325f
C11350 VPWR.n461 VGND 0.07978f
C11351 VPWR.t1193 VGND 0.08814f
C11352 VPWR.t911 VGND 0.05786f
C11353 VPWR.t831 VGND 0.06796f
C11354 VPWR.t1194 VGND 0.02456f
C11355 VPWR.t832 VGND 0.02183f
C11356 VPWR.n462 VGND 0.06746f
C11357 VPWR.n463 VGND 0.01325f
C11358 VPWR.n465 VGND 0.07978f
C11359 VPWR.t1247 VGND 0.08814f
C11360 VPWR.t919 VGND 0.05786f
C11361 VPWR.t1446 VGND 0.09829f
C11362 VPWR.n466 VGND 0.05616f
C11363 VPWR.n467 VGND 0.01325f
C11364 VPWR.n468 VGND 0.10257f
C11365 VPWR.n469 VGND 0.7488f
C11366 VPWR.n470 VGND 0.10257f
C11367 VPWR.t21 VGND 0.02456f
C11368 VPWR.t1562 VGND 0.02183f
C11369 VPWR.n471 VGND 0.06746f
C11370 VPWR.t1249 VGND 0.06796f
C11371 VPWR.t1006 VGND 0.02456f
C11372 VPWR.t1250 VGND 0.02183f
C11373 VPWR.n472 VGND 0.06746f
C11374 VPWR.n473 VGND 0.10257f
C11375 VPWR.n474 VGND 0.10257f
C11376 VPWR.t194 VGND 0.02456f
C11377 VPWR.t1014 VGND 0.02183f
C11378 VPWR.n475 VGND 0.06746f
C11379 VPWR.t1302 VGND 0.06796f
C11380 VPWR.t1868 VGND 0.02456f
C11381 VPWR.t1303 VGND 0.02183f
C11382 VPWR.n476 VGND 0.06746f
C11383 VPWR.n477 VGND 0.10257f
C11384 VPWR.n478 VGND 0.10257f
C11385 VPWR.t1202 VGND 0.02456f
C11386 VPWR.t1022 VGND 0.02183f
C11387 VPWR.n479 VGND 0.06746f
C11388 VPWR.t1205 VGND 0.06796f
C11389 VPWR.t335 VGND 0.02456f
C11390 VPWR.t1206 VGND 0.02183f
C11391 VPWR.n480 VGND 0.06746f
C11392 VPWR.n481 VGND 0.10257f
C11393 VPWR.n482 VGND 0.10257f
C11394 VPWR.t654 VGND 0.02456f
C11395 VPWR.t343 VGND 0.02183f
C11396 VPWR.n483 VGND 0.06746f
C11397 VPWR.t560 VGND 0.06796f
C11398 VPWR.t953 VGND 0.02456f
C11399 VPWR.t561 VGND 0.02183f
C11400 VPWR.n484 VGND 0.06746f
C11401 VPWR.n485 VGND 0.10257f
C11402 VPWR.n486 VGND 0.10257f
C11403 VPWR.t455 VGND 0.02456f
C11404 VPWR.t1930 VGND 0.02183f
C11405 VPWR.n487 VGND 0.06746f
C11406 VPWR.t458 VGND 0.06796f
C11407 VPWR.t859 VGND 0.02456f
C11408 VPWR.t459 VGND 0.02183f
C11409 VPWR.n488 VGND 0.06746f
C11410 VPWR.n489 VGND 0.10257f
C11411 VPWR.n490 VGND 0.10257f
C11412 VPWR.t1264 VGND 0.02456f
C11413 VPWR.t863 VGND 0.02183f
C11414 VPWR.n491 VGND 0.06746f
C11415 VPWR.t443 VGND 0.06796f
C11416 VPWR.t406 VGND 0.02456f
C11417 VPWR.t444 VGND 0.02183f
C11418 VPWR.n492 VGND 0.06746f
C11419 VPWR.n493 VGND 0.10257f
C11420 VPWR.n494 VGND 0.10257f
C11421 VPWR.t1094 VGND 0.02456f
C11422 VPWR.t692 VGND 0.02183f
C11423 VPWR.n495 VGND 0.06746f
C11424 VPWR.t1071 VGND 0.06796f
C11425 VPWR.t1919 VGND 0.02456f
C11426 VPWR.t1072 VGND 0.02183f
C11427 VPWR.n496 VGND 0.06746f
C11428 VPWR.n497 VGND 0.10257f
C11429 VPWR.n498 VGND 0.10257f
C11430 VPWR.t499 VGND 0.02456f
C11431 VPWR.t505 VGND 0.02183f
C11432 VPWR.n499 VGND 0.06746f
C11433 VPWR.t595 VGND 0.10698f
C11434 VPWR.t138 VGND 0.05786f
C11435 VPWR.t644 VGND 0.06796f
C11436 VPWR.t596 VGND 0.02456f
C11437 VPWR.t645 VGND 0.02183f
C11438 VPWR.n500 VGND 0.06746f
C11439 VPWR.t586 VGND 0.02456f
C11440 VPWR.t787 VGND 0.02183f
C11441 VPWR.n501 VGND 0.06746f
C11442 VPWR.t585 VGND 0.10698f
C11443 VPWR.t1879 VGND 0.05786f
C11444 VPWR.t786 VGND 0.06796f
C11445 VPWR.t1254 VGND 0.02456f
C11446 VPWR.t1780 VGND 0.02183f
C11447 VPWR.n502 VGND 0.06746f
C11448 VPWR.n503 VGND 0.01325f
C11449 VPWR.n504 VGND 0.05616f
C11450 VPWR.t1779 VGND 0.09829f
C11451 VPWR.t1221 VGND 0.05786f
C11452 VPWR.t1253 VGND 0.08814f
C11453 VPWR.t984 VGND 0.02456f
C11454 VPWR.t1224 VGND 0.02183f
C11455 VPWR.n505 VGND 0.06746f
C11456 VPWR.n506 VGND 0.01325f
C11457 VPWR.n508 VGND 0.07978f
C11458 VPWR.t1223 VGND 0.06796f
C11459 VPWR.t853 VGND 0.05786f
C11460 VPWR.t983 VGND 0.08814f
C11461 VPWR.t1305 VGND 0.02456f
C11462 VPWR.t990 VGND 0.02183f
C11463 VPWR.n509 VGND 0.06746f
C11464 VPWR.n510 VGND 0.01325f
C11465 VPWR.n512 VGND 0.07978f
C11466 VPWR.t989 VGND 0.06796f
C11467 VPWR.t1329 VGND 0.05786f
C11468 VPWR.t1304 VGND 0.08814f
C11469 VPWR.t67 VGND 0.02456f
C11470 VPWR.t975 VGND 0.02183f
C11471 VPWR.n513 VGND 0.06746f
C11472 VPWR.n514 VGND 0.01325f
C11473 VPWR.n516 VGND 0.07978f
C11474 VPWR.t974 VGND 0.06796f
C11475 VPWR.t1330 VGND 0.05786f
C11476 VPWR.t66 VGND 0.08814f
C11477 VPWR.t477 VGND 0.02456f
C11478 VPWR.t1024 VGND 0.02183f
C11479 VPWR.n517 VGND 0.06746f
C11480 VPWR.n518 VGND 0.01325f
C11481 VPWR.n520 VGND 0.07978f
C11482 VPWR.t1023 VGND 0.06796f
C11483 VPWR.t1880 VGND 0.05786f
C11484 VPWR.t476 VGND 0.08814f
C11485 VPWR.t386 VGND 0.02456f
C11486 VPWR.t481 VGND 0.02183f
C11487 VPWR.n521 VGND 0.06746f
C11488 VPWR.n522 VGND 0.01325f
C11489 VPWR.n524 VGND 0.07978f
C11490 VPWR.t480 VGND 0.06796f
C11491 VPWR.t1881 VGND 0.05786f
C11492 VPWR.t385 VGND 0.08814f
C11493 VPWR.t666 VGND 0.02456f
C11494 VPWR.t359 VGND 0.02183f
C11495 VPWR.n525 VGND 0.06746f
C11496 VPWR.n526 VGND 0.01325f
C11497 VPWR.n528 VGND 0.07978f
C11498 VPWR.t358 VGND 0.06796f
C11499 VPWR.t1333 VGND 0.05786f
C11500 VPWR.t665 VGND 0.08814f
C11501 VPWR.t542 VGND 0.02456f
C11502 VPWR.t670 VGND 0.02183f
C11503 VPWR.n529 VGND 0.06746f
C11504 VPWR.n530 VGND 0.01325f
C11505 VPWR.n532 VGND 0.07978f
C11506 VPWR.t669 VGND 0.06796f
C11507 VPWR.t1222 VGND 0.05786f
C11508 VPWR.t541 VGND 0.08814f
C11509 VPWR.t1912 VGND 0.02456f
C11510 VPWR.t609 VGND 0.02183f
C11511 VPWR.n533 VGND 0.06746f
C11512 VPWR.n534 VGND 0.01325f
C11513 VPWR.n536 VGND 0.07978f
C11514 VPWR.t608 VGND 0.06796f
C11515 VPWR.t1877 VGND 0.05786f
C11516 VPWR.t1911 VGND 0.08814f
C11517 VPWR.t850 VGND 0.02456f
C11518 VPWR.t1379 VGND 0.02183f
C11519 VPWR.n537 VGND 0.06746f
C11520 VPWR.n538 VGND 0.01325f
C11521 VPWR.n540 VGND 0.07978f
C11522 VPWR.t1378 VGND 0.06796f
C11523 VPWR.t1331 VGND 0.05786f
C11524 VPWR.t849 VGND 0.08814f
C11525 VPWR.t1211 VGND 0.02456f
C11526 VPWR.t1818 VGND 0.02183f
C11527 VPWR.n541 VGND 0.06746f
C11528 VPWR.n542 VGND 0.01325f
C11529 VPWR.n544 VGND 0.07978f
C11530 VPWR.t1817 VGND 0.06796f
C11531 VPWR.t1332 VGND 0.05786f
C11532 VPWR.t1210 VGND 0.08814f
C11533 VPWR.t7 VGND 0.02456f
C11534 VPWR.t898 VGND 0.02183f
C11535 VPWR.n545 VGND 0.06746f
C11536 VPWR.n546 VGND 0.01325f
C11537 VPWR.n548 VGND 0.07978f
C11538 VPWR.t897 VGND 0.06796f
C11539 VPWR.t1878 VGND 0.05786f
C11540 VPWR.t6 VGND 0.08814f
C11541 VPWR.t1070 VGND 0.02456f
C11542 VPWR.t672 VGND 0.02183f
C11543 VPWR.n549 VGND 0.06746f
C11544 VPWR.n550 VGND 0.01325f
C11545 VPWR.n552 VGND 0.07978f
C11546 VPWR.t671 VGND 0.06796f
C11547 VPWR.t851 VGND 0.05786f
C11548 VPWR.t1069 VGND 0.08814f
C11549 VPWR.t1270 VGND 0.02456f
C11550 VPWR.t1046 VGND 0.02183f
C11551 VPWR.n553 VGND 0.06746f
C11552 VPWR.n554 VGND 0.01325f
C11553 VPWR.n556 VGND 0.07978f
C11554 VPWR.t1045 VGND 0.06796f
C11555 VPWR.t852 VGND 0.05786f
C11556 VPWR.t1269 VGND 0.08814f
C11557 VPWR.t840 VGND 0.02456f
C11558 VPWR.t1274 VGND 0.02183f
C11559 VPWR.n557 VGND 0.06746f
C11560 VPWR.n558 VGND 0.01325f
C11561 VPWR.n560 VGND 0.07978f
C11562 VPWR.t1273 VGND 0.06796f
C11563 VPWR.t1220 VGND 0.05786f
C11564 VPWR.t839 VGND 0.08814f
C11565 VPWR.n561 VGND 0.07978f
C11566 VPWR.n563 VGND 0.01325f
C11567 VPWR.n564 VGND 0.10257f
C11568 VPWR.n565 VGND 0.74411f
C11569 VPWR.n566 VGND 0.10257f
C11570 VPWR.t572 VGND 0.02456f
C11571 VPWR.t292 VGND 0.02183f
C11572 VPWR.n567 VGND 0.06746f
C11573 VPWR.t571 VGND 0.10698f
C11574 VPWR.t1353 VGND 0.05786f
C11575 VPWR.t291 VGND 0.06796f
C11576 VPWR.t1188 VGND 0.08814f
C11577 VPWR.t736 VGND 0.02456f
C11578 VPWR.t517 VGND 0.02183f
C11579 VPWR.n568 VGND 0.06746f
C11580 VPWR.n569 VGND 0.10257f
C11581 VPWR.n570 VGND 0.10257f
C11582 VPWR.t1189 VGND 0.02456f
C11583 VPWR.t1084 VGND 0.02183f
C11584 VPWR.n571 VGND 0.06746f
C11585 VPWR.t1338 VGND 0.05786f
C11586 VPWR.t1083 VGND 0.06796f
C11587 VPWR.t681 VGND 0.08814f
C11588 VPWR.t1048 VGND 0.02456f
C11589 VPWR.t414 VGND 0.02183f
C11590 VPWR.n572 VGND 0.06746f
C11591 VPWR.n573 VGND 0.10257f
C11592 VPWR.n574 VGND 0.10257f
C11593 VPWR.t682 VGND 0.02456f
C11594 VPWR.t153 VGND 0.02183f
C11595 VPWR.n575 VGND 0.06746f
C11596 VPWR.t1352 VGND 0.05786f
C11597 VPWR.t152 VGND 0.06796f
C11598 VPWR.t52 VGND 0.08814f
C11599 VPWR.t145 VGND 0.02456f
C11600 VPWR.t61 VGND 0.02183f
C11601 VPWR.n576 VGND 0.06746f
C11602 VPWR.n577 VGND 0.10257f
C11603 VPWR.n578 VGND 0.10257f
C11604 VPWR.t53 VGND 0.02456f
C11605 VPWR.t723 VGND 0.02183f
C11606 VPWR.n579 VGND 0.06746f
C11607 VPWR.t1342 VGND 0.05786f
C11608 VPWR.t722 VGND 0.06796f
C11609 VPWR.t930 VGND 0.08814f
C11610 VPWR.t715 VGND 0.02456f
C11611 VPWR.t219 VGND 0.02183f
C11612 VPWR.n580 VGND 0.06746f
C11613 VPWR.n581 VGND 0.10257f
C11614 VPWR.n582 VGND 0.10257f
C11615 VPWR.t931 VGND 0.02456f
C11616 VPWR.t527 VGND 0.02183f
C11617 VPWR.n583 VGND 0.06746f
C11618 VPWR.t1350 VGND 0.05786f
C11619 VPWR.t526 VGND 0.06796f
C11620 VPWR.t322 VGND 0.08814f
C11621 VPWR.t47 VGND 0.02456f
C11622 VPWR.t331 VGND 0.02183f
C11623 VPWR.n584 VGND 0.06746f
C11624 VPWR.n585 VGND 0.10257f
C11625 VPWR.n586 VGND 0.10257f
C11626 VPWR.t323 VGND 0.02456f
C11627 VPWR.t555 VGND 0.02183f
C11628 VPWR.n587 VGND 0.06746f
C11629 VPWR.t867 VGND 0.05786f
C11630 VPWR.t554 VGND 0.06796f
C11631 VPWR.t1873 VGND 0.08814f
C11632 VPWR.t781 VGND 0.02456f
C11633 VPWR.t1864 VGND 0.02183f
C11634 VPWR.n588 VGND 0.06746f
C11635 VPWR.n589 VGND 0.10257f
C11636 VPWR.n590 VGND 0.10257f
C11637 VPWR.t1874 VGND 0.02456f
C11638 VPWR.t251 VGND 0.02183f
C11639 VPWR.n591 VGND 0.06746f
C11640 VPWR.t1341 VGND 0.05786f
C11641 VPWR.t250 VGND 0.06796f
C11642 VPWR.t530 VGND 0.08814f
C11643 VPWR.t180 VGND 0.02456f
C11644 VPWR.t641 VGND 0.02183f
C11645 VPWR.n592 VGND 0.06746f
C11646 VPWR.n593 VGND 0.10257f
C11647 VPWR.n594 VGND 0.10257f
C11648 VPWR.t531 VGND 0.02456f
C11649 VPWR.t13 VGND 0.02183f
C11650 VPWR.n595 VGND 0.06746f
C11651 VPWR.t1339 VGND 0.05786f
C11652 VPWR.t12 VGND 0.06796f
C11653 VPWR.t1234 VGND 0.02456f
C11654 VPWR.t1629 VGND 0.02183f
C11655 VPWR.n596 VGND 0.06746f
C11656 VPWR.t824 VGND 0.02456f
C11657 VPWR.t1740 VGND 0.02183f
C11658 VPWR.n597 VGND 0.06746f
C11659 VPWR.t579 VGND 0.10698f
C11660 VPWR.t303 VGND 0.05786f
C11661 VPWR.t792 VGND 0.06796f
C11662 VPWR.t580 VGND 0.02456f
C11663 VPWR.t793 VGND 0.02183f
C11664 VPWR.n598 VGND 0.06746f
C11665 VPWR.n599 VGND 0.01325f
C11666 VPWR.n601 VGND 0.07978f
C11667 VPWR.t782 VGND 0.08814f
C11668 VPWR.t437 VGND 0.05786f
C11669 VPWR.t909 VGND 0.06796f
C11670 VPWR.t783 VGND 0.02456f
C11671 VPWR.t910 VGND 0.02183f
C11672 VPWR.n602 VGND 0.06746f
C11673 VPWR.n603 VGND 0.01325f
C11674 VPWR.n605 VGND 0.07978f
C11675 VPWR.t1114 VGND 0.08814f
C11676 VPWR.t440 VGND 0.05786f
C11677 VPWR.t1037 VGND 0.06796f
C11678 VPWR.t1115 VGND 0.02456f
C11679 VPWR.t1038 VGND 0.02183f
C11680 VPWR.n606 VGND 0.06746f
C11681 VPWR.n607 VGND 0.01325f
C11682 VPWR.n609 VGND 0.07978f
C11683 VPWR.t1061 VGND 0.08814f
C11684 VPWR.t439 VGND 0.05786f
C11685 VPWR.t683 VGND 0.06796f
C11686 VPWR.t1062 VGND 0.02456f
C11687 VPWR.t684 VGND 0.02183f
C11688 VPWR.n610 VGND 0.06746f
C11689 VPWR.n611 VGND 0.01325f
C11690 VPWR.n613 VGND 0.07978f
C11691 VPWR.t749 VGND 0.08814f
C11692 VPWR.t302 VGND 0.05786f
C11693 VPWR.t1143 VGND 0.06796f
C11694 VPWR.t750 VGND 0.02456f
C11695 VPWR.t1144 VGND 0.02183f
C11696 VPWR.n614 VGND 0.06746f
C11697 VPWR.n615 VGND 0.01325f
C11698 VPWR.n617 VGND 0.07978f
C11699 VPWR.t903 VGND 0.08814f
C11700 VPWR.t435 VGND 0.05786f
C11701 VPWR.t1799 VGND 0.06796f
C11702 VPWR.t904 VGND 0.02456f
C11703 VPWR.t1800 VGND 0.02183f
C11704 VPWR.n618 VGND 0.06746f
C11705 VPWR.n619 VGND 0.01325f
C11706 VPWR.n621 VGND 0.07978f
C11707 VPWR.t1823 VGND 0.08814f
C11708 VPWR.t434 VGND 0.05786f
C11709 VPWR.t1390 VGND 0.06796f
C11710 VPWR.t1824 VGND 0.02456f
C11711 VPWR.t1391 VGND 0.02183f
C11712 VPWR.n622 VGND 0.06746f
C11713 VPWR.n623 VGND 0.01325f
C11714 VPWR.n625 VGND 0.07978f
C11715 VPWR.t1384 VGND 0.08814f
C11716 VPWR.t301 VGND 0.05786f
C11717 VPWR.t936 VGND 0.06796f
C11718 VPWR.t1385 VGND 0.02456f
C11719 VPWR.t937 VGND 0.02183f
C11720 VPWR.n626 VGND 0.06746f
C11721 VPWR.n627 VGND 0.01325f
C11722 VPWR.n629 VGND 0.07978f
C11723 VPWR.t236 VGND 0.08814f
C11724 VPWR.t300 VGND 0.05786f
C11725 VPWR.t1287 VGND 0.06796f
C11726 VPWR.t237 VGND 0.02456f
C11727 VPWR.t1288 VGND 0.02183f
C11728 VPWR.n630 VGND 0.06746f
C11729 VPWR.n631 VGND 0.01325f
C11730 VPWR.n633 VGND 0.07978f
C11731 VPWR.t1281 VGND 0.08814f
C11732 VPWR.t436 VGND 0.05786f
C11733 VPWR.t364 VGND 0.06796f
C11734 VPWR.t1282 VGND 0.02456f
C11735 VPWR.t365 VGND 0.02183f
C11736 VPWR.n634 VGND 0.06746f
C11737 VPWR.n635 VGND 0.01325f
C11738 VPWR.n637 VGND 0.07978f
C11739 VPWR.t354 VGND 0.08814f
C11740 VPWR.t305 VGND 0.05786f
C11741 VPWR.t1841 VGND 0.06796f
C11742 VPWR.t355 VGND 0.02456f
C11743 VPWR.t1842 VGND 0.02183f
C11744 VPWR.n638 VGND 0.06746f
C11745 VPWR.n639 VGND 0.01325f
C11746 VPWR.n641 VGND 0.07978f
C11747 VPWR.t486 VGND 0.08814f
C11748 VPWR.t304 VGND 0.05786f
C11749 VPWR.t1029 VGND 0.06796f
C11750 VPWR.t487 VGND 0.02456f
C11751 VPWR.t1030 VGND 0.02183f
C11752 VPWR.n642 VGND 0.06746f
C11753 VPWR.n643 VGND 0.01325f
C11754 VPWR.n645 VGND 0.07978f
C11755 VPWR.t630 VGND 0.08814f
C11756 VPWR.t433 VGND 0.05786f
C11757 VPWR.t185 VGND 0.06796f
C11758 VPWR.t631 VGND 0.02456f
C11759 VPWR.t186 VGND 0.02183f
C11760 VPWR.n646 VGND 0.06746f
C11761 VPWR.n647 VGND 0.01325f
C11762 VPWR.n649 VGND 0.07978f
C11763 VPWR.t1312 VGND 0.08814f
C11764 VPWR.t432 VGND 0.05786f
C11765 VPWR.t995 VGND 0.06796f
C11766 VPWR.t1313 VGND 0.02456f
C11767 VPWR.t996 VGND 0.02183f
C11768 VPWR.n650 VGND 0.06746f
C11769 VPWR.n651 VGND 0.01325f
C11770 VPWR.n653 VGND 0.07978f
C11771 VPWR.t601 VGND 0.08814f
C11772 VPWR.t431 VGND 0.05786f
C11773 VPWR.t1235 VGND 0.06796f
C11774 VPWR.t602 VGND 0.02456f
C11775 VPWR.t1236 VGND 0.02183f
C11776 VPWR.n654 VGND 0.06746f
C11777 VPWR.n655 VGND 0.01325f
C11778 VPWR.n657 VGND 0.07978f
C11779 VPWR.t823 VGND 0.08814f
C11780 VPWR.t438 VGND 0.05786f
C11781 VPWR.t1739 VGND 0.09829f
C11782 VPWR.n658 VGND 0.05616f
C11783 VPWR.n659 VGND 0.01325f
C11784 VPWR.n660 VGND 0.10257f
C11785 VPWR.n661 VGND 0.7488f
C11786 VPWR.n662 VGND 0.10257f
C11787 VPWR.t17 VGND 0.02456f
C11788 VPWR.t1463 VGND 0.02183f
C11789 VPWR.n663 VGND 0.06746f
C11790 VPWR.t825 VGND 0.06796f
C11791 VPWR.t1000 VGND 0.02456f
C11792 VPWR.t826 VGND 0.02183f
C11793 VPWR.n664 VGND 0.06746f
C11794 VPWR.n665 VGND 0.10257f
C11795 VPWR.n666 VGND 0.10257f
C11796 VPWR.t255 VGND 0.02456f
C11797 VPWR.t1196 VGND 0.02183f
C11798 VPWR.n667 VGND 0.06746f
C11799 VPWR.t1316 VGND 0.06796f
C11800 VPWR.t1164 VGND 0.02456f
C11801 VPWR.t1317 VGND 0.02183f
C11802 VPWR.n668 VGND 0.06746f
C11803 VPWR.n669 VGND 0.10257f
C11804 VPWR.n670 VGND 0.10257f
C11805 VPWR.t1410 VGND 0.02456f
C11806 VPWR.t1810 VGND 0.02183f
C11807 VPWR.n671 VGND 0.06746f
C11808 VPWR.t1122 VGND 0.06796f
C11809 VPWR.t347 VGND 0.02456f
C11810 VPWR.t1123 VGND 0.02183f
C11811 VPWR.n672 VGND 0.06746f
C11812 VPWR.n673 VGND 0.10257f
C11813 VPWR.n674 VGND 0.10257f
C11814 VPWR.t795 VGND 0.02456f
C11815 VPWR.t353 VGND 0.02183f
C11816 VPWR.n675 VGND 0.06746f
C11817 VPWR.t800 VGND 0.06796f
C11818 VPWR.t223 VGND 0.02456f
C11819 VPWR.t801 VGND 0.02183f
C11820 VPWR.n676 VGND 0.06746f
C11821 VPWR.n677 VGND 0.10257f
C11822 VPWR.n678 VGND 0.10257f
C11823 VPWR.t1900 VGND 0.02456f
C11824 VPWR.t241 VGND 0.02183f
C11825 VPWR.n679 VGND 0.06746f
C11826 VPWR.t1905 VGND 0.06796f
C11827 VPWR.t1100 VGND 0.02456f
C11828 VPWR.t1906 VGND 0.02183f
C11829 VPWR.n680 VGND 0.06746f
C11830 VPWR.n681 VGND 0.10257f
C11831 VPWR.n682 VGND 0.10257f
C11832 VPWR.t1324 VGND 0.02456f
C11833 VPWR.t844 VGND 0.02183f
C11834 VPWR.n683 VGND 0.06746f
C11835 VPWR.t1178 VGND 0.06796f
C11836 VPWR.t418 VGND 0.02456f
C11837 VPWR.t1179 VGND 0.02183f
C11838 VPWR.n684 VGND 0.06746f
C11839 VPWR.n685 VGND 0.10257f
C11840 VPWR.n686 VGND 0.10257f
C11841 VPWR.t1082 VGND 0.02456f
C11842 VPWR.t752 VGND 0.02183f
C11843 VPWR.n687 VGND 0.06746f
C11844 VPWR.t1057 VGND 0.06796f
C11845 VPWR.t1152 VGND 0.02456f
C11846 VPWR.t1058 VGND 0.02183f
C11847 VPWR.n688 VGND 0.06746f
C11848 VPWR.n689 VGND 0.10257f
C11849 VPWR.n690 VGND 0.10257f
C11850 VPWR.t71 VGND 0.02456f
C11851 VPWR.t1158 VGND 0.02183f
C11852 VPWR.n691 VGND 0.06746f
C11853 VPWR.t591 VGND 0.10698f
C11854 VPWR.t702 VGND 0.05786f
C11855 VPWR.t648 VGND 0.06796f
C11856 VPWR.t592 VGND 0.02456f
C11857 VPWR.t649 VGND 0.02183f
C11858 VPWR.n692 VGND 0.06746f
C11859 VPWR.t598 VGND 0.02456f
C11860 VPWR.t503 VGND 0.02183f
C11861 VPWR.n693 VGND 0.06746f
C11862 VPWR.t597 VGND 0.10698f
C11863 VPWR.t1265 VGND 0.05786f
C11864 VPWR.t502 VGND 0.06796f
C11865 VPWR.t19 VGND 0.02456f
C11866 VPWR.t1570 VGND 0.02183f
C11867 VPWR.n694 VGND 0.06746f
C11868 VPWR.n695 VGND 0.01325f
C11869 VPWR.n696 VGND 0.05616f
C11870 VPWR.t1569 VGND 0.09829f
C11871 VPWR.t1192 VGND 0.05786f
C11872 VPWR.t18 VGND 0.08814f
C11873 VPWR.t1004 VGND 0.02456f
C11874 VPWR.t1246 VGND 0.02183f
C11875 VPWR.n697 VGND 0.06746f
C11876 VPWR.n698 VGND 0.01325f
C11877 VPWR.n700 VGND 0.07978f
C11878 VPWR.t1245 VGND 0.06796f
C11879 VPWR.t1375 VGND 0.05786f
C11880 VPWR.t1003 VGND 0.08814f
C11881 VPWR.t192 VGND 0.02456f
C11882 VPWR.t1010 VGND 0.02183f
C11883 VPWR.n701 VGND 0.06746f
C11884 VPWR.n702 VGND 0.01325f
C11885 VPWR.n704 VGND 0.07978f
C11886 VPWR.t1009 VGND 0.06796f
C11887 VPWR.t869 VGND 0.05786f
C11888 VPWR.t191 VGND 0.08814f
C11889 VPWR.t1866 VGND 0.02456f
C11890 VPWR.t1301 VGND 0.02183f
C11891 VPWR.n705 VGND 0.06746f
C11892 VPWR.n706 VGND 0.01325f
C11893 VPWR.n708 VGND 0.07978f
C11894 VPWR.t1300 VGND 0.06796f
C11895 VPWR.t870 VGND 0.05786f
C11896 VPWR.t1865 VGND 0.08814f
C11897 VPWR.t559 VGND 0.02456f
C11898 VPWR.t1018 VGND 0.02183f
C11899 VPWR.n709 VGND 0.06746f
C11900 VPWR.n710 VGND 0.01325f
C11901 VPWR.n712 VGND 0.07978f
C11902 VPWR.t1017 VGND 0.06796f
C11903 VPWR.t1266 VGND 0.05786f
C11904 VPWR.t558 VGND 0.08814f
C11905 VPWR.t333 VGND 0.02456f
C11906 VPWR.t1204 VGND 0.02183f
C11907 VPWR.n713 VGND 0.06746f
C11908 VPWR.n714 VGND 0.01325f
C11909 VPWR.n716 VGND 0.07978f
C11910 VPWR.t1203 VGND 0.06796f
C11911 VPWR.t1267 VGND 0.05786f
C11912 VPWR.t332 VGND 0.08814f
C11913 VPWR.t652 VGND 0.02456f
C11914 VPWR.t339 VGND 0.02183f
C11915 VPWR.n717 VGND 0.06746f
C11916 VPWR.n718 VGND 0.01325f
C11917 VPWR.n720 VGND 0.07978f
C11918 VPWR.t338 VGND 0.06796f
C11919 VPWR.t873 VGND 0.05786f
C11920 VPWR.t651 VGND 0.08814f
C11921 VPWR.t951 VGND 0.02456f
C11922 VPWR.t656 VGND 0.02183f
C11923 VPWR.n721 VGND 0.06746f
C11924 VPWR.n722 VGND 0.01325f
C11925 VPWR.n724 VGND 0.07978f
C11926 VPWR.t655 VGND 0.06796f
C11927 VPWR.t547 VGND 0.05786f
C11928 VPWR.t950 VGND 0.08814f
C11929 VPWR.t453 VGND 0.02456f
C11930 VPWR.t1928 VGND 0.02183f
C11931 VPWR.n725 VGND 0.06746f
C11932 VPWR.n726 VGND 0.01325f
C11933 VPWR.n728 VGND 0.07978f
C11934 VPWR.t1927 VGND 0.06796f
C11935 VPWR.t1149 VGND 0.05786f
C11936 VPWR.t452 VGND 0.08814f
C11937 VPWR.t65 VGND 0.02456f
C11938 VPWR.t457 VGND 0.02183f
C11939 VPWR.n729 VGND 0.06746f
C11940 VPWR.n730 VGND 0.01325f
C11941 VPWR.n732 VGND 0.07978f
C11942 VPWR.t456 VGND 0.06796f
C11943 VPWR.t871 VGND 0.05786f
C11944 VPWR.t64 VGND 0.08814f
C11945 VPWR.t1262 VGND 0.02456f
C11946 VPWR.t861 VGND 0.02183f
C11947 VPWR.n733 VGND 0.06746f
C11948 VPWR.n734 VGND 0.01325f
C11949 VPWR.n736 VGND 0.07978f
C11950 VPWR.t860 VGND 0.06796f
C11951 VPWR.t872 VGND 0.05786f
C11952 VPWR.t1261 VGND 0.08814f
C11953 VPWR.t1403 VGND 0.02456f
C11954 VPWR.t442 VGND 0.02183f
C11955 VPWR.n737 VGND 0.06746f
C11956 VPWR.n738 VGND 0.01325f
C11957 VPWR.n740 VGND 0.07978f
C11958 VPWR.t441 VGND 0.06796f
C11959 VPWR.t1150 VGND 0.05786f
C11960 VPWR.t1402 VGND 0.08814f
C11961 VPWR.t1096 VGND 0.02456f
C11962 VPWR.t688 VGND 0.02183f
C11963 VPWR.n741 VGND 0.06746f
C11964 VPWR.n742 VGND 0.01325f
C11965 VPWR.n744 VGND 0.07978f
C11966 VPWR.t687 VGND 0.06796f
C11967 VPWR.t1373 VGND 0.05786f
C11968 VPWR.t1095 VGND 0.08814f
C11969 VPWR.t1917 VGND 0.02456f
C11970 VPWR.t1074 VGND 0.02183f
C11971 VPWR.n745 VGND 0.06746f
C11972 VPWR.n746 VGND 0.01325f
C11973 VPWR.n748 VGND 0.07978f
C11974 VPWR.t1073 VGND 0.06796f
C11975 VPWR.t1374 VGND 0.05786f
C11976 VPWR.t1916 VGND 0.08814f
C11977 VPWR.t294 VGND 0.02456f
C11978 VPWR.t1921 VGND 0.02183f
C11979 VPWR.n749 VGND 0.06746f
C11980 VPWR.n750 VGND 0.01325f
C11981 VPWR.n752 VGND 0.07978f
C11982 VPWR.t1920 VGND 0.06796f
C11983 VPWR.t1191 VGND 0.05786f
C11984 VPWR.t293 VGND 0.08814f
C11985 VPWR.n753 VGND 0.07978f
C11986 VPWR.n755 VGND 0.01325f
C11987 VPWR.n756 VGND 0.10257f
C11988 VPWR.n757 VGND 0.74411f
C11989 VPWR.n758 VGND 0.10257f
C11990 VPWR.t594 VGND 0.02456f
C11991 VPWR.t647 VGND 0.02183f
C11992 VPWR.n759 VGND 0.06746f
C11993 VPWR.t593 VGND 0.10698f
C11994 VPWR.t808 VGND 0.05786f
C11995 VPWR.t646 VGND 0.06796f
C11996 VPWR.t506 VGND 0.08814f
C11997 VPWR.t643 VGND 0.02456f
C11998 VPWR.t509 VGND 0.02183f
C11999 VPWR.n760 VGND 0.06746f
C12000 VPWR.n761 VGND 0.10257f
C12001 VPWR.n762 VGND 0.10257f
C12002 VPWR.t507 VGND 0.02456f
C12003 VPWR.t1066 VGND 0.02183f
C12004 VPWR.n763 VGND 0.06746f
C12005 VPWR.t968 VGND 0.05786f
C12006 VPWR.t1065 VGND 0.06796f
C12007 VPWR.t407 VGND 0.08814f
C12008 VPWR.t1090 VGND 0.02456f
C12009 VPWR.t5 VGND 0.02183f
C12010 VPWR.n764 VGND 0.06746f
C12011 VPWR.n765 VGND 0.10257f
C12012 VPWR.n766 VGND 0.10257f
C12013 VPWR.t408 VGND 0.02456f
C12014 VPWR.t448 VGND 0.02183f
C12015 VPWR.n767 VGND 0.06746f
C12016 VPWR.t807 VGND 0.05786f
C12017 VPWR.t447 VGND 0.06796f
C12018 VPWR.t864 VGND 0.08814f
C12019 VPWR.t446 VGND 0.02456f
C12020 VPWR.t1098 VGND 0.02183f
C12021 VPWR.n768 VGND 0.06746f
C12022 VPWR.n769 VGND 0.10257f
C12023 VPWR.n770 VGND 0.10257f
C12024 VPWR.t865 VGND 0.02456f
C12025 VPWR.t463 VGND 0.02183f
C12026 VPWR.n771 VGND 0.06746f
C12027 VPWR.t1031 VGND 0.05786f
C12028 VPWR.t462 VGND 0.06796f
C12029 VPWR.t226 VGND 0.08814f
C12030 VPWR.t461 VGND 0.02456f
C12031 VPWR.t544 VGND 0.02183f
C12032 VPWR.n772 VGND 0.06746f
C12033 VPWR.n773 VGND 0.10257f
C12034 VPWR.n774 VGND 0.10257f
C12035 VPWR.t227 VGND 0.02456f
C12036 VPWR.t565 VGND 0.02183f
C12037 VPWR.n775 VGND 0.06746f
C12038 VPWR.t805 VGND 0.05786f
C12039 VPWR.t564 VGND 0.06796f
C12040 VPWR.t340 VGND 0.08814f
C12041 VPWR.t563 VGND 0.02456f
C12042 VPWR.t345 VGND 0.02183f
C12043 VPWR.n776 VGND 0.06746f
C12044 VPWR.n777 VGND 0.10257f
C12045 VPWR.n778 VGND 0.10257f
C12046 VPWR.t341 VGND 0.02456f
C12047 VPWR.t1408 VGND 0.02183f
C12048 VPWR.n779 VGND 0.06746f
C12049 VPWR.t966 VGND 0.05786f
C12050 VPWR.t1407 VGND 0.06796f
C12051 VPWR.t1019 VGND 0.08814f
C12052 VPWR.t533 VGND 0.02456f
C12053 VPWR.t1162 VGND 0.02183f
C12054 VPWR.n780 VGND 0.06746f
C12055 VPWR.n781 VGND 0.10257f
C12056 VPWR.n782 VGND 0.10257f
C12057 VPWR.t1020 VGND 0.02456f
C12058 VPWR.t1307 VGND 0.02183f
C12059 VPWR.n783 VGND 0.06746f
C12060 VPWR.t971 VGND 0.05786f
C12061 VPWR.t1306 VGND 0.06796f
C12062 VPWR.t1011 VGND 0.08814f
C12063 VPWR.t245 VGND 0.02456f
C12064 VPWR.t998 VGND 0.02183f
C12065 VPWR.n784 VGND 0.06746f
C12066 VPWR.n785 VGND 0.10257f
C12067 VPWR.n786 VGND 0.10257f
C12068 VPWR.t1012 VGND 0.02456f
C12069 VPWR.t1252 VGND 0.02183f
C12070 VPWR.n787 VGND 0.06746f
C12071 VPWR.t969 VGND 0.05786f
C12072 VPWR.t1251 VGND 0.06796f
C12073 VPWR.t23 VGND 0.02456f
C12074 VPWR.t1530 VGND 0.02183f
C12075 VPWR.n788 VGND 0.06746f
C12076 VPWR.t1230 VGND 0.02456f
C12077 VPWR.t1635 VGND 0.02183f
C12078 VPWR.n789 VGND 0.06746f
C12079 VPWR.t573 VGND 0.10698f
C12080 VPWR.t396 VGND 0.05786f
C12081 VPWR.t289 VGND 0.06796f
C12082 VPWR.t574 VGND 0.02456f
C12083 VPWR.t290 VGND 0.02183f
C12084 VPWR.n790 VGND 0.06746f
C12085 VPWR.n791 VGND 0.01325f
C12086 VPWR.n793 VGND 0.07978f
C12087 VPWR.t733 VGND 0.08814f
C12088 VPWR.t391 VGND 0.05786f
C12089 VPWR.t512 VGND 0.06796f
C12090 VPWR.t734 VGND 0.02456f
C12091 VPWR.t513 VGND 0.02183f
C12092 VPWR.n794 VGND 0.06746f
C12093 VPWR.n795 VGND 0.01325f
C12094 VPWR.n797 VGND 0.07978f
C12095 VPWR.t1186 VGND 0.08814f
C12096 VPWR.t1849 VGND 0.05786f
C12097 VPWR.t1085 VGND 0.06796f
C12098 VPWR.t1187 VGND 0.02456f
C12099 VPWR.t1086 VGND 0.02183f
C12100 VPWR.n798 VGND 0.06746f
C12101 VPWR.n799 VGND 0.01325f
C12102 VPWR.n801 VGND 0.07978f
C12103 VPWR.t1049 VGND 0.08814f
C12104 VPWR.t1848 VGND 0.05786f
C12105 VPWR.t411 VGND 0.06796f
C12106 VPWR.t1050 VGND 0.02456f
C12107 VPWR.t412 VGND 0.02183f
C12108 VPWR.n802 VGND 0.06746f
C12109 VPWR.n803 VGND 0.01325f
C12110 VPWR.n805 VGND 0.07978f
C12111 VPWR.t677 VGND 0.08814f
C12112 VPWR.t395 VGND 0.05786f
C12113 VPWR.t148 VGND 0.06796f
C12114 VPWR.t678 VGND 0.02456f
C12115 VPWR.t149 VGND 0.02183f
C12116 VPWR.n806 VGND 0.06746f
C12117 VPWR.n807 VGND 0.01325f
C12118 VPWR.n809 VGND 0.07978f
C12119 VPWR.t142 VGND 0.08814f
C12120 VPWR.t1854 VGND 0.05786f
C12121 VPWR.t56 VGND 0.06796f
C12122 VPWR.t143 VGND 0.02456f
C12123 VPWR.t57 VGND 0.02183f
C12124 VPWR.n810 VGND 0.06746f
C12125 VPWR.n811 VGND 0.01325f
C12126 VPWR.n813 VGND 0.07978f
C12127 VPWR.t50 VGND 0.08814f
C12128 VPWR.t1853 VGND 0.05786f
C12129 VPWR.t718 VGND 0.06796f
C12130 VPWR.t51 VGND 0.02456f
C12131 VPWR.t719 VGND 0.02183f
C12132 VPWR.n814 VGND 0.06746f
C12133 VPWR.n815 VGND 0.01325f
C12134 VPWR.n817 VGND 0.07978f
C12135 VPWR.t712 VGND 0.08814f
C12136 VPWR.t394 VGND 0.05786f
C12137 VPWR.t230 VGND 0.06796f
C12138 VPWR.t713 VGND 0.02456f
C12139 VPWR.t231 VGND 0.02183f
C12140 VPWR.n818 VGND 0.06746f
C12141 VPWR.n819 VGND 0.01325f
C12142 VPWR.n821 VGND 0.07978f
C12143 VPWR.t610 VGND 0.08814f
C12144 VPWR.t393 VGND 0.05786f
C12145 VPWR.t522 VGND 0.06796f
C12146 VPWR.t611 VGND 0.02456f
C12147 VPWR.t523 VGND 0.02183f
C12148 VPWR.n822 VGND 0.06746f
C12149 VPWR.n823 VGND 0.01325f
C12150 VPWR.n825 VGND 0.07978f
C12151 VPWR.t44 VGND 0.08814f
C12152 VPWR.t1855 VGND 0.05786f
C12153 VPWR.t328 VGND 0.06796f
C12154 VPWR.t45 VGND 0.02456f
C12155 VPWR.t329 VGND 0.02183f
C12156 VPWR.n826 VGND 0.06746f
C12157 VPWR.n827 VGND 0.01325f
C12158 VPWR.n829 VGND 0.07978f
C12159 VPWR.t2 VGND 0.08814f
C12160 VPWR.t1847 VGND 0.05786f
C12161 VPWR.t550 VGND 0.06796f
C12162 VPWR.t3 VGND 0.02456f
C12163 VPWR.t551 VGND 0.02183f
C12164 VPWR.n830 VGND 0.06746f
C12165 VPWR.n831 VGND 0.01325f
C12166 VPWR.n833 VGND 0.07978f
C12167 VPWR.t778 VGND 0.08814f
C12168 VPWR.t321 VGND 0.05786f
C12169 VPWR.t1861 VGND 0.06796f
C12170 VPWR.t779 VGND 0.02456f
C12171 VPWR.t1862 VGND 0.02183f
C12172 VPWR.n834 VGND 0.06746f
C12173 VPWR.n835 VGND 0.01325f
C12174 VPWR.n837 VGND 0.07978f
C12175 VPWR.t1871 VGND 0.08814f
C12176 VPWR.t1852 VGND 0.05786f
C12177 VPWR.t248 VGND 0.06796f
C12178 VPWR.t1872 VGND 0.02456f
C12179 VPWR.t249 VGND 0.02183f
C12180 VPWR.n838 VGND 0.06746f
C12181 VPWR.n839 VGND 0.01325f
C12182 VPWR.n841 VGND 0.07978f
C12183 VPWR.t976 VGND 0.08814f
C12184 VPWR.t1851 VGND 0.05786f
C12185 VPWR.t638 VGND 0.06796f
C12186 VPWR.t977 VGND 0.02456f
C12187 VPWR.t639 VGND 0.02183f
C12188 VPWR.n842 VGND 0.06746f
C12189 VPWR.n843 VGND 0.01325f
C12190 VPWR.n845 VGND 0.07978f
C12191 VPWR.t40 VGND 0.08814f
C12192 VPWR.t1850 VGND 0.05786f
C12193 VPWR.t26 VGND 0.06796f
C12194 VPWR.t41 VGND 0.02456f
C12195 VPWR.t27 VGND 0.02183f
C12196 VPWR.n846 VGND 0.06746f
C12197 VPWR.n847 VGND 0.01325f
C12198 VPWR.n849 VGND 0.07978f
C12199 VPWR.t1229 VGND 0.08814f
C12200 VPWR.t392 VGND 0.05786f
C12201 VPWR.t1634 VGND 0.09829f
C12202 VPWR.n850 VGND 0.05616f
C12203 VPWR.n851 VGND 0.01325f
C12204 VPWR.n852 VGND 0.10257f
C12205 VPWR.n853 VGND 0.7488f
C12206 VPWR.n854 VGND 0.10257f
C12207 VPWR.t1244 VGND 0.02456f
C12208 VPWR.t1455 VGND 0.02183f
C12209 VPWR.n855 VGND 0.06746f
C12210 VPWR.t829 VGND 0.06796f
C12211 VPWR.t1002 VGND 0.02456f
C12212 VPWR.t830 VGND 0.02183f
C12213 VPWR.n856 VGND 0.06746f
C12214 VPWR.n857 VGND 0.10257f
C12215 VPWR.n858 VGND 0.10257f
C12216 VPWR.t257 VGND 0.02456f
C12217 VPWR.t1198 VGND 0.02183f
C12218 VPWR.n859 VGND 0.06746f
C12219 VPWR.t397 VGND 0.06796f
C12220 VPWR.t1806 VGND 0.02456f
C12221 VPWR.t398 VGND 0.02183f
C12222 VPWR.n860 VGND 0.06746f
C12223 VPWR.n861 VGND 0.10257f
C12224 VPWR.n862 VGND 0.10257f
C12225 VPWR.t1412 VGND 0.02456f
C12226 VPWR.t1812 VGND 0.02183f
C12227 VPWR.n863 VGND 0.06746f
C12228 VPWR.t1124 VGND 0.06796f
C12229 VPWR.t349 VGND 0.02456f
C12230 VPWR.t1125 VGND 0.02183f
C12231 VPWR.n864 VGND 0.06746f
C12232 VPWR.n865 VGND 0.10257f
C12233 VPWR.n866 VGND 0.10257f
C12234 VPWR.t797 VGND 0.02456f
C12235 VPWR.t382 VGND 0.02183f
C12236 VPWR.n867 VGND 0.06746f
C12237 VPWR.t802 VGND 0.06796f
C12238 VPWR.t225 VGND 0.02456f
C12239 VPWR.t803 VGND 0.02183f
C12240 VPWR.n868 VGND 0.06746f
C12241 VPWR.n869 VGND 0.10257f
C12242 VPWR.n870 VGND 0.10257f
C12243 VPWR.t1902 VGND 0.02456f
C12244 VPWR.t243 VGND 0.02183f
C12245 VPWR.n871 VGND 0.06746f
C12246 VPWR.t1907 VGND 0.06796f
C12247 VPWR.t1102 VGND 0.02456f
C12248 VPWR.t1908 VGND 0.02183f
C12249 VPWR.n872 VGND 0.06746f
C12250 VPWR.n873 VGND 0.10257f
C12251 VPWR.n874 VGND 0.10257f
C12252 VPWR.t1326 VGND 0.02456f
C12253 VPWR.t846 VGND 0.02183f
C12254 VPWR.n875 VGND 0.06746f
C12255 VPWR.t1180 VGND 0.06796f
C12256 VPWR.t686 VGND 0.02456f
C12257 VPWR.t1181 VGND 0.02183f
C12258 VPWR.n876 VGND 0.06746f
C12259 VPWR.n877 VGND 0.10257f
C12260 VPWR.n878 VGND 0.10257f
C12261 VPWR.t1080 VGND 0.02456f
C12262 VPWR.t756 VGND 0.02183f
C12263 VPWR.n879 VGND 0.06746f
C12264 VPWR.t1055 VGND 0.06796f
C12265 VPWR.t1154 VGND 0.02456f
C12266 VPWR.t1056 VGND 0.02183f
C12267 VPWR.n880 VGND 0.06746f
C12268 VPWR.n881 VGND 0.10257f
C12269 VPWR.n882 VGND 0.10257f
C12270 VPWR.t73 VGND 0.02456f
C12271 VPWR.t1160 VGND 0.02183f
C12272 VPWR.n883 VGND 0.06746f
C12273 VPWR.t589 VGND 0.10698f
C12274 VPWR.t538 VGND 0.05786f
C12275 VPWR.t835 VGND 0.06796f
C12276 VPWR.t590 VGND 0.02456f
C12277 VPWR.t836 VGND 0.02183f
C12278 VPWR.n884 VGND 0.06746f
C12279 VPWR.t576 VGND 0.02456f
C12280 VPWR.t288 VGND 0.02183f
C12281 VPWR.n885 VGND 0.06746f
C12282 VPWR.t575 VGND 0.10698f
C12283 VPWR.t217 VGND 0.05786f
C12284 VPWR.t287 VGND 0.06796f
C12285 VPWR.t1228 VGND 0.02456f
C12286 VPWR.t1642 VGND 0.02183f
C12287 VPWR.n886 VGND 0.06746f
C12288 VPWR.n887 VGND 0.01325f
C12289 VPWR.n888 VGND 0.05616f
C12290 VPWR.t1641 VGND 0.09829f
C12291 VPWR.t213 VGND 0.05786f
C12292 VPWR.t1227 VGND 0.08814f
C12293 VPWR.t39 VGND 0.02456f
C12294 VPWR.t25 VGND 0.02183f
C12295 VPWR.n889 VGND 0.06746f
C12296 VPWR.n890 VGND 0.01325f
C12297 VPWR.n892 VGND 0.07978f
C12298 VPWR.t24 VGND 0.06796f
C12299 VPWR.t955 VGND 0.05786f
C12300 VPWR.t38 VGND 0.08814f
C12301 VPWR.t973 VGND 0.02456f
C12302 VPWR.t637 VGND 0.02183f
C12303 VPWR.n893 VGND 0.06746f
C12304 VPWR.n894 VGND 0.01325f
C12305 VPWR.n896 VGND 0.07978f
C12306 VPWR.t636 VGND 0.06796f
C12307 VPWR.t956 VGND 0.05786f
C12308 VPWR.t972 VGND 0.08814f
C12309 VPWR.t1870 VGND 0.02456f
C12310 VPWR.t247 VGND 0.02183f
C12311 VPWR.n897 VGND 0.06746f
C12312 VPWR.n898 VGND 0.01325f
C12313 VPWR.n900 VGND 0.07978f
C12314 VPWR.t246 VGND 0.06796f
C12315 VPWR.t957 VGND 0.05786f
C12316 VPWR.t1869 VGND 0.08814f
C12317 VPWR.t777 VGND 0.02456f
C12318 VPWR.t1860 VGND 0.02183f
C12319 VPWR.n901 VGND 0.06746f
C12320 VPWR.n902 VGND 0.01325f
C12321 VPWR.n904 VGND 0.07978f
C12322 VPWR.t1859 VGND 0.06796f
C12323 VPWR.t1913 VGND 0.05786f
C12324 VPWR.t776 VGND 0.08814f
C12325 VPWR.t1 VGND 0.02456f
C12326 VPWR.t549 VGND 0.02183f
C12327 VPWR.n905 VGND 0.06746f
C12328 VPWR.n906 VGND 0.01325f
C12329 VPWR.n908 VGND 0.07978f
C12330 VPWR.t548 VGND 0.06796f
C12331 VPWR.t1914 VGND 0.05786f
C12332 VPWR.t0 VGND 0.08814f
C12333 VPWR.t43 VGND 0.02456f
C12334 VPWR.t327 VGND 0.02183f
C12335 VPWR.n909 VGND 0.06746f
C12336 VPWR.n910 VGND 0.01325f
C12337 VPWR.n912 VGND 0.07978f
C12338 VPWR.t326 VGND 0.06796f
C12339 VPWR.t960 VGND 0.05786f
C12340 VPWR.t42 VGND 0.08814f
C12341 VPWR.t607 VGND 0.02456f
C12342 VPWR.t521 VGND 0.02183f
C12343 VPWR.n913 VGND 0.06746f
C12344 VPWR.n914 VGND 0.01325f
C12345 VPWR.n916 VGND 0.07978f
C12346 VPWR.t520 VGND 0.06796f
C12347 VPWR.t214 VGND 0.05786f
C12348 VPWR.t606 VGND 0.08814f
C12349 VPWR.t711 VGND 0.02456f
C12350 VPWR.t229 VGND 0.02183f
C12351 VPWR.n917 VGND 0.06746f
C12352 VPWR.n918 VGND 0.01325f
C12353 VPWR.n920 VGND 0.07978f
C12354 VPWR.t228 VGND 0.06796f
C12355 VPWR.t215 VGND 0.05786f
C12356 VPWR.t710 VGND 0.08814f
C12357 VPWR.t49 VGND 0.02456f
C12358 VPWR.t717 VGND 0.02183f
C12359 VPWR.n921 VGND 0.06746f
C12360 VPWR.n922 VGND 0.01325f
C12361 VPWR.n924 VGND 0.07978f
C12362 VPWR.t716 VGND 0.06796f
C12363 VPWR.t958 VGND 0.05786f
C12364 VPWR.t48 VGND 0.08814f
C12365 VPWR.t929 VGND 0.02456f
C12366 VPWR.t55 VGND 0.02183f
C12367 VPWR.n925 VGND 0.06746f
C12368 VPWR.n926 VGND 0.01325f
C12369 VPWR.n928 VGND 0.07978f
C12370 VPWR.t54 VGND 0.06796f
C12371 VPWR.t959 VGND 0.05786f
C12372 VPWR.t928 VGND 0.08814f
C12373 VPWR.t676 VGND 0.02456f
C12374 VPWR.t147 VGND 0.02183f
C12375 VPWR.n929 VGND 0.06746f
C12376 VPWR.n930 VGND 0.01325f
C12377 VPWR.n932 VGND 0.07978f
C12378 VPWR.t146 VGND 0.06796f
C12379 VPWR.t216 VGND 0.05786f
C12380 VPWR.t675 VGND 0.08814f
C12381 VPWR.t1052 VGND 0.02456f
C12382 VPWR.t410 VGND 0.02183f
C12383 VPWR.n933 VGND 0.06746f
C12384 VPWR.n934 VGND 0.01325f
C12385 VPWR.n936 VGND 0.07978f
C12386 VPWR.t409 VGND 0.06796f
C12387 VPWR.t1915 VGND 0.05786f
C12388 VPWR.t1051 VGND 0.08814f
C12389 VPWR.t1185 VGND 0.02456f
C12390 VPWR.t1088 VGND 0.02183f
C12391 VPWR.n937 VGND 0.06746f
C12392 VPWR.n938 VGND 0.01325f
C12393 VPWR.n940 VGND 0.07978f
C12394 VPWR.t1087 VGND 0.06796f
C12395 VPWR.t954 VGND 0.05786f
C12396 VPWR.t1184 VGND 0.08814f
C12397 VPWR.t732 VGND 0.02456f
C12398 VPWR.t511 VGND 0.02183f
C12399 VPWR.n941 VGND 0.06746f
C12400 VPWR.n942 VGND 0.01325f
C12401 VPWR.n944 VGND 0.07978f
C12402 VPWR.t510 VGND 0.06796f
C12403 VPWR.t212 VGND 0.05786f
C12404 VPWR.t731 VGND 0.08814f
C12405 VPWR.n945 VGND 0.07978f
C12406 VPWR.n947 VGND 0.01325f
C12407 VPWR.n948 VGND 0.10257f
C12408 VPWR.n949 VGND 0.74411f
C12409 VPWR.n950 VGND 0.10257f
C12410 VPWR.t582 VGND 0.02456f
C12411 VPWR.t791 VGND 0.02183f
C12412 VPWR.n951 VGND 0.06746f
C12413 VPWR.t581 VGND 0.10698f
C12414 VPWR.t1133 VGND 0.05786f
C12415 VPWR.t790 VGND 0.06796f
C12416 VPWR.t1275 VGND 0.08814f
C12417 VPWR.t1129 VGND 0.02456f
C12418 VPWR.t1119 VGND 0.02183f
C12419 VPWR.n952 VGND 0.06746f
C12420 VPWR.n953 VGND 0.10257f
C12421 VPWR.n954 VGND 0.10257f
C12422 VPWR.t1276 VGND 0.02456f
C12423 VPWR.t1040 VGND 0.02183f
C12424 VPWR.n955 VGND 0.06746f
C12425 VPWR.t1137 VGND 0.05786f
C12426 VPWR.t1039 VGND 0.06796f
C12427 VPWR.t10 VGND 0.08814f
C12428 VPWR.t1064 VGND 0.02456f
C12429 VPWR.t680 VGND 0.02183f
C12430 VPWR.n956 VGND 0.06746f
C12431 VPWR.n957 VGND 0.10257f
C12432 VPWR.n958 VGND 0.10257f
C12433 VPWR.t11 VGND 0.02456f
C12434 VPWR.t908 VGND 0.02183f
C12435 VPWR.n959 VGND 0.06746f
C12436 VPWR.t1132 VGND 0.05786f
C12437 VPWR.t907 VGND 0.06796f
C12438 VPWR.t1819 VGND 0.08814f
C12439 VPWR.t900 VGND 0.02456f
C12440 VPWR.t1828 VGND 0.02183f
C12441 VPWR.n960 VGND 0.06746f
C12442 VPWR.n961 VGND 0.10257f
C12443 VPWR.n962 VGND 0.10257f
C12444 VPWR.t1820 VGND 0.02456f
C12445 VPWR.t1389 VGND 0.02183f
C12446 VPWR.n963 VGND 0.06746f
C12447 VPWR.t173 VGND 0.05786f
C12448 VPWR.t1388 VGND 0.06796f
C12449 VPWR.t234 VGND 0.08814f
C12450 VPWR.t1381 VGND 0.02456f
C12451 VPWR.t933 VGND 0.02183f
C12452 VPWR.n964 VGND 0.06746f
C12453 VPWR.n965 VGND 0.10257f
C12454 VPWR.n966 VGND 0.10257f
C12455 VPWR.t235 VGND 0.02456f
C12456 VPWR.t1286 VGND 0.02183f
C12457 VPWR.n967 VGND 0.06746f
C12458 VPWR.t1357 VGND 0.05786f
C12459 VPWR.t1285 VGND 0.06796f
C12460 VPWR.t389 VGND 0.08814f
C12461 VPWR.t1278 VGND 0.02456f
C12462 VPWR.t363 VGND 0.02183f
C12463 VPWR.n968 VGND 0.06746f
C12464 VPWR.n969 VGND 0.10257f
C12465 VPWR.n970 VGND 0.10257f
C12466 VPWR.t390 VGND 0.02456f
C12467 VPWR.t1840 VGND 0.02183f
C12468 VPWR.n971 VGND 0.06746f
C12469 VPWR.t1135 VGND 0.05786f
C12470 VPWR.t1839 VGND 0.06796f
C12471 VPWR.t628 VGND 0.08814f
C12472 VPWR.t483 VGND 0.02456f
C12473 VPWR.t1028 VGND 0.02183f
C12474 VPWR.n972 VGND 0.06746f
C12475 VPWR.n973 VGND 0.10257f
C12476 VPWR.n974 VGND 0.10257f
C12477 VPWR.t629 VGND 0.02456f
C12478 VPWR.t182 VGND 0.02183f
C12479 VPWR.n975 VGND 0.06746f
C12480 VPWR.t172 VGND 0.05786f
C12481 VPWR.t181 VGND 0.06796f
C12482 VPWR.t599 VGND 0.08814f
C12483 VPWR.t1311 VGND 0.02456f
C12484 VPWR.t994 VGND 0.02183f
C12485 VPWR.n976 VGND 0.06746f
C12486 VPWR.n977 VGND 0.10257f
C12487 VPWR.n978 VGND 0.10257f
C12488 VPWR.t600 VGND 0.02456f
C12489 VPWR.t1232 VGND 0.02183f
C12490 VPWR.n979 VGND 0.06746f
C12491 VPWR.t170 VGND 0.05786f
C12492 VPWR.t1231 VGND 0.06796f
C12493 VPWR.t822 VGND 0.02456f
C12494 VPWR.t1750 VGND 0.02183f
C12495 VPWR.n980 VGND 0.06746f
C12496 VPWR.t1240 VGND 0.02456f
C12497 VPWR.t1602 VGND 0.02183f
C12498 VPWR.n981 VGND 0.06746f
C12499 VPWR.t566 VGND 0.10698f
C12500 VPWR.t1292 VGND 0.05786f
C12501 VPWR.t500 VGND 0.06796f
C12502 VPWR.t567 VGND 0.02456f
C12503 VPWR.t501 VGND 0.02183f
C12504 VPWR.n982 VGND 0.06746f
C12505 VPWR.n983 VGND 0.01325f
C12506 VPWR.n985 VGND 0.07978f
C12507 VPWR.t285 VGND 0.08814f
C12508 VPWR.t1289 VGND 0.05786f
C12509 VPWR.t518 VGND 0.06796f
C12510 VPWR.t286 VGND 0.02456f
C12511 VPWR.t519 VGND 0.02183f
C12512 VPWR.n986 VGND 0.06746f
C12513 VPWR.n987 VGND 0.01325f
C12514 VPWR.n989 VGND 0.07978f
C12515 VPWR.t514 VGND 0.08814f
C12516 VPWR.t96 VGND 0.05786f
C12517 VPWR.t1075 VGND 0.06796f
C12518 VPWR.t515 VGND 0.02456f
C12519 VPWR.t1076 VGND 0.02183f
C12520 VPWR.n990 VGND 0.06746f
C12521 VPWR.n991 VGND 0.01325f
C12522 VPWR.n993 VGND 0.07978f
C12523 VPWR.t1041 VGND 0.08814f
C12524 VPWR.t95 VGND 0.05786f
C12525 VPWR.t415 VGND 0.06796f
C12526 VPWR.t1042 VGND 0.02456f
C12527 VPWR.t416 VGND 0.02183f
C12528 VPWR.n994 VGND 0.06746f
C12529 VPWR.n995 VGND 0.01325f
C12530 VPWR.n997 VGND 0.07978f
C12531 VPWR.t1398 VGND 0.08814f
C12532 VPWR.t492 VGND 0.05786f
C12533 VPWR.t1259 VGND 0.06796f
C12534 VPWR.t1399 VGND 0.02456f
C12535 VPWR.t1260 VGND 0.02183f
C12536 VPWR.n998 VGND 0.06746f
C12537 VPWR.n999 VGND 0.01325f
C12538 VPWR.n1001 VGND 0.07978f
C12539 VPWR.t150 VGND 0.08814f
C12540 VPWR.t1298 VGND 0.05786f
C12541 VPWR.t62 VGND 0.06796f
C12542 VPWR.t151 VGND 0.02456f
C12543 VPWR.t63 VGND 0.02183f
C12544 VPWR.n1002 VGND 0.06746f
C12545 VPWR.n1003 VGND 0.01325f
C12546 VPWR.n1005 VGND 0.07978f
C12547 VPWR.t58 VGND 0.08814f
C12548 VPWR.t1297 VGND 0.05786f
C12549 VPWR.t724 VGND 0.06796f
C12550 VPWR.t59 VGND 0.02456f
C12551 VPWR.t725 VGND 0.02183f
C12552 VPWR.n1006 VGND 0.06746f
C12553 VPWR.n1007 VGND 0.01325f
C12554 VPWR.n1009 VGND 0.07978f
C12555 VPWR.t720 VGND 0.08814f
C12556 VPWR.t491 VGND 0.05786f
C12557 VPWR.t220 VGND 0.06796f
C12558 VPWR.t721 VGND 0.02456f
C12559 VPWR.t221 VGND 0.02183f
C12560 VPWR.n1010 VGND 0.06746f
C12561 VPWR.n1011 VGND 0.01325f
C12562 VPWR.n1013 VGND 0.07978f
C12563 VPWR.t934 VGND 0.08814f
C12564 VPWR.t1291 VGND 0.05786f
C12565 VPWR.t528 VGND 0.06796f
C12566 VPWR.t935 VGND 0.02456f
C12567 VPWR.t529 VGND 0.02183f
C12568 VPWR.n1014 VGND 0.06746f
C12569 VPWR.n1015 VGND 0.01325f
C12570 VPWR.n1017 VGND 0.07978f
C12571 VPWR.t524 VGND 0.08814f
C12572 VPWR.t1299 VGND 0.05786f
C12573 VPWR.t336 VGND 0.06796f
C12574 VPWR.t525 VGND 0.02456f
C12575 VPWR.t337 VGND 0.02183f
C12576 VPWR.n1018 VGND 0.06746f
C12577 VPWR.n1019 VGND 0.01325f
C12578 VPWR.n1021 VGND 0.07978f
C12579 VPWR.t324 VGND 0.08814f
C12580 VPWR.t94 VGND 0.05786f
C12581 VPWR.t556 VGND 0.06796f
C12582 VPWR.t325 VGND 0.02456f
C12583 VPWR.t557 VGND 0.02183f
C12584 VPWR.n1022 VGND 0.06746f
C12585 VPWR.n1023 VGND 0.01325f
C12586 VPWR.n1025 VGND 0.07978f
C12587 VPWR.t552 VGND 0.08814f
C12588 VPWR.t1293 VGND 0.05786f
C12589 VPWR.t1015 VGND 0.06796f
C12590 VPWR.t553 VGND 0.02456f
C12591 VPWR.t1016 VGND 0.02183f
C12592 VPWR.n1026 VGND 0.06746f
C12593 VPWR.n1027 VGND 0.01325f
C12594 VPWR.n1029 VGND 0.07978f
C12595 VPWR.t1875 VGND 0.08814f
C12596 VPWR.t1296 VGND 0.05786f
C12597 VPWR.t252 VGND 0.06796f
C12598 VPWR.t1876 VGND 0.02456f
C12599 VPWR.t253 VGND 0.02183f
C12600 VPWR.n1030 VGND 0.06746f
C12601 VPWR.n1031 VGND 0.01325f
C12602 VPWR.n1033 VGND 0.07978f
C12603 VPWR.t183 VGND 0.08814f
C12604 VPWR.t1295 VGND 0.05786f
C12605 VPWR.t1007 VGND 0.06796f
C12606 VPWR.t184 VGND 0.02456f
C12607 VPWR.t1008 VGND 0.02183f
C12608 VPWR.n1034 VGND 0.06746f
C12609 VPWR.n1035 VGND 0.01325f
C12610 VPWR.n1037 VGND 0.07978f
C12611 VPWR.t634 VGND 0.08814f
C12612 VPWR.t97 VGND 0.05786f
C12613 VPWR.t14 VGND 0.06796f
C12614 VPWR.t635 VGND 0.02456f
C12615 VPWR.t15 VGND 0.02183f
C12616 VPWR.n1038 VGND 0.06746f
C12617 VPWR.n1039 VGND 0.01325f
C12618 VPWR.n1041 VGND 0.07978f
C12619 VPWR.t1239 VGND 0.08814f
C12620 VPWR.t1290 VGND 0.05786f
C12621 VPWR.t1601 VGND 0.09829f
C12622 VPWR.n1042 VGND 0.05616f
C12623 VPWR.n1043 VGND 0.01325f
C12624 VPWR.n1044 VGND 0.10257f
C12625 VPWR.n1045 VGND 4.31033f
C12626 VPWR.n1046 VGND 0.04841f
C12627 VPWR.n1047 VGND -0.01375f
C12628 VPWR.n1048 VGND 0.02243f
C12629 VPWR.t1605 VGND 0.01975f
C12630 VPWR.n1050 VGND 0.04219f
C12631 VPWR.t1719 VGND 0.02183f
C12632 VPWR.n1051 VGND 0.03459f
C12633 VPWR.t1241 VGND 0.06796f
C12634 VPWR.n1052 VGND 0.02243f
C12635 VPWR.t1497 VGND 0.01975f
C12636 VPWR.n1054 VGND 0.04219f
C12637 VPWR.t1242 VGND 0.02183f
C12638 VPWR.n1055 VGND 0.03459f
C12639 VPWR.n1056 VGND -0.01375f
C12640 VPWR.n1057 VGND 0.04841f
C12641 VPWR.n1058 VGND 0.02041f
C12642 VPWR.n1059 VGND 0.01398f
C12643 VPWR.n1060 VGND 0.04603f
C12644 VPWR.n1061 VGND 0.07184f
C12645 VPWR.n1062 VGND 0.04011f
C12646 VPWR.n1063 VGND 0.04841f
C12647 VPWR.n1064 VGND -0.01375f
C12648 VPWR.n1065 VGND 0.02243f
C12649 VPWR.t1583 VGND 0.01975f
C12650 VPWR.n1067 VGND 0.04219f
C12651 VPWR.t1887 VGND 0.02183f
C12652 VPWR.n1068 VGND 0.03459f
C12653 VPWR.t1886 VGND 0.06796f
C12654 VPWR.t1459 VGND 0.08814f
C12655 VPWR.n1069 VGND 0.02243f
C12656 VPWR.t1624 VGND 0.01975f
C12657 VPWR.n1071 VGND 0.04219f
C12658 VPWR.t190 VGND 0.02183f
C12659 VPWR.n1072 VGND 0.03459f
C12660 VPWR.n1074 VGND 0.1428f
C12661 VPWR.n1075 VGND 0.06156f
C12662 VPWR.n1076 VGND 0.02534f
C12663 VPWR.t1680 VGND 0.02456f
C12664 VPWR.t1672 VGND 0.02183f
C12665 VPWR.n1077 VGND 0.06746f
C12666 VPWR.t1671 VGND 0.06796f
C12667 VPWR.t1424 VGND 0.08814f
C12668 VPWR.t1711 VGND 0.02456f
C12669 VPWR.t1703 VGND 0.02183f
C12670 VPWR.n1078 VGND 0.06746f
C12671 VPWR.t1425 VGND 0.02456f
C12672 VPWR.t1548 VGND 0.02183f
C12673 VPWR.n1080 VGND 0.06746f
C12674 VPWR.t1420 VGND 0.05786f
C12675 VPWR.t1547 VGND 0.09829f
C12676 VPWR.n1081 VGND 0.05613f
C12677 VPWR.n1082 VGND 0.01252f
C12678 VPWR.n1083 VGND 0.02206f
C12679 VPWR.n1084 VGND 0.02421f
C12680 VPWR.n1086 VGND 0.01343f
C12681 VPWR.n1087 VGND 0.12963f
C12682 VPWR.n1088 VGND 0.02206f
C12683 VPWR.n1089 VGND 0.02421f
C12684 VPWR.n1090 VGND 0.01264f
C12685 VPWR.n1093 VGND 0.01264f
C12686 VPWR.n1095 VGND 0.0204f
C12687 VPWR.n1096 VGND 0.02077f
C12688 VPWR.n1097 VGND 0.01343f
C12689 VPWR.n1098 VGND 0.12963f
C12690 VPWR.n1099 VGND 0.02206f
C12691 VPWR.n1100 VGND 0.02421f
C12692 VPWR.n1101 VGND 0.01264f
C12693 VPWR.n1103 VGND 0.01264f
C12694 VPWR.n1105 VGND 0.0204f
C12695 VPWR.n1106 VGND 0.02077f
C12696 VPWR.n1107 VGND 0.01343f
C12697 VPWR.n1108 VGND 0.12963f
C12698 VPWR.n1109 VGND 0.02206f
C12699 VPWR.n1110 VGND 0.02421f
C12700 VPWR.n1111 VGND 0.01264f
C12701 VPWR.n1113 VGND 0.01264f
C12702 VPWR.n1115 VGND 0.0204f
C12703 VPWR.n1116 VGND 0.02077f
C12704 VPWR.n1117 VGND 0.01343f
C12705 VPWR.n1118 VGND 0.12963f
C12706 VPWR.n1119 VGND 0.02206f
C12707 VPWR.n1120 VGND 0.02421f
C12708 VPWR.n1121 VGND 0.01264f
C12709 VPWR.n1123 VGND 0.01264f
C12710 VPWR.n1125 VGND 0.0204f
C12711 VPWR.n1126 VGND 0.02077f
C12712 VPWR.n1127 VGND 0.01343f
C12713 VPWR.n1128 VGND 0.01957f
C12714 VPWR.n1129 VGND 0.02206f
C12715 VPWR.n1130 VGND 0.02421f
C12716 VPWR.n1131 VGND 0.01343f
C12717 VPWR.n1133 VGND 0.02297f
C12718 VPWR.n1134 VGND 0.01452f
C12719 VPWR.n1135 VGND 0.0204f
C12720 VPWR.n1136 VGND 0.02077f
C12721 VPWR.n1137 VGND 0.01309f
C12722 VPWR.n1138 VGND 0.02206f
C12723 VPWR.n1139 VGND 0.02421f
C12724 VPWR.t1729 VGND 0.02456f
C12725 VPWR.t1444 VGND 0.02183f
C12726 VPWR.n1141 VGND 0.06746f
C12727 VPWR.t1728 VGND 0.10698f
C12728 VPWR.t1721 VGND 0.05786f
C12729 VPWR.t1443 VGND 0.06796f
C12730 VPWR.t1598 VGND 0.08814f
C12731 VPWR.t1494 VGND 0.02456f
C12732 VPWR.t1580 VGND 0.02183f
C12733 VPWR.n1142 VGND 0.06746f
C12734 VPWR.n1144 VGND 0.02297f
C12735 VPWR.n1145 VGND 0.02723f
C12736 VPWR.n1146 VGND 0.02534f
C12737 VPWR.n1147 VGND 0.10257f
C12738 VPWR.n1149 VGND 0.01325f
C12739 VPWR.n1150 VGND 0.04841f
C12740 VPWR.n1151 VGND 0.04011f
C12741 VPWR.n1152 VGND 0.02041f
C12742 VPWR.n1153 VGND 0.01398f
C12743 VPWR.n1154 VGND 0.04603f
C12744 VPWR.n1155 VGND 0.07184f
C12745 VPWR.n1156 VGND 0.04841f
C12746 VPWR.n1157 VGND 0.04841f
C12747 VPWR.n1158 VGND 0.04841f
C12748 VPWR.n1159 VGND 0.04841f
C12749 VPWR.n1160 VGND 0.04841f
C12750 VPWR.n1161 VGND 0.04841f
C12751 VPWR.n1162 VGND 0.04011f
C12752 VPWR.n1164 VGND -0.01375f
C12753 VPWR.n1165 VGND 0.02243f
C12754 VPWR.t1716 VGND 0.01975f
C12755 VPWR.n1167 VGND 0.04219f
C12756 VPWR.t369 VGND 0.02183f
C12757 VPWR.n1168 VGND 0.03459f
C12758 VPWR.t368 VGND 0.06796f
C12759 VPWR.t1452 VGND 0.05786f
C12760 VPWR.t1582 VGND 0.08814f
C12761 VPWR.n1169 VGND 0.02243f
C12762 VPWR.t1450 VGND 0.01975f
C12763 VPWR.n1171 VGND 0.04219f
C12764 VPWR.t1846 VGND 0.02183f
C12765 VPWR.n1172 VGND 0.03459f
C12766 VPWR.n1175 VGND 0.02243f
C12767 VPWR.t1694 VGND 0.01975f
C12768 VPWR.n1177 VGND 0.04219f
C12769 VPWR.t298 VGND 0.02183f
C12770 VPWR.n1178 VGND 0.03459f
C12771 VPWR.t948 VGND 0.06796f
C12772 VPWR.n1179 VGND 0.02243f
C12773 VPWR.t1553 VGND 0.01975f
C12774 VPWR.n1181 VGND 0.04219f
C12775 VPWR.t949 VGND 0.02183f
C12776 VPWR.n1182 VGND 0.03459f
C12777 VPWR.n1185 VGND 0.02243f
C12778 VPWR.t1431 VGND 0.01975f
C12779 VPWR.n1187 VGND 0.04219f
C12780 VPWR.t1395 VGND 0.02183f
C12781 VPWR.n1188 VGND 0.03459f
C12782 VPWR.t1803 VGND 0.06796f
C12783 VPWR.n1189 VGND 0.02243f
C12784 VPWR.t1683 VGND 0.01975f
C12785 VPWR.n1191 VGND 0.04219f
C12786 VPWR.t1804 VGND 0.02183f
C12787 VPWR.n1192 VGND 0.03459f
C12788 VPWR.n1195 VGND 0.02297f
C12789 VPWR.n1196 VGND 0.02723f
C12790 VPWR.n1197 VGND 0.02534f
C12791 VPWR.t1479 VGND 0.02456f
C12792 VPWR.t1474 VGND 0.02183f
C12793 VPWR.n1198 VGND 0.06746f
C12794 VPWR.t1585 VGND 0.05786f
C12795 VPWR.t1592 VGND 0.06796f
C12796 VPWR.t1599 VGND 0.02456f
C12797 VPWR.t1593 VGND 0.02183f
C12798 VPWR.n1199 VGND 0.06746f
C12799 VPWR.n1201 VGND 0.07978f
C12800 VPWR.t1760 VGND 0.08814f
C12801 VPWR.t1626 VGND 0.05786f
C12802 VPWR.t1755 VGND 0.06796f
C12803 VPWR.t1761 VGND 0.02456f
C12804 VPWR.t1756 VGND 0.02183f
C12805 VPWR.n1202 VGND 0.06746f
C12806 VPWR.n1204 VGND 0.07978f
C12807 VPWR.t1478 VGND 0.08814f
C12808 VPWR.t1737 VGND 0.05786f
C12809 VPWR.t1473 VGND 0.06796f
C12810 VPWR.t1550 VGND 0.05786f
C12811 VPWR.t1679 VGND 0.08814f
C12812 VPWR.t1439 VGND 0.02456f
C12813 VPWR.t1540 VGND 0.02183f
C12814 VPWR.n1205 VGND 0.06746f
C12815 VPWR.n1207 VGND 0.07978f
C12816 VPWR.t1539 VGND 0.06796f
C12817 VPWR.t1524 VGND 0.05786f
C12818 VPWR.t1438 VGND 0.08814f
C12819 VPWR.t1418 VGND 0.02456f
C12820 VPWR.t1796 VGND 0.02183f
C12821 VPWR.n1208 VGND 0.06746f
C12822 VPWR.n1210 VGND 0.07978f
C12823 VPWR.t1795 VGND 0.06796f
C12824 VPWR.t1677 VGND 0.05786f
C12825 VPWR.t1417 VGND 0.08814f
C12826 VPWR.t1667 VGND 0.02456f
C12827 VPWR.t1777 VGND 0.02183f
C12828 VPWR.n1211 VGND 0.06746f
C12829 VPWR.n1213 VGND 0.02297f
C12830 VPWR.n1214 VGND 0.02723f
C12831 VPWR.n1215 VGND 0.02534f
C12832 VPWR.n1216 VGND 0.01264f
C12833 VPWR.n1218 VGND 0.07978f
C12834 VPWR.t1776 VGND 0.06796f
C12835 VPWR.t1652 VGND 0.05786f
C12836 VPWR.t1666 VGND 0.08814f
C12837 VPWR.t1545 VGND 0.02456f
C12838 VPWR.t1618 VGND 0.02183f
C12839 VPWR.n1219 VGND 0.06746f
C12840 VPWR.n1221 VGND 0.07978f
C12841 VPWR.t1617 VGND 0.06796f
C12842 VPWR.t1499 VGND 0.05786f
C12843 VPWR.t1544 VGND 0.08814f
C12844 VPWR.t1519 VGND 0.02456f
C12845 VPWR.t1514 VGND 0.02183f
C12846 VPWR.n1222 VGND 0.06746f
C12847 VPWR.n1224 VGND 0.07978f
C12848 VPWR.t1513 VGND 0.06796f
C12849 VPWR.t1782 VGND 0.05786f
C12850 VPWR.t1518 VGND 0.08814f
C12851 VPWR.t1753 VGND 0.02456f
C12852 VPWR.t1769 VGND 0.02183f
C12853 VPWR.n1225 VGND 0.06746f
C12854 VPWR.n1227 VGND 0.02297f
C12855 VPWR.n1228 VGND 0.02723f
C12856 VPWR.n1229 VGND 0.02534f
C12857 VPWR.n1230 VGND 0.01264f
C12858 VPWR.n1232 VGND 0.07978f
C12859 VPWR.t1768 VGND 0.06796f
C12860 VPWR.t1742 VGND 0.05786f
C12861 VPWR.t1752 VGND 0.08814f
C12862 VPWR.t1650 VGND 0.02456f
C12863 VPWR.t1732 VGND 0.02183f
C12864 VPWR.n1233 VGND 0.06746f
C12865 VPWR.n1235 VGND 0.07978f
C12866 VPWR.t1731 VGND 0.06796f
C12867 VPWR.t1516 VGND 0.05786f
C12868 VPWR.t1649 VGND 0.08814f
C12869 VPWR.t1491 VGND 0.02456f
C12870 VPWR.t1621 VGND 0.02183f
C12871 VPWR.n1236 VGND 0.06746f
C12872 VPWR.n1238 VGND 0.07978f
C12873 VPWR.t1620 VGND 0.06796f
C12874 VPWR.t1501 VGND 0.05786f
C12875 VPWR.t1490 VGND 0.08814f
C12876 VPWR.n1239 VGND 0.07978f
C12877 VPWR.n1241 VGND 0.01264f
C12878 VPWR.n1243 VGND 0.02243f
C12879 VPWR.t1658 VGND 0.01975f
C12880 VPWR.n1245 VGND 0.04219f
C12881 VPWR.t1148 VGND 0.02183f
C12882 VPWR.n1246 VGND 0.03459f
C12883 VPWR.t1521 VGND 0.10698f
C12884 VPWR.t1506 VGND 0.05786f
C12885 VPWR.t663 VGND 0.06796f
C12886 VPWR.n1247 VGND 0.02243f
C12887 VPWR.t1522 VGND 0.01975f
C12888 VPWR.n1249 VGND 0.04219f
C12889 VPWR.t664 VGND 0.02183f
C12890 VPWR.n1250 VGND 0.03459f
C12891 VPWR.n1251 VGND -0.01375f
C12892 VPWR.n1252 VGND 0.03455f
C12893 VPWR.t28 VGND 0.71923f
C12894 VPWR.n1253 VGND 0.39227f
C12895 VPWR.t100 VGND 0.71923f
C12896 VPWR.n1254 VGND 0.30507f
C12897 VPWR.n1255 VGND 0.21437f
C12898 VPWR.t729 VGND 0.04214f
C12899 VPWR.t32 VGND 0.01056f
C12900 VPWR.t35 VGND 0.01056f
C12901 VPWR.n1257 VGND 0.02319f
C12902 VPWR.t36 VGND 0.01056f
C12903 VPWR.t29 VGND 0.01056f
C12904 VPWR.n1258 VGND 0.02315f
C12905 VPWR.t106 VGND 0.01056f
C12906 VPWR.t105 VGND 0.01056f
C12907 VPWR.n1259 VGND 0.02315f
C12908 VPWR.n1260 VGND 0.07682f
C12909 VPWR.n1261 VGND 0.13403f
C12910 VPWR.n1262 VGND 0.04244f
C12911 VPWR.n1263 VGND 0.03117f
C12912 VPWR.t101 VGND 0.01056f
C12913 VPWR.t107 VGND 0.01056f
C12914 VPWR.n1264 VGND 0.02319f
C12915 VPWR.n1265 VGND 0.09511f
C12916 VPWR.n1267 VGND 0.01202f
C12917 VPWR.n1268 VGND 0.01408f
C12918 VPWR.n1269 VGND 0.02065f
C12919 VPWR.t728 VGND 0.04214f
C12920 VPWR.n1270 VGND 0.11101f
C12921 VPWR.t1405 VGND 0.04212f
C12922 VPWR.t1882 VGND 0.04212f
C12923 VPWR.n1272 VGND 0.09912f
C12924 VPWR.n1273 VGND 0.24742f
C12925 VPWR.n1274 VGND 1.20965f
C12926 VPWR.n1275 VGND 0.03455f
C12927 VPWR.t158 VGND 0.71923f
C12928 VPWR.n1276 VGND 0.39227f
C12929 VPWR.t207 VGND 0.71923f
C12930 VPWR.n1277 VGND 0.30507f
C12931 VPWR.n1278 VGND 0.2163f
C12932 VPWR.t165 VGND 0.01056f
C12933 VPWR.t163 VGND 0.01056f
C12934 VPWR.n1280 VGND 0.02319f
C12935 VPWR.t162 VGND 0.01056f
C12936 VPWR.t159 VGND 0.01056f
C12937 VPWR.n1281 VGND 0.02315f
C12938 VPWR.t208 VGND 0.01056f
C12939 VPWR.t209 VGND 0.01056f
C12940 VPWR.n1282 VGND 0.02315f
C12941 VPWR.n1283 VGND 0.07682f
C12942 VPWR.n1284 VGND 0.13403f
C12943 VPWR.n1285 VGND 0.04244f
C12944 VPWR.n1286 VGND 0.03117f
C12945 VPWR.t1107 VGND 0.01056f
C12946 VPWR.t660 VGND 0.01056f
C12947 VPWR.n1287 VGND 0.02319f
C12948 VPWR.n1288 VGND 0.09511f
C12949 VPWR.n1290 VGND 0.01202f
C12950 VPWR.n1291 VGND 0.01408f
C12951 VPWR.n1292 VGND 0.02028f
C12952 VPWR.t730 VGND 0.04208f
C12953 VPWR.n1294 VGND 0.04498f
C12954 VPWR.t759 VGND 0.04217f
C12955 VPWR.n1296 VGND 0.06716f
C12956 VPWR.n1297 VGND 0.24742f
C12957 VPWR.n1298 VGND 1.20965f
C12958 VPWR.n1299 VGND 0.03455f
C12959 VPWR.t114 VGND 0.71923f
C12960 VPWR.n1300 VGND 0.39227f
C12961 VPWR.t316 VGND 0.71923f
C12962 VPWR.n1301 VGND 0.30507f
C12963 VPWR.n1302 VGND 0.2163f
C12964 VPWR.t119 VGND 0.01056f
C12965 VPWR.t117 VGND 0.01056f
C12966 VPWR.n1304 VGND 0.02319f
C12967 VPWR.t116 VGND 0.01056f
C12968 VPWR.t115 VGND 0.01056f
C12969 VPWR.n1305 VGND 0.02315f
C12970 VPWR.t762 VGND 0.01056f
C12971 VPWR.t769 VGND 0.01056f
C12972 VPWR.n1306 VGND 0.02315f
C12973 VPWR.n1307 VGND 0.07682f
C12974 VPWR.n1308 VGND 0.13403f
C12975 VPWR.n1309 VGND 0.04244f
C12976 VPWR.n1310 VGND 0.03117f
C12977 VPWR.t766 VGND 0.01056f
C12978 VPWR.t763 VGND 0.01056f
C12979 VPWR.n1311 VGND 0.02319f
C12980 VPWR.n1312 VGND 0.09511f
C12981 VPWR.n1314 VGND 0.01202f
C12982 VPWR.n1315 VGND 0.01408f
C12983 VPWR.n1316 VGND 0.02028f
C12984 VPWR.n1317 VGND 0.01031f
C12985 VPWR.t1406 VGND 0.04217f
C12986 VPWR.t1883 VGND 0.04217f
C12987 VPWR.n1319 VGND 0.12454f
C12988 VPWR.n1320 VGND 0.24742f
C12989 VPWR.n1321 VGND 1.20965f
C12990 VPWR.t469 VGND 0.0421f
C12991 VPWR.t918 VGND 0.04217f
C12992 VPWR.t471 VGND 0.04181f
C12993 VPWR.n1322 VGND 0.10841f
C12994 VPWR.t264 VGND 0.04133f
C12995 VPWR.n1323 VGND 0.04995f
C12996 VPWR.n1324 VGND 0.03455f
C12997 VPWR.t450 VGND 0.03979f
C12998 VPWR.n1325 VGND 0.03784f
C12999 VPWR.t1836 VGND 0.01056f
C13000 VPWR.t318 VGND 0.01056f
C13001 VPWR.n1326 VGND 0.02308f
C13002 VPWR.t1348 VGND 0.03697f
C13003 VPWR.n1327 VGND 0.05544f
C13004 VPWR.n1328 VGND 0.03455f
C13005 VPWR.t1371 VGND 0.04212f
C13006 VPWR.n1329 VGND 0.05303f
C13007 VPWR.n1330 VGND 0.02028f
C13008 VPWR.n1331 VGND 0.03455f
C13009 VPWR.t320 VGND 0.01056f
C13010 VPWR.t473 VGND 0.01056f
C13011 VPWR.n1333 VGND 0.02308f
C13012 VPWR.n1334 VGND 0.03382f
C13013 VPWR.n1336 VGND 0.02591f
C13014 VPWR.n1337 VGND 0.02591f
C13015 VPWR.n1338 VGND 0.03455f
C13016 VPWR.t1832 VGND 0.01056f
C13017 VPWR.t625 VGND 0.01056f
C13018 VPWR.n1340 VGND 0.02308f
C13019 VPWR.n1341 VGND 0.02657f
C13020 VPWR.t266 VGND 0.01056f
C13021 VPWR.t429 VGND 0.01056f
C13022 VPWR.n1342 VGND 0.02308f
C13023 VPWR.n1343 VGND 0.02937f
C13024 VPWR.n1345 VGND 0.03136f
C13025 VPWR.n1346 VGND 0.01183f
C13026 VPWR.t299 VGND 0.03543f
C13027 VPWR.t468 VGND 0.07971f
C13028 VPWR.t917 VGND 0.09299f
C13029 VPWR.t470 VGND 0.1727f
C13030 VPWR.t1370 VGND 0.09292f
C13031 VPWR.t472 VGND 0.10548f
C13032 VPWR.t319 VGND 0.10254f
C13033 VPWR.t317 VGND 0.164f
C13034 VPWR.t1835 VGND 0.13949f
C13035 VPWR.t1347 VGND 0.09299f
C13036 VPWR.t624 VGND 0.09299f
C13037 VPWR.t428 VGND 0.09299f
C13038 VPWR.t1831 VGND 0.09299f
C13039 VPWR.t265 VGND 0.09299f
C13040 VPWR.t449 VGND 0.09299f
C13041 VPWR.t263 VGND 0.09188f
C13042 VPWR.n1348 VGND 0.31603f
C13043 VPWR.n1349 VGND 0.12841f
C13044 VPWR.n1350 VGND 0.01408f
C13045 VPWR.n1351 VGND 0.02591f
C13046 VPWR.n1352 VGND 0.03117f
C13047 VPWR.n1354 VGND 0.04686f
C13048 VPWR.n1355 VGND 0.23333f
C13049 VPWR.n1356 VGND 1.20965f
C13050 VPWR.t1404 VGND 0.04142f
C13051 VPWR.t1318 VGND 0.0413f
C13052 VPWR.t605 VGND 0.04212f
C13053 VPWR.n1357 VGND 0.0587f
C13054 VPWR.t37 VGND 0.04022f
C13055 VPWR.t108 VGND 0.04022f
C13056 VPWR.n1358 VGND 0.07296f
C13057 VPWR.n1359 VGND 0.03455f
C13058 VPWR.n1361 VGND 0.03455f
C13059 VPWR.t33 VGND 0.01056f
C13060 VPWR.t403 VGND 0.01056f
C13061 VPWR.n1362 VGND 0.02308f
C13062 VPWR.t109 VGND 0.01056f
C13063 VPWR.t889 VGND 0.01056f
C13064 VPWR.n1363 VGND 0.02308f
C13065 VPWR.n1364 VGND 0.04703f
C13066 VPWR.t891 VGND 0.04212f
C13067 VPWR.t474 VGND 0.04212f
C13068 VPWR.n1365 VGND 0.09708f
C13069 VPWR.n1366 VGND 0.02028f
C13070 VPWR.n1367 VGND 0.03455f
C13071 VPWR.t260 VGND 0.01056f
C13072 VPWR.t1367 VGND 0.01056f
C13073 VPWR.n1369 VGND 0.02308f
C13074 VPWR.t894 VGND 0.01056f
C13075 VPWR.t277 VGND 0.01056f
C13076 VPWR.n1370 VGND 0.02308f
C13077 VPWR.n1371 VGND 0.05314f
C13078 VPWR.n1373 VGND 0.03455f
C13079 VPWR.n1374 VGND 0.03455f
C13080 VPWR.n1375 VGND 0.03455f
C13081 VPWR.t31 VGND 0.01056f
C13082 VPWR.t34 VGND 0.01056f
C13083 VPWR.n1377 VGND 0.02308f
C13084 VPWR.t104 VGND 0.01056f
C13085 VPWR.t103 VGND 0.01056f
C13086 VPWR.n1378 VGND 0.02308f
C13087 VPWR.n1379 VGND 0.04703f
C13088 VPWR.n1382 VGND 0.03455f
C13089 VPWR.n1383 VGND 0.02591f
C13090 VPWR.t30 VGND 0.71923f
C13091 VPWR.n1385 VGND 0.39227f
C13092 VPWR.t102 VGND 0.71923f
C13093 VPWR.n1386 VGND 0.30507f
C13094 VPWR.n1387 VGND 0.21437f
C13095 VPWR.n1388 VGND 0.01408f
C13096 VPWR.n1389 VGND 0.02591f
C13097 VPWR.n1390 VGND 0.03136f
C13098 VPWR.n1392 VGND 0.04296f
C13099 VPWR.n1393 VGND 0.05819f
C13100 VPWR.n1394 VGND 0.23314f
C13101 VPWR.n1395 VGND 1.20965f
C13102 VPWR.t707 VGND 0.04208f
C13103 VPWR.t1268 VGND 0.04208f
C13104 VPWR.n1396 VGND 0.01031f
C13105 VPWR.t161 VGND 0.04022f
C13106 VPWR.t659 VGND 0.04022f
C13107 VPWR.n1397 VGND 0.07296f
C13108 VPWR.n1398 VGND 0.03455f
C13109 VPWR.n1400 VGND 0.03455f
C13110 VPWR.t166 VGND 0.01056f
C13111 VPWR.t892 VGND 0.01056f
C13112 VPWR.n1401 VGND 0.02308f
C13113 VPWR.t1105 VGND 0.01056f
C13114 VPWR.t475 VGND 0.01056f
C13115 VPWR.n1402 VGND 0.02308f
C13116 VPWR.n1403 VGND 0.04703f
C13117 VPWR.t401 VGND 0.04212f
C13118 VPWR.t269 VGND 0.04212f
C13119 VPWR.n1404 VGND 0.09708f
C13120 VPWR.n1405 VGND 0.02028f
C13121 VPWR.n1406 VGND 0.03455f
C13122 VPWR.t896 VGND 0.01056f
C13123 VPWR.t278 VGND 0.01056f
C13124 VPWR.n1408 VGND 0.02308f
C13125 VPWR.t402 VGND 0.01056f
C13126 VPWR.t262 VGND 0.01056f
C13127 VPWR.n1409 VGND 0.02308f
C13128 VPWR.n1410 VGND 0.05314f
C13129 VPWR.n1412 VGND 0.03455f
C13130 VPWR.n1413 VGND 0.03455f
C13131 VPWR.n1414 VGND 0.03455f
C13132 VPWR.t167 VGND 0.01056f
C13133 VPWR.t164 VGND 0.01056f
C13134 VPWR.n1416 VGND 0.02308f
C13135 VPWR.t211 VGND 0.01056f
C13136 VPWR.t1106 VGND 0.01056f
C13137 VPWR.n1417 VGND 0.02308f
C13138 VPWR.n1418 VGND 0.04703f
C13139 VPWR.n1421 VGND 0.03455f
C13140 VPWR.n1422 VGND 0.02591f
C13141 VPWR.t160 VGND 0.71923f
C13142 VPWR.n1424 VGND 0.39227f
C13143 VPWR.t210 VGND 0.71923f
C13144 VPWR.n1425 VGND 0.30507f
C13145 VPWR.n1426 VGND 0.2163f
C13146 VPWR.n1427 VGND 0.01408f
C13147 VPWR.n1428 VGND 0.02591f
C13148 VPWR.n1429 VGND 0.03136f
C13149 VPWR.n1431 VGND 0.08505f
C13150 VPWR.n1432 VGND 0.2369f
C13151 VPWR.n1433 VGND 1.20965f
C13152 VPWR.t118 VGND 0.04022f
C13153 VPWR.t764 VGND 0.04022f
C13154 VPWR.n1434 VGND 0.07296f
C13155 VPWR.n1435 VGND 0.03455f
C13156 VPWR.n1437 VGND 0.03455f
C13157 VPWR.t112 VGND 0.01056f
C13158 VPWR.t404 VGND 0.01056f
C13159 VPWR.n1438 VGND 0.02308f
C13160 VPWR.t765 VGND 0.01056f
C13161 VPWR.t1369 VGND 0.01056f
C13162 VPWR.n1439 VGND 0.02308f
C13163 VPWR.n1440 VGND 0.04703f
C13164 VPWR.t893 VGND 0.04212f
C13165 VPWR.t430 VGND 0.04212f
C13166 VPWR.n1441 VGND 0.09708f
C13167 VPWR.n1442 VGND 0.02028f
C13168 VPWR.n1443 VGND 0.03455f
C13169 VPWR.t261 VGND 0.01056f
C13170 VPWR.t1368 VGND 0.01056f
C13171 VPWR.n1445 VGND 0.02308f
C13172 VPWR.t1372 VGND 0.01056f
C13173 VPWR.t268 VGND 0.01056f
C13174 VPWR.n1446 VGND 0.02308f
C13175 VPWR.n1447 VGND 0.05314f
C13176 VPWR.n1449 VGND 0.03455f
C13177 VPWR.n1450 VGND 0.03455f
C13178 VPWR.n1451 VGND 0.03455f
C13179 VPWR.t113 VGND 0.01056f
C13180 VPWR.t111 VGND 0.01056f
C13181 VPWR.n1453 VGND 0.02308f
C13182 VPWR.t768 VGND 0.01056f
C13183 VPWR.t767 VGND 0.01056f
C13184 VPWR.n1454 VGND 0.02308f
C13185 VPWR.n1455 VGND 0.04703f
C13186 VPWR.n1458 VGND 0.03455f
C13187 VPWR.n1459 VGND 0.02591f
C13188 VPWR.t110 VGND 0.55172f
C13189 VPWR.n1461 VGND 0.31566f
C13190 VPWR.t267 VGND 0.55172f
C13191 VPWR.n1462 VGND 0.24735f
C13192 VPWR.n1463 VGND 0.20736f
C13193 VPWR.n1464 VGND 0.31701f
C13194 VPWR.n1465 VGND 4.60935f
C13195 VPWR.n1466 VGND 6.74793f
C13196 VPWR.n1467 VGND 0.06156f
C13197 VPWR.n1468 VGND 0.81081f
C13198 VPWR.n1469 VGND 0.74411f
C13199 VPWR.n1470 VGND 0.04779f
C13200 VPWR.n1471 VGND 0.04011f
C13201 VPWR.n1472 VGND 0.02041f
C13202 VPWR.n1473 VGND 0.01398f
C13203 VPWR.n1474 VGND 0.04603f
C13204 VPWR.n1475 VGND 0.05722f
C13205 VPWR.n1476 VGND 0.06763f
C13206 VPWR.n1477 VGND 0.02041f
C13207 VPWR.n1478 VGND 0.01398f
C13208 VPWR.n1479 VGND 0.04603f
C13209 VPWR.n1480 VGND 0.07184f
C13210 VPWR.n1481 VGND 0.06763f
C13211 VPWR.n1482 VGND 0.04841f
C13212 VPWR.n1483 VGND 0.04011f
C13213 VPWR.n1484 VGND 0.10257f
C13214 VPWR.n1485 VGND 0.01325f
C13215 VPWR.n1487 VGND 0.07978f
C13216 VPWR.t1674 VGND 0.08814f
C13217 VPWR.t1637 VGND 0.05786f
C13218 VPWR.t1336 VGND 0.06796f
C13219 VPWR.n1488 VGND 0.02243f
C13220 VPWR.t1675 VGND 0.01975f
C13221 VPWR.n1490 VGND 0.04219f
C13222 VPWR.t1337 VGND 0.02183f
C13223 VPWR.n1491 VGND 0.03459f
C13224 VPWR.n1492 VGND 0.01325f
C13225 VPWR.n1494 VGND 0.07978f
C13226 VPWR.t1784 VGND 0.08814f
C13227 VPWR.t1766 VGND 0.05786f
C13228 VPWR.t1091 VGND 0.06796f
C13229 VPWR.n1495 VGND 0.02243f
C13230 VPWR.t1785 VGND 0.01975f
C13231 VPWR.n1497 VGND 0.04219f
C13232 VPWR.t1092 VGND 0.02183f
C13233 VPWR.n1498 VGND 0.03459f
C13234 VPWR.n1500 VGND 0.07978f
C13235 VPWR.t1555 VGND 0.08814f
C13236 VPWR.t1422 VGND 0.05786f
C13237 VPWR.t1400 VGND 0.06796f
C13238 VPWR.n1501 VGND 0.02243f
C13239 VPWR.t1556 VGND 0.01975f
C13240 VPWR.n1503 VGND 0.04219f
C13241 VPWR.t1401 VGND 0.02183f
C13242 VPWR.n1504 VGND 0.03459f
C13243 VPWR.n1506 VGND 0.06156f
C13244 VPWR.n1507 VGND -0.01375f
C13245 VPWR.n1508 VGND 0.10257f
C13246 VPWR.n1509 VGND 0.01325f
C13247 VPWR.n1511 VGND 0.07978f
C13248 VPWR.t1657 VGND 0.08814f
C13249 VPWR.t1532 VGND 0.05786f
C13250 VPWR.t1147 VGND 0.06796f
C13251 VPWR.t1687 VGND 0.05786f
C13252 VPWR.t1682 VGND 0.08814f
C13253 VPWR.n1512 VGND 0.07978f
C13254 VPWR.n1514 VGND 0.01325f
C13255 VPWR.n1515 VGND 0.04011f
C13256 VPWR.n1516 VGND 0.10257f
C13257 VPWR.n1517 VGND -0.01375f
C13258 VPWR.n1518 VGND 0.06156f
C13259 VPWR.n1519 VGND 0.06156f
C13260 VPWR.n1520 VGND -0.01375f
C13261 VPWR.n1521 VGND 0.04011f
C13262 VPWR.n1522 VGND 0.10257f
C13263 VPWR.n1523 VGND 0.01325f
C13264 VPWR.n1525 VGND 0.07978f
C13265 VPWR.t1430 VGND 0.08814f
C13266 VPWR.t1689 VGND 0.05786f
C13267 VPWR.t1394 VGND 0.06796f
C13268 VPWR.t1537 VGND 0.05786f
C13269 VPWR.t1552 VGND 0.08814f
C13270 VPWR.n1526 VGND 0.07978f
C13271 VPWR.n1528 VGND 0.01325f
C13272 VPWR.n1529 VGND 0.04011f
C13273 VPWR.n1530 VGND 0.10257f
C13274 VPWR.n1531 VGND -0.01375f
C13275 VPWR.n1532 VGND 0.06156f
C13276 VPWR.n1533 VGND 0.06156f
C13277 VPWR.n1534 VGND -0.01375f
C13278 VPWR.n1535 VGND 0.04011f
C13279 VPWR.n1536 VGND 0.10257f
C13280 VPWR.n1537 VGND 0.01325f
C13281 VPWR.n1539 VGND 0.07978f
C13282 VPWR.t1693 VGND 0.08814f
C13283 VPWR.t1567 VGND 0.05786f
C13284 VPWR.t297 VGND 0.06796f
C13285 VPWR.t1685 VGND 0.05786f
C13286 VPWR.t1715 VGND 0.08814f
C13287 VPWR.n1540 VGND 0.07978f
C13288 VPWR.n1542 VGND 0.01325f
C13289 VPWR.n1543 VGND 0.04011f
C13290 VPWR.n1544 VGND 0.10257f
C13291 VPWR.n1545 VGND -0.01375f
C13292 VPWR.n1546 VGND 0.06156f
C13293 VPWR.n1547 VGND 0.06156f
C13294 VPWR.n1548 VGND 0.06156f
C13295 VPWR.n1549 VGND 0.06156f
C13296 VPWR.n1550 VGND -0.01375f
C13297 VPWR.n1551 VGND 0.10257f
C13298 VPWR.n1552 VGND 0.01325f
C13299 VPWR.n1554 VGND 0.07978f
C13300 VPWR.t1845 VGND 0.06796f
C13301 VPWR.t1436 VGND 0.05786f
C13302 VPWR.t1449 VGND 0.08814f
C13303 VPWR.n1555 VGND 0.07978f
C13304 VPWR.n1557 VGND 0.01325f
C13305 VPWR.n1558 VGND 0.10257f
C13306 VPWR.n1559 VGND 0.04011f
C13307 VPWR.n1560 VGND 0.04841f
C13308 VPWR.n1561 VGND 0.06763f
C13309 VPWR.n1562 VGND 0.02041f
C13310 VPWR.n1563 VGND 0.01398f
C13311 VPWR.n1564 VGND 0.04603f
C13312 VPWR.n1565 VGND 0.07184f
C13313 VPWR.n1566 VGND 0.06763f
C13314 VPWR.n1567 VGND 0.02041f
C13315 VPWR.n1568 VGND 0.01398f
C13316 VPWR.n1569 VGND 0.04603f
C13317 VPWR.n1570 VGND 0.07184f
C13318 VPWR.n1571 VGND 0.06763f
C13319 VPWR.n1572 VGND 0.02041f
C13320 VPWR.n1573 VGND 0.01398f
C13321 VPWR.n1574 VGND 0.04603f
C13322 VPWR.n1575 VGND 0.07184f
C13323 VPWR.n1576 VGND 0.06763f
C13324 VPWR.n1577 VGND 0.02041f
C13325 VPWR.n1578 VGND 0.01398f
C13326 VPWR.n1579 VGND 0.04603f
C13327 VPWR.n1580 VGND 0.07184f
C13328 VPWR.n1581 VGND 0.06763f
C13329 VPWR.n1582 VGND 0.02041f
C13330 VPWR.n1583 VGND 0.01398f
C13331 VPWR.n1584 VGND 0.04603f
C13332 VPWR.n1585 VGND 0.07184f
C13333 VPWR.n1586 VGND 0.06763f
C13334 VPWR.n1587 VGND 0.02041f
C13335 VPWR.n1588 VGND 0.01398f
C13336 VPWR.n1589 VGND 0.04603f
C13337 VPWR.n1590 VGND 0.07184f
C13338 VPWR.n1591 VGND 0.06763f
C13339 VPWR.n1592 VGND 0.02041f
C13340 VPWR.n1593 VGND 0.01398f
C13341 VPWR.n1594 VGND 0.04603f
C13342 VPWR.n1595 VGND 0.07184f
C13343 VPWR.n1596 VGND 0.06763f
C13344 VPWR.n1597 VGND 0.02041f
C13345 VPWR.n1598 VGND 0.01398f
C13346 VPWR.n1599 VGND 0.04603f
C13347 VPWR.n1600 VGND 0.07184f
C13348 VPWR.n1601 VGND 0.06763f
C13349 VPWR.n1602 VGND 0.04841f
C13350 VPWR.n1603 VGND 0.04011f
C13351 VPWR.n1604 VGND 0.10257f
C13352 VPWR.n1605 VGND -0.01375f
C13353 VPWR.n1606 VGND 0.06156f
C13354 VPWR.n1607 VGND 0.06156f
C13355 VPWR.n1608 VGND -0.01375f
C13356 VPWR.n1610 VGND 0.01264f
C13357 VPWR.n1612 VGND 0.07978f
C13358 VPWR.t1579 VGND 0.06796f
C13359 VPWR.t1457 VGND 0.05786f
C13360 VPWR.t1493 VGND 0.08814f
C13361 VPWR.n1613 VGND 0.07978f
C13362 VPWR.n1615 VGND 0.01264f
C13363 VPWR.n1616 VGND 0.02534f
C13364 VPWR.n1617 VGND 0.02297f
C13365 VPWR.n1618 VGND 0.02723f
C13366 VPWR.n1620 VGND 0.0204f
C13367 VPWR.n1621 VGND 0.02077f
C13368 VPWR.n1622 VGND 0.01309f
C13369 VPWR.n1624 VGND 0.01343f
C13370 VPWR.n1625 VGND 0.01757f
C13371 VPWR.n1626 VGND 0.17489f
C13372 VPWR.n1627 VGND 0.12963f
C13373 VPWR.n1628 VGND 0.01757f
C13374 VPWR.n1629 VGND 0.01309f
C13375 VPWR.n1630 VGND 0.02206f
C13376 VPWR.n1631 VGND 0.02421f
C13377 VPWR.n1632 VGND 0.02534f
C13378 VPWR.n1633 VGND 0.02297f
C13379 VPWR.n1634 VGND 0.02723f
C13380 VPWR.n1636 VGND 0.0204f
C13381 VPWR.n1637 VGND 0.02077f
C13382 VPWR.n1638 VGND 0.01343f
C13383 VPWR.n1639 VGND 0.01757f
C13384 VPWR.n1640 VGND 0.01309f
C13385 VPWR.n1641 VGND 0.02206f
C13386 VPWR.n1642 VGND 0.02421f
C13387 VPWR.n1643 VGND 0.02534f
C13388 VPWR.n1644 VGND 0.02297f
C13389 VPWR.n1645 VGND 0.02723f
C13390 VPWR.n1647 VGND 0.0204f
C13391 VPWR.n1648 VGND 0.02077f
C13392 VPWR.n1649 VGND 0.01309f
C13393 VPWR.n1651 VGND 0.01343f
C13394 VPWR.n1652 VGND 0.01757f
C13395 VPWR.n1653 VGND 0.12963f
C13396 VPWR.n1654 VGND 0.12963f
C13397 VPWR.n1655 VGND 0.01757f
C13398 VPWR.n1656 VGND 0.01309f
C13399 VPWR.n1657 VGND 0.02206f
C13400 VPWR.n1658 VGND 0.02421f
C13401 VPWR.n1659 VGND 0.02534f
C13402 VPWR.n1660 VGND 0.02297f
C13403 VPWR.n1661 VGND 0.02723f
C13404 VPWR.n1663 VGND 0.0204f
C13405 VPWR.n1664 VGND 0.02077f
C13406 VPWR.n1665 VGND 0.01343f
C13407 VPWR.n1666 VGND 0.01757f
C13408 VPWR.n1667 VGND 0.01309f
C13409 VPWR.n1668 VGND 0.02206f
C13410 VPWR.n1669 VGND 0.02421f
C13411 VPWR.n1670 VGND 0.02534f
C13412 VPWR.n1671 VGND 0.02297f
C13413 VPWR.n1672 VGND 0.02723f
C13414 VPWR.n1674 VGND 0.0204f
C13415 VPWR.n1675 VGND 0.02077f
C13416 VPWR.n1676 VGND 0.01309f
C13417 VPWR.n1678 VGND 0.01343f
C13418 VPWR.n1679 VGND 0.01757f
C13419 VPWR.n1680 VGND 0.12963f
C13420 VPWR.n1681 VGND 0.12963f
C13421 VPWR.n1682 VGND 0.01757f
C13422 VPWR.n1683 VGND 0.01309f
C13423 VPWR.n1684 VGND 0.02206f
C13424 VPWR.n1685 VGND 0.02421f
C13425 VPWR.n1686 VGND 0.02534f
C13426 VPWR.n1687 VGND 0.02297f
C13427 VPWR.n1688 VGND 0.02723f
C13428 VPWR.n1690 VGND 0.0204f
C13429 VPWR.n1691 VGND 0.02077f
C13430 VPWR.n1692 VGND 0.01343f
C13431 VPWR.n1693 VGND 0.01757f
C13432 VPWR.n1694 VGND 0.01309f
C13433 VPWR.n1695 VGND 0.02206f
C13434 VPWR.n1696 VGND 0.02421f
C13435 VPWR.n1697 VGND 0.02534f
C13436 VPWR.n1698 VGND 0.02297f
C13437 VPWR.n1699 VGND 0.02723f
C13438 VPWR.n1701 VGND 0.0204f
C13439 VPWR.n1702 VGND 0.02077f
C13440 VPWR.n1703 VGND 0.01309f
C13441 VPWR.n1705 VGND 0.01343f
C13442 VPWR.n1706 VGND 0.01757f
C13443 VPWR.n1707 VGND 0.12963f
C13444 VPWR.n1708 VGND 0.12963f
C13445 VPWR.n1709 VGND 0.01757f
C13446 VPWR.n1710 VGND 0.01309f
C13447 VPWR.n1711 VGND 0.02206f
C13448 VPWR.n1712 VGND 0.02421f
C13449 VPWR.n1713 VGND 0.02534f
C13450 VPWR.n1714 VGND 0.02297f
C13451 VPWR.n1715 VGND 0.02723f
C13452 VPWR.n1717 VGND 0.0204f
C13453 VPWR.n1718 VGND 0.02077f
C13454 VPWR.n1719 VGND 0.01343f
C13455 VPWR.n1720 VGND 0.01757f
C13456 VPWR.n1721 VGND 0.01309f
C13457 VPWR.n1722 VGND 0.02206f
C13458 VPWR.n1723 VGND 0.02421f
C13459 VPWR.n1724 VGND 0.02534f
C13460 VPWR.n1725 VGND 0.02297f
C13461 VPWR.n1726 VGND 0.02723f
C13462 VPWR.n1728 VGND 0.0204f
C13463 VPWR.n1729 VGND 0.02077f
C13464 VPWR.n1730 VGND 0.01309f
C13465 VPWR.n1732 VGND 0.01343f
C13466 VPWR.n1733 VGND 0.01757f
C13467 VPWR.n1734 VGND 0.12963f
C13468 VPWR.n1735 VGND 0.02206f
C13469 VPWR.n1736 VGND 0.02421f
C13470 VPWR.n1737 VGND 0.02297f
C13471 VPWR.n1738 VGND 0.02723f
C13472 VPWR.n1740 VGND 0.0204f
C13473 VPWR.n1741 VGND 0.02077f
C13474 VPWR.n1742 VGND 0.01309f
C13475 VPWR.n1744 VGND 0.01343f
C13476 VPWR.n1745 VGND 0.01757f
C13477 VPWR.n1746 VGND 0.15601f
C13478 VPWR.n1747 VGND 0.01873f
C13479 VPWR.n1748 VGND 0.01309f
C13480 VPWR.n1749 VGND 0.0204f
C13481 VPWR.n1750 VGND 0.02077f
C13482 VPWR.n1752 VGND 0.02297f
C13483 VPWR.n1753 VGND 0.02723f
C13484 VPWR.n1754 VGND 0.02534f
C13485 VPWR.n1756 VGND 0.01264f
C13486 VPWR.n1758 VGND 0.07978f
C13487 VPWR.t1702 VGND 0.06796f
C13488 VPWR.t1575 VGND 0.05786f
C13489 VPWR.t1710 VGND 0.08814f
C13490 VPWR.n1759 VGND 0.07978f
C13491 VPWR.n1761 VGND 0.01264f
C13492 VPWR.n1763 VGND 0.04011f
C13493 VPWR.n1764 VGND 0.02243f
C13494 VPWR.t1460 VGND 0.01975f
C13495 VPWR.n1766 VGND 0.04219f
C13496 VPWR.t982 VGND 0.02183f
C13497 VPWR.n1767 VGND 0.03459f
C13498 VPWR.t1723 VGND 0.05786f
C13499 VPWR.t981 VGND 0.06796f
C13500 VPWR.t1758 VGND 0.05786f
C13501 VPWR.t1496 VGND 0.08814f
C13502 VPWR.n1768 VGND 0.07978f
C13503 VPWR.n1770 VGND 0.01325f
C13504 VPWR.n1771 VGND 0.10257f
C13505 VPWR.n1772 VGND -0.01375f
C13506 VPWR.n1773 VGND 0.06156f
C13507 VPWR.n1774 VGND 0.06156f
C13508 VPWR.n1775 VGND -0.01375f
C13509 VPWR.n1776 VGND 0.10257f
C13510 VPWR.n1777 VGND 0.01325f
C13511 VPWR.n1779 VGND 0.07978f
C13512 VPWR.t189 VGND 0.06796f
C13513 VPWR.t1705 VGND 0.05786f
C13514 VPWR.t1623 VGND 0.08814f
C13515 VPWR.n1780 VGND 0.07978f
C13516 VPWR.n1782 VGND 0.01325f
C13517 VPWR.n1783 VGND 0.10257f
C13518 VPWR.n1784 VGND 0.04011f
C13519 VPWR.n1785 VGND 0.04841f
C13520 VPWR.n1786 VGND 0.06763f
C13521 VPWR.n1787 VGND 0.02041f
C13522 VPWR.n1788 VGND 0.01398f
C13523 VPWR.n1789 VGND 0.04603f
C13524 VPWR.n1790 VGND 0.07184f
C13525 VPWR.n1791 VGND 0.06763f
C13526 VPWR.n1792 VGND 0.02041f
C13527 VPWR.n1793 VGND 0.01398f
C13528 VPWR.n1794 VGND 0.04603f
C13529 VPWR.n1795 VGND 0.07184f
C13530 VPWR.n1796 VGND 0.02041f
C13531 VPWR.n1797 VGND 0.01398f
C13532 VPWR.n1798 VGND 0.04602f
C13533 VPWR.n1799 VGND 0.03788f
C13534 VPWR.n1800 VGND 0.02041f
C13535 VPWR.n1801 VGND 0.01398f
C13536 VPWR.n1802 VGND 0.04603f
C13537 VPWR.n1803 VGND 0.07184f
C13538 VPWR.n1804 VGND 0.06763f
C13539 VPWR.n1805 VGND 0.04841f
C13540 VPWR.n1806 VGND 0.04011f
C13541 VPWR.n1807 VGND 0.10257f
C13542 VPWR.n1808 VGND 0.01325f
C13543 VPWR.n1810 VGND 0.07978f
C13544 VPWR.t1604 VGND 0.08814f
C13545 VPWR.t1587 VGND 0.05786f
C13546 VPWR.t1718 VGND 0.09829f
C13547 VPWR.n1811 VGND 0.05616f
C13548 VPWR.n1812 VGND 0.01325f
C13549 VPWR.n1813 VGND 0.10257f
C13550 VPWR.n1814 VGND 0.12134f
C13551 VPWR.n1815 VGND 0.7488f
C13552 VPWR.n1816 VGND 0.06156f
C13553 VPWR.n1817 VGND 0.06156f
C13554 VPWR.n1818 VGND 0.06156f
C13555 VPWR.n1819 VGND 0.06156f
C13556 VPWR.n1820 VGND 0.06156f
C13557 VPWR.n1821 VGND 0.06156f
C13558 VPWR.n1822 VGND 0.06156f
C13559 VPWR.n1823 VGND 0.06156f
C13560 VPWR.n1824 VGND 0.06156f
C13561 VPWR.n1825 VGND 0.06156f
C13562 VPWR.n1826 VGND 0.06156f
C13563 VPWR.n1827 VGND 0.06156f
C13564 VPWR.n1828 VGND 0.06156f
C13565 VPWR.n1829 VGND 0.06156f
C13566 VPWR.n1830 VGND 0.06156f
C13567 VPWR.n1831 VGND 0.1428f
C13568 VPWR.n1832 VGND 0.7488f
C13569 VPWR.n1833 VGND 0.7488f
C13570 VPWR.n1834 VGND 0.1428f
C13571 VPWR.n1835 VGND 0.10257f
C13572 VPWR.n1836 VGND 0.01325f
C13573 VPWR.n1837 VGND 0.05616f
C13574 VPWR.t1749 VGND 0.09829f
C13575 VPWR.t1356 VGND 0.05786f
C13576 VPWR.t821 VGND 0.08814f
C13577 VPWR.n1838 VGND 0.07978f
C13578 VPWR.n1840 VGND 0.01325f
C13579 VPWR.n1841 VGND 0.10257f
C13580 VPWR.n1842 VGND 0.06156f
C13581 VPWR.n1843 VGND 0.06156f
C13582 VPWR.n1844 VGND 0.10257f
C13583 VPWR.n1845 VGND 0.01325f
C13584 VPWR.n1847 VGND 0.07978f
C13585 VPWR.t993 VGND 0.06796f
C13586 VPWR.t171 VGND 0.05786f
C13587 VPWR.t1310 VGND 0.08814f
C13588 VPWR.n1848 VGND 0.07978f
C13589 VPWR.n1850 VGND 0.01325f
C13590 VPWR.n1851 VGND 0.10257f
C13591 VPWR.n1852 VGND 0.06156f
C13592 VPWR.n1853 VGND 0.06156f
C13593 VPWR.n1854 VGND 0.10257f
C13594 VPWR.n1855 VGND 0.01325f
C13595 VPWR.n1857 VGND 0.07978f
C13596 VPWR.t1027 VGND 0.06796f
C13597 VPWR.t1134 VGND 0.05786f
C13598 VPWR.t482 VGND 0.08814f
C13599 VPWR.n1858 VGND 0.07978f
C13600 VPWR.n1860 VGND 0.01325f
C13601 VPWR.n1861 VGND 0.10257f
C13602 VPWR.n1862 VGND 0.06156f
C13603 VPWR.n1863 VGND 0.06156f
C13604 VPWR.n1864 VGND 0.10257f
C13605 VPWR.n1865 VGND 0.01325f
C13606 VPWR.n1867 VGND 0.07978f
C13607 VPWR.t362 VGND 0.06796f
C13608 VPWR.t1354 VGND 0.05786f
C13609 VPWR.t1277 VGND 0.08814f
C13610 VPWR.n1868 VGND 0.07978f
C13611 VPWR.n1870 VGND 0.01325f
C13612 VPWR.n1871 VGND 0.10257f
C13613 VPWR.n1872 VGND 0.06156f
C13614 VPWR.n1873 VGND 0.06156f
C13615 VPWR.n1874 VGND 0.10257f
C13616 VPWR.n1875 VGND 0.01325f
C13617 VPWR.n1877 VGND 0.07978f
C13618 VPWR.t932 VGND 0.06796f
C13619 VPWR.t1358 VGND 0.05786f
C13620 VPWR.t1380 VGND 0.08814f
C13621 VPWR.n1878 VGND 0.07978f
C13622 VPWR.n1880 VGND 0.01325f
C13623 VPWR.n1881 VGND 0.10257f
C13624 VPWR.n1882 VGND 0.06156f
C13625 VPWR.n1883 VGND 0.06156f
C13626 VPWR.n1884 VGND 0.10257f
C13627 VPWR.n1885 VGND 0.01325f
C13628 VPWR.n1887 VGND 0.07978f
C13629 VPWR.t1827 VGND 0.06796f
C13630 VPWR.t174 VGND 0.05786f
C13631 VPWR.t899 VGND 0.08814f
C13632 VPWR.n1888 VGND 0.07978f
C13633 VPWR.n1890 VGND 0.01325f
C13634 VPWR.n1891 VGND 0.10257f
C13635 VPWR.n1892 VGND 0.06156f
C13636 VPWR.n1893 VGND 0.06156f
C13637 VPWR.n1894 VGND 0.10257f
C13638 VPWR.n1895 VGND 0.01325f
C13639 VPWR.n1897 VGND 0.07978f
C13640 VPWR.t679 VGND 0.06796f
C13641 VPWR.t1136 VGND 0.05786f
C13642 VPWR.t1063 VGND 0.08814f
C13643 VPWR.n1898 VGND 0.07978f
C13644 VPWR.n1900 VGND 0.01325f
C13645 VPWR.n1901 VGND 0.10257f
C13646 VPWR.n1902 VGND 0.06156f
C13647 VPWR.n1903 VGND 0.06156f
C13648 VPWR.n1904 VGND 0.10257f
C13649 VPWR.n1905 VGND 0.01325f
C13650 VPWR.n1907 VGND 0.07978f
C13651 VPWR.t1118 VGND 0.06796f
C13652 VPWR.t1355 VGND 0.05786f
C13653 VPWR.t1128 VGND 0.08814f
C13654 VPWR.n1908 VGND 0.07978f
C13655 VPWR.n1910 VGND 0.01325f
C13656 VPWR.n1911 VGND 0.10257f
C13657 VPWR.n1912 VGND 0.06156f
C13658 VPWR.n1913 VGND 0.74411f
C13659 VPWR.n1914 VGND 0.1428f
C13660 VPWR.n1915 VGND 0.06156f
C13661 VPWR.n1916 VGND 0.06156f
C13662 VPWR.n1917 VGND 0.06156f
C13663 VPWR.n1918 VGND 0.06156f
C13664 VPWR.n1919 VGND 0.06156f
C13665 VPWR.n1920 VGND 0.06156f
C13666 VPWR.n1921 VGND 0.06156f
C13667 VPWR.n1922 VGND 0.06156f
C13668 VPWR.n1923 VGND 0.06156f
C13669 VPWR.n1924 VGND 0.06156f
C13670 VPWR.n1925 VGND 0.06156f
C13671 VPWR.n1926 VGND 0.06156f
C13672 VPWR.n1927 VGND 0.06156f
C13673 VPWR.n1928 VGND 0.06156f
C13674 VPWR.n1929 VGND 0.06156f
C13675 VPWR.n1930 VGND 0.74411f
C13676 VPWR.n1931 VGND 0.74411f
C13677 VPWR.n1932 VGND 0.06156f
C13678 VPWR.n1933 VGND 0.10257f
C13679 VPWR.n1934 VGND 0.01325f
C13680 VPWR.n1936 VGND 0.07978f
C13681 VPWR.t72 VGND 0.08814f
C13682 VPWR.t451 VGND 0.05786f
C13683 VPWR.t1159 VGND 0.06796f
C13684 VPWR.t814 VGND 0.05786f
C13685 VPWR.t1153 VGND 0.08814f
C13686 VPWR.n1937 VGND 0.07978f
C13687 VPWR.n1939 VGND 0.01325f
C13688 VPWR.n1940 VGND 0.10257f
C13689 VPWR.n1941 VGND 0.06156f
C13690 VPWR.n1942 VGND 0.06156f
C13691 VPWR.n1943 VGND 0.10257f
C13692 VPWR.n1944 VGND 0.01325f
C13693 VPWR.n1946 VGND 0.07978f
C13694 VPWR.t1079 VGND 0.08814f
C13695 VPWR.t813 VGND 0.05786f
C13696 VPWR.t755 VGND 0.06796f
C13697 VPWR.t537 VGND 0.05786f
C13698 VPWR.t685 VGND 0.08814f
C13699 VPWR.n1947 VGND 0.07978f
C13700 VPWR.n1949 VGND 0.01325f
C13701 VPWR.n1950 VGND 0.10257f
C13702 VPWR.n1951 VGND 0.06156f
C13703 VPWR.n1952 VGND 0.06156f
C13704 VPWR.n1953 VGND 0.10257f
C13705 VPWR.n1954 VGND 0.01325f
C13706 VPWR.n1956 VGND 0.07978f
C13707 VPWR.t1325 VGND 0.08814f
C13708 VPWR.t819 VGND 0.05786f
C13709 VPWR.t845 VGND 0.06796f
C13710 VPWR.t818 VGND 0.05786f
C13711 VPWR.t1101 VGND 0.08814f
C13712 VPWR.n1957 VGND 0.07978f
C13713 VPWR.n1959 VGND 0.01325f
C13714 VPWR.n1960 VGND 0.10257f
C13715 VPWR.n1961 VGND 0.06156f
C13716 VPWR.n1962 VGND 0.06156f
C13717 VPWR.n1963 VGND 0.10257f
C13718 VPWR.n1964 VGND 0.01325f
C13719 VPWR.n1966 VGND 0.07978f
C13720 VPWR.t1901 VGND 0.08814f
C13721 VPWR.t536 VGND 0.05786f
C13722 VPWR.t242 VGND 0.06796f
C13723 VPWR.t535 VGND 0.05786f
C13724 VPWR.t224 VGND 0.08814f
C13725 VPWR.n1967 VGND 0.07978f
C13726 VPWR.n1969 VGND 0.01325f
C13727 VPWR.n1970 VGND 0.10257f
C13728 VPWR.n1971 VGND 0.06156f
C13729 VPWR.n1972 VGND 0.06156f
C13730 VPWR.n1973 VGND 0.10257f
C13731 VPWR.n1974 VGND 0.01325f
C13732 VPWR.n1976 VGND 0.07978f
C13733 VPWR.t796 VGND 0.08814f
C13734 VPWR.t820 VGND 0.05786f
C13735 VPWR.t381 VGND 0.06796f
C13736 VPWR.t540 VGND 0.05786f
C13737 VPWR.t348 VGND 0.08814f
C13738 VPWR.n1977 VGND 0.07978f
C13739 VPWR.n1979 VGND 0.01325f
C13740 VPWR.n1980 VGND 0.10257f
C13741 VPWR.n1981 VGND 0.06156f
C13742 VPWR.n1982 VGND 0.06156f
C13743 VPWR.n1983 VGND 0.10257f
C13744 VPWR.n1984 VGND 0.01325f
C13745 VPWR.n1986 VGND 0.07978f
C13746 VPWR.t1411 VGND 0.08814f
C13747 VPWR.t539 VGND 0.05786f
C13748 VPWR.t1811 VGND 0.06796f
C13749 VPWR.t817 VGND 0.05786f
C13750 VPWR.t1805 VGND 0.08814f
C13751 VPWR.n1987 VGND 0.07978f
C13752 VPWR.n1989 VGND 0.01325f
C13753 VPWR.n1990 VGND 0.10257f
C13754 VPWR.n1991 VGND 0.06156f
C13755 VPWR.n1992 VGND 0.06156f
C13756 VPWR.n1993 VGND 0.10257f
C13757 VPWR.n1994 VGND 0.01325f
C13758 VPWR.n1996 VGND 0.07978f
C13759 VPWR.t256 VGND 0.08814f
C13760 VPWR.t816 VGND 0.05786f
C13761 VPWR.t1197 VGND 0.06796f
C13762 VPWR.t815 VGND 0.05786f
C13763 VPWR.t1001 VGND 0.08814f
C13764 VPWR.n1997 VGND 0.07978f
C13765 VPWR.n1999 VGND 0.01325f
C13766 VPWR.n2000 VGND 0.10257f
C13767 VPWR.n2001 VGND 0.06156f
C13768 VPWR.n2002 VGND 0.06156f
C13769 VPWR.n2003 VGND 0.10257f
C13770 VPWR.n2004 VGND 0.01325f
C13771 VPWR.n2006 VGND 0.07978f
C13772 VPWR.t1243 VGND 0.08814f
C13773 VPWR.t534 VGND 0.05786f
C13774 VPWR.t1454 VGND 0.09829f
C13775 VPWR.n2007 VGND 0.05616f
C13776 VPWR.n2008 VGND 0.01325f
C13777 VPWR.n2009 VGND 0.10257f
C13778 VPWR.n2010 VGND 0.1428f
C13779 VPWR.n2011 VGND 0.7488f
C13780 VPWR.n2012 VGND 0.06156f
C13781 VPWR.n2013 VGND 0.06156f
C13782 VPWR.n2014 VGND 0.06156f
C13783 VPWR.n2015 VGND 0.06156f
C13784 VPWR.n2016 VGND 0.06156f
C13785 VPWR.n2017 VGND 0.06156f
C13786 VPWR.n2018 VGND 0.06156f
C13787 VPWR.n2019 VGND 0.06156f
C13788 VPWR.n2020 VGND 0.06156f
C13789 VPWR.n2021 VGND 0.06156f
C13790 VPWR.n2022 VGND 0.06156f
C13791 VPWR.n2023 VGND 0.06156f
C13792 VPWR.n2024 VGND 0.06156f
C13793 VPWR.n2025 VGND 0.06156f
C13794 VPWR.n2026 VGND 0.06156f
C13795 VPWR.n2027 VGND 0.1428f
C13796 VPWR.n2028 VGND 0.7488f
C13797 VPWR.n2029 VGND 0.7488f
C13798 VPWR.n2030 VGND 0.1428f
C13799 VPWR.n2031 VGND 0.10257f
C13800 VPWR.n2032 VGND 0.01325f
C13801 VPWR.n2033 VGND 0.05616f
C13802 VPWR.t1529 VGND 0.09829f
C13803 VPWR.t804 VGND 0.05786f
C13804 VPWR.t22 VGND 0.08814f
C13805 VPWR.n2034 VGND 0.07978f
C13806 VPWR.n2036 VGND 0.01325f
C13807 VPWR.n2037 VGND 0.10257f
C13808 VPWR.n2038 VGND 0.06156f
C13809 VPWR.n2039 VGND 0.06156f
C13810 VPWR.n2040 VGND 0.10257f
C13811 VPWR.n2041 VGND 0.01325f
C13812 VPWR.n2043 VGND 0.07978f
C13813 VPWR.t997 VGND 0.06796f
C13814 VPWR.t970 VGND 0.05786f
C13815 VPWR.t244 VGND 0.08814f
C13816 VPWR.n2044 VGND 0.07978f
C13817 VPWR.n2046 VGND 0.01325f
C13818 VPWR.n2047 VGND 0.10257f
C13819 VPWR.n2048 VGND 0.06156f
C13820 VPWR.n2049 VGND 0.06156f
C13821 VPWR.n2050 VGND 0.10257f
C13822 VPWR.n2051 VGND 0.01325f
C13823 VPWR.n2053 VGND 0.07978f
C13824 VPWR.t1161 VGND 0.06796f
C13825 VPWR.t965 VGND 0.05786f
C13826 VPWR.t532 VGND 0.08814f
C13827 VPWR.n2054 VGND 0.07978f
C13828 VPWR.n2056 VGND 0.01325f
C13829 VPWR.n2057 VGND 0.10257f
C13830 VPWR.n2058 VGND 0.06156f
C13831 VPWR.n2059 VGND 0.06156f
C13832 VPWR.n2060 VGND 0.10257f
C13833 VPWR.n2061 VGND 0.01325f
C13834 VPWR.n2063 VGND 0.07978f
C13835 VPWR.t344 VGND 0.06796f
C13836 VPWR.t1033 VGND 0.05786f
C13837 VPWR.t562 VGND 0.08814f
C13838 VPWR.n2064 VGND 0.07978f
C13839 VPWR.n2066 VGND 0.01325f
C13840 VPWR.n2067 VGND 0.10257f
C13841 VPWR.n2068 VGND 0.06156f
C13842 VPWR.n2069 VGND 0.06156f
C13843 VPWR.n2070 VGND 0.10257f
C13844 VPWR.n2071 VGND 0.01325f
C13845 VPWR.n2073 VGND 0.07978f
C13846 VPWR.t543 VGND 0.06796f
C13847 VPWR.t806 VGND 0.05786f
C13848 VPWR.t460 VGND 0.08814f
C13849 VPWR.n2074 VGND 0.07978f
C13850 VPWR.n2076 VGND 0.01325f
C13851 VPWR.n2077 VGND 0.10257f
C13852 VPWR.n2078 VGND 0.06156f
C13853 VPWR.n2079 VGND 0.06156f
C13854 VPWR.n2080 VGND 0.10257f
C13855 VPWR.n2081 VGND 0.01325f
C13856 VPWR.n2083 VGND 0.07978f
C13857 VPWR.t1097 VGND 0.06796f
C13858 VPWR.t1032 VGND 0.05786f
C13859 VPWR.t445 VGND 0.08814f
C13860 VPWR.n2084 VGND 0.07978f
C13861 VPWR.n2086 VGND 0.01325f
C13862 VPWR.n2087 VGND 0.10257f
C13863 VPWR.n2088 VGND 0.06156f
C13864 VPWR.n2089 VGND 0.06156f
C13865 VPWR.n2090 VGND 0.10257f
C13866 VPWR.n2091 VGND 0.01325f
C13867 VPWR.n2093 VGND 0.07978f
C13868 VPWR.t4 VGND 0.06796f
C13869 VPWR.t967 VGND 0.05786f
C13870 VPWR.t1089 VGND 0.08814f
C13871 VPWR.n2094 VGND 0.07978f
C13872 VPWR.n2096 VGND 0.01325f
C13873 VPWR.n2097 VGND 0.10257f
C13874 VPWR.n2098 VGND 0.06156f
C13875 VPWR.n2099 VGND 0.06156f
C13876 VPWR.n2100 VGND 0.10257f
C13877 VPWR.n2101 VGND 0.01325f
C13878 VPWR.n2103 VGND 0.07978f
C13879 VPWR.t508 VGND 0.06796f
C13880 VPWR.t1034 VGND 0.05786f
C13881 VPWR.t642 VGND 0.08814f
C13882 VPWR.n2104 VGND 0.07978f
C13883 VPWR.n2106 VGND 0.01325f
C13884 VPWR.n2107 VGND 0.10257f
C13885 VPWR.n2108 VGND 0.06156f
C13886 VPWR.n2109 VGND 0.74411f
C13887 VPWR.n2110 VGND 0.1428f
C13888 VPWR.n2111 VGND 0.06156f
C13889 VPWR.n2112 VGND 0.06156f
C13890 VPWR.n2113 VGND 0.06156f
C13891 VPWR.n2114 VGND 0.06156f
C13892 VPWR.n2115 VGND 0.06156f
C13893 VPWR.n2116 VGND 0.06156f
C13894 VPWR.n2117 VGND 0.06156f
C13895 VPWR.n2118 VGND 0.06156f
C13896 VPWR.n2119 VGND 0.06156f
C13897 VPWR.n2120 VGND 0.06156f
C13898 VPWR.n2121 VGND 0.06156f
C13899 VPWR.n2122 VGND 0.06156f
C13900 VPWR.n2123 VGND 0.06156f
C13901 VPWR.n2124 VGND 0.06156f
C13902 VPWR.n2125 VGND 0.06156f
C13903 VPWR.n2126 VGND 0.74411f
C13904 VPWR.n2127 VGND 0.74411f
C13905 VPWR.n2128 VGND 0.06156f
C13906 VPWR.n2129 VGND 0.10257f
C13907 VPWR.n2130 VGND 0.01325f
C13908 VPWR.n2132 VGND 0.07978f
C13909 VPWR.t70 VGND 0.08814f
C13910 VPWR.t1257 VGND 0.05786f
C13911 VPWR.t1157 VGND 0.06796f
C13912 VPWR.t603 VGND 0.05786f
C13913 VPWR.t1151 VGND 0.08814f
C13914 VPWR.n2133 VGND 0.07978f
C13915 VPWR.n2135 VGND 0.01325f
C13916 VPWR.n2136 VGND 0.10257f
C13917 VPWR.n2137 VGND 0.06156f
C13918 VPWR.n2138 VGND 0.06156f
C13919 VPWR.n2139 VGND 0.10257f
C13920 VPWR.n2140 VGND 0.01325f
C13921 VPWR.n2142 VGND 0.07978f
C13922 VPWR.t1081 VGND 0.08814f
C13923 VPWR.t497 VGND 0.05786f
C13924 VPWR.t751 VGND 0.06796f
C13925 VPWR.t701 VGND 0.05786f
C13926 VPWR.t417 VGND 0.08814f
C13927 VPWR.n2143 VGND 0.07978f
C13928 VPWR.n2145 VGND 0.01325f
C13929 VPWR.n2146 VGND 0.10257f
C13930 VPWR.n2147 VGND 0.06156f
C13931 VPWR.n2148 VGND 0.06156f
C13932 VPWR.n2149 VGND 0.10257f
C13933 VPWR.n2150 VGND 0.01325f
C13934 VPWR.n2152 VGND 0.07978f
C13935 VPWR.t1323 VGND 0.08814f
C13936 VPWR.t1141 VGND 0.05786f
C13937 VPWR.t843 VGND 0.06796f
C13938 VPWR.t1140 VGND 0.05786f
C13939 VPWR.t1099 VGND 0.08814f
C13940 VPWR.n2153 VGND 0.07978f
C13941 VPWR.n2155 VGND 0.01325f
C13942 VPWR.n2156 VGND 0.10257f
C13943 VPWR.n2157 VGND 0.06156f
C13944 VPWR.n2158 VGND 0.06156f
C13945 VPWR.n2159 VGND 0.10257f
C13946 VPWR.n2160 VGND 0.01325f
C13947 VPWR.n2162 VGND 0.07978f
C13948 VPWR.t1899 VGND 0.08814f
C13949 VPWR.t700 VGND 0.05786f
C13950 VPWR.t240 VGND 0.06796f
C13951 VPWR.t699 VGND 0.05786f
C13952 VPWR.t222 VGND 0.08814f
C13953 VPWR.n2163 VGND 0.07978f
C13954 VPWR.n2165 VGND 0.01325f
C13955 VPWR.n2166 VGND 0.10257f
C13956 VPWR.n2167 VGND 0.06156f
C13957 VPWR.n2168 VGND 0.06156f
C13958 VPWR.n2169 VGND 0.10257f
C13959 VPWR.n2170 VGND 0.01325f
C13960 VPWR.n2172 VGND 0.07978f
C13961 VPWR.t794 VGND 0.08814f
C13962 VPWR.t1142 VGND 0.05786f
C13963 VPWR.t352 VGND 0.06796f
C13964 VPWR.t496 VGND 0.05786f
C13965 VPWR.t346 VGND 0.08814f
C13966 VPWR.n2173 VGND 0.07978f
C13967 VPWR.n2175 VGND 0.01325f
C13968 VPWR.n2176 VGND 0.10257f
C13969 VPWR.n2177 VGND 0.06156f
C13970 VPWR.n2178 VGND 0.06156f
C13971 VPWR.n2179 VGND 0.10257f
C13972 VPWR.n2180 VGND 0.01325f
C13973 VPWR.n2182 VGND 0.07978f
C13974 VPWR.t1409 VGND 0.08814f
C13975 VPWR.t495 VGND 0.05786f
C13976 VPWR.t1809 VGND 0.06796f
C13977 VPWR.t1139 VGND 0.05786f
C13978 VPWR.t1163 VGND 0.08814f
C13979 VPWR.n2183 VGND 0.07978f
C13980 VPWR.n2185 VGND 0.01325f
C13981 VPWR.n2186 VGND 0.10257f
C13982 VPWR.n2187 VGND 0.06156f
C13983 VPWR.n2188 VGND 0.06156f
C13984 VPWR.n2189 VGND 0.10257f
C13985 VPWR.n2190 VGND 0.01325f
C13986 VPWR.n2192 VGND 0.07978f
C13987 VPWR.t254 VGND 0.08814f
C13988 VPWR.t1138 VGND 0.05786f
C13989 VPWR.t1195 VGND 0.06796f
C13990 VPWR.t604 VGND 0.05786f
C13991 VPWR.t999 VGND 0.08814f
C13992 VPWR.n2193 VGND 0.07978f
C13993 VPWR.n2195 VGND 0.01325f
C13994 VPWR.n2196 VGND 0.10257f
C13995 VPWR.n2197 VGND 0.06156f
C13996 VPWR.n2198 VGND 0.06156f
C13997 VPWR.n2199 VGND 0.10257f
C13998 VPWR.n2200 VGND 0.01325f
C13999 VPWR.n2202 VGND 0.07978f
C14000 VPWR.t16 VGND 0.08814f
C14001 VPWR.t1258 VGND 0.05786f
C14002 VPWR.t1462 VGND 0.09829f
C14003 VPWR.n2203 VGND 0.05616f
C14004 VPWR.n2204 VGND 0.01325f
C14005 VPWR.n2205 VGND 0.10257f
C14006 VPWR.n2206 VGND 0.1428f
C14007 VPWR.n2207 VGND 0.7488f
C14008 VPWR.n2208 VGND 0.06156f
C14009 VPWR.n2209 VGND 0.06156f
C14010 VPWR.n2210 VGND 0.06156f
C14011 VPWR.n2211 VGND 0.06156f
C14012 VPWR.n2212 VGND 0.06156f
C14013 VPWR.n2213 VGND 0.06156f
C14014 VPWR.n2214 VGND 0.06156f
C14015 VPWR.n2215 VGND 0.06156f
C14016 VPWR.n2216 VGND 0.06156f
C14017 VPWR.n2217 VGND 0.06156f
C14018 VPWR.n2218 VGND 0.06156f
C14019 VPWR.n2219 VGND 0.06156f
C14020 VPWR.n2220 VGND 0.06156f
C14021 VPWR.n2221 VGND 0.06156f
C14022 VPWR.n2222 VGND 0.06156f
C14023 VPWR.n2223 VGND 0.1428f
C14024 VPWR.n2224 VGND 0.7488f
C14025 VPWR.n2225 VGND 0.7488f
C14026 VPWR.n2226 VGND 0.1428f
C14027 VPWR.n2227 VGND 0.10257f
C14028 VPWR.n2228 VGND 0.01325f
C14029 VPWR.n2229 VGND 0.05616f
C14030 VPWR.t1628 VGND 0.09829f
C14031 VPWR.t1349 VGND 0.05786f
C14032 VPWR.t1233 VGND 0.08814f
C14033 VPWR.n2230 VGND 0.07978f
C14034 VPWR.n2232 VGND 0.01325f
C14035 VPWR.n2233 VGND 0.10257f
C14036 VPWR.n2234 VGND 0.06156f
C14037 VPWR.n2235 VGND 0.06156f
C14038 VPWR.n2236 VGND 0.10257f
C14039 VPWR.n2237 VGND 0.01325f
C14040 VPWR.n2239 VGND 0.07978f
C14041 VPWR.t640 VGND 0.06796f
C14042 VPWR.t1340 VGND 0.05786f
C14043 VPWR.t179 VGND 0.08814f
C14044 VPWR.n2240 VGND 0.07978f
C14045 VPWR.n2242 VGND 0.01325f
C14046 VPWR.n2243 VGND 0.10257f
C14047 VPWR.n2244 VGND 0.06156f
C14048 VPWR.n2245 VGND 0.06156f
C14049 VPWR.n2246 VGND 0.10257f
C14050 VPWR.n2247 VGND 0.01325f
C14051 VPWR.n2249 VGND 0.07978f
C14052 VPWR.t1863 VGND 0.06796f
C14053 VPWR.t866 VGND 0.05786f
C14054 VPWR.t780 VGND 0.08814f
C14055 VPWR.n2250 VGND 0.07978f
C14056 VPWR.n2252 VGND 0.01325f
C14057 VPWR.n2253 VGND 0.10257f
C14058 VPWR.n2254 VGND 0.06156f
C14059 VPWR.n2255 VGND 0.06156f
C14060 VPWR.n2256 VGND 0.10257f
C14061 VPWR.n2257 VGND 0.01325f
C14062 VPWR.n2259 VGND 0.07978f
C14063 VPWR.t330 VGND 0.06796f
C14064 VPWR.t1344 VGND 0.05786f
C14065 VPWR.t46 VGND 0.08814f
C14066 VPWR.n2260 VGND 0.07978f
C14067 VPWR.n2262 VGND 0.01325f
C14068 VPWR.n2263 VGND 0.10257f
C14069 VPWR.n2264 VGND 0.06156f
C14070 VPWR.n2265 VGND 0.06156f
C14071 VPWR.n2266 VGND 0.10257f
C14072 VPWR.n2267 VGND 0.01325f
C14073 VPWR.n2269 VGND 0.07978f
C14074 VPWR.t218 VGND 0.06796f
C14075 VPWR.t1351 VGND 0.05786f
C14076 VPWR.t714 VGND 0.08814f
C14077 VPWR.n2270 VGND 0.07978f
C14078 VPWR.n2272 VGND 0.01325f
C14079 VPWR.n2273 VGND 0.10257f
C14080 VPWR.n2274 VGND 0.06156f
C14081 VPWR.n2275 VGND 0.06156f
C14082 VPWR.n2276 VGND 0.10257f
C14083 VPWR.n2277 VGND 0.01325f
C14084 VPWR.n2279 VGND 0.07978f
C14085 VPWR.t60 VGND 0.06796f
C14086 VPWR.t1343 VGND 0.05786f
C14087 VPWR.t144 VGND 0.08814f
C14088 VPWR.n2280 VGND 0.07978f
C14089 VPWR.n2282 VGND 0.01325f
C14090 VPWR.n2283 VGND 0.10257f
C14091 VPWR.n2284 VGND 0.06156f
C14092 VPWR.n2285 VGND 0.06156f
C14093 VPWR.n2286 VGND 0.10257f
C14094 VPWR.n2287 VGND 0.01325f
C14095 VPWR.n2289 VGND 0.07978f
C14096 VPWR.t413 VGND 0.06796f
C14097 VPWR.t868 VGND 0.05786f
C14098 VPWR.t1047 VGND 0.08814f
C14099 VPWR.n2290 VGND 0.07978f
C14100 VPWR.n2292 VGND 0.01325f
C14101 VPWR.n2293 VGND 0.10257f
C14102 VPWR.n2294 VGND 0.06156f
C14103 VPWR.n2295 VGND 0.06156f
C14104 VPWR.n2296 VGND 0.10257f
C14105 VPWR.n2297 VGND 0.01325f
C14106 VPWR.n2299 VGND 0.07978f
C14107 VPWR.t516 VGND 0.06796f
C14108 VPWR.t1345 VGND 0.05786f
C14109 VPWR.t735 VGND 0.08814f
C14110 VPWR.n2300 VGND 0.07978f
C14111 VPWR.n2302 VGND 0.01325f
C14112 VPWR.n2303 VGND 0.10257f
C14113 VPWR.n2304 VGND 0.06156f
C14114 VPWR.n2305 VGND 0.74411f
C14115 VPWR.n2306 VGND 0.1428f
C14116 VPWR.n2307 VGND 0.06156f
C14117 VPWR.n2308 VGND 0.06156f
C14118 VPWR.n2309 VGND 0.06156f
C14119 VPWR.n2310 VGND 0.06156f
C14120 VPWR.n2311 VGND 0.06156f
C14121 VPWR.n2312 VGND 0.06156f
C14122 VPWR.n2313 VGND 0.06156f
C14123 VPWR.n2314 VGND 0.06156f
C14124 VPWR.n2315 VGND 0.06156f
C14125 VPWR.n2316 VGND 0.06156f
C14126 VPWR.n2317 VGND 0.06156f
C14127 VPWR.n2318 VGND 0.06156f
C14128 VPWR.n2319 VGND 0.06156f
C14129 VPWR.n2320 VGND 0.06156f
C14130 VPWR.n2321 VGND 0.06156f
C14131 VPWR.n2322 VGND 0.74411f
C14132 VPWR.n2323 VGND 0.74411f
C14133 VPWR.n2324 VGND 0.06156f
C14134 VPWR.n2325 VGND 0.10257f
C14135 VPWR.n2326 VGND 0.01325f
C14136 VPWR.n2328 VGND 0.07978f
C14137 VPWR.t498 VGND 0.08814f
C14138 VPWR.t1321 VGND 0.05786f
C14139 VPWR.t504 VGND 0.06796f
C14140 VPWR.t770 VGND 0.05786f
C14141 VPWR.t1918 VGND 0.08814f
C14142 VPWR.n2329 VGND 0.07978f
C14143 VPWR.n2331 VGND 0.01325f
C14144 VPWR.n2332 VGND 0.10257f
C14145 VPWR.n2333 VGND 0.06156f
C14146 VPWR.n2334 VGND 0.06156f
C14147 VPWR.n2335 VGND 0.10257f
C14148 VPWR.n2336 VGND 0.01325f
C14149 VPWR.n2338 VGND 0.07978f
C14150 VPWR.t1093 VGND 0.08814f
C14151 VPWR.t141 VGND 0.05786f
C14152 VPWR.t691 VGND 0.06796f
C14153 VPWR.t1838 VGND 0.05786f
C14154 VPWR.t405 VGND 0.08814f
C14155 VPWR.n2339 VGND 0.07978f
C14156 VPWR.n2341 VGND 0.01325f
C14157 VPWR.n2342 VGND 0.10257f
C14158 VPWR.n2343 VGND 0.06156f
C14159 VPWR.n2344 VGND 0.06156f
C14160 VPWR.n2345 VGND 0.10257f
C14161 VPWR.n2346 VGND 0.01325f
C14162 VPWR.n2348 VGND 0.07978f
C14163 VPWR.t1263 VGND 0.08814f
C14164 VPWR.t775 VGND 0.05786f
C14165 VPWR.t862 VGND 0.06796f
C14166 VPWR.t774 VGND 0.05786f
C14167 VPWR.t858 VGND 0.08814f
C14168 VPWR.n2349 VGND 0.07978f
C14169 VPWR.n2351 VGND 0.01325f
C14170 VPWR.n2352 VGND 0.10257f
C14171 VPWR.n2353 VGND 0.06156f
C14172 VPWR.n2354 VGND 0.06156f
C14173 VPWR.n2355 VGND 0.10257f
C14174 VPWR.n2356 VGND 0.01325f
C14175 VPWR.n2358 VGND 0.07978f
C14176 VPWR.t454 VGND 0.08814f
C14177 VPWR.t1837 VGND 0.05786f
C14178 VPWR.t1929 VGND 0.06796f
C14179 VPWR.t650 VGND 0.05786f
C14180 VPWR.t952 VGND 0.08814f
C14181 VPWR.n2359 VGND 0.07978f
C14182 VPWR.n2361 VGND 0.01325f
C14183 VPWR.n2362 VGND 0.10257f
C14184 VPWR.n2363 VGND 0.06156f
C14185 VPWR.n2364 VGND 0.06156f
C14186 VPWR.n2365 VGND 0.10257f
C14187 VPWR.n2366 VGND 0.01325f
C14188 VPWR.n2368 VGND 0.07978f
C14189 VPWR.t653 VGND 0.08814f
C14190 VPWR.t1320 VGND 0.05786f
C14191 VPWR.t342 VGND 0.06796f
C14192 VPWR.t140 VGND 0.05786f
C14193 VPWR.t334 VGND 0.08814f
C14194 VPWR.n2369 VGND 0.07978f
C14195 VPWR.n2371 VGND 0.01325f
C14196 VPWR.n2372 VGND 0.10257f
C14197 VPWR.n2373 VGND 0.06156f
C14198 VPWR.n2374 VGND 0.06156f
C14199 VPWR.n2375 VGND 0.10257f
C14200 VPWR.n2376 VGND 0.01325f
C14201 VPWR.n2378 VGND 0.07978f
C14202 VPWR.t1201 VGND 0.08814f
C14203 VPWR.t139 VGND 0.05786f
C14204 VPWR.t1021 VGND 0.06796f
C14205 VPWR.t773 VGND 0.05786f
C14206 VPWR.t1867 VGND 0.08814f
C14207 VPWR.n2379 VGND 0.07978f
C14208 VPWR.n2381 VGND 0.01325f
C14209 VPWR.n2382 VGND 0.10257f
C14210 VPWR.n2383 VGND 0.06156f
C14211 VPWR.n2384 VGND 0.06156f
C14212 VPWR.n2385 VGND 0.10257f
C14213 VPWR.n2386 VGND 0.01325f
C14214 VPWR.n2388 VGND 0.07978f
C14215 VPWR.t193 VGND 0.08814f
C14216 VPWR.t772 VGND 0.05786f
C14217 VPWR.t1013 VGND 0.06796f
C14218 VPWR.t771 VGND 0.05786f
C14219 VPWR.t1005 VGND 0.08814f
C14220 VPWR.n2389 VGND 0.07978f
C14221 VPWR.n2391 VGND 0.01325f
C14222 VPWR.n2392 VGND 0.10257f
C14223 VPWR.n2393 VGND 0.06156f
C14224 VPWR.n2394 VGND 0.06156f
C14225 VPWR.n2395 VGND 0.10257f
C14226 VPWR.n2396 VGND 0.01325f
C14227 VPWR.n2398 VGND 0.07978f
C14228 VPWR.t20 VGND 0.08814f
C14229 VPWR.t1322 VGND 0.05786f
C14230 VPWR.t1561 VGND 0.09829f
C14231 VPWR.n2399 VGND 0.05616f
C14232 VPWR.n2400 VGND 0.01325f
C14233 VPWR.n2401 VGND 0.10257f
C14234 VPWR.n2402 VGND 0.1428f
C14235 VPWR.n2403 VGND 0.7488f
C14236 VPWR.n2404 VGND 0.06156f
C14237 VPWR.n2405 VGND 0.06156f
C14238 VPWR.n2406 VGND 0.06156f
C14239 VPWR.n2407 VGND 0.06156f
C14240 VPWR.n2408 VGND 0.06156f
C14241 VPWR.n2409 VGND 0.06156f
C14242 VPWR.n2410 VGND 0.06156f
C14243 VPWR.n2411 VGND 0.06156f
C14244 VPWR.n2412 VGND 0.06156f
C14245 VPWR.n2413 VGND 0.06156f
C14246 VPWR.n2414 VGND 0.06156f
C14247 VPWR.n2415 VGND 0.06156f
C14248 VPWR.n2416 VGND 0.06156f
C14249 VPWR.n2417 VGND 0.06156f
C14250 VPWR.n2418 VGND 0.06156f
C14251 VPWR.n2419 VGND 0.1428f
C14252 VPWR.n2420 VGND 0.7488f
C14253 VPWR.n2421 VGND 0.7488f
C14254 VPWR.n2422 VGND 0.1428f
C14255 VPWR.n2423 VGND 0.10257f
C14256 VPWR.n2424 VGND 0.01325f
C14257 VPWR.n2425 VGND 0.05616f
C14258 VPWR.t1734 VGND 0.09829f
C14259 VPWR.t1365 VGND 0.05786f
C14260 VPWR.t827 VGND 0.08814f
C14261 VPWR.n2426 VGND 0.07978f
C14262 VPWR.n2428 VGND 0.01325f
C14263 VPWR.n2429 VGND 0.10257f
C14264 VPWR.n2430 VGND 0.06156f
C14265 VPWR.n2431 VGND 0.06156f
C14266 VPWR.n2432 VGND 0.10257f
C14267 VPWR.n2433 VGND 0.01325f
C14268 VPWR.n2435 VGND 0.07978f
C14269 VPWR.t979 VGND 0.06796f
C14270 VPWR.t885 VGND 0.05786f
C14271 VPWR.t1314 VGND 0.08814f
C14272 VPWR.n2436 VGND 0.07978f
C14273 VPWR.n2438 VGND 0.01325f
C14274 VPWR.n2439 VGND 0.10257f
C14275 VPWR.n2440 VGND 0.06156f
C14276 VPWR.n2441 VGND 0.06156f
C14277 VPWR.n2442 VGND 0.10257f
C14278 VPWR.n2443 VGND 0.01325f
C14279 VPWR.n2445 VGND 0.07978f
C14280 VPWR.t1884 VGND 0.06796f
C14281 VPWR.t1207 VGND 0.05786f
C14282 VPWR.t488 VGND 0.08814f
C14283 VPWR.n2446 VGND 0.07978f
C14284 VPWR.n2448 VGND 0.01325f
C14285 VPWR.n2449 VGND 0.10257f
C14286 VPWR.n2450 VGND 0.06156f
C14287 VPWR.n2451 VGND 0.06156f
C14288 VPWR.n2452 VGND 0.10257f
C14289 VPWR.n2453 VGND 0.01325f
C14290 VPWR.n2455 VGND 0.07978f
C14291 VPWR.t366 VGND 0.06796f
C14292 VPWR.t1363 VGND 0.05786f
C14293 VPWR.t1283 VGND 0.08814f
C14294 VPWR.n2456 VGND 0.07978f
C14295 VPWR.n2458 VGND 0.01325f
C14296 VPWR.n2459 VGND 0.10257f
C14297 VPWR.n2460 VGND 0.06156f
C14298 VPWR.n2461 VGND 0.06156f
C14299 VPWR.n2462 VGND 0.10257f
C14300 VPWR.n2463 VGND 0.01325f
C14301 VPWR.n2465 VGND 0.07978f
C14302 VPWR.t938 VGND 0.06796f
C14303 VPWR.t1360 VGND 0.05786f
C14304 VPWR.t1386 VGND 0.08814f
C14305 VPWR.n2466 VGND 0.07978f
C14306 VPWR.n2468 VGND 0.01325f
C14307 VPWR.n2469 VGND 0.10257f
C14308 VPWR.n2470 VGND 0.06156f
C14309 VPWR.n2471 VGND 0.06156f
C14310 VPWR.n2472 VGND 0.10257f
C14311 VPWR.n2473 VGND 0.01325f
C14312 VPWR.n2475 VGND 0.07978f
C14313 VPWR.t1801 VGND 0.06796f
C14314 VPWR.t888 VGND 0.05786f
C14315 VPWR.t905 VGND 0.08814f
C14316 VPWR.n2476 VGND 0.07978f
C14317 VPWR.n2478 VGND 0.01325f
C14318 VPWR.n2479 VGND 0.10257f
C14319 VPWR.n2480 VGND 0.06156f
C14320 VPWR.n2481 VGND 0.06156f
C14321 VPWR.n2482 VGND 0.10257f
C14322 VPWR.n2483 VGND 0.01325f
C14323 VPWR.n2485 VGND 0.07978f
C14324 VPWR.t1396 VGND 0.06796f
C14325 VPWR.t1209 VGND 0.05786f
C14326 VPWR.t1059 VGND 0.08814f
C14327 VPWR.n2486 VGND 0.07978f
C14328 VPWR.n2488 VGND 0.01325f
C14329 VPWR.n2489 VGND 0.10257f
C14330 VPWR.n2490 VGND 0.06156f
C14331 VPWR.n2491 VGND 0.06156f
C14332 VPWR.n2492 VGND 0.10257f
C14333 VPWR.n2493 VGND 0.01325f
C14334 VPWR.n2495 VGND 0.07978f
C14335 VPWR.t1334 VGND 0.06796f
C14336 VPWR.t1364 VGND 0.05786f
C14337 VPWR.t784 VGND 0.08814f
C14338 VPWR.n2496 VGND 0.07978f
C14339 VPWR.n2498 VGND 0.01325f
C14340 VPWR.n2499 VGND 0.10257f
C14341 VPWR.n2500 VGND 0.06156f
C14342 VPWR.n2501 VGND 0.74411f
C14343 VPWR.n2502 VGND 0.1428f
C14344 VPWR.n2503 VGND 0.06156f
C14345 VPWR.n2504 VGND 0.06156f
C14346 VPWR.n2505 VGND 0.06156f
C14347 VPWR.n2506 VGND 0.06156f
C14348 VPWR.n2507 VGND 0.06156f
C14349 VPWR.n2508 VGND 0.06156f
C14350 VPWR.n2509 VGND 0.06156f
C14351 VPWR.n2510 VGND 0.06156f
C14352 VPWR.n2511 VGND 0.06156f
C14353 VPWR.n2512 VGND 0.06156f
C14354 VPWR.n2513 VGND 0.06156f
C14355 VPWR.n2514 VGND 0.06156f
C14356 VPWR.n2515 VGND 0.06156f
C14357 VPWR.n2516 VGND 0.06156f
C14358 VPWR.n2517 VGND 0.06156f
C14359 VPWR.n2518 VGND 0.74411f
C14360 VPWR.n2519 VGND 0.42115f
C14361 VPWR.n2520 VGND 0.06156f
C14362 VPWR.n2521 VGND 0.06379f
C14363 VPWR.n2523 VGND 0.01264f
C14364 VPWR.n2525 VGND 0.07978f
C14365 VPWR.t1610 VGND 0.08814f
C14366 VPWR.t1577 VGND 0.05786f
C14367 VPWR.t1707 VGND 0.06796f
C14368 VPWR.t1713 VGND 0.05786f
C14369 VPWR.t1725 VGND 0.08814f
C14370 VPWR.n2526 VGND 0.07978f
C14371 VPWR.n2528 VGND 0.01264f
C14372 VPWR.n2530 VGND 0.06379f
C14373 VPWR.n2531 VGND 0.06156f
C14374 VPWR.n2532 VGND 0.06156f
C14375 VPWR.n2533 VGND 0.06379f
C14376 VPWR.n2535 VGND 0.01264f
C14377 VPWR.n2537 VGND 0.07978f
C14378 VPWR.t1487 VGND 0.08814f
C14379 VPWR.t1747 VGND 0.05786f
C14380 VPWR.t1481 VGND 0.06796f
C14381 VPWR.t1471 VGND 0.05786f
C14382 VPWR.t1595 VGND 0.08814f
C14383 VPWR.n2538 VGND 0.07978f
C14384 VPWR.n2540 VGND 0.01264f
C14385 VPWR.n2542 VGND 0.06379f
C14386 VPWR.n2543 VGND 0.06156f
C14387 VPWR.n2544 VGND 0.06156f
C14388 VPWR.n2545 VGND 0.06379f
C14389 VPWR.n2547 VGND 0.01264f
C14390 VPWR.n2549 VGND 0.07978f
C14391 VPWR.t1607 VGND 0.08814f
C14392 VPWR.t1615 VGND 0.05786f
C14393 VPWR.t1744 VGND 0.06796f
C14394 VPWR.t1639 VGND 0.05786f
C14395 VPWR.t1763 VGND 0.08814f
C14396 VPWR.n2550 VGND 0.07978f
C14397 VPWR.n2552 VGND 0.01264f
C14398 VPWR.n2554 VGND 0.06379f
C14399 VPWR.n2555 VGND 0.06156f
C14400 VPWR.n2556 VGND 0.06156f
C14401 VPWR.n2557 VGND 0.06379f
C14402 VPWR.n2559 VGND 0.01264f
C14403 VPWR.n2561 VGND 0.07978f
C14404 VPWR.t1484 VGND 0.08814f
C14405 VPWR.t1476 VGND 0.05786f
C14406 VPWR.t1503 VGND 0.06796f
C14407 VPWR.t1511 VGND 0.05786f
C14408 VPWR.t1644 VGND 0.08814f
C14409 VPWR.n2562 VGND 0.07978f
C14410 VPWR.n2564 VGND 0.01264f
C14411 VPWR.n2566 VGND 0.06379f
C14412 VPWR.n2567 VGND 0.06156f
C14413 VPWR.n2568 VGND 0.06156f
C14414 VPWR.n2569 VGND 0.06379f
C14415 VPWR.n2571 VGND 0.01264f
C14416 VPWR.n2573 VGND 0.07978f
C14417 VPWR.t1660 VGND 0.08814f
C14418 VPWR.t1613 VGND 0.05786f
C14419 VPWR.t1696 VGND 0.06796f
C14420 VPWR.t1774 VGND 0.05786f
C14421 VPWR.t1790 VGND 0.08814f
C14422 VPWR.n2574 VGND 0.07978f
C14423 VPWR.n2576 VGND 0.01264f
C14424 VPWR.n2578 VGND 0.06379f
C14425 VPWR.n2579 VGND 0.06156f
C14426 VPWR.n2580 VGND 0.06156f
C14427 VPWR.n2581 VGND 0.06379f
C14428 VPWR.n2583 VGND 0.01264f
C14429 VPWR.n2585 VGND 0.07978f
C14430 VPWR.t1534 VGND 0.08814f
C14431 VPWR.t1793 VGND 0.05786f
C14432 VPWR.t1526 VGND 0.06796f
C14433 VPWR.t1647 VGND 0.05786f
C14434 VPWR.t1564 VGND 0.08814f
C14435 VPWR.n2586 VGND 0.07978f
C14436 VPWR.n2588 VGND 0.01264f
C14437 VPWR.n2590 VGND 0.06379f
C14438 VPWR.n2591 VGND 0.06156f
C14439 VPWR.n2592 VGND 0.06156f
C14440 VPWR.n2593 VGND 0.06379f
C14441 VPWR.n2595 VGND 0.01264f
C14442 VPWR.n2597 VGND 0.07978f
C14443 VPWR.t1414 VGND 0.08814f
C14444 VPWR.t1669 VGND 0.05786f
C14445 VPWR.t1787 VGND 0.06796f
C14446 VPWR.t1691 VGND 0.05786f
C14447 VPWR.t1433 VGND 0.08814f
C14448 VPWR.n2598 VGND 0.07978f
C14449 VPWR.n2600 VGND 0.01264f
C14450 VPWR.n2602 VGND 0.06379f
C14451 VPWR.n2603 VGND 0.06156f
C14452 VPWR.n2604 VGND 0.06156f
C14453 VPWR.n2605 VGND 0.06379f
C14454 VPWR.n2607 VGND 0.01264f
C14455 VPWR.n2609 VGND 0.07978f
C14456 VPWR.t1558 VGND 0.08814f
C14457 VPWR.t1542 VGND 0.05786f
C14458 VPWR.t1663 VGND 0.09829f
C14459 VPWR.n2610 VGND 0.05613f
C14460 VPWR.n2611 VGND 0.01252f
C14461 VPWR.n2613 VGND 0.08001f
C14462 VPWR.n2614 VGND 0.1428f
C14463 VPWR.n2615 VGND 1.96285f
C14464 VPWR.n2616 VGND 0.79936f
C14465 VPWR.n2617 VGND 0.33493f
C14466 VPWR.t123 VGND 0.04022f
C14467 VPWR.t942 VGND 0.04022f
C14468 VPWR.n2618 VGND 0.07296f
C14469 VPWR.n2619 VGND 0.03455f
C14470 VPWR.t121 VGND 0.01056f
C14471 VPWR.t129 VGND 0.01056f
C14472 VPWR.n2620 VGND 0.02267f
C14473 VPWR.t947 VGND 0.01056f
C14474 VPWR.t941 VGND 0.01056f
C14475 VPWR.n2621 VGND 0.02267f
C14476 VPWR.n2623 VGND 0.03455f
C14477 VPWR.t697 VGND 0.01056f
C14478 VPWR.t426 VGND 0.01056f
C14479 VPWR.n2624 VGND 0.02267f
C14480 VPWR.t315 VGND 0.01056f
C14481 VPWR.t307 VGND 0.01056f
C14482 VPWR.n2625 VGND 0.02267f
C14483 VPWR.t199 VGND 0.04212f
C14484 VPWR.t274 VGND 0.04212f
C14485 VPWR.n2626 VGND 0.09713f
C14486 VPWR.n2627 VGND 0.03117f
C14487 VPWR.n2628 VGND 0.01004f
C14488 VPWR.n2629 VGND 0.04558f
C14489 VPWR.t273 VGND 0.01056f
C14490 VPWR.t127 VGND 0.01056f
C14491 VPWR.n2631 VGND 0.02267f
C14492 VPWR.t201 VGND 0.01056f
C14493 VPWR.t945 VGND 0.01056f
C14494 VPWR.n2632 VGND 0.02267f
C14495 VPWR.n2633 VGND 0.04558f
C14496 VPWR.n2634 VGND 0.01051f
C14497 VPWR.n2635 VGND 0.03455f
C14498 VPWR.n2636 VGND 0.03455f
C14499 VPWR.n2637 VGND 0.03455f
C14500 VPWR.n2639 VGND 0.04558f
C14501 VPWR.n2642 VGND 0.03455f
C14502 VPWR.n2643 VGND 0.02591f
C14503 VPWR.t198 VGND 0.1262f
C14504 VPWR.t314 VGND 0.18598f
C14505 VPWR.t306 VGND 0.18598f
C14506 VPWR.t200 VGND 0.18598f
C14507 VPWR.t126 VGND 0.18598f
C14508 VPWR.t120 VGND 0.18598f
C14509 VPWR.t128 VGND 0.18598f
C14510 VPWR.t122 VGND 0.41406f
C14511 VPWR.n2645 VGND 0.45194f
C14512 VPWR.n2646 VGND 0.01314f
C14513 VPWR.n2647 VGND 0.7927f
C14514 VPWR.n2648 VGND 0.03455f
C14515 VPWR.t275 VGND 0.1262f
C14516 VPWR.t310 VGND 0.18598f
C14517 VPWR.t271 VGND 0.18598f
C14518 VPWR.t376 VGND 0.18598f
C14519 VPWR.t76 VGND 0.18598f
C14520 VPWR.t86 VGND 0.18598f
C14521 VPWR.t78 VGND 0.18598f
C14522 VPWR.t88 VGND 0.30554f
C14523 VPWR.t168 VGND 0.32436f
C14524 VPWR.n2649 VGND 0.45773f
C14525 VPWR.n2650 VGND 0.13021f
C14526 VPWR.n2651 VGND 0.03455f
C14527 VPWR.t87 VGND 0.01056f
C14528 VPWR.t79 VGND 0.01056f
C14529 VPWR.n2652 VGND 0.02267f
C14530 VPWR.t1892 VGND 0.01056f
C14531 VPWR.t1898 VGND 0.01056f
C14532 VPWR.n2653 VGND 0.02267f
C14533 VPWR.n2654 VGND 0.04558f
C14534 VPWR.n2655 VGND 0.03455f
C14535 VPWR.t694 VGND 0.01056f
C14536 VPWR.t77 VGND 0.01056f
C14537 VPWR.n2656 VGND 0.02267f
C14538 VPWR.t377 VGND 0.01056f
C14539 VPWR.t1896 VGND 0.01056f
C14540 VPWR.n2657 VGND 0.02267f
C14541 VPWR.t276 VGND 0.04212f
C14542 VPWR.t695 VGND 0.04212f
C14543 VPWR.n2659 VGND 0.09713f
C14544 VPWR.t423 VGND 0.01056f
C14545 VPWR.t272 VGND 0.01056f
C14546 VPWR.n2660 VGND 0.02267f
C14547 VPWR.t311 VGND 0.01056f
C14548 VPWR.t1858 VGND 0.01056f
C14549 VPWR.n2661 VGND 0.02267f
C14550 VPWR.n2662 VGND 0.04558f
C14551 VPWR.n2663 VGND 0.01004f
C14552 VPWR.n2664 VGND 0.03117f
C14553 VPWR.n2665 VGND 0.03455f
C14554 VPWR.n2666 VGND 0.03455f
C14555 VPWR.n2667 VGND 0.01051f
C14556 VPWR.n2668 VGND 0.04558f
C14557 VPWR.n2671 VGND 0.03455f
C14558 VPWR.n2672 VGND 0.03455f
C14559 VPWR.t89 VGND 0.04022f
C14560 VPWR.t1894 VGND 0.04022f
C14561 VPWR.n2675 VGND 0.07296f
C14562 VPWR.n2677 VGND 0.02591f
C14563 VPWR.n2678 VGND 0.01314f
C14564 VPWR.n2679 VGND 0.02591f
C14565 VPWR.n2680 VGND 0.01031f
C14566 VPWR.t169 VGND 0.04208f
C14567 VPWR.t1798 VGND 0.04208f
C14568 VPWR.n2682 VGND 0.08505f
C14569 VPWR.n2683 VGND 0.02404f
C14570 VPWR.n2684 VGND 1.20645f
C14571 VPWR.n2685 VGND 0.03455f
C14572 VPWR.t155 VGND 0.0413f
C14573 VPWR.t419 VGND 0.1262f
C14574 VPWR.t312 VGND 0.18598f
C14575 VPWR.t374 VGND 0.18598f
C14576 VPWR.t205 VGND 0.18598f
C14577 VPWR.t657 VGND 0.18598f
C14578 VPWR.t1168 VGND 0.18598f
C14579 VPWR.t1174 VGND 0.18598f
C14580 VPWR.t1170 VGND 0.30554f
C14581 VPWR.t92 VGND 0.11735f
C14582 VPWR.t154 VGND 0.09299f
C14583 VPWR.t1108 VGND 0.20702f
C14584 VPWR.n2686 VGND 0.4057f
C14585 VPWR.n2687 VGND 0.12828f
C14586 VPWR.n2688 VGND 0.03455f
C14587 VPWR.t1169 VGND 0.01056f
C14588 VPWR.t1175 VGND 0.01056f
C14589 VPWR.n2689 VGND 0.02267f
C14590 VPWR.t1923 VGND 0.01056f
C14591 VPWR.t1319 VGND 0.01056f
C14592 VPWR.n2690 VGND 0.02267f
C14593 VPWR.n2691 VGND 0.04558f
C14594 VPWR.n2692 VGND 0.03455f
C14595 VPWR.t380 VGND 0.01056f
C14596 VPWR.t1173 VGND 0.01056f
C14597 VPWR.n2693 VGND 0.02267f
C14598 VPWR.t206 VGND 0.01056f
C14599 VPWR.t658 VGND 0.01056f
C14600 VPWR.n2694 VGND 0.02267f
C14601 VPWR.t696 VGND 0.04212f
C14602 VPWR.t420 VGND 0.04212f
C14603 VPWR.n2696 VGND 0.09713f
C14604 VPWR.t313 VGND 0.01056f
C14605 VPWR.t465 VGND 0.01056f
C14606 VPWR.n2697 VGND 0.02267f
C14607 VPWR.t1856 VGND 0.01056f
C14608 VPWR.t375 VGND 0.01056f
C14609 VPWR.n2698 VGND 0.02267f
C14610 VPWR.n2699 VGND 0.04558f
C14611 VPWR.n2700 VGND 0.01004f
C14612 VPWR.n2701 VGND 0.03117f
C14613 VPWR.n2702 VGND 0.03455f
C14614 VPWR.n2703 VGND 0.03455f
C14615 VPWR.n2704 VGND 0.01051f
C14616 VPWR.n2705 VGND 0.04558f
C14617 VPWR.n2708 VGND 0.03455f
C14618 VPWR.n2709 VGND 0.03455f
C14619 VPWR.t1171 VGND 0.04022f
C14620 VPWR.t1922 VGND 0.04022f
C14621 VPWR.n2712 VGND 0.07296f
C14622 VPWR.n2714 VGND 0.02591f
C14623 VPWR.n2715 VGND 0.01314f
C14624 VPWR.n2716 VGND 0.02591f
C14625 VPWR.t1109 VGND 0.04212f
C14626 VPWR.n2717 VGND 0.0587f
C14627 VPWR.n2719 VGND 0.04296f
C14628 VPWR.t93 VGND 0.04141f
C14629 VPWR.n2720 VGND 0.05367f
C14630 VPWR.n2721 VGND 0.02047f
C14631 VPWR.n2722 VGND 1.20645f
C14632 VPWR.n2723 VGND 0.03455f
C14633 VPWR.t378 VGND 0.07157f
C14634 VPWR.t283 VGND 0.10548f
C14635 VPWR.t372 VGND 0.10254f
C14636 VPWR.t203 VGND 0.164f
C14637 VPWR.t614 VGND 0.13949f
C14638 VPWR.t195 VGND 0.09299f
C14639 VPWR.t620 VGND 0.09299f
C14640 VPWR.t280 VGND 0.09299f
C14641 VPWR.t856 VGND 0.09299f
C14642 VPWR.t424 VGND 0.09299f
C14643 VPWR.t618 VGND 0.09299f
C14644 VPWR.t466 VGND 0.12952f
C14645 VPWR.t490 VGND 0.07306f
C14646 VPWR.t737 VGND 0.07971f
C14647 VPWR.t98 VGND 0.09299f
C14648 VPWR.t739 VGND 0.1727f
C14649 VPWR.n2724 VGND 0.27839f
C14650 VPWR.n2725 VGND 0.12841f
C14651 VPWR.t740 VGND 0.04181f
C14652 VPWR.n2726 VGND 0.03455f
C14653 VPWR.t467 VGND 0.04133f
C14654 VPWR.t619 VGND 0.03979f
C14655 VPWR.t281 VGND 0.01056f
C14656 VPWR.t425 VGND 0.01056f
C14657 VPWR.n2727 VGND 0.02267f
C14658 VPWR.t621 VGND 0.01056f
C14659 VPWR.t857 VGND 0.01056f
C14660 VPWR.n2728 VGND 0.02267f
C14661 VPWR.n2729 VGND 0.02585f
C14662 VPWR.n2730 VGND 0.03455f
C14663 VPWR.t204 VGND 0.01056f
C14664 VPWR.t615 VGND 0.01056f
C14665 VPWR.n2731 VGND 0.02267f
C14666 VPWR.t379 VGND 0.04212f
C14667 VPWR.n2733 VGND 0.05308f
C14668 VPWR.t284 VGND 0.01056f
C14669 VPWR.t373 VGND 0.01056f
C14670 VPWR.n2734 VGND 0.02267f
C14671 VPWR.n2735 VGND 0.02585f
C14672 VPWR.n2736 VGND 0.01004f
C14673 VPWR.n2737 VGND 0.03117f
C14674 VPWR.n2738 VGND 0.03455f
C14675 VPWR.n2739 VGND 0.03455f
C14676 VPWR.n2740 VGND 0.01051f
C14677 VPWR.n2741 VGND 0.02525f
C14678 VPWR.t196 VGND 0.03697f
C14679 VPWR.n2742 VGND 0.02947f
C14680 VPWR.n2744 VGND 0.03455f
C14681 VPWR.n2745 VGND 0.03455f
C14682 VPWR.n2746 VGND 0.02864f
C14683 VPWR.n2748 VGND 0.03791f
C14684 VPWR.n2749 VGND 0.04995f
C14685 VPWR.n2751 VGND 0.02047f
C14686 VPWR.n2752 VGND 0.01314f
C14687 VPWR.n2753 VGND 0.02591f
C14688 VPWR.t99 VGND 0.04217f
C14689 VPWR.n2754 VGND 0.10841f
C14690 VPWR.t738 VGND 0.0421f
C14691 VPWR.n2756 VGND 0.04686f
C14692 VPWR.n2757 VGND 0.02028f
C14693 VPWR.n2758 VGND 1.20645f
C14694 VPWR.n2759 VGND 0.03117f
C14695 VPWR.t422 VGND 0.49153f
C14696 VPWR.t464 VGND 0.18598f
C14697 VPWR.t202 VGND 0.18598f
C14698 VPWR.t282 VGND 0.18598f
C14699 VPWR.t130 VGND 0.18598f
C14700 VPWR.t124 VGND 0.18598f
C14701 VPWR.t132 VGND 0.18598f
C14702 VPWR.t134 VGND 0.16827f
C14703 VPWR.t961 VGND 0.40739f
C14704 VPWR.t876 VGND 0.11292f
C14705 VPWR.n2760 VGND 0.24407f
C14706 VPWR.n2761 VGND 0.13021f
C14707 VPWR.t131 VGND 0.01056f
C14708 VPWR.t125 VGND 0.01056f
C14709 VPWR.n2762 VGND 0.02315f
C14710 VPWR.t944 VGND 0.01056f
C14711 VPWR.t943 VGND 0.01056f
C14712 VPWR.n2763 VGND 0.02315f
C14713 VPWR.n2764 VGND 0.08787f
C14714 VPWR.n2765 VGND 0.07124f
C14715 VPWR.t133 VGND 0.01056f
C14716 VPWR.t135 VGND 0.01056f
C14717 VPWR.n2766 VGND 0.02319f
C14718 VPWR.t946 VGND 0.01056f
C14719 VPWR.t940 VGND 0.01056f
C14720 VPWR.n2767 VGND 0.02319f
C14721 VPWR.n2768 VGND 0.09631f
C14722 VPWR.n2770 VGND 0.27821f
C14723 VPWR.n2771 VGND 0.01314f
C14724 VPWR.n2772 VGND 0.01202f
C14725 VPWR.n2773 VGND 0.01031f
C14726 VPWR.t962 VGND 0.04217f
C14727 VPWR.t1890 VGND 0.04217f
C14728 VPWR.n2775 VGND 0.12454f
C14729 VPWR.n2776 VGND 0.02591f
C14730 VPWR.n2777 VGND 1.20645f
C14731 VPWR.n2778 VGND 0.03117f
C14732 VPWR.t308 VGND 0.49153f
C14733 VPWR.t371 VGND 0.18598f
C14734 VPWR.t279 VGND 0.18598f
C14735 VPWR.t698 VGND 0.18598f
C14736 VPWR.t80 VGND 0.18598f
C14737 VPWR.t90 VGND 0.18598f
C14738 VPWR.t82 VGND 0.18598f
C14739 VPWR.t84 VGND 0.16827f
C14740 VPWR.t926 VGND 0.362f
C14741 VPWR.t878 VGND 0.07971f
C14742 VPWR.t882 VGND 0.0786f
C14743 VPWR.n2779 VGND 0.24297f
C14744 VPWR.n2780 VGND 0.13021f
C14745 VPWR.t81 VGND 0.01056f
C14746 VPWR.t91 VGND 0.01056f
C14747 VPWR.n2781 VGND 0.02315f
C14748 VPWR.t1891 VGND 0.01056f
C14749 VPWR.t1897 VGND 0.01056f
C14750 VPWR.n2782 VGND 0.02315f
C14751 VPWR.n2783 VGND 0.08787f
C14752 VPWR.n2784 VGND 0.07124f
C14753 VPWR.t83 VGND 0.01056f
C14754 VPWR.t85 VGND 0.01056f
C14755 VPWR.n2785 VGND 0.02319f
C14756 VPWR.t1893 VGND 0.01056f
C14757 VPWR.t1895 VGND 0.01056f
C14758 VPWR.n2786 VGND 0.02319f
C14759 VPWR.n2787 VGND 0.09631f
C14760 VPWR.n2789 VGND 0.27821f
C14761 VPWR.n2790 VGND 0.01314f
C14762 VPWR.n2791 VGND 0.01183f
C14763 VPWR.t879 VGND 0.04208f
C14764 VPWR.n2793 VGND 0.04498f
C14765 VPWR.t927 VGND 0.04217f
C14766 VPWR.n2795 VGND 0.06716f
C14767 VPWR.n2796 VGND 0.02591f
C14768 VPWR.n2797 VGND 1.20645f
C14769 VPWR.n2798 VGND 0.03154f
C14770 VPWR.t370 VGND 0.49153f
C14771 VPWR.t197 VGND 0.18598f
C14772 VPWR.t421 VGND 0.18598f
C14773 VPWR.t270 VGND 0.18598f
C14774 VPWR.t1176 VGND 0.18598f
C14775 VPWR.t1110 VGND 0.18598f
C14776 VPWR.t136 VGND 0.18598f
C14777 VPWR.t1166 VGND 0.16827f
C14778 VPWR.t963 VGND 0.38525f
C14779 VPWR.t874 VGND 0.13284f
C14780 VPWR.n2799 VGND 0.24186f
C14781 VPWR.n2800 VGND 0.12828f
C14782 VPWR.t877 VGND 0.04214f
C14783 VPWR.t1177 VGND 0.01056f
C14784 VPWR.t1172 VGND 0.01056f
C14785 VPWR.n2801 VGND 0.02315f
C14786 VPWR.t1888 VGND 0.01056f
C14787 VPWR.t1111 VGND 0.01056f
C14788 VPWR.n2802 VGND 0.02315f
C14789 VPWR.n2803 VGND 0.08787f
C14790 VPWR.n2804 VGND 0.07124f
C14791 VPWR.t1165 VGND 0.01056f
C14792 VPWR.t1167 VGND 0.01056f
C14793 VPWR.n2805 VGND 0.02319f
C14794 VPWR.t137 VGND 0.01056f
C14795 VPWR.t1924 VGND 0.01056f
C14796 VPWR.n2806 VGND 0.02319f
C14797 VPWR.n2807 VGND 0.09631f
C14798 VPWR.n2809 VGND 0.27821f
C14799 VPWR.n2810 VGND 0.01314f
C14800 VPWR.n2811 VGND 0.01164f
C14801 VPWR.t875 VGND 0.04214f
C14802 VPWR.n2812 VGND 0.11101f
C14803 VPWR.t964 VGND 0.04212f
C14804 VPWR.t1889 VGND 0.04212f
C14805 VPWR.n2814 VGND 0.09912f
C14806 VPWR.n2815 VGND 0.02591f
C14807 VPWR.n2816 VGND 1.20645f
C14808 VPWR.n2817 VGND 0.03154f
C14809 VPWR.t925 VGND 0.04212f
C14810 VPWR.n2818 VGND 0.01164f
C14811 VPWR.t881 VGND 0.04214f
C14812 VPWR.n2819 VGND 0.01314f
C14813 VPWR.t427 VGND 0.27876f
C14814 VPWR.t693 VGND 0.10548f
C14815 VPWR.t309 VGND 0.10548f
C14816 VPWR.t1857 VGND 0.10548f
C14817 VPWR.t616 VGND 0.10548f
C14818 VPWR.t1130 VGND 0.10548f
C14819 VPWR.t854 VGND 0.10548f
C14820 VPWR.t175 VGND 0.09543f
C14821 VPWR.t924 VGND 0.21849f
C14822 VPWR.t880 VGND 0.07534f
C14823 VPWR.n2820 VGND 0.1346f
C14824 VPWR.t855 VGND 0.01056f
C14825 VPWR.t176 VGND 0.01056f
C14826 VPWR.n2821 VGND 0.02319f
C14827 VPWR.n2822 VGND 0.05707f
C14828 VPWR.t617 VGND 0.01056f
C14829 VPWR.t1131 VGND 0.01056f
C14830 VPWR.n2823 VGND 0.02413f
C14831 VPWR.n2824 VGND 0.12886f
C14832 VPWR.n2825 VGND 0.27821f
C14833 VPWR.n2827 VGND 0.07122f
C14834 VPWR.n2828 VGND 0.06252f
C14835 VPWR.n2830 VGND 0.05418f
C14836 VPWR.n2831 VGND 0.02591f
C14837 VPWR.n2832 VGND 1.04215f
C14838 VPWR.n2833 VGND 1.2177f
C14839 VPWR.n2834 VGND 0.07719f
C14840 VPWR.t747 VGND 1.35171f
C14841 VPWR.t833 VGND 0.81507f
C14842 VPWR.n2835 VGND 1.02838f
C14843 VPWR.t568 VGND 1.76037f
C14844 VPWR.n2836 VGND 0.07719f
C14845 VPWR.t569 VGND 0.03559f
C14846 VPWR.n2837 VGND 0.22076f
C14847 VPWR.n2838 VGND 0.13668f
C14848 VPWR.n2839 VGND 0.97674f
C14849 VPWR.n2840 VGND 0.13668f
C14850 VPWR.n2841 VGND 0.07719f
C14851 VPWR.t570 VGND 0.03559f
C14852 VPWR.n2842 VGND 0.22076f
C14853 VPWR.n2843 VGND 0.155f
C14854 VPWR.n2844 VGND 0.29302f
C14855 VPWR.n2845 VGND 0.08697f
C14856 VPWR.n2846 VGND 0.16539f
C14857 VPWR.n2847 VGND 0.09048f
C14858 VPWR.n2848 VGND 0.0964f
C14859 VPWR.n2849 VGND 0.13668f
C14860 VPWR.n2850 VGND 0.63993f
C14861 VPWR.n2851 VGND 0.13668f
C14862 VPWR.n2852 VGND 0.0964f
C14863 VPWR.n2853 VGND 0.07971f
C14864 VPWR.n2854 VGND 0.01995f
C14865 VPWR.n2855 VGND 0.01662f
C14866 VPWR.n2856 VGND 0.01648f
C14867 VPWR.n2857 VGND 0.08751f
C14868 VPWR.n2858 VGND 0.26519f
C14869 VPWR.n2859 VGND 0.28412f
C14870 VPWR.n2860 VGND 0.29979f
C14871 VPWR.n2861 VGND 1.87026f
C14872 XThR.Tn[2].t5 VGND 0.01796f
C14873 XThR.Tn[2].t3 VGND 0.01796f
C14874 XThR.Tn[2].n0 VGND 0.03626f
C14875 XThR.Tn[2].t6 VGND 0.01796f
C14876 XThR.Tn[2].t2 VGND 0.01796f
C14877 XThR.Tn[2].n1 VGND 0.04242f
C14878 XThR.Tn[2].n2 VGND 0.12726f
C14879 XThR.Tn[2].t1 VGND 0.01168f
C14880 XThR.Tn[2].t8 VGND 0.01168f
C14881 XThR.Tn[2].n3 VGND 0.02659f
C14882 XThR.Tn[2].t4 VGND 0.01168f
C14883 XThR.Tn[2].t10 VGND 0.01168f
C14884 XThR.Tn[2].n4 VGND 0.02659f
C14885 XThR.Tn[2].t7 VGND 0.01168f
C14886 XThR.Tn[2].t9 VGND 0.01168f
C14887 XThR.Tn[2].n5 VGND 0.0443f
C14888 XThR.Tn[2].t0 VGND 0.01168f
C14889 XThR.Tn[2].t11 VGND 0.01168f
C14890 XThR.Tn[2].n6 VGND 0.02659f
C14891 XThR.Tn[2].n7 VGND 0.12662f
C14892 XThR.Tn[2].n8 VGND 0.07828f
C14893 XThR.Tn[2].n9 VGND 0.08834f
C14894 XThR.Tn[2].t21 VGND 0.01404f
C14895 XThR.Tn[2].t14 VGND 0.01537f
C14896 XThR.Tn[2].n10 VGND 0.03754f
C14897 XThR.Tn[2].n11 VGND 0.07211f
C14898 XThR.Tn[2].t40 VGND 0.01404f
C14899 XThR.Tn[2].t31 VGND 0.01537f
C14900 XThR.Tn[2].n12 VGND 0.03754f
C14901 XThR.Tn[2].t55 VGND 0.01399f
C14902 XThR.Tn[2].t66 VGND 0.01532f
C14903 XThR.Tn[2].n13 VGND 0.03906f
C14904 XThR.Tn[2].n14 VGND 0.02744f
C14905 XThR.Tn[2].n16 VGND 0.08806f
C14906 XThR.Tn[2].t15 VGND 0.01404f
C14907 XThR.Tn[2].t67 VGND 0.01537f
C14908 XThR.Tn[2].n17 VGND 0.03754f
C14909 XThR.Tn[2].t30 VGND 0.01399f
C14910 XThR.Tn[2].t43 VGND 0.01532f
C14911 XThR.Tn[2].n18 VGND 0.03906f
C14912 XThR.Tn[2].n19 VGND 0.02744f
C14913 XThR.Tn[2].n21 VGND 0.08806f
C14914 XThR.Tn[2].t32 VGND 0.01404f
C14915 XThR.Tn[2].t23 VGND 0.01537f
C14916 XThR.Tn[2].n22 VGND 0.03754f
C14917 XThR.Tn[2].t47 VGND 0.01399f
C14918 XThR.Tn[2].t60 VGND 0.01532f
C14919 XThR.Tn[2].n23 VGND 0.03906f
C14920 XThR.Tn[2].n24 VGND 0.02744f
C14921 XThR.Tn[2].n26 VGND 0.08806f
C14922 XThR.Tn[2].t58 VGND 0.01404f
C14923 XThR.Tn[2].t50 VGND 0.01537f
C14924 XThR.Tn[2].n27 VGND 0.03754f
C14925 XThR.Tn[2].t16 VGND 0.01399f
C14926 XThR.Tn[2].t28 VGND 0.01532f
C14927 XThR.Tn[2].n28 VGND 0.03906f
C14928 XThR.Tn[2].n29 VGND 0.02744f
C14929 XThR.Tn[2].n31 VGND 0.08806f
C14930 XThR.Tn[2].t34 VGND 0.01404f
C14931 XThR.Tn[2].t25 VGND 0.01537f
C14932 XThR.Tn[2].n32 VGND 0.03754f
C14933 XThR.Tn[2].t48 VGND 0.01399f
C14934 XThR.Tn[2].t62 VGND 0.01532f
C14935 XThR.Tn[2].n33 VGND 0.03906f
C14936 XThR.Tn[2].n34 VGND 0.02744f
C14937 XThR.Tn[2].n36 VGND 0.08806f
C14938 XThR.Tn[2].t70 VGND 0.01404f
C14939 XThR.Tn[2].t41 VGND 0.01537f
C14940 XThR.Tn[2].n37 VGND 0.03754f
C14941 XThR.Tn[2].t22 VGND 0.01399f
C14942 XThR.Tn[2].t20 VGND 0.01532f
C14943 XThR.Tn[2].n38 VGND 0.03906f
C14944 XThR.Tn[2].n39 VGND 0.02744f
C14945 XThR.Tn[2].n41 VGND 0.08806f
C14946 XThR.Tn[2].t39 VGND 0.01404f
C14947 XThR.Tn[2].t35 VGND 0.01537f
C14948 XThR.Tn[2].n42 VGND 0.03754f
C14949 XThR.Tn[2].t54 VGND 0.01399f
C14950 XThR.Tn[2].t12 VGND 0.01532f
C14951 XThR.Tn[2].n43 VGND 0.03906f
C14952 XThR.Tn[2].n44 VGND 0.02744f
C14953 XThR.Tn[2].n46 VGND 0.08806f
C14954 XThR.Tn[2].t44 VGND 0.01404f
C14955 XThR.Tn[2].t49 VGND 0.01537f
C14956 XThR.Tn[2].n47 VGND 0.03754f
C14957 XThR.Tn[2].t57 VGND 0.01399f
C14958 XThR.Tn[2].t27 VGND 0.01532f
C14959 XThR.Tn[2].n48 VGND 0.03906f
C14960 XThR.Tn[2].n49 VGND 0.02744f
C14961 XThR.Tn[2].n51 VGND 0.08806f
C14962 XThR.Tn[2].t61 VGND 0.01404f
C14963 XThR.Tn[2].t69 VGND 0.01537f
C14964 XThR.Tn[2].n52 VGND 0.03754f
C14965 XThR.Tn[2].t18 VGND 0.01399f
C14966 XThR.Tn[2].t45 VGND 0.01532f
C14967 XThR.Tn[2].n53 VGND 0.03906f
C14968 XThR.Tn[2].n54 VGND 0.02744f
C14969 XThR.Tn[2].n56 VGND 0.08806f
C14970 XThR.Tn[2].t52 VGND 0.01404f
C14971 XThR.Tn[2].t26 VGND 0.01537f
C14972 XThR.Tn[2].n57 VGND 0.03754f
C14973 XThR.Tn[2].t68 VGND 0.01399f
C14974 XThR.Tn[2].t63 VGND 0.01532f
C14975 XThR.Tn[2].n58 VGND 0.03906f
C14976 XThR.Tn[2].n59 VGND 0.02744f
C14977 XThR.Tn[2].n61 VGND 0.08806f
C14978 XThR.Tn[2].t73 VGND 0.01404f
C14979 XThR.Tn[2].t64 VGND 0.01537f
C14980 XThR.Tn[2].n62 VGND 0.03754f
C14981 XThR.Tn[2].t24 VGND 0.01399f
C14982 XThR.Tn[2].t37 VGND 0.01532f
C14983 XThR.Tn[2].n63 VGND 0.03906f
C14984 XThR.Tn[2].n64 VGND 0.02744f
C14985 XThR.Tn[2].n66 VGND 0.08806f
C14986 XThR.Tn[2].t42 VGND 0.01404f
C14987 XThR.Tn[2].t36 VGND 0.01537f
C14988 XThR.Tn[2].n67 VGND 0.03754f
C14989 XThR.Tn[2].t56 VGND 0.01399f
C14990 XThR.Tn[2].t13 VGND 0.01532f
C14991 XThR.Tn[2].n68 VGND 0.03906f
C14992 XThR.Tn[2].n69 VGND 0.02744f
C14993 XThR.Tn[2].n71 VGND 0.08806f
C14994 XThR.Tn[2].t59 VGND 0.01404f
C14995 XThR.Tn[2].t51 VGND 0.01537f
C14996 XThR.Tn[2].n72 VGND 0.03754f
C14997 XThR.Tn[2].t17 VGND 0.01399f
C14998 XThR.Tn[2].t29 VGND 0.01532f
C14999 XThR.Tn[2].n73 VGND 0.03906f
C15000 XThR.Tn[2].n74 VGND 0.02744f
C15001 XThR.Tn[2].n76 VGND 0.08806f
C15002 XThR.Tn[2].t19 VGND 0.01404f
C15003 XThR.Tn[2].t72 VGND 0.01537f
C15004 XThR.Tn[2].n77 VGND 0.03754f
C15005 XThR.Tn[2].t33 VGND 0.01399f
C15006 XThR.Tn[2].t46 VGND 0.01532f
C15007 XThR.Tn[2].n78 VGND 0.03906f
C15008 XThR.Tn[2].n79 VGND 0.02744f
C15009 XThR.Tn[2].n81 VGND 0.08806f
C15010 XThR.Tn[2].t53 VGND 0.01404f
C15011 XThR.Tn[2].t65 VGND 0.01537f
C15012 XThR.Tn[2].n82 VGND 0.03754f
C15013 XThR.Tn[2].t71 VGND 0.01399f
C15014 XThR.Tn[2].t38 VGND 0.01532f
C15015 XThR.Tn[2].n83 VGND 0.03906f
C15016 XThR.Tn[2].n84 VGND 0.02744f
C15017 XThR.Tn[2].n86 VGND 0.08806f
C15018 XThR.Tn[2].n87 VGND 0.08002f
C15019 XThR.Tn[2].n88 VGND 0.17341f
.ends

