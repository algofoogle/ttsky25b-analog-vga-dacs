magic
tech sky130A
magscale 1 2
timestamp 1757957546
<< metal1 >>
rect 10676 38319 10756 38324
rect 6845 38314 10756 38319
rect 6845 38256 10688 38314
rect 10746 38256 10756 38314
rect 6845 38249 10756 38256
rect 6860 37812 6900 38249
rect 10676 38244 10756 38249
rect 7450 38170 10756 38180
rect 7450 38112 10688 38170
rect 10746 38112 10756 38170
rect 7450 38100 10756 38112
rect 7470 37808 7510 38100
rect 10676 38029 10756 38038
rect 9026 38028 10756 38029
rect 9026 37970 10688 38028
rect 10746 37970 10756 38028
rect 9026 37968 10756 37970
rect 9036 37812 9076 37968
rect 10676 37958 10756 37968
rect 10676 37889 10756 37898
rect 9108 37888 10756 37889
rect 9108 37830 10688 37888
rect 10746 37830 10756 37888
rect 9108 37828 10756 37830
rect 9118 37812 9158 37828
rect 10676 37818 10756 37828
rect 18744 30729 18824 30734
rect 18734 30724 18824 30729
rect 18734 30666 18756 30724
rect 18814 30666 18824 30724
rect 18734 30659 18824 30666
rect 18744 30654 18824 30659
rect 18734 30580 18824 30590
rect 18734 30522 18756 30580
rect 18814 30522 18824 30580
rect 18734 30510 18824 30522
rect 18744 29039 18824 29048
rect 18734 29038 18824 29039
rect 18734 28980 18756 29038
rect 18814 28980 18824 29038
rect 18734 28978 18824 28980
rect 18744 28968 18824 28978
rect 18744 28487 18824 28496
rect 18734 28486 18824 28487
rect 18734 28428 18756 28486
rect 18814 28428 18824 28486
rect 18734 28426 18824 28428
rect 18744 28416 18824 28426
rect 10676 25605 10756 25610
rect 6845 25600 10756 25605
rect 6845 25542 10688 25600
rect 10746 25542 10756 25600
rect 6845 25535 10756 25542
rect 6860 25098 6900 25535
rect 10676 25530 10756 25535
rect 7450 25456 10756 25466
rect 7450 25398 10688 25456
rect 10746 25398 10756 25456
rect 7450 25386 10756 25398
rect 7470 25094 7510 25386
rect 10676 25315 10756 25324
rect 9026 25314 10756 25315
rect 9026 25256 10688 25314
rect 10746 25256 10756 25314
rect 9026 25254 10756 25256
rect 9036 25098 9076 25254
rect 10676 25244 10756 25254
rect 10676 25175 10756 25184
rect 9108 25174 10756 25175
rect 9108 25116 10688 25174
rect 10746 25116 10756 25174
rect 9108 25114 10756 25116
rect 9118 25098 9158 25114
rect 10676 25104 10756 25114
rect 18744 18015 18824 18020
rect 18734 18010 18824 18015
rect 18734 17952 18756 18010
rect 18814 17952 18824 18010
rect 18734 17945 18824 17952
rect 18744 17940 18824 17945
rect 18734 17866 18824 17876
rect 18734 17808 18756 17866
rect 18814 17808 18824 17866
rect 18734 17796 18824 17808
rect 18744 16325 18824 16334
rect 18734 16324 18824 16325
rect 18734 16266 18756 16324
rect 18814 16266 18824 16324
rect 18734 16264 18824 16266
rect 18744 16254 18824 16264
rect 18744 15773 18824 15782
rect 18734 15772 18824 15773
rect 18734 15714 18756 15772
rect 18814 15714 18824 15772
rect 18734 15712 18824 15714
rect 18744 15702 18824 15712
rect 10676 12891 10756 12896
rect 6845 12886 10756 12891
rect 6845 12828 10688 12886
rect 10746 12828 10756 12886
rect 6845 12821 10756 12828
rect 6860 12384 6900 12821
rect 10676 12816 10756 12821
rect 7450 12742 10756 12752
rect 7450 12684 10688 12742
rect 10746 12684 10756 12742
rect 7450 12672 10756 12684
rect 7470 12380 7510 12672
rect 10676 12601 10756 12610
rect 9026 12600 10756 12601
rect 9026 12542 10688 12600
rect 10746 12542 10756 12600
rect 9026 12540 10756 12542
rect 9036 12384 9076 12540
rect 10676 12530 10756 12540
rect 10676 12461 10756 12470
rect 9108 12460 10756 12461
rect 9108 12402 10688 12460
rect 10746 12402 10756 12460
rect 9108 12400 10756 12402
rect 9118 12384 9158 12400
rect 10676 12390 10756 12400
rect 18744 5301 18824 5306
rect 18734 5296 18824 5301
rect 18734 5238 18756 5296
rect 18814 5238 18824 5296
rect 18734 5231 18824 5238
rect 18744 5226 18824 5231
rect 18734 5152 18824 5162
rect 18734 5094 18756 5152
rect 18814 5094 18824 5152
rect 18734 5082 18824 5094
rect 18744 3611 18824 3620
rect 18734 3610 18824 3611
rect 18734 3552 18756 3610
rect 18814 3552 18824 3610
rect 18734 3550 18824 3552
rect 18744 3540 18824 3550
rect 18744 3059 18824 3068
rect 18734 3058 18824 3059
rect 18734 3000 18756 3058
rect 18814 3000 18824 3058
rect 18734 2998 18824 3000
rect 18744 2988 18824 2998
<< via1 >>
rect 10688 38256 10746 38314
rect 10688 38112 10746 38170
rect 10688 37970 10746 38028
rect 10688 37830 10746 37888
rect 18756 30666 18814 30724
rect 18756 30522 18814 30580
rect 18756 28980 18814 29038
rect 18756 28428 18814 28486
rect 10688 25542 10746 25600
rect 10688 25398 10746 25456
rect 10688 25256 10746 25314
rect 10688 25116 10746 25174
rect 18756 17952 18814 18010
rect 18756 17808 18814 17866
rect 18756 16266 18814 16324
rect 18756 15714 18814 15772
rect 10688 12828 10746 12886
rect 10688 12684 10746 12742
rect 10688 12542 10746 12600
rect 10688 12402 10746 12460
rect 18756 5238 18814 5296
rect 18756 5094 18814 5152
rect 18756 3552 18814 3610
rect 18756 3000 18814 3058
<< metal2 >>
rect 21028 44902 21112 44912
rect 21028 44800 21038 44902
rect 21102 44800 21112 44902
rect 21028 44790 21112 44800
rect 21580 44902 21664 44912
rect 21580 44800 21590 44902
rect 21654 44800 21664 44902
rect 21580 44790 21664 44800
rect 22132 44902 22216 44912
rect 22132 44800 22142 44902
rect 22206 44800 22216 44902
rect 22132 44790 22216 44800
rect 22684 44902 22768 44912
rect 22684 44800 22694 44902
rect 22758 44800 22768 44902
rect 22684 44790 22768 44800
rect 23236 44902 23320 44912
rect 23236 44800 23246 44902
rect 23310 44800 23320 44902
rect 23236 44790 23320 44800
rect 23788 44902 23872 44912
rect 23788 44800 23798 44902
rect 23862 44800 23872 44902
rect 23788 44790 23872 44800
rect 24340 44902 24424 44912
rect 24340 44800 24350 44902
rect 24414 44800 24424 44902
rect 24340 44790 24424 44800
rect 24892 44902 24976 44912
rect 24892 44800 24902 44902
rect 24966 44800 24976 44902
rect 24892 44790 24976 44800
rect 25444 44902 25528 44912
rect 25444 44800 25454 44902
rect 25518 44800 25528 44902
rect 25444 44790 25528 44800
rect 25996 44902 26080 44912
rect 25996 44800 26006 44902
rect 26070 44800 26080 44902
rect 25996 44790 26080 44800
rect 26548 44902 26632 44912
rect 26548 44800 26558 44902
rect 26622 44800 26632 44902
rect 26548 44790 26632 44800
rect 27100 44902 27184 44912
rect 27100 44800 27110 44902
rect 27174 44800 27184 44902
rect 27100 44790 27184 44800
rect 27652 44902 27736 44912
rect 27652 44800 27662 44902
rect 27726 44800 27736 44902
rect 27652 44790 27736 44800
rect 28204 44902 28288 44912
rect 28204 44800 28214 44902
rect 28278 44800 28288 44902
rect 28204 44790 28288 44800
rect 28756 44902 28840 44912
rect 28756 44800 28766 44902
rect 28830 44800 28840 44902
rect 28756 44790 28840 44800
rect 29308 44902 29392 44912
rect 29308 44800 29318 44902
rect 29382 44800 29392 44902
rect 29308 44790 29392 44800
rect 21038 44758 21102 44790
rect 21590 44758 21654 44790
rect 22142 44758 22206 44790
rect 22694 44758 22758 44790
rect 23246 44758 23310 44790
rect 23798 44758 23862 44790
rect 24350 44758 24414 44790
rect 24902 44758 24966 44790
rect 25454 44758 25518 44790
rect 26006 44758 26070 44790
rect 26558 44758 26622 44790
rect 27110 44758 27174 44790
rect 27662 44758 27726 44790
rect 28214 44758 28278 44790
rect 28766 44758 28830 44790
rect 29318 44758 29382 44790
rect 10676 38314 10756 38324
rect 10676 38256 10688 38314
rect 10746 38256 10756 38314
rect 10676 38244 10756 38256
rect 10676 38170 10756 38180
rect 10676 38112 10688 38170
rect 10746 38112 10756 38170
rect 10676 38100 10756 38112
rect 10676 38028 10756 38038
rect 10676 37970 10688 38028
rect 10746 37970 10756 38028
rect 10676 37958 10756 37970
rect 10676 37888 10756 37898
rect 10676 37830 10688 37888
rect 10746 37830 10756 37888
rect 10676 37818 10756 37830
rect 19072 36972 19148 36982
rect 19072 36966 19082 36972
rect 18748 36920 19082 36966
rect 19072 36916 19082 36920
rect 19138 36916 19148 36972
rect 19072 36906 19148 36916
rect 19072 36698 19148 36708
rect 19072 36694 19082 36698
rect 18748 36648 19082 36694
rect 19072 36642 19082 36648
rect 19138 36642 19148 36698
rect 19072 36632 19148 36642
rect 19072 36426 19148 36436
rect 19072 36422 19082 36426
rect 18748 36376 19082 36422
rect 19072 36370 19082 36376
rect 19138 36370 19148 36426
rect 19072 36360 19148 36370
rect 18744 30724 18824 30734
rect 18744 30666 18756 30724
rect 18814 30666 18824 30724
rect 18744 30654 18824 30666
rect 18744 30580 18824 30590
rect 18744 30522 18756 30580
rect 18814 30522 18824 30580
rect 18744 30510 18824 30522
rect 18744 29038 18824 29048
rect 18744 28980 18756 29038
rect 18814 28980 18824 29038
rect 18744 28968 18824 28980
rect 18744 28486 18824 28496
rect 18744 28428 18756 28486
rect 18814 28428 18824 28486
rect 18744 28416 18824 28428
rect 10676 25600 10756 25610
rect 10676 25542 10688 25600
rect 10746 25542 10756 25600
rect 10676 25530 10756 25542
rect 10676 25456 10756 25466
rect 10676 25398 10688 25456
rect 10746 25398 10756 25456
rect 10676 25386 10756 25398
rect 10676 25314 10756 25324
rect 10676 25256 10688 25314
rect 10746 25256 10756 25314
rect 10676 25244 10756 25256
rect 10676 25174 10756 25184
rect 10676 25116 10688 25174
rect 10746 25116 10756 25174
rect 10676 25104 10756 25116
rect 19072 24258 19148 24268
rect 19072 24252 19082 24258
rect 18748 24206 19082 24252
rect 19072 24202 19082 24206
rect 19138 24202 19148 24258
rect 19072 24192 19148 24202
rect 19072 23984 19148 23994
rect 19072 23980 19082 23984
rect 18748 23934 19082 23980
rect 19072 23928 19082 23934
rect 19138 23928 19148 23984
rect 19072 23918 19148 23928
rect 19072 23712 19148 23722
rect 19072 23708 19082 23712
rect 18748 23662 19082 23708
rect 19072 23656 19082 23662
rect 19138 23656 19148 23712
rect 19072 23646 19148 23656
rect 18744 18010 18824 18020
rect 18744 17952 18756 18010
rect 18814 17952 18824 18010
rect 18744 17940 18824 17952
rect 18744 17866 18824 17876
rect 18744 17808 18756 17866
rect 18814 17808 18824 17866
rect 18744 17796 18824 17808
rect 18744 16324 18824 16334
rect 18744 16266 18756 16324
rect 18814 16266 18824 16324
rect 18744 16254 18824 16266
rect 18744 15772 18824 15782
rect 18744 15714 18756 15772
rect 18814 15714 18824 15772
rect 18744 15702 18824 15714
rect 10676 12886 10756 12896
rect 10676 12828 10688 12886
rect 10746 12828 10756 12886
rect 10676 12816 10756 12828
rect 10676 12742 10756 12752
rect 10676 12684 10688 12742
rect 10746 12684 10756 12742
rect 10676 12672 10756 12684
rect 10676 12600 10756 12610
rect 10676 12542 10688 12600
rect 10746 12542 10756 12600
rect 10676 12530 10756 12542
rect 10676 12460 10756 12470
rect 10676 12402 10688 12460
rect 10746 12402 10756 12460
rect 10676 12390 10756 12402
rect 19072 11544 19148 11554
rect 19072 11538 19082 11544
rect 18748 11492 19082 11538
rect 19072 11488 19082 11492
rect 19138 11488 19148 11544
rect 19072 11478 19148 11488
rect 19072 11270 19148 11280
rect 19072 11266 19082 11270
rect 18748 11220 19082 11266
rect 19072 11214 19082 11220
rect 19138 11214 19148 11270
rect 19072 11204 19148 11214
rect 19072 10998 19148 11008
rect 19072 10994 19082 10998
rect 18748 10948 19082 10994
rect 19072 10942 19082 10948
rect 19138 10942 19148 10998
rect 19072 10932 19148 10942
rect 18744 5296 18824 5306
rect 18744 5238 18756 5296
rect 18814 5238 18824 5296
rect 18744 5226 18824 5238
rect 18744 5152 18824 5162
rect 18744 5094 18756 5152
rect 18814 5094 18824 5152
rect 18744 5082 18824 5094
rect 18744 3610 18824 3620
rect 18744 3552 18756 3610
rect 18814 3552 18824 3610
rect 18744 3540 18824 3552
rect 18744 3058 18824 3068
rect 18744 3000 18756 3058
rect 18814 3000 18824 3058
rect 18744 2988 18824 3000
<< via2 >>
rect 21038 44800 21102 44902
rect 21590 44800 21654 44902
rect 22142 44800 22206 44902
rect 22694 44800 22758 44902
rect 23246 44800 23310 44902
rect 23798 44800 23862 44902
rect 24350 44800 24414 44902
rect 24902 44800 24966 44902
rect 25454 44800 25518 44902
rect 26006 44800 26070 44902
rect 26558 44800 26622 44902
rect 27110 44800 27174 44902
rect 27662 44800 27726 44902
rect 28214 44800 28278 44902
rect 28766 44800 28830 44902
rect 29318 44800 29382 44902
rect 10688 38256 10746 38314
rect 10688 38112 10746 38170
rect 10688 37970 10746 38028
rect 10688 37830 10746 37888
rect 19082 36916 19138 36972
rect 19082 36642 19138 36698
rect 19082 36370 19138 36426
rect 18756 30666 18814 30724
rect 18756 30522 18814 30580
rect 18756 28980 18814 29038
rect 18756 28428 18814 28486
rect 10688 25542 10746 25600
rect 10688 25398 10746 25456
rect 10688 25256 10746 25314
rect 10688 25116 10746 25174
rect 19082 24202 19138 24258
rect 19082 23928 19138 23984
rect 19082 23656 19138 23712
rect 18756 17952 18814 18010
rect 18756 17808 18814 17866
rect 18756 16266 18814 16324
rect 18756 15714 18814 15772
rect 10688 12828 10746 12886
rect 10688 12684 10746 12742
rect 10688 12542 10746 12600
rect 10688 12402 10746 12460
rect 19082 11488 19138 11544
rect 19082 11214 19138 11270
rect 19082 10942 19138 10998
rect 18756 5238 18814 5296
rect 18756 5094 18814 5152
rect 18756 3552 18814 3610
rect 18756 3000 18814 3058
<< metal3 >>
rect 9722 44846 9728 44910
rect 9792 44846 9798 44910
rect 21028 44906 21112 44912
rect 740 43980 746 44044
rect 810 44042 816 44044
rect 9730 44042 9790 44846
rect 21028 44796 21034 44906
rect 21106 44796 21112 44906
rect 21028 44790 21112 44796
rect 21580 44906 21664 44912
rect 21580 44796 21586 44906
rect 21658 44796 21664 44906
rect 21580 44790 21664 44796
rect 22132 44906 22216 44912
rect 22132 44796 22138 44906
rect 22210 44796 22216 44906
rect 22132 44790 22216 44796
rect 22684 44906 22768 44912
rect 22684 44796 22690 44906
rect 22762 44796 22768 44906
rect 22684 44790 22768 44796
rect 23236 44906 23320 44912
rect 23236 44796 23242 44906
rect 23314 44796 23320 44906
rect 23236 44790 23320 44796
rect 23788 44906 23872 44912
rect 23788 44796 23794 44906
rect 23866 44796 23872 44906
rect 23788 44790 23872 44796
rect 24340 44906 24424 44912
rect 24340 44796 24346 44906
rect 24418 44796 24424 44906
rect 24340 44790 24424 44796
rect 24892 44906 24976 44912
rect 24892 44796 24898 44906
rect 24970 44796 24976 44906
rect 24892 44790 24976 44796
rect 25444 44906 25528 44912
rect 25444 44796 25450 44906
rect 25522 44796 25528 44906
rect 25444 44790 25528 44796
rect 25996 44906 26080 44912
rect 25996 44796 26002 44906
rect 26074 44796 26080 44906
rect 25996 44790 26080 44796
rect 26548 44906 26632 44912
rect 26548 44796 26554 44906
rect 26626 44796 26632 44906
rect 26548 44790 26632 44796
rect 27100 44906 27184 44912
rect 27100 44796 27106 44906
rect 27178 44796 27184 44906
rect 27100 44790 27184 44796
rect 27652 44906 27736 44912
rect 27652 44796 27658 44906
rect 27730 44796 27736 44906
rect 27652 44790 27736 44796
rect 28204 44906 28288 44912
rect 28204 44796 28210 44906
rect 28282 44796 28288 44906
rect 28204 44790 28288 44796
rect 28756 44906 28840 44912
rect 28756 44796 28762 44906
rect 28834 44796 28840 44906
rect 28756 44790 28840 44796
rect 29308 44906 29392 44912
rect 29308 44796 29314 44906
rect 29386 44796 29392 44906
rect 29308 44790 29392 44796
rect 810 43982 9790 44042
rect 810 43980 816 43982
rect 13798 42640 20540 42644
rect 13798 42528 18794 42640
rect 18926 42528 20540 42640
rect 13798 42524 20540 42528
rect 13798 42368 20540 42372
rect 13798 42256 18242 42368
rect 18374 42256 20540 42368
rect 13798 42252 20540 42256
rect 13798 42096 20540 42100
rect 13798 41984 17690 42096
rect 17822 41984 20540 42096
rect 13798 41980 20540 41984
rect 13798 41824 20540 41828
rect 13798 41712 17138 41824
rect 17270 41712 20540 41824
rect 13798 41708 20540 41712
rect 13798 41552 20540 41556
rect 13798 41440 16586 41552
rect 16718 41440 20540 41552
rect 13798 41436 20540 41440
rect 13798 41280 20540 41284
rect 13798 41168 16034 41280
rect 16166 41168 20540 41280
rect 13798 41164 20540 41168
rect 13798 41008 20540 41012
rect 13798 40896 15482 41008
rect 15614 40896 20540 41008
rect 13798 40892 20540 40896
rect 13798 40736 20540 40740
rect 13798 40624 14930 40736
rect 15062 40624 20540 40736
rect 13798 40620 20540 40624
rect 13798 40464 20540 40468
rect 13798 40352 14378 40464
rect 14510 40352 20540 40464
rect 13798 40348 20540 40352
rect 13798 40192 20540 40196
rect 13798 40080 13826 40192
rect 13958 40080 20540 40192
rect 13798 40076 20540 40080
rect 10676 38316 10756 38324
rect 10676 38314 20549 38316
rect 10676 38256 10688 38314
rect 10746 38256 20549 38314
rect 10676 38254 20549 38256
rect 10676 38244 10756 38254
rect 10676 38172 10756 38180
rect 10676 38170 20379 38172
rect 10676 38112 10688 38170
rect 10746 38112 20379 38170
rect 10676 38110 20379 38112
rect 10676 38100 10756 38110
rect 10676 38030 10756 38038
rect 10676 38028 20209 38030
rect 10676 37970 10688 38028
rect 10746 37970 20209 38028
rect 10676 37968 20209 37970
rect 10676 37958 10756 37968
rect 10676 37890 10756 37898
rect 10676 37888 19956 37890
rect 10676 37830 10688 37888
rect 10746 37830 19956 37888
rect 10676 37828 19956 37830
rect 10676 37818 10756 37828
rect 200 37744 2380 37754
rect 200 36940 210 37744
rect 910 36940 2380 37744
rect 19894 37179 19956 37828
rect 20147 37453 20209 37968
rect 20317 37737 20379 38110
rect 20487 37933 20549 38254
rect 20317 37675 20547 37737
rect 20147 37391 20531 37453
rect 19894 37117 20551 37179
rect 19072 36980 19148 36982
rect 19072 36972 20344 36980
rect 19072 36916 19082 36972
rect 19138 36916 20344 36972
rect 19072 36908 20344 36916
rect 19072 36906 19148 36908
rect 19072 36706 19148 36708
rect 19072 36698 20154 36706
rect 19072 36642 19082 36698
rect 19138 36642 20154 36698
rect 19072 36634 20154 36642
rect 19072 36632 19148 36634
rect 19072 36434 19148 36436
rect 19072 36426 19934 36434
rect 19072 36370 19082 36426
rect 19138 36370 19934 36426
rect 19072 36362 19934 36370
rect 19072 36360 19148 36362
rect 200 34946 210 35960
rect 910 34946 2380 35960
rect 19023 35652 19201 35657
rect 17672 35472 17678 35652
rect 17856 35651 19202 35652
rect 17856 35473 19023 35651
rect 19201 35473 19202 35651
rect 17856 35472 19202 35473
rect 19023 35467 19201 35472
rect 19862 35272 19934 36362
rect 20082 35542 20154 36634
rect 20272 35812 20344 36908
rect 20272 35740 20556 35812
rect 20082 35470 20532 35542
rect 19862 35200 20538 35272
rect 200 34936 2380 34946
rect 18744 30726 18824 30734
rect 18744 30724 20541 30726
rect 18744 30666 18756 30724
rect 18814 30666 20541 30724
rect 18744 30664 20541 30666
rect 18744 30654 18824 30664
rect 18744 30582 18824 30590
rect 18744 30580 20389 30582
rect 18744 30522 18756 30580
rect 18814 30522 20389 30580
rect 18744 30520 20389 30522
rect 18744 30510 18824 30520
rect 20327 29551 20389 30520
rect 20479 29765 20541 30664
rect 20327 29489 20513 29551
rect 20123 29213 20521 29275
rect 18744 29040 18824 29048
rect 20123 29040 20185 29213
rect 18744 29038 20185 29040
rect 18744 28980 18756 29038
rect 18814 28980 20185 29038
rect 18744 28978 20185 28980
rect 18744 28968 18824 28978
rect 20327 28951 20537 29013
rect 18744 28488 18824 28496
rect 20327 28488 20389 28951
rect 18744 28486 20389 28488
rect 18744 28428 18756 28486
rect 18814 28428 20389 28486
rect 18744 28426 20389 28428
rect 18744 28416 18824 28426
rect 19829 26722 20007 26727
rect 17594 26542 17600 26722
rect 17778 26721 20008 26722
rect 17778 26543 19829 26721
rect 20007 26543 20008 26721
rect 17778 26542 20008 26543
rect 19829 26537 20007 26542
rect 10676 25602 10756 25610
rect 10676 25600 20545 25602
rect 10676 25542 10688 25600
rect 10746 25542 20545 25600
rect 10676 25540 20545 25542
rect 10676 25530 10756 25540
rect 10676 25458 10756 25466
rect 10676 25456 20377 25458
rect 10676 25398 10688 25456
rect 10746 25398 20377 25456
rect 10676 25396 20377 25398
rect 10676 25386 10756 25396
rect 10676 25316 10756 25324
rect 10676 25314 20219 25316
rect 10676 25256 10688 25314
rect 10746 25256 20219 25314
rect 10676 25254 20219 25256
rect 10676 25244 10756 25254
rect 10676 25176 10756 25184
rect 10676 25174 20049 25176
rect 10676 25116 10688 25174
rect 10746 25116 20049 25174
rect 10676 25114 20049 25116
rect 10676 25104 10756 25114
rect 200 25030 2380 25040
rect 200 24120 210 25030
rect 910 24120 2380 25030
rect 19987 24461 20049 25114
rect 20157 24655 20219 25254
rect 20315 24927 20377 25396
rect 20483 25149 20545 25540
rect 20315 24865 20547 24927
rect 20157 24593 20539 24655
rect 19987 24399 20247 24461
rect 20185 24387 20247 24399
rect 20185 24325 20559 24387
rect 19072 24266 19148 24268
rect 19072 24258 20056 24266
rect 19072 24202 19082 24258
rect 19138 24202 20056 24258
rect 19072 24194 20056 24202
rect 19072 24192 19148 24194
rect 19984 24120 20056 24194
rect 19984 24048 20542 24120
rect 19072 23992 19148 23994
rect 19072 23984 19870 23992
rect 19072 23928 19082 23984
rect 19138 23928 19870 23984
rect 19072 23920 19870 23928
rect 19072 23918 19148 23920
rect 19798 23850 19870 23920
rect 19798 23778 20550 23850
rect 19072 23720 19148 23722
rect 19072 23712 19644 23720
rect 19072 23656 19082 23712
rect 19138 23656 19644 23712
rect 19072 23648 19644 23656
rect 19072 23646 19148 23648
rect 19572 23582 19644 23648
rect 19572 23510 20526 23582
rect 200 22232 210 23140
rect 910 22232 2380 23140
rect 200 22222 2380 22232
rect 20241 18071 20561 18133
rect 18744 18012 18824 18020
rect 20241 18012 20303 18071
rect 18744 18010 20303 18012
rect 18744 17952 18756 18010
rect 18814 17952 20303 18010
rect 18744 17950 20303 17952
rect 18744 17940 18824 17950
rect 18744 17868 18824 17876
rect 18744 17866 20531 17868
rect 18744 17808 18756 17866
rect 18814 17808 20531 17866
rect 18744 17806 20531 17808
rect 18744 17796 18824 17806
rect 20331 17519 20541 17581
rect 18744 16326 18824 16334
rect 20331 16326 20393 17519
rect 18744 16324 20393 16326
rect 18744 16266 18756 16324
rect 18814 16266 20393 16324
rect 18744 16264 20393 16266
rect 18744 16254 18824 16264
rect 18744 15774 18824 15782
rect 20493 15774 20555 17317
rect 18744 15772 20555 15774
rect 18744 15714 18756 15772
rect 18814 15714 20555 15772
rect 18744 15712 20555 15714
rect 18744 15702 18824 15712
rect 19570 13998 19950 14010
rect 17860 13818 17866 13998
rect 18044 13997 19950 13998
rect 18044 13819 19577 13997
rect 19755 13819 19950 13997
rect 18044 13818 19950 13819
rect 19570 13810 19950 13818
rect 18514 13447 20533 13509
rect 10676 12888 10756 12896
rect 18514 12888 18576 13447
rect 10676 12886 18576 12888
rect 10676 12828 10688 12886
rect 10746 12828 18576 12886
rect 10676 12826 18576 12828
rect 18657 13175 20555 13237
rect 10676 12816 10756 12826
rect 10676 12744 10756 12752
rect 18657 12744 18719 13175
rect 10676 12742 18719 12744
rect 10676 12684 10688 12742
rect 10746 12684 18719 12742
rect 10676 12682 18719 12684
rect 18801 12905 20535 12967
rect 10676 12672 10756 12682
rect 10676 12602 10756 12610
rect 18801 12602 18863 12905
rect 10676 12600 18863 12602
rect 10676 12542 10688 12600
rect 10746 12542 18863 12600
rect 10676 12540 18863 12542
rect 18971 12631 20539 12693
rect 10676 12530 10756 12540
rect 10676 12462 10756 12470
rect 18971 12462 19033 12631
rect 10676 12460 19033 12462
rect 10676 12402 10688 12460
rect 10746 12402 19033 12460
rect 10676 12400 19033 12402
rect 10676 12390 10756 12400
rect 20034 12356 20534 12428
rect 200 12316 2380 12326
rect 200 11380 210 12316
rect 910 11380 2380 12316
rect 19072 11552 19148 11554
rect 20034 11552 20106 12356
rect 19072 11544 20106 11552
rect 19072 11488 19082 11544
rect 19138 11488 20106 11544
rect 19072 11480 20106 11488
rect 20282 12078 20550 12150
rect 19072 11478 19148 11480
rect 19072 11278 19148 11280
rect 20282 11278 20354 12078
rect 19072 11270 20354 11278
rect 19072 11214 19082 11270
rect 19138 11214 20354 11270
rect 19072 11206 20354 11214
rect 19072 11204 19148 11206
rect 19072 11006 19148 11008
rect 20502 11006 20574 11878
rect 19072 10998 20574 11006
rect 19072 10942 19082 10998
rect 19138 10942 20574 10998
rect 19072 10934 20574 10942
rect 19072 10932 19148 10934
rect 200 9518 210 10400
rect 910 9518 2380 10400
rect 200 9508 2380 9518
rect 19785 6373 20557 6435
rect 18744 5298 18824 5306
rect 19785 5298 19847 6373
rect 18744 5296 19847 5298
rect 18744 5238 18756 5296
rect 18814 5238 19847 5296
rect 18744 5236 19847 5238
rect 19951 6101 20547 6163
rect 18744 5226 18824 5236
rect 18744 5154 18824 5162
rect 19951 5154 20013 6101
rect 18744 5152 20013 5154
rect 18744 5094 18756 5152
rect 18814 5094 20013 5152
rect 18744 5092 20013 5094
rect 20133 5833 20547 5895
rect 18744 5082 18824 5092
rect 18744 3612 18824 3620
rect 20133 3612 20195 5833
rect 18744 3610 20195 3612
rect 18744 3552 18756 3610
rect 18814 3552 20195 3610
rect 18744 3550 20195 3552
rect 20329 5561 20551 5623
rect 18744 3540 18824 3550
rect 18744 3060 18824 3068
rect 20329 3060 20391 5561
rect 18744 3058 20391 3060
rect 18744 3000 18756 3058
rect 18814 3000 20391 3058
rect 18744 2998 20391 3000
rect 18744 2988 18824 2998
rect 19022 2786 19202 2792
rect 19022 830 19202 2608
rect 18770 829 19202 830
rect 18765 651 18771 829
rect 18949 651 19202 829
rect 18770 650 19202 651
<< via3 >>
rect 9728 44846 9792 44910
rect 746 43980 810 44044
rect 21034 44902 21106 44906
rect 21034 44800 21038 44902
rect 21038 44800 21102 44902
rect 21102 44800 21106 44902
rect 21034 44796 21106 44800
rect 21586 44902 21658 44906
rect 21586 44800 21590 44902
rect 21590 44800 21654 44902
rect 21654 44800 21658 44902
rect 21586 44796 21658 44800
rect 22138 44902 22210 44906
rect 22138 44800 22142 44902
rect 22142 44800 22206 44902
rect 22206 44800 22210 44902
rect 22138 44796 22210 44800
rect 22690 44902 22762 44906
rect 22690 44800 22694 44902
rect 22694 44800 22758 44902
rect 22758 44800 22762 44902
rect 22690 44796 22762 44800
rect 23242 44902 23314 44906
rect 23242 44800 23246 44902
rect 23246 44800 23310 44902
rect 23310 44800 23314 44902
rect 23242 44796 23314 44800
rect 23794 44902 23866 44906
rect 23794 44800 23798 44902
rect 23798 44800 23862 44902
rect 23862 44800 23866 44902
rect 23794 44796 23866 44800
rect 24346 44902 24418 44906
rect 24346 44800 24350 44902
rect 24350 44800 24414 44902
rect 24414 44800 24418 44902
rect 24346 44796 24418 44800
rect 24898 44902 24970 44906
rect 24898 44800 24902 44902
rect 24902 44800 24966 44902
rect 24966 44800 24970 44902
rect 24898 44796 24970 44800
rect 25450 44902 25522 44906
rect 25450 44800 25454 44902
rect 25454 44800 25518 44902
rect 25518 44800 25522 44902
rect 25450 44796 25522 44800
rect 26002 44902 26074 44906
rect 26002 44800 26006 44902
rect 26006 44800 26070 44902
rect 26070 44800 26074 44902
rect 26002 44796 26074 44800
rect 26554 44902 26626 44906
rect 26554 44800 26558 44902
rect 26558 44800 26622 44902
rect 26622 44800 26626 44902
rect 26554 44796 26626 44800
rect 27106 44902 27178 44906
rect 27106 44800 27110 44902
rect 27110 44800 27174 44902
rect 27174 44800 27178 44902
rect 27106 44796 27178 44800
rect 27658 44902 27730 44906
rect 27658 44800 27662 44902
rect 27662 44800 27726 44902
rect 27726 44800 27730 44902
rect 27658 44796 27730 44800
rect 28210 44902 28282 44906
rect 28210 44800 28214 44902
rect 28214 44800 28278 44902
rect 28278 44800 28282 44902
rect 28210 44796 28282 44800
rect 28762 44902 28834 44906
rect 28762 44800 28766 44902
rect 28766 44800 28830 44902
rect 28830 44800 28834 44902
rect 28762 44796 28834 44800
rect 29314 44902 29386 44906
rect 29314 44800 29318 44902
rect 29318 44800 29382 44902
rect 29382 44800 29386 44902
rect 29314 44796 29386 44800
rect 18794 42528 18926 42640
rect 18242 42256 18374 42368
rect 17690 41984 17822 42096
rect 17138 41712 17270 41824
rect 16586 41440 16718 41552
rect 16034 41168 16166 41280
rect 15482 40896 15614 41008
rect 14930 40624 15062 40736
rect 14378 40352 14510 40464
rect 13826 40080 13958 40192
rect 210 36940 910 37744
rect 210 34946 910 35960
rect 17678 35472 17856 35652
rect 19023 35473 19201 35651
rect 17600 26542 17778 26722
rect 19829 26543 20007 26721
rect 210 24120 910 25030
rect 210 22232 910 23140
rect 17866 13818 18044 13998
rect 19577 13819 19755 13997
rect 210 11380 910 12316
rect 210 9518 910 10400
rect 19022 2608 19202 2786
rect 18771 651 18949 829
<< metal4 >>
rect 6134 44804 6194 45152
rect 6686 44804 6746 45152
rect 7238 44804 7298 45152
rect 7790 44804 7850 45152
rect 8342 44804 8402 45152
rect 8894 44804 8954 45152
rect 9446 44908 9506 45152
rect 9727 44910 9793 44911
rect 9727 44908 9728 44910
rect 9446 44848 9728 44908
rect 9727 44846 9728 44848
rect 9792 44908 9793 44910
rect 9998 44908 10058 45152
rect 9792 44848 10058 44908
rect 9792 44846 9793 44848
rect 9727 44845 9793 44846
rect 10550 44804 10610 45152
rect 11102 44804 11162 45152
rect 11654 44804 11714 45152
rect 12206 44804 12266 45152
rect 12758 44804 12818 45152
rect 13310 44804 13370 45152
rect 13862 44858 13922 45152
rect 14414 44858 14474 45152
rect 14966 44858 15026 45152
rect 15518 44858 15578 45152
rect 16070 44858 16130 45152
rect 16622 44858 16682 45152
rect 17174 44858 17234 45152
rect 17726 44858 17786 45152
rect 18278 44858 18338 45152
rect 18830 44858 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44912 21098 45152
rect 21590 44912 21650 45152
rect 22142 44912 22202 45152
rect 22694 44912 22754 45152
rect 23246 44912 23306 45152
rect 23798 44912 23858 45152
rect 24350 44912 24410 45152
rect 24902 44912 24962 45152
rect 25454 44912 25514 45152
rect 26006 44912 26066 45152
rect 26558 44912 26618 45152
rect 27110 44912 27170 45152
rect 27662 44912 27722 45152
rect 28214 44912 28274 45152
rect 28766 44912 28826 45152
rect 29318 44912 29378 45152
rect 21028 44906 21112 44912
rect 1120 44704 9360 44804
rect 10144 44704 13440 44804
rect 1120 44556 13440 44704
rect 200 44044 920 44152
rect 200 43980 746 44044
rect 810 43980 920 44044
rect 200 37744 920 43980
rect 200 36940 210 37744
rect 910 36940 920 37744
rect 200 35960 920 36940
rect 200 34946 210 35960
rect 910 34946 920 35960
rect 200 25030 920 34946
rect 200 24120 210 25030
rect 910 24120 920 25030
rect 200 23140 920 24120
rect 200 22232 210 23140
rect 910 22232 920 23140
rect 200 12316 920 22232
rect 200 11380 210 12316
rect 910 11380 920 12316
rect 200 10400 920 11380
rect 200 9518 210 10400
rect 910 9518 920 10400
rect 200 1000 920 9518
rect 1120 1000 1840 44556
rect 13822 40192 13962 44858
rect 13822 40080 13826 40192
rect 13958 40080 13962 40192
rect 13822 40028 13962 40080
rect 14374 40464 14514 44858
rect 14374 40352 14378 40464
rect 14510 40352 14514 40464
rect 14374 40028 14514 40352
rect 14926 40736 15066 44858
rect 14926 40624 14930 40736
rect 15062 40624 15066 40736
rect 14926 40028 15066 40624
rect 15478 41008 15618 44858
rect 15478 40896 15482 41008
rect 15614 40896 15618 41008
rect 15478 40028 15618 40896
rect 16030 41280 16170 44858
rect 16030 41168 16034 41280
rect 16166 41168 16170 41280
rect 16030 40028 16170 41168
rect 16582 41552 16722 44858
rect 16582 41440 16586 41552
rect 16718 41440 16722 41552
rect 16582 40028 16722 41440
rect 17134 41824 17274 44858
rect 17134 41712 17138 41824
rect 17270 41712 17274 41824
rect 17134 40028 17274 41712
rect 17686 42096 17826 44858
rect 17686 41984 17690 42096
rect 17822 41984 17826 42096
rect 17686 40028 17826 41984
rect 18238 42368 18378 44858
rect 18238 42256 18242 42368
rect 18374 42256 18378 42368
rect 18238 40028 18378 42256
rect 18790 42640 18930 44858
rect 21028 44796 21034 44906
rect 21106 44796 21112 44906
rect 21028 44790 21112 44796
rect 21580 44906 21664 44912
rect 21580 44796 21586 44906
rect 21658 44796 21664 44906
rect 21580 44790 21664 44796
rect 22132 44906 22216 44912
rect 22132 44796 22138 44906
rect 22210 44796 22216 44906
rect 22132 44790 22216 44796
rect 22684 44906 22768 44912
rect 22684 44796 22690 44906
rect 22762 44796 22768 44906
rect 22684 44790 22768 44796
rect 23236 44906 23320 44912
rect 23236 44796 23242 44906
rect 23314 44796 23320 44906
rect 23236 44790 23320 44796
rect 23788 44906 23872 44912
rect 23788 44796 23794 44906
rect 23866 44796 23872 44906
rect 23788 44790 23872 44796
rect 24340 44906 24424 44912
rect 24340 44796 24346 44906
rect 24418 44796 24424 44906
rect 24340 44790 24424 44796
rect 24892 44906 24976 44912
rect 24892 44796 24898 44906
rect 24970 44796 24976 44906
rect 24892 44790 24976 44796
rect 25444 44906 25528 44912
rect 25444 44796 25450 44906
rect 25522 44796 25528 44906
rect 25444 44790 25528 44796
rect 25996 44906 26080 44912
rect 25996 44796 26002 44906
rect 26074 44796 26080 44906
rect 25996 44790 26080 44796
rect 26548 44906 26632 44912
rect 26548 44796 26554 44906
rect 26626 44796 26632 44906
rect 26548 44790 26632 44796
rect 27100 44906 27184 44912
rect 27100 44796 27106 44906
rect 27178 44796 27184 44906
rect 27100 44790 27184 44796
rect 27652 44906 27736 44912
rect 27652 44796 27658 44906
rect 27730 44796 27736 44906
rect 27652 44790 27736 44796
rect 28204 44906 28288 44912
rect 28204 44796 28210 44906
rect 28282 44796 28288 44906
rect 28204 44790 28288 44796
rect 28756 44906 28840 44912
rect 28756 44796 28762 44906
rect 28834 44796 28840 44906
rect 28756 44790 28840 44796
rect 29308 44906 29392 44912
rect 29308 44796 29314 44906
rect 29386 44796 29392 44906
rect 29308 44790 29392 44796
rect 18790 42528 18794 42640
rect 18926 42528 18930 42640
rect 18790 40028 18930 42528
rect 17677 35652 17857 35653
rect 15663 35613 17569 35626
rect 17677 35613 17678 35652
rect 15663 35536 17678 35613
rect 17513 35511 17678 35536
rect 17677 35472 17678 35511
rect 17856 35472 17857 35652
rect 17677 35471 17857 35472
rect 19022 35651 19202 35652
rect 19022 35473 19023 35651
rect 19201 35473 19202 35651
rect 17599 26722 17779 26723
rect 15482 26542 17600 26722
rect 17778 26542 17779 26722
rect 17599 26541 17779 26542
rect 17865 13998 18045 13999
rect 15482 13818 17866 13998
rect 18044 13818 18045 13998
rect 17865 13817 18045 13818
rect 19022 2787 19202 35473
rect 19828 26721 20308 26722
rect 19828 26543 19829 26721
rect 20007 26543 20308 26721
rect 19828 26542 20308 26543
rect 19570 13998 19950 14010
rect 19570 13997 19956 13998
rect 19570 13819 19577 13997
rect 19755 13819 19956 13997
rect 19570 13810 19956 13819
rect 19021 2786 19203 2787
rect 19021 2608 19022 2786
rect 19202 2608 19203 2786
rect 19021 2607 19203 2608
rect 15486 1112 19556 1292
rect 18770 829 18950 830
rect 18770 651 18771 829
rect 18949 651 18950 829
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 651
rect 19376 674 19556 1112
rect 19776 996 19956 13810
rect 20128 1308 20308 26542
rect 20128 1128 23796 1308
rect 19776 816 23484 996
rect 19376 494 22814 674
rect 22634 0 22814 494
rect 23304 610 23484 816
rect 23616 894 23796 1128
rect 24124 1000 24444 44200
rect 24784 1000 25104 44200
rect 30524 1000 30844 44200
rect 31184 1000 31504 44200
rect 23616 714 30542 894
rect 23304 430 26678 610
rect 26498 0 26678 430
rect 30362 0 30542 714
use controller_wrapper  controller_wrapper_0
timestamp 1757954071
transform 1 0 20468 0 1 900
box 0 496 11394 43900
use csdac255  dac_blue
timestamp 1757954071
transform -1 0 16648 0 1 1000
box -2130 0 14828 11424
use csdac255  dac_green
timestamp 1757954071
transform -1 0 16648 0 1 13714
box -2130 0 14828 11424
use csdac255  dac_red
timestamp 1757954071
transform -1 0 16648 0 1 26428
box -2130 0 14828 11424
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 920 44152 0 FreeSans 3200 90 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 1120 1000 1840 44152 0 FreeSans 3200 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 24124 1000 24444 44200 0 FreeSans 1600 90 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 24784 1000 25104 44200 0 FreeSans 1600 90 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 30524 1000 30844 44200 0 FreeSans 1600 90 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 31184 1000 31504 44200 0 FreeSans 1600 90 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
